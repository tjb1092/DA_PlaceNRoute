magic
tech scmos
timestamp 1555018311 
<< pdiffusion >>
rect 1 -26 7 -20
rect 8 -26 14 -20
rect 15 -26 21 -20
rect 22 -26 28 -20
rect 29 -26 35 -20
rect 36 -26 42 -20
rect 43 -26 49 -20
rect 50 -26 56 -20
rect 211 -26 217 -20
rect 253 -26 256 -20
rect 351 -26 354 -20
rect 393 -26 399 -20
rect 414 -26 420 -20
rect 421 -26 424 -20
rect 428 -26 434 -20
rect 442 -26 448 -20
rect 484 -26 487 -20
rect 547 -26 550 -20
rect 554 -26 560 -20
rect 568 -26 574 -20
rect 575 -26 578 -20
rect 582 -26 585 -20
rect 603 -26 606 -20
rect 610 -26 616 -20
rect 617 -26 620 -20
rect 624 -26 627 -20
rect 631 -26 637 -20
rect 638 -26 641 -20
rect 645 -26 648 -20
rect 652 -26 658 -20
rect 659 -26 665 -20
rect 680 -26 686 -20
rect 687 -26 690 -20
rect 701 -26 707 -20
rect 708 -26 711 -20
rect 715 -26 718 -20
rect 729 -26 732 -20
rect 764 -26 770 -20
rect 771 -26 774 -20
rect 792 -26 798 -20
rect 799 -26 805 -20
rect 806 -26 812 -20
rect 813 -26 816 -20
rect 820 -26 826 -20
rect 827 -26 830 -20
rect 834 -26 837 -20
rect 841 -26 847 -20
rect 848 -26 854 -20
rect 855 -26 861 -20
rect 862 -26 868 -20
rect 869 -26 872 -20
rect 883 -26 889 -20
rect 890 -26 893 -20
rect 897 -26 903 -20
rect 911 -26 917 -20
rect 918 -26 921 -20
rect 960 -26 963 -20
rect 967 -26 973 -20
rect 974 -26 980 -20
rect 981 -26 984 -20
rect 988 -26 991 -20
rect 1037 -26 1040 -20
rect 1072 -26 1075 -20
rect 1086 -26 1089 -20
rect 1093 -26 1096 -20
rect 1121 -26 1127 -20
rect 1128 -26 1134 -20
rect 1205 -26 1208 -20
rect 1436 -26 1442 -20
rect 1625 -26 1631 -20
rect 1 -73 7 -67
rect 8 -73 14 -67
rect 15 -73 21 -67
rect 22 -73 28 -67
rect 29 -73 35 -67
rect 36 -73 42 -67
rect 43 -73 49 -67
rect 50 -73 56 -67
rect 57 -73 63 -67
rect 183 -73 186 -67
rect 197 -73 200 -67
rect 239 -73 242 -67
rect 274 -73 277 -67
rect 295 -73 298 -67
rect 309 -73 315 -67
rect 316 -73 319 -67
rect 351 -73 357 -67
rect 393 -73 396 -67
rect 400 -73 406 -67
rect 407 -73 413 -67
rect 414 -73 417 -67
rect 421 -73 424 -67
rect 463 -73 466 -67
rect 470 -73 473 -67
rect 477 -73 480 -67
rect 484 -73 487 -67
rect 491 -73 494 -67
rect 498 -73 501 -67
rect 505 -73 508 -67
rect 519 -73 522 -67
rect 533 -73 536 -67
rect 540 -73 546 -67
rect 547 -73 550 -67
rect 561 -73 567 -67
rect 568 -73 571 -67
rect 582 -73 588 -67
rect 589 -73 592 -67
rect 596 -73 599 -67
rect 603 -73 606 -67
rect 610 -73 613 -67
rect 617 -73 620 -67
rect 638 -73 641 -67
rect 645 -73 648 -67
rect 652 -73 658 -67
rect 659 -73 662 -67
rect 666 -73 669 -67
rect 673 -73 679 -67
rect 680 -73 683 -67
rect 687 -73 690 -67
rect 694 -73 700 -67
rect 701 -73 704 -67
rect 708 -73 711 -67
rect 715 -73 718 -67
rect 722 -73 725 -67
rect 729 -73 732 -67
rect 736 -73 742 -67
rect 743 -73 746 -67
rect 750 -73 753 -67
rect 757 -73 760 -67
rect 764 -73 767 -67
rect 771 -73 774 -67
rect 778 -73 781 -67
rect 785 -73 791 -67
rect 792 -73 795 -67
rect 799 -73 805 -67
rect 806 -73 809 -67
rect 813 -73 816 -67
rect 820 -73 823 -67
rect 827 -73 830 -67
rect 834 -73 837 -67
rect 841 -73 844 -67
rect 848 -73 854 -67
rect 855 -73 861 -67
rect 862 -73 865 -67
rect 869 -73 872 -67
rect 876 -73 879 -67
rect 883 -73 889 -67
rect 890 -73 893 -67
rect 897 -73 903 -67
rect 904 -73 910 -67
rect 911 -73 914 -67
rect 918 -73 921 -67
rect 925 -73 928 -67
rect 932 -73 935 -67
rect 939 -73 945 -67
rect 946 -73 949 -67
rect 953 -73 959 -67
rect 960 -73 963 -67
rect 967 -73 970 -67
rect 974 -73 977 -67
rect 981 -73 984 -67
rect 988 -73 991 -67
rect 995 -73 1001 -67
rect 1002 -73 1005 -67
rect 1009 -73 1012 -67
rect 1016 -73 1019 -67
rect 1023 -73 1029 -67
rect 1030 -73 1033 -67
rect 1037 -73 1040 -67
rect 1044 -73 1047 -67
rect 1051 -73 1054 -67
rect 1058 -73 1061 -67
rect 1065 -73 1071 -67
rect 1072 -73 1075 -67
rect 1079 -73 1082 -67
rect 1086 -73 1089 -67
rect 1093 -73 1096 -67
rect 1100 -73 1103 -67
rect 1107 -73 1113 -67
rect 1114 -73 1120 -67
rect 1121 -73 1127 -67
rect 1149 -73 1152 -67
rect 1163 -73 1169 -67
rect 1177 -73 1180 -67
rect 1212 -73 1215 -67
rect 1219 -73 1222 -67
rect 1226 -73 1232 -67
rect 1233 -73 1239 -67
rect 1289 -73 1292 -67
rect 1317 -73 1323 -67
rect 1331 -73 1334 -67
rect 1359 -73 1362 -67
rect 1485 -73 1488 -67
rect 1632 -73 1635 -67
rect 1758 -73 1761 -67
rect 1 -150 7 -144
rect 8 -150 14 -144
rect 57 -150 60 -144
rect 64 -150 67 -144
rect 71 -150 74 -144
rect 78 -150 81 -144
rect 85 -150 88 -144
rect 92 -150 95 -144
rect 99 -150 102 -144
rect 106 -150 109 -144
rect 113 -150 116 -144
rect 120 -150 126 -144
rect 127 -150 130 -144
rect 134 -150 137 -144
rect 141 -150 147 -144
rect 148 -150 154 -144
rect 155 -150 158 -144
rect 162 -150 165 -144
rect 169 -150 172 -144
rect 176 -150 179 -144
rect 183 -150 186 -144
rect 190 -150 193 -144
rect 197 -150 200 -144
rect 204 -150 207 -144
rect 211 -150 214 -144
rect 218 -150 221 -144
rect 225 -150 231 -144
rect 232 -150 238 -144
rect 239 -150 242 -144
rect 246 -150 249 -144
rect 253 -150 259 -144
rect 260 -150 266 -144
rect 267 -150 273 -144
rect 274 -150 277 -144
rect 281 -150 284 -144
rect 288 -150 291 -144
rect 295 -150 298 -144
rect 302 -150 305 -144
rect 309 -150 312 -144
rect 316 -150 319 -144
rect 323 -150 326 -144
rect 330 -150 333 -144
rect 337 -150 340 -144
rect 344 -150 347 -144
rect 351 -150 354 -144
rect 358 -150 361 -144
rect 365 -150 368 -144
rect 372 -150 375 -144
rect 379 -150 382 -144
rect 386 -150 392 -144
rect 393 -150 396 -144
rect 400 -150 403 -144
rect 407 -150 410 -144
rect 414 -150 417 -144
rect 421 -150 424 -144
rect 428 -150 431 -144
rect 435 -150 438 -144
rect 442 -150 448 -144
rect 449 -150 452 -144
rect 456 -150 462 -144
rect 463 -150 469 -144
rect 470 -150 476 -144
rect 477 -150 480 -144
rect 484 -150 487 -144
rect 491 -150 494 -144
rect 498 -150 501 -144
rect 505 -150 508 -144
rect 512 -150 515 -144
rect 519 -150 525 -144
rect 526 -150 532 -144
rect 533 -150 536 -144
rect 540 -150 543 -144
rect 547 -150 550 -144
rect 554 -150 557 -144
rect 561 -150 567 -144
rect 568 -150 571 -144
rect 575 -150 578 -144
rect 582 -150 585 -144
rect 589 -150 592 -144
rect 596 -150 602 -144
rect 603 -150 606 -144
rect 610 -150 613 -144
rect 617 -150 620 -144
rect 624 -150 627 -144
rect 631 -150 634 -144
rect 638 -150 641 -144
rect 645 -150 651 -144
rect 652 -150 655 -144
rect 659 -150 662 -144
rect 666 -150 669 -144
rect 673 -150 679 -144
rect 680 -150 686 -144
rect 687 -150 690 -144
rect 694 -150 700 -144
rect 701 -150 704 -144
rect 708 -150 711 -144
rect 715 -150 718 -144
rect 722 -150 725 -144
rect 729 -150 735 -144
rect 736 -150 742 -144
rect 743 -150 746 -144
rect 750 -150 753 -144
rect 757 -150 760 -144
rect 764 -150 770 -144
rect 771 -150 777 -144
rect 778 -150 781 -144
rect 785 -150 788 -144
rect 792 -150 795 -144
rect 799 -150 805 -144
rect 806 -150 809 -144
rect 813 -150 816 -144
rect 820 -150 823 -144
rect 827 -150 830 -144
rect 834 -150 840 -144
rect 841 -150 844 -144
rect 848 -150 851 -144
rect 855 -150 858 -144
rect 862 -150 865 -144
rect 869 -150 872 -144
rect 876 -150 879 -144
rect 883 -150 886 -144
rect 890 -150 893 -144
rect 897 -150 900 -144
rect 904 -150 907 -144
rect 911 -150 914 -144
rect 918 -150 921 -144
rect 925 -150 931 -144
rect 932 -150 938 -144
rect 939 -150 942 -144
rect 946 -150 952 -144
rect 953 -150 956 -144
rect 960 -150 966 -144
rect 967 -150 970 -144
rect 974 -150 980 -144
rect 981 -150 984 -144
rect 988 -150 991 -144
rect 995 -150 998 -144
rect 1002 -150 1005 -144
rect 1009 -150 1012 -144
rect 1016 -150 1019 -144
rect 1023 -150 1026 -144
rect 1030 -150 1033 -144
rect 1037 -150 1040 -144
rect 1044 -150 1047 -144
rect 1051 -150 1054 -144
rect 1058 -150 1061 -144
rect 1065 -150 1068 -144
rect 1072 -150 1078 -144
rect 1079 -150 1082 -144
rect 1086 -150 1092 -144
rect 1093 -150 1096 -144
rect 1100 -150 1103 -144
rect 1107 -150 1110 -144
rect 1114 -150 1117 -144
rect 1121 -150 1124 -144
rect 1128 -150 1131 -144
rect 1135 -150 1138 -144
rect 1142 -150 1148 -144
rect 1149 -150 1152 -144
rect 1156 -150 1159 -144
rect 1163 -150 1166 -144
rect 1170 -150 1176 -144
rect 1177 -150 1180 -144
rect 1184 -150 1187 -144
rect 1191 -150 1194 -144
rect 1198 -150 1201 -144
rect 1205 -150 1208 -144
rect 1212 -150 1215 -144
rect 1219 -150 1222 -144
rect 1226 -150 1229 -144
rect 1233 -150 1236 -144
rect 1240 -150 1243 -144
rect 1247 -150 1250 -144
rect 1254 -150 1257 -144
rect 1261 -150 1267 -144
rect 1268 -150 1271 -144
rect 1275 -150 1278 -144
rect 1282 -150 1285 -144
rect 1289 -150 1292 -144
rect 1296 -150 1299 -144
rect 1303 -150 1306 -144
rect 1310 -150 1313 -144
rect 1317 -150 1320 -144
rect 1324 -150 1327 -144
rect 1352 -150 1355 -144
rect 1359 -150 1362 -144
rect 1373 -150 1376 -144
rect 1422 -150 1425 -144
rect 1506 -150 1509 -144
rect 1513 -150 1516 -144
rect 1639 -150 1642 -144
rect 1884 -150 1887 -144
rect 1 -253 7 -247
rect 8 -253 14 -247
rect 15 -253 18 -247
rect 22 -253 25 -247
rect 29 -253 32 -247
rect 36 -253 39 -247
rect 43 -253 46 -247
rect 50 -253 53 -247
rect 57 -253 60 -247
rect 64 -253 70 -247
rect 71 -253 74 -247
rect 78 -253 84 -247
rect 85 -253 91 -247
rect 92 -253 95 -247
rect 99 -253 102 -247
rect 106 -253 109 -247
rect 113 -253 119 -247
rect 120 -253 123 -247
rect 127 -253 130 -247
rect 134 -253 140 -247
rect 141 -253 144 -247
rect 148 -253 151 -247
rect 155 -253 161 -247
rect 162 -253 165 -247
rect 169 -253 172 -247
rect 176 -253 179 -247
rect 183 -253 186 -247
rect 190 -253 196 -247
rect 197 -253 203 -247
rect 204 -253 210 -247
rect 211 -253 217 -247
rect 218 -253 221 -247
rect 225 -253 228 -247
rect 232 -253 235 -247
rect 239 -253 245 -247
rect 246 -253 249 -247
rect 253 -253 256 -247
rect 260 -253 263 -247
rect 267 -253 273 -247
rect 274 -253 277 -247
rect 281 -253 284 -247
rect 288 -253 291 -247
rect 295 -253 301 -247
rect 302 -253 305 -247
rect 309 -253 315 -247
rect 316 -253 319 -247
rect 323 -253 326 -247
rect 330 -253 333 -247
rect 337 -253 340 -247
rect 344 -253 347 -247
rect 351 -253 354 -247
rect 358 -253 361 -247
rect 365 -253 368 -247
rect 372 -253 375 -247
rect 379 -253 382 -247
rect 386 -253 389 -247
rect 393 -253 396 -247
rect 400 -253 403 -247
rect 407 -253 410 -247
rect 414 -253 417 -247
rect 421 -253 424 -247
rect 428 -253 431 -247
rect 435 -253 441 -247
rect 442 -253 445 -247
rect 449 -253 452 -247
rect 456 -253 459 -247
rect 463 -253 469 -247
rect 470 -253 473 -247
rect 477 -253 480 -247
rect 484 -253 487 -247
rect 491 -253 494 -247
rect 498 -253 501 -247
rect 505 -253 508 -247
rect 512 -253 515 -247
rect 519 -253 525 -247
rect 526 -253 529 -247
rect 533 -253 539 -247
rect 540 -253 543 -247
rect 547 -253 550 -247
rect 554 -253 557 -247
rect 561 -253 564 -247
rect 568 -253 571 -247
rect 575 -253 578 -247
rect 582 -253 585 -247
rect 589 -253 595 -247
rect 596 -253 599 -247
rect 603 -253 606 -247
rect 610 -253 613 -247
rect 617 -253 623 -247
rect 624 -253 627 -247
rect 631 -253 634 -247
rect 638 -253 641 -247
rect 645 -253 648 -247
rect 652 -253 655 -247
rect 659 -253 662 -247
rect 666 -253 669 -247
rect 673 -253 676 -247
rect 680 -253 683 -247
rect 687 -253 690 -247
rect 694 -253 697 -247
rect 701 -253 707 -247
rect 708 -253 714 -247
rect 715 -253 718 -247
rect 722 -253 725 -247
rect 729 -253 732 -247
rect 736 -253 739 -247
rect 743 -253 746 -247
rect 750 -253 753 -247
rect 757 -253 760 -247
rect 764 -253 767 -247
rect 771 -253 774 -247
rect 778 -253 781 -247
rect 785 -253 788 -247
rect 792 -253 795 -247
rect 799 -253 802 -247
rect 806 -253 809 -247
rect 813 -253 816 -247
rect 820 -253 823 -247
rect 827 -253 830 -247
rect 834 -253 837 -247
rect 841 -253 844 -247
rect 848 -253 851 -247
rect 855 -253 858 -247
rect 862 -253 865 -247
rect 869 -253 872 -247
rect 876 -253 879 -247
rect 883 -253 889 -247
rect 890 -253 896 -247
rect 897 -253 900 -247
rect 904 -253 907 -247
rect 911 -253 917 -247
rect 918 -253 921 -247
rect 925 -253 928 -247
rect 932 -253 935 -247
rect 939 -253 942 -247
rect 946 -253 949 -247
rect 953 -253 956 -247
rect 960 -253 963 -247
rect 967 -253 970 -247
rect 974 -253 977 -247
rect 981 -253 984 -247
rect 988 -253 994 -247
rect 995 -253 1001 -247
rect 1002 -253 1005 -247
rect 1009 -253 1015 -247
rect 1016 -253 1019 -247
rect 1023 -253 1026 -247
rect 1030 -253 1033 -247
rect 1037 -253 1040 -247
rect 1044 -253 1047 -247
rect 1051 -253 1054 -247
rect 1058 -253 1061 -247
rect 1065 -253 1068 -247
rect 1072 -253 1075 -247
rect 1079 -253 1082 -247
rect 1086 -253 1089 -247
rect 1093 -253 1096 -247
rect 1100 -253 1103 -247
rect 1107 -253 1110 -247
rect 1114 -253 1117 -247
rect 1121 -253 1124 -247
rect 1128 -253 1131 -247
rect 1135 -253 1138 -247
rect 1142 -253 1145 -247
rect 1149 -253 1155 -247
rect 1156 -253 1159 -247
rect 1163 -253 1166 -247
rect 1170 -253 1173 -247
rect 1177 -253 1183 -247
rect 1184 -253 1187 -247
rect 1191 -253 1194 -247
rect 1198 -253 1204 -247
rect 1205 -253 1208 -247
rect 1212 -253 1218 -247
rect 1219 -253 1222 -247
rect 1226 -253 1229 -247
rect 1233 -253 1236 -247
rect 1240 -253 1243 -247
rect 1247 -253 1250 -247
rect 1254 -253 1257 -247
rect 1261 -253 1264 -247
rect 1268 -253 1271 -247
rect 1275 -253 1278 -247
rect 1282 -253 1285 -247
rect 1289 -253 1292 -247
rect 1296 -253 1299 -247
rect 1303 -253 1306 -247
rect 1310 -253 1313 -247
rect 1317 -253 1320 -247
rect 1324 -253 1330 -247
rect 1331 -253 1334 -247
rect 1338 -253 1341 -247
rect 1345 -253 1348 -247
rect 1352 -253 1355 -247
rect 1359 -253 1362 -247
rect 1366 -253 1369 -247
rect 1373 -253 1376 -247
rect 1380 -253 1383 -247
rect 1387 -253 1390 -247
rect 1394 -253 1397 -247
rect 1401 -253 1404 -247
rect 1408 -253 1411 -247
rect 1415 -253 1418 -247
rect 1422 -253 1425 -247
rect 1429 -253 1432 -247
rect 1436 -253 1439 -247
rect 1443 -253 1446 -247
rect 1450 -253 1453 -247
rect 1457 -253 1460 -247
rect 1464 -253 1467 -247
rect 1471 -253 1474 -247
rect 1478 -253 1481 -247
rect 1485 -253 1488 -247
rect 1492 -253 1495 -247
rect 1499 -253 1502 -247
rect 1506 -253 1509 -247
rect 1513 -253 1516 -247
rect 1520 -253 1523 -247
rect 1527 -253 1530 -247
rect 1534 -253 1537 -247
rect 1541 -253 1547 -247
rect 1548 -253 1554 -247
rect 1555 -253 1558 -247
rect 1562 -253 1568 -247
rect 1569 -253 1572 -247
rect 1576 -253 1579 -247
rect 1583 -253 1586 -247
rect 1590 -253 1593 -247
rect 1611 -253 1617 -247
rect 1625 -253 1628 -247
rect 1632 -253 1635 -247
rect 1667 -253 1670 -247
rect 1814 -253 1817 -247
rect 1940 -253 1943 -247
rect 1 -378 7 -372
rect 8 -378 14 -372
rect 15 -378 18 -372
rect 22 -378 25 -372
rect 29 -378 32 -372
rect 36 -378 39 -372
rect 43 -378 49 -372
rect 50 -378 56 -372
rect 57 -378 60 -372
rect 64 -378 67 -372
rect 71 -378 74 -372
rect 78 -378 81 -372
rect 85 -378 88 -372
rect 92 -378 98 -372
rect 99 -378 102 -372
rect 106 -378 109 -372
rect 113 -378 116 -372
rect 120 -378 123 -372
rect 127 -378 130 -372
rect 134 -378 140 -372
rect 141 -378 144 -372
rect 148 -378 151 -372
rect 155 -378 158 -372
rect 162 -378 168 -372
rect 169 -378 172 -372
rect 176 -378 179 -372
rect 183 -378 189 -372
rect 190 -378 196 -372
rect 197 -378 200 -372
rect 204 -378 207 -372
rect 211 -378 214 -372
rect 218 -378 221 -372
rect 225 -378 228 -372
rect 232 -378 235 -372
rect 239 -378 245 -372
rect 246 -378 249 -372
rect 253 -378 256 -372
rect 260 -378 263 -372
rect 267 -378 270 -372
rect 274 -378 277 -372
rect 281 -378 284 -372
rect 288 -378 291 -372
rect 295 -378 298 -372
rect 302 -378 305 -372
rect 309 -378 312 -372
rect 316 -378 319 -372
rect 323 -378 326 -372
rect 330 -378 333 -372
rect 337 -378 340 -372
rect 344 -378 347 -372
rect 351 -378 354 -372
rect 358 -378 361 -372
rect 365 -378 368 -372
rect 372 -378 375 -372
rect 379 -378 382 -372
rect 386 -378 389 -372
rect 393 -378 396 -372
rect 400 -378 406 -372
rect 407 -378 410 -372
rect 414 -378 417 -372
rect 421 -378 424 -372
rect 428 -378 434 -372
rect 435 -378 438 -372
rect 442 -378 448 -372
rect 449 -378 452 -372
rect 456 -378 459 -372
rect 463 -378 466 -372
rect 470 -378 473 -372
rect 477 -378 483 -372
rect 484 -378 487 -372
rect 491 -378 494 -372
rect 498 -378 501 -372
rect 505 -378 508 -372
rect 512 -378 515 -372
rect 519 -378 522 -372
rect 526 -378 529 -372
rect 533 -378 536 -372
rect 540 -378 543 -372
rect 547 -378 550 -372
rect 554 -378 557 -372
rect 561 -378 564 -372
rect 568 -378 571 -372
rect 575 -378 578 -372
rect 582 -378 585 -372
rect 589 -378 592 -372
rect 596 -378 599 -372
rect 603 -378 606 -372
rect 610 -378 613 -372
rect 617 -378 620 -372
rect 624 -378 630 -372
rect 631 -378 637 -372
rect 638 -378 641 -372
rect 645 -378 651 -372
rect 652 -378 655 -372
rect 659 -378 662 -372
rect 666 -378 669 -372
rect 673 -378 676 -372
rect 680 -378 683 -372
rect 687 -378 690 -372
rect 694 -378 697 -372
rect 701 -378 704 -372
rect 708 -378 711 -372
rect 715 -378 718 -372
rect 722 -378 725 -372
rect 729 -378 732 -372
rect 736 -378 739 -372
rect 743 -378 749 -372
rect 750 -378 753 -372
rect 757 -378 763 -372
rect 764 -378 767 -372
rect 771 -378 777 -372
rect 778 -378 781 -372
rect 785 -378 788 -372
rect 792 -378 798 -372
rect 799 -378 805 -372
rect 806 -378 812 -372
rect 813 -378 816 -372
rect 820 -378 823 -372
rect 827 -378 830 -372
rect 834 -378 840 -372
rect 841 -378 847 -372
rect 848 -378 851 -372
rect 855 -378 858 -372
rect 862 -378 865 -372
rect 869 -378 872 -372
rect 876 -378 882 -372
rect 883 -378 886 -372
rect 890 -378 896 -372
rect 897 -378 900 -372
rect 904 -378 907 -372
rect 911 -378 914 -372
rect 918 -378 921 -372
rect 925 -378 928 -372
rect 932 -378 935 -372
rect 939 -378 942 -372
rect 946 -378 949 -372
rect 953 -378 956 -372
rect 960 -378 963 -372
rect 967 -378 970 -372
rect 974 -378 980 -372
rect 981 -378 984 -372
rect 988 -378 994 -372
rect 995 -378 998 -372
rect 1002 -378 1005 -372
rect 1009 -378 1012 -372
rect 1016 -378 1022 -372
rect 1023 -378 1029 -372
rect 1030 -378 1033 -372
rect 1037 -378 1040 -372
rect 1044 -378 1047 -372
rect 1051 -378 1054 -372
rect 1058 -378 1061 -372
rect 1065 -378 1068 -372
rect 1072 -378 1078 -372
rect 1079 -378 1085 -372
rect 1086 -378 1089 -372
rect 1093 -378 1096 -372
rect 1100 -378 1106 -372
rect 1107 -378 1110 -372
rect 1114 -378 1117 -372
rect 1121 -378 1124 -372
rect 1128 -378 1131 -372
rect 1135 -378 1138 -372
rect 1142 -378 1145 -372
rect 1149 -378 1152 -372
rect 1156 -378 1159 -372
rect 1163 -378 1166 -372
rect 1170 -378 1173 -372
rect 1177 -378 1183 -372
rect 1184 -378 1187 -372
rect 1191 -378 1194 -372
rect 1198 -378 1201 -372
rect 1205 -378 1208 -372
rect 1212 -378 1215 -372
rect 1219 -378 1222 -372
rect 1226 -378 1229 -372
rect 1233 -378 1236 -372
rect 1240 -378 1243 -372
rect 1247 -378 1250 -372
rect 1254 -378 1257 -372
rect 1261 -378 1264 -372
rect 1268 -378 1271 -372
rect 1275 -378 1278 -372
rect 1282 -378 1285 -372
rect 1289 -378 1292 -372
rect 1296 -378 1299 -372
rect 1303 -378 1306 -372
rect 1310 -378 1313 -372
rect 1317 -378 1320 -372
rect 1324 -378 1330 -372
rect 1331 -378 1334 -372
rect 1338 -378 1341 -372
rect 1345 -378 1348 -372
rect 1352 -378 1358 -372
rect 1359 -378 1362 -372
rect 1366 -378 1369 -372
rect 1373 -378 1376 -372
rect 1380 -378 1383 -372
rect 1387 -378 1390 -372
rect 1394 -378 1397 -372
rect 1401 -378 1404 -372
rect 1408 -378 1411 -372
rect 1415 -378 1418 -372
rect 1422 -378 1425 -372
rect 1429 -378 1432 -372
rect 1436 -378 1439 -372
rect 1443 -378 1446 -372
rect 1450 -378 1453 -372
rect 1457 -378 1460 -372
rect 1464 -378 1467 -372
rect 1471 -378 1474 -372
rect 1478 -378 1481 -372
rect 1485 -378 1488 -372
rect 1492 -378 1495 -372
rect 1499 -378 1502 -372
rect 1506 -378 1509 -372
rect 1513 -378 1516 -372
rect 1520 -378 1523 -372
rect 1527 -378 1530 -372
rect 1534 -378 1537 -372
rect 1541 -378 1544 -372
rect 1548 -378 1551 -372
rect 1555 -378 1558 -372
rect 1562 -378 1565 -372
rect 1569 -378 1572 -372
rect 1576 -378 1579 -372
rect 1583 -378 1586 -372
rect 1590 -378 1593 -372
rect 1597 -378 1600 -372
rect 1604 -378 1607 -372
rect 1611 -378 1617 -372
rect 1618 -378 1621 -372
rect 1625 -378 1628 -372
rect 1632 -378 1635 -372
rect 1639 -378 1642 -372
rect 1646 -378 1649 -372
rect 1653 -378 1656 -372
rect 1660 -378 1663 -372
rect 1667 -378 1670 -372
rect 1674 -378 1677 -372
rect 1681 -378 1684 -372
rect 1688 -378 1691 -372
rect 1695 -378 1698 -372
rect 1702 -378 1705 -372
rect 1709 -378 1712 -372
rect 1716 -378 1719 -372
rect 1723 -378 1726 -372
rect 1730 -378 1733 -372
rect 1737 -378 1740 -372
rect 1744 -378 1747 -372
rect 1751 -378 1754 -372
rect 1758 -378 1761 -372
rect 1765 -378 1768 -372
rect 1772 -378 1775 -372
rect 1779 -378 1782 -372
rect 1786 -378 1789 -372
rect 1793 -378 1796 -372
rect 1800 -378 1803 -372
rect 1807 -378 1810 -372
rect 1814 -378 1817 -372
rect 1821 -378 1824 -372
rect 1828 -378 1831 -372
rect 1835 -378 1838 -372
rect 1842 -378 1845 -372
rect 1926 -378 1929 -372
rect 1961 -378 1967 -372
rect 1968 -378 1971 -372
rect 1982 -378 1985 -372
rect 2003 -378 2006 -372
rect 2192 -378 2195 -372
rect 1 -507 4 -501
rect 8 -507 14 -501
rect 15 -507 18 -501
rect 22 -507 25 -501
rect 29 -507 35 -501
rect 36 -507 42 -501
rect 43 -507 46 -501
rect 50 -507 53 -501
rect 57 -507 63 -501
rect 64 -507 67 -501
rect 71 -507 74 -501
rect 78 -507 81 -501
rect 85 -507 88 -501
rect 92 -507 95 -501
rect 99 -507 102 -501
rect 106 -507 109 -501
rect 113 -507 119 -501
rect 120 -507 123 -501
rect 127 -507 130 -501
rect 134 -507 137 -501
rect 141 -507 144 -501
rect 148 -507 151 -501
rect 155 -507 158 -501
rect 162 -507 168 -501
rect 169 -507 175 -501
rect 176 -507 179 -501
rect 183 -507 186 -501
rect 190 -507 193 -501
rect 197 -507 200 -501
rect 204 -507 207 -501
rect 211 -507 217 -501
rect 218 -507 224 -501
rect 225 -507 228 -501
rect 232 -507 238 -501
rect 239 -507 242 -501
rect 246 -507 249 -501
rect 253 -507 256 -501
rect 260 -507 263 -501
rect 267 -507 270 -501
rect 274 -507 277 -501
rect 281 -507 284 -501
rect 288 -507 291 -501
rect 295 -507 298 -501
rect 302 -507 305 -501
rect 309 -507 312 -501
rect 316 -507 319 -501
rect 323 -507 326 -501
rect 330 -507 333 -501
rect 337 -507 340 -501
rect 344 -507 347 -501
rect 351 -507 354 -501
rect 358 -507 361 -501
rect 365 -507 368 -501
rect 372 -507 375 -501
rect 379 -507 382 -501
rect 386 -507 389 -501
rect 393 -507 396 -501
rect 400 -507 403 -501
rect 407 -507 410 -501
rect 414 -507 417 -501
rect 421 -507 424 -501
rect 428 -507 431 -501
rect 435 -507 438 -501
rect 442 -507 445 -501
rect 449 -507 452 -501
rect 456 -507 459 -501
rect 463 -507 466 -501
rect 470 -507 473 -501
rect 477 -507 480 -501
rect 484 -507 487 -501
rect 491 -507 497 -501
rect 498 -507 501 -501
rect 505 -507 508 -501
rect 512 -507 515 -501
rect 519 -507 522 -501
rect 526 -507 529 -501
rect 533 -507 539 -501
rect 540 -507 543 -501
rect 547 -507 550 -501
rect 554 -507 557 -501
rect 561 -507 564 -501
rect 568 -507 571 -501
rect 575 -507 578 -501
rect 582 -507 585 -501
rect 589 -507 592 -501
rect 596 -507 602 -501
rect 603 -507 606 -501
rect 610 -507 613 -501
rect 617 -507 623 -501
rect 624 -507 627 -501
rect 631 -507 637 -501
rect 638 -507 641 -501
rect 645 -507 648 -501
rect 652 -507 658 -501
rect 659 -507 662 -501
rect 666 -507 669 -501
rect 673 -507 676 -501
rect 680 -507 683 -501
rect 687 -507 690 -501
rect 694 -507 697 -501
rect 701 -507 704 -501
rect 708 -507 711 -501
rect 715 -507 721 -501
rect 722 -507 728 -501
rect 729 -507 732 -501
rect 736 -507 742 -501
rect 743 -507 746 -501
rect 750 -507 753 -501
rect 757 -507 760 -501
rect 764 -507 767 -501
rect 771 -507 774 -501
rect 778 -507 781 -501
rect 785 -507 788 -501
rect 792 -507 795 -501
rect 799 -507 802 -501
rect 806 -507 809 -501
rect 813 -507 816 -501
rect 820 -507 823 -501
rect 827 -507 830 -501
rect 834 -507 837 -501
rect 841 -507 844 -501
rect 848 -507 854 -501
rect 855 -507 858 -501
rect 862 -507 865 -501
rect 869 -507 872 -501
rect 876 -507 879 -501
rect 883 -507 889 -501
rect 890 -507 893 -501
rect 897 -507 900 -501
rect 904 -507 907 -501
rect 911 -507 917 -501
rect 918 -507 921 -501
rect 925 -507 928 -501
rect 932 -507 938 -501
rect 939 -507 942 -501
rect 946 -507 949 -501
rect 953 -507 959 -501
rect 960 -507 963 -501
rect 967 -507 973 -501
rect 974 -507 980 -501
rect 981 -507 987 -501
rect 988 -507 994 -501
rect 995 -507 998 -501
rect 1002 -507 1008 -501
rect 1009 -507 1012 -501
rect 1016 -507 1019 -501
rect 1023 -507 1029 -501
rect 1030 -507 1033 -501
rect 1037 -507 1040 -501
rect 1044 -507 1047 -501
rect 1051 -507 1054 -501
rect 1058 -507 1061 -501
rect 1065 -507 1068 -501
rect 1072 -507 1075 -501
rect 1079 -507 1085 -501
rect 1086 -507 1089 -501
rect 1093 -507 1096 -501
rect 1100 -507 1103 -501
rect 1107 -507 1110 -501
rect 1114 -507 1117 -501
rect 1121 -507 1127 -501
rect 1128 -507 1131 -501
rect 1135 -507 1138 -501
rect 1142 -507 1145 -501
rect 1149 -507 1152 -501
rect 1156 -507 1159 -501
rect 1163 -507 1169 -501
rect 1170 -507 1173 -501
rect 1177 -507 1180 -501
rect 1184 -507 1187 -501
rect 1191 -507 1194 -501
rect 1198 -507 1201 -501
rect 1205 -507 1208 -501
rect 1212 -507 1215 -501
rect 1219 -507 1222 -501
rect 1226 -507 1229 -501
rect 1233 -507 1236 -501
rect 1240 -507 1243 -501
rect 1247 -507 1250 -501
rect 1254 -507 1257 -501
rect 1261 -507 1264 -501
rect 1268 -507 1271 -501
rect 1275 -507 1278 -501
rect 1282 -507 1285 -501
rect 1289 -507 1292 -501
rect 1296 -507 1299 -501
rect 1303 -507 1306 -501
rect 1310 -507 1313 -501
rect 1317 -507 1320 -501
rect 1324 -507 1327 -501
rect 1331 -507 1334 -501
rect 1338 -507 1341 -501
rect 1345 -507 1348 -501
rect 1352 -507 1355 -501
rect 1359 -507 1362 -501
rect 1366 -507 1369 -501
rect 1373 -507 1376 -501
rect 1380 -507 1383 -501
rect 1387 -507 1390 -501
rect 1394 -507 1397 -501
rect 1401 -507 1404 -501
rect 1408 -507 1411 -501
rect 1415 -507 1418 -501
rect 1422 -507 1425 -501
rect 1429 -507 1432 -501
rect 1436 -507 1442 -501
rect 1443 -507 1446 -501
rect 1450 -507 1453 -501
rect 1457 -507 1460 -501
rect 1464 -507 1467 -501
rect 1471 -507 1474 -501
rect 1478 -507 1481 -501
rect 1485 -507 1488 -501
rect 1492 -507 1495 -501
rect 1499 -507 1502 -501
rect 1506 -507 1509 -501
rect 1513 -507 1516 -501
rect 1520 -507 1523 -501
rect 1527 -507 1530 -501
rect 1534 -507 1537 -501
rect 1541 -507 1544 -501
rect 1548 -507 1551 -501
rect 1555 -507 1558 -501
rect 1562 -507 1565 -501
rect 1569 -507 1572 -501
rect 1576 -507 1579 -501
rect 1583 -507 1586 -501
rect 1590 -507 1593 -501
rect 1597 -507 1600 -501
rect 1604 -507 1607 -501
rect 1611 -507 1614 -501
rect 1618 -507 1621 -501
rect 1625 -507 1628 -501
rect 1632 -507 1635 -501
rect 1639 -507 1642 -501
rect 1646 -507 1649 -501
rect 1653 -507 1656 -501
rect 1660 -507 1663 -501
rect 1667 -507 1670 -501
rect 1674 -507 1677 -501
rect 1681 -507 1684 -501
rect 1688 -507 1691 -501
rect 1695 -507 1698 -501
rect 1702 -507 1705 -501
rect 1709 -507 1712 -501
rect 1716 -507 1719 -501
rect 1723 -507 1726 -501
rect 1730 -507 1733 -501
rect 1737 -507 1740 -501
rect 1744 -507 1747 -501
rect 1751 -507 1754 -501
rect 1758 -507 1761 -501
rect 1765 -507 1768 -501
rect 1772 -507 1775 -501
rect 1779 -507 1782 -501
rect 1786 -507 1789 -501
rect 1793 -507 1796 -501
rect 1800 -507 1803 -501
rect 1807 -507 1810 -501
rect 1814 -507 1817 -501
rect 1821 -507 1824 -501
rect 1828 -507 1831 -501
rect 1835 -507 1838 -501
rect 1842 -507 1845 -501
rect 1849 -507 1852 -501
rect 1856 -507 1859 -501
rect 1863 -507 1866 -501
rect 1870 -507 1873 -501
rect 1877 -507 1880 -501
rect 1884 -507 1887 -501
rect 1891 -507 1894 -501
rect 1898 -507 1901 -501
rect 1905 -507 1908 -501
rect 1912 -507 1915 -501
rect 1919 -507 1922 -501
rect 1926 -507 1929 -501
rect 1933 -507 1936 -501
rect 1940 -507 1943 -501
rect 1947 -507 1950 -501
rect 1954 -507 1960 -501
rect 1961 -507 1964 -501
rect 1968 -507 1971 -501
rect 1975 -507 1981 -501
rect 1982 -507 1985 -501
rect 1989 -507 1992 -501
rect 1996 -507 1999 -501
rect 2003 -507 2009 -501
rect 2010 -507 2016 -501
rect 2017 -507 2023 -501
rect 2038 -507 2041 -501
rect 2087 -507 2090 -501
rect 2115 -507 2118 -501
rect 2143 -507 2146 -501
rect 2262 -507 2265 -501
rect 2283 -507 2286 -501
rect 1 -640 7 -634
rect 8 -640 11 -634
rect 15 -640 18 -634
rect 22 -640 25 -634
rect 29 -640 32 -634
rect 36 -640 39 -634
rect 43 -640 46 -634
rect 50 -640 53 -634
rect 57 -640 63 -634
rect 64 -640 67 -634
rect 71 -640 77 -634
rect 78 -640 81 -634
rect 85 -640 88 -634
rect 92 -640 95 -634
rect 99 -640 105 -634
rect 106 -640 109 -634
rect 113 -640 116 -634
rect 120 -640 123 -634
rect 127 -640 130 -634
rect 134 -640 140 -634
rect 141 -640 144 -634
rect 148 -640 151 -634
rect 155 -640 158 -634
rect 162 -640 165 -634
rect 169 -640 175 -634
rect 176 -640 179 -634
rect 183 -640 186 -634
rect 190 -640 193 -634
rect 197 -640 200 -634
rect 204 -640 210 -634
rect 211 -640 214 -634
rect 218 -640 221 -634
rect 225 -640 228 -634
rect 232 -640 235 -634
rect 239 -640 242 -634
rect 246 -640 252 -634
rect 253 -640 256 -634
rect 260 -640 263 -634
rect 267 -640 273 -634
rect 274 -640 277 -634
rect 281 -640 284 -634
rect 288 -640 291 -634
rect 295 -640 298 -634
rect 302 -640 305 -634
rect 309 -640 312 -634
rect 316 -640 319 -634
rect 323 -640 326 -634
rect 330 -640 333 -634
rect 337 -640 340 -634
rect 344 -640 347 -634
rect 351 -640 354 -634
rect 358 -640 361 -634
rect 365 -640 368 -634
rect 372 -640 375 -634
rect 379 -640 382 -634
rect 386 -640 389 -634
rect 393 -640 396 -634
rect 400 -640 403 -634
rect 407 -640 410 -634
rect 414 -640 417 -634
rect 421 -640 424 -634
rect 428 -640 434 -634
rect 435 -640 438 -634
rect 442 -640 445 -634
rect 449 -640 452 -634
rect 456 -640 459 -634
rect 463 -640 466 -634
rect 470 -640 473 -634
rect 477 -640 480 -634
rect 484 -640 487 -634
rect 491 -640 494 -634
rect 498 -640 501 -634
rect 505 -640 508 -634
rect 512 -640 515 -634
rect 519 -640 522 -634
rect 526 -640 529 -634
rect 533 -640 539 -634
rect 540 -640 543 -634
rect 547 -640 550 -634
rect 554 -640 557 -634
rect 561 -640 567 -634
rect 568 -640 571 -634
rect 575 -640 578 -634
rect 582 -640 588 -634
rect 589 -640 595 -634
rect 596 -640 599 -634
rect 603 -640 606 -634
rect 610 -640 613 -634
rect 617 -640 620 -634
rect 624 -640 627 -634
rect 631 -640 634 -634
rect 638 -640 641 -634
rect 645 -640 651 -634
rect 652 -640 655 -634
rect 659 -640 665 -634
rect 666 -640 669 -634
rect 673 -640 676 -634
rect 680 -640 683 -634
rect 687 -640 690 -634
rect 694 -640 697 -634
rect 701 -640 704 -634
rect 708 -640 711 -634
rect 715 -640 718 -634
rect 722 -640 725 -634
rect 729 -640 735 -634
rect 736 -640 739 -634
rect 743 -640 749 -634
rect 750 -640 753 -634
rect 757 -640 760 -634
rect 764 -640 767 -634
rect 771 -640 774 -634
rect 778 -640 781 -634
rect 785 -640 791 -634
rect 792 -640 795 -634
rect 799 -640 802 -634
rect 806 -640 812 -634
rect 813 -640 816 -634
rect 820 -640 826 -634
rect 827 -640 830 -634
rect 834 -640 837 -634
rect 841 -640 844 -634
rect 848 -640 854 -634
rect 855 -640 858 -634
rect 862 -640 865 -634
rect 869 -640 872 -634
rect 876 -640 879 -634
rect 883 -640 886 -634
rect 890 -640 893 -634
rect 897 -640 900 -634
rect 904 -640 907 -634
rect 911 -640 914 -634
rect 918 -640 921 -634
rect 925 -640 931 -634
rect 932 -640 935 -634
rect 939 -640 945 -634
rect 946 -640 949 -634
rect 953 -640 956 -634
rect 960 -640 963 -634
rect 967 -640 970 -634
rect 974 -640 977 -634
rect 981 -640 987 -634
rect 988 -640 991 -634
rect 995 -640 998 -634
rect 1002 -640 1005 -634
rect 1009 -640 1015 -634
rect 1016 -640 1019 -634
rect 1023 -640 1026 -634
rect 1030 -640 1036 -634
rect 1037 -640 1040 -634
rect 1044 -640 1047 -634
rect 1051 -640 1054 -634
rect 1058 -640 1064 -634
rect 1065 -640 1068 -634
rect 1072 -640 1075 -634
rect 1079 -640 1085 -634
rect 1086 -640 1089 -634
rect 1093 -640 1099 -634
rect 1100 -640 1103 -634
rect 1107 -640 1110 -634
rect 1114 -640 1117 -634
rect 1121 -640 1124 -634
rect 1128 -640 1131 -634
rect 1135 -640 1138 -634
rect 1142 -640 1148 -634
rect 1149 -640 1155 -634
rect 1156 -640 1159 -634
rect 1163 -640 1166 -634
rect 1170 -640 1173 -634
rect 1177 -640 1180 -634
rect 1184 -640 1187 -634
rect 1191 -640 1194 -634
rect 1198 -640 1204 -634
rect 1205 -640 1208 -634
rect 1212 -640 1218 -634
rect 1219 -640 1222 -634
rect 1226 -640 1229 -634
rect 1233 -640 1236 -634
rect 1240 -640 1243 -634
rect 1247 -640 1250 -634
rect 1254 -640 1257 -634
rect 1261 -640 1264 -634
rect 1268 -640 1271 -634
rect 1275 -640 1278 -634
rect 1282 -640 1285 -634
rect 1289 -640 1292 -634
rect 1296 -640 1302 -634
rect 1303 -640 1306 -634
rect 1310 -640 1313 -634
rect 1317 -640 1320 -634
rect 1324 -640 1327 -634
rect 1331 -640 1334 -634
rect 1338 -640 1341 -634
rect 1345 -640 1348 -634
rect 1352 -640 1355 -634
rect 1359 -640 1362 -634
rect 1366 -640 1369 -634
rect 1373 -640 1376 -634
rect 1380 -640 1383 -634
rect 1387 -640 1390 -634
rect 1394 -640 1397 -634
rect 1401 -640 1404 -634
rect 1408 -640 1411 -634
rect 1415 -640 1418 -634
rect 1422 -640 1425 -634
rect 1429 -640 1432 -634
rect 1436 -640 1439 -634
rect 1443 -640 1446 -634
rect 1450 -640 1453 -634
rect 1457 -640 1460 -634
rect 1464 -640 1467 -634
rect 1471 -640 1474 -634
rect 1478 -640 1481 -634
rect 1485 -640 1491 -634
rect 1492 -640 1495 -634
rect 1499 -640 1502 -634
rect 1506 -640 1509 -634
rect 1513 -640 1516 -634
rect 1520 -640 1523 -634
rect 1527 -640 1530 -634
rect 1534 -640 1537 -634
rect 1541 -640 1544 -634
rect 1548 -640 1551 -634
rect 1555 -640 1558 -634
rect 1562 -640 1565 -634
rect 1569 -640 1572 -634
rect 1576 -640 1579 -634
rect 1583 -640 1586 -634
rect 1590 -640 1593 -634
rect 1597 -640 1600 -634
rect 1604 -640 1607 -634
rect 1611 -640 1614 -634
rect 1618 -640 1621 -634
rect 1625 -640 1628 -634
rect 1632 -640 1635 -634
rect 1639 -640 1642 -634
rect 1646 -640 1649 -634
rect 1653 -640 1656 -634
rect 1660 -640 1663 -634
rect 1667 -640 1670 -634
rect 1674 -640 1677 -634
rect 1681 -640 1684 -634
rect 1688 -640 1691 -634
rect 1695 -640 1698 -634
rect 1702 -640 1705 -634
rect 1709 -640 1712 -634
rect 1716 -640 1719 -634
rect 1723 -640 1726 -634
rect 1730 -640 1733 -634
rect 1737 -640 1740 -634
rect 1744 -640 1747 -634
rect 1751 -640 1754 -634
rect 1758 -640 1761 -634
rect 1765 -640 1768 -634
rect 1772 -640 1775 -634
rect 1779 -640 1782 -634
rect 1786 -640 1789 -634
rect 1793 -640 1796 -634
rect 1800 -640 1803 -634
rect 1807 -640 1810 -634
rect 1814 -640 1817 -634
rect 1821 -640 1824 -634
rect 1828 -640 1831 -634
rect 1835 -640 1838 -634
rect 1842 -640 1845 -634
rect 1849 -640 1852 -634
rect 1856 -640 1859 -634
rect 1863 -640 1866 -634
rect 1870 -640 1873 -634
rect 1877 -640 1880 -634
rect 1884 -640 1887 -634
rect 1891 -640 1894 -634
rect 1898 -640 1901 -634
rect 1905 -640 1908 -634
rect 1912 -640 1915 -634
rect 1919 -640 1922 -634
rect 1926 -640 1929 -634
rect 1933 -640 1936 -634
rect 1940 -640 1943 -634
rect 1947 -640 1950 -634
rect 1954 -640 1957 -634
rect 1961 -640 1964 -634
rect 1968 -640 1971 -634
rect 1975 -640 1978 -634
rect 1982 -640 1985 -634
rect 1989 -640 1992 -634
rect 1996 -640 1999 -634
rect 2003 -640 2006 -634
rect 2010 -640 2013 -634
rect 2017 -640 2020 -634
rect 2024 -640 2027 -634
rect 2031 -640 2034 -634
rect 2038 -640 2041 -634
rect 2045 -640 2048 -634
rect 2052 -640 2055 -634
rect 2059 -640 2062 -634
rect 2066 -640 2069 -634
rect 2073 -640 2076 -634
rect 2080 -640 2083 -634
rect 2087 -640 2090 -634
rect 2094 -640 2097 -634
rect 2101 -640 2104 -634
rect 2108 -640 2111 -634
rect 2115 -640 2118 -634
rect 2122 -640 2125 -634
rect 2129 -640 2132 -634
rect 2136 -640 2139 -634
rect 2143 -640 2146 -634
rect 2150 -640 2153 -634
rect 2157 -640 2160 -634
rect 2164 -640 2167 -634
rect 2171 -640 2174 -634
rect 2178 -640 2181 -634
rect 2185 -640 2188 -634
rect 2192 -640 2195 -634
rect 2199 -640 2202 -634
rect 2206 -640 2212 -634
rect 2213 -640 2219 -634
rect 2220 -640 2226 -634
rect 2290 -640 2293 -634
rect 2325 -640 2328 -634
rect 2360 -640 2363 -634
rect 1 -817 4 -811
rect 8 -817 14 -811
rect 15 -817 21 -811
rect 22 -817 25 -811
rect 29 -817 32 -811
rect 36 -817 39 -811
rect 43 -817 49 -811
rect 50 -817 53 -811
rect 57 -817 60 -811
rect 64 -817 70 -811
rect 71 -817 74 -811
rect 78 -817 84 -811
rect 85 -817 88 -811
rect 92 -817 95 -811
rect 99 -817 102 -811
rect 106 -817 109 -811
rect 113 -817 116 -811
rect 120 -817 126 -811
rect 127 -817 133 -811
rect 134 -817 137 -811
rect 141 -817 147 -811
rect 148 -817 151 -811
rect 155 -817 158 -811
rect 162 -817 165 -811
rect 169 -817 172 -811
rect 176 -817 179 -811
rect 183 -817 189 -811
rect 190 -817 193 -811
rect 197 -817 200 -811
rect 204 -817 210 -811
rect 211 -817 214 -811
rect 218 -817 224 -811
rect 225 -817 228 -811
rect 232 -817 238 -811
rect 239 -817 242 -811
rect 246 -817 249 -811
rect 253 -817 256 -811
rect 260 -817 263 -811
rect 267 -817 270 -811
rect 274 -817 277 -811
rect 281 -817 284 -811
rect 288 -817 291 -811
rect 295 -817 298 -811
rect 302 -817 305 -811
rect 309 -817 312 -811
rect 316 -817 319 -811
rect 323 -817 326 -811
rect 330 -817 333 -811
rect 337 -817 340 -811
rect 344 -817 347 -811
rect 351 -817 354 -811
rect 358 -817 364 -811
rect 365 -817 368 -811
rect 372 -817 375 -811
rect 379 -817 382 -811
rect 386 -817 389 -811
rect 393 -817 396 -811
rect 400 -817 403 -811
rect 407 -817 410 -811
rect 414 -817 417 -811
rect 421 -817 424 -811
rect 428 -817 431 -811
rect 435 -817 438 -811
rect 442 -817 445 -811
rect 449 -817 452 -811
rect 456 -817 459 -811
rect 463 -817 466 -811
rect 470 -817 473 -811
rect 477 -817 480 -811
rect 484 -817 487 -811
rect 491 -817 494 -811
rect 498 -817 501 -811
rect 505 -817 508 -811
rect 512 -817 515 -811
rect 519 -817 525 -811
rect 526 -817 529 -811
rect 533 -817 536 -811
rect 540 -817 543 -811
rect 547 -817 550 -811
rect 554 -817 557 -811
rect 561 -817 564 -811
rect 568 -817 571 -811
rect 575 -817 578 -811
rect 582 -817 588 -811
rect 589 -817 595 -811
rect 596 -817 599 -811
rect 603 -817 606 -811
rect 610 -817 613 -811
rect 617 -817 620 -811
rect 624 -817 627 -811
rect 631 -817 634 -811
rect 638 -817 641 -811
rect 645 -817 648 -811
rect 652 -817 655 -811
rect 659 -817 662 -811
rect 666 -817 669 -811
rect 673 -817 676 -811
rect 680 -817 686 -811
rect 687 -817 690 -811
rect 694 -817 700 -811
rect 701 -817 704 -811
rect 708 -817 711 -811
rect 715 -817 718 -811
rect 722 -817 728 -811
rect 729 -817 732 -811
rect 736 -817 739 -811
rect 743 -817 749 -811
rect 750 -817 756 -811
rect 757 -817 760 -811
rect 764 -817 767 -811
rect 771 -817 774 -811
rect 778 -817 781 -811
rect 785 -817 788 -811
rect 792 -817 795 -811
rect 799 -817 802 -811
rect 806 -817 809 -811
rect 813 -817 816 -811
rect 820 -817 823 -811
rect 827 -817 833 -811
rect 834 -817 837 -811
rect 841 -817 844 -811
rect 848 -817 851 -811
rect 855 -817 858 -811
rect 862 -817 865 -811
rect 869 -817 872 -811
rect 876 -817 882 -811
rect 883 -817 886 -811
rect 890 -817 893 -811
rect 897 -817 900 -811
rect 904 -817 907 -811
rect 911 -817 914 -811
rect 918 -817 921 -811
rect 925 -817 928 -811
rect 932 -817 935 -811
rect 939 -817 942 -811
rect 946 -817 949 -811
rect 953 -817 959 -811
rect 960 -817 963 -811
rect 967 -817 970 -811
rect 974 -817 977 -811
rect 981 -817 984 -811
rect 988 -817 991 -811
rect 995 -817 998 -811
rect 1002 -817 1005 -811
rect 1009 -817 1015 -811
rect 1016 -817 1019 -811
rect 1023 -817 1026 -811
rect 1030 -817 1033 -811
rect 1037 -817 1040 -811
rect 1044 -817 1047 -811
rect 1051 -817 1054 -811
rect 1058 -817 1061 -811
rect 1065 -817 1068 -811
rect 1072 -817 1075 -811
rect 1079 -817 1082 -811
rect 1086 -817 1089 -811
rect 1093 -817 1099 -811
rect 1100 -817 1103 -811
rect 1107 -817 1113 -811
rect 1114 -817 1117 -811
rect 1121 -817 1124 -811
rect 1128 -817 1134 -811
rect 1135 -817 1141 -811
rect 1142 -817 1148 -811
rect 1149 -817 1152 -811
rect 1156 -817 1162 -811
rect 1163 -817 1166 -811
rect 1170 -817 1176 -811
rect 1177 -817 1180 -811
rect 1184 -817 1187 -811
rect 1191 -817 1194 -811
rect 1198 -817 1201 -811
rect 1205 -817 1211 -811
rect 1212 -817 1218 -811
rect 1219 -817 1225 -811
rect 1226 -817 1229 -811
rect 1233 -817 1236 -811
rect 1240 -817 1243 -811
rect 1247 -817 1250 -811
rect 1254 -817 1257 -811
rect 1261 -817 1264 -811
rect 1268 -817 1271 -811
rect 1275 -817 1278 -811
rect 1282 -817 1285 -811
rect 1289 -817 1292 -811
rect 1296 -817 1299 -811
rect 1303 -817 1306 -811
rect 1310 -817 1313 -811
rect 1317 -817 1320 -811
rect 1324 -817 1327 -811
rect 1331 -817 1337 -811
rect 1338 -817 1341 -811
rect 1345 -817 1348 -811
rect 1352 -817 1355 -811
rect 1359 -817 1365 -811
rect 1366 -817 1372 -811
rect 1373 -817 1376 -811
rect 1380 -817 1383 -811
rect 1387 -817 1390 -811
rect 1394 -817 1397 -811
rect 1401 -817 1404 -811
rect 1408 -817 1411 -811
rect 1415 -817 1418 -811
rect 1422 -817 1425 -811
rect 1429 -817 1432 -811
rect 1436 -817 1439 -811
rect 1443 -817 1446 -811
rect 1450 -817 1453 -811
rect 1457 -817 1460 -811
rect 1464 -817 1467 -811
rect 1471 -817 1474 -811
rect 1478 -817 1481 -811
rect 1485 -817 1488 -811
rect 1492 -817 1495 -811
rect 1499 -817 1502 -811
rect 1506 -817 1509 -811
rect 1513 -817 1516 -811
rect 1520 -817 1523 -811
rect 1527 -817 1530 -811
rect 1534 -817 1540 -811
rect 1541 -817 1544 -811
rect 1548 -817 1551 -811
rect 1555 -817 1558 -811
rect 1562 -817 1565 -811
rect 1569 -817 1572 -811
rect 1576 -817 1579 -811
rect 1583 -817 1586 -811
rect 1590 -817 1593 -811
rect 1597 -817 1600 -811
rect 1604 -817 1607 -811
rect 1611 -817 1614 -811
rect 1618 -817 1621 -811
rect 1625 -817 1628 -811
rect 1632 -817 1635 -811
rect 1639 -817 1642 -811
rect 1646 -817 1649 -811
rect 1653 -817 1656 -811
rect 1660 -817 1663 -811
rect 1667 -817 1670 -811
rect 1674 -817 1677 -811
rect 1681 -817 1684 -811
rect 1688 -817 1691 -811
rect 1695 -817 1698 -811
rect 1702 -817 1705 -811
rect 1709 -817 1712 -811
rect 1716 -817 1719 -811
rect 1723 -817 1726 -811
rect 1730 -817 1733 -811
rect 1737 -817 1740 -811
rect 1744 -817 1747 -811
rect 1751 -817 1754 -811
rect 1758 -817 1761 -811
rect 1765 -817 1768 -811
rect 1772 -817 1775 -811
rect 1779 -817 1782 -811
rect 1786 -817 1789 -811
rect 1793 -817 1796 -811
rect 1800 -817 1803 -811
rect 1807 -817 1810 -811
rect 1814 -817 1817 -811
rect 1821 -817 1824 -811
rect 1828 -817 1831 -811
rect 1835 -817 1838 -811
rect 1842 -817 1845 -811
rect 1849 -817 1852 -811
rect 1856 -817 1859 -811
rect 1863 -817 1866 -811
rect 1870 -817 1873 -811
rect 1877 -817 1880 -811
rect 1884 -817 1887 -811
rect 1891 -817 1894 -811
rect 1898 -817 1901 -811
rect 1905 -817 1908 -811
rect 1912 -817 1915 -811
rect 1919 -817 1922 -811
rect 1926 -817 1929 -811
rect 1933 -817 1936 -811
rect 1940 -817 1943 -811
rect 1947 -817 1950 -811
rect 1954 -817 1957 -811
rect 1961 -817 1964 -811
rect 1968 -817 1971 -811
rect 1975 -817 1978 -811
rect 1982 -817 1985 -811
rect 1989 -817 1992 -811
rect 1996 -817 1999 -811
rect 2003 -817 2006 -811
rect 2010 -817 2013 -811
rect 2017 -817 2020 -811
rect 2024 -817 2027 -811
rect 2031 -817 2034 -811
rect 2038 -817 2041 -811
rect 2045 -817 2048 -811
rect 2052 -817 2055 -811
rect 2059 -817 2062 -811
rect 2066 -817 2069 -811
rect 2073 -817 2076 -811
rect 2080 -817 2083 -811
rect 2087 -817 2090 -811
rect 2094 -817 2097 -811
rect 2101 -817 2104 -811
rect 2108 -817 2111 -811
rect 2115 -817 2118 -811
rect 2122 -817 2125 -811
rect 2129 -817 2132 -811
rect 2136 -817 2139 -811
rect 2143 -817 2146 -811
rect 2150 -817 2153 -811
rect 2157 -817 2160 -811
rect 2164 -817 2167 -811
rect 2171 -817 2174 -811
rect 2178 -817 2181 -811
rect 2185 -817 2188 -811
rect 2192 -817 2195 -811
rect 2199 -817 2202 -811
rect 2206 -817 2209 -811
rect 2213 -817 2216 -811
rect 2220 -817 2223 -811
rect 2227 -817 2230 -811
rect 2234 -817 2237 -811
rect 2241 -817 2244 -811
rect 2248 -817 2251 -811
rect 2255 -817 2258 -811
rect 2262 -817 2265 -811
rect 2269 -817 2272 -811
rect 2276 -817 2279 -811
rect 2283 -817 2286 -811
rect 2290 -817 2293 -811
rect 2297 -817 2300 -811
rect 2304 -817 2307 -811
rect 2311 -817 2314 -811
rect 2318 -817 2321 -811
rect 2325 -817 2328 -811
rect 2346 -817 2349 -811
rect 2402 -817 2405 -811
rect 1 -1006 4 -1000
rect 8 -1006 11 -1000
rect 15 -1006 18 -1000
rect 22 -1006 25 -1000
rect 29 -1006 32 -1000
rect 36 -1006 39 -1000
rect 43 -1006 46 -1000
rect 50 -1006 53 -1000
rect 57 -1006 60 -1000
rect 64 -1006 67 -1000
rect 71 -1006 74 -1000
rect 78 -1006 81 -1000
rect 85 -1006 88 -1000
rect 92 -1006 98 -1000
rect 99 -1006 105 -1000
rect 106 -1006 109 -1000
rect 113 -1006 116 -1000
rect 120 -1006 123 -1000
rect 127 -1006 130 -1000
rect 134 -1006 140 -1000
rect 141 -1006 144 -1000
rect 148 -1006 151 -1000
rect 155 -1006 158 -1000
rect 162 -1006 165 -1000
rect 169 -1006 172 -1000
rect 176 -1006 182 -1000
rect 183 -1006 189 -1000
rect 190 -1006 193 -1000
rect 197 -1006 200 -1000
rect 204 -1006 207 -1000
rect 211 -1006 214 -1000
rect 218 -1006 224 -1000
rect 225 -1006 228 -1000
rect 232 -1006 235 -1000
rect 239 -1006 242 -1000
rect 246 -1006 249 -1000
rect 253 -1006 256 -1000
rect 260 -1006 263 -1000
rect 267 -1006 273 -1000
rect 274 -1006 277 -1000
rect 281 -1006 284 -1000
rect 288 -1006 291 -1000
rect 295 -1006 298 -1000
rect 302 -1006 305 -1000
rect 309 -1006 312 -1000
rect 316 -1006 319 -1000
rect 323 -1006 326 -1000
rect 330 -1006 333 -1000
rect 337 -1006 340 -1000
rect 344 -1006 347 -1000
rect 351 -1006 354 -1000
rect 358 -1006 361 -1000
rect 365 -1006 368 -1000
rect 372 -1006 378 -1000
rect 379 -1006 382 -1000
rect 386 -1006 392 -1000
rect 393 -1006 396 -1000
rect 400 -1006 403 -1000
rect 407 -1006 410 -1000
rect 414 -1006 417 -1000
rect 421 -1006 424 -1000
rect 428 -1006 431 -1000
rect 435 -1006 438 -1000
rect 442 -1006 445 -1000
rect 449 -1006 452 -1000
rect 456 -1006 459 -1000
rect 463 -1006 466 -1000
rect 470 -1006 473 -1000
rect 477 -1006 480 -1000
rect 484 -1006 487 -1000
rect 491 -1006 494 -1000
rect 498 -1006 501 -1000
rect 505 -1006 508 -1000
rect 512 -1006 515 -1000
rect 519 -1006 522 -1000
rect 526 -1006 532 -1000
rect 533 -1006 536 -1000
rect 540 -1006 543 -1000
rect 547 -1006 550 -1000
rect 554 -1006 557 -1000
rect 561 -1006 564 -1000
rect 568 -1006 571 -1000
rect 575 -1006 578 -1000
rect 582 -1006 585 -1000
rect 589 -1006 592 -1000
rect 596 -1006 599 -1000
rect 603 -1006 606 -1000
rect 610 -1006 616 -1000
rect 617 -1006 620 -1000
rect 624 -1006 630 -1000
rect 631 -1006 637 -1000
rect 638 -1006 641 -1000
rect 645 -1006 648 -1000
rect 652 -1006 655 -1000
rect 659 -1006 662 -1000
rect 666 -1006 669 -1000
rect 673 -1006 676 -1000
rect 680 -1006 683 -1000
rect 687 -1006 690 -1000
rect 694 -1006 697 -1000
rect 701 -1006 704 -1000
rect 708 -1006 711 -1000
rect 715 -1006 721 -1000
rect 722 -1006 725 -1000
rect 729 -1006 732 -1000
rect 736 -1006 739 -1000
rect 743 -1006 746 -1000
rect 750 -1006 753 -1000
rect 757 -1006 760 -1000
rect 764 -1006 767 -1000
rect 771 -1006 777 -1000
rect 778 -1006 784 -1000
rect 785 -1006 788 -1000
rect 792 -1006 798 -1000
rect 799 -1006 802 -1000
rect 806 -1006 809 -1000
rect 813 -1006 819 -1000
rect 820 -1006 823 -1000
rect 827 -1006 833 -1000
rect 834 -1006 837 -1000
rect 841 -1006 844 -1000
rect 848 -1006 851 -1000
rect 855 -1006 858 -1000
rect 862 -1006 865 -1000
rect 869 -1006 872 -1000
rect 876 -1006 879 -1000
rect 883 -1006 886 -1000
rect 890 -1006 893 -1000
rect 897 -1006 900 -1000
rect 904 -1006 907 -1000
rect 911 -1006 914 -1000
rect 918 -1006 921 -1000
rect 925 -1006 928 -1000
rect 932 -1006 938 -1000
rect 939 -1006 942 -1000
rect 946 -1006 949 -1000
rect 953 -1006 959 -1000
rect 960 -1006 963 -1000
rect 967 -1006 970 -1000
rect 974 -1006 977 -1000
rect 981 -1006 984 -1000
rect 988 -1006 991 -1000
rect 995 -1006 998 -1000
rect 1002 -1006 1005 -1000
rect 1009 -1006 1012 -1000
rect 1016 -1006 1022 -1000
rect 1023 -1006 1026 -1000
rect 1030 -1006 1033 -1000
rect 1037 -1006 1043 -1000
rect 1044 -1006 1047 -1000
rect 1051 -1006 1057 -1000
rect 1058 -1006 1064 -1000
rect 1065 -1006 1068 -1000
rect 1072 -1006 1075 -1000
rect 1079 -1006 1082 -1000
rect 1086 -1006 1089 -1000
rect 1093 -1006 1096 -1000
rect 1100 -1006 1103 -1000
rect 1107 -1006 1110 -1000
rect 1114 -1006 1117 -1000
rect 1121 -1006 1127 -1000
rect 1128 -1006 1131 -1000
rect 1135 -1006 1138 -1000
rect 1142 -1006 1145 -1000
rect 1149 -1006 1152 -1000
rect 1156 -1006 1159 -1000
rect 1163 -1006 1166 -1000
rect 1170 -1006 1176 -1000
rect 1177 -1006 1180 -1000
rect 1184 -1006 1187 -1000
rect 1191 -1006 1197 -1000
rect 1198 -1006 1201 -1000
rect 1205 -1006 1208 -1000
rect 1212 -1006 1215 -1000
rect 1219 -1006 1222 -1000
rect 1226 -1006 1229 -1000
rect 1233 -1006 1236 -1000
rect 1240 -1006 1246 -1000
rect 1247 -1006 1250 -1000
rect 1254 -1006 1257 -1000
rect 1261 -1006 1264 -1000
rect 1268 -1006 1274 -1000
rect 1275 -1006 1278 -1000
rect 1282 -1006 1288 -1000
rect 1289 -1006 1292 -1000
rect 1296 -1006 1299 -1000
rect 1303 -1006 1306 -1000
rect 1310 -1006 1316 -1000
rect 1317 -1006 1320 -1000
rect 1324 -1006 1327 -1000
rect 1331 -1006 1334 -1000
rect 1338 -1006 1341 -1000
rect 1345 -1006 1348 -1000
rect 1352 -1006 1355 -1000
rect 1359 -1006 1362 -1000
rect 1366 -1006 1369 -1000
rect 1373 -1006 1376 -1000
rect 1380 -1006 1383 -1000
rect 1387 -1006 1390 -1000
rect 1394 -1006 1400 -1000
rect 1401 -1006 1404 -1000
rect 1408 -1006 1411 -1000
rect 1415 -1006 1418 -1000
rect 1422 -1006 1425 -1000
rect 1429 -1006 1432 -1000
rect 1436 -1006 1439 -1000
rect 1443 -1006 1446 -1000
rect 1450 -1006 1453 -1000
rect 1457 -1006 1460 -1000
rect 1464 -1006 1467 -1000
rect 1471 -1006 1474 -1000
rect 1478 -1006 1481 -1000
rect 1485 -1006 1488 -1000
rect 1492 -1006 1495 -1000
rect 1499 -1006 1502 -1000
rect 1506 -1006 1509 -1000
rect 1513 -1006 1519 -1000
rect 1520 -1006 1523 -1000
rect 1527 -1006 1530 -1000
rect 1534 -1006 1537 -1000
rect 1541 -1006 1544 -1000
rect 1548 -1006 1551 -1000
rect 1555 -1006 1558 -1000
rect 1562 -1006 1565 -1000
rect 1569 -1006 1575 -1000
rect 1576 -1006 1582 -1000
rect 1583 -1006 1586 -1000
rect 1590 -1006 1593 -1000
rect 1597 -1006 1600 -1000
rect 1604 -1006 1607 -1000
rect 1611 -1006 1614 -1000
rect 1618 -1006 1621 -1000
rect 1625 -1006 1628 -1000
rect 1632 -1006 1635 -1000
rect 1639 -1006 1642 -1000
rect 1646 -1006 1649 -1000
rect 1653 -1006 1656 -1000
rect 1660 -1006 1663 -1000
rect 1667 -1006 1670 -1000
rect 1674 -1006 1677 -1000
rect 1681 -1006 1684 -1000
rect 1688 -1006 1691 -1000
rect 1695 -1006 1698 -1000
rect 1702 -1006 1705 -1000
rect 1709 -1006 1712 -1000
rect 1716 -1006 1719 -1000
rect 1723 -1006 1726 -1000
rect 1730 -1006 1733 -1000
rect 1737 -1006 1740 -1000
rect 1744 -1006 1747 -1000
rect 1751 -1006 1754 -1000
rect 1758 -1006 1761 -1000
rect 1765 -1006 1768 -1000
rect 1772 -1006 1775 -1000
rect 1779 -1006 1782 -1000
rect 1786 -1006 1789 -1000
rect 1793 -1006 1796 -1000
rect 1800 -1006 1803 -1000
rect 1807 -1006 1810 -1000
rect 1814 -1006 1817 -1000
rect 1821 -1006 1824 -1000
rect 1828 -1006 1831 -1000
rect 1835 -1006 1838 -1000
rect 1842 -1006 1845 -1000
rect 1849 -1006 1852 -1000
rect 1856 -1006 1859 -1000
rect 1863 -1006 1866 -1000
rect 1870 -1006 1873 -1000
rect 1877 -1006 1880 -1000
rect 1884 -1006 1887 -1000
rect 1891 -1006 1894 -1000
rect 1898 -1006 1901 -1000
rect 1905 -1006 1908 -1000
rect 1912 -1006 1915 -1000
rect 1919 -1006 1922 -1000
rect 1926 -1006 1929 -1000
rect 1933 -1006 1936 -1000
rect 1940 -1006 1943 -1000
rect 1947 -1006 1950 -1000
rect 1954 -1006 1957 -1000
rect 1961 -1006 1964 -1000
rect 1968 -1006 1971 -1000
rect 1975 -1006 1978 -1000
rect 1982 -1006 1985 -1000
rect 1989 -1006 1992 -1000
rect 1996 -1006 1999 -1000
rect 2003 -1006 2006 -1000
rect 2010 -1006 2013 -1000
rect 2017 -1006 2020 -1000
rect 2024 -1006 2027 -1000
rect 2031 -1006 2034 -1000
rect 2038 -1006 2041 -1000
rect 2045 -1006 2048 -1000
rect 2052 -1006 2055 -1000
rect 2059 -1006 2062 -1000
rect 2066 -1006 2069 -1000
rect 2073 -1006 2076 -1000
rect 2080 -1006 2083 -1000
rect 2087 -1006 2090 -1000
rect 2094 -1006 2097 -1000
rect 2101 -1006 2104 -1000
rect 2108 -1006 2111 -1000
rect 2115 -1006 2118 -1000
rect 2122 -1006 2125 -1000
rect 2129 -1006 2132 -1000
rect 2136 -1006 2139 -1000
rect 2143 -1006 2146 -1000
rect 2150 -1006 2153 -1000
rect 2157 -1006 2160 -1000
rect 2164 -1006 2167 -1000
rect 2171 -1006 2174 -1000
rect 2178 -1006 2181 -1000
rect 2185 -1006 2188 -1000
rect 2192 -1006 2195 -1000
rect 2199 -1006 2202 -1000
rect 2206 -1006 2209 -1000
rect 2213 -1006 2216 -1000
rect 2220 -1006 2223 -1000
rect 2227 -1006 2230 -1000
rect 2234 -1006 2237 -1000
rect 2241 -1006 2244 -1000
rect 2248 -1006 2251 -1000
rect 2255 -1006 2258 -1000
rect 2262 -1006 2265 -1000
rect 2269 -1006 2272 -1000
rect 2276 -1006 2279 -1000
rect 2283 -1006 2286 -1000
rect 2290 -1006 2293 -1000
rect 2297 -1006 2300 -1000
rect 2304 -1006 2307 -1000
rect 2311 -1006 2314 -1000
rect 2318 -1006 2321 -1000
rect 2325 -1006 2328 -1000
rect 2332 -1006 2338 -1000
rect 2339 -1006 2345 -1000
rect 2346 -1006 2352 -1000
rect 2353 -1006 2356 -1000
rect 2360 -1006 2363 -1000
rect 2367 -1006 2370 -1000
rect 2374 -1006 2377 -1000
rect 2402 -1006 2405 -1000
rect 2416 -1006 2419 -1000
rect 1 -1173 7 -1167
rect 8 -1173 11 -1167
rect 15 -1173 18 -1167
rect 22 -1173 25 -1167
rect 29 -1173 32 -1167
rect 36 -1173 39 -1167
rect 43 -1173 46 -1167
rect 50 -1173 53 -1167
rect 57 -1173 60 -1167
rect 64 -1173 67 -1167
rect 71 -1173 74 -1167
rect 78 -1173 81 -1167
rect 85 -1173 91 -1167
rect 92 -1173 95 -1167
rect 99 -1173 102 -1167
rect 106 -1173 112 -1167
rect 113 -1173 119 -1167
rect 120 -1173 123 -1167
rect 127 -1173 130 -1167
rect 134 -1173 140 -1167
rect 141 -1173 147 -1167
rect 148 -1173 151 -1167
rect 155 -1173 158 -1167
rect 162 -1173 165 -1167
rect 169 -1173 172 -1167
rect 176 -1173 179 -1167
rect 183 -1173 186 -1167
rect 190 -1173 193 -1167
rect 197 -1173 200 -1167
rect 204 -1173 207 -1167
rect 211 -1173 214 -1167
rect 218 -1173 221 -1167
rect 225 -1173 228 -1167
rect 232 -1173 235 -1167
rect 239 -1173 245 -1167
rect 246 -1173 249 -1167
rect 253 -1173 256 -1167
rect 260 -1173 263 -1167
rect 267 -1173 270 -1167
rect 274 -1173 277 -1167
rect 281 -1173 284 -1167
rect 288 -1173 291 -1167
rect 295 -1173 298 -1167
rect 302 -1173 305 -1167
rect 309 -1173 312 -1167
rect 316 -1173 319 -1167
rect 323 -1173 326 -1167
rect 330 -1173 333 -1167
rect 337 -1173 340 -1167
rect 344 -1173 347 -1167
rect 351 -1173 354 -1167
rect 358 -1173 361 -1167
rect 365 -1173 368 -1167
rect 372 -1173 375 -1167
rect 379 -1173 382 -1167
rect 386 -1173 389 -1167
rect 393 -1173 396 -1167
rect 400 -1173 403 -1167
rect 407 -1173 410 -1167
rect 414 -1173 417 -1167
rect 421 -1173 427 -1167
rect 428 -1173 434 -1167
rect 435 -1173 438 -1167
rect 442 -1173 445 -1167
rect 449 -1173 452 -1167
rect 456 -1173 459 -1167
rect 463 -1173 466 -1167
rect 470 -1173 473 -1167
rect 477 -1173 480 -1167
rect 484 -1173 487 -1167
rect 491 -1173 494 -1167
rect 498 -1173 501 -1167
rect 505 -1173 511 -1167
rect 512 -1173 515 -1167
rect 519 -1173 522 -1167
rect 526 -1173 529 -1167
rect 533 -1173 536 -1167
rect 540 -1173 543 -1167
rect 547 -1173 550 -1167
rect 554 -1173 557 -1167
rect 561 -1173 564 -1167
rect 568 -1173 571 -1167
rect 575 -1173 578 -1167
rect 582 -1173 585 -1167
rect 589 -1173 595 -1167
rect 596 -1173 599 -1167
rect 603 -1173 609 -1167
rect 610 -1173 613 -1167
rect 617 -1173 620 -1167
rect 624 -1173 627 -1167
rect 631 -1173 634 -1167
rect 638 -1173 641 -1167
rect 645 -1173 648 -1167
rect 652 -1173 658 -1167
rect 659 -1173 662 -1167
rect 666 -1173 669 -1167
rect 673 -1173 676 -1167
rect 680 -1173 683 -1167
rect 687 -1173 690 -1167
rect 694 -1173 697 -1167
rect 701 -1173 704 -1167
rect 708 -1173 711 -1167
rect 715 -1173 718 -1167
rect 722 -1173 725 -1167
rect 729 -1173 735 -1167
rect 736 -1173 739 -1167
rect 743 -1173 746 -1167
rect 750 -1173 753 -1167
rect 757 -1173 763 -1167
rect 764 -1173 767 -1167
rect 771 -1173 777 -1167
rect 778 -1173 781 -1167
rect 785 -1173 788 -1167
rect 792 -1173 795 -1167
rect 799 -1173 802 -1167
rect 806 -1173 809 -1167
rect 813 -1173 816 -1167
rect 820 -1173 826 -1167
rect 827 -1173 830 -1167
rect 834 -1173 837 -1167
rect 841 -1173 844 -1167
rect 848 -1173 854 -1167
rect 855 -1173 858 -1167
rect 862 -1173 868 -1167
rect 869 -1173 872 -1167
rect 876 -1173 882 -1167
rect 883 -1173 886 -1167
rect 890 -1173 893 -1167
rect 897 -1173 900 -1167
rect 904 -1173 910 -1167
rect 911 -1173 914 -1167
rect 918 -1173 921 -1167
rect 925 -1173 928 -1167
rect 932 -1173 935 -1167
rect 939 -1173 942 -1167
rect 946 -1173 952 -1167
rect 953 -1173 959 -1167
rect 960 -1173 966 -1167
rect 967 -1173 970 -1167
rect 974 -1173 977 -1167
rect 981 -1173 984 -1167
rect 988 -1173 991 -1167
rect 995 -1173 998 -1167
rect 1002 -1173 1008 -1167
rect 1009 -1173 1012 -1167
rect 1016 -1173 1019 -1167
rect 1023 -1173 1026 -1167
rect 1030 -1173 1033 -1167
rect 1037 -1173 1040 -1167
rect 1044 -1173 1050 -1167
rect 1051 -1173 1054 -1167
rect 1058 -1173 1061 -1167
rect 1065 -1173 1068 -1167
rect 1072 -1173 1075 -1167
rect 1079 -1173 1082 -1167
rect 1086 -1173 1089 -1167
rect 1093 -1173 1096 -1167
rect 1100 -1173 1103 -1167
rect 1107 -1173 1110 -1167
rect 1114 -1173 1117 -1167
rect 1121 -1173 1124 -1167
rect 1128 -1173 1131 -1167
rect 1135 -1173 1138 -1167
rect 1142 -1173 1145 -1167
rect 1149 -1173 1152 -1167
rect 1156 -1173 1162 -1167
rect 1163 -1173 1169 -1167
rect 1170 -1173 1173 -1167
rect 1177 -1173 1183 -1167
rect 1184 -1173 1187 -1167
rect 1191 -1173 1194 -1167
rect 1198 -1173 1204 -1167
rect 1205 -1173 1208 -1167
rect 1212 -1173 1215 -1167
rect 1219 -1173 1225 -1167
rect 1226 -1173 1229 -1167
rect 1233 -1173 1239 -1167
rect 1240 -1173 1243 -1167
rect 1247 -1173 1250 -1167
rect 1254 -1173 1257 -1167
rect 1261 -1173 1264 -1167
rect 1268 -1173 1271 -1167
rect 1275 -1173 1278 -1167
rect 1282 -1173 1285 -1167
rect 1289 -1173 1292 -1167
rect 1296 -1173 1299 -1167
rect 1303 -1173 1309 -1167
rect 1310 -1173 1313 -1167
rect 1317 -1173 1320 -1167
rect 1324 -1173 1327 -1167
rect 1331 -1173 1337 -1167
rect 1338 -1173 1341 -1167
rect 1345 -1173 1348 -1167
rect 1352 -1173 1355 -1167
rect 1359 -1173 1362 -1167
rect 1366 -1173 1369 -1167
rect 1373 -1173 1376 -1167
rect 1380 -1173 1383 -1167
rect 1387 -1173 1390 -1167
rect 1394 -1173 1397 -1167
rect 1401 -1173 1404 -1167
rect 1408 -1173 1411 -1167
rect 1415 -1173 1418 -1167
rect 1422 -1173 1425 -1167
rect 1429 -1173 1432 -1167
rect 1436 -1173 1439 -1167
rect 1443 -1173 1449 -1167
rect 1450 -1173 1453 -1167
rect 1457 -1173 1460 -1167
rect 1464 -1173 1467 -1167
rect 1471 -1173 1474 -1167
rect 1478 -1173 1481 -1167
rect 1485 -1173 1488 -1167
rect 1492 -1173 1495 -1167
rect 1499 -1173 1502 -1167
rect 1506 -1173 1509 -1167
rect 1513 -1173 1516 -1167
rect 1520 -1173 1523 -1167
rect 1527 -1173 1530 -1167
rect 1534 -1173 1537 -1167
rect 1541 -1173 1544 -1167
rect 1548 -1173 1554 -1167
rect 1555 -1173 1558 -1167
rect 1562 -1173 1565 -1167
rect 1569 -1173 1572 -1167
rect 1576 -1173 1579 -1167
rect 1583 -1173 1586 -1167
rect 1590 -1173 1593 -1167
rect 1597 -1173 1600 -1167
rect 1604 -1173 1607 -1167
rect 1611 -1173 1614 -1167
rect 1618 -1173 1621 -1167
rect 1625 -1173 1628 -1167
rect 1632 -1173 1635 -1167
rect 1639 -1173 1642 -1167
rect 1646 -1173 1649 -1167
rect 1653 -1173 1656 -1167
rect 1660 -1173 1663 -1167
rect 1667 -1173 1670 -1167
rect 1674 -1173 1677 -1167
rect 1681 -1173 1684 -1167
rect 1688 -1173 1691 -1167
rect 1695 -1173 1698 -1167
rect 1702 -1173 1705 -1167
rect 1709 -1173 1712 -1167
rect 1716 -1173 1719 -1167
rect 1723 -1173 1726 -1167
rect 1730 -1173 1733 -1167
rect 1737 -1173 1743 -1167
rect 1744 -1173 1747 -1167
rect 1751 -1173 1754 -1167
rect 1758 -1173 1761 -1167
rect 1765 -1173 1768 -1167
rect 1772 -1173 1775 -1167
rect 1779 -1173 1782 -1167
rect 1786 -1173 1789 -1167
rect 1793 -1173 1796 -1167
rect 1800 -1173 1803 -1167
rect 1807 -1173 1810 -1167
rect 1814 -1173 1817 -1167
rect 1821 -1173 1824 -1167
rect 1828 -1173 1831 -1167
rect 1835 -1173 1838 -1167
rect 1842 -1173 1845 -1167
rect 1849 -1173 1852 -1167
rect 1856 -1173 1859 -1167
rect 1863 -1173 1866 -1167
rect 1870 -1173 1873 -1167
rect 1877 -1173 1880 -1167
rect 1884 -1173 1887 -1167
rect 1891 -1173 1894 -1167
rect 1898 -1173 1901 -1167
rect 1905 -1173 1908 -1167
rect 1912 -1173 1915 -1167
rect 1919 -1173 1922 -1167
rect 1926 -1173 1929 -1167
rect 1933 -1173 1936 -1167
rect 1940 -1173 1943 -1167
rect 1947 -1173 1950 -1167
rect 1954 -1173 1957 -1167
rect 1961 -1173 1964 -1167
rect 1968 -1173 1971 -1167
rect 1975 -1173 1978 -1167
rect 1982 -1173 1985 -1167
rect 1989 -1173 1992 -1167
rect 1996 -1173 1999 -1167
rect 2003 -1173 2006 -1167
rect 2010 -1173 2013 -1167
rect 2017 -1173 2020 -1167
rect 2024 -1173 2027 -1167
rect 2031 -1173 2034 -1167
rect 2038 -1173 2041 -1167
rect 2045 -1173 2048 -1167
rect 2052 -1173 2055 -1167
rect 2059 -1173 2062 -1167
rect 2066 -1173 2069 -1167
rect 2073 -1173 2076 -1167
rect 2080 -1173 2083 -1167
rect 2087 -1173 2090 -1167
rect 2094 -1173 2097 -1167
rect 2101 -1173 2104 -1167
rect 2108 -1173 2111 -1167
rect 2115 -1173 2118 -1167
rect 2122 -1173 2125 -1167
rect 2129 -1173 2132 -1167
rect 2136 -1173 2139 -1167
rect 2143 -1173 2146 -1167
rect 2150 -1173 2153 -1167
rect 2157 -1173 2160 -1167
rect 2164 -1173 2167 -1167
rect 2171 -1173 2174 -1167
rect 2178 -1173 2181 -1167
rect 2185 -1173 2188 -1167
rect 2192 -1173 2195 -1167
rect 2199 -1173 2202 -1167
rect 2206 -1173 2209 -1167
rect 2213 -1173 2216 -1167
rect 2220 -1173 2223 -1167
rect 2227 -1173 2230 -1167
rect 2234 -1173 2237 -1167
rect 2241 -1173 2244 -1167
rect 2248 -1173 2251 -1167
rect 2255 -1173 2258 -1167
rect 2262 -1173 2265 -1167
rect 2269 -1173 2272 -1167
rect 2276 -1173 2279 -1167
rect 2283 -1173 2286 -1167
rect 2290 -1173 2293 -1167
rect 2297 -1173 2300 -1167
rect 2304 -1173 2307 -1167
rect 2311 -1173 2314 -1167
rect 2318 -1173 2321 -1167
rect 2325 -1173 2328 -1167
rect 2332 -1173 2335 -1167
rect 2339 -1173 2342 -1167
rect 2346 -1173 2349 -1167
rect 2353 -1173 2356 -1167
rect 2360 -1173 2363 -1167
rect 2367 -1173 2370 -1167
rect 2374 -1173 2377 -1167
rect 2381 -1173 2384 -1167
rect 2388 -1173 2394 -1167
rect 2395 -1173 2401 -1167
rect 2402 -1173 2405 -1167
rect 2423 -1173 2426 -1167
rect 2430 -1173 2433 -1167
rect 2437 -1173 2440 -1167
rect 1 -1356 7 -1350
rect 8 -1356 11 -1350
rect 15 -1356 21 -1350
rect 22 -1356 25 -1350
rect 29 -1356 32 -1350
rect 36 -1356 39 -1350
rect 43 -1356 46 -1350
rect 50 -1356 53 -1350
rect 57 -1356 60 -1350
rect 64 -1356 67 -1350
rect 71 -1356 74 -1350
rect 78 -1356 84 -1350
rect 85 -1356 88 -1350
rect 92 -1356 95 -1350
rect 99 -1356 102 -1350
rect 106 -1356 109 -1350
rect 113 -1356 116 -1350
rect 120 -1356 126 -1350
rect 127 -1356 130 -1350
rect 134 -1356 137 -1350
rect 141 -1356 144 -1350
rect 148 -1356 151 -1350
rect 155 -1356 158 -1350
rect 162 -1356 165 -1350
rect 169 -1356 172 -1350
rect 176 -1356 179 -1350
rect 183 -1356 186 -1350
rect 190 -1356 193 -1350
rect 197 -1356 200 -1350
rect 204 -1356 210 -1350
rect 211 -1356 214 -1350
rect 218 -1356 221 -1350
rect 225 -1356 231 -1350
rect 232 -1356 235 -1350
rect 239 -1356 242 -1350
rect 246 -1356 252 -1350
rect 253 -1356 259 -1350
rect 260 -1356 263 -1350
rect 267 -1356 273 -1350
rect 274 -1356 277 -1350
rect 281 -1356 284 -1350
rect 288 -1356 291 -1350
rect 295 -1356 298 -1350
rect 302 -1356 305 -1350
rect 309 -1356 312 -1350
rect 316 -1356 319 -1350
rect 323 -1356 326 -1350
rect 330 -1356 333 -1350
rect 337 -1356 340 -1350
rect 344 -1356 347 -1350
rect 351 -1356 354 -1350
rect 358 -1356 361 -1350
rect 365 -1356 368 -1350
rect 372 -1356 375 -1350
rect 379 -1356 382 -1350
rect 386 -1356 389 -1350
rect 393 -1356 396 -1350
rect 400 -1356 403 -1350
rect 407 -1356 410 -1350
rect 414 -1356 417 -1350
rect 421 -1356 424 -1350
rect 428 -1356 431 -1350
rect 435 -1356 438 -1350
rect 442 -1356 445 -1350
rect 449 -1356 452 -1350
rect 456 -1356 459 -1350
rect 463 -1356 466 -1350
rect 470 -1356 473 -1350
rect 477 -1356 480 -1350
rect 484 -1356 487 -1350
rect 491 -1356 494 -1350
rect 498 -1356 501 -1350
rect 505 -1356 508 -1350
rect 512 -1356 515 -1350
rect 519 -1356 522 -1350
rect 526 -1356 529 -1350
rect 533 -1356 536 -1350
rect 540 -1356 543 -1350
rect 547 -1356 550 -1350
rect 554 -1356 557 -1350
rect 561 -1356 564 -1350
rect 568 -1356 571 -1350
rect 575 -1356 578 -1350
rect 582 -1356 585 -1350
rect 589 -1356 592 -1350
rect 596 -1356 599 -1350
rect 603 -1356 609 -1350
rect 610 -1356 613 -1350
rect 617 -1356 620 -1350
rect 624 -1356 627 -1350
rect 631 -1356 634 -1350
rect 638 -1356 644 -1350
rect 645 -1356 648 -1350
rect 652 -1356 655 -1350
rect 659 -1356 662 -1350
rect 666 -1356 669 -1350
rect 673 -1356 679 -1350
rect 680 -1356 683 -1350
rect 687 -1356 690 -1350
rect 694 -1356 697 -1350
rect 701 -1356 704 -1350
rect 708 -1356 711 -1350
rect 715 -1356 718 -1350
rect 722 -1356 728 -1350
rect 729 -1356 732 -1350
rect 736 -1356 739 -1350
rect 743 -1356 746 -1350
rect 750 -1356 753 -1350
rect 757 -1356 760 -1350
rect 764 -1356 767 -1350
rect 771 -1356 774 -1350
rect 778 -1356 784 -1350
rect 785 -1356 791 -1350
rect 792 -1356 798 -1350
rect 799 -1356 802 -1350
rect 806 -1356 809 -1350
rect 813 -1356 816 -1350
rect 820 -1356 823 -1350
rect 827 -1356 833 -1350
rect 834 -1356 840 -1350
rect 841 -1356 844 -1350
rect 848 -1356 851 -1350
rect 855 -1356 858 -1350
rect 862 -1356 868 -1350
rect 869 -1356 872 -1350
rect 876 -1356 882 -1350
rect 883 -1356 886 -1350
rect 890 -1356 896 -1350
rect 897 -1356 900 -1350
rect 904 -1356 907 -1350
rect 911 -1356 914 -1350
rect 918 -1356 921 -1350
rect 925 -1356 928 -1350
rect 932 -1356 935 -1350
rect 939 -1356 942 -1350
rect 946 -1356 949 -1350
rect 953 -1356 959 -1350
rect 960 -1356 963 -1350
rect 967 -1356 970 -1350
rect 974 -1356 977 -1350
rect 981 -1356 987 -1350
rect 988 -1356 994 -1350
rect 995 -1356 1001 -1350
rect 1002 -1356 1008 -1350
rect 1009 -1356 1015 -1350
rect 1016 -1356 1019 -1350
rect 1023 -1356 1026 -1350
rect 1030 -1356 1033 -1350
rect 1037 -1356 1043 -1350
rect 1044 -1356 1047 -1350
rect 1051 -1356 1054 -1350
rect 1058 -1356 1061 -1350
rect 1065 -1356 1068 -1350
rect 1072 -1356 1075 -1350
rect 1079 -1356 1082 -1350
rect 1086 -1356 1089 -1350
rect 1093 -1356 1096 -1350
rect 1100 -1356 1106 -1350
rect 1107 -1356 1110 -1350
rect 1114 -1356 1117 -1350
rect 1121 -1356 1124 -1350
rect 1128 -1356 1131 -1350
rect 1135 -1356 1138 -1350
rect 1142 -1356 1145 -1350
rect 1149 -1356 1155 -1350
rect 1156 -1356 1159 -1350
rect 1163 -1356 1166 -1350
rect 1170 -1356 1173 -1350
rect 1177 -1356 1180 -1350
rect 1184 -1356 1187 -1350
rect 1191 -1356 1194 -1350
rect 1198 -1356 1201 -1350
rect 1205 -1356 1208 -1350
rect 1212 -1356 1218 -1350
rect 1219 -1356 1222 -1350
rect 1226 -1356 1229 -1350
rect 1233 -1356 1236 -1350
rect 1240 -1356 1243 -1350
rect 1247 -1356 1250 -1350
rect 1254 -1356 1257 -1350
rect 1261 -1356 1264 -1350
rect 1268 -1356 1271 -1350
rect 1275 -1356 1278 -1350
rect 1282 -1356 1285 -1350
rect 1289 -1356 1292 -1350
rect 1296 -1356 1299 -1350
rect 1303 -1356 1306 -1350
rect 1310 -1356 1313 -1350
rect 1317 -1356 1320 -1350
rect 1324 -1356 1327 -1350
rect 1331 -1356 1334 -1350
rect 1338 -1356 1341 -1350
rect 1345 -1356 1348 -1350
rect 1352 -1356 1355 -1350
rect 1359 -1356 1362 -1350
rect 1366 -1356 1372 -1350
rect 1373 -1356 1376 -1350
rect 1380 -1356 1386 -1350
rect 1387 -1356 1390 -1350
rect 1394 -1356 1397 -1350
rect 1401 -1356 1404 -1350
rect 1408 -1356 1411 -1350
rect 1415 -1356 1421 -1350
rect 1422 -1356 1425 -1350
rect 1429 -1356 1435 -1350
rect 1436 -1356 1439 -1350
rect 1443 -1356 1449 -1350
rect 1450 -1356 1453 -1350
rect 1457 -1356 1460 -1350
rect 1464 -1356 1467 -1350
rect 1471 -1356 1474 -1350
rect 1478 -1356 1481 -1350
rect 1485 -1356 1488 -1350
rect 1492 -1356 1495 -1350
rect 1499 -1356 1502 -1350
rect 1506 -1356 1512 -1350
rect 1513 -1356 1516 -1350
rect 1520 -1356 1523 -1350
rect 1527 -1356 1530 -1350
rect 1534 -1356 1537 -1350
rect 1541 -1356 1544 -1350
rect 1548 -1356 1551 -1350
rect 1555 -1356 1558 -1350
rect 1562 -1356 1565 -1350
rect 1569 -1356 1572 -1350
rect 1576 -1356 1579 -1350
rect 1583 -1356 1586 -1350
rect 1590 -1356 1593 -1350
rect 1597 -1356 1600 -1350
rect 1604 -1356 1607 -1350
rect 1611 -1356 1614 -1350
rect 1618 -1356 1621 -1350
rect 1625 -1356 1628 -1350
rect 1632 -1356 1635 -1350
rect 1639 -1356 1642 -1350
rect 1646 -1356 1649 -1350
rect 1653 -1356 1656 -1350
rect 1660 -1356 1663 -1350
rect 1667 -1356 1670 -1350
rect 1674 -1356 1680 -1350
rect 1681 -1356 1684 -1350
rect 1688 -1356 1691 -1350
rect 1695 -1356 1698 -1350
rect 1702 -1356 1705 -1350
rect 1709 -1356 1712 -1350
rect 1716 -1356 1719 -1350
rect 1723 -1356 1726 -1350
rect 1730 -1356 1733 -1350
rect 1737 -1356 1740 -1350
rect 1744 -1356 1747 -1350
rect 1751 -1356 1754 -1350
rect 1758 -1356 1761 -1350
rect 1765 -1356 1768 -1350
rect 1772 -1356 1775 -1350
rect 1779 -1356 1782 -1350
rect 1786 -1356 1789 -1350
rect 1793 -1356 1796 -1350
rect 1800 -1356 1803 -1350
rect 1807 -1356 1810 -1350
rect 1814 -1356 1817 -1350
rect 1821 -1356 1824 -1350
rect 1828 -1356 1831 -1350
rect 1835 -1356 1838 -1350
rect 1842 -1356 1845 -1350
rect 1849 -1356 1852 -1350
rect 1856 -1356 1859 -1350
rect 1863 -1356 1866 -1350
rect 1870 -1356 1873 -1350
rect 1877 -1356 1880 -1350
rect 1884 -1356 1887 -1350
rect 1891 -1356 1894 -1350
rect 1898 -1356 1901 -1350
rect 1905 -1356 1908 -1350
rect 1912 -1356 1915 -1350
rect 1919 -1356 1922 -1350
rect 1926 -1356 1929 -1350
rect 1933 -1356 1936 -1350
rect 1940 -1356 1943 -1350
rect 1947 -1356 1950 -1350
rect 1954 -1356 1957 -1350
rect 1961 -1356 1964 -1350
rect 1968 -1356 1971 -1350
rect 1975 -1356 1978 -1350
rect 1982 -1356 1985 -1350
rect 1989 -1356 1992 -1350
rect 1996 -1356 1999 -1350
rect 2003 -1356 2006 -1350
rect 2010 -1356 2013 -1350
rect 2017 -1356 2020 -1350
rect 2024 -1356 2027 -1350
rect 2031 -1356 2034 -1350
rect 2038 -1356 2041 -1350
rect 2045 -1356 2048 -1350
rect 2052 -1356 2055 -1350
rect 2059 -1356 2062 -1350
rect 2066 -1356 2069 -1350
rect 2073 -1356 2076 -1350
rect 2080 -1356 2083 -1350
rect 2087 -1356 2090 -1350
rect 2094 -1356 2097 -1350
rect 2101 -1356 2104 -1350
rect 2108 -1356 2111 -1350
rect 2115 -1356 2118 -1350
rect 2122 -1356 2125 -1350
rect 2129 -1356 2132 -1350
rect 2136 -1356 2139 -1350
rect 2143 -1356 2146 -1350
rect 2150 -1356 2153 -1350
rect 2157 -1356 2160 -1350
rect 2164 -1356 2167 -1350
rect 2171 -1356 2174 -1350
rect 2178 -1356 2181 -1350
rect 2185 -1356 2188 -1350
rect 2192 -1356 2195 -1350
rect 2199 -1356 2202 -1350
rect 2206 -1356 2209 -1350
rect 2213 -1356 2216 -1350
rect 2220 -1356 2223 -1350
rect 2227 -1356 2230 -1350
rect 2234 -1356 2237 -1350
rect 2241 -1356 2244 -1350
rect 2248 -1356 2251 -1350
rect 2255 -1356 2258 -1350
rect 2262 -1356 2265 -1350
rect 2269 -1356 2272 -1350
rect 2276 -1356 2279 -1350
rect 2283 -1356 2286 -1350
rect 2290 -1356 2293 -1350
rect 2297 -1356 2300 -1350
rect 2304 -1356 2307 -1350
rect 2311 -1356 2314 -1350
rect 2318 -1356 2321 -1350
rect 2325 -1356 2328 -1350
rect 2332 -1356 2335 -1350
rect 2339 -1356 2345 -1350
rect 2346 -1356 2349 -1350
rect 2353 -1356 2356 -1350
rect 2360 -1356 2363 -1350
rect 2367 -1356 2370 -1350
rect 2374 -1356 2377 -1350
rect 2381 -1356 2384 -1350
rect 2388 -1356 2391 -1350
rect 2395 -1356 2398 -1350
rect 2402 -1356 2405 -1350
rect 2409 -1356 2412 -1350
rect 2416 -1356 2419 -1350
rect 2423 -1356 2426 -1350
rect 2430 -1356 2433 -1350
rect 2437 -1356 2440 -1350
rect 2444 -1356 2447 -1350
rect 2451 -1356 2454 -1350
rect 2458 -1356 2461 -1350
rect 2465 -1356 2468 -1350
rect 2472 -1356 2475 -1350
rect 2479 -1356 2482 -1350
rect 2486 -1356 2489 -1350
rect 2493 -1356 2496 -1350
rect 2500 -1356 2503 -1350
rect 2507 -1356 2510 -1350
rect 2514 -1356 2517 -1350
rect 2521 -1356 2524 -1350
rect 2528 -1356 2531 -1350
rect 2535 -1356 2538 -1350
rect 2542 -1356 2545 -1350
rect 2549 -1356 2552 -1350
rect 2556 -1356 2559 -1350
rect 2563 -1356 2566 -1350
rect 2570 -1356 2573 -1350
rect 2577 -1356 2580 -1350
rect 1 -1533 4 -1527
rect 8 -1533 11 -1527
rect 15 -1533 21 -1527
rect 22 -1533 28 -1527
rect 29 -1533 32 -1527
rect 36 -1533 42 -1527
rect 43 -1533 49 -1527
rect 50 -1533 56 -1527
rect 57 -1533 60 -1527
rect 64 -1533 67 -1527
rect 71 -1533 74 -1527
rect 78 -1533 81 -1527
rect 85 -1533 91 -1527
rect 92 -1533 95 -1527
rect 99 -1533 102 -1527
rect 106 -1533 112 -1527
rect 113 -1533 119 -1527
rect 120 -1533 123 -1527
rect 127 -1533 130 -1527
rect 134 -1533 137 -1527
rect 141 -1533 144 -1527
rect 148 -1533 151 -1527
rect 155 -1533 158 -1527
rect 162 -1533 165 -1527
rect 169 -1533 172 -1527
rect 176 -1533 179 -1527
rect 183 -1533 186 -1527
rect 190 -1533 193 -1527
rect 197 -1533 203 -1527
rect 204 -1533 210 -1527
rect 211 -1533 214 -1527
rect 218 -1533 221 -1527
rect 225 -1533 228 -1527
rect 232 -1533 238 -1527
rect 239 -1533 242 -1527
rect 246 -1533 249 -1527
rect 253 -1533 256 -1527
rect 260 -1533 263 -1527
rect 267 -1533 270 -1527
rect 274 -1533 277 -1527
rect 281 -1533 284 -1527
rect 288 -1533 291 -1527
rect 295 -1533 298 -1527
rect 302 -1533 305 -1527
rect 309 -1533 312 -1527
rect 316 -1533 319 -1527
rect 323 -1533 326 -1527
rect 330 -1533 333 -1527
rect 337 -1533 340 -1527
rect 344 -1533 347 -1527
rect 351 -1533 354 -1527
rect 358 -1533 361 -1527
rect 365 -1533 368 -1527
rect 372 -1533 375 -1527
rect 379 -1533 382 -1527
rect 386 -1533 389 -1527
rect 393 -1533 396 -1527
rect 400 -1533 403 -1527
rect 407 -1533 410 -1527
rect 414 -1533 417 -1527
rect 421 -1533 424 -1527
rect 428 -1533 431 -1527
rect 435 -1533 438 -1527
rect 442 -1533 445 -1527
rect 449 -1533 452 -1527
rect 456 -1533 459 -1527
rect 463 -1533 466 -1527
rect 470 -1533 473 -1527
rect 477 -1533 480 -1527
rect 484 -1533 487 -1527
rect 491 -1533 494 -1527
rect 498 -1533 501 -1527
rect 505 -1533 508 -1527
rect 512 -1533 518 -1527
rect 519 -1533 522 -1527
rect 526 -1533 529 -1527
rect 533 -1533 536 -1527
rect 540 -1533 543 -1527
rect 547 -1533 550 -1527
rect 554 -1533 557 -1527
rect 561 -1533 564 -1527
rect 568 -1533 571 -1527
rect 575 -1533 578 -1527
rect 582 -1533 585 -1527
rect 589 -1533 595 -1527
rect 596 -1533 599 -1527
rect 603 -1533 606 -1527
rect 610 -1533 613 -1527
rect 617 -1533 620 -1527
rect 624 -1533 630 -1527
rect 631 -1533 634 -1527
rect 638 -1533 644 -1527
rect 645 -1533 648 -1527
rect 652 -1533 655 -1527
rect 659 -1533 662 -1527
rect 666 -1533 669 -1527
rect 673 -1533 676 -1527
rect 680 -1533 683 -1527
rect 687 -1533 693 -1527
rect 694 -1533 697 -1527
rect 701 -1533 704 -1527
rect 708 -1533 711 -1527
rect 715 -1533 718 -1527
rect 722 -1533 725 -1527
rect 729 -1533 732 -1527
rect 736 -1533 742 -1527
rect 743 -1533 746 -1527
rect 750 -1533 753 -1527
rect 757 -1533 760 -1527
rect 764 -1533 767 -1527
rect 771 -1533 774 -1527
rect 778 -1533 781 -1527
rect 785 -1533 788 -1527
rect 792 -1533 798 -1527
rect 799 -1533 802 -1527
rect 806 -1533 812 -1527
rect 813 -1533 816 -1527
rect 820 -1533 826 -1527
rect 827 -1533 830 -1527
rect 834 -1533 837 -1527
rect 841 -1533 844 -1527
rect 848 -1533 851 -1527
rect 855 -1533 858 -1527
rect 862 -1533 868 -1527
rect 869 -1533 872 -1527
rect 876 -1533 882 -1527
rect 883 -1533 889 -1527
rect 890 -1533 893 -1527
rect 897 -1533 900 -1527
rect 904 -1533 910 -1527
rect 911 -1533 914 -1527
rect 918 -1533 921 -1527
rect 925 -1533 928 -1527
rect 932 -1533 935 -1527
rect 939 -1533 945 -1527
rect 946 -1533 949 -1527
rect 953 -1533 956 -1527
rect 960 -1533 966 -1527
rect 967 -1533 970 -1527
rect 974 -1533 977 -1527
rect 981 -1533 984 -1527
rect 988 -1533 991 -1527
rect 995 -1533 998 -1527
rect 1002 -1533 1005 -1527
rect 1009 -1533 1012 -1527
rect 1016 -1533 1022 -1527
rect 1023 -1533 1026 -1527
rect 1030 -1533 1033 -1527
rect 1037 -1533 1040 -1527
rect 1044 -1533 1047 -1527
rect 1051 -1533 1054 -1527
rect 1058 -1533 1061 -1527
rect 1065 -1533 1068 -1527
rect 1072 -1533 1075 -1527
rect 1079 -1533 1082 -1527
rect 1086 -1533 1092 -1527
rect 1093 -1533 1096 -1527
rect 1100 -1533 1103 -1527
rect 1107 -1533 1110 -1527
rect 1114 -1533 1117 -1527
rect 1121 -1533 1124 -1527
rect 1128 -1533 1131 -1527
rect 1135 -1533 1138 -1527
rect 1142 -1533 1145 -1527
rect 1149 -1533 1155 -1527
rect 1156 -1533 1162 -1527
rect 1163 -1533 1166 -1527
rect 1170 -1533 1173 -1527
rect 1177 -1533 1180 -1527
rect 1184 -1533 1187 -1527
rect 1191 -1533 1194 -1527
rect 1198 -1533 1201 -1527
rect 1205 -1533 1208 -1527
rect 1212 -1533 1215 -1527
rect 1219 -1533 1222 -1527
rect 1226 -1533 1229 -1527
rect 1233 -1533 1236 -1527
rect 1240 -1533 1243 -1527
rect 1247 -1533 1253 -1527
rect 1254 -1533 1260 -1527
rect 1261 -1533 1267 -1527
rect 1268 -1533 1271 -1527
rect 1275 -1533 1278 -1527
rect 1282 -1533 1288 -1527
rect 1289 -1533 1292 -1527
rect 1296 -1533 1299 -1527
rect 1303 -1533 1306 -1527
rect 1310 -1533 1313 -1527
rect 1317 -1533 1320 -1527
rect 1324 -1533 1327 -1527
rect 1331 -1533 1334 -1527
rect 1338 -1533 1341 -1527
rect 1345 -1533 1351 -1527
rect 1352 -1533 1355 -1527
rect 1359 -1533 1362 -1527
rect 1366 -1533 1369 -1527
rect 1373 -1533 1376 -1527
rect 1380 -1533 1383 -1527
rect 1387 -1533 1390 -1527
rect 1394 -1533 1397 -1527
rect 1401 -1533 1404 -1527
rect 1408 -1533 1411 -1527
rect 1415 -1533 1418 -1527
rect 1422 -1533 1428 -1527
rect 1429 -1533 1432 -1527
rect 1436 -1533 1439 -1527
rect 1443 -1533 1446 -1527
rect 1450 -1533 1453 -1527
rect 1457 -1533 1460 -1527
rect 1464 -1533 1467 -1527
rect 1471 -1533 1474 -1527
rect 1478 -1533 1484 -1527
rect 1485 -1533 1491 -1527
rect 1492 -1533 1495 -1527
rect 1499 -1533 1505 -1527
rect 1506 -1533 1509 -1527
rect 1513 -1533 1516 -1527
rect 1520 -1533 1523 -1527
rect 1527 -1533 1530 -1527
rect 1534 -1533 1537 -1527
rect 1541 -1533 1544 -1527
rect 1548 -1533 1551 -1527
rect 1555 -1533 1558 -1527
rect 1562 -1533 1565 -1527
rect 1569 -1533 1572 -1527
rect 1576 -1533 1579 -1527
rect 1583 -1533 1586 -1527
rect 1590 -1533 1593 -1527
rect 1597 -1533 1600 -1527
rect 1604 -1533 1607 -1527
rect 1611 -1533 1614 -1527
rect 1618 -1533 1621 -1527
rect 1625 -1533 1628 -1527
rect 1632 -1533 1635 -1527
rect 1639 -1533 1642 -1527
rect 1646 -1533 1649 -1527
rect 1653 -1533 1656 -1527
rect 1660 -1533 1663 -1527
rect 1667 -1533 1670 -1527
rect 1674 -1533 1677 -1527
rect 1681 -1533 1684 -1527
rect 1688 -1533 1691 -1527
rect 1695 -1533 1698 -1527
rect 1702 -1533 1705 -1527
rect 1709 -1533 1712 -1527
rect 1716 -1533 1719 -1527
rect 1723 -1533 1726 -1527
rect 1730 -1533 1733 -1527
rect 1737 -1533 1740 -1527
rect 1744 -1533 1747 -1527
rect 1751 -1533 1754 -1527
rect 1758 -1533 1761 -1527
rect 1765 -1533 1768 -1527
rect 1772 -1533 1775 -1527
rect 1779 -1533 1782 -1527
rect 1786 -1533 1789 -1527
rect 1793 -1533 1796 -1527
rect 1800 -1533 1803 -1527
rect 1807 -1533 1810 -1527
rect 1814 -1533 1817 -1527
rect 1821 -1533 1824 -1527
rect 1828 -1533 1831 -1527
rect 1835 -1533 1838 -1527
rect 1842 -1533 1845 -1527
rect 1849 -1533 1852 -1527
rect 1856 -1533 1859 -1527
rect 1863 -1533 1866 -1527
rect 1870 -1533 1873 -1527
rect 1877 -1533 1880 -1527
rect 1884 -1533 1887 -1527
rect 1891 -1533 1894 -1527
rect 1898 -1533 1901 -1527
rect 1905 -1533 1908 -1527
rect 1912 -1533 1915 -1527
rect 1919 -1533 1922 -1527
rect 1926 -1533 1929 -1527
rect 1933 -1533 1936 -1527
rect 1940 -1533 1943 -1527
rect 1947 -1533 1950 -1527
rect 1954 -1533 1957 -1527
rect 1961 -1533 1964 -1527
rect 1968 -1533 1971 -1527
rect 1975 -1533 1978 -1527
rect 1982 -1533 1985 -1527
rect 1989 -1533 1992 -1527
rect 1996 -1533 1999 -1527
rect 2003 -1533 2006 -1527
rect 2010 -1533 2013 -1527
rect 2017 -1533 2020 -1527
rect 2024 -1533 2027 -1527
rect 2031 -1533 2034 -1527
rect 2038 -1533 2041 -1527
rect 2045 -1533 2048 -1527
rect 2052 -1533 2055 -1527
rect 2059 -1533 2062 -1527
rect 2066 -1533 2069 -1527
rect 2073 -1533 2076 -1527
rect 2080 -1533 2083 -1527
rect 2087 -1533 2090 -1527
rect 2094 -1533 2097 -1527
rect 2101 -1533 2104 -1527
rect 2108 -1533 2111 -1527
rect 2115 -1533 2118 -1527
rect 2122 -1533 2125 -1527
rect 2129 -1533 2132 -1527
rect 2136 -1533 2139 -1527
rect 2143 -1533 2146 -1527
rect 2150 -1533 2153 -1527
rect 2157 -1533 2160 -1527
rect 2164 -1533 2167 -1527
rect 2171 -1533 2174 -1527
rect 2178 -1533 2181 -1527
rect 2185 -1533 2188 -1527
rect 2192 -1533 2195 -1527
rect 2199 -1533 2202 -1527
rect 2206 -1533 2209 -1527
rect 2213 -1533 2216 -1527
rect 2220 -1533 2223 -1527
rect 2227 -1533 2230 -1527
rect 2234 -1533 2237 -1527
rect 2241 -1533 2244 -1527
rect 2248 -1533 2251 -1527
rect 2255 -1533 2258 -1527
rect 2262 -1533 2265 -1527
rect 2269 -1533 2272 -1527
rect 2276 -1533 2279 -1527
rect 2283 -1533 2286 -1527
rect 2290 -1533 2293 -1527
rect 2297 -1533 2300 -1527
rect 2304 -1533 2307 -1527
rect 2311 -1533 2314 -1527
rect 2318 -1533 2321 -1527
rect 2325 -1533 2328 -1527
rect 2332 -1533 2335 -1527
rect 2339 -1533 2342 -1527
rect 2346 -1533 2349 -1527
rect 2353 -1533 2356 -1527
rect 2360 -1533 2363 -1527
rect 2367 -1533 2370 -1527
rect 2374 -1533 2377 -1527
rect 2381 -1533 2384 -1527
rect 2388 -1533 2391 -1527
rect 2395 -1533 2398 -1527
rect 2402 -1533 2405 -1527
rect 2409 -1533 2412 -1527
rect 2416 -1533 2419 -1527
rect 2423 -1533 2426 -1527
rect 2430 -1533 2433 -1527
rect 2437 -1533 2440 -1527
rect 2444 -1533 2447 -1527
rect 2451 -1533 2454 -1527
rect 2458 -1533 2461 -1527
rect 2465 -1533 2468 -1527
rect 2472 -1533 2475 -1527
rect 2479 -1533 2482 -1527
rect 2486 -1533 2489 -1527
rect 2493 -1533 2496 -1527
rect 2500 -1533 2503 -1527
rect 2507 -1533 2510 -1527
rect 2514 -1533 2517 -1527
rect 2521 -1533 2524 -1527
rect 2528 -1533 2531 -1527
rect 2535 -1533 2538 -1527
rect 2542 -1533 2545 -1527
rect 2549 -1533 2552 -1527
rect 2556 -1533 2559 -1527
rect 1 -1706 7 -1700
rect 8 -1706 14 -1700
rect 15 -1706 18 -1700
rect 22 -1706 25 -1700
rect 29 -1706 32 -1700
rect 36 -1706 39 -1700
rect 43 -1706 46 -1700
rect 50 -1706 53 -1700
rect 57 -1706 60 -1700
rect 64 -1706 67 -1700
rect 71 -1706 74 -1700
rect 78 -1706 81 -1700
rect 85 -1706 88 -1700
rect 92 -1706 98 -1700
rect 99 -1706 102 -1700
rect 106 -1706 109 -1700
rect 113 -1706 116 -1700
rect 120 -1706 123 -1700
rect 127 -1706 130 -1700
rect 134 -1706 137 -1700
rect 141 -1706 144 -1700
rect 148 -1706 151 -1700
rect 155 -1706 158 -1700
rect 162 -1706 165 -1700
rect 169 -1706 172 -1700
rect 176 -1706 182 -1700
rect 183 -1706 186 -1700
rect 190 -1706 196 -1700
rect 197 -1706 200 -1700
rect 204 -1706 207 -1700
rect 211 -1706 217 -1700
rect 218 -1706 221 -1700
rect 225 -1706 231 -1700
rect 232 -1706 238 -1700
rect 239 -1706 242 -1700
rect 246 -1706 252 -1700
rect 253 -1706 256 -1700
rect 260 -1706 263 -1700
rect 267 -1706 270 -1700
rect 274 -1706 277 -1700
rect 281 -1706 284 -1700
rect 288 -1706 291 -1700
rect 295 -1706 298 -1700
rect 302 -1706 305 -1700
rect 309 -1706 312 -1700
rect 316 -1706 319 -1700
rect 323 -1706 326 -1700
rect 330 -1706 333 -1700
rect 337 -1706 340 -1700
rect 344 -1706 347 -1700
rect 351 -1706 354 -1700
rect 358 -1706 361 -1700
rect 365 -1706 368 -1700
rect 372 -1706 375 -1700
rect 379 -1706 382 -1700
rect 386 -1706 389 -1700
rect 393 -1706 396 -1700
rect 400 -1706 403 -1700
rect 407 -1706 410 -1700
rect 414 -1706 417 -1700
rect 421 -1706 424 -1700
rect 428 -1706 431 -1700
rect 435 -1706 438 -1700
rect 442 -1706 445 -1700
rect 449 -1706 455 -1700
rect 456 -1706 462 -1700
rect 463 -1706 466 -1700
rect 470 -1706 473 -1700
rect 477 -1706 483 -1700
rect 484 -1706 487 -1700
rect 491 -1706 494 -1700
rect 498 -1706 501 -1700
rect 505 -1706 508 -1700
rect 512 -1706 515 -1700
rect 519 -1706 522 -1700
rect 526 -1706 529 -1700
rect 533 -1706 536 -1700
rect 540 -1706 543 -1700
rect 547 -1706 550 -1700
rect 554 -1706 557 -1700
rect 561 -1706 564 -1700
rect 568 -1706 571 -1700
rect 575 -1706 581 -1700
rect 582 -1706 585 -1700
rect 589 -1706 592 -1700
rect 596 -1706 599 -1700
rect 603 -1706 606 -1700
rect 610 -1706 613 -1700
rect 617 -1706 620 -1700
rect 624 -1706 627 -1700
rect 631 -1706 634 -1700
rect 638 -1706 644 -1700
rect 645 -1706 648 -1700
rect 652 -1706 655 -1700
rect 659 -1706 662 -1700
rect 666 -1706 669 -1700
rect 673 -1706 676 -1700
rect 680 -1706 683 -1700
rect 687 -1706 690 -1700
rect 694 -1706 700 -1700
rect 701 -1706 704 -1700
rect 708 -1706 711 -1700
rect 715 -1706 721 -1700
rect 722 -1706 725 -1700
rect 729 -1706 732 -1700
rect 736 -1706 739 -1700
rect 743 -1706 746 -1700
rect 750 -1706 753 -1700
rect 757 -1706 760 -1700
rect 764 -1706 767 -1700
rect 771 -1706 774 -1700
rect 778 -1706 781 -1700
rect 785 -1706 788 -1700
rect 792 -1706 795 -1700
rect 799 -1706 802 -1700
rect 806 -1706 809 -1700
rect 813 -1706 816 -1700
rect 820 -1706 823 -1700
rect 827 -1706 830 -1700
rect 834 -1706 837 -1700
rect 841 -1706 844 -1700
rect 848 -1706 851 -1700
rect 855 -1706 861 -1700
rect 862 -1706 865 -1700
rect 869 -1706 872 -1700
rect 876 -1706 879 -1700
rect 883 -1706 886 -1700
rect 890 -1706 893 -1700
rect 897 -1706 900 -1700
rect 904 -1706 907 -1700
rect 911 -1706 914 -1700
rect 918 -1706 921 -1700
rect 925 -1706 928 -1700
rect 932 -1706 938 -1700
rect 939 -1706 942 -1700
rect 946 -1706 949 -1700
rect 953 -1706 956 -1700
rect 960 -1706 963 -1700
rect 967 -1706 973 -1700
rect 974 -1706 977 -1700
rect 981 -1706 984 -1700
rect 988 -1706 991 -1700
rect 995 -1706 998 -1700
rect 1002 -1706 1005 -1700
rect 1009 -1706 1012 -1700
rect 1016 -1706 1022 -1700
rect 1023 -1706 1026 -1700
rect 1030 -1706 1036 -1700
rect 1037 -1706 1040 -1700
rect 1044 -1706 1047 -1700
rect 1051 -1706 1054 -1700
rect 1058 -1706 1061 -1700
rect 1065 -1706 1068 -1700
rect 1072 -1706 1078 -1700
rect 1079 -1706 1082 -1700
rect 1086 -1706 1089 -1700
rect 1093 -1706 1096 -1700
rect 1100 -1706 1103 -1700
rect 1107 -1706 1113 -1700
rect 1114 -1706 1117 -1700
rect 1121 -1706 1124 -1700
rect 1128 -1706 1131 -1700
rect 1135 -1706 1138 -1700
rect 1142 -1706 1145 -1700
rect 1149 -1706 1155 -1700
rect 1156 -1706 1159 -1700
rect 1163 -1706 1166 -1700
rect 1170 -1706 1173 -1700
rect 1177 -1706 1180 -1700
rect 1184 -1706 1187 -1700
rect 1191 -1706 1194 -1700
rect 1198 -1706 1201 -1700
rect 1205 -1706 1208 -1700
rect 1212 -1706 1215 -1700
rect 1219 -1706 1222 -1700
rect 1226 -1706 1229 -1700
rect 1233 -1706 1236 -1700
rect 1240 -1706 1243 -1700
rect 1247 -1706 1250 -1700
rect 1254 -1706 1257 -1700
rect 1261 -1706 1267 -1700
rect 1268 -1706 1271 -1700
rect 1275 -1706 1281 -1700
rect 1282 -1706 1285 -1700
rect 1289 -1706 1295 -1700
rect 1296 -1706 1299 -1700
rect 1303 -1706 1306 -1700
rect 1310 -1706 1313 -1700
rect 1317 -1706 1320 -1700
rect 1324 -1706 1327 -1700
rect 1331 -1706 1334 -1700
rect 1338 -1706 1341 -1700
rect 1345 -1706 1348 -1700
rect 1352 -1706 1355 -1700
rect 1359 -1706 1365 -1700
rect 1366 -1706 1369 -1700
rect 1373 -1706 1376 -1700
rect 1380 -1706 1383 -1700
rect 1387 -1706 1390 -1700
rect 1394 -1706 1397 -1700
rect 1401 -1706 1404 -1700
rect 1408 -1706 1411 -1700
rect 1415 -1706 1418 -1700
rect 1422 -1706 1425 -1700
rect 1429 -1706 1432 -1700
rect 1436 -1706 1442 -1700
rect 1443 -1706 1446 -1700
rect 1450 -1706 1453 -1700
rect 1457 -1706 1460 -1700
rect 1464 -1706 1470 -1700
rect 1471 -1706 1474 -1700
rect 1478 -1706 1481 -1700
rect 1485 -1706 1488 -1700
rect 1492 -1706 1498 -1700
rect 1499 -1706 1502 -1700
rect 1506 -1706 1512 -1700
rect 1513 -1706 1516 -1700
rect 1520 -1706 1523 -1700
rect 1527 -1706 1533 -1700
rect 1534 -1706 1540 -1700
rect 1541 -1706 1544 -1700
rect 1548 -1706 1551 -1700
rect 1555 -1706 1558 -1700
rect 1562 -1706 1565 -1700
rect 1569 -1706 1572 -1700
rect 1576 -1706 1579 -1700
rect 1583 -1706 1586 -1700
rect 1590 -1706 1593 -1700
rect 1597 -1706 1600 -1700
rect 1604 -1706 1607 -1700
rect 1611 -1706 1614 -1700
rect 1618 -1706 1621 -1700
rect 1625 -1706 1628 -1700
rect 1632 -1706 1635 -1700
rect 1639 -1706 1642 -1700
rect 1646 -1706 1649 -1700
rect 1653 -1706 1656 -1700
rect 1660 -1706 1663 -1700
rect 1667 -1706 1670 -1700
rect 1674 -1706 1677 -1700
rect 1681 -1706 1684 -1700
rect 1688 -1706 1691 -1700
rect 1695 -1706 1698 -1700
rect 1702 -1706 1708 -1700
rect 1709 -1706 1712 -1700
rect 1716 -1706 1719 -1700
rect 1723 -1706 1726 -1700
rect 1730 -1706 1733 -1700
rect 1737 -1706 1740 -1700
rect 1744 -1706 1747 -1700
rect 1751 -1706 1754 -1700
rect 1758 -1706 1761 -1700
rect 1765 -1706 1768 -1700
rect 1772 -1706 1775 -1700
rect 1779 -1706 1782 -1700
rect 1786 -1706 1789 -1700
rect 1793 -1706 1796 -1700
rect 1800 -1706 1803 -1700
rect 1807 -1706 1813 -1700
rect 1814 -1706 1817 -1700
rect 1821 -1706 1824 -1700
rect 1828 -1706 1831 -1700
rect 1835 -1706 1838 -1700
rect 1842 -1706 1845 -1700
rect 1849 -1706 1852 -1700
rect 1856 -1706 1859 -1700
rect 1863 -1706 1866 -1700
rect 1870 -1706 1873 -1700
rect 1877 -1706 1880 -1700
rect 1884 -1706 1887 -1700
rect 1891 -1706 1894 -1700
rect 1898 -1706 1901 -1700
rect 1905 -1706 1908 -1700
rect 1912 -1706 1915 -1700
rect 1919 -1706 1922 -1700
rect 1926 -1706 1929 -1700
rect 1933 -1706 1936 -1700
rect 1940 -1706 1943 -1700
rect 1947 -1706 1950 -1700
rect 1954 -1706 1957 -1700
rect 1961 -1706 1964 -1700
rect 1968 -1706 1971 -1700
rect 1975 -1706 1978 -1700
rect 1982 -1706 1985 -1700
rect 1989 -1706 1992 -1700
rect 1996 -1706 1999 -1700
rect 2003 -1706 2006 -1700
rect 2010 -1706 2013 -1700
rect 2017 -1706 2020 -1700
rect 2024 -1706 2027 -1700
rect 2031 -1706 2034 -1700
rect 2038 -1706 2041 -1700
rect 2045 -1706 2048 -1700
rect 2052 -1706 2055 -1700
rect 2059 -1706 2062 -1700
rect 2066 -1706 2069 -1700
rect 2073 -1706 2076 -1700
rect 2080 -1706 2083 -1700
rect 2087 -1706 2090 -1700
rect 2094 -1706 2097 -1700
rect 2101 -1706 2104 -1700
rect 2108 -1706 2111 -1700
rect 2115 -1706 2118 -1700
rect 2122 -1706 2125 -1700
rect 2129 -1706 2132 -1700
rect 2136 -1706 2139 -1700
rect 2143 -1706 2146 -1700
rect 2150 -1706 2153 -1700
rect 2157 -1706 2160 -1700
rect 2164 -1706 2167 -1700
rect 2171 -1706 2174 -1700
rect 2178 -1706 2181 -1700
rect 2185 -1706 2188 -1700
rect 2192 -1706 2195 -1700
rect 2199 -1706 2202 -1700
rect 2206 -1706 2209 -1700
rect 2213 -1706 2216 -1700
rect 2220 -1706 2223 -1700
rect 2227 -1706 2230 -1700
rect 2234 -1706 2237 -1700
rect 2241 -1706 2244 -1700
rect 2248 -1706 2251 -1700
rect 2255 -1706 2258 -1700
rect 2262 -1706 2265 -1700
rect 2269 -1706 2272 -1700
rect 2276 -1706 2279 -1700
rect 2283 -1706 2286 -1700
rect 2290 -1706 2293 -1700
rect 2297 -1706 2300 -1700
rect 2304 -1706 2307 -1700
rect 2311 -1706 2314 -1700
rect 2318 -1706 2321 -1700
rect 2325 -1706 2328 -1700
rect 2332 -1706 2335 -1700
rect 2339 -1706 2342 -1700
rect 2346 -1706 2349 -1700
rect 2353 -1706 2356 -1700
rect 2360 -1706 2363 -1700
rect 2367 -1706 2370 -1700
rect 2374 -1706 2377 -1700
rect 2381 -1706 2384 -1700
rect 2388 -1706 2391 -1700
rect 2395 -1706 2398 -1700
rect 2402 -1706 2405 -1700
rect 2409 -1706 2412 -1700
rect 2416 -1706 2419 -1700
rect 2423 -1706 2429 -1700
rect 2430 -1706 2436 -1700
rect 2437 -1706 2443 -1700
rect 2444 -1706 2447 -1700
rect 2451 -1706 2454 -1700
rect 2493 -1706 2496 -1700
rect 1 -1857 4 -1851
rect 8 -1857 11 -1851
rect 15 -1857 18 -1851
rect 22 -1857 25 -1851
rect 29 -1857 32 -1851
rect 36 -1857 39 -1851
rect 43 -1857 49 -1851
rect 50 -1857 53 -1851
rect 57 -1857 60 -1851
rect 64 -1857 67 -1851
rect 71 -1857 74 -1851
rect 78 -1857 81 -1851
rect 85 -1857 88 -1851
rect 92 -1857 95 -1851
rect 99 -1857 102 -1851
rect 106 -1857 109 -1851
rect 113 -1857 116 -1851
rect 120 -1857 126 -1851
rect 127 -1857 130 -1851
rect 134 -1857 137 -1851
rect 141 -1857 144 -1851
rect 148 -1857 151 -1851
rect 155 -1857 161 -1851
rect 162 -1857 165 -1851
rect 169 -1857 172 -1851
rect 176 -1857 179 -1851
rect 183 -1857 189 -1851
rect 190 -1857 193 -1851
rect 197 -1857 203 -1851
rect 204 -1857 207 -1851
rect 211 -1857 214 -1851
rect 218 -1857 221 -1851
rect 225 -1857 231 -1851
rect 232 -1857 238 -1851
rect 239 -1857 242 -1851
rect 246 -1857 252 -1851
rect 253 -1857 256 -1851
rect 260 -1857 263 -1851
rect 267 -1857 270 -1851
rect 274 -1857 277 -1851
rect 281 -1857 284 -1851
rect 288 -1857 291 -1851
rect 295 -1857 298 -1851
rect 302 -1857 305 -1851
rect 309 -1857 312 -1851
rect 316 -1857 319 -1851
rect 323 -1857 326 -1851
rect 330 -1857 333 -1851
rect 337 -1857 340 -1851
rect 344 -1857 347 -1851
rect 351 -1857 354 -1851
rect 358 -1857 361 -1851
rect 365 -1857 368 -1851
rect 372 -1857 375 -1851
rect 379 -1857 382 -1851
rect 386 -1857 389 -1851
rect 393 -1857 396 -1851
rect 400 -1857 403 -1851
rect 407 -1857 410 -1851
rect 414 -1857 417 -1851
rect 421 -1857 424 -1851
rect 428 -1857 434 -1851
rect 435 -1857 438 -1851
rect 442 -1857 448 -1851
rect 449 -1857 452 -1851
rect 456 -1857 459 -1851
rect 463 -1857 466 -1851
rect 470 -1857 473 -1851
rect 477 -1857 480 -1851
rect 484 -1857 487 -1851
rect 491 -1857 494 -1851
rect 498 -1857 501 -1851
rect 505 -1857 508 -1851
rect 512 -1857 518 -1851
rect 519 -1857 522 -1851
rect 526 -1857 529 -1851
rect 533 -1857 536 -1851
rect 540 -1857 543 -1851
rect 547 -1857 550 -1851
rect 554 -1857 557 -1851
rect 561 -1857 567 -1851
rect 568 -1857 571 -1851
rect 575 -1857 578 -1851
rect 582 -1857 585 -1851
rect 589 -1857 592 -1851
rect 596 -1857 599 -1851
rect 603 -1857 606 -1851
rect 610 -1857 616 -1851
rect 617 -1857 620 -1851
rect 624 -1857 627 -1851
rect 631 -1857 637 -1851
rect 638 -1857 641 -1851
rect 645 -1857 651 -1851
rect 652 -1857 655 -1851
rect 659 -1857 662 -1851
rect 666 -1857 669 -1851
rect 673 -1857 676 -1851
rect 680 -1857 683 -1851
rect 687 -1857 690 -1851
rect 694 -1857 697 -1851
rect 701 -1857 704 -1851
rect 708 -1857 711 -1851
rect 715 -1857 718 -1851
rect 722 -1857 728 -1851
rect 729 -1857 735 -1851
rect 736 -1857 742 -1851
rect 743 -1857 746 -1851
rect 750 -1857 753 -1851
rect 757 -1857 760 -1851
rect 764 -1857 767 -1851
rect 771 -1857 774 -1851
rect 778 -1857 781 -1851
rect 785 -1857 788 -1851
rect 792 -1857 795 -1851
rect 799 -1857 805 -1851
rect 806 -1857 809 -1851
rect 813 -1857 816 -1851
rect 820 -1857 823 -1851
rect 827 -1857 830 -1851
rect 834 -1857 837 -1851
rect 841 -1857 844 -1851
rect 848 -1857 854 -1851
rect 855 -1857 858 -1851
rect 862 -1857 865 -1851
rect 869 -1857 872 -1851
rect 876 -1857 879 -1851
rect 883 -1857 886 -1851
rect 890 -1857 896 -1851
rect 897 -1857 900 -1851
rect 904 -1857 910 -1851
rect 911 -1857 914 -1851
rect 918 -1857 921 -1851
rect 925 -1857 928 -1851
rect 932 -1857 935 -1851
rect 939 -1857 945 -1851
rect 946 -1857 949 -1851
rect 953 -1857 959 -1851
rect 960 -1857 963 -1851
rect 967 -1857 970 -1851
rect 974 -1857 977 -1851
rect 981 -1857 984 -1851
rect 988 -1857 991 -1851
rect 995 -1857 998 -1851
rect 1002 -1857 1005 -1851
rect 1009 -1857 1012 -1851
rect 1016 -1857 1019 -1851
rect 1023 -1857 1026 -1851
rect 1030 -1857 1033 -1851
rect 1037 -1857 1040 -1851
rect 1044 -1857 1047 -1851
rect 1051 -1857 1054 -1851
rect 1058 -1857 1061 -1851
rect 1065 -1857 1068 -1851
rect 1072 -1857 1075 -1851
rect 1079 -1857 1082 -1851
rect 1086 -1857 1089 -1851
rect 1093 -1857 1096 -1851
rect 1100 -1857 1103 -1851
rect 1107 -1857 1110 -1851
rect 1114 -1857 1117 -1851
rect 1121 -1857 1124 -1851
rect 1128 -1857 1131 -1851
rect 1135 -1857 1141 -1851
rect 1142 -1857 1145 -1851
rect 1149 -1857 1152 -1851
rect 1156 -1857 1159 -1851
rect 1163 -1857 1166 -1851
rect 1170 -1857 1173 -1851
rect 1177 -1857 1183 -1851
rect 1184 -1857 1187 -1851
rect 1191 -1857 1194 -1851
rect 1198 -1857 1201 -1851
rect 1205 -1857 1211 -1851
rect 1212 -1857 1215 -1851
rect 1219 -1857 1222 -1851
rect 1226 -1857 1229 -1851
rect 1233 -1857 1236 -1851
rect 1240 -1857 1243 -1851
rect 1247 -1857 1250 -1851
rect 1254 -1857 1257 -1851
rect 1261 -1857 1264 -1851
rect 1268 -1857 1271 -1851
rect 1275 -1857 1281 -1851
rect 1282 -1857 1285 -1851
rect 1289 -1857 1295 -1851
rect 1296 -1857 1299 -1851
rect 1303 -1857 1309 -1851
rect 1310 -1857 1313 -1851
rect 1317 -1857 1320 -1851
rect 1324 -1857 1327 -1851
rect 1331 -1857 1334 -1851
rect 1338 -1857 1341 -1851
rect 1345 -1857 1348 -1851
rect 1352 -1857 1355 -1851
rect 1359 -1857 1362 -1851
rect 1366 -1857 1369 -1851
rect 1373 -1857 1376 -1851
rect 1380 -1857 1383 -1851
rect 1387 -1857 1390 -1851
rect 1394 -1857 1397 -1851
rect 1401 -1857 1404 -1851
rect 1408 -1857 1411 -1851
rect 1415 -1857 1418 -1851
rect 1422 -1857 1425 -1851
rect 1429 -1857 1432 -1851
rect 1436 -1857 1442 -1851
rect 1443 -1857 1446 -1851
rect 1450 -1857 1453 -1851
rect 1457 -1857 1460 -1851
rect 1464 -1857 1470 -1851
rect 1471 -1857 1474 -1851
rect 1478 -1857 1481 -1851
rect 1485 -1857 1488 -1851
rect 1492 -1857 1495 -1851
rect 1499 -1857 1502 -1851
rect 1506 -1857 1512 -1851
rect 1513 -1857 1516 -1851
rect 1520 -1857 1523 -1851
rect 1527 -1857 1530 -1851
rect 1534 -1857 1537 -1851
rect 1541 -1857 1544 -1851
rect 1548 -1857 1551 -1851
rect 1555 -1857 1558 -1851
rect 1562 -1857 1565 -1851
rect 1569 -1857 1572 -1851
rect 1576 -1857 1579 -1851
rect 1583 -1857 1586 -1851
rect 1590 -1857 1593 -1851
rect 1597 -1857 1600 -1851
rect 1604 -1857 1607 -1851
rect 1611 -1857 1614 -1851
rect 1618 -1857 1621 -1851
rect 1625 -1857 1631 -1851
rect 1632 -1857 1635 -1851
rect 1639 -1857 1642 -1851
rect 1646 -1857 1649 -1851
rect 1653 -1857 1656 -1851
rect 1660 -1857 1666 -1851
rect 1667 -1857 1670 -1851
rect 1674 -1857 1677 -1851
rect 1681 -1857 1684 -1851
rect 1688 -1857 1691 -1851
rect 1695 -1857 1698 -1851
rect 1702 -1857 1705 -1851
rect 1709 -1857 1712 -1851
rect 1716 -1857 1719 -1851
rect 1723 -1857 1726 -1851
rect 1730 -1857 1733 -1851
rect 1737 -1857 1740 -1851
rect 1744 -1857 1747 -1851
rect 1751 -1857 1754 -1851
rect 1758 -1857 1761 -1851
rect 1765 -1857 1768 -1851
rect 1772 -1857 1775 -1851
rect 1779 -1857 1782 -1851
rect 1786 -1857 1789 -1851
rect 1793 -1857 1796 -1851
rect 1800 -1857 1803 -1851
rect 1807 -1857 1810 -1851
rect 1814 -1857 1817 -1851
rect 1821 -1857 1824 -1851
rect 1828 -1857 1831 -1851
rect 1835 -1857 1838 -1851
rect 1842 -1857 1845 -1851
rect 1849 -1857 1855 -1851
rect 1856 -1857 1859 -1851
rect 1863 -1857 1869 -1851
rect 1870 -1857 1873 -1851
rect 1877 -1857 1880 -1851
rect 1884 -1857 1887 -1851
rect 1891 -1857 1894 -1851
rect 1898 -1857 1901 -1851
rect 1905 -1857 1908 -1851
rect 1912 -1857 1915 -1851
rect 1919 -1857 1922 -1851
rect 1926 -1857 1929 -1851
rect 1933 -1857 1936 -1851
rect 1940 -1857 1943 -1851
rect 1947 -1857 1950 -1851
rect 1954 -1857 1957 -1851
rect 1961 -1857 1964 -1851
rect 1968 -1857 1971 -1851
rect 1975 -1857 1978 -1851
rect 1982 -1857 1985 -1851
rect 1989 -1857 1992 -1851
rect 1996 -1857 1999 -1851
rect 2003 -1857 2006 -1851
rect 2010 -1857 2013 -1851
rect 2017 -1857 2020 -1851
rect 2024 -1857 2027 -1851
rect 2031 -1857 2034 -1851
rect 2038 -1857 2041 -1851
rect 2045 -1857 2048 -1851
rect 2052 -1857 2055 -1851
rect 2059 -1857 2062 -1851
rect 2066 -1857 2069 -1851
rect 2073 -1857 2076 -1851
rect 2080 -1857 2083 -1851
rect 2087 -1857 2090 -1851
rect 2094 -1857 2097 -1851
rect 2101 -1857 2104 -1851
rect 2108 -1857 2111 -1851
rect 2115 -1857 2118 -1851
rect 2122 -1857 2125 -1851
rect 2129 -1857 2132 -1851
rect 2136 -1857 2139 -1851
rect 2143 -1857 2146 -1851
rect 2150 -1857 2153 -1851
rect 2157 -1857 2160 -1851
rect 2164 -1857 2167 -1851
rect 2171 -1857 2174 -1851
rect 2178 -1857 2181 -1851
rect 2185 -1857 2188 -1851
rect 2192 -1857 2195 -1851
rect 2199 -1857 2202 -1851
rect 2206 -1857 2209 -1851
rect 2213 -1857 2216 -1851
rect 2220 -1857 2223 -1851
rect 2227 -1857 2230 -1851
rect 2234 -1857 2237 -1851
rect 2241 -1857 2244 -1851
rect 2248 -1857 2251 -1851
rect 2255 -1857 2258 -1851
rect 2262 -1857 2265 -1851
rect 2269 -1857 2272 -1851
rect 2276 -1857 2279 -1851
rect 2283 -1857 2286 -1851
rect 2290 -1857 2293 -1851
rect 2297 -1857 2300 -1851
rect 2304 -1857 2307 -1851
rect 2311 -1857 2314 -1851
rect 2318 -1857 2321 -1851
rect 2325 -1857 2328 -1851
rect 2332 -1857 2335 -1851
rect 2339 -1857 2342 -1851
rect 2346 -1857 2349 -1851
rect 2353 -1857 2356 -1851
rect 2360 -1857 2363 -1851
rect 2367 -1857 2370 -1851
rect 2374 -1857 2377 -1851
rect 2381 -1857 2384 -1851
rect 2388 -1857 2391 -1851
rect 2395 -1857 2398 -1851
rect 2402 -1857 2405 -1851
rect 2409 -1857 2412 -1851
rect 2416 -1857 2419 -1851
rect 2423 -1857 2426 -1851
rect 2430 -1857 2433 -1851
rect 2437 -1857 2440 -1851
rect 2444 -1857 2447 -1851
rect 2451 -1857 2454 -1851
rect 2458 -1857 2461 -1851
rect 2465 -1857 2471 -1851
rect 2472 -1857 2478 -1851
rect 1 -2032 4 -2026
rect 8 -2032 11 -2026
rect 15 -2032 18 -2026
rect 22 -2032 25 -2026
rect 29 -2032 32 -2026
rect 36 -2032 39 -2026
rect 43 -2032 46 -2026
rect 50 -2032 56 -2026
rect 57 -2032 60 -2026
rect 64 -2032 67 -2026
rect 71 -2032 74 -2026
rect 78 -2032 81 -2026
rect 85 -2032 91 -2026
rect 92 -2032 95 -2026
rect 99 -2032 105 -2026
rect 106 -2032 109 -2026
rect 113 -2032 116 -2026
rect 120 -2032 123 -2026
rect 127 -2032 133 -2026
rect 134 -2032 137 -2026
rect 141 -2032 144 -2026
rect 148 -2032 151 -2026
rect 155 -2032 161 -2026
rect 162 -2032 165 -2026
rect 169 -2032 175 -2026
rect 176 -2032 179 -2026
rect 183 -2032 186 -2026
rect 190 -2032 196 -2026
rect 197 -2032 200 -2026
rect 204 -2032 207 -2026
rect 211 -2032 217 -2026
rect 218 -2032 221 -2026
rect 225 -2032 228 -2026
rect 232 -2032 235 -2026
rect 239 -2032 242 -2026
rect 246 -2032 249 -2026
rect 253 -2032 256 -2026
rect 260 -2032 263 -2026
rect 267 -2032 270 -2026
rect 274 -2032 277 -2026
rect 281 -2032 284 -2026
rect 288 -2032 291 -2026
rect 295 -2032 298 -2026
rect 302 -2032 305 -2026
rect 309 -2032 312 -2026
rect 316 -2032 319 -2026
rect 323 -2032 326 -2026
rect 330 -2032 333 -2026
rect 337 -2032 340 -2026
rect 344 -2032 347 -2026
rect 351 -2032 354 -2026
rect 358 -2032 361 -2026
rect 365 -2032 368 -2026
rect 372 -2032 375 -2026
rect 379 -2032 382 -2026
rect 386 -2032 389 -2026
rect 393 -2032 396 -2026
rect 400 -2032 403 -2026
rect 407 -2032 410 -2026
rect 414 -2032 417 -2026
rect 421 -2032 424 -2026
rect 428 -2032 431 -2026
rect 435 -2032 438 -2026
rect 442 -2032 445 -2026
rect 449 -2032 452 -2026
rect 456 -2032 459 -2026
rect 463 -2032 466 -2026
rect 470 -2032 473 -2026
rect 477 -2032 480 -2026
rect 484 -2032 487 -2026
rect 491 -2032 494 -2026
rect 498 -2032 501 -2026
rect 505 -2032 508 -2026
rect 512 -2032 515 -2026
rect 519 -2032 522 -2026
rect 526 -2032 529 -2026
rect 533 -2032 536 -2026
rect 540 -2032 546 -2026
rect 547 -2032 550 -2026
rect 554 -2032 557 -2026
rect 561 -2032 564 -2026
rect 568 -2032 571 -2026
rect 575 -2032 578 -2026
rect 582 -2032 588 -2026
rect 589 -2032 592 -2026
rect 596 -2032 599 -2026
rect 603 -2032 606 -2026
rect 610 -2032 613 -2026
rect 617 -2032 620 -2026
rect 624 -2032 627 -2026
rect 631 -2032 637 -2026
rect 638 -2032 641 -2026
rect 645 -2032 648 -2026
rect 652 -2032 655 -2026
rect 659 -2032 662 -2026
rect 666 -2032 669 -2026
rect 673 -2032 676 -2026
rect 680 -2032 683 -2026
rect 687 -2032 690 -2026
rect 694 -2032 697 -2026
rect 701 -2032 704 -2026
rect 708 -2032 711 -2026
rect 715 -2032 718 -2026
rect 722 -2032 725 -2026
rect 729 -2032 732 -2026
rect 736 -2032 742 -2026
rect 743 -2032 746 -2026
rect 750 -2032 753 -2026
rect 757 -2032 760 -2026
rect 764 -2032 767 -2026
rect 771 -2032 774 -2026
rect 778 -2032 784 -2026
rect 785 -2032 788 -2026
rect 792 -2032 795 -2026
rect 799 -2032 805 -2026
rect 806 -2032 809 -2026
rect 813 -2032 816 -2026
rect 820 -2032 823 -2026
rect 827 -2032 833 -2026
rect 834 -2032 837 -2026
rect 841 -2032 844 -2026
rect 848 -2032 851 -2026
rect 855 -2032 858 -2026
rect 862 -2032 865 -2026
rect 869 -2032 872 -2026
rect 876 -2032 879 -2026
rect 883 -2032 886 -2026
rect 890 -2032 893 -2026
rect 897 -2032 900 -2026
rect 904 -2032 907 -2026
rect 911 -2032 914 -2026
rect 918 -2032 924 -2026
rect 925 -2032 928 -2026
rect 932 -2032 935 -2026
rect 939 -2032 942 -2026
rect 946 -2032 949 -2026
rect 953 -2032 959 -2026
rect 960 -2032 963 -2026
rect 967 -2032 970 -2026
rect 974 -2032 980 -2026
rect 981 -2032 984 -2026
rect 988 -2032 991 -2026
rect 995 -2032 998 -2026
rect 1002 -2032 1005 -2026
rect 1009 -2032 1012 -2026
rect 1016 -2032 1019 -2026
rect 1023 -2032 1026 -2026
rect 1030 -2032 1033 -2026
rect 1037 -2032 1040 -2026
rect 1044 -2032 1047 -2026
rect 1051 -2032 1054 -2026
rect 1058 -2032 1064 -2026
rect 1065 -2032 1068 -2026
rect 1072 -2032 1075 -2026
rect 1079 -2032 1082 -2026
rect 1086 -2032 1089 -2026
rect 1093 -2032 1096 -2026
rect 1100 -2032 1103 -2026
rect 1107 -2032 1113 -2026
rect 1114 -2032 1117 -2026
rect 1121 -2032 1127 -2026
rect 1128 -2032 1131 -2026
rect 1135 -2032 1138 -2026
rect 1142 -2032 1145 -2026
rect 1149 -2032 1155 -2026
rect 1156 -2032 1159 -2026
rect 1163 -2032 1169 -2026
rect 1170 -2032 1173 -2026
rect 1177 -2032 1180 -2026
rect 1184 -2032 1190 -2026
rect 1191 -2032 1194 -2026
rect 1198 -2032 1201 -2026
rect 1205 -2032 1208 -2026
rect 1212 -2032 1215 -2026
rect 1219 -2032 1222 -2026
rect 1226 -2032 1232 -2026
rect 1233 -2032 1236 -2026
rect 1240 -2032 1243 -2026
rect 1247 -2032 1250 -2026
rect 1254 -2032 1257 -2026
rect 1261 -2032 1264 -2026
rect 1268 -2032 1271 -2026
rect 1275 -2032 1278 -2026
rect 1282 -2032 1285 -2026
rect 1289 -2032 1292 -2026
rect 1296 -2032 1302 -2026
rect 1303 -2032 1306 -2026
rect 1310 -2032 1313 -2026
rect 1317 -2032 1320 -2026
rect 1324 -2032 1327 -2026
rect 1331 -2032 1334 -2026
rect 1338 -2032 1341 -2026
rect 1345 -2032 1348 -2026
rect 1352 -2032 1355 -2026
rect 1359 -2032 1365 -2026
rect 1366 -2032 1369 -2026
rect 1373 -2032 1376 -2026
rect 1380 -2032 1383 -2026
rect 1387 -2032 1390 -2026
rect 1394 -2032 1397 -2026
rect 1401 -2032 1404 -2026
rect 1408 -2032 1411 -2026
rect 1415 -2032 1418 -2026
rect 1422 -2032 1425 -2026
rect 1429 -2032 1432 -2026
rect 1436 -2032 1442 -2026
rect 1443 -2032 1446 -2026
rect 1450 -2032 1453 -2026
rect 1457 -2032 1460 -2026
rect 1464 -2032 1467 -2026
rect 1471 -2032 1477 -2026
rect 1478 -2032 1481 -2026
rect 1485 -2032 1491 -2026
rect 1492 -2032 1498 -2026
rect 1499 -2032 1502 -2026
rect 1506 -2032 1509 -2026
rect 1513 -2032 1516 -2026
rect 1520 -2032 1526 -2026
rect 1527 -2032 1530 -2026
rect 1534 -2032 1540 -2026
rect 1541 -2032 1544 -2026
rect 1548 -2032 1554 -2026
rect 1555 -2032 1558 -2026
rect 1562 -2032 1565 -2026
rect 1569 -2032 1572 -2026
rect 1576 -2032 1579 -2026
rect 1583 -2032 1586 -2026
rect 1590 -2032 1593 -2026
rect 1597 -2032 1600 -2026
rect 1604 -2032 1607 -2026
rect 1611 -2032 1614 -2026
rect 1618 -2032 1624 -2026
rect 1625 -2032 1628 -2026
rect 1632 -2032 1638 -2026
rect 1639 -2032 1642 -2026
rect 1646 -2032 1649 -2026
rect 1653 -2032 1656 -2026
rect 1660 -2032 1666 -2026
rect 1667 -2032 1670 -2026
rect 1674 -2032 1677 -2026
rect 1681 -2032 1684 -2026
rect 1688 -2032 1691 -2026
rect 1695 -2032 1698 -2026
rect 1702 -2032 1705 -2026
rect 1709 -2032 1712 -2026
rect 1716 -2032 1719 -2026
rect 1723 -2032 1726 -2026
rect 1730 -2032 1736 -2026
rect 1737 -2032 1740 -2026
rect 1744 -2032 1747 -2026
rect 1751 -2032 1754 -2026
rect 1758 -2032 1761 -2026
rect 1765 -2032 1768 -2026
rect 1772 -2032 1775 -2026
rect 1779 -2032 1782 -2026
rect 1786 -2032 1789 -2026
rect 1793 -2032 1796 -2026
rect 1800 -2032 1803 -2026
rect 1807 -2032 1810 -2026
rect 1814 -2032 1817 -2026
rect 1821 -2032 1824 -2026
rect 1828 -2032 1831 -2026
rect 1835 -2032 1838 -2026
rect 1842 -2032 1845 -2026
rect 1849 -2032 1852 -2026
rect 1856 -2032 1859 -2026
rect 1863 -2032 1866 -2026
rect 1870 -2032 1873 -2026
rect 1877 -2032 1880 -2026
rect 1884 -2032 1887 -2026
rect 1891 -2032 1894 -2026
rect 1898 -2032 1901 -2026
rect 1905 -2032 1908 -2026
rect 1912 -2032 1915 -2026
rect 1919 -2032 1922 -2026
rect 1926 -2032 1929 -2026
rect 1933 -2032 1936 -2026
rect 1940 -2032 1943 -2026
rect 1947 -2032 1950 -2026
rect 1954 -2032 1957 -2026
rect 1961 -2032 1964 -2026
rect 1968 -2032 1971 -2026
rect 1975 -2032 1978 -2026
rect 1982 -2032 1985 -2026
rect 1989 -2032 1992 -2026
rect 1996 -2032 1999 -2026
rect 2003 -2032 2006 -2026
rect 2010 -2032 2013 -2026
rect 2017 -2032 2020 -2026
rect 2024 -2032 2027 -2026
rect 2031 -2032 2034 -2026
rect 2038 -2032 2041 -2026
rect 2045 -2032 2048 -2026
rect 2052 -2032 2055 -2026
rect 2059 -2032 2062 -2026
rect 2066 -2032 2069 -2026
rect 2073 -2032 2076 -2026
rect 2080 -2032 2083 -2026
rect 2087 -2032 2090 -2026
rect 2094 -2032 2097 -2026
rect 2101 -2032 2104 -2026
rect 2108 -2032 2111 -2026
rect 2115 -2032 2118 -2026
rect 2122 -2032 2125 -2026
rect 2129 -2032 2132 -2026
rect 2136 -2032 2139 -2026
rect 2143 -2032 2146 -2026
rect 2150 -2032 2153 -2026
rect 2157 -2032 2160 -2026
rect 2164 -2032 2167 -2026
rect 2171 -2032 2174 -2026
rect 2178 -2032 2181 -2026
rect 2185 -2032 2188 -2026
rect 2192 -2032 2195 -2026
rect 2199 -2032 2202 -2026
rect 2206 -2032 2209 -2026
rect 2213 -2032 2216 -2026
rect 2220 -2032 2223 -2026
rect 2227 -2032 2230 -2026
rect 2234 -2032 2237 -2026
rect 2241 -2032 2244 -2026
rect 2248 -2032 2251 -2026
rect 2255 -2032 2258 -2026
rect 2262 -2032 2265 -2026
rect 2269 -2032 2272 -2026
rect 2276 -2032 2279 -2026
rect 2283 -2032 2286 -2026
rect 2290 -2032 2293 -2026
rect 2297 -2032 2300 -2026
rect 2304 -2032 2307 -2026
rect 2311 -2032 2314 -2026
rect 2318 -2032 2321 -2026
rect 2325 -2032 2328 -2026
rect 2332 -2032 2335 -2026
rect 2339 -2032 2342 -2026
rect 2346 -2032 2349 -2026
rect 2353 -2032 2356 -2026
rect 2360 -2032 2363 -2026
rect 2367 -2032 2370 -2026
rect 2374 -2032 2377 -2026
rect 2381 -2032 2384 -2026
rect 2388 -2032 2391 -2026
rect 2395 -2032 2398 -2026
rect 2402 -2032 2405 -2026
rect 2409 -2032 2412 -2026
rect 2416 -2032 2422 -2026
rect 2423 -2032 2426 -2026
rect 1 -2183 7 -2177
rect 8 -2183 11 -2177
rect 15 -2183 18 -2177
rect 22 -2183 25 -2177
rect 29 -2183 32 -2177
rect 36 -2183 42 -2177
rect 43 -2183 46 -2177
rect 50 -2183 56 -2177
rect 57 -2183 60 -2177
rect 64 -2183 67 -2177
rect 71 -2183 74 -2177
rect 78 -2183 81 -2177
rect 85 -2183 88 -2177
rect 92 -2183 98 -2177
rect 99 -2183 102 -2177
rect 106 -2183 109 -2177
rect 113 -2183 116 -2177
rect 120 -2183 126 -2177
rect 127 -2183 133 -2177
rect 134 -2183 140 -2177
rect 141 -2183 144 -2177
rect 148 -2183 151 -2177
rect 155 -2183 158 -2177
rect 162 -2183 165 -2177
rect 169 -2183 172 -2177
rect 176 -2183 179 -2177
rect 183 -2183 186 -2177
rect 190 -2183 193 -2177
rect 197 -2183 200 -2177
rect 204 -2183 207 -2177
rect 211 -2183 214 -2177
rect 218 -2183 221 -2177
rect 225 -2183 228 -2177
rect 232 -2183 238 -2177
rect 239 -2183 245 -2177
rect 246 -2183 249 -2177
rect 253 -2183 259 -2177
rect 260 -2183 263 -2177
rect 267 -2183 270 -2177
rect 274 -2183 277 -2177
rect 281 -2183 284 -2177
rect 288 -2183 291 -2177
rect 295 -2183 298 -2177
rect 302 -2183 305 -2177
rect 309 -2183 312 -2177
rect 316 -2183 319 -2177
rect 323 -2183 326 -2177
rect 330 -2183 333 -2177
rect 337 -2183 340 -2177
rect 344 -2183 347 -2177
rect 351 -2183 354 -2177
rect 358 -2183 361 -2177
rect 365 -2183 368 -2177
rect 372 -2183 375 -2177
rect 379 -2183 382 -2177
rect 386 -2183 389 -2177
rect 393 -2183 396 -2177
rect 400 -2183 406 -2177
rect 407 -2183 410 -2177
rect 414 -2183 417 -2177
rect 421 -2183 424 -2177
rect 428 -2183 431 -2177
rect 435 -2183 438 -2177
rect 442 -2183 445 -2177
rect 449 -2183 452 -2177
rect 456 -2183 459 -2177
rect 463 -2183 466 -2177
rect 470 -2183 473 -2177
rect 477 -2183 480 -2177
rect 484 -2183 487 -2177
rect 491 -2183 497 -2177
rect 498 -2183 501 -2177
rect 505 -2183 508 -2177
rect 512 -2183 518 -2177
rect 519 -2183 522 -2177
rect 526 -2183 529 -2177
rect 533 -2183 536 -2177
rect 540 -2183 543 -2177
rect 547 -2183 550 -2177
rect 554 -2183 557 -2177
rect 561 -2183 564 -2177
rect 568 -2183 571 -2177
rect 575 -2183 578 -2177
rect 582 -2183 585 -2177
rect 589 -2183 592 -2177
rect 596 -2183 599 -2177
rect 603 -2183 606 -2177
rect 610 -2183 613 -2177
rect 617 -2183 620 -2177
rect 624 -2183 627 -2177
rect 631 -2183 634 -2177
rect 638 -2183 641 -2177
rect 645 -2183 648 -2177
rect 652 -2183 658 -2177
rect 659 -2183 662 -2177
rect 666 -2183 672 -2177
rect 673 -2183 676 -2177
rect 680 -2183 683 -2177
rect 687 -2183 690 -2177
rect 694 -2183 697 -2177
rect 701 -2183 704 -2177
rect 708 -2183 711 -2177
rect 715 -2183 718 -2177
rect 722 -2183 725 -2177
rect 729 -2183 732 -2177
rect 736 -2183 739 -2177
rect 743 -2183 749 -2177
rect 750 -2183 753 -2177
rect 757 -2183 763 -2177
rect 764 -2183 767 -2177
rect 771 -2183 774 -2177
rect 778 -2183 781 -2177
rect 785 -2183 791 -2177
rect 792 -2183 795 -2177
rect 799 -2183 802 -2177
rect 806 -2183 809 -2177
rect 813 -2183 816 -2177
rect 820 -2183 823 -2177
rect 827 -2183 830 -2177
rect 834 -2183 837 -2177
rect 841 -2183 844 -2177
rect 848 -2183 851 -2177
rect 855 -2183 858 -2177
rect 862 -2183 865 -2177
rect 869 -2183 872 -2177
rect 876 -2183 879 -2177
rect 883 -2183 886 -2177
rect 890 -2183 893 -2177
rect 897 -2183 900 -2177
rect 904 -2183 907 -2177
rect 911 -2183 914 -2177
rect 918 -2183 921 -2177
rect 925 -2183 928 -2177
rect 932 -2183 935 -2177
rect 939 -2183 942 -2177
rect 946 -2183 949 -2177
rect 953 -2183 956 -2177
rect 960 -2183 963 -2177
rect 967 -2183 970 -2177
rect 974 -2183 980 -2177
rect 981 -2183 984 -2177
rect 988 -2183 991 -2177
rect 995 -2183 998 -2177
rect 1002 -2183 1005 -2177
rect 1009 -2183 1012 -2177
rect 1016 -2183 1019 -2177
rect 1023 -2183 1026 -2177
rect 1030 -2183 1033 -2177
rect 1037 -2183 1040 -2177
rect 1044 -2183 1047 -2177
rect 1051 -2183 1057 -2177
rect 1058 -2183 1061 -2177
rect 1065 -2183 1068 -2177
rect 1072 -2183 1075 -2177
rect 1079 -2183 1082 -2177
rect 1086 -2183 1089 -2177
rect 1093 -2183 1096 -2177
rect 1100 -2183 1103 -2177
rect 1107 -2183 1110 -2177
rect 1114 -2183 1117 -2177
rect 1121 -2183 1124 -2177
rect 1128 -2183 1131 -2177
rect 1135 -2183 1138 -2177
rect 1142 -2183 1145 -2177
rect 1149 -2183 1155 -2177
rect 1156 -2183 1159 -2177
rect 1163 -2183 1166 -2177
rect 1170 -2183 1173 -2177
rect 1177 -2183 1180 -2177
rect 1184 -2183 1190 -2177
rect 1191 -2183 1194 -2177
rect 1198 -2183 1204 -2177
rect 1205 -2183 1208 -2177
rect 1212 -2183 1215 -2177
rect 1219 -2183 1225 -2177
rect 1226 -2183 1232 -2177
rect 1233 -2183 1236 -2177
rect 1240 -2183 1243 -2177
rect 1247 -2183 1250 -2177
rect 1254 -2183 1260 -2177
rect 1261 -2183 1264 -2177
rect 1268 -2183 1271 -2177
rect 1275 -2183 1278 -2177
rect 1282 -2183 1285 -2177
rect 1289 -2183 1292 -2177
rect 1296 -2183 1299 -2177
rect 1303 -2183 1309 -2177
rect 1310 -2183 1313 -2177
rect 1317 -2183 1320 -2177
rect 1324 -2183 1327 -2177
rect 1331 -2183 1337 -2177
rect 1338 -2183 1344 -2177
rect 1345 -2183 1348 -2177
rect 1352 -2183 1355 -2177
rect 1359 -2183 1362 -2177
rect 1366 -2183 1372 -2177
rect 1373 -2183 1376 -2177
rect 1380 -2183 1386 -2177
rect 1387 -2183 1390 -2177
rect 1394 -2183 1397 -2177
rect 1401 -2183 1407 -2177
rect 1408 -2183 1411 -2177
rect 1415 -2183 1418 -2177
rect 1422 -2183 1425 -2177
rect 1429 -2183 1432 -2177
rect 1436 -2183 1439 -2177
rect 1443 -2183 1446 -2177
rect 1450 -2183 1453 -2177
rect 1457 -2183 1460 -2177
rect 1464 -2183 1467 -2177
rect 1471 -2183 1474 -2177
rect 1478 -2183 1481 -2177
rect 1485 -2183 1491 -2177
rect 1492 -2183 1495 -2177
rect 1499 -2183 1502 -2177
rect 1506 -2183 1509 -2177
rect 1513 -2183 1516 -2177
rect 1520 -2183 1523 -2177
rect 1527 -2183 1530 -2177
rect 1534 -2183 1537 -2177
rect 1541 -2183 1544 -2177
rect 1548 -2183 1551 -2177
rect 1555 -2183 1558 -2177
rect 1562 -2183 1565 -2177
rect 1569 -2183 1572 -2177
rect 1576 -2183 1582 -2177
rect 1583 -2183 1586 -2177
rect 1590 -2183 1593 -2177
rect 1597 -2183 1600 -2177
rect 1604 -2183 1607 -2177
rect 1611 -2183 1614 -2177
rect 1618 -2183 1621 -2177
rect 1625 -2183 1628 -2177
rect 1632 -2183 1635 -2177
rect 1639 -2183 1642 -2177
rect 1646 -2183 1652 -2177
rect 1653 -2183 1656 -2177
rect 1660 -2183 1663 -2177
rect 1667 -2183 1670 -2177
rect 1674 -2183 1677 -2177
rect 1681 -2183 1684 -2177
rect 1688 -2183 1691 -2177
rect 1695 -2183 1698 -2177
rect 1702 -2183 1705 -2177
rect 1709 -2183 1715 -2177
rect 1716 -2183 1719 -2177
rect 1723 -2183 1726 -2177
rect 1730 -2183 1733 -2177
rect 1737 -2183 1740 -2177
rect 1744 -2183 1747 -2177
rect 1751 -2183 1754 -2177
rect 1758 -2183 1761 -2177
rect 1765 -2183 1768 -2177
rect 1772 -2183 1775 -2177
rect 1779 -2183 1782 -2177
rect 1786 -2183 1789 -2177
rect 1793 -2183 1796 -2177
rect 1800 -2183 1803 -2177
rect 1807 -2183 1810 -2177
rect 1814 -2183 1817 -2177
rect 1821 -2183 1824 -2177
rect 1828 -2183 1831 -2177
rect 1835 -2183 1841 -2177
rect 1842 -2183 1845 -2177
rect 1849 -2183 1852 -2177
rect 1856 -2183 1862 -2177
rect 1863 -2183 1866 -2177
rect 1870 -2183 1873 -2177
rect 1877 -2183 1880 -2177
rect 1884 -2183 1887 -2177
rect 1891 -2183 1894 -2177
rect 1898 -2183 1901 -2177
rect 1905 -2183 1908 -2177
rect 1912 -2183 1915 -2177
rect 1919 -2183 1922 -2177
rect 1926 -2183 1929 -2177
rect 1933 -2183 1936 -2177
rect 1940 -2183 1943 -2177
rect 1947 -2183 1950 -2177
rect 1954 -2183 1960 -2177
rect 1961 -2183 1964 -2177
rect 1968 -2183 1971 -2177
rect 1975 -2183 1978 -2177
rect 1982 -2183 1985 -2177
rect 1989 -2183 1992 -2177
rect 1996 -2183 1999 -2177
rect 2003 -2183 2006 -2177
rect 2010 -2183 2013 -2177
rect 2017 -2183 2020 -2177
rect 2024 -2183 2027 -2177
rect 2031 -2183 2034 -2177
rect 2038 -2183 2041 -2177
rect 2045 -2183 2048 -2177
rect 2052 -2183 2055 -2177
rect 2059 -2183 2062 -2177
rect 2066 -2183 2069 -2177
rect 2073 -2183 2076 -2177
rect 2080 -2183 2083 -2177
rect 2087 -2183 2090 -2177
rect 2094 -2183 2097 -2177
rect 2101 -2183 2104 -2177
rect 2108 -2183 2111 -2177
rect 2115 -2183 2118 -2177
rect 2122 -2183 2125 -2177
rect 2129 -2183 2132 -2177
rect 2136 -2183 2139 -2177
rect 2143 -2183 2146 -2177
rect 2150 -2183 2153 -2177
rect 2157 -2183 2160 -2177
rect 2164 -2183 2167 -2177
rect 2171 -2183 2174 -2177
rect 2178 -2183 2181 -2177
rect 2185 -2183 2188 -2177
rect 2192 -2183 2195 -2177
rect 2199 -2183 2202 -2177
rect 2206 -2183 2209 -2177
rect 2213 -2183 2216 -2177
rect 2220 -2183 2223 -2177
rect 2227 -2183 2230 -2177
rect 2234 -2183 2237 -2177
rect 2241 -2183 2244 -2177
rect 2248 -2183 2251 -2177
rect 2255 -2183 2258 -2177
rect 2262 -2183 2265 -2177
rect 2269 -2183 2272 -2177
rect 2276 -2183 2279 -2177
rect 2283 -2183 2286 -2177
rect 2290 -2183 2293 -2177
rect 2297 -2183 2300 -2177
rect 2304 -2183 2307 -2177
rect 2311 -2183 2314 -2177
rect 2318 -2183 2321 -2177
rect 2325 -2183 2328 -2177
rect 2332 -2183 2335 -2177
rect 2339 -2183 2342 -2177
rect 2346 -2183 2349 -2177
rect 2353 -2183 2356 -2177
rect 2360 -2183 2363 -2177
rect 2367 -2183 2370 -2177
rect 2374 -2183 2377 -2177
rect 2381 -2183 2384 -2177
rect 2388 -2183 2391 -2177
rect 2395 -2183 2398 -2177
rect 2402 -2183 2405 -2177
rect 2409 -2183 2412 -2177
rect 2416 -2183 2419 -2177
rect 2423 -2183 2426 -2177
rect 1 -2332 4 -2326
rect 8 -2332 14 -2326
rect 15 -2332 18 -2326
rect 22 -2332 25 -2326
rect 29 -2332 35 -2326
rect 36 -2332 39 -2326
rect 43 -2332 46 -2326
rect 50 -2332 53 -2326
rect 57 -2332 60 -2326
rect 64 -2332 67 -2326
rect 71 -2332 74 -2326
rect 78 -2332 81 -2326
rect 85 -2332 88 -2326
rect 92 -2332 98 -2326
rect 99 -2332 102 -2326
rect 106 -2332 109 -2326
rect 113 -2332 116 -2326
rect 120 -2332 123 -2326
rect 127 -2332 130 -2326
rect 134 -2332 137 -2326
rect 141 -2332 147 -2326
rect 148 -2332 151 -2326
rect 155 -2332 158 -2326
rect 162 -2332 168 -2326
rect 169 -2332 172 -2326
rect 176 -2332 179 -2326
rect 183 -2332 186 -2326
rect 190 -2332 193 -2326
rect 197 -2332 200 -2326
rect 204 -2332 207 -2326
rect 211 -2332 214 -2326
rect 218 -2332 221 -2326
rect 225 -2332 228 -2326
rect 232 -2332 235 -2326
rect 239 -2332 245 -2326
rect 246 -2332 252 -2326
rect 253 -2332 256 -2326
rect 260 -2332 263 -2326
rect 267 -2332 270 -2326
rect 274 -2332 277 -2326
rect 281 -2332 284 -2326
rect 288 -2332 291 -2326
rect 295 -2332 298 -2326
rect 302 -2332 305 -2326
rect 309 -2332 312 -2326
rect 316 -2332 319 -2326
rect 323 -2332 326 -2326
rect 330 -2332 333 -2326
rect 337 -2332 340 -2326
rect 344 -2332 347 -2326
rect 351 -2332 354 -2326
rect 358 -2332 361 -2326
rect 365 -2332 368 -2326
rect 372 -2332 375 -2326
rect 379 -2332 382 -2326
rect 386 -2332 389 -2326
rect 393 -2332 396 -2326
rect 400 -2332 403 -2326
rect 407 -2332 410 -2326
rect 414 -2332 417 -2326
rect 421 -2332 424 -2326
rect 428 -2332 434 -2326
rect 435 -2332 438 -2326
rect 442 -2332 445 -2326
rect 449 -2332 452 -2326
rect 456 -2332 459 -2326
rect 463 -2332 466 -2326
rect 470 -2332 473 -2326
rect 477 -2332 480 -2326
rect 484 -2332 487 -2326
rect 491 -2332 494 -2326
rect 498 -2332 501 -2326
rect 505 -2332 508 -2326
rect 512 -2332 515 -2326
rect 519 -2332 522 -2326
rect 526 -2332 529 -2326
rect 533 -2332 536 -2326
rect 540 -2332 543 -2326
rect 547 -2332 550 -2326
rect 554 -2332 557 -2326
rect 561 -2332 564 -2326
rect 568 -2332 571 -2326
rect 575 -2332 578 -2326
rect 582 -2332 585 -2326
rect 589 -2332 595 -2326
rect 596 -2332 599 -2326
rect 603 -2332 606 -2326
rect 610 -2332 613 -2326
rect 617 -2332 623 -2326
rect 624 -2332 630 -2326
rect 631 -2332 634 -2326
rect 638 -2332 641 -2326
rect 645 -2332 648 -2326
rect 652 -2332 655 -2326
rect 659 -2332 665 -2326
rect 666 -2332 672 -2326
rect 673 -2332 676 -2326
rect 680 -2332 683 -2326
rect 687 -2332 690 -2326
rect 694 -2332 697 -2326
rect 701 -2332 707 -2326
rect 708 -2332 711 -2326
rect 715 -2332 718 -2326
rect 722 -2332 728 -2326
rect 729 -2332 732 -2326
rect 736 -2332 739 -2326
rect 743 -2332 746 -2326
rect 750 -2332 753 -2326
rect 757 -2332 760 -2326
rect 764 -2332 770 -2326
rect 771 -2332 774 -2326
rect 778 -2332 784 -2326
rect 785 -2332 788 -2326
rect 792 -2332 795 -2326
rect 799 -2332 802 -2326
rect 806 -2332 809 -2326
rect 813 -2332 816 -2326
rect 820 -2332 823 -2326
rect 827 -2332 830 -2326
rect 834 -2332 837 -2326
rect 841 -2332 844 -2326
rect 848 -2332 851 -2326
rect 855 -2332 861 -2326
rect 862 -2332 865 -2326
rect 869 -2332 872 -2326
rect 876 -2332 879 -2326
rect 883 -2332 886 -2326
rect 890 -2332 893 -2326
rect 897 -2332 900 -2326
rect 904 -2332 907 -2326
rect 911 -2332 914 -2326
rect 918 -2332 924 -2326
rect 925 -2332 928 -2326
rect 932 -2332 938 -2326
rect 939 -2332 942 -2326
rect 946 -2332 949 -2326
rect 953 -2332 956 -2326
rect 960 -2332 963 -2326
rect 967 -2332 970 -2326
rect 974 -2332 980 -2326
rect 981 -2332 984 -2326
rect 988 -2332 994 -2326
rect 995 -2332 998 -2326
rect 1002 -2332 1005 -2326
rect 1009 -2332 1012 -2326
rect 1016 -2332 1019 -2326
rect 1023 -2332 1026 -2326
rect 1030 -2332 1033 -2326
rect 1037 -2332 1043 -2326
rect 1044 -2332 1047 -2326
rect 1051 -2332 1054 -2326
rect 1058 -2332 1061 -2326
rect 1065 -2332 1068 -2326
rect 1072 -2332 1075 -2326
rect 1079 -2332 1082 -2326
rect 1086 -2332 1089 -2326
rect 1093 -2332 1096 -2326
rect 1100 -2332 1103 -2326
rect 1107 -2332 1110 -2326
rect 1114 -2332 1117 -2326
rect 1121 -2332 1124 -2326
rect 1128 -2332 1131 -2326
rect 1135 -2332 1141 -2326
rect 1142 -2332 1145 -2326
rect 1149 -2332 1152 -2326
rect 1156 -2332 1159 -2326
rect 1163 -2332 1166 -2326
rect 1170 -2332 1173 -2326
rect 1177 -2332 1180 -2326
rect 1184 -2332 1187 -2326
rect 1191 -2332 1194 -2326
rect 1198 -2332 1201 -2326
rect 1205 -2332 1208 -2326
rect 1212 -2332 1215 -2326
rect 1219 -2332 1222 -2326
rect 1226 -2332 1229 -2326
rect 1233 -2332 1236 -2326
rect 1240 -2332 1243 -2326
rect 1247 -2332 1253 -2326
rect 1254 -2332 1257 -2326
rect 1261 -2332 1264 -2326
rect 1268 -2332 1271 -2326
rect 1275 -2332 1278 -2326
rect 1282 -2332 1285 -2326
rect 1289 -2332 1295 -2326
rect 1296 -2332 1299 -2326
rect 1303 -2332 1306 -2326
rect 1310 -2332 1313 -2326
rect 1317 -2332 1323 -2326
rect 1324 -2332 1327 -2326
rect 1331 -2332 1334 -2326
rect 1338 -2332 1341 -2326
rect 1345 -2332 1348 -2326
rect 1352 -2332 1355 -2326
rect 1359 -2332 1362 -2326
rect 1366 -2332 1369 -2326
rect 1373 -2332 1376 -2326
rect 1380 -2332 1383 -2326
rect 1387 -2332 1390 -2326
rect 1394 -2332 1400 -2326
rect 1401 -2332 1404 -2326
rect 1408 -2332 1411 -2326
rect 1415 -2332 1418 -2326
rect 1422 -2332 1425 -2326
rect 1429 -2332 1432 -2326
rect 1436 -2332 1439 -2326
rect 1443 -2332 1446 -2326
rect 1450 -2332 1453 -2326
rect 1457 -2332 1460 -2326
rect 1464 -2332 1467 -2326
rect 1471 -2332 1474 -2326
rect 1478 -2332 1481 -2326
rect 1485 -2332 1488 -2326
rect 1492 -2332 1498 -2326
rect 1499 -2332 1505 -2326
rect 1506 -2332 1509 -2326
rect 1513 -2332 1519 -2326
rect 1520 -2332 1523 -2326
rect 1527 -2332 1530 -2326
rect 1534 -2332 1537 -2326
rect 1541 -2332 1547 -2326
rect 1548 -2332 1551 -2326
rect 1555 -2332 1558 -2326
rect 1562 -2332 1565 -2326
rect 1569 -2332 1572 -2326
rect 1576 -2332 1579 -2326
rect 1583 -2332 1586 -2326
rect 1590 -2332 1593 -2326
rect 1597 -2332 1600 -2326
rect 1604 -2332 1607 -2326
rect 1611 -2332 1614 -2326
rect 1618 -2332 1621 -2326
rect 1625 -2332 1631 -2326
rect 1632 -2332 1635 -2326
rect 1639 -2332 1642 -2326
rect 1646 -2332 1649 -2326
rect 1653 -2332 1656 -2326
rect 1660 -2332 1663 -2326
rect 1667 -2332 1670 -2326
rect 1674 -2332 1677 -2326
rect 1681 -2332 1687 -2326
rect 1688 -2332 1691 -2326
rect 1695 -2332 1698 -2326
rect 1702 -2332 1705 -2326
rect 1709 -2332 1712 -2326
rect 1716 -2332 1719 -2326
rect 1723 -2332 1726 -2326
rect 1730 -2332 1733 -2326
rect 1737 -2332 1740 -2326
rect 1744 -2332 1747 -2326
rect 1751 -2332 1754 -2326
rect 1758 -2332 1761 -2326
rect 1765 -2332 1768 -2326
rect 1772 -2332 1775 -2326
rect 1779 -2332 1782 -2326
rect 1786 -2332 1789 -2326
rect 1793 -2332 1796 -2326
rect 1800 -2332 1803 -2326
rect 1807 -2332 1810 -2326
rect 1814 -2332 1817 -2326
rect 1821 -2332 1824 -2326
rect 1828 -2332 1831 -2326
rect 1835 -2332 1838 -2326
rect 1842 -2332 1845 -2326
rect 1849 -2332 1852 -2326
rect 1856 -2332 1859 -2326
rect 1863 -2332 1866 -2326
rect 1870 -2332 1873 -2326
rect 1877 -2332 1880 -2326
rect 1884 -2332 1887 -2326
rect 1891 -2332 1897 -2326
rect 1898 -2332 1901 -2326
rect 1905 -2332 1908 -2326
rect 1912 -2332 1915 -2326
rect 1919 -2332 1922 -2326
rect 1926 -2332 1929 -2326
rect 1933 -2332 1939 -2326
rect 1940 -2332 1943 -2326
rect 1947 -2332 1950 -2326
rect 1954 -2332 1957 -2326
rect 1961 -2332 1964 -2326
rect 1968 -2332 1971 -2326
rect 1975 -2332 1981 -2326
rect 1982 -2332 1985 -2326
rect 1989 -2332 1992 -2326
rect 1996 -2332 1999 -2326
rect 2003 -2332 2006 -2326
rect 2010 -2332 2013 -2326
rect 2017 -2332 2020 -2326
rect 2024 -2332 2027 -2326
rect 2031 -2332 2034 -2326
rect 2038 -2332 2041 -2326
rect 2045 -2332 2048 -2326
rect 2052 -2332 2055 -2326
rect 2059 -2332 2062 -2326
rect 2066 -2332 2069 -2326
rect 2073 -2332 2076 -2326
rect 2080 -2332 2083 -2326
rect 2087 -2332 2090 -2326
rect 2094 -2332 2097 -2326
rect 2101 -2332 2104 -2326
rect 2108 -2332 2111 -2326
rect 2115 -2332 2118 -2326
rect 2122 -2332 2125 -2326
rect 2129 -2332 2132 -2326
rect 2136 -2332 2139 -2326
rect 2143 -2332 2146 -2326
rect 2150 -2332 2153 -2326
rect 2157 -2332 2160 -2326
rect 2164 -2332 2167 -2326
rect 2171 -2332 2174 -2326
rect 2178 -2332 2181 -2326
rect 2185 -2332 2188 -2326
rect 2192 -2332 2195 -2326
rect 2199 -2332 2202 -2326
rect 2206 -2332 2209 -2326
rect 2213 -2332 2216 -2326
rect 2220 -2332 2223 -2326
rect 2227 -2332 2230 -2326
rect 2234 -2332 2237 -2326
rect 2241 -2332 2244 -2326
rect 2248 -2332 2251 -2326
rect 2255 -2332 2258 -2326
rect 2262 -2332 2265 -2326
rect 2269 -2332 2272 -2326
rect 2276 -2332 2279 -2326
rect 2283 -2332 2286 -2326
rect 2290 -2332 2293 -2326
rect 2297 -2332 2300 -2326
rect 2304 -2332 2307 -2326
rect 2311 -2332 2314 -2326
rect 2318 -2332 2321 -2326
rect 2325 -2332 2328 -2326
rect 2332 -2332 2338 -2326
rect 2339 -2332 2345 -2326
rect 2346 -2332 2349 -2326
rect 1 -2505 7 -2499
rect 8 -2505 14 -2499
rect 15 -2505 21 -2499
rect 22 -2505 25 -2499
rect 29 -2505 35 -2499
rect 36 -2505 42 -2499
rect 43 -2505 46 -2499
rect 50 -2505 53 -2499
rect 57 -2505 63 -2499
rect 64 -2505 67 -2499
rect 71 -2505 74 -2499
rect 78 -2505 81 -2499
rect 85 -2505 88 -2499
rect 92 -2505 98 -2499
rect 99 -2505 102 -2499
rect 106 -2505 112 -2499
rect 113 -2505 116 -2499
rect 120 -2505 123 -2499
rect 127 -2505 130 -2499
rect 134 -2505 137 -2499
rect 141 -2505 144 -2499
rect 148 -2505 151 -2499
rect 155 -2505 158 -2499
rect 162 -2505 168 -2499
rect 169 -2505 172 -2499
rect 176 -2505 179 -2499
rect 183 -2505 186 -2499
rect 190 -2505 193 -2499
rect 197 -2505 200 -2499
rect 204 -2505 207 -2499
rect 211 -2505 214 -2499
rect 218 -2505 221 -2499
rect 225 -2505 228 -2499
rect 232 -2505 235 -2499
rect 239 -2505 242 -2499
rect 246 -2505 249 -2499
rect 253 -2505 256 -2499
rect 260 -2505 263 -2499
rect 267 -2505 270 -2499
rect 274 -2505 277 -2499
rect 281 -2505 284 -2499
rect 288 -2505 291 -2499
rect 295 -2505 298 -2499
rect 302 -2505 305 -2499
rect 309 -2505 312 -2499
rect 316 -2505 319 -2499
rect 323 -2505 326 -2499
rect 330 -2505 333 -2499
rect 337 -2505 340 -2499
rect 344 -2505 347 -2499
rect 351 -2505 354 -2499
rect 358 -2505 361 -2499
rect 365 -2505 368 -2499
rect 372 -2505 375 -2499
rect 379 -2505 382 -2499
rect 386 -2505 389 -2499
rect 393 -2505 396 -2499
rect 400 -2505 403 -2499
rect 407 -2505 410 -2499
rect 414 -2505 417 -2499
rect 421 -2505 424 -2499
rect 428 -2505 431 -2499
rect 435 -2505 438 -2499
rect 442 -2505 445 -2499
rect 449 -2505 452 -2499
rect 456 -2505 459 -2499
rect 463 -2505 466 -2499
rect 470 -2505 473 -2499
rect 477 -2505 483 -2499
rect 484 -2505 487 -2499
rect 491 -2505 494 -2499
rect 498 -2505 501 -2499
rect 505 -2505 508 -2499
rect 512 -2505 515 -2499
rect 519 -2505 522 -2499
rect 526 -2505 529 -2499
rect 533 -2505 536 -2499
rect 540 -2505 543 -2499
rect 547 -2505 550 -2499
rect 554 -2505 557 -2499
rect 561 -2505 564 -2499
rect 568 -2505 571 -2499
rect 575 -2505 578 -2499
rect 582 -2505 585 -2499
rect 589 -2505 592 -2499
rect 596 -2505 599 -2499
rect 603 -2505 609 -2499
rect 610 -2505 613 -2499
rect 617 -2505 620 -2499
rect 624 -2505 627 -2499
rect 631 -2505 634 -2499
rect 638 -2505 641 -2499
rect 645 -2505 648 -2499
rect 652 -2505 655 -2499
rect 659 -2505 662 -2499
rect 666 -2505 672 -2499
rect 673 -2505 676 -2499
rect 680 -2505 683 -2499
rect 687 -2505 690 -2499
rect 694 -2505 697 -2499
rect 701 -2505 704 -2499
rect 708 -2505 711 -2499
rect 715 -2505 718 -2499
rect 722 -2505 725 -2499
rect 729 -2505 732 -2499
rect 736 -2505 742 -2499
rect 743 -2505 746 -2499
rect 750 -2505 753 -2499
rect 757 -2505 760 -2499
rect 764 -2505 767 -2499
rect 771 -2505 777 -2499
rect 778 -2505 781 -2499
rect 785 -2505 788 -2499
rect 792 -2505 798 -2499
rect 799 -2505 802 -2499
rect 806 -2505 809 -2499
rect 813 -2505 816 -2499
rect 820 -2505 823 -2499
rect 827 -2505 830 -2499
rect 834 -2505 837 -2499
rect 841 -2505 844 -2499
rect 848 -2505 851 -2499
rect 855 -2505 861 -2499
rect 862 -2505 865 -2499
rect 869 -2505 875 -2499
rect 876 -2505 879 -2499
rect 883 -2505 886 -2499
rect 890 -2505 893 -2499
rect 897 -2505 900 -2499
rect 904 -2505 907 -2499
rect 911 -2505 914 -2499
rect 918 -2505 924 -2499
rect 925 -2505 928 -2499
rect 932 -2505 935 -2499
rect 939 -2505 942 -2499
rect 946 -2505 949 -2499
rect 953 -2505 959 -2499
rect 960 -2505 963 -2499
rect 967 -2505 970 -2499
rect 974 -2505 980 -2499
rect 981 -2505 984 -2499
rect 988 -2505 994 -2499
rect 995 -2505 998 -2499
rect 1002 -2505 1005 -2499
rect 1009 -2505 1015 -2499
rect 1016 -2505 1022 -2499
rect 1023 -2505 1026 -2499
rect 1030 -2505 1033 -2499
rect 1037 -2505 1040 -2499
rect 1044 -2505 1047 -2499
rect 1051 -2505 1057 -2499
rect 1058 -2505 1061 -2499
rect 1065 -2505 1068 -2499
rect 1072 -2505 1078 -2499
rect 1079 -2505 1085 -2499
rect 1086 -2505 1089 -2499
rect 1093 -2505 1096 -2499
rect 1100 -2505 1103 -2499
rect 1107 -2505 1110 -2499
rect 1114 -2505 1117 -2499
rect 1121 -2505 1124 -2499
rect 1128 -2505 1131 -2499
rect 1135 -2505 1138 -2499
rect 1142 -2505 1145 -2499
rect 1149 -2505 1152 -2499
rect 1156 -2505 1159 -2499
rect 1163 -2505 1166 -2499
rect 1170 -2505 1176 -2499
rect 1177 -2505 1180 -2499
rect 1184 -2505 1187 -2499
rect 1191 -2505 1194 -2499
rect 1198 -2505 1201 -2499
rect 1205 -2505 1208 -2499
rect 1212 -2505 1218 -2499
rect 1219 -2505 1222 -2499
rect 1226 -2505 1229 -2499
rect 1233 -2505 1236 -2499
rect 1240 -2505 1243 -2499
rect 1247 -2505 1250 -2499
rect 1254 -2505 1257 -2499
rect 1261 -2505 1264 -2499
rect 1268 -2505 1274 -2499
rect 1275 -2505 1278 -2499
rect 1282 -2505 1285 -2499
rect 1289 -2505 1295 -2499
rect 1296 -2505 1299 -2499
rect 1303 -2505 1306 -2499
rect 1310 -2505 1313 -2499
rect 1317 -2505 1320 -2499
rect 1324 -2505 1327 -2499
rect 1331 -2505 1337 -2499
rect 1338 -2505 1341 -2499
rect 1345 -2505 1348 -2499
rect 1352 -2505 1358 -2499
rect 1359 -2505 1365 -2499
rect 1366 -2505 1369 -2499
rect 1373 -2505 1379 -2499
rect 1380 -2505 1383 -2499
rect 1387 -2505 1390 -2499
rect 1394 -2505 1397 -2499
rect 1401 -2505 1404 -2499
rect 1408 -2505 1411 -2499
rect 1415 -2505 1418 -2499
rect 1422 -2505 1425 -2499
rect 1429 -2505 1432 -2499
rect 1436 -2505 1439 -2499
rect 1443 -2505 1446 -2499
rect 1450 -2505 1453 -2499
rect 1457 -2505 1460 -2499
rect 1464 -2505 1467 -2499
rect 1471 -2505 1474 -2499
rect 1478 -2505 1481 -2499
rect 1485 -2505 1488 -2499
rect 1492 -2505 1495 -2499
rect 1499 -2505 1502 -2499
rect 1506 -2505 1509 -2499
rect 1513 -2505 1516 -2499
rect 1520 -2505 1523 -2499
rect 1527 -2505 1530 -2499
rect 1534 -2505 1537 -2499
rect 1541 -2505 1544 -2499
rect 1548 -2505 1551 -2499
rect 1555 -2505 1558 -2499
rect 1562 -2505 1565 -2499
rect 1569 -2505 1572 -2499
rect 1576 -2505 1582 -2499
rect 1583 -2505 1586 -2499
rect 1590 -2505 1593 -2499
rect 1597 -2505 1603 -2499
rect 1604 -2505 1607 -2499
rect 1611 -2505 1614 -2499
rect 1618 -2505 1621 -2499
rect 1625 -2505 1628 -2499
rect 1632 -2505 1635 -2499
rect 1639 -2505 1642 -2499
rect 1646 -2505 1649 -2499
rect 1653 -2505 1656 -2499
rect 1660 -2505 1663 -2499
rect 1667 -2505 1670 -2499
rect 1674 -2505 1680 -2499
rect 1681 -2505 1684 -2499
rect 1688 -2505 1691 -2499
rect 1695 -2505 1698 -2499
rect 1702 -2505 1705 -2499
rect 1709 -2505 1712 -2499
rect 1716 -2505 1719 -2499
rect 1723 -2505 1726 -2499
rect 1730 -2505 1733 -2499
rect 1737 -2505 1740 -2499
rect 1744 -2505 1747 -2499
rect 1751 -2505 1754 -2499
rect 1758 -2505 1761 -2499
rect 1765 -2505 1768 -2499
rect 1772 -2505 1775 -2499
rect 1779 -2505 1782 -2499
rect 1786 -2505 1789 -2499
rect 1793 -2505 1796 -2499
rect 1800 -2505 1806 -2499
rect 1807 -2505 1810 -2499
rect 1814 -2505 1817 -2499
rect 1821 -2505 1824 -2499
rect 1828 -2505 1831 -2499
rect 1835 -2505 1838 -2499
rect 1842 -2505 1845 -2499
rect 1849 -2505 1852 -2499
rect 1856 -2505 1859 -2499
rect 1863 -2505 1866 -2499
rect 1870 -2505 1873 -2499
rect 1877 -2505 1880 -2499
rect 1884 -2505 1887 -2499
rect 1891 -2505 1894 -2499
rect 1898 -2505 1901 -2499
rect 1905 -2505 1908 -2499
rect 1912 -2505 1915 -2499
rect 1919 -2505 1922 -2499
rect 1926 -2505 1929 -2499
rect 1933 -2505 1936 -2499
rect 1940 -2505 1943 -2499
rect 1947 -2505 1950 -2499
rect 1954 -2505 1957 -2499
rect 1961 -2505 1964 -2499
rect 1968 -2505 1971 -2499
rect 1975 -2505 1978 -2499
rect 1982 -2505 1985 -2499
rect 1989 -2505 1992 -2499
rect 1996 -2505 1999 -2499
rect 2003 -2505 2006 -2499
rect 2010 -2505 2013 -2499
rect 2017 -2505 2020 -2499
rect 2024 -2505 2027 -2499
rect 2031 -2505 2034 -2499
rect 2038 -2505 2041 -2499
rect 2045 -2505 2048 -2499
rect 2052 -2505 2055 -2499
rect 2059 -2505 2062 -2499
rect 2066 -2505 2069 -2499
rect 2073 -2505 2076 -2499
rect 2080 -2505 2083 -2499
rect 2087 -2505 2090 -2499
rect 2094 -2505 2097 -2499
rect 2101 -2505 2104 -2499
rect 2108 -2505 2111 -2499
rect 2115 -2505 2118 -2499
rect 2122 -2505 2125 -2499
rect 2129 -2505 2132 -2499
rect 2136 -2505 2139 -2499
rect 2143 -2505 2146 -2499
rect 2150 -2505 2153 -2499
rect 2157 -2505 2160 -2499
rect 2164 -2505 2167 -2499
rect 2171 -2505 2174 -2499
rect 2178 -2505 2181 -2499
rect 2185 -2505 2188 -2499
rect 2192 -2505 2195 -2499
rect 2199 -2505 2202 -2499
rect 2206 -2505 2209 -2499
rect 2213 -2505 2216 -2499
rect 2220 -2505 2223 -2499
rect 2227 -2505 2230 -2499
rect 2234 -2505 2237 -2499
rect 2241 -2505 2244 -2499
rect 2248 -2505 2251 -2499
rect 2255 -2505 2258 -2499
rect 2262 -2505 2265 -2499
rect 2269 -2505 2272 -2499
rect 2276 -2505 2282 -2499
rect 2283 -2505 2286 -2499
rect 2290 -2505 2293 -2499
rect 2297 -2505 2300 -2499
rect 2304 -2505 2307 -2499
rect 2311 -2505 2314 -2499
rect 1 -2678 7 -2672
rect 8 -2678 11 -2672
rect 15 -2678 18 -2672
rect 22 -2678 28 -2672
rect 29 -2678 32 -2672
rect 36 -2678 39 -2672
rect 43 -2678 46 -2672
rect 50 -2678 56 -2672
rect 57 -2678 60 -2672
rect 64 -2678 70 -2672
rect 71 -2678 77 -2672
rect 78 -2678 81 -2672
rect 85 -2678 88 -2672
rect 92 -2678 95 -2672
rect 99 -2678 105 -2672
rect 106 -2678 109 -2672
rect 113 -2678 116 -2672
rect 120 -2678 123 -2672
rect 127 -2678 133 -2672
rect 134 -2678 137 -2672
rect 141 -2678 144 -2672
rect 148 -2678 151 -2672
rect 155 -2678 158 -2672
rect 162 -2678 165 -2672
rect 169 -2678 172 -2672
rect 176 -2678 179 -2672
rect 183 -2678 186 -2672
rect 190 -2678 193 -2672
rect 197 -2678 203 -2672
rect 204 -2678 207 -2672
rect 211 -2678 214 -2672
rect 218 -2678 221 -2672
rect 225 -2678 228 -2672
rect 232 -2678 235 -2672
rect 239 -2678 245 -2672
rect 246 -2678 249 -2672
rect 253 -2678 256 -2672
rect 260 -2678 263 -2672
rect 267 -2678 270 -2672
rect 274 -2678 277 -2672
rect 281 -2678 284 -2672
rect 288 -2678 291 -2672
rect 295 -2678 298 -2672
rect 302 -2678 305 -2672
rect 309 -2678 312 -2672
rect 316 -2678 319 -2672
rect 323 -2678 326 -2672
rect 330 -2678 333 -2672
rect 337 -2678 340 -2672
rect 344 -2678 347 -2672
rect 351 -2678 354 -2672
rect 358 -2678 361 -2672
rect 365 -2678 368 -2672
rect 372 -2678 375 -2672
rect 379 -2678 382 -2672
rect 386 -2678 389 -2672
rect 393 -2678 396 -2672
rect 400 -2678 403 -2672
rect 407 -2678 413 -2672
rect 414 -2678 417 -2672
rect 421 -2678 424 -2672
rect 428 -2678 431 -2672
rect 435 -2678 438 -2672
rect 442 -2678 445 -2672
rect 449 -2678 452 -2672
rect 456 -2678 459 -2672
rect 463 -2678 466 -2672
rect 470 -2678 473 -2672
rect 477 -2678 480 -2672
rect 484 -2678 487 -2672
rect 491 -2678 494 -2672
rect 498 -2678 501 -2672
rect 505 -2678 508 -2672
rect 512 -2678 515 -2672
rect 519 -2678 522 -2672
rect 526 -2678 529 -2672
rect 533 -2678 536 -2672
rect 540 -2678 543 -2672
rect 547 -2678 550 -2672
rect 554 -2678 560 -2672
rect 561 -2678 564 -2672
rect 568 -2678 571 -2672
rect 575 -2678 578 -2672
rect 582 -2678 585 -2672
rect 589 -2678 592 -2672
rect 596 -2678 599 -2672
rect 603 -2678 606 -2672
rect 610 -2678 613 -2672
rect 617 -2678 620 -2672
rect 624 -2678 627 -2672
rect 631 -2678 634 -2672
rect 638 -2678 641 -2672
rect 645 -2678 648 -2672
rect 652 -2678 655 -2672
rect 659 -2678 662 -2672
rect 666 -2678 669 -2672
rect 673 -2678 676 -2672
rect 680 -2678 683 -2672
rect 687 -2678 690 -2672
rect 694 -2678 697 -2672
rect 701 -2678 704 -2672
rect 708 -2678 711 -2672
rect 715 -2678 718 -2672
rect 722 -2678 728 -2672
rect 729 -2678 732 -2672
rect 736 -2678 739 -2672
rect 743 -2678 746 -2672
rect 750 -2678 753 -2672
rect 757 -2678 760 -2672
rect 764 -2678 767 -2672
rect 771 -2678 774 -2672
rect 778 -2678 781 -2672
rect 785 -2678 791 -2672
rect 792 -2678 795 -2672
rect 799 -2678 802 -2672
rect 806 -2678 812 -2672
rect 813 -2678 819 -2672
rect 820 -2678 826 -2672
rect 827 -2678 830 -2672
rect 834 -2678 837 -2672
rect 841 -2678 844 -2672
rect 848 -2678 851 -2672
rect 855 -2678 858 -2672
rect 862 -2678 865 -2672
rect 869 -2678 872 -2672
rect 876 -2678 879 -2672
rect 883 -2678 886 -2672
rect 890 -2678 896 -2672
rect 897 -2678 900 -2672
rect 904 -2678 907 -2672
rect 911 -2678 914 -2672
rect 918 -2678 924 -2672
rect 925 -2678 928 -2672
rect 932 -2678 935 -2672
rect 939 -2678 942 -2672
rect 946 -2678 952 -2672
rect 953 -2678 959 -2672
rect 960 -2678 963 -2672
rect 967 -2678 970 -2672
rect 974 -2678 977 -2672
rect 981 -2678 984 -2672
rect 988 -2678 991 -2672
rect 995 -2678 998 -2672
rect 1002 -2678 1008 -2672
rect 1009 -2678 1015 -2672
rect 1016 -2678 1019 -2672
rect 1023 -2678 1026 -2672
rect 1030 -2678 1033 -2672
rect 1037 -2678 1043 -2672
rect 1044 -2678 1047 -2672
rect 1051 -2678 1054 -2672
rect 1058 -2678 1061 -2672
rect 1065 -2678 1068 -2672
rect 1072 -2678 1075 -2672
rect 1079 -2678 1082 -2672
rect 1086 -2678 1089 -2672
rect 1093 -2678 1096 -2672
rect 1100 -2678 1103 -2672
rect 1107 -2678 1110 -2672
rect 1114 -2678 1117 -2672
rect 1121 -2678 1127 -2672
rect 1128 -2678 1131 -2672
rect 1135 -2678 1141 -2672
rect 1142 -2678 1145 -2672
rect 1149 -2678 1152 -2672
rect 1156 -2678 1159 -2672
rect 1163 -2678 1166 -2672
rect 1170 -2678 1173 -2672
rect 1177 -2678 1180 -2672
rect 1184 -2678 1190 -2672
rect 1191 -2678 1197 -2672
rect 1198 -2678 1201 -2672
rect 1205 -2678 1208 -2672
rect 1212 -2678 1215 -2672
rect 1219 -2678 1222 -2672
rect 1226 -2678 1229 -2672
rect 1233 -2678 1239 -2672
rect 1240 -2678 1246 -2672
rect 1247 -2678 1250 -2672
rect 1254 -2678 1257 -2672
rect 1261 -2678 1264 -2672
rect 1268 -2678 1271 -2672
rect 1275 -2678 1278 -2672
rect 1282 -2678 1285 -2672
rect 1289 -2678 1292 -2672
rect 1296 -2678 1299 -2672
rect 1303 -2678 1306 -2672
rect 1310 -2678 1316 -2672
rect 1317 -2678 1320 -2672
rect 1324 -2678 1330 -2672
rect 1331 -2678 1334 -2672
rect 1338 -2678 1341 -2672
rect 1345 -2678 1348 -2672
rect 1352 -2678 1355 -2672
rect 1359 -2678 1362 -2672
rect 1366 -2678 1369 -2672
rect 1373 -2678 1376 -2672
rect 1380 -2678 1383 -2672
rect 1387 -2678 1390 -2672
rect 1394 -2678 1400 -2672
rect 1401 -2678 1404 -2672
rect 1408 -2678 1414 -2672
rect 1415 -2678 1418 -2672
rect 1422 -2678 1425 -2672
rect 1429 -2678 1435 -2672
rect 1436 -2678 1442 -2672
rect 1443 -2678 1449 -2672
rect 1450 -2678 1453 -2672
rect 1457 -2678 1460 -2672
rect 1464 -2678 1467 -2672
rect 1471 -2678 1474 -2672
rect 1478 -2678 1481 -2672
rect 1485 -2678 1488 -2672
rect 1492 -2678 1495 -2672
rect 1499 -2678 1502 -2672
rect 1506 -2678 1512 -2672
rect 1513 -2678 1516 -2672
rect 1520 -2678 1523 -2672
rect 1527 -2678 1530 -2672
rect 1534 -2678 1537 -2672
rect 1541 -2678 1544 -2672
rect 1548 -2678 1551 -2672
rect 1555 -2678 1558 -2672
rect 1562 -2678 1565 -2672
rect 1569 -2678 1572 -2672
rect 1576 -2678 1582 -2672
rect 1583 -2678 1586 -2672
rect 1590 -2678 1593 -2672
rect 1597 -2678 1600 -2672
rect 1604 -2678 1607 -2672
rect 1611 -2678 1614 -2672
rect 1618 -2678 1621 -2672
rect 1625 -2678 1628 -2672
rect 1632 -2678 1635 -2672
rect 1639 -2678 1642 -2672
rect 1646 -2678 1649 -2672
rect 1653 -2678 1656 -2672
rect 1660 -2678 1663 -2672
rect 1667 -2678 1670 -2672
rect 1674 -2678 1677 -2672
rect 1681 -2678 1684 -2672
rect 1688 -2678 1691 -2672
rect 1695 -2678 1698 -2672
rect 1702 -2678 1705 -2672
rect 1709 -2678 1712 -2672
rect 1716 -2678 1719 -2672
rect 1723 -2678 1726 -2672
rect 1730 -2678 1733 -2672
rect 1737 -2678 1740 -2672
rect 1744 -2678 1747 -2672
rect 1751 -2678 1757 -2672
rect 1758 -2678 1761 -2672
rect 1765 -2678 1768 -2672
rect 1772 -2678 1775 -2672
rect 1779 -2678 1782 -2672
rect 1786 -2678 1789 -2672
rect 1793 -2678 1796 -2672
rect 1800 -2678 1803 -2672
rect 1807 -2678 1810 -2672
rect 1814 -2678 1817 -2672
rect 1821 -2678 1824 -2672
rect 1828 -2678 1831 -2672
rect 1835 -2678 1838 -2672
rect 1842 -2678 1845 -2672
rect 1849 -2678 1852 -2672
rect 1856 -2678 1859 -2672
rect 1863 -2678 1866 -2672
rect 1870 -2678 1873 -2672
rect 1877 -2678 1880 -2672
rect 1884 -2678 1887 -2672
rect 1891 -2678 1894 -2672
rect 1898 -2678 1901 -2672
rect 1905 -2678 1908 -2672
rect 1912 -2678 1915 -2672
rect 1919 -2678 1922 -2672
rect 1926 -2678 1929 -2672
rect 1933 -2678 1936 -2672
rect 1940 -2678 1943 -2672
rect 1947 -2678 1950 -2672
rect 1954 -2678 1957 -2672
rect 1961 -2678 1964 -2672
rect 1968 -2678 1971 -2672
rect 1975 -2678 1978 -2672
rect 1982 -2678 1985 -2672
rect 1989 -2678 1992 -2672
rect 1996 -2678 1999 -2672
rect 2003 -2678 2006 -2672
rect 2010 -2678 2013 -2672
rect 2017 -2678 2020 -2672
rect 2024 -2678 2027 -2672
rect 2031 -2678 2034 -2672
rect 2038 -2678 2041 -2672
rect 2045 -2678 2048 -2672
rect 2052 -2678 2055 -2672
rect 2059 -2678 2062 -2672
rect 2066 -2678 2069 -2672
rect 2073 -2678 2076 -2672
rect 2080 -2678 2083 -2672
rect 2087 -2678 2090 -2672
rect 2094 -2678 2097 -2672
rect 2101 -2678 2104 -2672
rect 2108 -2678 2111 -2672
rect 2115 -2678 2118 -2672
rect 2122 -2678 2125 -2672
rect 2129 -2678 2132 -2672
rect 2136 -2678 2139 -2672
rect 2143 -2678 2146 -2672
rect 2150 -2678 2153 -2672
rect 2157 -2678 2160 -2672
rect 2164 -2678 2167 -2672
rect 2171 -2678 2174 -2672
rect 2178 -2678 2181 -2672
rect 2185 -2678 2188 -2672
rect 2192 -2678 2195 -2672
rect 2199 -2678 2202 -2672
rect 2206 -2678 2209 -2672
rect 2213 -2678 2216 -2672
rect 2220 -2678 2223 -2672
rect 2227 -2678 2230 -2672
rect 2234 -2678 2237 -2672
rect 2241 -2678 2244 -2672
rect 2262 -2678 2265 -2672
rect 2269 -2678 2272 -2672
rect 1 -2841 4 -2835
rect 8 -2841 11 -2835
rect 15 -2841 18 -2835
rect 22 -2841 25 -2835
rect 29 -2841 32 -2835
rect 36 -2841 39 -2835
rect 43 -2841 46 -2835
rect 50 -2841 56 -2835
rect 57 -2841 60 -2835
rect 64 -2841 67 -2835
rect 71 -2841 74 -2835
rect 78 -2841 84 -2835
rect 85 -2841 88 -2835
rect 92 -2841 95 -2835
rect 99 -2841 102 -2835
rect 106 -2841 112 -2835
rect 113 -2841 116 -2835
rect 120 -2841 123 -2835
rect 127 -2841 130 -2835
rect 134 -2841 137 -2835
rect 141 -2841 144 -2835
rect 148 -2841 151 -2835
rect 155 -2841 158 -2835
rect 162 -2841 165 -2835
rect 169 -2841 172 -2835
rect 176 -2841 179 -2835
rect 183 -2841 186 -2835
rect 190 -2841 193 -2835
rect 197 -2841 200 -2835
rect 204 -2841 207 -2835
rect 211 -2841 214 -2835
rect 218 -2841 224 -2835
rect 225 -2841 228 -2835
rect 232 -2841 238 -2835
rect 239 -2841 242 -2835
rect 246 -2841 252 -2835
rect 253 -2841 256 -2835
rect 260 -2841 263 -2835
rect 267 -2841 270 -2835
rect 274 -2841 277 -2835
rect 281 -2841 284 -2835
rect 288 -2841 291 -2835
rect 295 -2841 298 -2835
rect 302 -2841 305 -2835
rect 309 -2841 312 -2835
rect 316 -2841 319 -2835
rect 323 -2841 326 -2835
rect 330 -2841 333 -2835
rect 337 -2841 340 -2835
rect 344 -2841 347 -2835
rect 351 -2841 354 -2835
rect 358 -2841 361 -2835
rect 365 -2841 368 -2835
rect 372 -2841 375 -2835
rect 379 -2841 382 -2835
rect 386 -2841 389 -2835
rect 393 -2841 396 -2835
rect 400 -2841 403 -2835
rect 407 -2841 410 -2835
rect 414 -2841 417 -2835
rect 421 -2841 424 -2835
rect 428 -2841 434 -2835
rect 435 -2841 438 -2835
rect 442 -2841 445 -2835
rect 449 -2841 452 -2835
rect 456 -2841 462 -2835
rect 463 -2841 466 -2835
rect 470 -2841 473 -2835
rect 477 -2841 480 -2835
rect 484 -2841 487 -2835
rect 491 -2841 494 -2835
rect 498 -2841 501 -2835
rect 505 -2841 508 -2835
rect 512 -2841 515 -2835
rect 519 -2841 522 -2835
rect 526 -2841 529 -2835
rect 533 -2841 536 -2835
rect 540 -2841 546 -2835
rect 547 -2841 550 -2835
rect 554 -2841 557 -2835
rect 561 -2841 564 -2835
rect 568 -2841 571 -2835
rect 575 -2841 578 -2835
rect 582 -2841 585 -2835
rect 589 -2841 592 -2835
rect 596 -2841 599 -2835
rect 603 -2841 606 -2835
rect 610 -2841 613 -2835
rect 617 -2841 623 -2835
rect 624 -2841 627 -2835
rect 631 -2841 634 -2835
rect 638 -2841 641 -2835
rect 645 -2841 648 -2835
rect 652 -2841 655 -2835
rect 659 -2841 665 -2835
rect 666 -2841 669 -2835
rect 673 -2841 676 -2835
rect 680 -2841 683 -2835
rect 687 -2841 690 -2835
rect 694 -2841 697 -2835
rect 701 -2841 707 -2835
rect 708 -2841 711 -2835
rect 715 -2841 718 -2835
rect 722 -2841 725 -2835
rect 729 -2841 735 -2835
rect 736 -2841 739 -2835
rect 743 -2841 749 -2835
rect 750 -2841 753 -2835
rect 757 -2841 760 -2835
rect 764 -2841 767 -2835
rect 771 -2841 774 -2835
rect 778 -2841 781 -2835
rect 785 -2841 791 -2835
rect 792 -2841 795 -2835
rect 799 -2841 802 -2835
rect 806 -2841 809 -2835
rect 813 -2841 816 -2835
rect 820 -2841 823 -2835
rect 827 -2841 830 -2835
rect 834 -2841 840 -2835
rect 841 -2841 844 -2835
rect 848 -2841 851 -2835
rect 855 -2841 858 -2835
rect 862 -2841 868 -2835
rect 869 -2841 872 -2835
rect 876 -2841 879 -2835
rect 883 -2841 886 -2835
rect 890 -2841 893 -2835
rect 897 -2841 900 -2835
rect 904 -2841 907 -2835
rect 911 -2841 917 -2835
rect 918 -2841 921 -2835
rect 925 -2841 928 -2835
rect 932 -2841 935 -2835
rect 939 -2841 945 -2835
rect 946 -2841 949 -2835
rect 953 -2841 956 -2835
rect 960 -2841 966 -2835
rect 967 -2841 970 -2835
rect 974 -2841 980 -2835
rect 981 -2841 984 -2835
rect 988 -2841 991 -2835
rect 995 -2841 998 -2835
rect 1002 -2841 1005 -2835
rect 1009 -2841 1012 -2835
rect 1016 -2841 1019 -2835
rect 1023 -2841 1026 -2835
rect 1030 -2841 1033 -2835
rect 1037 -2841 1040 -2835
rect 1044 -2841 1047 -2835
rect 1051 -2841 1057 -2835
rect 1058 -2841 1064 -2835
rect 1065 -2841 1068 -2835
rect 1072 -2841 1075 -2835
rect 1079 -2841 1082 -2835
rect 1086 -2841 1089 -2835
rect 1093 -2841 1099 -2835
rect 1100 -2841 1103 -2835
rect 1107 -2841 1110 -2835
rect 1114 -2841 1117 -2835
rect 1121 -2841 1124 -2835
rect 1128 -2841 1131 -2835
rect 1135 -2841 1138 -2835
rect 1142 -2841 1145 -2835
rect 1149 -2841 1152 -2835
rect 1156 -2841 1159 -2835
rect 1163 -2841 1166 -2835
rect 1170 -2841 1173 -2835
rect 1177 -2841 1180 -2835
rect 1184 -2841 1187 -2835
rect 1191 -2841 1194 -2835
rect 1198 -2841 1201 -2835
rect 1205 -2841 1208 -2835
rect 1212 -2841 1215 -2835
rect 1219 -2841 1222 -2835
rect 1226 -2841 1229 -2835
rect 1233 -2841 1236 -2835
rect 1240 -2841 1243 -2835
rect 1247 -2841 1250 -2835
rect 1254 -2841 1260 -2835
rect 1261 -2841 1264 -2835
rect 1268 -2841 1271 -2835
rect 1275 -2841 1278 -2835
rect 1282 -2841 1288 -2835
rect 1289 -2841 1292 -2835
rect 1296 -2841 1299 -2835
rect 1303 -2841 1306 -2835
rect 1310 -2841 1316 -2835
rect 1317 -2841 1320 -2835
rect 1324 -2841 1327 -2835
rect 1331 -2841 1334 -2835
rect 1338 -2841 1341 -2835
rect 1345 -2841 1351 -2835
rect 1352 -2841 1355 -2835
rect 1359 -2841 1362 -2835
rect 1366 -2841 1369 -2835
rect 1373 -2841 1376 -2835
rect 1380 -2841 1383 -2835
rect 1387 -2841 1393 -2835
rect 1394 -2841 1397 -2835
rect 1401 -2841 1404 -2835
rect 1408 -2841 1411 -2835
rect 1415 -2841 1418 -2835
rect 1422 -2841 1425 -2835
rect 1429 -2841 1435 -2835
rect 1436 -2841 1439 -2835
rect 1443 -2841 1446 -2835
rect 1450 -2841 1456 -2835
rect 1457 -2841 1460 -2835
rect 1464 -2841 1467 -2835
rect 1471 -2841 1474 -2835
rect 1478 -2841 1481 -2835
rect 1485 -2841 1491 -2835
rect 1492 -2841 1498 -2835
rect 1499 -2841 1502 -2835
rect 1506 -2841 1509 -2835
rect 1513 -2841 1516 -2835
rect 1520 -2841 1523 -2835
rect 1527 -2841 1530 -2835
rect 1534 -2841 1537 -2835
rect 1541 -2841 1544 -2835
rect 1548 -2841 1551 -2835
rect 1555 -2841 1558 -2835
rect 1562 -2841 1568 -2835
rect 1569 -2841 1572 -2835
rect 1576 -2841 1579 -2835
rect 1583 -2841 1586 -2835
rect 1590 -2841 1593 -2835
rect 1597 -2841 1600 -2835
rect 1604 -2841 1607 -2835
rect 1611 -2841 1614 -2835
rect 1618 -2841 1621 -2835
rect 1625 -2841 1628 -2835
rect 1632 -2841 1635 -2835
rect 1639 -2841 1642 -2835
rect 1646 -2841 1649 -2835
rect 1653 -2841 1656 -2835
rect 1660 -2841 1663 -2835
rect 1667 -2841 1670 -2835
rect 1674 -2841 1677 -2835
rect 1681 -2841 1687 -2835
rect 1688 -2841 1691 -2835
rect 1695 -2841 1698 -2835
rect 1702 -2841 1708 -2835
rect 1709 -2841 1712 -2835
rect 1716 -2841 1719 -2835
rect 1723 -2841 1726 -2835
rect 1730 -2841 1733 -2835
rect 1737 -2841 1740 -2835
rect 1744 -2841 1747 -2835
rect 1751 -2841 1757 -2835
rect 1758 -2841 1761 -2835
rect 1765 -2841 1768 -2835
rect 1772 -2841 1775 -2835
rect 1779 -2841 1782 -2835
rect 1786 -2841 1789 -2835
rect 1793 -2841 1796 -2835
rect 1800 -2841 1803 -2835
rect 1807 -2841 1810 -2835
rect 1814 -2841 1817 -2835
rect 1821 -2841 1824 -2835
rect 1828 -2841 1831 -2835
rect 1835 -2841 1838 -2835
rect 1842 -2841 1845 -2835
rect 1849 -2841 1852 -2835
rect 1856 -2841 1859 -2835
rect 1863 -2841 1866 -2835
rect 1870 -2841 1873 -2835
rect 1877 -2841 1880 -2835
rect 1884 -2841 1887 -2835
rect 1891 -2841 1894 -2835
rect 1898 -2841 1901 -2835
rect 1905 -2841 1908 -2835
rect 1912 -2841 1915 -2835
rect 1919 -2841 1922 -2835
rect 1926 -2841 1929 -2835
rect 1933 -2841 1936 -2835
rect 1940 -2841 1943 -2835
rect 1947 -2841 1950 -2835
rect 1954 -2841 1957 -2835
rect 1961 -2841 1964 -2835
rect 1968 -2841 1971 -2835
rect 1975 -2841 1978 -2835
rect 1982 -2841 1985 -2835
rect 1989 -2841 1992 -2835
rect 1996 -2841 1999 -2835
rect 2003 -2841 2006 -2835
rect 2010 -2841 2013 -2835
rect 2017 -2841 2020 -2835
rect 2024 -2841 2027 -2835
rect 2031 -2841 2034 -2835
rect 2038 -2841 2041 -2835
rect 2045 -2841 2048 -2835
rect 2052 -2841 2055 -2835
rect 2059 -2841 2062 -2835
rect 2066 -2841 2069 -2835
rect 2073 -2841 2076 -2835
rect 2080 -2841 2083 -2835
rect 2087 -2841 2090 -2835
rect 2094 -2841 2097 -2835
rect 2101 -2841 2104 -2835
rect 2108 -2841 2111 -2835
rect 2115 -2841 2118 -2835
rect 2122 -2841 2125 -2835
rect 2129 -2841 2132 -2835
rect 2136 -2841 2139 -2835
rect 2143 -2841 2146 -2835
rect 2150 -2841 2153 -2835
rect 2157 -2841 2160 -2835
rect 2164 -2841 2167 -2835
rect 2171 -2841 2174 -2835
rect 2178 -2841 2181 -2835
rect 2185 -2841 2188 -2835
rect 2192 -2841 2195 -2835
rect 2199 -2841 2202 -2835
rect 2206 -2841 2209 -2835
rect 2213 -2841 2216 -2835
rect 2220 -2841 2226 -2835
rect 2227 -2841 2230 -2835
rect 2234 -2841 2237 -2835
rect 2241 -2841 2244 -2835
rect 2248 -2841 2251 -2835
rect 2255 -2841 2261 -2835
rect 2262 -2841 2265 -2835
rect 2269 -2841 2272 -2835
rect 1 -2986 7 -2980
rect 8 -2986 14 -2980
rect 15 -2986 18 -2980
rect 22 -2986 25 -2980
rect 29 -2986 32 -2980
rect 36 -2986 39 -2980
rect 43 -2986 46 -2980
rect 50 -2986 56 -2980
rect 57 -2986 60 -2980
rect 64 -2986 67 -2980
rect 71 -2986 74 -2980
rect 78 -2986 81 -2980
rect 85 -2986 88 -2980
rect 92 -2986 95 -2980
rect 99 -2986 105 -2980
rect 106 -2986 112 -2980
rect 113 -2986 119 -2980
rect 120 -2986 126 -2980
rect 127 -2986 130 -2980
rect 134 -2986 137 -2980
rect 141 -2986 144 -2980
rect 148 -2986 151 -2980
rect 155 -2986 161 -2980
rect 162 -2986 165 -2980
rect 169 -2986 172 -2980
rect 176 -2986 179 -2980
rect 183 -2986 186 -2980
rect 190 -2986 193 -2980
rect 197 -2986 200 -2980
rect 204 -2986 207 -2980
rect 211 -2986 217 -2980
rect 218 -2986 221 -2980
rect 225 -2986 228 -2980
rect 232 -2986 235 -2980
rect 239 -2986 242 -2980
rect 246 -2986 249 -2980
rect 253 -2986 259 -2980
rect 260 -2986 263 -2980
rect 267 -2986 270 -2980
rect 274 -2986 277 -2980
rect 281 -2986 284 -2980
rect 288 -2986 291 -2980
rect 295 -2986 298 -2980
rect 302 -2986 305 -2980
rect 309 -2986 312 -2980
rect 316 -2986 319 -2980
rect 323 -2986 326 -2980
rect 330 -2986 333 -2980
rect 337 -2986 340 -2980
rect 344 -2986 347 -2980
rect 351 -2986 354 -2980
rect 358 -2986 361 -2980
rect 365 -2986 368 -2980
rect 372 -2986 375 -2980
rect 379 -2986 382 -2980
rect 386 -2986 389 -2980
rect 393 -2986 396 -2980
rect 400 -2986 403 -2980
rect 407 -2986 410 -2980
rect 414 -2986 417 -2980
rect 421 -2986 424 -2980
rect 428 -2986 431 -2980
rect 435 -2986 438 -2980
rect 442 -2986 445 -2980
rect 449 -2986 452 -2980
rect 456 -2986 459 -2980
rect 463 -2986 469 -2980
rect 470 -2986 473 -2980
rect 477 -2986 480 -2980
rect 484 -2986 487 -2980
rect 491 -2986 494 -2980
rect 498 -2986 501 -2980
rect 505 -2986 508 -2980
rect 512 -2986 515 -2980
rect 519 -2986 522 -2980
rect 526 -2986 529 -2980
rect 533 -2986 536 -2980
rect 540 -2986 546 -2980
rect 547 -2986 550 -2980
rect 554 -2986 557 -2980
rect 561 -2986 567 -2980
rect 568 -2986 574 -2980
rect 575 -2986 578 -2980
rect 582 -2986 585 -2980
rect 589 -2986 592 -2980
rect 596 -2986 599 -2980
rect 603 -2986 606 -2980
rect 610 -2986 613 -2980
rect 617 -2986 620 -2980
rect 624 -2986 627 -2980
rect 631 -2986 634 -2980
rect 638 -2986 644 -2980
rect 645 -2986 648 -2980
rect 652 -2986 655 -2980
rect 659 -2986 665 -2980
rect 666 -2986 669 -2980
rect 673 -2986 676 -2980
rect 680 -2986 683 -2980
rect 687 -2986 690 -2980
rect 694 -2986 697 -2980
rect 701 -2986 704 -2980
rect 708 -2986 711 -2980
rect 715 -2986 718 -2980
rect 722 -2986 725 -2980
rect 729 -2986 732 -2980
rect 736 -2986 742 -2980
rect 743 -2986 746 -2980
rect 750 -2986 753 -2980
rect 757 -2986 760 -2980
rect 764 -2986 767 -2980
rect 771 -2986 774 -2980
rect 778 -2986 781 -2980
rect 785 -2986 788 -2980
rect 792 -2986 795 -2980
rect 799 -2986 802 -2980
rect 806 -2986 809 -2980
rect 813 -2986 816 -2980
rect 820 -2986 823 -2980
rect 827 -2986 830 -2980
rect 834 -2986 837 -2980
rect 841 -2986 844 -2980
rect 848 -2986 851 -2980
rect 855 -2986 858 -2980
rect 862 -2986 865 -2980
rect 869 -2986 872 -2980
rect 876 -2986 882 -2980
rect 883 -2986 886 -2980
rect 890 -2986 893 -2980
rect 897 -2986 900 -2980
rect 904 -2986 907 -2980
rect 911 -2986 917 -2980
rect 918 -2986 924 -2980
rect 925 -2986 928 -2980
rect 932 -2986 935 -2980
rect 939 -2986 942 -2980
rect 946 -2986 949 -2980
rect 953 -2986 956 -2980
rect 960 -2986 966 -2980
rect 967 -2986 970 -2980
rect 974 -2986 977 -2980
rect 981 -2986 987 -2980
rect 988 -2986 991 -2980
rect 995 -2986 998 -2980
rect 1002 -2986 1005 -2980
rect 1009 -2986 1012 -2980
rect 1016 -2986 1019 -2980
rect 1023 -2986 1026 -2980
rect 1030 -2986 1036 -2980
rect 1037 -2986 1043 -2980
rect 1044 -2986 1047 -2980
rect 1051 -2986 1057 -2980
rect 1058 -2986 1064 -2980
rect 1065 -2986 1071 -2980
rect 1072 -2986 1075 -2980
rect 1079 -2986 1082 -2980
rect 1086 -2986 1089 -2980
rect 1093 -2986 1099 -2980
rect 1100 -2986 1103 -2980
rect 1107 -2986 1110 -2980
rect 1114 -2986 1117 -2980
rect 1121 -2986 1127 -2980
rect 1128 -2986 1131 -2980
rect 1135 -2986 1141 -2980
rect 1142 -2986 1145 -2980
rect 1149 -2986 1152 -2980
rect 1156 -2986 1162 -2980
rect 1163 -2986 1166 -2980
rect 1170 -2986 1173 -2980
rect 1177 -2986 1180 -2980
rect 1184 -2986 1187 -2980
rect 1191 -2986 1194 -2980
rect 1198 -2986 1204 -2980
rect 1205 -2986 1211 -2980
rect 1212 -2986 1215 -2980
rect 1219 -2986 1222 -2980
rect 1226 -2986 1229 -2980
rect 1233 -2986 1236 -2980
rect 1240 -2986 1243 -2980
rect 1247 -2986 1250 -2980
rect 1254 -2986 1257 -2980
rect 1261 -2986 1264 -2980
rect 1268 -2986 1271 -2980
rect 1275 -2986 1278 -2980
rect 1282 -2986 1285 -2980
rect 1289 -2986 1292 -2980
rect 1296 -2986 1299 -2980
rect 1303 -2986 1306 -2980
rect 1310 -2986 1316 -2980
rect 1317 -2986 1320 -2980
rect 1324 -2986 1327 -2980
rect 1331 -2986 1334 -2980
rect 1338 -2986 1341 -2980
rect 1345 -2986 1348 -2980
rect 1352 -2986 1355 -2980
rect 1359 -2986 1365 -2980
rect 1366 -2986 1369 -2980
rect 1373 -2986 1376 -2980
rect 1380 -2986 1383 -2980
rect 1387 -2986 1390 -2980
rect 1394 -2986 1397 -2980
rect 1401 -2986 1404 -2980
rect 1408 -2986 1411 -2980
rect 1415 -2986 1421 -2980
rect 1422 -2986 1425 -2980
rect 1429 -2986 1432 -2980
rect 1436 -2986 1439 -2980
rect 1443 -2986 1446 -2980
rect 1450 -2986 1453 -2980
rect 1457 -2986 1460 -2980
rect 1464 -2986 1467 -2980
rect 1471 -2986 1474 -2980
rect 1478 -2986 1481 -2980
rect 1485 -2986 1488 -2980
rect 1492 -2986 1495 -2980
rect 1499 -2986 1502 -2980
rect 1506 -2986 1509 -2980
rect 1513 -2986 1516 -2980
rect 1520 -2986 1523 -2980
rect 1527 -2986 1530 -2980
rect 1534 -2986 1537 -2980
rect 1541 -2986 1544 -2980
rect 1548 -2986 1551 -2980
rect 1555 -2986 1558 -2980
rect 1562 -2986 1565 -2980
rect 1569 -2986 1575 -2980
rect 1576 -2986 1579 -2980
rect 1583 -2986 1586 -2980
rect 1590 -2986 1593 -2980
rect 1597 -2986 1600 -2980
rect 1604 -2986 1607 -2980
rect 1611 -2986 1614 -2980
rect 1618 -2986 1621 -2980
rect 1625 -2986 1628 -2980
rect 1632 -2986 1635 -2980
rect 1639 -2986 1642 -2980
rect 1646 -2986 1649 -2980
rect 1653 -2986 1656 -2980
rect 1660 -2986 1663 -2980
rect 1667 -2986 1670 -2980
rect 1674 -2986 1677 -2980
rect 1681 -2986 1684 -2980
rect 1688 -2986 1691 -2980
rect 1695 -2986 1698 -2980
rect 1702 -2986 1705 -2980
rect 1709 -2986 1712 -2980
rect 1716 -2986 1719 -2980
rect 1723 -2986 1726 -2980
rect 1730 -2986 1733 -2980
rect 1737 -2986 1740 -2980
rect 1744 -2986 1747 -2980
rect 1751 -2986 1754 -2980
rect 1758 -2986 1761 -2980
rect 1765 -2986 1771 -2980
rect 1772 -2986 1775 -2980
rect 1779 -2986 1782 -2980
rect 1786 -2986 1789 -2980
rect 1793 -2986 1796 -2980
rect 1800 -2986 1803 -2980
rect 1807 -2986 1810 -2980
rect 1814 -2986 1817 -2980
rect 1821 -2986 1824 -2980
rect 1828 -2986 1831 -2980
rect 1835 -2986 1838 -2980
rect 1842 -2986 1845 -2980
rect 1849 -2986 1852 -2980
rect 1856 -2986 1859 -2980
rect 1863 -2986 1866 -2980
rect 1870 -2986 1873 -2980
rect 1877 -2986 1880 -2980
rect 1884 -2986 1887 -2980
rect 1891 -2986 1894 -2980
rect 1898 -2986 1901 -2980
rect 1905 -2986 1908 -2980
rect 1912 -2986 1915 -2980
rect 1919 -2986 1922 -2980
rect 1926 -2986 1929 -2980
rect 1933 -2986 1936 -2980
rect 1940 -2986 1943 -2980
rect 1947 -2986 1950 -2980
rect 1954 -2986 1957 -2980
rect 1961 -2986 1964 -2980
rect 1968 -2986 1971 -2980
rect 1975 -2986 1978 -2980
rect 1982 -2986 1985 -2980
rect 1989 -2986 1992 -2980
rect 1996 -2986 1999 -2980
rect 2003 -2986 2006 -2980
rect 2010 -2986 2013 -2980
rect 2017 -2986 2020 -2980
rect 2024 -2986 2027 -2980
rect 2031 -2986 2034 -2980
rect 2038 -2986 2041 -2980
rect 2045 -2986 2048 -2980
rect 2052 -2986 2055 -2980
rect 2059 -2986 2062 -2980
rect 2066 -2986 2069 -2980
rect 2073 -2986 2076 -2980
rect 2080 -2986 2083 -2980
rect 2087 -2986 2090 -2980
rect 2094 -2986 2100 -2980
rect 2101 -2986 2104 -2980
rect 2108 -2986 2111 -2980
rect 2115 -2986 2118 -2980
rect 2122 -2986 2125 -2980
rect 2129 -2986 2132 -2980
rect 2136 -2986 2139 -2980
rect 2143 -2986 2146 -2980
rect 2150 -2986 2153 -2980
rect 1 -3101 7 -3095
rect 8 -3101 14 -3095
rect 15 -3101 21 -3095
rect 22 -3101 25 -3095
rect 29 -3101 32 -3095
rect 36 -3101 39 -3095
rect 43 -3101 49 -3095
rect 50 -3101 56 -3095
rect 57 -3101 60 -3095
rect 64 -3101 67 -3095
rect 71 -3101 74 -3095
rect 78 -3101 84 -3095
rect 85 -3101 88 -3095
rect 92 -3101 98 -3095
rect 99 -3101 102 -3095
rect 106 -3101 109 -3095
rect 113 -3101 116 -3095
rect 120 -3101 123 -3095
rect 127 -3101 133 -3095
rect 134 -3101 140 -3095
rect 141 -3101 144 -3095
rect 148 -3101 151 -3095
rect 155 -3101 158 -3095
rect 162 -3101 168 -3095
rect 169 -3101 175 -3095
rect 176 -3101 179 -3095
rect 183 -3101 186 -3095
rect 190 -3101 193 -3095
rect 197 -3101 200 -3095
rect 204 -3101 210 -3095
rect 211 -3101 214 -3095
rect 218 -3101 221 -3095
rect 225 -3101 228 -3095
rect 232 -3101 238 -3095
rect 239 -3101 242 -3095
rect 246 -3101 249 -3095
rect 253 -3101 256 -3095
rect 260 -3101 263 -3095
rect 267 -3101 270 -3095
rect 274 -3101 277 -3095
rect 281 -3101 284 -3095
rect 288 -3101 291 -3095
rect 295 -3101 298 -3095
rect 302 -3101 305 -3095
rect 309 -3101 312 -3095
rect 316 -3101 319 -3095
rect 323 -3101 326 -3095
rect 330 -3101 333 -3095
rect 337 -3101 340 -3095
rect 344 -3101 347 -3095
rect 351 -3101 354 -3095
rect 358 -3101 361 -3095
rect 365 -3101 368 -3095
rect 372 -3101 375 -3095
rect 379 -3101 382 -3095
rect 386 -3101 389 -3095
rect 393 -3101 396 -3095
rect 400 -3101 403 -3095
rect 407 -3101 410 -3095
rect 414 -3101 417 -3095
rect 421 -3101 424 -3095
rect 428 -3101 431 -3095
rect 435 -3101 438 -3095
rect 442 -3101 445 -3095
rect 449 -3101 452 -3095
rect 456 -3101 462 -3095
rect 463 -3101 466 -3095
rect 470 -3101 473 -3095
rect 477 -3101 480 -3095
rect 484 -3101 487 -3095
rect 491 -3101 494 -3095
rect 498 -3101 501 -3095
rect 505 -3101 508 -3095
rect 512 -3101 515 -3095
rect 519 -3101 522 -3095
rect 526 -3101 532 -3095
rect 533 -3101 536 -3095
rect 540 -3101 543 -3095
rect 547 -3101 550 -3095
rect 554 -3101 557 -3095
rect 561 -3101 564 -3095
rect 568 -3101 571 -3095
rect 575 -3101 578 -3095
rect 582 -3101 585 -3095
rect 589 -3101 592 -3095
rect 596 -3101 599 -3095
rect 603 -3101 606 -3095
rect 610 -3101 616 -3095
rect 617 -3101 620 -3095
rect 624 -3101 627 -3095
rect 631 -3101 634 -3095
rect 638 -3101 641 -3095
rect 645 -3101 648 -3095
rect 652 -3101 655 -3095
rect 659 -3101 662 -3095
rect 666 -3101 669 -3095
rect 673 -3101 676 -3095
rect 680 -3101 683 -3095
rect 687 -3101 690 -3095
rect 694 -3101 697 -3095
rect 701 -3101 704 -3095
rect 708 -3101 711 -3095
rect 715 -3101 718 -3095
rect 722 -3101 725 -3095
rect 729 -3101 732 -3095
rect 736 -3101 739 -3095
rect 743 -3101 746 -3095
rect 750 -3101 753 -3095
rect 757 -3101 760 -3095
rect 764 -3101 767 -3095
rect 771 -3101 774 -3095
rect 778 -3101 781 -3095
rect 785 -3101 788 -3095
rect 792 -3101 795 -3095
rect 799 -3101 802 -3095
rect 806 -3101 809 -3095
rect 813 -3101 819 -3095
rect 820 -3101 823 -3095
rect 827 -3101 830 -3095
rect 834 -3101 837 -3095
rect 841 -3101 844 -3095
rect 848 -3101 851 -3095
rect 855 -3101 858 -3095
rect 862 -3101 868 -3095
rect 869 -3101 872 -3095
rect 876 -3101 882 -3095
rect 883 -3101 886 -3095
rect 890 -3101 896 -3095
rect 897 -3101 900 -3095
rect 904 -3101 907 -3095
rect 911 -3101 917 -3095
rect 918 -3101 921 -3095
rect 925 -3101 928 -3095
rect 932 -3101 935 -3095
rect 939 -3101 942 -3095
rect 946 -3101 949 -3095
rect 953 -3101 956 -3095
rect 960 -3101 963 -3095
rect 967 -3101 970 -3095
rect 974 -3101 977 -3095
rect 981 -3101 984 -3095
rect 988 -3101 991 -3095
rect 995 -3101 998 -3095
rect 1002 -3101 1005 -3095
rect 1009 -3101 1012 -3095
rect 1016 -3101 1019 -3095
rect 1023 -3101 1026 -3095
rect 1030 -3101 1033 -3095
rect 1037 -3101 1040 -3095
rect 1044 -3101 1047 -3095
rect 1051 -3101 1057 -3095
rect 1058 -3101 1061 -3095
rect 1065 -3101 1068 -3095
rect 1072 -3101 1078 -3095
rect 1079 -3101 1085 -3095
rect 1086 -3101 1089 -3095
rect 1093 -3101 1096 -3095
rect 1100 -3101 1103 -3095
rect 1107 -3101 1110 -3095
rect 1114 -3101 1117 -3095
rect 1121 -3101 1127 -3095
rect 1128 -3101 1131 -3095
rect 1135 -3101 1138 -3095
rect 1142 -3101 1145 -3095
rect 1149 -3101 1152 -3095
rect 1156 -3101 1162 -3095
rect 1163 -3101 1166 -3095
rect 1170 -3101 1173 -3095
rect 1177 -3101 1180 -3095
rect 1184 -3101 1187 -3095
rect 1191 -3101 1194 -3095
rect 1198 -3101 1201 -3095
rect 1205 -3101 1208 -3095
rect 1212 -3101 1218 -3095
rect 1219 -3101 1222 -3095
rect 1226 -3101 1229 -3095
rect 1233 -3101 1239 -3095
rect 1240 -3101 1243 -3095
rect 1247 -3101 1253 -3095
rect 1254 -3101 1257 -3095
rect 1261 -3101 1264 -3095
rect 1268 -3101 1271 -3095
rect 1275 -3101 1281 -3095
rect 1282 -3101 1285 -3095
rect 1289 -3101 1292 -3095
rect 1296 -3101 1299 -3095
rect 1303 -3101 1306 -3095
rect 1310 -3101 1316 -3095
rect 1317 -3101 1320 -3095
rect 1324 -3101 1327 -3095
rect 1331 -3101 1334 -3095
rect 1338 -3101 1341 -3095
rect 1345 -3101 1348 -3095
rect 1352 -3101 1355 -3095
rect 1359 -3101 1362 -3095
rect 1366 -3101 1369 -3095
rect 1373 -3101 1376 -3095
rect 1380 -3101 1383 -3095
rect 1387 -3101 1390 -3095
rect 1394 -3101 1400 -3095
rect 1401 -3101 1407 -3095
rect 1408 -3101 1411 -3095
rect 1415 -3101 1418 -3095
rect 1422 -3101 1425 -3095
rect 1429 -3101 1432 -3095
rect 1436 -3101 1439 -3095
rect 1443 -3101 1449 -3095
rect 1450 -3101 1453 -3095
rect 1457 -3101 1460 -3095
rect 1464 -3101 1467 -3095
rect 1471 -3101 1474 -3095
rect 1478 -3101 1481 -3095
rect 1485 -3101 1488 -3095
rect 1492 -3101 1495 -3095
rect 1499 -3101 1502 -3095
rect 1506 -3101 1509 -3095
rect 1513 -3101 1516 -3095
rect 1520 -3101 1523 -3095
rect 1527 -3101 1530 -3095
rect 1534 -3101 1537 -3095
rect 1541 -3101 1544 -3095
rect 1548 -3101 1551 -3095
rect 1555 -3101 1561 -3095
rect 1562 -3101 1568 -3095
rect 1569 -3101 1572 -3095
rect 1576 -3101 1579 -3095
rect 1583 -3101 1586 -3095
rect 1590 -3101 1593 -3095
rect 1597 -3101 1600 -3095
rect 1604 -3101 1607 -3095
rect 1611 -3101 1614 -3095
rect 1618 -3101 1621 -3095
rect 1625 -3101 1628 -3095
rect 1632 -3101 1635 -3095
rect 1639 -3101 1642 -3095
rect 1646 -3101 1649 -3095
rect 1653 -3101 1656 -3095
rect 1660 -3101 1663 -3095
rect 1667 -3101 1670 -3095
rect 1674 -3101 1677 -3095
rect 1681 -3101 1687 -3095
rect 1688 -3101 1691 -3095
rect 1695 -3101 1698 -3095
rect 1702 -3101 1705 -3095
rect 1709 -3101 1712 -3095
rect 1716 -3101 1719 -3095
rect 1723 -3101 1726 -3095
rect 1730 -3101 1733 -3095
rect 1737 -3101 1740 -3095
rect 1744 -3101 1747 -3095
rect 1751 -3101 1754 -3095
rect 1758 -3101 1761 -3095
rect 1765 -3101 1768 -3095
rect 1772 -3101 1775 -3095
rect 1779 -3101 1782 -3095
rect 1786 -3101 1789 -3095
rect 1793 -3101 1796 -3095
rect 1800 -3101 1803 -3095
rect 1807 -3101 1810 -3095
rect 1814 -3101 1817 -3095
rect 1821 -3101 1824 -3095
rect 1828 -3101 1831 -3095
rect 1835 -3101 1838 -3095
rect 1842 -3101 1845 -3095
rect 1849 -3101 1852 -3095
rect 1856 -3101 1859 -3095
rect 1863 -3101 1866 -3095
rect 1870 -3101 1873 -3095
rect 1877 -3101 1883 -3095
rect 1884 -3101 1887 -3095
rect 1891 -3101 1894 -3095
rect 1898 -3101 1901 -3095
rect 1905 -3101 1908 -3095
rect 1912 -3101 1915 -3095
rect 1919 -3101 1922 -3095
rect 1926 -3101 1929 -3095
rect 1933 -3101 1936 -3095
rect 1940 -3101 1943 -3095
rect 1947 -3101 1950 -3095
rect 1954 -3101 1957 -3095
rect 1961 -3101 1967 -3095
rect 1968 -3101 1971 -3095
rect 1975 -3101 1978 -3095
rect 1982 -3101 1985 -3095
rect 1989 -3101 1992 -3095
rect 1996 -3101 1999 -3095
rect 2003 -3101 2006 -3095
rect 2031 -3101 2034 -3095
rect 2045 -3101 2048 -3095
rect 2073 -3101 2076 -3095
rect 1 -3232 7 -3226
rect 8 -3232 14 -3226
rect 15 -3232 21 -3226
rect 92 -3232 95 -3226
rect 99 -3232 102 -3226
rect 106 -3232 109 -3226
rect 113 -3232 119 -3226
rect 120 -3232 123 -3226
rect 127 -3232 130 -3226
rect 134 -3232 137 -3226
rect 141 -3232 144 -3226
rect 148 -3232 151 -3226
rect 155 -3232 158 -3226
rect 162 -3232 165 -3226
rect 169 -3232 175 -3226
rect 176 -3232 179 -3226
rect 183 -3232 189 -3226
rect 190 -3232 196 -3226
rect 197 -3232 200 -3226
rect 204 -3232 210 -3226
rect 211 -3232 214 -3226
rect 218 -3232 221 -3226
rect 225 -3232 228 -3226
rect 232 -3232 235 -3226
rect 239 -3232 242 -3226
rect 246 -3232 249 -3226
rect 253 -3232 256 -3226
rect 260 -3232 263 -3226
rect 267 -3232 270 -3226
rect 274 -3232 277 -3226
rect 281 -3232 284 -3226
rect 288 -3232 291 -3226
rect 295 -3232 298 -3226
rect 302 -3232 305 -3226
rect 309 -3232 312 -3226
rect 316 -3232 319 -3226
rect 323 -3232 326 -3226
rect 330 -3232 333 -3226
rect 337 -3232 340 -3226
rect 344 -3232 347 -3226
rect 351 -3232 354 -3226
rect 358 -3232 361 -3226
rect 365 -3232 368 -3226
rect 372 -3232 375 -3226
rect 379 -3232 382 -3226
rect 386 -3232 389 -3226
rect 393 -3232 396 -3226
rect 400 -3232 406 -3226
rect 407 -3232 410 -3226
rect 414 -3232 420 -3226
rect 421 -3232 427 -3226
rect 428 -3232 431 -3226
rect 435 -3232 438 -3226
rect 442 -3232 445 -3226
rect 449 -3232 452 -3226
rect 456 -3232 459 -3226
rect 463 -3232 466 -3226
rect 470 -3232 473 -3226
rect 477 -3232 480 -3226
rect 484 -3232 487 -3226
rect 491 -3232 497 -3226
rect 498 -3232 501 -3226
rect 505 -3232 508 -3226
rect 512 -3232 515 -3226
rect 519 -3232 522 -3226
rect 526 -3232 529 -3226
rect 533 -3232 536 -3226
rect 540 -3232 543 -3226
rect 547 -3232 550 -3226
rect 554 -3232 557 -3226
rect 561 -3232 564 -3226
rect 568 -3232 571 -3226
rect 575 -3232 581 -3226
rect 582 -3232 585 -3226
rect 589 -3232 592 -3226
rect 596 -3232 599 -3226
rect 603 -3232 606 -3226
rect 610 -3232 616 -3226
rect 617 -3232 620 -3226
rect 624 -3232 627 -3226
rect 631 -3232 634 -3226
rect 638 -3232 641 -3226
rect 645 -3232 648 -3226
rect 652 -3232 655 -3226
rect 659 -3232 662 -3226
rect 666 -3232 669 -3226
rect 673 -3232 679 -3226
rect 680 -3232 683 -3226
rect 687 -3232 690 -3226
rect 694 -3232 697 -3226
rect 701 -3232 704 -3226
rect 708 -3232 711 -3226
rect 715 -3232 721 -3226
rect 722 -3232 725 -3226
rect 729 -3232 732 -3226
rect 736 -3232 739 -3226
rect 743 -3232 749 -3226
rect 750 -3232 753 -3226
rect 757 -3232 760 -3226
rect 764 -3232 770 -3226
rect 771 -3232 774 -3226
rect 778 -3232 781 -3226
rect 785 -3232 788 -3226
rect 792 -3232 795 -3226
rect 799 -3232 805 -3226
rect 806 -3232 809 -3226
rect 813 -3232 819 -3226
rect 820 -3232 823 -3226
rect 827 -3232 830 -3226
rect 834 -3232 837 -3226
rect 841 -3232 844 -3226
rect 848 -3232 851 -3226
rect 855 -3232 858 -3226
rect 862 -3232 865 -3226
rect 869 -3232 875 -3226
rect 876 -3232 879 -3226
rect 883 -3232 886 -3226
rect 890 -3232 893 -3226
rect 897 -3232 900 -3226
rect 904 -3232 907 -3226
rect 911 -3232 914 -3226
rect 918 -3232 921 -3226
rect 925 -3232 928 -3226
rect 932 -3232 935 -3226
rect 939 -3232 945 -3226
rect 946 -3232 949 -3226
rect 953 -3232 959 -3226
rect 960 -3232 963 -3226
rect 967 -3232 970 -3226
rect 974 -3232 977 -3226
rect 981 -3232 987 -3226
rect 988 -3232 991 -3226
rect 995 -3232 998 -3226
rect 1002 -3232 1005 -3226
rect 1009 -3232 1012 -3226
rect 1016 -3232 1019 -3226
rect 1023 -3232 1026 -3226
rect 1030 -3232 1033 -3226
rect 1037 -3232 1040 -3226
rect 1044 -3232 1047 -3226
rect 1051 -3232 1054 -3226
rect 1058 -3232 1061 -3226
rect 1065 -3232 1068 -3226
rect 1072 -3232 1075 -3226
rect 1079 -3232 1082 -3226
rect 1086 -3232 1089 -3226
rect 1093 -3232 1096 -3226
rect 1100 -3232 1103 -3226
rect 1107 -3232 1113 -3226
rect 1114 -3232 1117 -3226
rect 1121 -3232 1124 -3226
rect 1128 -3232 1131 -3226
rect 1135 -3232 1138 -3226
rect 1142 -3232 1145 -3226
rect 1149 -3232 1152 -3226
rect 1156 -3232 1159 -3226
rect 1163 -3232 1169 -3226
rect 1170 -3232 1173 -3226
rect 1177 -3232 1180 -3226
rect 1184 -3232 1187 -3226
rect 1191 -3232 1194 -3226
rect 1198 -3232 1201 -3226
rect 1205 -3232 1208 -3226
rect 1212 -3232 1218 -3226
rect 1219 -3232 1222 -3226
rect 1226 -3232 1229 -3226
rect 1233 -3232 1239 -3226
rect 1240 -3232 1243 -3226
rect 1247 -3232 1250 -3226
rect 1254 -3232 1260 -3226
rect 1261 -3232 1264 -3226
rect 1268 -3232 1271 -3226
rect 1275 -3232 1278 -3226
rect 1282 -3232 1285 -3226
rect 1289 -3232 1292 -3226
rect 1296 -3232 1299 -3226
rect 1303 -3232 1306 -3226
rect 1310 -3232 1313 -3226
rect 1317 -3232 1320 -3226
rect 1324 -3232 1327 -3226
rect 1331 -3232 1334 -3226
rect 1338 -3232 1341 -3226
rect 1345 -3232 1348 -3226
rect 1352 -3232 1358 -3226
rect 1359 -3232 1362 -3226
rect 1366 -3232 1369 -3226
rect 1373 -3232 1376 -3226
rect 1380 -3232 1383 -3226
rect 1387 -3232 1390 -3226
rect 1394 -3232 1397 -3226
rect 1401 -3232 1404 -3226
rect 1408 -3232 1411 -3226
rect 1415 -3232 1418 -3226
rect 1422 -3232 1425 -3226
rect 1429 -3232 1432 -3226
rect 1436 -3232 1439 -3226
rect 1443 -3232 1446 -3226
rect 1450 -3232 1453 -3226
rect 1457 -3232 1463 -3226
rect 1464 -3232 1467 -3226
rect 1471 -3232 1474 -3226
rect 1478 -3232 1481 -3226
rect 1485 -3232 1488 -3226
rect 1492 -3232 1495 -3226
rect 1499 -3232 1502 -3226
rect 1506 -3232 1509 -3226
rect 1513 -3232 1516 -3226
rect 1520 -3232 1523 -3226
rect 1527 -3232 1530 -3226
rect 1534 -3232 1537 -3226
rect 1541 -3232 1544 -3226
rect 1548 -3232 1551 -3226
rect 1555 -3232 1558 -3226
rect 1562 -3232 1565 -3226
rect 1569 -3232 1572 -3226
rect 1576 -3232 1582 -3226
rect 1583 -3232 1586 -3226
rect 1590 -3232 1593 -3226
rect 1597 -3232 1600 -3226
rect 1604 -3232 1607 -3226
rect 1611 -3232 1614 -3226
rect 1618 -3232 1621 -3226
rect 1625 -3232 1628 -3226
rect 1632 -3232 1635 -3226
rect 1639 -3232 1645 -3226
rect 1646 -3232 1652 -3226
rect 1653 -3232 1659 -3226
rect 1660 -3232 1663 -3226
rect 1667 -3232 1673 -3226
rect 1674 -3232 1677 -3226
rect 1681 -3232 1687 -3226
rect 1688 -3232 1691 -3226
rect 1695 -3232 1698 -3226
rect 1702 -3232 1705 -3226
rect 1709 -3232 1712 -3226
rect 1716 -3232 1719 -3226
rect 1723 -3232 1726 -3226
rect 1730 -3232 1733 -3226
rect 1737 -3232 1740 -3226
rect 1744 -3232 1747 -3226
rect 1751 -3232 1754 -3226
rect 1758 -3232 1761 -3226
rect 1765 -3232 1768 -3226
rect 1772 -3232 1775 -3226
rect 1779 -3232 1782 -3226
rect 1807 -3232 1810 -3226
rect 1814 -3232 1817 -3226
rect 1821 -3232 1824 -3226
rect 1849 -3232 1855 -3226
rect 1856 -3232 1859 -3226
rect 1863 -3232 1866 -3226
rect 1877 -3232 1880 -3226
rect 1884 -3232 1887 -3226
rect 1891 -3232 1894 -3226
rect 1905 -3232 1908 -3226
rect 1919 -3232 1922 -3226
rect 1961 -3232 1967 -3226
rect 1968 -3232 1971 -3226
rect 1975 -3232 1978 -3226
rect 1982 -3232 1985 -3226
rect 2017 -3232 2020 -3226
rect 2045 -3232 2048 -3226
rect 1 -3335 7 -3329
rect 8 -3335 14 -3329
rect 15 -3335 21 -3329
rect 22 -3335 28 -3329
rect 29 -3335 35 -3329
rect 36 -3335 42 -3329
rect 141 -3335 144 -3329
rect 162 -3335 165 -3329
rect 169 -3335 172 -3329
rect 176 -3335 179 -3329
rect 183 -3335 186 -3329
rect 190 -3335 193 -3329
rect 197 -3335 200 -3329
rect 204 -3335 207 -3329
rect 211 -3335 217 -3329
rect 218 -3335 221 -3329
rect 225 -3335 231 -3329
rect 232 -3335 238 -3329
rect 239 -3335 242 -3329
rect 246 -3335 249 -3329
rect 253 -3335 259 -3329
rect 260 -3335 263 -3329
rect 267 -3335 270 -3329
rect 274 -3335 277 -3329
rect 281 -3335 284 -3329
rect 288 -3335 291 -3329
rect 295 -3335 298 -3329
rect 302 -3335 305 -3329
rect 309 -3335 312 -3329
rect 316 -3335 319 -3329
rect 323 -3335 326 -3329
rect 330 -3335 333 -3329
rect 337 -3335 340 -3329
rect 344 -3335 347 -3329
rect 351 -3335 354 -3329
rect 358 -3335 361 -3329
rect 365 -3335 368 -3329
rect 372 -3335 375 -3329
rect 379 -3335 385 -3329
rect 386 -3335 389 -3329
rect 393 -3335 396 -3329
rect 400 -3335 403 -3329
rect 407 -3335 410 -3329
rect 414 -3335 420 -3329
rect 421 -3335 424 -3329
rect 428 -3335 431 -3329
rect 435 -3335 438 -3329
rect 442 -3335 445 -3329
rect 449 -3335 452 -3329
rect 456 -3335 459 -3329
rect 463 -3335 466 -3329
rect 470 -3335 473 -3329
rect 477 -3335 480 -3329
rect 484 -3335 487 -3329
rect 491 -3335 494 -3329
rect 498 -3335 501 -3329
rect 505 -3335 508 -3329
rect 512 -3335 515 -3329
rect 519 -3335 522 -3329
rect 526 -3335 529 -3329
rect 533 -3335 539 -3329
rect 540 -3335 543 -3329
rect 547 -3335 550 -3329
rect 554 -3335 557 -3329
rect 561 -3335 564 -3329
rect 568 -3335 571 -3329
rect 575 -3335 578 -3329
rect 582 -3335 585 -3329
rect 589 -3335 592 -3329
rect 596 -3335 602 -3329
rect 603 -3335 606 -3329
rect 610 -3335 613 -3329
rect 617 -3335 620 -3329
rect 624 -3335 627 -3329
rect 631 -3335 634 -3329
rect 638 -3335 644 -3329
rect 645 -3335 648 -3329
rect 652 -3335 655 -3329
rect 659 -3335 662 -3329
rect 666 -3335 669 -3329
rect 673 -3335 676 -3329
rect 680 -3335 683 -3329
rect 687 -3335 690 -3329
rect 694 -3335 697 -3329
rect 701 -3335 704 -3329
rect 708 -3335 711 -3329
rect 715 -3335 718 -3329
rect 722 -3335 728 -3329
rect 729 -3335 735 -3329
rect 736 -3335 739 -3329
rect 743 -3335 746 -3329
rect 750 -3335 753 -3329
rect 757 -3335 760 -3329
rect 764 -3335 767 -3329
rect 771 -3335 774 -3329
rect 778 -3335 784 -3329
rect 785 -3335 788 -3329
rect 792 -3335 795 -3329
rect 799 -3335 802 -3329
rect 806 -3335 809 -3329
rect 813 -3335 816 -3329
rect 820 -3335 823 -3329
rect 827 -3335 830 -3329
rect 834 -3335 837 -3329
rect 841 -3335 844 -3329
rect 848 -3335 854 -3329
rect 855 -3335 858 -3329
rect 862 -3335 865 -3329
rect 869 -3335 872 -3329
rect 876 -3335 879 -3329
rect 883 -3335 886 -3329
rect 890 -3335 893 -3329
rect 897 -3335 900 -3329
rect 904 -3335 907 -3329
rect 911 -3335 914 -3329
rect 918 -3335 921 -3329
rect 925 -3335 931 -3329
rect 932 -3335 935 -3329
rect 939 -3335 942 -3329
rect 946 -3335 949 -3329
rect 953 -3335 959 -3329
rect 960 -3335 963 -3329
rect 967 -3335 973 -3329
rect 974 -3335 980 -3329
rect 981 -3335 984 -3329
rect 988 -3335 994 -3329
rect 995 -3335 998 -3329
rect 1002 -3335 1005 -3329
rect 1009 -3335 1012 -3329
rect 1016 -3335 1019 -3329
rect 1023 -3335 1026 -3329
rect 1030 -3335 1033 -3329
rect 1037 -3335 1040 -3329
rect 1044 -3335 1047 -3329
rect 1051 -3335 1054 -3329
rect 1058 -3335 1061 -3329
rect 1065 -3335 1071 -3329
rect 1072 -3335 1075 -3329
rect 1079 -3335 1085 -3329
rect 1086 -3335 1089 -3329
rect 1093 -3335 1099 -3329
rect 1100 -3335 1106 -3329
rect 1107 -3335 1110 -3329
rect 1114 -3335 1117 -3329
rect 1121 -3335 1124 -3329
rect 1128 -3335 1131 -3329
rect 1135 -3335 1138 -3329
rect 1142 -3335 1145 -3329
rect 1149 -3335 1152 -3329
rect 1156 -3335 1159 -3329
rect 1163 -3335 1166 -3329
rect 1170 -3335 1173 -3329
rect 1177 -3335 1180 -3329
rect 1184 -3335 1187 -3329
rect 1191 -3335 1194 -3329
rect 1198 -3335 1201 -3329
rect 1205 -3335 1208 -3329
rect 1212 -3335 1218 -3329
rect 1219 -3335 1222 -3329
rect 1226 -3335 1229 -3329
rect 1233 -3335 1239 -3329
rect 1240 -3335 1243 -3329
rect 1247 -3335 1250 -3329
rect 1254 -3335 1257 -3329
rect 1261 -3335 1264 -3329
rect 1268 -3335 1274 -3329
rect 1275 -3335 1278 -3329
rect 1282 -3335 1285 -3329
rect 1289 -3335 1292 -3329
rect 1296 -3335 1299 -3329
rect 1303 -3335 1306 -3329
rect 1310 -3335 1313 -3329
rect 1317 -3335 1320 -3329
rect 1324 -3335 1327 -3329
rect 1331 -3335 1334 -3329
rect 1338 -3335 1344 -3329
rect 1345 -3335 1348 -3329
rect 1352 -3335 1355 -3329
rect 1359 -3335 1362 -3329
rect 1366 -3335 1372 -3329
rect 1373 -3335 1376 -3329
rect 1380 -3335 1386 -3329
rect 1387 -3335 1390 -3329
rect 1394 -3335 1397 -3329
rect 1401 -3335 1404 -3329
rect 1408 -3335 1411 -3329
rect 1415 -3335 1421 -3329
rect 1422 -3335 1425 -3329
rect 1429 -3335 1432 -3329
rect 1436 -3335 1439 -3329
rect 1443 -3335 1446 -3329
rect 1450 -3335 1453 -3329
rect 1457 -3335 1460 -3329
rect 1464 -3335 1467 -3329
rect 1471 -3335 1474 -3329
rect 1478 -3335 1481 -3329
rect 1485 -3335 1488 -3329
rect 1492 -3335 1495 -3329
rect 1499 -3335 1502 -3329
rect 1506 -3335 1509 -3329
rect 1513 -3335 1516 -3329
rect 1520 -3335 1523 -3329
rect 1527 -3335 1530 -3329
rect 1555 -3335 1558 -3329
rect 1562 -3335 1565 -3329
rect 1590 -3335 1593 -3329
rect 1597 -3335 1600 -3329
rect 1604 -3335 1610 -3329
rect 1625 -3335 1628 -3329
rect 1653 -3335 1656 -3329
rect 1660 -3335 1663 -3329
rect 1667 -3335 1670 -3329
rect 1716 -3335 1719 -3329
rect 1723 -3335 1729 -3329
rect 1730 -3335 1733 -3329
rect 1737 -3335 1740 -3329
rect 1744 -3335 1747 -3329
rect 1751 -3335 1754 -3329
rect 1765 -3335 1768 -3329
rect 1779 -3335 1782 -3329
rect 1786 -3335 1789 -3329
rect 1793 -3335 1796 -3329
rect 1800 -3335 1803 -3329
rect 1814 -3335 1817 -3329
rect 1835 -3335 1838 -3329
rect 1842 -3335 1845 -3329
rect 1849 -3335 1855 -3329
rect 1856 -3335 1859 -3329
rect 1863 -3335 1866 -3329
rect 1870 -3335 1873 -3329
rect 1877 -3335 1880 -3329
rect 1884 -3335 1890 -3329
rect 1891 -3335 1894 -3329
rect 1905 -3335 1908 -3329
rect 1961 -3335 1964 -3329
rect 1968 -3335 1971 -3329
rect 2024 -3335 2027 -3329
rect 2031 -3335 2034 -3329
rect 1 -3422 7 -3416
rect 8 -3422 14 -3416
rect 15 -3422 21 -3416
rect 22 -3422 28 -3416
rect 29 -3422 35 -3416
rect 36 -3422 42 -3416
rect 43 -3422 49 -3416
rect 50 -3422 56 -3416
rect 169 -3422 175 -3416
rect 176 -3422 182 -3416
rect 295 -3422 298 -3416
rect 309 -3422 312 -3416
rect 316 -3422 322 -3416
rect 330 -3422 333 -3416
rect 337 -3422 340 -3416
rect 344 -3422 347 -3416
rect 358 -3422 361 -3416
rect 372 -3422 375 -3416
rect 379 -3422 382 -3416
rect 386 -3422 392 -3416
rect 393 -3422 396 -3416
rect 400 -3422 406 -3416
rect 407 -3422 410 -3416
rect 421 -3422 424 -3416
rect 428 -3422 431 -3416
rect 435 -3422 441 -3416
rect 442 -3422 445 -3416
rect 449 -3422 452 -3416
rect 456 -3422 459 -3416
rect 463 -3422 466 -3416
rect 470 -3422 476 -3416
rect 477 -3422 480 -3416
rect 484 -3422 490 -3416
rect 491 -3422 494 -3416
rect 498 -3422 501 -3416
rect 505 -3422 508 -3416
rect 512 -3422 515 -3416
rect 519 -3422 522 -3416
rect 526 -3422 529 -3416
rect 533 -3422 536 -3416
rect 540 -3422 543 -3416
rect 547 -3422 550 -3416
rect 554 -3422 560 -3416
rect 561 -3422 564 -3416
rect 568 -3422 571 -3416
rect 575 -3422 578 -3416
rect 582 -3422 585 -3416
rect 589 -3422 592 -3416
rect 596 -3422 599 -3416
rect 603 -3422 606 -3416
rect 610 -3422 613 -3416
rect 617 -3422 620 -3416
rect 624 -3422 627 -3416
rect 631 -3422 634 -3416
rect 638 -3422 641 -3416
rect 645 -3422 648 -3416
rect 652 -3422 655 -3416
rect 659 -3422 662 -3416
rect 666 -3422 672 -3416
rect 673 -3422 676 -3416
rect 680 -3422 683 -3416
rect 687 -3422 690 -3416
rect 694 -3422 697 -3416
rect 701 -3422 704 -3416
rect 708 -3422 711 -3416
rect 715 -3422 718 -3416
rect 722 -3422 728 -3416
rect 729 -3422 732 -3416
rect 736 -3422 739 -3416
rect 743 -3422 746 -3416
rect 750 -3422 753 -3416
rect 757 -3422 760 -3416
rect 764 -3422 767 -3416
rect 771 -3422 774 -3416
rect 778 -3422 781 -3416
rect 785 -3422 788 -3416
rect 792 -3422 795 -3416
rect 799 -3422 805 -3416
rect 806 -3422 809 -3416
rect 813 -3422 816 -3416
rect 820 -3422 823 -3416
rect 827 -3422 830 -3416
rect 834 -3422 837 -3416
rect 841 -3422 847 -3416
rect 848 -3422 851 -3416
rect 855 -3422 861 -3416
rect 862 -3422 865 -3416
rect 869 -3422 872 -3416
rect 876 -3422 879 -3416
rect 883 -3422 886 -3416
rect 890 -3422 893 -3416
rect 897 -3422 903 -3416
rect 904 -3422 907 -3416
rect 911 -3422 914 -3416
rect 918 -3422 924 -3416
rect 925 -3422 928 -3416
rect 932 -3422 938 -3416
rect 939 -3422 942 -3416
rect 946 -3422 949 -3416
rect 953 -3422 956 -3416
rect 960 -3422 963 -3416
rect 967 -3422 970 -3416
rect 974 -3422 977 -3416
rect 981 -3422 984 -3416
rect 988 -3422 994 -3416
rect 995 -3422 998 -3416
rect 1002 -3422 1005 -3416
rect 1009 -3422 1012 -3416
rect 1016 -3422 1019 -3416
rect 1023 -3422 1029 -3416
rect 1030 -3422 1036 -3416
rect 1037 -3422 1040 -3416
rect 1044 -3422 1047 -3416
rect 1051 -3422 1054 -3416
rect 1058 -3422 1061 -3416
rect 1065 -3422 1071 -3416
rect 1072 -3422 1075 -3416
rect 1079 -3422 1082 -3416
rect 1086 -3422 1089 -3416
rect 1093 -3422 1096 -3416
rect 1100 -3422 1103 -3416
rect 1107 -3422 1110 -3416
rect 1114 -3422 1117 -3416
rect 1121 -3422 1127 -3416
rect 1135 -3422 1138 -3416
rect 1142 -3422 1145 -3416
rect 1156 -3422 1162 -3416
rect 1170 -3422 1173 -3416
rect 1177 -3422 1180 -3416
rect 1184 -3422 1187 -3416
rect 1191 -3422 1194 -3416
rect 1198 -3422 1201 -3416
rect 1205 -3422 1211 -3416
rect 1212 -3422 1215 -3416
rect 1219 -3422 1222 -3416
rect 1226 -3422 1229 -3416
rect 1233 -3422 1236 -3416
rect 1240 -3422 1243 -3416
rect 1247 -3422 1250 -3416
rect 1254 -3422 1257 -3416
rect 1261 -3422 1264 -3416
rect 1268 -3422 1271 -3416
rect 1275 -3422 1281 -3416
rect 1282 -3422 1285 -3416
rect 1289 -3422 1292 -3416
rect 1296 -3422 1299 -3416
rect 1303 -3422 1309 -3416
rect 1331 -3422 1334 -3416
rect 1345 -3422 1348 -3416
rect 1359 -3422 1362 -3416
rect 1366 -3422 1369 -3416
rect 1373 -3422 1379 -3416
rect 1380 -3422 1383 -3416
rect 1450 -3422 1453 -3416
rect 1457 -3422 1460 -3416
rect 1464 -3422 1467 -3416
rect 1471 -3422 1474 -3416
rect 1499 -3422 1502 -3416
rect 1520 -3422 1523 -3416
rect 1527 -3422 1530 -3416
rect 1548 -3422 1554 -3416
rect 1583 -3422 1589 -3416
rect 1611 -3422 1614 -3416
rect 1646 -3422 1649 -3416
rect 1653 -3422 1656 -3416
rect 1723 -3422 1726 -3416
rect 1730 -3422 1733 -3416
rect 1737 -3422 1740 -3416
rect 1758 -3422 1761 -3416
rect 1765 -3422 1771 -3416
rect 1779 -3422 1782 -3416
rect 1786 -3422 1789 -3416
rect 1800 -3422 1803 -3416
rect 1807 -3422 1813 -3416
rect 1821 -3422 1824 -3416
rect 1828 -3422 1831 -3416
rect 1835 -3422 1838 -3416
rect 1842 -3422 1845 -3416
rect 1849 -3422 1852 -3416
rect 1856 -3422 1859 -3416
rect 1863 -3422 1866 -3416
rect 1870 -3422 1873 -3416
rect 1954 -3422 1957 -3416
rect 1961 -3422 1964 -3416
rect 2024 -3422 2027 -3416
rect 2031 -3422 2034 -3416
rect 1 -3467 7 -3461
rect 8 -3467 14 -3461
rect 15 -3467 21 -3461
rect 22 -3467 28 -3461
rect 29 -3467 35 -3461
rect 36 -3467 42 -3461
rect 43 -3467 49 -3461
rect 50 -3467 56 -3461
rect 57 -3467 63 -3461
rect 64 -3467 70 -3461
rect 71 -3467 77 -3461
rect 169 -3467 175 -3461
rect 267 -3467 273 -3461
rect 323 -3467 326 -3461
rect 379 -3467 382 -3461
rect 414 -3467 417 -3461
rect 421 -3467 424 -3461
rect 435 -3467 441 -3461
rect 442 -3467 445 -3461
rect 456 -3467 459 -3461
rect 463 -3467 469 -3461
rect 484 -3467 487 -3461
rect 491 -3467 494 -3461
rect 498 -3467 501 -3461
rect 505 -3467 508 -3461
rect 512 -3467 515 -3461
rect 519 -3467 525 -3461
rect 533 -3467 536 -3461
rect 540 -3467 543 -3461
rect 547 -3467 553 -3461
rect 554 -3467 557 -3461
rect 561 -3467 564 -3461
rect 568 -3467 571 -3461
rect 575 -3467 581 -3461
rect 582 -3467 585 -3461
rect 589 -3467 595 -3461
rect 596 -3467 599 -3461
rect 603 -3467 606 -3461
rect 610 -3467 613 -3461
rect 617 -3467 623 -3461
rect 624 -3467 630 -3461
rect 631 -3467 634 -3461
rect 638 -3467 644 -3461
rect 645 -3467 648 -3461
rect 652 -3467 655 -3461
rect 659 -3467 662 -3461
rect 666 -3467 669 -3461
rect 673 -3467 676 -3461
rect 680 -3467 686 -3461
rect 687 -3467 690 -3461
rect 694 -3467 697 -3461
rect 701 -3467 707 -3461
rect 708 -3467 711 -3461
rect 715 -3467 718 -3461
rect 722 -3467 725 -3461
rect 729 -3467 735 -3461
rect 736 -3467 739 -3461
rect 743 -3467 746 -3461
rect 750 -3467 753 -3461
rect 757 -3467 760 -3461
rect 778 -3467 781 -3461
rect 792 -3467 795 -3461
rect 799 -3467 802 -3461
rect 806 -3467 809 -3461
rect 813 -3467 816 -3461
rect 820 -3467 823 -3461
rect 827 -3467 830 -3461
rect 834 -3467 837 -3461
rect 841 -3467 844 -3461
rect 848 -3467 851 -3461
rect 876 -3467 879 -3461
rect 883 -3467 886 -3461
rect 911 -3467 917 -3461
rect 918 -3467 924 -3461
rect 953 -3467 956 -3461
rect 974 -3467 977 -3461
rect 995 -3467 998 -3461
rect 1002 -3467 1005 -3461
rect 1009 -3467 1012 -3461
rect 1016 -3467 1019 -3461
rect 1023 -3467 1026 -3461
rect 1030 -3467 1033 -3461
rect 1037 -3467 1040 -3461
rect 1044 -3467 1047 -3461
rect 1051 -3467 1054 -3461
rect 1058 -3467 1064 -3461
rect 1065 -3467 1068 -3461
rect 1072 -3467 1075 -3461
rect 1079 -3467 1085 -3461
rect 1086 -3467 1089 -3461
rect 1093 -3467 1096 -3461
rect 1100 -3467 1103 -3461
rect 1107 -3467 1110 -3461
rect 1121 -3467 1127 -3461
rect 1128 -3467 1131 -3461
rect 1156 -3467 1159 -3461
rect 1163 -3467 1166 -3461
rect 1170 -3467 1173 -3461
rect 1177 -3467 1183 -3461
rect 1184 -3467 1187 -3461
rect 1191 -3467 1194 -3461
rect 1198 -3467 1201 -3461
rect 1205 -3467 1208 -3461
rect 1212 -3467 1215 -3461
rect 1219 -3467 1222 -3461
rect 1226 -3467 1229 -3461
rect 1233 -3467 1236 -3461
rect 1240 -3467 1243 -3461
rect 1247 -3467 1250 -3461
rect 1282 -3467 1288 -3461
rect 1289 -3467 1292 -3461
rect 1303 -3467 1309 -3461
rect 1310 -3467 1313 -3461
rect 1317 -3467 1323 -3461
rect 1324 -3467 1327 -3461
rect 1331 -3467 1334 -3461
rect 1359 -3467 1362 -3461
rect 1436 -3467 1439 -3461
rect 1443 -3467 1446 -3461
rect 1450 -3467 1453 -3461
rect 1457 -3467 1463 -3461
rect 1464 -3467 1467 -3461
rect 1492 -3467 1495 -3461
rect 1499 -3467 1502 -3461
rect 1513 -3467 1516 -3461
rect 1520 -3467 1523 -3461
rect 1625 -3467 1631 -3461
rect 1639 -3467 1642 -3461
rect 1723 -3467 1726 -3461
rect 1730 -3467 1733 -3461
rect 1744 -3467 1750 -3461
rect 1765 -3467 1768 -3461
rect 1779 -3467 1782 -3461
rect 1793 -3467 1796 -3461
rect 1821 -3467 1824 -3461
rect 1828 -3467 1831 -3461
rect 1835 -3467 1841 -3461
rect 1842 -3467 1845 -3461
rect 1849 -3467 1852 -3461
rect 1856 -3467 1862 -3461
rect 1863 -3467 1866 -3461
rect 1870 -3467 1873 -3461
rect 1954 -3467 1957 -3461
rect 1961 -3467 1964 -3461
rect 2024 -3467 2027 -3461
rect 2031 -3467 2034 -3461
rect 1 -3496 7 -3490
rect 8 -3496 14 -3490
rect 15 -3496 21 -3490
rect 22 -3496 28 -3490
rect 29 -3496 35 -3490
rect 36 -3496 42 -3490
rect 43 -3496 49 -3490
rect 50 -3496 56 -3490
rect 57 -3496 63 -3490
rect 64 -3496 70 -3490
rect 71 -3496 77 -3490
rect 78 -3496 84 -3490
rect 85 -3496 91 -3490
rect 92 -3496 98 -3490
rect 99 -3496 105 -3490
rect 106 -3496 112 -3490
rect 113 -3496 119 -3490
rect 120 -3496 126 -3490
rect 127 -3496 133 -3490
rect 134 -3496 140 -3490
rect 141 -3496 147 -3490
rect 148 -3496 154 -3490
rect 330 -3496 333 -3490
rect 365 -3496 371 -3490
rect 386 -3496 389 -3490
rect 393 -3496 396 -3490
rect 428 -3496 434 -3490
rect 463 -3496 466 -3490
rect 470 -3496 473 -3490
rect 477 -3496 480 -3490
rect 484 -3496 487 -3490
rect 519 -3496 525 -3490
rect 533 -3496 536 -3490
rect 540 -3496 543 -3490
rect 568 -3496 571 -3490
rect 582 -3496 585 -3490
rect 589 -3496 592 -3490
rect 603 -3496 606 -3490
rect 610 -3496 613 -3490
rect 617 -3496 620 -3490
rect 631 -3496 634 -3490
rect 638 -3496 641 -3490
rect 645 -3496 648 -3490
rect 652 -3496 658 -3490
rect 680 -3496 683 -3490
rect 715 -3496 718 -3490
rect 736 -3496 739 -3490
rect 743 -3496 746 -3490
rect 750 -3496 753 -3490
rect 757 -3496 760 -3490
rect 764 -3496 767 -3490
rect 771 -3496 774 -3490
rect 778 -3496 781 -3490
rect 785 -3496 791 -3490
rect 792 -3496 795 -3490
rect 813 -3496 816 -3490
rect 827 -3496 830 -3490
rect 841 -3496 844 -3490
rect 862 -3496 868 -3490
rect 869 -3496 872 -3490
rect 883 -3496 889 -3490
rect 897 -3496 900 -3490
rect 974 -3496 977 -3490
rect 995 -3496 998 -3490
rect 1009 -3496 1012 -3490
rect 1016 -3496 1019 -3490
rect 1023 -3496 1026 -3490
rect 1030 -3496 1033 -3490
rect 1037 -3496 1040 -3490
rect 1044 -3496 1047 -3490
rect 1051 -3496 1054 -3490
rect 1058 -3496 1061 -3490
rect 1065 -3496 1068 -3490
rect 1079 -3496 1082 -3490
rect 1142 -3496 1145 -3490
rect 1177 -3496 1180 -3490
rect 1191 -3496 1194 -3490
rect 1233 -3496 1236 -3490
rect 1240 -3496 1243 -3490
rect 1247 -3496 1253 -3490
rect 1254 -3496 1257 -3490
rect 1261 -3496 1267 -3490
rect 1268 -3496 1274 -3490
rect 1275 -3496 1278 -3490
rect 1282 -3496 1288 -3490
rect 1289 -3496 1292 -3490
rect 1303 -3496 1306 -3490
rect 1310 -3496 1316 -3490
rect 1359 -3496 1362 -3490
rect 1429 -3496 1435 -3490
rect 1436 -3496 1439 -3490
rect 1492 -3496 1495 -3490
rect 1499 -3496 1505 -3490
rect 1506 -3496 1509 -3490
rect 1513 -3496 1516 -3490
rect 1520 -3496 1523 -3490
rect 1569 -3496 1572 -3490
rect 1639 -3496 1642 -3490
rect 1723 -3496 1729 -3490
rect 1730 -3496 1733 -3490
rect 1779 -3496 1782 -3490
rect 1786 -3496 1792 -3490
rect 1842 -3496 1845 -3490
rect 1849 -3496 1852 -3490
rect 1863 -3496 1866 -3490
rect 1954 -3496 1960 -3490
rect 2024 -3496 2027 -3490
rect 2031 -3496 2034 -3490
rect 1 -3519 7 -3513
rect 8 -3519 14 -3513
rect 15 -3519 21 -3513
rect 22 -3519 28 -3513
rect 29 -3519 35 -3513
rect 36 -3519 42 -3513
rect 43 -3519 49 -3513
rect 50 -3519 56 -3513
rect 57 -3519 63 -3513
rect 64 -3519 70 -3513
rect 71 -3519 77 -3513
rect 78 -3519 84 -3513
rect 85 -3519 91 -3513
rect 92 -3519 98 -3513
rect 99 -3519 105 -3513
rect 106 -3519 112 -3513
rect 113 -3519 119 -3513
rect 120 -3519 126 -3513
rect 127 -3519 133 -3513
rect 134 -3519 140 -3513
rect 141 -3519 147 -3513
rect 148 -3519 154 -3513
rect 155 -3519 161 -3513
rect 162 -3519 168 -3513
rect 169 -3519 175 -3513
rect 176 -3519 182 -3513
rect 183 -3519 189 -3513
rect 190 -3519 196 -3513
rect 197 -3519 203 -3513
rect 204 -3519 210 -3513
rect 211 -3519 217 -3513
rect 337 -3519 343 -3513
rect 393 -3519 396 -3513
rect 428 -3519 431 -3513
rect 463 -3519 466 -3513
rect 477 -3519 480 -3513
rect 540 -3519 543 -3513
rect 547 -3519 550 -3513
rect 575 -3519 578 -3513
rect 582 -3519 585 -3513
rect 603 -3519 606 -3513
rect 610 -3519 613 -3513
rect 617 -3519 620 -3513
rect 624 -3519 627 -3513
rect 631 -3519 634 -3513
rect 638 -3519 641 -3513
rect 708 -3519 711 -3513
rect 729 -3519 732 -3513
rect 736 -3519 739 -3513
rect 743 -3519 746 -3513
rect 750 -3519 753 -3513
rect 757 -3519 760 -3513
rect 764 -3519 767 -3513
rect 771 -3519 777 -3513
rect 778 -3519 781 -3513
rect 785 -3519 791 -3513
rect 792 -3519 795 -3513
rect 799 -3519 802 -3513
rect 806 -3519 812 -3513
rect 890 -3519 893 -3513
rect 967 -3519 970 -3513
rect 1002 -3519 1005 -3513
rect 1009 -3519 1012 -3513
rect 1016 -3519 1019 -3513
rect 1023 -3519 1026 -3513
rect 1030 -3519 1033 -3513
rect 1037 -3519 1040 -3513
rect 1044 -3519 1047 -3513
rect 1051 -3519 1054 -3513
rect 1058 -3519 1064 -3513
rect 1065 -3519 1068 -3513
rect 1121 -3519 1124 -3513
rect 1149 -3519 1152 -3513
rect 1156 -3519 1162 -3513
rect 1205 -3519 1208 -3513
rect 1233 -3519 1236 -3513
rect 1359 -3519 1362 -3513
rect 1366 -3519 1372 -3513
rect 1506 -3519 1509 -3513
rect 1513 -3519 1516 -3513
rect 1520 -3519 1523 -3513
rect 1611 -3519 1614 -3513
rect 1639 -3519 1642 -3513
rect 1849 -3519 1852 -3513
rect 1856 -3519 1862 -3513
rect 2024 -3519 2027 -3513
rect 2031 -3519 2034 -3513
rect 1 -3538 7 -3532
rect 8 -3538 14 -3532
rect 15 -3538 21 -3532
rect 22 -3538 28 -3532
rect 29 -3538 35 -3532
rect 36 -3538 42 -3532
rect 43 -3538 49 -3532
rect 50 -3538 56 -3532
rect 57 -3538 63 -3532
rect 64 -3538 70 -3532
rect 71 -3538 77 -3532
rect 78 -3538 84 -3532
rect 85 -3538 91 -3532
rect 92 -3538 98 -3532
rect 99 -3538 105 -3532
rect 106 -3538 112 -3532
rect 113 -3538 119 -3532
rect 120 -3538 126 -3532
rect 127 -3538 133 -3532
rect 134 -3538 140 -3532
rect 141 -3538 147 -3532
rect 148 -3538 154 -3532
rect 155 -3538 161 -3532
rect 162 -3538 168 -3532
rect 169 -3538 175 -3532
rect 176 -3538 182 -3532
rect 183 -3538 189 -3532
rect 190 -3538 196 -3532
rect 197 -3538 203 -3532
rect 204 -3538 210 -3532
rect 211 -3538 217 -3532
rect 393 -3538 396 -3532
rect 407 -3538 410 -3532
rect 463 -3538 466 -3532
rect 470 -3538 476 -3532
rect 477 -3538 480 -3532
rect 540 -3538 543 -3532
rect 547 -3538 550 -3532
rect 575 -3538 578 -3532
rect 582 -3538 585 -3532
rect 603 -3538 606 -3532
rect 610 -3538 613 -3532
rect 617 -3538 620 -3532
rect 624 -3538 630 -3532
rect 631 -3538 637 -3532
rect 638 -3538 641 -3532
rect 645 -3538 648 -3532
rect 708 -3538 711 -3532
rect 715 -3538 718 -3532
rect 722 -3538 725 -3532
rect 729 -3538 732 -3532
rect 736 -3538 742 -3532
rect 743 -3538 746 -3532
rect 764 -3538 767 -3532
rect 785 -3538 788 -3532
rect 792 -3538 795 -3532
rect 925 -3538 928 -3532
rect 967 -3538 973 -3532
rect 1009 -3538 1012 -3532
rect 1023 -3538 1029 -3532
rect 1030 -3538 1033 -3532
rect 1037 -3538 1043 -3532
rect 1044 -3538 1047 -3532
rect 1058 -3538 1061 -3532
rect 1065 -3538 1068 -3532
rect 1212 -3538 1215 -3532
rect 1219 -3538 1225 -3532
rect 1506 -3538 1509 -3532
rect 1513 -3538 1516 -3532
rect 1520 -3538 1523 -3532
rect 1632 -3538 1635 -3532
rect 1639 -3538 1642 -3532
rect 2024 -3538 2027 -3532
rect 2031 -3538 2034 -3532
rect 1 -3553 7 -3547
rect 8 -3553 14 -3547
rect 15 -3553 21 -3547
rect 22 -3553 28 -3547
rect 29 -3553 35 -3547
rect 36 -3553 42 -3547
rect 43 -3553 49 -3547
rect 50 -3553 56 -3547
rect 57 -3553 63 -3547
rect 64 -3553 70 -3547
rect 71 -3553 77 -3547
rect 78 -3553 84 -3547
rect 85 -3553 91 -3547
rect 92 -3553 98 -3547
rect 99 -3553 105 -3547
rect 106 -3553 112 -3547
rect 113 -3553 119 -3547
rect 120 -3553 126 -3547
rect 127 -3553 133 -3547
rect 134 -3553 140 -3547
rect 141 -3553 147 -3547
rect 148 -3553 154 -3547
rect 155 -3553 161 -3547
rect 162 -3553 168 -3547
rect 169 -3553 175 -3547
rect 176 -3553 182 -3547
rect 183 -3553 189 -3547
rect 190 -3553 196 -3547
rect 197 -3553 203 -3547
rect 204 -3553 210 -3547
rect 211 -3553 217 -3547
rect 218 -3553 224 -3547
rect 225 -3553 231 -3547
rect 232 -3553 238 -3547
rect 239 -3553 245 -3547
rect 400 -3553 403 -3547
rect 407 -3553 410 -3547
rect 540 -3553 543 -3547
rect 547 -3553 553 -3547
rect 554 -3553 557 -3547
rect 582 -3553 588 -3547
rect 589 -3553 592 -3547
rect 603 -3553 606 -3547
rect 610 -3553 613 -3547
rect 617 -3553 620 -3547
rect 645 -3553 648 -3547
rect 701 -3553 704 -3547
rect 715 -3553 718 -3547
rect 722 -3553 725 -3547
rect 729 -3553 732 -3547
rect 757 -3553 760 -3547
rect 785 -3553 791 -3547
rect 792 -3553 795 -3547
rect 1016 -3553 1022 -3547
rect 1037 -3553 1040 -3547
rect 1058 -3553 1061 -3547
rect 1506 -3553 1509 -3547
rect 1513 -3553 1516 -3547
rect 1520 -3553 1523 -3547
rect 1639 -3553 1642 -3547
rect 1646 -3553 1649 -3547
rect 2024 -3553 2027 -3547
rect 2031 -3553 2034 -3547
rect 1 -3568 7 -3562
rect 8 -3568 14 -3562
rect 15 -3568 21 -3562
rect 22 -3568 28 -3562
rect 29 -3568 35 -3562
rect 36 -3568 42 -3562
rect 43 -3568 49 -3562
rect 50 -3568 56 -3562
rect 57 -3568 63 -3562
rect 64 -3568 70 -3562
rect 71 -3568 77 -3562
rect 78 -3568 84 -3562
rect 85 -3568 91 -3562
rect 92 -3568 98 -3562
rect 99 -3568 105 -3562
rect 106 -3568 112 -3562
rect 113 -3568 119 -3562
rect 120 -3568 126 -3562
rect 127 -3568 133 -3562
rect 134 -3568 140 -3562
rect 141 -3568 147 -3562
rect 148 -3568 154 -3562
rect 155 -3568 161 -3562
rect 162 -3568 168 -3562
rect 169 -3568 175 -3562
rect 176 -3568 182 -3562
rect 183 -3568 189 -3562
rect 190 -3568 196 -3562
rect 197 -3568 203 -3562
rect 204 -3568 210 -3562
rect 211 -3568 217 -3562
rect 218 -3568 224 -3562
rect 225 -3568 231 -3562
rect 232 -3568 238 -3562
rect 239 -3568 245 -3562
rect 400 -3568 403 -3562
rect 407 -3568 410 -3562
rect 603 -3568 606 -3562
rect 610 -3568 613 -3562
rect 617 -3568 620 -3562
rect 645 -3568 651 -3562
rect 701 -3568 704 -3562
rect 715 -3568 718 -3562
rect 722 -3568 725 -3562
rect 729 -3568 732 -3562
rect 757 -3568 760 -3562
rect 1058 -3568 1064 -3562
rect 1065 -3568 1068 -3562
rect 1513 -3568 1519 -3562
rect 1520 -3568 1523 -3562
rect 1639 -3568 1642 -3562
rect 1646 -3568 1649 -3562
rect 2024 -3568 2030 -3562
rect 1 -3583 7 -3577
rect 8 -3583 14 -3577
rect 15 -3583 21 -3577
rect 22 -3583 28 -3577
rect 29 -3583 35 -3577
rect 36 -3583 42 -3577
rect 43 -3583 49 -3577
rect 50 -3583 56 -3577
rect 57 -3583 63 -3577
rect 64 -3583 70 -3577
rect 71 -3583 77 -3577
rect 78 -3583 84 -3577
rect 85 -3583 91 -3577
rect 92 -3583 98 -3577
rect 99 -3583 105 -3577
rect 106 -3583 112 -3577
rect 113 -3583 119 -3577
rect 120 -3583 126 -3577
rect 127 -3583 133 -3577
rect 134 -3583 140 -3577
rect 141 -3583 147 -3577
rect 148 -3583 154 -3577
rect 155 -3583 161 -3577
rect 162 -3583 168 -3577
rect 169 -3583 175 -3577
rect 176 -3583 182 -3577
rect 183 -3583 189 -3577
rect 190 -3583 196 -3577
rect 197 -3583 203 -3577
rect 204 -3583 210 -3577
rect 211 -3583 217 -3577
rect 218 -3583 224 -3577
rect 225 -3583 231 -3577
rect 232 -3583 238 -3577
rect 239 -3583 245 -3577
rect 246 -3583 252 -3577
rect 253 -3583 259 -3577
rect 260 -3583 266 -3577
rect 267 -3583 273 -3577
rect 400 -3583 403 -3577
rect 407 -3583 410 -3577
rect 603 -3583 606 -3577
rect 610 -3583 613 -3577
rect 617 -3583 620 -3577
rect 701 -3583 704 -3577
rect 715 -3583 718 -3577
rect 722 -3583 725 -3577
rect 729 -3583 732 -3577
rect 757 -3583 760 -3577
rect 1639 -3583 1642 -3577
rect 1646 -3583 1649 -3577
rect 1 -3596 7 -3590
rect 8 -3596 14 -3590
rect 15 -3596 21 -3590
rect 22 -3596 28 -3590
rect 29 -3596 35 -3590
rect 36 -3596 42 -3590
rect 43 -3596 49 -3590
rect 50 -3596 56 -3590
rect 57 -3596 63 -3590
rect 64 -3596 70 -3590
rect 71 -3596 77 -3590
rect 78 -3596 84 -3590
rect 85 -3596 91 -3590
rect 92 -3596 98 -3590
rect 99 -3596 105 -3590
rect 106 -3596 112 -3590
rect 113 -3596 119 -3590
rect 120 -3596 126 -3590
rect 127 -3596 133 -3590
rect 134 -3596 140 -3590
rect 141 -3596 147 -3590
rect 148 -3596 154 -3590
rect 155 -3596 161 -3590
rect 162 -3596 168 -3590
rect 169 -3596 175 -3590
rect 176 -3596 182 -3590
rect 183 -3596 189 -3590
rect 190 -3596 196 -3590
rect 197 -3596 203 -3590
rect 204 -3596 210 -3590
rect 211 -3596 217 -3590
rect 218 -3596 224 -3590
rect 225 -3596 231 -3590
rect 232 -3596 238 -3590
rect 239 -3596 245 -3590
rect 246 -3596 252 -3590
rect 393 -3596 396 -3590
rect 400 -3596 403 -3590
rect 603 -3596 606 -3590
rect 610 -3596 613 -3590
rect 617 -3596 623 -3590
rect 701 -3596 704 -3590
rect 722 -3596 728 -3590
rect 729 -3596 732 -3590
rect 757 -3596 760 -3590
rect 1639 -3596 1642 -3590
rect 1646 -3596 1649 -3590
rect 1 -3607 7 -3601
rect 8 -3607 14 -3601
rect 15 -3607 21 -3601
rect 22 -3607 28 -3601
rect 29 -3607 35 -3601
rect 36 -3607 42 -3601
rect 43 -3607 49 -3601
rect 50 -3607 56 -3601
rect 57 -3607 63 -3601
rect 64 -3607 70 -3601
rect 71 -3607 77 -3601
rect 78 -3607 84 -3601
rect 85 -3607 91 -3601
rect 92 -3607 98 -3601
rect 99 -3607 105 -3601
rect 106 -3607 112 -3601
rect 113 -3607 119 -3601
rect 120 -3607 126 -3601
rect 127 -3607 133 -3601
rect 134 -3607 140 -3601
rect 141 -3607 147 -3601
rect 148 -3607 154 -3601
rect 155 -3607 161 -3601
rect 162 -3607 168 -3601
rect 169 -3607 175 -3601
rect 176 -3607 182 -3601
rect 183 -3607 189 -3601
rect 190 -3607 196 -3601
rect 197 -3607 203 -3601
rect 204 -3607 210 -3601
rect 211 -3607 217 -3601
rect 218 -3607 224 -3601
rect 225 -3607 231 -3601
rect 232 -3607 238 -3601
rect 239 -3607 245 -3601
rect 246 -3607 252 -3601
rect 393 -3607 396 -3601
rect 400 -3607 403 -3601
rect 603 -3607 606 -3601
rect 610 -3607 613 -3601
rect 701 -3607 707 -3601
rect 757 -3607 760 -3601
rect 1639 -3607 1642 -3601
rect 1646 -3607 1649 -3601
rect 1 -3618 7 -3612
rect 8 -3618 14 -3612
rect 15 -3618 21 -3612
rect 22 -3618 28 -3612
rect 29 -3618 35 -3612
rect 36 -3618 42 -3612
rect 43 -3618 49 -3612
rect 50 -3618 56 -3612
rect 57 -3618 63 -3612
rect 64 -3618 70 -3612
rect 71 -3618 77 -3612
rect 78 -3618 84 -3612
rect 85 -3618 91 -3612
rect 92 -3618 98 -3612
rect 99 -3618 105 -3612
rect 106 -3618 112 -3612
rect 113 -3618 119 -3612
rect 120 -3618 126 -3612
rect 127 -3618 133 -3612
rect 134 -3618 140 -3612
rect 141 -3618 147 -3612
rect 148 -3618 154 -3612
rect 155 -3618 161 -3612
rect 162 -3618 168 -3612
rect 169 -3618 175 -3612
rect 176 -3618 182 -3612
rect 183 -3618 189 -3612
rect 190 -3618 196 -3612
rect 197 -3618 203 -3612
rect 204 -3618 210 -3612
rect 211 -3618 217 -3612
rect 218 -3618 224 -3612
rect 225 -3618 231 -3612
rect 232 -3618 238 -3612
rect 239 -3618 245 -3612
rect 393 -3618 396 -3612
rect 400 -3618 403 -3612
rect 603 -3618 606 -3612
rect 610 -3618 613 -3612
rect 694 -3618 697 -3612
rect 757 -3618 760 -3612
rect 1639 -3618 1645 -3612
rect 1646 -3618 1649 -3612
rect 1 -3629 7 -3623
rect 8 -3629 14 -3623
rect 15 -3629 21 -3623
rect 22 -3629 28 -3623
rect 29 -3629 35 -3623
rect 36 -3629 42 -3623
rect 43 -3629 49 -3623
rect 50 -3629 56 -3623
rect 57 -3629 63 -3623
rect 64 -3629 70 -3623
rect 71 -3629 77 -3623
rect 78 -3629 84 -3623
rect 85 -3629 91 -3623
rect 92 -3629 98 -3623
rect 99 -3629 105 -3623
rect 106 -3629 112 -3623
rect 113 -3629 119 -3623
rect 120 -3629 126 -3623
rect 127 -3629 133 -3623
rect 134 -3629 140 -3623
rect 141 -3629 147 -3623
rect 148 -3629 154 -3623
rect 155 -3629 161 -3623
rect 162 -3629 168 -3623
rect 169 -3629 175 -3623
rect 176 -3629 182 -3623
rect 183 -3629 189 -3623
rect 190 -3629 196 -3623
rect 197 -3629 203 -3623
rect 204 -3629 210 -3623
rect 211 -3629 217 -3623
rect 218 -3629 224 -3623
rect 225 -3629 231 -3623
rect 232 -3629 238 -3623
rect 393 -3629 396 -3623
rect 400 -3629 403 -3623
rect 603 -3629 606 -3623
rect 610 -3629 613 -3623
rect 694 -3629 697 -3623
rect 757 -3629 763 -3623
rect 764 -3629 767 -3623
rect 1 -3640 7 -3634
rect 8 -3640 14 -3634
rect 15 -3640 21 -3634
rect 22 -3640 28 -3634
rect 29 -3640 35 -3634
rect 36 -3640 42 -3634
rect 43 -3640 49 -3634
rect 50 -3640 56 -3634
rect 57 -3640 63 -3634
rect 64 -3640 70 -3634
rect 71 -3640 77 -3634
rect 78 -3640 84 -3634
rect 85 -3640 91 -3634
rect 92 -3640 98 -3634
rect 99 -3640 105 -3634
rect 106 -3640 112 -3634
rect 113 -3640 119 -3634
rect 120 -3640 126 -3634
rect 127 -3640 133 -3634
rect 134 -3640 140 -3634
rect 141 -3640 147 -3634
rect 148 -3640 154 -3634
rect 155 -3640 161 -3634
rect 162 -3640 168 -3634
rect 169 -3640 175 -3634
rect 176 -3640 182 -3634
rect 183 -3640 189 -3634
rect 190 -3640 196 -3634
rect 197 -3640 203 -3634
rect 204 -3640 210 -3634
rect 211 -3640 217 -3634
rect 218 -3640 224 -3634
rect 225 -3640 231 -3634
rect 232 -3640 238 -3634
rect 393 -3640 396 -3634
rect 400 -3640 403 -3634
rect 603 -3640 606 -3634
rect 610 -3640 613 -3634
rect 694 -3640 697 -3634
rect 1 -3651 7 -3645
rect 8 -3651 14 -3645
rect 15 -3651 21 -3645
rect 22 -3651 28 -3645
rect 29 -3651 35 -3645
rect 36 -3651 42 -3645
rect 43 -3651 49 -3645
rect 50 -3651 56 -3645
rect 57 -3651 63 -3645
rect 64 -3651 70 -3645
rect 71 -3651 77 -3645
rect 78 -3651 84 -3645
rect 85 -3651 91 -3645
rect 92 -3651 98 -3645
rect 99 -3651 105 -3645
rect 106 -3651 112 -3645
rect 113 -3651 119 -3645
rect 120 -3651 126 -3645
rect 127 -3651 133 -3645
rect 134 -3651 140 -3645
rect 141 -3651 147 -3645
rect 148 -3651 154 -3645
rect 155 -3651 161 -3645
rect 162 -3651 168 -3645
rect 169 -3651 175 -3645
rect 176 -3651 182 -3645
rect 183 -3651 189 -3645
rect 190 -3651 196 -3645
rect 197 -3651 203 -3645
rect 204 -3651 210 -3645
rect 211 -3651 217 -3645
rect 218 -3651 224 -3645
rect 225 -3651 231 -3645
rect 232 -3651 238 -3645
rect 239 -3651 245 -3645
rect 246 -3651 252 -3645
rect 253 -3651 259 -3645
rect 260 -3651 266 -3645
rect 267 -3651 273 -3645
rect 393 -3651 396 -3645
rect 400 -3651 403 -3645
rect 603 -3651 606 -3645
rect 610 -3651 613 -3645
rect 694 -3651 697 -3645
rect 1 -3666 7 -3660
rect 8 -3666 14 -3660
rect 15 -3666 21 -3660
rect 22 -3666 28 -3660
rect 29 -3666 35 -3660
rect 36 -3666 42 -3660
rect 43 -3666 49 -3660
rect 50 -3666 56 -3660
rect 57 -3666 63 -3660
rect 64 -3666 70 -3660
rect 71 -3666 77 -3660
rect 78 -3666 84 -3660
rect 85 -3666 91 -3660
rect 92 -3666 98 -3660
rect 99 -3666 105 -3660
rect 106 -3666 112 -3660
rect 113 -3666 119 -3660
rect 120 -3666 126 -3660
rect 127 -3666 133 -3660
rect 134 -3666 140 -3660
rect 141 -3666 147 -3660
rect 148 -3666 154 -3660
rect 155 -3666 161 -3660
rect 162 -3666 168 -3660
rect 169 -3666 175 -3660
rect 176 -3666 182 -3660
rect 183 -3666 189 -3660
rect 190 -3666 196 -3660
rect 197 -3666 203 -3660
rect 204 -3666 210 -3660
rect 393 -3666 399 -3660
rect 400 -3666 403 -3660
rect 603 -3666 606 -3660
rect 610 -3666 616 -3660
rect 694 -3666 700 -3660
<< polysilicon >>
rect 212 -27 213 -25
rect 254 -21 255 -19
rect 254 -27 255 -25
rect 352 -21 353 -19
rect 352 -27 353 -25
rect 397 -21 398 -19
rect 397 -27 398 -25
rect 415 -21 416 -19
rect 422 -21 423 -19
rect 422 -27 423 -25
rect 432 -21 433 -19
rect 432 -27 433 -25
rect 446 -27 447 -25
rect 485 -21 486 -19
rect 485 -27 486 -25
rect 548 -21 549 -19
rect 548 -27 549 -25
rect 555 -21 556 -19
rect 572 -21 573 -19
rect 569 -27 570 -25
rect 572 -27 573 -25
rect 576 -21 577 -19
rect 576 -27 577 -25
rect 583 -21 584 -19
rect 583 -27 584 -25
rect 604 -21 605 -19
rect 604 -27 605 -25
rect 611 -21 612 -19
rect 611 -27 612 -25
rect 618 -21 619 -19
rect 618 -27 619 -25
rect 625 -21 626 -19
rect 625 -27 626 -25
rect 632 -21 633 -19
rect 635 -21 636 -19
rect 639 -21 640 -19
rect 639 -27 640 -25
rect 646 -21 647 -19
rect 646 -27 647 -25
rect 653 -27 654 -25
rect 656 -27 657 -25
rect 663 -21 664 -19
rect 660 -27 661 -25
rect 681 -21 682 -19
rect 681 -27 682 -25
rect 688 -21 689 -19
rect 688 -27 689 -25
rect 705 -21 706 -19
rect 702 -27 703 -25
rect 709 -21 710 -19
rect 709 -27 710 -25
rect 716 -21 717 -19
rect 716 -27 717 -25
rect 730 -21 731 -19
rect 730 -27 731 -25
rect 765 -21 766 -19
rect 768 -27 769 -25
rect 772 -21 773 -19
rect 772 -27 773 -25
rect 796 -21 797 -19
rect 800 -21 801 -19
rect 803 -21 804 -19
rect 810 -21 811 -19
rect 807 -27 808 -25
rect 810 -27 811 -25
rect 814 -21 815 -19
rect 814 -27 815 -25
rect 821 -21 822 -19
rect 824 -21 825 -19
rect 828 -21 829 -19
rect 828 -27 829 -25
rect 835 -21 836 -19
rect 835 -27 836 -25
rect 842 -21 843 -19
rect 845 -21 846 -19
rect 842 -27 843 -25
rect 852 -21 853 -19
rect 849 -27 850 -25
rect 859 -21 860 -19
rect 863 -21 864 -19
rect 863 -27 864 -25
rect 870 -21 871 -19
rect 870 -27 871 -25
rect 884 -21 885 -19
rect 887 -21 888 -19
rect 887 -27 888 -25
rect 891 -21 892 -19
rect 891 -27 892 -25
rect 898 -27 899 -25
rect 915 -21 916 -19
rect 912 -27 913 -25
rect 915 -27 916 -25
rect 919 -21 920 -19
rect 919 -27 920 -25
rect 961 -21 962 -19
rect 961 -27 962 -25
rect 968 -21 969 -19
rect 968 -27 969 -25
rect 978 -21 979 -19
rect 978 -27 979 -25
rect 982 -21 983 -19
rect 982 -27 983 -25
rect 989 -21 990 -19
rect 989 -27 990 -25
rect 1038 -21 1039 -19
rect 1038 -27 1039 -25
rect 1073 -21 1074 -19
rect 1073 -27 1074 -25
rect 1087 -21 1088 -19
rect 1087 -27 1088 -25
rect 1094 -21 1095 -19
rect 1094 -27 1095 -25
rect 1125 -21 1126 -19
rect 1129 -21 1130 -19
rect 1132 -27 1133 -25
rect 1206 -21 1207 -19
rect 1206 -27 1207 -25
rect 1437 -21 1438 -19
rect 1437 -27 1438 -25
rect 1440 -27 1441 -25
rect 1629 -27 1630 -25
rect 184 -68 185 -66
rect 184 -74 185 -72
rect 198 -68 199 -66
rect 198 -74 199 -72
rect 240 -68 241 -66
rect 240 -74 241 -72
rect 275 -68 276 -66
rect 275 -74 276 -72
rect 296 -68 297 -66
rect 296 -74 297 -72
rect 313 -68 314 -66
rect 310 -74 311 -72
rect 317 -68 318 -66
rect 317 -74 318 -72
rect 355 -68 356 -66
rect 352 -74 353 -72
rect 394 -68 395 -66
rect 394 -74 395 -72
rect 404 -68 405 -66
rect 401 -74 402 -72
rect 404 -74 405 -72
rect 408 -74 409 -72
rect 411 -74 412 -72
rect 415 -68 416 -66
rect 415 -74 416 -72
rect 422 -68 423 -66
rect 422 -74 423 -72
rect 464 -68 465 -66
rect 464 -74 465 -72
rect 471 -68 472 -66
rect 471 -74 472 -72
rect 478 -68 479 -66
rect 478 -74 479 -72
rect 485 -68 486 -66
rect 485 -74 486 -72
rect 492 -68 493 -66
rect 492 -74 493 -72
rect 499 -68 500 -66
rect 499 -74 500 -72
rect 506 -68 507 -66
rect 506 -74 507 -72
rect 520 -68 521 -66
rect 520 -74 521 -72
rect 534 -68 535 -66
rect 534 -74 535 -72
rect 541 -74 542 -72
rect 544 -74 545 -72
rect 548 -68 549 -66
rect 548 -74 549 -72
rect 565 -68 566 -66
rect 565 -74 566 -72
rect 569 -68 570 -66
rect 569 -74 570 -72
rect 583 -68 584 -66
rect 583 -74 584 -72
rect 590 -68 591 -66
rect 590 -74 591 -72
rect 597 -68 598 -66
rect 597 -74 598 -72
rect 604 -68 605 -66
rect 604 -74 605 -72
rect 611 -68 612 -66
rect 611 -74 612 -72
rect 618 -68 619 -66
rect 618 -74 619 -72
rect 639 -68 640 -66
rect 639 -74 640 -72
rect 646 -68 647 -66
rect 646 -74 647 -72
rect 653 -68 654 -66
rect 656 -74 657 -72
rect 660 -68 661 -66
rect 660 -74 661 -72
rect 667 -68 668 -66
rect 667 -74 668 -72
rect 674 -68 675 -66
rect 677 -68 678 -66
rect 677 -74 678 -72
rect 681 -68 682 -66
rect 681 -74 682 -72
rect 688 -68 689 -66
rect 688 -74 689 -72
rect 695 -68 696 -66
rect 702 -68 703 -66
rect 702 -74 703 -72
rect 709 -68 710 -66
rect 709 -74 710 -72
rect 716 -68 717 -66
rect 716 -74 717 -72
rect 723 -68 724 -66
rect 723 -74 724 -72
rect 730 -68 731 -66
rect 730 -74 731 -72
rect 737 -68 738 -66
rect 740 -68 741 -66
rect 744 -68 745 -66
rect 744 -74 745 -72
rect 751 -68 752 -66
rect 751 -74 752 -72
rect 758 -68 759 -66
rect 758 -74 759 -72
rect 765 -68 766 -66
rect 765 -74 766 -72
rect 772 -68 773 -66
rect 772 -74 773 -72
rect 779 -68 780 -66
rect 779 -74 780 -72
rect 789 -74 790 -72
rect 793 -68 794 -66
rect 793 -74 794 -72
rect 800 -68 801 -66
rect 803 -68 804 -66
rect 800 -74 801 -72
rect 807 -68 808 -66
rect 807 -74 808 -72
rect 814 -68 815 -66
rect 814 -74 815 -72
rect 821 -68 822 -66
rect 821 -74 822 -72
rect 828 -68 829 -66
rect 828 -74 829 -72
rect 835 -68 836 -66
rect 835 -74 836 -72
rect 842 -68 843 -66
rect 842 -74 843 -72
rect 849 -68 850 -66
rect 852 -68 853 -66
rect 852 -74 853 -72
rect 856 -68 857 -66
rect 856 -74 857 -72
rect 859 -74 860 -72
rect 863 -68 864 -66
rect 863 -74 864 -72
rect 870 -68 871 -66
rect 870 -74 871 -72
rect 877 -68 878 -66
rect 877 -74 878 -72
rect 884 -68 885 -66
rect 887 -68 888 -66
rect 891 -68 892 -66
rect 891 -74 892 -72
rect 901 -68 902 -66
rect 898 -74 899 -72
rect 908 -68 909 -66
rect 908 -74 909 -72
rect 912 -68 913 -66
rect 912 -74 913 -72
rect 919 -68 920 -66
rect 919 -74 920 -72
rect 926 -68 927 -66
rect 926 -74 927 -72
rect 933 -68 934 -66
rect 933 -74 934 -72
rect 940 -68 941 -66
rect 943 -74 944 -72
rect 947 -68 948 -66
rect 947 -74 948 -72
rect 954 -74 955 -72
rect 957 -74 958 -72
rect 961 -68 962 -66
rect 961 -74 962 -72
rect 968 -68 969 -66
rect 968 -74 969 -72
rect 975 -68 976 -66
rect 975 -74 976 -72
rect 982 -68 983 -66
rect 982 -74 983 -72
rect 989 -68 990 -66
rect 989 -74 990 -72
rect 996 -74 997 -72
rect 999 -74 1000 -72
rect 1003 -68 1004 -66
rect 1003 -74 1004 -72
rect 1010 -68 1011 -66
rect 1010 -74 1011 -72
rect 1017 -68 1018 -66
rect 1017 -74 1018 -72
rect 1024 -68 1025 -66
rect 1024 -74 1025 -72
rect 1027 -74 1028 -72
rect 1031 -68 1032 -66
rect 1031 -74 1032 -72
rect 1038 -68 1039 -66
rect 1038 -74 1039 -72
rect 1045 -68 1046 -66
rect 1045 -74 1046 -72
rect 1052 -68 1053 -66
rect 1052 -74 1053 -72
rect 1059 -68 1060 -66
rect 1059 -74 1060 -72
rect 1066 -68 1067 -66
rect 1069 -68 1070 -66
rect 1073 -68 1074 -66
rect 1073 -74 1074 -72
rect 1080 -68 1081 -66
rect 1080 -74 1081 -72
rect 1087 -68 1088 -66
rect 1087 -74 1088 -72
rect 1094 -68 1095 -66
rect 1094 -74 1095 -72
rect 1101 -68 1102 -66
rect 1101 -74 1102 -72
rect 1108 -68 1109 -66
rect 1111 -74 1112 -72
rect 1115 -68 1116 -66
rect 1118 -74 1119 -72
rect 1125 -68 1126 -66
rect 1125 -74 1126 -72
rect 1150 -68 1151 -66
rect 1150 -74 1151 -72
rect 1167 -74 1168 -72
rect 1178 -68 1179 -66
rect 1178 -74 1179 -72
rect 1213 -68 1214 -66
rect 1213 -74 1214 -72
rect 1220 -68 1221 -66
rect 1220 -74 1221 -72
rect 1227 -74 1228 -72
rect 1234 -68 1235 -66
rect 1234 -74 1235 -72
rect 1237 -74 1238 -72
rect 1290 -68 1291 -66
rect 1290 -74 1291 -72
rect 1321 -68 1322 -66
rect 1321 -74 1322 -72
rect 1332 -68 1333 -66
rect 1332 -74 1333 -72
rect 1360 -68 1361 -66
rect 1360 -74 1361 -72
rect 1486 -68 1487 -66
rect 1486 -74 1487 -72
rect 1633 -68 1634 -66
rect 1633 -74 1634 -72
rect 1759 -68 1760 -66
rect 1759 -74 1760 -72
rect 58 -145 59 -143
rect 58 -151 59 -149
rect 65 -145 66 -143
rect 65 -151 66 -149
rect 72 -145 73 -143
rect 72 -151 73 -149
rect 79 -145 80 -143
rect 79 -151 80 -149
rect 86 -145 87 -143
rect 86 -151 87 -149
rect 93 -145 94 -143
rect 93 -151 94 -149
rect 100 -145 101 -143
rect 100 -151 101 -149
rect 107 -145 108 -143
rect 107 -151 108 -149
rect 114 -145 115 -143
rect 114 -151 115 -149
rect 121 -145 122 -143
rect 124 -145 125 -143
rect 124 -151 125 -149
rect 128 -145 129 -143
rect 128 -151 129 -149
rect 135 -145 136 -143
rect 135 -151 136 -149
rect 142 -145 143 -143
rect 145 -151 146 -149
rect 149 -145 150 -143
rect 152 -145 153 -143
rect 152 -151 153 -149
rect 156 -145 157 -143
rect 156 -151 157 -149
rect 163 -145 164 -143
rect 163 -151 164 -149
rect 170 -145 171 -143
rect 170 -151 171 -149
rect 177 -145 178 -143
rect 177 -151 178 -149
rect 184 -145 185 -143
rect 184 -151 185 -149
rect 191 -145 192 -143
rect 191 -151 192 -149
rect 198 -145 199 -143
rect 198 -151 199 -149
rect 205 -145 206 -143
rect 205 -151 206 -149
rect 212 -145 213 -143
rect 212 -151 213 -149
rect 219 -145 220 -143
rect 219 -151 220 -149
rect 226 -145 227 -143
rect 229 -145 230 -143
rect 226 -151 227 -149
rect 233 -145 234 -143
rect 236 -145 237 -143
rect 240 -145 241 -143
rect 240 -151 241 -149
rect 247 -145 248 -143
rect 247 -151 248 -149
rect 254 -151 255 -149
rect 257 -151 258 -149
rect 261 -145 262 -143
rect 264 -145 265 -143
rect 261 -151 262 -149
rect 268 -151 269 -149
rect 275 -145 276 -143
rect 275 -151 276 -149
rect 282 -145 283 -143
rect 282 -151 283 -149
rect 289 -145 290 -143
rect 289 -151 290 -149
rect 296 -145 297 -143
rect 296 -151 297 -149
rect 303 -145 304 -143
rect 303 -151 304 -149
rect 310 -145 311 -143
rect 310 -151 311 -149
rect 317 -145 318 -143
rect 317 -151 318 -149
rect 324 -145 325 -143
rect 324 -151 325 -149
rect 331 -145 332 -143
rect 331 -151 332 -149
rect 338 -145 339 -143
rect 338 -151 339 -149
rect 345 -145 346 -143
rect 345 -151 346 -149
rect 352 -145 353 -143
rect 352 -151 353 -149
rect 359 -145 360 -143
rect 359 -151 360 -149
rect 366 -145 367 -143
rect 366 -151 367 -149
rect 373 -145 374 -143
rect 373 -151 374 -149
rect 380 -145 381 -143
rect 380 -151 381 -149
rect 387 -145 388 -143
rect 390 -145 391 -143
rect 390 -151 391 -149
rect 394 -145 395 -143
rect 394 -151 395 -149
rect 401 -145 402 -143
rect 401 -151 402 -149
rect 408 -145 409 -143
rect 408 -151 409 -149
rect 415 -145 416 -143
rect 415 -151 416 -149
rect 422 -145 423 -143
rect 422 -151 423 -149
rect 429 -145 430 -143
rect 429 -151 430 -149
rect 436 -145 437 -143
rect 436 -151 437 -149
rect 443 -145 444 -143
rect 446 -145 447 -143
rect 450 -145 451 -143
rect 450 -151 451 -149
rect 457 -145 458 -143
rect 460 -145 461 -143
rect 460 -151 461 -149
rect 467 -145 468 -143
rect 467 -151 468 -149
rect 471 -145 472 -143
rect 474 -145 475 -143
rect 478 -145 479 -143
rect 478 -151 479 -149
rect 485 -145 486 -143
rect 485 -151 486 -149
rect 492 -145 493 -143
rect 492 -151 493 -149
rect 499 -145 500 -143
rect 499 -151 500 -149
rect 506 -145 507 -143
rect 506 -151 507 -149
rect 513 -145 514 -143
rect 513 -151 514 -149
rect 523 -145 524 -143
rect 520 -151 521 -149
rect 523 -151 524 -149
rect 527 -145 528 -143
rect 530 -145 531 -143
rect 527 -151 528 -149
rect 530 -151 531 -149
rect 534 -145 535 -143
rect 534 -151 535 -149
rect 541 -145 542 -143
rect 541 -151 542 -149
rect 548 -145 549 -143
rect 548 -151 549 -149
rect 555 -145 556 -143
rect 555 -151 556 -149
rect 562 -145 563 -143
rect 565 -145 566 -143
rect 565 -151 566 -149
rect 569 -145 570 -143
rect 569 -151 570 -149
rect 576 -145 577 -143
rect 576 -151 577 -149
rect 583 -145 584 -143
rect 583 -151 584 -149
rect 590 -145 591 -143
rect 590 -151 591 -149
rect 597 -145 598 -143
rect 600 -145 601 -143
rect 600 -151 601 -149
rect 604 -145 605 -143
rect 604 -151 605 -149
rect 611 -145 612 -143
rect 611 -151 612 -149
rect 618 -145 619 -143
rect 618 -151 619 -149
rect 625 -145 626 -143
rect 625 -151 626 -149
rect 632 -145 633 -143
rect 632 -151 633 -149
rect 639 -145 640 -143
rect 639 -151 640 -149
rect 649 -145 650 -143
rect 649 -151 650 -149
rect 653 -145 654 -143
rect 653 -151 654 -149
rect 660 -145 661 -143
rect 660 -151 661 -149
rect 667 -145 668 -143
rect 667 -151 668 -149
rect 674 -145 675 -143
rect 674 -151 675 -149
rect 681 -145 682 -143
rect 684 -151 685 -149
rect 688 -145 689 -143
rect 688 -151 689 -149
rect 698 -145 699 -143
rect 695 -151 696 -149
rect 698 -151 699 -149
rect 702 -145 703 -143
rect 702 -151 703 -149
rect 709 -145 710 -143
rect 709 -151 710 -149
rect 716 -145 717 -143
rect 716 -151 717 -149
rect 723 -145 724 -143
rect 723 -151 724 -149
rect 730 -145 731 -143
rect 733 -151 734 -149
rect 737 -145 738 -143
rect 740 -145 741 -143
rect 737 -151 738 -149
rect 744 -145 745 -143
rect 744 -151 745 -149
rect 751 -145 752 -143
rect 751 -151 752 -149
rect 758 -145 759 -143
rect 758 -151 759 -149
rect 765 -145 766 -143
rect 765 -151 766 -149
rect 768 -151 769 -149
rect 772 -145 773 -143
rect 772 -151 773 -149
rect 779 -145 780 -143
rect 779 -151 780 -149
rect 786 -145 787 -143
rect 786 -151 787 -149
rect 793 -145 794 -143
rect 793 -151 794 -149
rect 803 -145 804 -143
rect 800 -151 801 -149
rect 803 -151 804 -149
rect 807 -145 808 -143
rect 807 -151 808 -149
rect 814 -145 815 -143
rect 814 -151 815 -149
rect 821 -145 822 -143
rect 821 -151 822 -149
rect 828 -145 829 -143
rect 828 -151 829 -149
rect 835 -145 836 -143
rect 835 -151 836 -149
rect 838 -151 839 -149
rect 842 -145 843 -143
rect 842 -151 843 -149
rect 849 -145 850 -143
rect 849 -151 850 -149
rect 856 -145 857 -143
rect 856 -151 857 -149
rect 863 -145 864 -143
rect 863 -151 864 -149
rect 870 -145 871 -143
rect 870 -151 871 -149
rect 877 -145 878 -143
rect 877 -151 878 -149
rect 884 -145 885 -143
rect 884 -151 885 -149
rect 891 -145 892 -143
rect 891 -151 892 -149
rect 898 -145 899 -143
rect 898 -151 899 -149
rect 905 -145 906 -143
rect 905 -151 906 -149
rect 912 -145 913 -143
rect 912 -151 913 -149
rect 919 -145 920 -143
rect 919 -151 920 -149
rect 929 -151 930 -149
rect 933 -145 934 -143
rect 936 -151 937 -149
rect 940 -145 941 -143
rect 940 -151 941 -149
rect 947 -145 948 -143
rect 947 -151 948 -149
rect 950 -151 951 -149
rect 954 -145 955 -143
rect 954 -151 955 -149
rect 961 -151 962 -149
rect 968 -145 969 -143
rect 968 -151 969 -149
rect 975 -145 976 -143
rect 975 -151 976 -149
rect 982 -145 983 -143
rect 982 -151 983 -149
rect 989 -145 990 -143
rect 989 -151 990 -149
rect 996 -145 997 -143
rect 996 -151 997 -149
rect 1003 -145 1004 -143
rect 1003 -151 1004 -149
rect 1010 -145 1011 -143
rect 1010 -151 1011 -149
rect 1017 -145 1018 -143
rect 1017 -151 1018 -149
rect 1024 -145 1025 -143
rect 1024 -151 1025 -149
rect 1031 -145 1032 -143
rect 1031 -151 1032 -149
rect 1038 -145 1039 -143
rect 1038 -151 1039 -149
rect 1045 -145 1046 -143
rect 1045 -151 1046 -149
rect 1052 -145 1053 -143
rect 1052 -151 1053 -149
rect 1059 -145 1060 -143
rect 1059 -151 1060 -149
rect 1066 -145 1067 -143
rect 1066 -151 1067 -149
rect 1076 -145 1077 -143
rect 1073 -151 1074 -149
rect 1076 -151 1077 -149
rect 1080 -145 1081 -143
rect 1080 -151 1081 -149
rect 1087 -145 1088 -143
rect 1087 -151 1088 -149
rect 1090 -151 1091 -149
rect 1094 -145 1095 -143
rect 1094 -151 1095 -149
rect 1101 -145 1102 -143
rect 1101 -151 1102 -149
rect 1108 -145 1109 -143
rect 1108 -151 1109 -149
rect 1115 -145 1116 -143
rect 1115 -151 1116 -149
rect 1122 -145 1123 -143
rect 1122 -151 1123 -149
rect 1129 -145 1130 -143
rect 1129 -151 1130 -149
rect 1136 -145 1137 -143
rect 1136 -151 1137 -149
rect 1143 -145 1144 -143
rect 1143 -151 1144 -149
rect 1146 -151 1147 -149
rect 1150 -145 1151 -143
rect 1150 -151 1151 -149
rect 1157 -145 1158 -143
rect 1157 -151 1158 -149
rect 1164 -145 1165 -143
rect 1164 -151 1165 -149
rect 1171 -145 1172 -143
rect 1171 -151 1172 -149
rect 1174 -151 1175 -149
rect 1178 -145 1179 -143
rect 1178 -151 1179 -149
rect 1185 -145 1186 -143
rect 1185 -151 1186 -149
rect 1192 -145 1193 -143
rect 1192 -151 1193 -149
rect 1199 -145 1200 -143
rect 1199 -151 1200 -149
rect 1206 -145 1207 -143
rect 1206 -151 1207 -149
rect 1213 -145 1214 -143
rect 1213 -151 1214 -149
rect 1220 -145 1221 -143
rect 1220 -151 1221 -149
rect 1227 -145 1228 -143
rect 1227 -151 1228 -149
rect 1234 -145 1235 -143
rect 1234 -151 1235 -149
rect 1241 -145 1242 -143
rect 1241 -151 1242 -149
rect 1248 -145 1249 -143
rect 1248 -151 1249 -149
rect 1255 -145 1256 -143
rect 1255 -151 1256 -149
rect 1262 -151 1263 -149
rect 1265 -151 1266 -149
rect 1269 -145 1270 -143
rect 1269 -151 1270 -149
rect 1276 -145 1277 -143
rect 1276 -151 1277 -149
rect 1283 -145 1284 -143
rect 1283 -151 1284 -149
rect 1290 -145 1291 -143
rect 1290 -151 1291 -149
rect 1297 -145 1298 -143
rect 1297 -151 1298 -149
rect 1304 -145 1305 -143
rect 1304 -151 1305 -149
rect 1311 -145 1312 -143
rect 1311 -151 1312 -149
rect 1318 -145 1319 -143
rect 1318 -151 1319 -149
rect 1325 -145 1326 -143
rect 1325 -151 1326 -149
rect 1353 -145 1354 -143
rect 1353 -151 1354 -149
rect 1360 -145 1361 -143
rect 1360 -151 1361 -149
rect 1374 -145 1375 -143
rect 1374 -151 1375 -149
rect 1423 -145 1424 -143
rect 1423 -151 1424 -149
rect 1507 -145 1508 -143
rect 1507 -151 1508 -149
rect 1514 -145 1515 -143
rect 1514 -151 1515 -149
rect 1640 -145 1641 -143
rect 1640 -151 1641 -149
rect 1885 -145 1886 -143
rect 1885 -151 1886 -149
rect 16 -248 17 -246
rect 16 -254 17 -252
rect 23 -248 24 -246
rect 23 -254 24 -252
rect 30 -248 31 -246
rect 30 -254 31 -252
rect 37 -248 38 -246
rect 37 -254 38 -252
rect 44 -248 45 -246
rect 44 -254 45 -252
rect 51 -248 52 -246
rect 51 -254 52 -252
rect 58 -248 59 -246
rect 58 -254 59 -252
rect 72 -248 73 -246
rect 72 -254 73 -252
rect 79 -248 80 -246
rect 79 -254 80 -252
rect 89 -248 90 -246
rect 89 -254 90 -252
rect 93 -248 94 -246
rect 93 -254 94 -252
rect 100 -248 101 -246
rect 100 -254 101 -252
rect 107 -248 108 -246
rect 107 -254 108 -252
rect 117 -248 118 -246
rect 117 -254 118 -252
rect 121 -248 122 -246
rect 121 -254 122 -252
rect 128 -248 129 -246
rect 128 -254 129 -252
rect 135 -248 136 -246
rect 135 -254 136 -252
rect 138 -254 139 -252
rect 142 -248 143 -246
rect 142 -254 143 -252
rect 149 -248 150 -246
rect 149 -254 150 -252
rect 156 -248 157 -246
rect 159 -248 160 -246
rect 156 -254 157 -252
rect 163 -248 164 -246
rect 163 -254 164 -252
rect 170 -248 171 -246
rect 170 -254 171 -252
rect 177 -248 178 -246
rect 177 -254 178 -252
rect 184 -248 185 -246
rect 184 -254 185 -252
rect 194 -248 195 -246
rect 194 -254 195 -252
rect 198 -248 199 -246
rect 201 -248 202 -246
rect 205 -254 206 -252
rect 208 -254 209 -252
rect 212 -248 213 -246
rect 212 -254 213 -252
rect 219 -248 220 -246
rect 219 -254 220 -252
rect 226 -248 227 -246
rect 226 -254 227 -252
rect 233 -248 234 -246
rect 233 -254 234 -252
rect 240 -248 241 -246
rect 243 -248 244 -246
rect 240 -254 241 -252
rect 247 -248 248 -246
rect 247 -254 248 -252
rect 254 -248 255 -246
rect 254 -254 255 -252
rect 261 -248 262 -246
rect 261 -254 262 -252
rect 271 -248 272 -246
rect 268 -254 269 -252
rect 271 -254 272 -252
rect 275 -248 276 -246
rect 275 -254 276 -252
rect 282 -248 283 -246
rect 282 -254 283 -252
rect 289 -248 290 -246
rect 289 -254 290 -252
rect 296 -248 297 -246
rect 299 -254 300 -252
rect 303 -248 304 -246
rect 303 -254 304 -252
rect 310 -248 311 -246
rect 310 -254 311 -252
rect 313 -254 314 -252
rect 317 -248 318 -246
rect 317 -254 318 -252
rect 324 -248 325 -246
rect 324 -254 325 -252
rect 331 -248 332 -246
rect 331 -254 332 -252
rect 338 -248 339 -246
rect 338 -254 339 -252
rect 345 -248 346 -246
rect 345 -254 346 -252
rect 352 -248 353 -246
rect 352 -254 353 -252
rect 359 -248 360 -246
rect 359 -254 360 -252
rect 366 -248 367 -246
rect 366 -254 367 -252
rect 373 -248 374 -246
rect 373 -254 374 -252
rect 380 -248 381 -246
rect 380 -254 381 -252
rect 387 -248 388 -246
rect 387 -254 388 -252
rect 394 -248 395 -246
rect 394 -254 395 -252
rect 401 -248 402 -246
rect 401 -254 402 -252
rect 408 -248 409 -246
rect 408 -254 409 -252
rect 415 -248 416 -246
rect 415 -254 416 -252
rect 422 -248 423 -246
rect 422 -254 423 -252
rect 429 -248 430 -246
rect 429 -254 430 -252
rect 436 -248 437 -246
rect 439 -248 440 -246
rect 436 -254 437 -252
rect 439 -254 440 -252
rect 443 -248 444 -246
rect 443 -254 444 -252
rect 450 -248 451 -246
rect 450 -254 451 -252
rect 457 -248 458 -246
rect 457 -254 458 -252
rect 464 -254 465 -252
rect 467 -254 468 -252
rect 471 -248 472 -246
rect 471 -254 472 -252
rect 478 -248 479 -246
rect 478 -254 479 -252
rect 485 -248 486 -246
rect 485 -254 486 -252
rect 492 -248 493 -246
rect 492 -254 493 -252
rect 499 -248 500 -246
rect 499 -254 500 -252
rect 506 -248 507 -246
rect 506 -254 507 -252
rect 513 -248 514 -246
rect 513 -254 514 -252
rect 520 -248 521 -246
rect 523 -248 524 -246
rect 523 -254 524 -252
rect 527 -248 528 -246
rect 527 -254 528 -252
rect 534 -248 535 -246
rect 537 -248 538 -246
rect 534 -254 535 -252
rect 537 -254 538 -252
rect 541 -248 542 -246
rect 541 -254 542 -252
rect 548 -248 549 -246
rect 548 -254 549 -252
rect 555 -248 556 -246
rect 555 -254 556 -252
rect 562 -248 563 -246
rect 562 -254 563 -252
rect 569 -248 570 -246
rect 569 -254 570 -252
rect 576 -248 577 -246
rect 576 -254 577 -252
rect 583 -248 584 -246
rect 583 -254 584 -252
rect 593 -248 594 -246
rect 590 -254 591 -252
rect 597 -248 598 -246
rect 597 -254 598 -252
rect 604 -248 605 -246
rect 604 -254 605 -252
rect 611 -248 612 -246
rect 611 -254 612 -252
rect 621 -248 622 -246
rect 618 -254 619 -252
rect 621 -254 622 -252
rect 625 -248 626 -246
rect 625 -254 626 -252
rect 632 -248 633 -246
rect 632 -254 633 -252
rect 639 -248 640 -246
rect 639 -254 640 -252
rect 646 -248 647 -246
rect 646 -254 647 -252
rect 653 -248 654 -246
rect 653 -254 654 -252
rect 660 -248 661 -246
rect 660 -254 661 -252
rect 667 -248 668 -246
rect 667 -254 668 -252
rect 674 -248 675 -246
rect 674 -254 675 -252
rect 681 -248 682 -246
rect 681 -254 682 -252
rect 688 -248 689 -246
rect 688 -254 689 -252
rect 695 -248 696 -246
rect 695 -254 696 -252
rect 705 -248 706 -246
rect 702 -254 703 -252
rect 705 -254 706 -252
rect 709 -248 710 -246
rect 712 -248 713 -246
rect 709 -254 710 -252
rect 712 -254 713 -252
rect 716 -248 717 -246
rect 716 -254 717 -252
rect 723 -248 724 -246
rect 723 -254 724 -252
rect 730 -248 731 -246
rect 730 -254 731 -252
rect 737 -248 738 -246
rect 737 -254 738 -252
rect 744 -248 745 -246
rect 744 -254 745 -252
rect 751 -248 752 -246
rect 751 -254 752 -252
rect 758 -248 759 -246
rect 758 -254 759 -252
rect 765 -248 766 -246
rect 765 -254 766 -252
rect 772 -248 773 -246
rect 772 -254 773 -252
rect 779 -248 780 -246
rect 779 -254 780 -252
rect 786 -248 787 -246
rect 786 -254 787 -252
rect 793 -248 794 -246
rect 793 -254 794 -252
rect 800 -248 801 -246
rect 800 -254 801 -252
rect 807 -248 808 -246
rect 807 -254 808 -252
rect 814 -248 815 -246
rect 814 -254 815 -252
rect 821 -248 822 -246
rect 821 -254 822 -252
rect 828 -248 829 -246
rect 828 -254 829 -252
rect 835 -248 836 -246
rect 835 -254 836 -252
rect 842 -248 843 -246
rect 842 -254 843 -252
rect 849 -248 850 -246
rect 849 -254 850 -252
rect 856 -248 857 -246
rect 856 -254 857 -252
rect 863 -248 864 -246
rect 863 -254 864 -252
rect 870 -248 871 -246
rect 870 -254 871 -252
rect 877 -248 878 -246
rect 877 -254 878 -252
rect 884 -248 885 -246
rect 887 -248 888 -246
rect 887 -254 888 -252
rect 894 -248 895 -246
rect 894 -254 895 -252
rect 898 -248 899 -246
rect 898 -254 899 -252
rect 905 -248 906 -246
rect 905 -254 906 -252
rect 915 -248 916 -246
rect 912 -254 913 -252
rect 915 -254 916 -252
rect 919 -248 920 -246
rect 919 -254 920 -252
rect 926 -248 927 -246
rect 926 -254 927 -252
rect 933 -248 934 -246
rect 933 -254 934 -252
rect 940 -248 941 -246
rect 940 -254 941 -252
rect 947 -248 948 -246
rect 947 -254 948 -252
rect 954 -248 955 -246
rect 954 -254 955 -252
rect 961 -248 962 -246
rect 961 -254 962 -252
rect 968 -248 969 -246
rect 968 -254 969 -252
rect 975 -248 976 -246
rect 975 -254 976 -252
rect 982 -248 983 -246
rect 982 -254 983 -252
rect 989 -248 990 -246
rect 992 -254 993 -252
rect 999 -248 1000 -246
rect 996 -254 997 -252
rect 1003 -248 1004 -246
rect 1003 -254 1004 -252
rect 1010 -248 1011 -246
rect 1013 -248 1014 -246
rect 1010 -254 1011 -252
rect 1017 -248 1018 -246
rect 1017 -254 1018 -252
rect 1024 -248 1025 -246
rect 1024 -254 1025 -252
rect 1031 -248 1032 -246
rect 1031 -254 1032 -252
rect 1038 -248 1039 -246
rect 1038 -254 1039 -252
rect 1045 -248 1046 -246
rect 1045 -254 1046 -252
rect 1052 -248 1053 -246
rect 1052 -254 1053 -252
rect 1059 -248 1060 -246
rect 1059 -254 1060 -252
rect 1066 -248 1067 -246
rect 1066 -254 1067 -252
rect 1073 -248 1074 -246
rect 1073 -254 1074 -252
rect 1080 -248 1081 -246
rect 1080 -254 1081 -252
rect 1087 -248 1088 -246
rect 1087 -254 1088 -252
rect 1094 -248 1095 -246
rect 1094 -254 1095 -252
rect 1101 -248 1102 -246
rect 1101 -254 1102 -252
rect 1108 -248 1109 -246
rect 1108 -254 1109 -252
rect 1115 -248 1116 -246
rect 1115 -254 1116 -252
rect 1122 -248 1123 -246
rect 1122 -254 1123 -252
rect 1129 -248 1130 -246
rect 1129 -254 1130 -252
rect 1136 -248 1137 -246
rect 1136 -254 1137 -252
rect 1143 -248 1144 -246
rect 1143 -254 1144 -252
rect 1150 -248 1151 -246
rect 1150 -254 1151 -252
rect 1153 -254 1154 -252
rect 1157 -248 1158 -246
rect 1157 -254 1158 -252
rect 1164 -248 1165 -246
rect 1164 -254 1165 -252
rect 1171 -248 1172 -246
rect 1171 -254 1172 -252
rect 1178 -248 1179 -246
rect 1178 -254 1179 -252
rect 1185 -248 1186 -246
rect 1185 -254 1186 -252
rect 1192 -248 1193 -246
rect 1192 -254 1193 -252
rect 1199 -248 1200 -246
rect 1202 -248 1203 -246
rect 1206 -248 1207 -246
rect 1206 -254 1207 -252
rect 1213 -248 1214 -246
rect 1216 -248 1217 -246
rect 1213 -254 1214 -252
rect 1220 -248 1221 -246
rect 1220 -254 1221 -252
rect 1227 -248 1228 -246
rect 1227 -254 1228 -252
rect 1234 -248 1235 -246
rect 1234 -254 1235 -252
rect 1241 -248 1242 -246
rect 1241 -254 1242 -252
rect 1248 -248 1249 -246
rect 1248 -254 1249 -252
rect 1255 -248 1256 -246
rect 1255 -254 1256 -252
rect 1262 -248 1263 -246
rect 1262 -254 1263 -252
rect 1269 -248 1270 -246
rect 1269 -254 1270 -252
rect 1276 -248 1277 -246
rect 1276 -254 1277 -252
rect 1283 -248 1284 -246
rect 1283 -254 1284 -252
rect 1290 -248 1291 -246
rect 1290 -254 1291 -252
rect 1297 -248 1298 -246
rect 1297 -254 1298 -252
rect 1304 -248 1305 -246
rect 1304 -254 1305 -252
rect 1311 -248 1312 -246
rect 1311 -254 1312 -252
rect 1318 -248 1319 -246
rect 1318 -254 1319 -252
rect 1325 -248 1326 -246
rect 1328 -248 1329 -246
rect 1332 -248 1333 -246
rect 1332 -254 1333 -252
rect 1339 -248 1340 -246
rect 1339 -254 1340 -252
rect 1346 -248 1347 -246
rect 1346 -254 1347 -252
rect 1353 -248 1354 -246
rect 1353 -254 1354 -252
rect 1360 -248 1361 -246
rect 1360 -254 1361 -252
rect 1367 -248 1368 -246
rect 1367 -254 1368 -252
rect 1374 -248 1375 -246
rect 1374 -254 1375 -252
rect 1381 -248 1382 -246
rect 1381 -254 1382 -252
rect 1388 -248 1389 -246
rect 1388 -254 1389 -252
rect 1395 -248 1396 -246
rect 1395 -254 1396 -252
rect 1402 -248 1403 -246
rect 1402 -254 1403 -252
rect 1409 -248 1410 -246
rect 1409 -254 1410 -252
rect 1416 -248 1417 -246
rect 1416 -254 1417 -252
rect 1423 -248 1424 -246
rect 1423 -254 1424 -252
rect 1430 -248 1431 -246
rect 1430 -254 1431 -252
rect 1437 -248 1438 -246
rect 1437 -254 1438 -252
rect 1444 -248 1445 -246
rect 1444 -254 1445 -252
rect 1451 -248 1452 -246
rect 1451 -254 1452 -252
rect 1458 -248 1459 -246
rect 1458 -254 1459 -252
rect 1465 -248 1466 -246
rect 1465 -254 1466 -252
rect 1472 -248 1473 -246
rect 1472 -254 1473 -252
rect 1479 -248 1480 -246
rect 1479 -254 1480 -252
rect 1486 -248 1487 -246
rect 1486 -254 1487 -252
rect 1493 -248 1494 -246
rect 1493 -254 1494 -252
rect 1500 -248 1501 -246
rect 1500 -254 1501 -252
rect 1507 -248 1508 -246
rect 1507 -254 1508 -252
rect 1514 -248 1515 -246
rect 1514 -254 1515 -252
rect 1521 -248 1522 -246
rect 1521 -254 1522 -252
rect 1528 -248 1529 -246
rect 1528 -254 1529 -252
rect 1535 -248 1536 -246
rect 1535 -254 1536 -252
rect 1542 -248 1543 -246
rect 1542 -254 1543 -252
rect 1545 -254 1546 -252
rect 1549 -248 1550 -246
rect 1552 -254 1553 -252
rect 1556 -248 1557 -246
rect 1556 -254 1557 -252
rect 1566 -248 1567 -246
rect 1563 -254 1564 -252
rect 1570 -248 1571 -246
rect 1570 -254 1571 -252
rect 1577 -248 1578 -246
rect 1577 -254 1578 -252
rect 1584 -248 1585 -246
rect 1584 -254 1585 -252
rect 1591 -248 1592 -246
rect 1591 -254 1592 -252
rect 1612 -248 1613 -246
rect 1615 -248 1616 -246
rect 1612 -254 1613 -252
rect 1626 -248 1627 -246
rect 1626 -254 1627 -252
rect 1633 -248 1634 -246
rect 1633 -254 1634 -252
rect 1668 -248 1669 -246
rect 1668 -254 1669 -252
rect 1815 -248 1816 -246
rect 1815 -254 1816 -252
rect 1941 -248 1942 -246
rect 1941 -254 1942 -252
rect 16 -373 17 -371
rect 16 -379 17 -377
rect 23 -373 24 -371
rect 23 -379 24 -377
rect 30 -373 31 -371
rect 30 -379 31 -377
rect 37 -373 38 -371
rect 37 -379 38 -377
rect 47 -373 48 -371
rect 44 -379 45 -377
rect 51 -373 52 -371
rect 54 -373 55 -371
rect 54 -379 55 -377
rect 58 -373 59 -371
rect 58 -379 59 -377
rect 65 -373 66 -371
rect 65 -379 66 -377
rect 72 -373 73 -371
rect 72 -379 73 -377
rect 79 -373 80 -371
rect 79 -379 80 -377
rect 86 -373 87 -371
rect 86 -379 87 -377
rect 93 -373 94 -371
rect 93 -379 94 -377
rect 96 -379 97 -377
rect 100 -373 101 -371
rect 100 -379 101 -377
rect 107 -373 108 -371
rect 107 -379 108 -377
rect 114 -373 115 -371
rect 114 -379 115 -377
rect 121 -373 122 -371
rect 121 -379 122 -377
rect 128 -373 129 -371
rect 128 -379 129 -377
rect 135 -373 136 -371
rect 138 -373 139 -371
rect 142 -373 143 -371
rect 142 -379 143 -377
rect 149 -373 150 -371
rect 149 -379 150 -377
rect 156 -373 157 -371
rect 156 -379 157 -377
rect 163 -373 164 -371
rect 166 -373 167 -371
rect 163 -379 164 -377
rect 166 -379 167 -377
rect 170 -373 171 -371
rect 170 -379 171 -377
rect 177 -373 178 -371
rect 177 -379 178 -377
rect 187 -373 188 -371
rect 184 -379 185 -377
rect 187 -379 188 -377
rect 191 -373 192 -371
rect 191 -379 192 -377
rect 198 -373 199 -371
rect 198 -379 199 -377
rect 205 -373 206 -371
rect 205 -379 206 -377
rect 212 -373 213 -371
rect 212 -379 213 -377
rect 219 -373 220 -371
rect 219 -379 220 -377
rect 226 -373 227 -371
rect 226 -379 227 -377
rect 233 -373 234 -371
rect 233 -379 234 -377
rect 240 -373 241 -371
rect 243 -373 244 -371
rect 240 -379 241 -377
rect 247 -373 248 -371
rect 247 -379 248 -377
rect 254 -373 255 -371
rect 254 -379 255 -377
rect 261 -373 262 -371
rect 261 -379 262 -377
rect 268 -373 269 -371
rect 268 -379 269 -377
rect 275 -373 276 -371
rect 275 -379 276 -377
rect 282 -373 283 -371
rect 282 -379 283 -377
rect 289 -373 290 -371
rect 289 -379 290 -377
rect 296 -373 297 -371
rect 296 -379 297 -377
rect 303 -373 304 -371
rect 303 -379 304 -377
rect 310 -373 311 -371
rect 310 -379 311 -377
rect 317 -373 318 -371
rect 317 -379 318 -377
rect 324 -373 325 -371
rect 324 -379 325 -377
rect 331 -373 332 -371
rect 331 -379 332 -377
rect 338 -373 339 -371
rect 338 -379 339 -377
rect 345 -373 346 -371
rect 345 -379 346 -377
rect 352 -373 353 -371
rect 352 -379 353 -377
rect 359 -373 360 -371
rect 359 -379 360 -377
rect 366 -373 367 -371
rect 366 -379 367 -377
rect 373 -373 374 -371
rect 373 -379 374 -377
rect 380 -373 381 -371
rect 380 -379 381 -377
rect 387 -373 388 -371
rect 387 -379 388 -377
rect 394 -373 395 -371
rect 394 -379 395 -377
rect 401 -373 402 -371
rect 404 -373 405 -371
rect 401 -379 402 -377
rect 408 -373 409 -371
rect 408 -379 409 -377
rect 415 -373 416 -371
rect 415 -379 416 -377
rect 422 -373 423 -371
rect 422 -379 423 -377
rect 432 -373 433 -371
rect 429 -379 430 -377
rect 432 -379 433 -377
rect 436 -373 437 -371
rect 436 -379 437 -377
rect 443 -373 444 -371
rect 443 -379 444 -377
rect 446 -379 447 -377
rect 450 -373 451 -371
rect 450 -379 451 -377
rect 457 -373 458 -371
rect 457 -379 458 -377
rect 464 -373 465 -371
rect 464 -379 465 -377
rect 471 -373 472 -371
rect 471 -379 472 -377
rect 478 -373 479 -371
rect 481 -373 482 -371
rect 478 -379 479 -377
rect 481 -379 482 -377
rect 485 -373 486 -371
rect 485 -379 486 -377
rect 492 -373 493 -371
rect 492 -379 493 -377
rect 499 -373 500 -371
rect 499 -379 500 -377
rect 506 -373 507 -371
rect 506 -379 507 -377
rect 513 -373 514 -371
rect 513 -379 514 -377
rect 520 -373 521 -371
rect 520 -379 521 -377
rect 527 -373 528 -371
rect 527 -379 528 -377
rect 534 -373 535 -371
rect 534 -379 535 -377
rect 541 -373 542 -371
rect 541 -379 542 -377
rect 548 -373 549 -371
rect 548 -379 549 -377
rect 555 -373 556 -371
rect 555 -379 556 -377
rect 562 -373 563 -371
rect 562 -379 563 -377
rect 569 -373 570 -371
rect 569 -379 570 -377
rect 576 -373 577 -371
rect 576 -379 577 -377
rect 583 -373 584 -371
rect 583 -379 584 -377
rect 590 -373 591 -371
rect 590 -379 591 -377
rect 597 -373 598 -371
rect 597 -379 598 -377
rect 604 -373 605 -371
rect 604 -379 605 -377
rect 611 -373 612 -371
rect 611 -379 612 -377
rect 618 -373 619 -371
rect 618 -379 619 -377
rect 625 -373 626 -371
rect 628 -373 629 -371
rect 625 -379 626 -377
rect 632 -373 633 -371
rect 632 -379 633 -377
rect 635 -379 636 -377
rect 639 -373 640 -371
rect 639 -379 640 -377
rect 646 -373 647 -371
rect 649 -379 650 -377
rect 653 -373 654 -371
rect 653 -379 654 -377
rect 660 -373 661 -371
rect 660 -379 661 -377
rect 667 -373 668 -371
rect 667 -379 668 -377
rect 674 -373 675 -371
rect 674 -379 675 -377
rect 681 -373 682 -371
rect 681 -379 682 -377
rect 688 -373 689 -371
rect 688 -379 689 -377
rect 695 -373 696 -371
rect 695 -379 696 -377
rect 702 -373 703 -371
rect 702 -379 703 -377
rect 709 -373 710 -371
rect 709 -379 710 -377
rect 716 -373 717 -371
rect 716 -379 717 -377
rect 723 -373 724 -371
rect 723 -379 724 -377
rect 730 -373 731 -371
rect 730 -379 731 -377
rect 737 -373 738 -371
rect 737 -379 738 -377
rect 747 -373 748 -371
rect 744 -379 745 -377
rect 747 -379 748 -377
rect 751 -373 752 -371
rect 751 -379 752 -377
rect 761 -373 762 -371
rect 758 -379 759 -377
rect 761 -379 762 -377
rect 765 -373 766 -371
rect 765 -379 766 -377
rect 772 -373 773 -371
rect 772 -379 773 -377
rect 775 -379 776 -377
rect 779 -373 780 -371
rect 779 -379 780 -377
rect 786 -373 787 -371
rect 786 -379 787 -377
rect 793 -373 794 -371
rect 796 -373 797 -371
rect 793 -379 794 -377
rect 796 -379 797 -377
rect 800 -373 801 -371
rect 803 -379 804 -377
rect 810 -373 811 -371
rect 807 -379 808 -377
rect 810 -379 811 -377
rect 814 -373 815 -371
rect 814 -379 815 -377
rect 821 -373 822 -371
rect 821 -379 822 -377
rect 828 -373 829 -371
rect 828 -379 829 -377
rect 835 -373 836 -371
rect 838 -373 839 -371
rect 835 -379 836 -377
rect 842 -373 843 -371
rect 845 -373 846 -371
rect 842 -379 843 -377
rect 845 -379 846 -377
rect 849 -373 850 -371
rect 849 -379 850 -377
rect 856 -373 857 -371
rect 856 -379 857 -377
rect 863 -373 864 -371
rect 863 -379 864 -377
rect 870 -373 871 -371
rect 870 -379 871 -377
rect 877 -373 878 -371
rect 880 -373 881 -371
rect 877 -379 878 -377
rect 884 -373 885 -371
rect 884 -379 885 -377
rect 891 -373 892 -371
rect 894 -373 895 -371
rect 891 -379 892 -377
rect 898 -373 899 -371
rect 898 -379 899 -377
rect 905 -373 906 -371
rect 905 -379 906 -377
rect 912 -373 913 -371
rect 912 -379 913 -377
rect 919 -373 920 -371
rect 919 -379 920 -377
rect 926 -373 927 -371
rect 926 -379 927 -377
rect 933 -373 934 -371
rect 933 -379 934 -377
rect 940 -373 941 -371
rect 940 -379 941 -377
rect 947 -373 948 -371
rect 947 -379 948 -377
rect 954 -373 955 -371
rect 954 -379 955 -377
rect 961 -373 962 -371
rect 961 -379 962 -377
rect 968 -373 969 -371
rect 968 -379 969 -377
rect 975 -379 976 -377
rect 978 -379 979 -377
rect 982 -373 983 -371
rect 982 -379 983 -377
rect 989 -373 990 -371
rect 989 -379 990 -377
rect 992 -379 993 -377
rect 996 -373 997 -371
rect 996 -379 997 -377
rect 1003 -373 1004 -371
rect 1003 -379 1004 -377
rect 1010 -373 1011 -371
rect 1010 -379 1011 -377
rect 1017 -373 1018 -371
rect 1020 -373 1021 -371
rect 1017 -379 1018 -377
rect 1020 -379 1021 -377
rect 1024 -373 1025 -371
rect 1027 -373 1028 -371
rect 1027 -379 1028 -377
rect 1031 -373 1032 -371
rect 1031 -379 1032 -377
rect 1038 -373 1039 -371
rect 1038 -379 1039 -377
rect 1045 -373 1046 -371
rect 1045 -379 1046 -377
rect 1052 -373 1053 -371
rect 1052 -379 1053 -377
rect 1059 -373 1060 -371
rect 1059 -379 1060 -377
rect 1066 -373 1067 -371
rect 1066 -379 1067 -377
rect 1073 -373 1074 -371
rect 1076 -373 1077 -371
rect 1073 -379 1074 -377
rect 1076 -379 1077 -377
rect 1083 -373 1084 -371
rect 1080 -379 1081 -377
rect 1083 -379 1084 -377
rect 1087 -373 1088 -371
rect 1087 -379 1088 -377
rect 1094 -373 1095 -371
rect 1094 -379 1095 -377
rect 1104 -373 1105 -371
rect 1101 -379 1102 -377
rect 1104 -379 1105 -377
rect 1108 -373 1109 -371
rect 1108 -379 1109 -377
rect 1115 -373 1116 -371
rect 1115 -379 1116 -377
rect 1122 -373 1123 -371
rect 1122 -379 1123 -377
rect 1129 -373 1130 -371
rect 1129 -379 1130 -377
rect 1136 -373 1137 -371
rect 1136 -379 1137 -377
rect 1143 -373 1144 -371
rect 1143 -379 1144 -377
rect 1150 -373 1151 -371
rect 1150 -379 1151 -377
rect 1157 -373 1158 -371
rect 1157 -379 1158 -377
rect 1164 -373 1165 -371
rect 1164 -379 1165 -377
rect 1171 -373 1172 -371
rect 1171 -379 1172 -377
rect 1181 -373 1182 -371
rect 1178 -379 1179 -377
rect 1181 -379 1182 -377
rect 1185 -373 1186 -371
rect 1185 -379 1186 -377
rect 1192 -373 1193 -371
rect 1192 -379 1193 -377
rect 1199 -373 1200 -371
rect 1199 -379 1200 -377
rect 1206 -373 1207 -371
rect 1206 -379 1207 -377
rect 1213 -373 1214 -371
rect 1213 -379 1214 -377
rect 1220 -373 1221 -371
rect 1220 -379 1221 -377
rect 1227 -373 1228 -371
rect 1227 -379 1228 -377
rect 1234 -373 1235 -371
rect 1234 -379 1235 -377
rect 1241 -373 1242 -371
rect 1241 -379 1242 -377
rect 1248 -373 1249 -371
rect 1248 -379 1249 -377
rect 1255 -373 1256 -371
rect 1255 -379 1256 -377
rect 1262 -373 1263 -371
rect 1262 -379 1263 -377
rect 1269 -373 1270 -371
rect 1269 -379 1270 -377
rect 1276 -373 1277 -371
rect 1276 -379 1277 -377
rect 1283 -373 1284 -371
rect 1283 -379 1284 -377
rect 1290 -373 1291 -371
rect 1290 -379 1291 -377
rect 1297 -373 1298 -371
rect 1297 -379 1298 -377
rect 1304 -373 1305 -371
rect 1304 -379 1305 -377
rect 1311 -373 1312 -371
rect 1311 -379 1312 -377
rect 1318 -373 1319 -371
rect 1318 -379 1319 -377
rect 1325 -373 1326 -371
rect 1328 -373 1329 -371
rect 1328 -379 1329 -377
rect 1332 -373 1333 -371
rect 1332 -379 1333 -377
rect 1339 -373 1340 -371
rect 1339 -379 1340 -377
rect 1346 -373 1347 -371
rect 1346 -379 1347 -377
rect 1353 -379 1354 -377
rect 1356 -379 1357 -377
rect 1360 -373 1361 -371
rect 1360 -379 1361 -377
rect 1367 -373 1368 -371
rect 1367 -379 1368 -377
rect 1374 -373 1375 -371
rect 1374 -379 1375 -377
rect 1381 -373 1382 -371
rect 1381 -379 1382 -377
rect 1388 -373 1389 -371
rect 1388 -379 1389 -377
rect 1395 -373 1396 -371
rect 1395 -379 1396 -377
rect 1402 -373 1403 -371
rect 1402 -379 1403 -377
rect 1409 -373 1410 -371
rect 1409 -379 1410 -377
rect 1416 -373 1417 -371
rect 1416 -379 1417 -377
rect 1423 -373 1424 -371
rect 1423 -379 1424 -377
rect 1430 -373 1431 -371
rect 1430 -379 1431 -377
rect 1437 -373 1438 -371
rect 1437 -379 1438 -377
rect 1444 -373 1445 -371
rect 1444 -379 1445 -377
rect 1451 -373 1452 -371
rect 1451 -379 1452 -377
rect 1458 -373 1459 -371
rect 1458 -379 1459 -377
rect 1465 -373 1466 -371
rect 1465 -379 1466 -377
rect 1472 -373 1473 -371
rect 1472 -379 1473 -377
rect 1479 -373 1480 -371
rect 1479 -379 1480 -377
rect 1486 -373 1487 -371
rect 1486 -379 1487 -377
rect 1493 -373 1494 -371
rect 1493 -379 1494 -377
rect 1500 -373 1501 -371
rect 1500 -379 1501 -377
rect 1507 -373 1508 -371
rect 1507 -379 1508 -377
rect 1514 -373 1515 -371
rect 1514 -379 1515 -377
rect 1521 -373 1522 -371
rect 1521 -379 1522 -377
rect 1528 -373 1529 -371
rect 1528 -379 1529 -377
rect 1535 -373 1536 -371
rect 1535 -379 1536 -377
rect 1542 -373 1543 -371
rect 1542 -379 1543 -377
rect 1549 -373 1550 -371
rect 1549 -379 1550 -377
rect 1556 -373 1557 -371
rect 1556 -379 1557 -377
rect 1563 -373 1564 -371
rect 1563 -379 1564 -377
rect 1570 -373 1571 -371
rect 1570 -379 1571 -377
rect 1577 -373 1578 -371
rect 1577 -379 1578 -377
rect 1584 -373 1585 -371
rect 1584 -379 1585 -377
rect 1591 -373 1592 -371
rect 1591 -379 1592 -377
rect 1598 -373 1599 -371
rect 1598 -379 1599 -377
rect 1605 -373 1606 -371
rect 1605 -379 1606 -377
rect 1612 -373 1613 -371
rect 1615 -373 1616 -371
rect 1612 -379 1613 -377
rect 1619 -373 1620 -371
rect 1619 -379 1620 -377
rect 1626 -373 1627 -371
rect 1626 -379 1627 -377
rect 1633 -373 1634 -371
rect 1633 -379 1634 -377
rect 1640 -373 1641 -371
rect 1640 -379 1641 -377
rect 1647 -373 1648 -371
rect 1647 -379 1648 -377
rect 1654 -373 1655 -371
rect 1654 -379 1655 -377
rect 1661 -373 1662 -371
rect 1661 -379 1662 -377
rect 1668 -373 1669 -371
rect 1668 -379 1669 -377
rect 1675 -373 1676 -371
rect 1675 -379 1676 -377
rect 1682 -373 1683 -371
rect 1682 -379 1683 -377
rect 1689 -373 1690 -371
rect 1689 -379 1690 -377
rect 1696 -373 1697 -371
rect 1696 -379 1697 -377
rect 1703 -373 1704 -371
rect 1703 -379 1704 -377
rect 1710 -373 1711 -371
rect 1710 -379 1711 -377
rect 1717 -373 1718 -371
rect 1717 -379 1718 -377
rect 1724 -373 1725 -371
rect 1724 -379 1725 -377
rect 1731 -373 1732 -371
rect 1731 -379 1732 -377
rect 1738 -373 1739 -371
rect 1738 -379 1739 -377
rect 1745 -373 1746 -371
rect 1745 -379 1746 -377
rect 1752 -373 1753 -371
rect 1752 -379 1753 -377
rect 1759 -373 1760 -371
rect 1759 -379 1760 -377
rect 1766 -373 1767 -371
rect 1766 -379 1767 -377
rect 1773 -373 1774 -371
rect 1773 -379 1774 -377
rect 1780 -373 1781 -371
rect 1780 -379 1781 -377
rect 1787 -373 1788 -371
rect 1787 -379 1788 -377
rect 1794 -373 1795 -371
rect 1794 -379 1795 -377
rect 1801 -373 1802 -371
rect 1801 -379 1802 -377
rect 1808 -373 1809 -371
rect 1808 -379 1809 -377
rect 1815 -373 1816 -371
rect 1815 -379 1816 -377
rect 1822 -373 1823 -371
rect 1822 -379 1823 -377
rect 1829 -373 1830 -371
rect 1829 -379 1830 -377
rect 1836 -373 1837 -371
rect 1836 -379 1837 -377
rect 1843 -373 1844 -371
rect 1843 -379 1844 -377
rect 1927 -373 1928 -371
rect 1927 -379 1928 -377
rect 1962 -373 1963 -371
rect 1962 -379 1963 -377
rect 1969 -373 1970 -371
rect 1969 -379 1970 -377
rect 1983 -373 1984 -371
rect 1983 -379 1984 -377
rect 2004 -373 2005 -371
rect 2004 -379 2005 -377
rect 2193 -373 2194 -371
rect 2193 -379 2194 -377
rect 2 -502 3 -500
rect 2 -508 3 -506
rect 9 -508 10 -506
rect 16 -502 17 -500
rect 16 -508 17 -506
rect 23 -502 24 -500
rect 23 -508 24 -506
rect 44 -502 45 -500
rect 44 -508 45 -506
rect 51 -502 52 -500
rect 51 -508 52 -506
rect 61 -502 62 -500
rect 61 -508 62 -506
rect 65 -502 66 -500
rect 65 -508 66 -506
rect 72 -502 73 -500
rect 72 -508 73 -506
rect 79 -502 80 -500
rect 79 -508 80 -506
rect 86 -502 87 -500
rect 86 -508 87 -506
rect 93 -502 94 -500
rect 93 -508 94 -506
rect 100 -502 101 -500
rect 100 -508 101 -506
rect 107 -502 108 -500
rect 107 -508 108 -506
rect 114 -508 115 -506
rect 117 -508 118 -506
rect 121 -502 122 -500
rect 121 -508 122 -506
rect 128 -502 129 -500
rect 128 -508 129 -506
rect 135 -502 136 -500
rect 135 -508 136 -506
rect 142 -502 143 -500
rect 142 -508 143 -506
rect 149 -502 150 -500
rect 149 -508 150 -506
rect 156 -502 157 -500
rect 156 -508 157 -506
rect 163 -502 164 -500
rect 166 -502 167 -500
rect 166 -508 167 -506
rect 173 -502 174 -500
rect 170 -508 171 -506
rect 173 -508 174 -506
rect 177 -502 178 -500
rect 177 -508 178 -506
rect 184 -502 185 -500
rect 184 -508 185 -506
rect 191 -502 192 -500
rect 191 -508 192 -506
rect 198 -502 199 -500
rect 198 -508 199 -506
rect 205 -502 206 -500
rect 205 -508 206 -506
rect 212 -502 213 -500
rect 215 -502 216 -500
rect 215 -508 216 -506
rect 219 -502 220 -500
rect 222 -502 223 -500
rect 219 -508 220 -506
rect 222 -508 223 -506
rect 226 -502 227 -500
rect 226 -508 227 -506
rect 233 -502 234 -500
rect 233 -508 234 -506
rect 236 -508 237 -506
rect 240 -502 241 -500
rect 240 -508 241 -506
rect 247 -502 248 -500
rect 247 -508 248 -506
rect 254 -502 255 -500
rect 254 -508 255 -506
rect 261 -502 262 -500
rect 261 -508 262 -506
rect 268 -502 269 -500
rect 268 -508 269 -506
rect 275 -502 276 -500
rect 275 -508 276 -506
rect 282 -502 283 -500
rect 282 -508 283 -506
rect 289 -502 290 -500
rect 289 -508 290 -506
rect 296 -502 297 -500
rect 296 -508 297 -506
rect 303 -502 304 -500
rect 303 -508 304 -506
rect 310 -502 311 -500
rect 310 -508 311 -506
rect 317 -502 318 -500
rect 317 -508 318 -506
rect 324 -502 325 -500
rect 324 -508 325 -506
rect 331 -502 332 -500
rect 331 -508 332 -506
rect 338 -502 339 -500
rect 338 -508 339 -506
rect 345 -502 346 -500
rect 345 -508 346 -506
rect 352 -502 353 -500
rect 352 -508 353 -506
rect 359 -502 360 -500
rect 359 -508 360 -506
rect 366 -502 367 -500
rect 366 -508 367 -506
rect 373 -502 374 -500
rect 373 -508 374 -506
rect 380 -502 381 -500
rect 380 -508 381 -506
rect 387 -502 388 -500
rect 387 -508 388 -506
rect 394 -502 395 -500
rect 394 -508 395 -506
rect 401 -502 402 -500
rect 401 -508 402 -506
rect 408 -502 409 -500
rect 408 -508 409 -506
rect 415 -502 416 -500
rect 415 -508 416 -506
rect 422 -502 423 -500
rect 422 -508 423 -506
rect 429 -502 430 -500
rect 429 -508 430 -506
rect 436 -502 437 -500
rect 436 -508 437 -506
rect 443 -502 444 -500
rect 443 -508 444 -506
rect 450 -502 451 -500
rect 450 -508 451 -506
rect 457 -502 458 -500
rect 457 -508 458 -506
rect 464 -502 465 -500
rect 464 -508 465 -506
rect 471 -502 472 -500
rect 471 -508 472 -506
rect 478 -502 479 -500
rect 478 -508 479 -506
rect 485 -502 486 -500
rect 485 -508 486 -506
rect 492 -502 493 -500
rect 495 -502 496 -500
rect 492 -508 493 -506
rect 495 -508 496 -506
rect 499 -502 500 -500
rect 499 -508 500 -506
rect 506 -502 507 -500
rect 506 -508 507 -506
rect 513 -502 514 -500
rect 513 -508 514 -506
rect 520 -502 521 -500
rect 520 -508 521 -506
rect 527 -502 528 -500
rect 527 -508 528 -506
rect 534 -502 535 -500
rect 534 -508 535 -506
rect 537 -508 538 -506
rect 541 -502 542 -500
rect 541 -508 542 -506
rect 548 -502 549 -500
rect 548 -508 549 -506
rect 555 -502 556 -500
rect 555 -508 556 -506
rect 562 -502 563 -500
rect 562 -508 563 -506
rect 569 -502 570 -500
rect 569 -508 570 -506
rect 576 -502 577 -500
rect 576 -508 577 -506
rect 583 -502 584 -500
rect 583 -508 584 -506
rect 590 -502 591 -500
rect 590 -508 591 -506
rect 597 -502 598 -500
rect 600 -502 601 -500
rect 600 -508 601 -506
rect 604 -502 605 -500
rect 604 -508 605 -506
rect 611 -502 612 -500
rect 611 -508 612 -506
rect 618 -502 619 -500
rect 621 -502 622 -500
rect 618 -508 619 -506
rect 621 -508 622 -506
rect 625 -502 626 -500
rect 625 -508 626 -506
rect 632 -502 633 -500
rect 635 -508 636 -506
rect 639 -502 640 -500
rect 639 -508 640 -506
rect 646 -502 647 -500
rect 646 -508 647 -506
rect 653 -502 654 -500
rect 653 -508 654 -506
rect 656 -508 657 -506
rect 660 -502 661 -500
rect 660 -508 661 -506
rect 667 -502 668 -500
rect 667 -508 668 -506
rect 674 -502 675 -500
rect 674 -508 675 -506
rect 681 -502 682 -500
rect 681 -508 682 -506
rect 688 -502 689 -500
rect 688 -508 689 -506
rect 695 -502 696 -500
rect 695 -508 696 -506
rect 702 -502 703 -500
rect 702 -508 703 -506
rect 709 -502 710 -500
rect 709 -508 710 -506
rect 716 -502 717 -500
rect 719 -502 720 -500
rect 716 -508 717 -506
rect 723 -502 724 -500
rect 726 -502 727 -500
rect 723 -508 724 -506
rect 726 -508 727 -506
rect 730 -502 731 -500
rect 730 -508 731 -506
rect 737 -502 738 -500
rect 740 -502 741 -500
rect 737 -508 738 -506
rect 740 -508 741 -506
rect 744 -502 745 -500
rect 744 -508 745 -506
rect 751 -502 752 -500
rect 751 -508 752 -506
rect 758 -502 759 -500
rect 758 -508 759 -506
rect 765 -502 766 -500
rect 765 -508 766 -506
rect 772 -502 773 -500
rect 772 -508 773 -506
rect 779 -502 780 -500
rect 779 -508 780 -506
rect 786 -502 787 -500
rect 786 -508 787 -506
rect 793 -502 794 -500
rect 793 -508 794 -506
rect 800 -502 801 -500
rect 800 -508 801 -506
rect 807 -502 808 -500
rect 807 -508 808 -506
rect 814 -502 815 -500
rect 814 -508 815 -506
rect 821 -502 822 -500
rect 821 -508 822 -506
rect 828 -502 829 -500
rect 828 -508 829 -506
rect 835 -502 836 -500
rect 835 -508 836 -506
rect 842 -502 843 -500
rect 842 -508 843 -506
rect 849 -502 850 -500
rect 852 -502 853 -500
rect 849 -508 850 -506
rect 856 -502 857 -500
rect 856 -508 857 -506
rect 863 -502 864 -500
rect 863 -508 864 -506
rect 870 -502 871 -500
rect 870 -508 871 -506
rect 877 -502 878 -500
rect 877 -508 878 -506
rect 887 -502 888 -500
rect 887 -508 888 -506
rect 891 -502 892 -500
rect 891 -508 892 -506
rect 898 -502 899 -500
rect 898 -508 899 -506
rect 905 -502 906 -500
rect 905 -508 906 -506
rect 912 -502 913 -500
rect 912 -508 913 -506
rect 915 -508 916 -506
rect 919 -502 920 -500
rect 919 -508 920 -506
rect 926 -502 927 -500
rect 926 -508 927 -506
rect 933 -502 934 -500
rect 933 -508 934 -506
rect 936 -508 937 -506
rect 940 -502 941 -500
rect 940 -508 941 -506
rect 947 -502 948 -500
rect 947 -508 948 -506
rect 954 -502 955 -500
rect 957 -502 958 -500
rect 954 -508 955 -506
rect 961 -502 962 -500
rect 961 -508 962 -506
rect 968 -502 969 -500
rect 971 -502 972 -500
rect 968 -508 969 -506
rect 971 -508 972 -506
rect 978 -502 979 -500
rect 975 -508 976 -506
rect 978 -508 979 -506
rect 982 -502 983 -500
rect 985 -502 986 -500
rect 982 -508 983 -506
rect 985 -508 986 -506
rect 989 -502 990 -500
rect 989 -508 990 -506
rect 992 -508 993 -506
rect 996 -502 997 -500
rect 996 -508 997 -506
rect 1006 -502 1007 -500
rect 1003 -508 1004 -506
rect 1006 -508 1007 -506
rect 1010 -502 1011 -500
rect 1010 -508 1011 -506
rect 1017 -502 1018 -500
rect 1017 -508 1018 -506
rect 1024 -502 1025 -500
rect 1027 -502 1028 -500
rect 1031 -502 1032 -500
rect 1031 -508 1032 -506
rect 1038 -502 1039 -500
rect 1038 -508 1039 -506
rect 1045 -502 1046 -500
rect 1045 -508 1046 -506
rect 1052 -502 1053 -500
rect 1052 -508 1053 -506
rect 1059 -502 1060 -500
rect 1059 -508 1060 -506
rect 1066 -502 1067 -500
rect 1066 -508 1067 -506
rect 1073 -502 1074 -500
rect 1073 -508 1074 -506
rect 1080 -502 1081 -500
rect 1083 -502 1084 -500
rect 1080 -508 1081 -506
rect 1083 -508 1084 -506
rect 1087 -502 1088 -500
rect 1087 -508 1088 -506
rect 1094 -502 1095 -500
rect 1094 -508 1095 -506
rect 1101 -502 1102 -500
rect 1101 -508 1102 -506
rect 1108 -502 1109 -500
rect 1108 -508 1109 -506
rect 1115 -502 1116 -500
rect 1115 -508 1116 -506
rect 1122 -502 1123 -500
rect 1125 -502 1126 -500
rect 1125 -508 1126 -506
rect 1129 -502 1130 -500
rect 1129 -508 1130 -506
rect 1136 -502 1137 -500
rect 1136 -508 1137 -506
rect 1143 -502 1144 -500
rect 1143 -508 1144 -506
rect 1150 -502 1151 -500
rect 1150 -508 1151 -506
rect 1157 -502 1158 -500
rect 1157 -508 1158 -506
rect 1167 -502 1168 -500
rect 1164 -508 1165 -506
rect 1167 -508 1168 -506
rect 1171 -502 1172 -500
rect 1171 -508 1172 -506
rect 1178 -502 1179 -500
rect 1178 -508 1179 -506
rect 1185 -502 1186 -500
rect 1185 -508 1186 -506
rect 1192 -502 1193 -500
rect 1192 -508 1193 -506
rect 1199 -502 1200 -500
rect 1199 -508 1200 -506
rect 1206 -502 1207 -500
rect 1206 -508 1207 -506
rect 1213 -502 1214 -500
rect 1213 -508 1214 -506
rect 1220 -502 1221 -500
rect 1220 -508 1221 -506
rect 1227 -502 1228 -500
rect 1227 -508 1228 -506
rect 1234 -502 1235 -500
rect 1234 -508 1235 -506
rect 1241 -502 1242 -500
rect 1241 -508 1242 -506
rect 1248 -502 1249 -500
rect 1248 -508 1249 -506
rect 1255 -502 1256 -500
rect 1255 -508 1256 -506
rect 1262 -502 1263 -500
rect 1262 -508 1263 -506
rect 1269 -502 1270 -500
rect 1269 -508 1270 -506
rect 1276 -502 1277 -500
rect 1276 -508 1277 -506
rect 1283 -502 1284 -500
rect 1283 -508 1284 -506
rect 1290 -502 1291 -500
rect 1290 -508 1291 -506
rect 1297 -502 1298 -500
rect 1297 -508 1298 -506
rect 1304 -502 1305 -500
rect 1304 -508 1305 -506
rect 1311 -502 1312 -500
rect 1311 -508 1312 -506
rect 1318 -502 1319 -500
rect 1318 -508 1319 -506
rect 1325 -502 1326 -500
rect 1325 -508 1326 -506
rect 1332 -502 1333 -500
rect 1332 -508 1333 -506
rect 1339 -502 1340 -500
rect 1339 -508 1340 -506
rect 1346 -502 1347 -500
rect 1346 -508 1347 -506
rect 1353 -502 1354 -500
rect 1353 -508 1354 -506
rect 1360 -502 1361 -500
rect 1360 -508 1361 -506
rect 1367 -502 1368 -500
rect 1367 -508 1368 -506
rect 1374 -502 1375 -500
rect 1374 -508 1375 -506
rect 1381 -502 1382 -500
rect 1381 -508 1382 -506
rect 1388 -502 1389 -500
rect 1388 -508 1389 -506
rect 1395 -502 1396 -500
rect 1395 -508 1396 -506
rect 1402 -502 1403 -500
rect 1402 -508 1403 -506
rect 1409 -502 1410 -500
rect 1409 -508 1410 -506
rect 1416 -502 1417 -500
rect 1416 -508 1417 -506
rect 1423 -502 1424 -500
rect 1423 -508 1424 -506
rect 1430 -502 1431 -500
rect 1430 -508 1431 -506
rect 1440 -502 1441 -500
rect 1437 -508 1438 -506
rect 1440 -508 1441 -506
rect 1444 -502 1445 -500
rect 1444 -508 1445 -506
rect 1451 -502 1452 -500
rect 1451 -508 1452 -506
rect 1458 -502 1459 -500
rect 1458 -508 1459 -506
rect 1465 -502 1466 -500
rect 1465 -508 1466 -506
rect 1472 -502 1473 -500
rect 1472 -508 1473 -506
rect 1479 -502 1480 -500
rect 1479 -508 1480 -506
rect 1486 -502 1487 -500
rect 1486 -508 1487 -506
rect 1493 -502 1494 -500
rect 1493 -508 1494 -506
rect 1500 -502 1501 -500
rect 1500 -508 1501 -506
rect 1507 -502 1508 -500
rect 1507 -508 1508 -506
rect 1514 -502 1515 -500
rect 1514 -508 1515 -506
rect 1521 -502 1522 -500
rect 1521 -508 1522 -506
rect 1528 -502 1529 -500
rect 1528 -508 1529 -506
rect 1535 -502 1536 -500
rect 1535 -508 1536 -506
rect 1542 -502 1543 -500
rect 1542 -508 1543 -506
rect 1549 -502 1550 -500
rect 1549 -508 1550 -506
rect 1556 -502 1557 -500
rect 1556 -508 1557 -506
rect 1563 -502 1564 -500
rect 1563 -508 1564 -506
rect 1570 -502 1571 -500
rect 1570 -508 1571 -506
rect 1577 -502 1578 -500
rect 1577 -508 1578 -506
rect 1584 -502 1585 -500
rect 1584 -508 1585 -506
rect 1591 -502 1592 -500
rect 1591 -508 1592 -506
rect 1598 -502 1599 -500
rect 1598 -508 1599 -506
rect 1605 -502 1606 -500
rect 1605 -508 1606 -506
rect 1612 -502 1613 -500
rect 1612 -508 1613 -506
rect 1619 -502 1620 -500
rect 1619 -508 1620 -506
rect 1626 -502 1627 -500
rect 1626 -508 1627 -506
rect 1633 -502 1634 -500
rect 1633 -508 1634 -506
rect 1640 -502 1641 -500
rect 1640 -508 1641 -506
rect 1647 -502 1648 -500
rect 1647 -508 1648 -506
rect 1654 -502 1655 -500
rect 1654 -508 1655 -506
rect 1661 -502 1662 -500
rect 1661 -508 1662 -506
rect 1668 -502 1669 -500
rect 1668 -508 1669 -506
rect 1675 -502 1676 -500
rect 1675 -508 1676 -506
rect 1682 -502 1683 -500
rect 1682 -508 1683 -506
rect 1689 -502 1690 -500
rect 1689 -508 1690 -506
rect 1696 -502 1697 -500
rect 1696 -508 1697 -506
rect 1703 -502 1704 -500
rect 1703 -508 1704 -506
rect 1710 -502 1711 -500
rect 1710 -508 1711 -506
rect 1717 -502 1718 -500
rect 1717 -508 1718 -506
rect 1724 -502 1725 -500
rect 1724 -508 1725 -506
rect 1731 -502 1732 -500
rect 1731 -508 1732 -506
rect 1738 -502 1739 -500
rect 1738 -508 1739 -506
rect 1745 -502 1746 -500
rect 1745 -508 1746 -506
rect 1752 -502 1753 -500
rect 1752 -508 1753 -506
rect 1759 -502 1760 -500
rect 1759 -508 1760 -506
rect 1766 -502 1767 -500
rect 1766 -508 1767 -506
rect 1773 -502 1774 -500
rect 1773 -508 1774 -506
rect 1780 -502 1781 -500
rect 1780 -508 1781 -506
rect 1787 -502 1788 -500
rect 1787 -508 1788 -506
rect 1794 -502 1795 -500
rect 1794 -508 1795 -506
rect 1801 -502 1802 -500
rect 1801 -508 1802 -506
rect 1808 -502 1809 -500
rect 1808 -508 1809 -506
rect 1815 -502 1816 -500
rect 1815 -508 1816 -506
rect 1822 -502 1823 -500
rect 1822 -508 1823 -506
rect 1829 -502 1830 -500
rect 1829 -508 1830 -506
rect 1836 -502 1837 -500
rect 1836 -508 1837 -506
rect 1843 -502 1844 -500
rect 1843 -508 1844 -506
rect 1850 -502 1851 -500
rect 1850 -508 1851 -506
rect 1857 -502 1858 -500
rect 1857 -508 1858 -506
rect 1864 -502 1865 -500
rect 1864 -508 1865 -506
rect 1871 -502 1872 -500
rect 1871 -508 1872 -506
rect 1878 -502 1879 -500
rect 1878 -508 1879 -506
rect 1885 -502 1886 -500
rect 1885 -508 1886 -506
rect 1892 -502 1893 -500
rect 1892 -508 1893 -506
rect 1899 -502 1900 -500
rect 1899 -508 1900 -506
rect 1906 -502 1907 -500
rect 1906 -508 1907 -506
rect 1913 -502 1914 -500
rect 1913 -508 1914 -506
rect 1920 -502 1921 -500
rect 1920 -508 1921 -506
rect 1927 -502 1928 -500
rect 1927 -508 1928 -506
rect 1934 -502 1935 -500
rect 1934 -508 1935 -506
rect 1941 -502 1942 -500
rect 1941 -508 1942 -506
rect 1948 -502 1949 -500
rect 1948 -508 1949 -506
rect 1955 -502 1956 -500
rect 1958 -502 1959 -500
rect 1955 -508 1956 -506
rect 1958 -508 1959 -506
rect 1962 -502 1963 -500
rect 1962 -508 1963 -506
rect 1969 -502 1970 -500
rect 1969 -508 1970 -506
rect 1976 -502 1977 -500
rect 1976 -508 1977 -506
rect 1979 -508 1980 -506
rect 1983 -502 1984 -500
rect 1983 -508 1984 -506
rect 1990 -502 1991 -500
rect 1990 -508 1991 -506
rect 1997 -502 1998 -500
rect 1997 -508 1998 -506
rect 2007 -508 2008 -506
rect 2011 -502 2012 -500
rect 2011 -508 2012 -506
rect 2014 -508 2015 -506
rect 2018 -508 2019 -506
rect 2021 -508 2022 -506
rect 2039 -502 2040 -500
rect 2039 -508 2040 -506
rect 2088 -502 2089 -500
rect 2088 -508 2089 -506
rect 2116 -502 2117 -500
rect 2116 -508 2117 -506
rect 2144 -502 2145 -500
rect 2144 -508 2145 -506
rect 2263 -502 2264 -500
rect 2263 -508 2264 -506
rect 2284 -502 2285 -500
rect 2284 -508 2285 -506
rect 5 -641 6 -639
rect 9 -635 10 -633
rect 9 -641 10 -639
rect 16 -635 17 -633
rect 16 -641 17 -639
rect 23 -635 24 -633
rect 23 -641 24 -639
rect 30 -635 31 -633
rect 30 -641 31 -639
rect 37 -635 38 -633
rect 37 -641 38 -639
rect 44 -635 45 -633
rect 44 -641 45 -639
rect 51 -635 52 -633
rect 51 -641 52 -639
rect 58 -635 59 -633
rect 61 -635 62 -633
rect 58 -641 59 -639
rect 65 -635 66 -633
rect 65 -641 66 -639
rect 72 -635 73 -633
rect 75 -635 76 -633
rect 72 -641 73 -639
rect 75 -641 76 -639
rect 79 -635 80 -633
rect 79 -641 80 -639
rect 86 -635 87 -633
rect 86 -641 87 -639
rect 93 -635 94 -633
rect 93 -641 94 -639
rect 100 -635 101 -633
rect 103 -635 104 -633
rect 100 -641 101 -639
rect 107 -635 108 -633
rect 107 -641 108 -639
rect 114 -635 115 -633
rect 114 -641 115 -639
rect 121 -635 122 -633
rect 121 -641 122 -639
rect 128 -635 129 -633
rect 128 -641 129 -639
rect 135 -635 136 -633
rect 138 -635 139 -633
rect 135 -641 136 -639
rect 142 -635 143 -633
rect 142 -641 143 -639
rect 149 -635 150 -633
rect 149 -641 150 -639
rect 156 -635 157 -633
rect 156 -641 157 -639
rect 163 -635 164 -633
rect 163 -641 164 -639
rect 173 -635 174 -633
rect 173 -641 174 -639
rect 177 -635 178 -633
rect 177 -641 178 -639
rect 184 -635 185 -633
rect 184 -641 185 -639
rect 191 -635 192 -633
rect 191 -641 192 -639
rect 198 -635 199 -633
rect 198 -641 199 -639
rect 205 -635 206 -633
rect 205 -641 206 -639
rect 208 -641 209 -639
rect 212 -635 213 -633
rect 212 -641 213 -639
rect 219 -635 220 -633
rect 219 -641 220 -639
rect 226 -635 227 -633
rect 226 -641 227 -639
rect 233 -635 234 -633
rect 233 -641 234 -639
rect 240 -635 241 -633
rect 240 -641 241 -639
rect 247 -635 248 -633
rect 250 -635 251 -633
rect 250 -641 251 -639
rect 254 -635 255 -633
rect 254 -641 255 -639
rect 261 -635 262 -633
rect 261 -641 262 -639
rect 268 -635 269 -633
rect 268 -641 269 -639
rect 275 -635 276 -633
rect 275 -641 276 -639
rect 282 -635 283 -633
rect 282 -641 283 -639
rect 289 -635 290 -633
rect 289 -641 290 -639
rect 296 -635 297 -633
rect 296 -641 297 -639
rect 303 -635 304 -633
rect 303 -641 304 -639
rect 310 -635 311 -633
rect 310 -641 311 -639
rect 317 -635 318 -633
rect 317 -641 318 -639
rect 324 -635 325 -633
rect 324 -641 325 -639
rect 331 -635 332 -633
rect 331 -641 332 -639
rect 338 -635 339 -633
rect 338 -641 339 -639
rect 345 -635 346 -633
rect 345 -641 346 -639
rect 352 -635 353 -633
rect 352 -641 353 -639
rect 359 -635 360 -633
rect 359 -641 360 -639
rect 366 -635 367 -633
rect 366 -641 367 -639
rect 373 -635 374 -633
rect 373 -641 374 -639
rect 380 -635 381 -633
rect 380 -641 381 -639
rect 387 -635 388 -633
rect 387 -641 388 -639
rect 394 -635 395 -633
rect 394 -641 395 -639
rect 401 -635 402 -633
rect 401 -641 402 -639
rect 408 -635 409 -633
rect 408 -641 409 -639
rect 415 -635 416 -633
rect 415 -641 416 -639
rect 422 -635 423 -633
rect 422 -641 423 -639
rect 429 -635 430 -633
rect 432 -635 433 -633
rect 429 -641 430 -639
rect 432 -641 433 -639
rect 436 -635 437 -633
rect 436 -641 437 -639
rect 443 -635 444 -633
rect 443 -641 444 -639
rect 450 -635 451 -633
rect 450 -641 451 -639
rect 457 -635 458 -633
rect 457 -641 458 -639
rect 464 -635 465 -633
rect 464 -641 465 -639
rect 471 -635 472 -633
rect 471 -641 472 -639
rect 478 -635 479 -633
rect 478 -641 479 -639
rect 485 -635 486 -633
rect 485 -641 486 -639
rect 492 -635 493 -633
rect 492 -641 493 -639
rect 499 -635 500 -633
rect 499 -641 500 -639
rect 506 -635 507 -633
rect 506 -641 507 -639
rect 513 -635 514 -633
rect 513 -641 514 -639
rect 520 -635 521 -633
rect 520 -641 521 -639
rect 527 -635 528 -633
rect 527 -641 528 -639
rect 537 -635 538 -633
rect 534 -641 535 -639
rect 537 -641 538 -639
rect 541 -635 542 -633
rect 541 -641 542 -639
rect 548 -635 549 -633
rect 548 -641 549 -639
rect 555 -635 556 -633
rect 555 -641 556 -639
rect 562 -635 563 -633
rect 565 -635 566 -633
rect 562 -641 563 -639
rect 565 -641 566 -639
rect 569 -635 570 -633
rect 569 -641 570 -639
rect 576 -635 577 -633
rect 576 -641 577 -639
rect 583 -635 584 -633
rect 586 -635 587 -633
rect 583 -641 584 -639
rect 586 -641 587 -639
rect 590 -635 591 -633
rect 593 -635 594 -633
rect 590 -641 591 -639
rect 597 -635 598 -633
rect 597 -641 598 -639
rect 604 -635 605 -633
rect 604 -641 605 -639
rect 611 -635 612 -633
rect 611 -641 612 -639
rect 618 -635 619 -633
rect 618 -641 619 -639
rect 625 -635 626 -633
rect 625 -641 626 -639
rect 632 -635 633 -633
rect 632 -641 633 -639
rect 639 -635 640 -633
rect 639 -641 640 -639
rect 649 -635 650 -633
rect 646 -641 647 -639
rect 649 -641 650 -639
rect 653 -635 654 -633
rect 653 -641 654 -639
rect 660 -635 661 -633
rect 663 -635 664 -633
rect 660 -641 661 -639
rect 663 -641 664 -639
rect 667 -635 668 -633
rect 667 -641 668 -639
rect 674 -635 675 -633
rect 674 -641 675 -639
rect 681 -635 682 -633
rect 681 -641 682 -639
rect 688 -635 689 -633
rect 688 -641 689 -639
rect 695 -635 696 -633
rect 695 -641 696 -639
rect 702 -635 703 -633
rect 702 -641 703 -639
rect 709 -635 710 -633
rect 709 -641 710 -639
rect 716 -635 717 -633
rect 716 -641 717 -639
rect 723 -635 724 -633
rect 723 -641 724 -639
rect 730 -635 731 -633
rect 733 -635 734 -633
rect 730 -641 731 -639
rect 733 -641 734 -639
rect 737 -635 738 -633
rect 737 -641 738 -639
rect 744 -635 745 -633
rect 744 -641 745 -639
rect 747 -641 748 -639
rect 751 -635 752 -633
rect 751 -641 752 -639
rect 758 -635 759 -633
rect 758 -641 759 -639
rect 765 -635 766 -633
rect 765 -641 766 -639
rect 772 -635 773 -633
rect 772 -641 773 -639
rect 779 -635 780 -633
rect 779 -641 780 -639
rect 786 -635 787 -633
rect 789 -641 790 -639
rect 793 -635 794 -633
rect 793 -641 794 -639
rect 800 -635 801 -633
rect 800 -641 801 -639
rect 810 -635 811 -633
rect 807 -641 808 -639
rect 810 -641 811 -639
rect 814 -635 815 -633
rect 814 -641 815 -639
rect 821 -635 822 -633
rect 824 -635 825 -633
rect 821 -641 822 -639
rect 824 -641 825 -639
rect 828 -635 829 -633
rect 828 -641 829 -639
rect 835 -635 836 -633
rect 835 -641 836 -639
rect 842 -635 843 -633
rect 842 -641 843 -639
rect 849 -635 850 -633
rect 852 -635 853 -633
rect 849 -641 850 -639
rect 852 -641 853 -639
rect 856 -635 857 -633
rect 856 -641 857 -639
rect 863 -635 864 -633
rect 863 -641 864 -639
rect 870 -635 871 -633
rect 870 -641 871 -639
rect 877 -635 878 -633
rect 877 -641 878 -639
rect 884 -635 885 -633
rect 884 -641 885 -639
rect 891 -635 892 -633
rect 891 -641 892 -639
rect 898 -635 899 -633
rect 898 -641 899 -639
rect 905 -635 906 -633
rect 905 -641 906 -639
rect 912 -635 913 -633
rect 912 -641 913 -639
rect 919 -635 920 -633
rect 919 -641 920 -639
rect 926 -635 927 -633
rect 929 -635 930 -633
rect 926 -641 927 -639
rect 929 -641 930 -639
rect 933 -635 934 -633
rect 933 -641 934 -639
rect 940 -635 941 -633
rect 940 -641 941 -639
rect 943 -641 944 -639
rect 947 -635 948 -633
rect 947 -641 948 -639
rect 954 -635 955 -633
rect 954 -641 955 -639
rect 961 -635 962 -633
rect 961 -641 962 -639
rect 968 -635 969 -633
rect 968 -641 969 -639
rect 975 -635 976 -633
rect 975 -641 976 -639
rect 985 -635 986 -633
rect 985 -641 986 -639
rect 989 -635 990 -633
rect 989 -641 990 -639
rect 996 -635 997 -633
rect 996 -641 997 -639
rect 1003 -635 1004 -633
rect 1003 -641 1004 -639
rect 1010 -635 1011 -633
rect 1013 -635 1014 -633
rect 1010 -641 1011 -639
rect 1017 -635 1018 -633
rect 1017 -641 1018 -639
rect 1024 -635 1025 -633
rect 1024 -641 1025 -639
rect 1031 -635 1032 -633
rect 1034 -635 1035 -633
rect 1031 -641 1032 -639
rect 1038 -635 1039 -633
rect 1038 -641 1039 -639
rect 1045 -635 1046 -633
rect 1045 -641 1046 -639
rect 1052 -635 1053 -633
rect 1052 -641 1053 -639
rect 1059 -635 1060 -633
rect 1062 -635 1063 -633
rect 1059 -641 1060 -639
rect 1062 -641 1063 -639
rect 1066 -635 1067 -633
rect 1066 -641 1067 -639
rect 1073 -635 1074 -633
rect 1073 -641 1074 -639
rect 1080 -635 1081 -633
rect 1080 -641 1081 -639
rect 1083 -641 1084 -639
rect 1087 -635 1088 -633
rect 1087 -641 1088 -639
rect 1094 -635 1095 -633
rect 1094 -641 1095 -639
rect 1097 -641 1098 -639
rect 1101 -635 1102 -633
rect 1101 -641 1102 -639
rect 1108 -635 1109 -633
rect 1108 -641 1109 -639
rect 1115 -635 1116 -633
rect 1115 -641 1116 -639
rect 1122 -635 1123 -633
rect 1122 -641 1123 -639
rect 1129 -635 1130 -633
rect 1129 -641 1130 -639
rect 1136 -635 1137 -633
rect 1136 -641 1137 -639
rect 1143 -635 1144 -633
rect 1146 -635 1147 -633
rect 1143 -641 1144 -639
rect 1146 -641 1147 -639
rect 1150 -635 1151 -633
rect 1150 -641 1151 -639
rect 1153 -641 1154 -639
rect 1157 -635 1158 -633
rect 1157 -641 1158 -639
rect 1164 -635 1165 -633
rect 1164 -641 1165 -639
rect 1171 -635 1172 -633
rect 1171 -641 1172 -639
rect 1178 -635 1179 -633
rect 1178 -641 1179 -639
rect 1185 -635 1186 -633
rect 1185 -641 1186 -639
rect 1192 -635 1193 -633
rect 1192 -641 1193 -639
rect 1199 -635 1200 -633
rect 1202 -635 1203 -633
rect 1199 -641 1200 -639
rect 1202 -641 1203 -639
rect 1206 -635 1207 -633
rect 1206 -641 1207 -639
rect 1213 -635 1214 -633
rect 1216 -635 1217 -633
rect 1213 -641 1214 -639
rect 1216 -641 1217 -639
rect 1220 -635 1221 -633
rect 1220 -641 1221 -639
rect 1227 -635 1228 -633
rect 1227 -641 1228 -639
rect 1234 -635 1235 -633
rect 1234 -641 1235 -639
rect 1241 -635 1242 -633
rect 1241 -641 1242 -639
rect 1248 -635 1249 -633
rect 1248 -641 1249 -639
rect 1255 -635 1256 -633
rect 1255 -641 1256 -639
rect 1262 -635 1263 -633
rect 1262 -641 1263 -639
rect 1269 -635 1270 -633
rect 1269 -641 1270 -639
rect 1276 -635 1277 -633
rect 1276 -641 1277 -639
rect 1283 -635 1284 -633
rect 1283 -641 1284 -639
rect 1290 -635 1291 -633
rect 1290 -641 1291 -639
rect 1297 -635 1298 -633
rect 1297 -641 1298 -639
rect 1300 -641 1301 -639
rect 1304 -635 1305 -633
rect 1304 -641 1305 -639
rect 1311 -635 1312 -633
rect 1311 -641 1312 -639
rect 1318 -635 1319 -633
rect 1318 -641 1319 -639
rect 1325 -635 1326 -633
rect 1325 -641 1326 -639
rect 1332 -635 1333 -633
rect 1332 -641 1333 -639
rect 1339 -635 1340 -633
rect 1339 -641 1340 -639
rect 1346 -635 1347 -633
rect 1346 -641 1347 -639
rect 1353 -635 1354 -633
rect 1353 -641 1354 -639
rect 1360 -635 1361 -633
rect 1360 -641 1361 -639
rect 1367 -635 1368 -633
rect 1367 -641 1368 -639
rect 1374 -635 1375 -633
rect 1374 -641 1375 -639
rect 1381 -635 1382 -633
rect 1381 -641 1382 -639
rect 1388 -635 1389 -633
rect 1388 -641 1389 -639
rect 1395 -635 1396 -633
rect 1395 -641 1396 -639
rect 1402 -635 1403 -633
rect 1402 -641 1403 -639
rect 1409 -635 1410 -633
rect 1409 -641 1410 -639
rect 1416 -635 1417 -633
rect 1416 -641 1417 -639
rect 1423 -635 1424 -633
rect 1423 -641 1424 -639
rect 1430 -635 1431 -633
rect 1430 -641 1431 -639
rect 1437 -635 1438 -633
rect 1437 -641 1438 -639
rect 1444 -635 1445 -633
rect 1444 -641 1445 -639
rect 1451 -635 1452 -633
rect 1451 -641 1452 -639
rect 1458 -635 1459 -633
rect 1458 -641 1459 -639
rect 1465 -635 1466 -633
rect 1465 -641 1466 -639
rect 1472 -635 1473 -633
rect 1472 -641 1473 -639
rect 1479 -635 1480 -633
rect 1479 -641 1480 -639
rect 1489 -635 1490 -633
rect 1486 -641 1487 -639
rect 1493 -635 1494 -633
rect 1493 -641 1494 -639
rect 1500 -635 1501 -633
rect 1500 -641 1501 -639
rect 1507 -635 1508 -633
rect 1507 -641 1508 -639
rect 1514 -635 1515 -633
rect 1514 -641 1515 -639
rect 1521 -635 1522 -633
rect 1521 -641 1522 -639
rect 1528 -635 1529 -633
rect 1528 -641 1529 -639
rect 1535 -635 1536 -633
rect 1535 -641 1536 -639
rect 1542 -635 1543 -633
rect 1542 -641 1543 -639
rect 1549 -635 1550 -633
rect 1549 -641 1550 -639
rect 1556 -635 1557 -633
rect 1556 -641 1557 -639
rect 1563 -635 1564 -633
rect 1563 -641 1564 -639
rect 1570 -635 1571 -633
rect 1570 -641 1571 -639
rect 1577 -635 1578 -633
rect 1577 -641 1578 -639
rect 1584 -635 1585 -633
rect 1584 -641 1585 -639
rect 1591 -635 1592 -633
rect 1591 -641 1592 -639
rect 1598 -635 1599 -633
rect 1598 -641 1599 -639
rect 1605 -635 1606 -633
rect 1605 -641 1606 -639
rect 1612 -635 1613 -633
rect 1612 -641 1613 -639
rect 1619 -635 1620 -633
rect 1619 -641 1620 -639
rect 1626 -635 1627 -633
rect 1626 -641 1627 -639
rect 1633 -635 1634 -633
rect 1633 -641 1634 -639
rect 1640 -635 1641 -633
rect 1640 -641 1641 -639
rect 1647 -635 1648 -633
rect 1647 -641 1648 -639
rect 1654 -635 1655 -633
rect 1654 -641 1655 -639
rect 1661 -635 1662 -633
rect 1661 -641 1662 -639
rect 1668 -635 1669 -633
rect 1668 -641 1669 -639
rect 1675 -635 1676 -633
rect 1675 -641 1676 -639
rect 1682 -635 1683 -633
rect 1682 -641 1683 -639
rect 1689 -635 1690 -633
rect 1689 -641 1690 -639
rect 1696 -635 1697 -633
rect 1696 -641 1697 -639
rect 1703 -635 1704 -633
rect 1703 -641 1704 -639
rect 1710 -635 1711 -633
rect 1710 -641 1711 -639
rect 1717 -635 1718 -633
rect 1717 -641 1718 -639
rect 1724 -635 1725 -633
rect 1724 -641 1725 -639
rect 1731 -635 1732 -633
rect 1731 -641 1732 -639
rect 1738 -635 1739 -633
rect 1738 -641 1739 -639
rect 1745 -635 1746 -633
rect 1745 -641 1746 -639
rect 1752 -635 1753 -633
rect 1752 -641 1753 -639
rect 1759 -635 1760 -633
rect 1759 -641 1760 -639
rect 1766 -635 1767 -633
rect 1766 -641 1767 -639
rect 1773 -635 1774 -633
rect 1773 -641 1774 -639
rect 1780 -635 1781 -633
rect 1780 -641 1781 -639
rect 1787 -635 1788 -633
rect 1787 -641 1788 -639
rect 1794 -635 1795 -633
rect 1794 -641 1795 -639
rect 1801 -635 1802 -633
rect 1801 -641 1802 -639
rect 1808 -635 1809 -633
rect 1808 -641 1809 -639
rect 1815 -635 1816 -633
rect 1815 -641 1816 -639
rect 1822 -635 1823 -633
rect 1822 -641 1823 -639
rect 1829 -635 1830 -633
rect 1829 -641 1830 -639
rect 1836 -635 1837 -633
rect 1836 -641 1837 -639
rect 1843 -635 1844 -633
rect 1843 -641 1844 -639
rect 1850 -635 1851 -633
rect 1850 -641 1851 -639
rect 1857 -635 1858 -633
rect 1857 -641 1858 -639
rect 1864 -635 1865 -633
rect 1864 -641 1865 -639
rect 1871 -635 1872 -633
rect 1871 -641 1872 -639
rect 1878 -635 1879 -633
rect 1878 -641 1879 -639
rect 1885 -635 1886 -633
rect 1885 -641 1886 -639
rect 1892 -635 1893 -633
rect 1892 -641 1893 -639
rect 1899 -635 1900 -633
rect 1899 -641 1900 -639
rect 1906 -635 1907 -633
rect 1906 -641 1907 -639
rect 1913 -635 1914 -633
rect 1913 -641 1914 -639
rect 1920 -635 1921 -633
rect 1920 -641 1921 -639
rect 1927 -635 1928 -633
rect 1927 -641 1928 -639
rect 1934 -635 1935 -633
rect 1934 -641 1935 -639
rect 1941 -635 1942 -633
rect 1941 -641 1942 -639
rect 1948 -635 1949 -633
rect 1948 -641 1949 -639
rect 1955 -635 1956 -633
rect 1955 -641 1956 -639
rect 1962 -635 1963 -633
rect 1962 -641 1963 -639
rect 1969 -635 1970 -633
rect 1969 -641 1970 -639
rect 1976 -635 1977 -633
rect 1976 -641 1977 -639
rect 1983 -635 1984 -633
rect 1983 -641 1984 -639
rect 1990 -635 1991 -633
rect 1990 -641 1991 -639
rect 1997 -635 1998 -633
rect 1997 -641 1998 -639
rect 2004 -635 2005 -633
rect 2004 -641 2005 -639
rect 2011 -635 2012 -633
rect 2011 -641 2012 -639
rect 2018 -635 2019 -633
rect 2018 -641 2019 -639
rect 2025 -635 2026 -633
rect 2025 -641 2026 -639
rect 2032 -635 2033 -633
rect 2032 -641 2033 -639
rect 2039 -635 2040 -633
rect 2039 -641 2040 -639
rect 2046 -635 2047 -633
rect 2046 -641 2047 -639
rect 2053 -635 2054 -633
rect 2053 -641 2054 -639
rect 2060 -635 2061 -633
rect 2060 -641 2061 -639
rect 2067 -635 2068 -633
rect 2067 -641 2068 -639
rect 2074 -635 2075 -633
rect 2074 -641 2075 -639
rect 2081 -635 2082 -633
rect 2081 -641 2082 -639
rect 2088 -635 2089 -633
rect 2088 -641 2089 -639
rect 2095 -635 2096 -633
rect 2095 -641 2096 -639
rect 2102 -635 2103 -633
rect 2102 -641 2103 -639
rect 2109 -635 2110 -633
rect 2109 -641 2110 -639
rect 2116 -635 2117 -633
rect 2116 -641 2117 -639
rect 2123 -635 2124 -633
rect 2123 -641 2124 -639
rect 2130 -635 2131 -633
rect 2130 -641 2131 -639
rect 2137 -635 2138 -633
rect 2137 -641 2138 -639
rect 2144 -635 2145 -633
rect 2144 -641 2145 -639
rect 2151 -635 2152 -633
rect 2151 -641 2152 -639
rect 2158 -635 2159 -633
rect 2158 -641 2159 -639
rect 2165 -635 2166 -633
rect 2165 -641 2166 -639
rect 2172 -635 2173 -633
rect 2172 -641 2173 -639
rect 2179 -635 2180 -633
rect 2179 -641 2180 -639
rect 2186 -635 2187 -633
rect 2186 -641 2187 -639
rect 2193 -635 2194 -633
rect 2193 -641 2194 -639
rect 2200 -635 2201 -633
rect 2200 -641 2201 -639
rect 2207 -635 2208 -633
rect 2210 -635 2211 -633
rect 2207 -641 2208 -639
rect 2214 -635 2215 -633
rect 2214 -641 2215 -639
rect 2217 -641 2218 -639
rect 2221 -635 2222 -633
rect 2224 -635 2225 -633
rect 2224 -641 2225 -639
rect 2291 -635 2292 -633
rect 2291 -641 2292 -639
rect 2326 -635 2327 -633
rect 2326 -641 2327 -639
rect 2361 -635 2362 -633
rect 2361 -641 2362 -639
rect 2 -812 3 -810
rect 2 -818 3 -816
rect 12 -812 13 -810
rect 9 -818 10 -816
rect 19 -812 20 -810
rect 16 -818 17 -816
rect 19 -818 20 -816
rect 23 -812 24 -810
rect 23 -818 24 -816
rect 30 -812 31 -810
rect 30 -818 31 -816
rect 37 -812 38 -810
rect 37 -818 38 -816
rect 44 -812 45 -810
rect 47 -812 48 -810
rect 44 -818 45 -816
rect 47 -818 48 -816
rect 51 -812 52 -810
rect 51 -818 52 -816
rect 58 -812 59 -810
rect 58 -818 59 -816
rect 65 -812 66 -810
rect 68 -812 69 -810
rect 65 -818 66 -816
rect 72 -812 73 -810
rect 72 -818 73 -816
rect 79 -812 80 -810
rect 82 -812 83 -810
rect 79 -818 80 -816
rect 86 -812 87 -810
rect 86 -818 87 -816
rect 93 -812 94 -810
rect 93 -818 94 -816
rect 100 -812 101 -810
rect 100 -818 101 -816
rect 107 -812 108 -810
rect 107 -818 108 -816
rect 114 -812 115 -810
rect 114 -818 115 -816
rect 121 -818 122 -816
rect 124 -818 125 -816
rect 128 -812 129 -810
rect 131 -812 132 -810
rect 128 -818 129 -816
rect 135 -812 136 -810
rect 135 -818 136 -816
rect 142 -812 143 -810
rect 145 -812 146 -810
rect 145 -818 146 -816
rect 149 -812 150 -810
rect 149 -818 150 -816
rect 156 -812 157 -810
rect 156 -818 157 -816
rect 163 -812 164 -810
rect 163 -818 164 -816
rect 170 -812 171 -810
rect 170 -818 171 -816
rect 177 -812 178 -810
rect 177 -818 178 -816
rect 184 -812 185 -810
rect 187 -812 188 -810
rect 184 -818 185 -816
rect 187 -818 188 -816
rect 191 -812 192 -810
rect 191 -818 192 -816
rect 198 -812 199 -810
rect 198 -818 199 -816
rect 205 -812 206 -810
rect 208 -812 209 -810
rect 205 -818 206 -816
rect 212 -812 213 -810
rect 212 -818 213 -816
rect 219 -812 220 -810
rect 222 -812 223 -810
rect 222 -818 223 -816
rect 226 -812 227 -810
rect 226 -818 227 -816
rect 233 -812 234 -810
rect 236 -812 237 -810
rect 233 -818 234 -816
rect 240 -812 241 -810
rect 240 -818 241 -816
rect 247 -812 248 -810
rect 247 -818 248 -816
rect 254 -812 255 -810
rect 254 -818 255 -816
rect 261 -812 262 -810
rect 261 -818 262 -816
rect 268 -812 269 -810
rect 268 -818 269 -816
rect 275 -812 276 -810
rect 275 -818 276 -816
rect 282 -812 283 -810
rect 282 -818 283 -816
rect 289 -812 290 -810
rect 289 -818 290 -816
rect 296 -812 297 -810
rect 296 -818 297 -816
rect 303 -812 304 -810
rect 303 -818 304 -816
rect 310 -812 311 -810
rect 310 -818 311 -816
rect 317 -812 318 -810
rect 317 -818 318 -816
rect 324 -812 325 -810
rect 324 -818 325 -816
rect 331 -812 332 -810
rect 331 -818 332 -816
rect 338 -812 339 -810
rect 338 -818 339 -816
rect 345 -812 346 -810
rect 345 -818 346 -816
rect 352 -812 353 -810
rect 352 -818 353 -816
rect 359 -812 360 -810
rect 362 -812 363 -810
rect 359 -818 360 -816
rect 362 -818 363 -816
rect 366 -812 367 -810
rect 366 -818 367 -816
rect 373 -812 374 -810
rect 373 -818 374 -816
rect 380 -812 381 -810
rect 380 -818 381 -816
rect 387 -812 388 -810
rect 387 -818 388 -816
rect 394 -812 395 -810
rect 394 -818 395 -816
rect 401 -812 402 -810
rect 401 -818 402 -816
rect 408 -812 409 -810
rect 408 -818 409 -816
rect 415 -812 416 -810
rect 415 -818 416 -816
rect 422 -812 423 -810
rect 422 -818 423 -816
rect 429 -812 430 -810
rect 429 -818 430 -816
rect 436 -812 437 -810
rect 436 -818 437 -816
rect 443 -812 444 -810
rect 443 -818 444 -816
rect 450 -812 451 -810
rect 450 -818 451 -816
rect 457 -812 458 -810
rect 457 -818 458 -816
rect 464 -812 465 -810
rect 464 -818 465 -816
rect 471 -812 472 -810
rect 471 -818 472 -816
rect 478 -812 479 -810
rect 478 -818 479 -816
rect 485 -812 486 -810
rect 485 -818 486 -816
rect 492 -812 493 -810
rect 492 -818 493 -816
rect 499 -812 500 -810
rect 499 -818 500 -816
rect 506 -812 507 -810
rect 506 -818 507 -816
rect 513 -812 514 -810
rect 513 -818 514 -816
rect 520 -812 521 -810
rect 523 -812 524 -810
rect 520 -818 521 -816
rect 527 -812 528 -810
rect 527 -818 528 -816
rect 534 -812 535 -810
rect 534 -818 535 -816
rect 541 -812 542 -810
rect 541 -818 542 -816
rect 548 -812 549 -810
rect 548 -818 549 -816
rect 555 -812 556 -810
rect 555 -818 556 -816
rect 562 -812 563 -810
rect 562 -818 563 -816
rect 569 -812 570 -810
rect 569 -818 570 -816
rect 576 -812 577 -810
rect 576 -818 577 -816
rect 583 -812 584 -810
rect 586 -812 587 -810
rect 583 -818 584 -816
rect 586 -818 587 -816
rect 590 -812 591 -810
rect 590 -818 591 -816
rect 593 -818 594 -816
rect 597 -812 598 -810
rect 597 -818 598 -816
rect 604 -812 605 -810
rect 604 -818 605 -816
rect 611 -812 612 -810
rect 611 -818 612 -816
rect 618 -812 619 -810
rect 618 -818 619 -816
rect 625 -812 626 -810
rect 625 -818 626 -816
rect 632 -812 633 -810
rect 632 -818 633 -816
rect 639 -812 640 -810
rect 639 -818 640 -816
rect 646 -812 647 -810
rect 646 -818 647 -816
rect 653 -812 654 -810
rect 653 -818 654 -816
rect 660 -812 661 -810
rect 660 -818 661 -816
rect 667 -812 668 -810
rect 667 -818 668 -816
rect 674 -812 675 -810
rect 674 -818 675 -816
rect 681 -812 682 -810
rect 684 -812 685 -810
rect 684 -818 685 -816
rect 688 -812 689 -810
rect 688 -818 689 -816
rect 698 -812 699 -810
rect 695 -818 696 -816
rect 698 -818 699 -816
rect 702 -812 703 -810
rect 702 -818 703 -816
rect 709 -812 710 -810
rect 709 -818 710 -816
rect 716 -812 717 -810
rect 716 -818 717 -816
rect 726 -812 727 -810
rect 723 -818 724 -816
rect 726 -818 727 -816
rect 730 -812 731 -810
rect 730 -818 731 -816
rect 737 -812 738 -810
rect 737 -818 738 -816
rect 744 -812 745 -810
rect 747 -812 748 -810
rect 744 -818 745 -816
rect 747 -818 748 -816
rect 751 -812 752 -810
rect 754 -812 755 -810
rect 751 -818 752 -816
rect 754 -818 755 -816
rect 758 -812 759 -810
rect 758 -818 759 -816
rect 765 -812 766 -810
rect 765 -818 766 -816
rect 772 -812 773 -810
rect 772 -818 773 -816
rect 779 -812 780 -810
rect 779 -818 780 -816
rect 786 -812 787 -810
rect 786 -818 787 -816
rect 793 -812 794 -810
rect 793 -818 794 -816
rect 800 -812 801 -810
rect 800 -818 801 -816
rect 807 -812 808 -810
rect 807 -818 808 -816
rect 814 -812 815 -810
rect 814 -818 815 -816
rect 821 -812 822 -810
rect 821 -818 822 -816
rect 828 -812 829 -810
rect 828 -818 829 -816
rect 831 -818 832 -816
rect 835 -812 836 -810
rect 835 -818 836 -816
rect 842 -812 843 -810
rect 842 -818 843 -816
rect 849 -812 850 -810
rect 849 -818 850 -816
rect 856 -812 857 -810
rect 856 -818 857 -816
rect 863 -812 864 -810
rect 863 -818 864 -816
rect 870 -812 871 -810
rect 870 -818 871 -816
rect 880 -812 881 -810
rect 877 -818 878 -816
rect 884 -812 885 -810
rect 884 -818 885 -816
rect 891 -812 892 -810
rect 891 -818 892 -816
rect 898 -812 899 -810
rect 898 -818 899 -816
rect 905 -812 906 -810
rect 905 -818 906 -816
rect 912 -812 913 -810
rect 912 -818 913 -816
rect 919 -812 920 -810
rect 919 -818 920 -816
rect 926 -812 927 -810
rect 926 -818 927 -816
rect 933 -812 934 -810
rect 933 -818 934 -816
rect 940 -812 941 -810
rect 940 -818 941 -816
rect 947 -812 948 -810
rect 947 -818 948 -816
rect 954 -812 955 -810
rect 957 -812 958 -810
rect 954 -818 955 -816
rect 957 -818 958 -816
rect 961 -812 962 -810
rect 961 -818 962 -816
rect 968 -812 969 -810
rect 968 -818 969 -816
rect 975 -812 976 -810
rect 975 -818 976 -816
rect 982 -812 983 -810
rect 982 -818 983 -816
rect 989 -812 990 -810
rect 989 -818 990 -816
rect 996 -812 997 -810
rect 996 -818 997 -816
rect 1003 -812 1004 -810
rect 1003 -818 1004 -816
rect 1010 -812 1011 -810
rect 1010 -818 1011 -816
rect 1013 -818 1014 -816
rect 1017 -812 1018 -810
rect 1017 -818 1018 -816
rect 1024 -812 1025 -810
rect 1024 -818 1025 -816
rect 1031 -812 1032 -810
rect 1031 -818 1032 -816
rect 1038 -812 1039 -810
rect 1038 -818 1039 -816
rect 1045 -812 1046 -810
rect 1045 -818 1046 -816
rect 1052 -812 1053 -810
rect 1052 -818 1053 -816
rect 1059 -812 1060 -810
rect 1059 -818 1060 -816
rect 1066 -812 1067 -810
rect 1066 -818 1067 -816
rect 1073 -812 1074 -810
rect 1073 -818 1074 -816
rect 1080 -812 1081 -810
rect 1080 -818 1081 -816
rect 1087 -812 1088 -810
rect 1087 -818 1088 -816
rect 1094 -812 1095 -810
rect 1094 -818 1095 -816
rect 1101 -812 1102 -810
rect 1101 -818 1102 -816
rect 1108 -812 1109 -810
rect 1111 -812 1112 -810
rect 1108 -818 1109 -816
rect 1111 -818 1112 -816
rect 1115 -812 1116 -810
rect 1115 -818 1116 -816
rect 1122 -812 1123 -810
rect 1122 -818 1123 -816
rect 1129 -812 1130 -810
rect 1129 -818 1130 -816
rect 1132 -818 1133 -816
rect 1136 -812 1137 -810
rect 1139 -812 1140 -810
rect 1136 -818 1137 -816
rect 1139 -818 1140 -816
rect 1143 -812 1144 -810
rect 1146 -812 1147 -810
rect 1143 -818 1144 -816
rect 1146 -818 1147 -816
rect 1150 -812 1151 -810
rect 1150 -818 1151 -816
rect 1157 -812 1158 -810
rect 1157 -818 1158 -816
rect 1160 -818 1161 -816
rect 1164 -812 1165 -810
rect 1164 -818 1165 -816
rect 1171 -812 1172 -810
rect 1174 -812 1175 -810
rect 1171 -818 1172 -816
rect 1174 -818 1175 -816
rect 1178 -812 1179 -810
rect 1178 -818 1179 -816
rect 1185 -812 1186 -810
rect 1185 -818 1186 -816
rect 1192 -812 1193 -810
rect 1192 -818 1193 -816
rect 1199 -812 1200 -810
rect 1199 -818 1200 -816
rect 1206 -812 1207 -810
rect 1209 -812 1210 -810
rect 1206 -818 1207 -816
rect 1209 -818 1210 -816
rect 1213 -812 1214 -810
rect 1213 -818 1214 -816
rect 1216 -818 1217 -816
rect 1220 -812 1221 -810
rect 1223 -812 1224 -810
rect 1220 -818 1221 -816
rect 1223 -818 1224 -816
rect 1227 -812 1228 -810
rect 1227 -818 1228 -816
rect 1234 -812 1235 -810
rect 1234 -818 1235 -816
rect 1241 -812 1242 -810
rect 1241 -818 1242 -816
rect 1248 -812 1249 -810
rect 1248 -818 1249 -816
rect 1255 -812 1256 -810
rect 1255 -818 1256 -816
rect 1262 -812 1263 -810
rect 1262 -818 1263 -816
rect 1269 -812 1270 -810
rect 1269 -818 1270 -816
rect 1276 -812 1277 -810
rect 1276 -818 1277 -816
rect 1283 -812 1284 -810
rect 1283 -818 1284 -816
rect 1290 -812 1291 -810
rect 1290 -818 1291 -816
rect 1297 -812 1298 -810
rect 1297 -818 1298 -816
rect 1304 -812 1305 -810
rect 1304 -818 1305 -816
rect 1311 -812 1312 -810
rect 1311 -818 1312 -816
rect 1318 -812 1319 -810
rect 1318 -818 1319 -816
rect 1325 -812 1326 -810
rect 1325 -818 1326 -816
rect 1332 -812 1333 -810
rect 1335 -818 1336 -816
rect 1339 -812 1340 -810
rect 1339 -818 1340 -816
rect 1346 -812 1347 -810
rect 1346 -818 1347 -816
rect 1353 -812 1354 -810
rect 1353 -818 1354 -816
rect 1360 -812 1361 -810
rect 1360 -818 1361 -816
rect 1363 -818 1364 -816
rect 1370 -812 1371 -810
rect 1367 -818 1368 -816
rect 1370 -818 1371 -816
rect 1374 -812 1375 -810
rect 1374 -818 1375 -816
rect 1381 -812 1382 -810
rect 1381 -818 1382 -816
rect 1388 -812 1389 -810
rect 1388 -818 1389 -816
rect 1395 -812 1396 -810
rect 1395 -818 1396 -816
rect 1402 -812 1403 -810
rect 1402 -818 1403 -816
rect 1409 -812 1410 -810
rect 1409 -818 1410 -816
rect 1416 -812 1417 -810
rect 1416 -818 1417 -816
rect 1423 -812 1424 -810
rect 1423 -818 1424 -816
rect 1430 -812 1431 -810
rect 1430 -818 1431 -816
rect 1437 -812 1438 -810
rect 1437 -818 1438 -816
rect 1444 -812 1445 -810
rect 1444 -818 1445 -816
rect 1451 -812 1452 -810
rect 1451 -818 1452 -816
rect 1458 -812 1459 -810
rect 1458 -818 1459 -816
rect 1465 -812 1466 -810
rect 1465 -818 1466 -816
rect 1472 -812 1473 -810
rect 1472 -818 1473 -816
rect 1479 -812 1480 -810
rect 1479 -818 1480 -816
rect 1486 -812 1487 -810
rect 1486 -818 1487 -816
rect 1493 -812 1494 -810
rect 1493 -818 1494 -816
rect 1500 -812 1501 -810
rect 1500 -818 1501 -816
rect 1507 -812 1508 -810
rect 1507 -818 1508 -816
rect 1514 -812 1515 -810
rect 1514 -818 1515 -816
rect 1521 -812 1522 -810
rect 1521 -818 1522 -816
rect 1528 -812 1529 -810
rect 1528 -818 1529 -816
rect 1535 -812 1536 -810
rect 1538 -812 1539 -810
rect 1535 -818 1536 -816
rect 1538 -818 1539 -816
rect 1542 -812 1543 -810
rect 1542 -818 1543 -816
rect 1549 -812 1550 -810
rect 1549 -818 1550 -816
rect 1556 -812 1557 -810
rect 1556 -818 1557 -816
rect 1563 -812 1564 -810
rect 1563 -818 1564 -816
rect 1570 -812 1571 -810
rect 1570 -818 1571 -816
rect 1577 -812 1578 -810
rect 1577 -818 1578 -816
rect 1584 -812 1585 -810
rect 1584 -818 1585 -816
rect 1591 -812 1592 -810
rect 1591 -818 1592 -816
rect 1598 -812 1599 -810
rect 1598 -818 1599 -816
rect 1605 -812 1606 -810
rect 1605 -818 1606 -816
rect 1612 -812 1613 -810
rect 1612 -818 1613 -816
rect 1619 -812 1620 -810
rect 1619 -818 1620 -816
rect 1626 -812 1627 -810
rect 1626 -818 1627 -816
rect 1633 -812 1634 -810
rect 1633 -818 1634 -816
rect 1640 -812 1641 -810
rect 1640 -818 1641 -816
rect 1647 -812 1648 -810
rect 1647 -818 1648 -816
rect 1654 -812 1655 -810
rect 1654 -818 1655 -816
rect 1661 -812 1662 -810
rect 1661 -818 1662 -816
rect 1668 -812 1669 -810
rect 1668 -818 1669 -816
rect 1675 -812 1676 -810
rect 1675 -818 1676 -816
rect 1682 -812 1683 -810
rect 1682 -818 1683 -816
rect 1689 -812 1690 -810
rect 1689 -818 1690 -816
rect 1696 -812 1697 -810
rect 1696 -818 1697 -816
rect 1703 -812 1704 -810
rect 1703 -818 1704 -816
rect 1710 -812 1711 -810
rect 1710 -818 1711 -816
rect 1717 -812 1718 -810
rect 1717 -818 1718 -816
rect 1724 -812 1725 -810
rect 1724 -818 1725 -816
rect 1731 -812 1732 -810
rect 1731 -818 1732 -816
rect 1738 -812 1739 -810
rect 1738 -818 1739 -816
rect 1745 -812 1746 -810
rect 1745 -818 1746 -816
rect 1752 -812 1753 -810
rect 1752 -818 1753 -816
rect 1759 -812 1760 -810
rect 1759 -818 1760 -816
rect 1766 -812 1767 -810
rect 1766 -818 1767 -816
rect 1773 -812 1774 -810
rect 1773 -818 1774 -816
rect 1780 -812 1781 -810
rect 1780 -818 1781 -816
rect 1787 -812 1788 -810
rect 1787 -818 1788 -816
rect 1794 -812 1795 -810
rect 1794 -818 1795 -816
rect 1801 -812 1802 -810
rect 1801 -818 1802 -816
rect 1808 -812 1809 -810
rect 1808 -818 1809 -816
rect 1815 -812 1816 -810
rect 1815 -818 1816 -816
rect 1822 -812 1823 -810
rect 1822 -818 1823 -816
rect 1829 -812 1830 -810
rect 1829 -818 1830 -816
rect 1836 -812 1837 -810
rect 1836 -818 1837 -816
rect 1843 -812 1844 -810
rect 1843 -818 1844 -816
rect 1850 -812 1851 -810
rect 1850 -818 1851 -816
rect 1857 -812 1858 -810
rect 1857 -818 1858 -816
rect 1864 -812 1865 -810
rect 1864 -818 1865 -816
rect 1871 -812 1872 -810
rect 1871 -818 1872 -816
rect 1878 -812 1879 -810
rect 1878 -818 1879 -816
rect 1885 -812 1886 -810
rect 1885 -818 1886 -816
rect 1892 -812 1893 -810
rect 1892 -818 1893 -816
rect 1899 -812 1900 -810
rect 1899 -818 1900 -816
rect 1906 -812 1907 -810
rect 1906 -818 1907 -816
rect 1913 -812 1914 -810
rect 1913 -818 1914 -816
rect 1920 -812 1921 -810
rect 1920 -818 1921 -816
rect 1927 -812 1928 -810
rect 1927 -818 1928 -816
rect 1934 -812 1935 -810
rect 1934 -818 1935 -816
rect 1941 -812 1942 -810
rect 1941 -818 1942 -816
rect 1948 -812 1949 -810
rect 1948 -818 1949 -816
rect 1955 -812 1956 -810
rect 1955 -818 1956 -816
rect 1962 -812 1963 -810
rect 1962 -818 1963 -816
rect 1969 -812 1970 -810
rect 1969 -818 1970 -816
rect 1976 -812 1977 -810
rect 1976 -818 1977 -816
rect 1983 -812 1984 -810
rect 1983 -818 1984 -816
rect 1990 -812 1991 -810
rect 1990 -818 1991 -816
rect 1997 -812 1998 -810
rect 1997 -818 1998 -816
rect 2004 -812 2005 -810
rect 2004 -818 2005 -816
rect 2011 -812 2012 -810
rect 2011 -818 2012 -816
rect 2018 -812 2019 -810
rect 2018 -818 2019 -816
rect 2025 -812 2026 -810
rect 2025 -818 2026 -816
rect 2032 -812 2033 -810
rect 2032 -818 2033 -816
rect 2039 -812 2040 -810
rect 2039 -818 2040 -816
rect 2046 -812 2047 -810
rect 2046 -818 2047 -816
rect 2053 -812 2054 -810
rect 2053 -818 2054 -816
rect 2060 -812 2061 -810
rect 2060 -818 2061 -816
rect 2067 -812 2068 -810
rect 2067 -818 2068 -816
rect 2074 -812 2075 -810
rect 2074 -818 2075 -816
rect 2081 -812 2082 -810
rect 2081 -818 2082 -816
rect 2088 -812 2089 -810
rect 2088 -818 2089 -816
rect 2095 -812 2096 -810
rect 2095 -818 2096 -816
rect 2102 -812 2103 -810
rect 2102 -818 2103 -816
rect 2109 -812 2110 -810
rect 2109 -818 2110 -816
rect 2116 -812 2117 -810
rect 2116 -818 2117 -816
rect 2123 -812 2124 -810
rect 2123 -818 2124 -816
rect 2130 -812 2131 -810
rect 2130 -818 2131 -816
rect 2137 -812 2138 -810
rect 2137 -818 2138 -816
rect 2144 -812 2145 -810
rect 2144 -818 2145 -816
rect 2151 -812 2152 -810
rect 2151 -818 2152 -816
rect 2158 -812 2159 -810
rect 2158 -818 2159 -816
rect 2165 -812 2166 -810
rect 2165 -818 2166 -816
rect 2172 -812 2173 -810
rect 2172 -818 2173 -816
rect 2179 -812 2180 -810
rect 2179 -818 2180 -816
rect 2186 -812 2187 -810
rect 2186 -818 2187 -816
rect 2193 -812 2194 -810
rect 2193 -818 2194 -816
rect 2200 -812 2201 -810
rect 2200 -818 2201 -816
rect 2207 -812 2208 -810
rect 2207 -818 2208 -816
rect 2214 -812 2215 -810
rect 2214 -818 2215 -816
rect 2221 -812 2222 -810
rect 2221 -818 2222 -816
rect 2228 -812 2229 -810
rect 2228 -818 2229 -816
rect 2235 -812 2236 -810
rect 2235 -818 2236 -816
rect 2242 -812 2243 -810
rect 2242 -818 2243 -816
rect 2249 -812 2250 -810
rect 2249 -818 2250 -816
rect 2256 -812 2257 -810
rect 2256 -818 2257 -816
rect 2263 -812 2264 -810
rect 2263 -818 2264 -816
rect 2270 -812 2271 -810
rect 2270 -818 2271 -816
rect 2277 -812 2278 -810
rect 2277 -818 2278 -816
rect 2284 -812 2285 -810
rect 2284 -818 2285 -816
rect 2291 -812 2292 -810
rect 2291 -818 2292 -816
rect 2298 -812 2299 -810
rect 2298 -818 2299 -816
rect 2305 -812 2306 -810
rect 2305 -818 2306 -816
rect 2312 -812 2313 -810
rect 2312 -818 2313 -816
rect 2319 -812 2320 -810
rect 2319 -818 2320 -816
rect 2326 -812 2327 -810
rect 2326 -818 2327 -816
rect 2347 -812 2348 -810
rect 2347 -818 2348 -816
rect 2403 -812 2404 -810
rect 2403 -818 2404 -816
rect 2 -1001 3 -999
rect 2 -1007 3 -1005
rect 9 -1001 10 -999
rect 9 -1007 10 -1005
rect 16 -1001 17 -999
rect 16 -1007 17 -1005
rect 23 -1001 24 -999
rect 23 -1007 24 -1005
rect 30 -1001 31 -999
rect 30 -1007 31 -1005
rect 37 -1001 38 -999
rect 37 -1007 38 -1005
rect 44 -1001 45 -999
rect 44 -1007 45 -1005
rect 51 -1001 52 -999
rect 51 -1007 52 -1005
rect 58 -1001 59 -999
rect 58 -1007 59 -1005
rect 65 -1001 66 -999
rect 65 -1007 66 -1005
rect 72 -1001 73 -999
rect 72 -1007 73 -1005
rect 79 -1001 80 -999
rect 79 -1007 80 -1005
rect 86 -1001 87 -999
rect 86 -1007 87 -1005
rect 93 -1007 94 -1005
rect 96 -1007 97 -1005
rect 100 -1001 101 -999
rect 103 -1001 104 -999
rect 100 -1007 101 -1005
rect 103 -1007 104 -1005
rect 107 -1001 108 -999
rect 107 -1007 108 -1005
rect 114 -1001 115 -999
rect 114 -1007 115 -1005
rect 121 -1001 122 -999
rect 121 -1007 122 -1005
rect 128 -1001 129 -999
rect 128 -1007 129 -1005
rect 135 -1001 136 -999
rect 135 -1007 136 -1005
rect 138 -1007 139 -1005
rect 142 -1001 143 -999
rect 142 -1007 143 -1005
rect 149 -1001 150 -999
rect 149 -1007 150 -1005
rect 156 -1001 157 -999
rect 156 -1007 157 -1005
rect 163 -1001 164 -999
rect 163 -1007 164 -1005
rect 170 -1001 171 -999
rect 170 -1007 171 -1005
rect 177 -1001 178 -999
rect 180 -1001 181 -999
rect 177 -1007 178 -1005
rect 180 -1007 181 -1005
rect 184 -1001 185 -999
rect 187 -1001 188 -999
rect 187 -1007 188 -1005
rect 191 -1001 192 -999
rect 191 -1007 192 -1005
rect 198 -1001 199 -999
rect 198 -1007 199 -1005
rect 205 -1001 206 -999
rect 205 -1007 206 -1005
rect 212 -1001 213 -999
rect 212 -1007 213 -1005
rect 219 -1001 220 -999
rect 222 -1001 223 -999
rect 222 -1007 223 -1005
rect 226 -1001 227 -999
rect 226 -1007 227 -1005
rect 233 -1001 234 -999
rect 233 -1007 234 -1005
rect 240 -1001 241 -999
rect 240 -1007 241 -1005
rect 247 -1001 248 -999
rect 247 -1007 248 -1005
rect 254 -1001 255 -999
rect 254 -1007 255 -1005
rect 261 -1001 262 -999
rect 261 -1007 262 -1005
rect 268 -1001 269 -999
rect 271 -1001 272 -999
rect 271 -1007 272 -1005
rect 275 -1001 276 -999
rect 275 -1007 276 -1005
rect 282 -1001 283 -999
rect 282 -1007 283 -1005
rect 289 -1001 290 -999
rect 289 -1007 290 -1005
rect 296 -1001 297 -999
rect 296 -1007 297 -1005
rect 303 -1001 304 -999
rect 303 -1007 304 -1005
rect 310 -1001 311 -999
rect 310 -1007 311 -1005
rect 317 -1001 318 -999
rect 317 -1007 318 -1005
rect 324 -1001 325 -999
rect 324 -1007 325 -1005
rect 331 -1001 332 -999
rect 331 -1007 332 -1005
rect 338 -1001 339 -999
rect 338 -1007 339 -1005
rect 345 -1001 346 -999
rect 345 -1007 346 -1005
rect 352 -1001 353 -999
rect 352 -1007 353 -1005
rect 359 -1001 360 -999
rect 359 -1007 360 -1005
rect 366 -1001 367 -999
rect 366 -1007 367 -1005
rect 373 -1001 374 -999
rect 376 -1001 377 -999
rect 373 -1007 374 -1005
rect 376 -1007 377 -1005
rect 380 -1001 381 -999
rect 380 -1007 381 -1005
rect 387 -1001 388 -999
rect 390 -1001 391 -999
rect 390 -1007 391 -1005
rect 394 -1001 395 -999
rect 394 -1007 395 -1005
rect 401 -1001 402 -999
rect 401 -1007 402 -1005
rect 408 -1001 409 -999
rect 408 -1007 409 -1005
rect 415 -1001 416 -999
rect 415 -1007 416 -1005
rect 422 -1001 423 -999
rect 422 -1007 423 -1005
rect 429 -1001 430 -999
rect 429 -1007 430 -1005
rect 436 -1001 437 -999
rect 436 -1007 437 -1005
rect 443 -1001 444 -999
rect 443 -1007 444 -1005
rect 450 -1001 451 -999
rect 450 -1007 451 -1005
rect 457 -1001 458 -999
rect 457 -1007 458 -1005
rect 464 -1001 465 -999
rect 464 -1007 465 -1005
rect 471 -1001 472 -999
rect 471 -1007 472 -1005
rect 478 -1001 479 -999
rect 478 -1007 479 -1005
rect 485 -1001 486 -999
rect 485 -1007 486 -1005
rect 492 -1001 493 -999
rect 492 -1007 493 -1005
rect 499 -1001 500 -999
rect 499 -1007 500 -1005
rect 506 -1001 507 -999
rect 506 -1007 507 -1005
rect 513 -1001 514 -999
rect 513 -1007 514 -1005
rect 520 -1001 521 -999
rect 520 -1007 521 -1005
rect 527 -1001 528 -999
rect 530 -1001 531 -999
rect 534 -1001 535 -999
rect 534 -1007 535 -1005
rect 541 -1001 542 -999
rect 541 -1007 542 -1005
rect 548 -1001 549 -999
rect 548 -1007 549 -1005
rect 555 -1001 556 -999
rect 555 -1007 556 -1005
rect 562 -1001 563 -999
rect 562 -1007 563 -1005
rect 569 -1001 570 -999
rect 569 -1007 570 -1005
rect 576 -1001 577 -999
rect 576 -1007 577 -1005
rect 583 -1001 584 -999
rect 583 -1007 584 -1005
rect 590 -1001 591 -999
rect 590 -1007 591 -1005
rect 597 -1001 598 -999
rect 597 -1007 598 -1005
rect 604 -1001 605 -999
rect 604 -1007 605 -1005
rect 611 -1001 612 -999
rect 614 -1001 615 -999
rect 611 -1007 612 -1005
rect 618 -1001 619 -999
rect 618 -1007 619 -1005
rect 625 -1001 626 -999
rect 628 -1001 629 -999
rect 625 -1007 626 -1005
rect 628 -1007 629 -1005
rect 632 -1001 633 -999
rect 635 -1001 636 -999
rect 632 -1007 633 -1005
rect 635 -1007 636 -1005
rect 639 -1001 640 -999
rect 639 -1007 640 -1005
rect 646 -1001 647 -999
rect 646 -1007 647 -1005
rect 653 -1001 654 -999
rect 653 -1007 654 -1005
rect 660 -1001 661 -999
rect 660 -1007 661 -1005
rect 667 -1001 668 -999
rect 667 -1007 668 -1005
rect 674 -1001 675 -999
rect 674 -1007 675 -1005
rect 681 -1001 682 -999
rect 681 -1007 682 -1005
rect 688 -1001 689 -999
rect 688 -1007 689 -1005
rect 695 -1001 696 -999
rect 695 -1007 696 -1005
rect 702 -1001 703 -999
rect 702 -1007 703 -1005
rect 709 -1001 710 -999
rect 709 -1007 710 -1005
rect 716 -1001 717 -999
rect 719 -1001 720 -999
rect 719 -1007 720 -1005
rect 723 -1001 724 -999
rect 723 -1007 724 -1005
rect 730 -1001 731 -999
rect 730 -1007 731 -1005
rect 737 -1001 738 -999
rect 737 -1007 738 -1005
rect 744 -1001 745 -999
rect 744 -1007 745 -1005
rect 751 -1001 752 -999
rect 751 -1007 752 -1005
rect 758 -1001 759 -999
rect 758 -1007 759 -1005
rect 765 -1001 766 -999
rect 765 -1007 766 -1005
rect 772 -1001 773 -999
rect 775 -1001 776 -999
rect 772 -1007 773 -1005
rect 775 -1007 776 -1005
rect 782 -1001 783 -999
rect 779 -1007 780 -1005
rect 782 -1007 783 -1005
rect 786 -1001 787 -999
rect 786 -1007 787 -1005
rect 793 -1001 794 -999
rect 796 -1001 797 -999
rect 793 -1007 794 -1005
rect 796 -1007 797 -1005
rect 800 -1001 801 -999
rect 800 -1007 801 -1005
rect 807 -1001 808 -999
rect 807 -1007 808 -1005
rect 814 -1001 815 -999
rect 817 -1001 818 -999
rect 814 -1007 815 -1005
rect 817 -1007 818 -1005
rect 821 -1001 822 -999
rect 821 -1007 822 -1005
rect 828 -1001 829 -999
rect 828 -1007 829 -1005
rect 831 -1007 832 -1005
rect 835 -1001 836 -999
rect 835 -1007 836 -1005
rect 842 -1001 843 -999
rect 842 -1007 843 -1005
rect 849 -1001 850 -999
rect 849 -1007 850 -1005
rect 856 -1001 857 -999
rect 856 -1007 857 -1005
rect 863 -1001 864 -999
rect 863 -1007 864 -1005
rect 870 -1001 871 -999
rect 870 -1007 871 -1005
rect 877 -1001 878 -999
rect 877 -1007 878 -1005
rect 884 -1001 885 -999
rect 884 -1007 885 -1005
rect 891 -1001 892 -999
rect 891 -1007 892 -1005
rect 898 -1001 899 -999
rect 898 -1007 899 -1005
rect 905 -1001 906 -999
rect 905 -1007 906 -1005
rect 912 -1001 913 -999
rect 912 -1007 913 -1005
rect 919 -1001 920 -999
rect 919 -1007 920 -1005
rect 926 -1001 927 -999
rect 926 -1007 927 -1005
rect 933 -1001 934 -999
rect 936 -1001 937 -999
rect 936 -1007 937 -1005
rect 940 -1001 941 -999
rect 940 -1007 941 -1005
rect 947 -1001 948 -999
rect 947 -1007 948 -1005
rect 954 -1001 955 -999
rect 954 -1007 955 -1005
rect 957 -1007 958 -1005
rect 961 -1001 962 -999
rect 961 -1007 962 -1005
rect 968 -1001 969 -999
rect 968 -1007 969 -1005
rect 975 -1001 976 -999
rect 975 -1007 976 -1005
rect 982 -1001 983 -999
rect 982 -1007 983 -1005
rect 989 -1001 990 -999
rect 989 -1007 990 -1005
rect 996 -1001 997 -999
rect 996 -1007 997 -1005
rect 1003 -1001 1004 -999
rect 1003 -1007 1004 -1005
rect 1010 -1001 1011 -999
rect 1010 -1007 1011 -1005
rect 1017 -1001 1018 -999
rect 1020 -1001 1021 -999
rect 1017 -1007 1018 -1005
rect 1020 -1007 1021 -1005
rect 1024 -1001 1025 -999
rect 1024 -1007 1025 -1005
rect 1031 -1001 1032 -999
rect 1031 -1007 1032 -1005
rect 1041 -1001 1042 -999
rect 1038 -1007 1039 -1005
rect 1041 -1007 1042 -1005
rect 1045 -1001 1046 -999
rect 1045 -1007 1046 -1005
rect 1052 -1001 1053 -999
rect 1055 -1001 1056 -999
rect 1052 -1007 1053 -1005
rect 1055 -1007 1056 -1005
rect 1059 -1001 1060 -999
rect 1062 -1007 1063 -1005
rect 1066 -1001 1067 -999
rect 1066 -1007 1067 -1005
rect 1073 -1001 1074 -999
rect 1073 -1007 1074 -1005
rect 1080 -1001 1081 -999
rect 1080 -1007 1081 -1005
rect 1087 -1001 1088 -999
rect 1087 -1007 1088 -1005
rect 1094 -1001 1095 -999
rect 1094 -1007 1095 -1005
rect 1101 -1001 1102 -999
rect 1101 -1007 1102 -1005
rect 1108 -1001 1109 -999
rect 1108 -1007 1109 -1005
rect 1115 -1001 1116 -999
rect 1115 -1007 1116 -1005
rect 1122 -1001 1123 -999
rect 1125 -1001 1126 -999
rect 1122 -1007 1123 -1005
rect 1125 -1007 1126 -1005
rect 1129 -1001 1130 -999
rect 1129 -1007 1130 -1005
rect 1136 -1001 1137 -999
rect 1136 -1007 1137 -1005
rect 1143 -1001 1144 -999
rect 1143 -1007 1144 -1005
rect 1150 -1001 1151 -999
rect 1150 -1007 1151 -1005
rect 1157 -1001 1158 -999
rect 1157 -1007 1158 -1005
rect 1164 -1001 1165 -999
rect 1164 -1007 1165 -1005
rect 1171 -1001 1172 -999
rect 1174 -1001 1175 -999
rect 1171 -1007 1172 -1005
rect 1174 -1007 1175 -1005
rect 1178 -1001 1179 -999
rect 1178 -1007 1179 -1005
rect 1185 -1001 1186 -999
rect 1185 -1007 1186 -1005
rect 1192 -1001 1193 -999
rect 1195 -1001 1196 -999
rect 1192 -1007 1193 -1005
rect 1195 -1007 1196 -1005
rect 1199 -1001 1200 -999
rect 1199 -1007 1200 -1005
rect 1206 -1001 1207 -999
rect 1206 -1007 1207 -1005
rect 1213 -1001 1214 -999
rect 1213 -1007 1214 -1005
rect 1220 -1001 1221 -999
rect 1220 -1007 1221 -1005
rect 1227 -1001 1228 -999
rect 1227 -1007 1228 -1005
rect 1234 -1001 1235 -999
rect 1234 -1007 1235 -1005
rect 1241 -1001 1242 -999
rect 1244 -1001 1245 -999
rect 1241 -1007 1242 -1005
rect 1244 -1007 1245 -1005
rect 1248 -1001 1249 -999
rect 1248 -1007 1249 -1005
rect 1255 -1001 1256 -999
rect 1255 -1007 1256 -1005
rect 1262 -1001 1263 -999
rect 1262 -1007 1263 -1005
rect 1269 -1001 1270 -999
rect 1272 -1001 1273 -999
rect 1269 -1007 1270 -1005
rect 1272 -1007 1273 -1005
rect 1276 -1001 1277 -999
rect 1276 -1007 1277 -1005
rect 1283 -1001 1284 -999
rect 1286 -1001 1287 -999
rect 1283 -1007 1284 -1005
rect 1286 -1007 1287 -1005
rect 1290 -1001 1291 -999
rect 1290 -1007 1291 -1005
rect 1297 -1001 1298 -999
rect 1297 -1007 1298 -1005
rect 1304 -1001 1305 -999
rect 1304 -1007 1305 -1005
rect 1311 -1001 1312 -999
rect 1314 -1001 1315 -999
rect 1311 -1007 1312 -1005
rect 1314 -1007 1315 -1005
rect 1318 -1001 1319 -999
rect 1318 -1007 1319 -1005
rect 1325 -1001 1326 -999
rect 1325 -1007 1326 -1005
rect 1332 -1001 1333 -999
rect 1332 -1007 1333 -1005
rect 1339 -1001 1340 -999
rect 1339 -1007 1340 -1005
rect 1346 -1001 1347 -999
rect 1346 -1007 1347 -1005
rect 1353 -1001 1354 -999
rect 1353 -1007 1354 -1005
rect 1360 -1001 1361 -999
rect 1360 -1007 1361 -1005
rect 1367 -1001 1368 -999
rect 1367 -1007 1368 -1005
rect 1374 -1001 1375 -999
rect 1374 -1007 1375 -1005
rect 1381 -1001 1382 -999
rect 1381 -1007 1382 -1005
rect 1388 -1001 1389 -999
rect 1388 -1007 1389 -1005
rect 1395 -1001 1396 -999
rect 1398 -1001 1399 -999
rect 1395 -1007 1396 -1005
rect 1398 -1007 1399 -1005
rect 1402 -1001 1403 -999
rect 1402 -1007 1403 -1005
rect 1409 -1001 1410 -999
rect 1409 -1007 1410 -1005
rect 1416 -1001 1417 -999
rect 1416 -1007 1417 -1005
rect 1423 -1001 1424 -999
rect 1423 -1007 1424 -1005
rect 1430 -1001 1431 -999
rect 1430 -1007 1431 -1005
rect 1437 -1001 1438 -999
rect 1437 -1007 1438 -1005
rect 1444 -1001 1445 -999
rect 1444 -1007 1445 -1005
rect 1451 -1001 1452 -999
rect 1451 -1007 1452 -1005
rect 1458 -1001 1459 -999
rect 1458 -1007 1459 -1005
rect 1465 -1001 1466 -999
rect 1465 -1007 1466 -1005
rect 1472 -1001 1473 -999
rect 1472 -1007 1473 -1005
rect 1479 -1001 1480 -999
rect 1479 -1007 1480 -1005
rect 1486 -1001 1487 -999
rect 1486 -1007 1487 -1005
rect 1493 -1001 1494 -999
rect 1493 -1007 1494 -1005
rect 1500 -1001 1501 -999
rect 1500 -1007 1501 -1005
rect 1507 -1001 1508 -999
rect 1507 -1007 1508 -1005
rect 1514 -1001 1515 -999
rect 1517 -1001 1518 -999
rect 1514 -1007 1515 -1005
rect 1517 -1007 1518 -1005
rect 1521 -1001 1522 -999
rect 1521 -1007 1522 -1005
rect 1528 -1001 1529 -999
rect 1528 -1007 1529 -1005
rect 1535 -1001 1536 -999
rect 1535 -1007 1536 -1005
rect 1542 -1001 1543 -999
rect 1542 -1007 1543 -1005
rect 1549 -1001 1550 -999
rect 1549 -1007 1550 -1005
rect 1556 -1001 1557 -999
rect 1556 -1007 1557 -1005
rect 1563 -1001 1564 -999
rect 1563 -1007 1564 -1005
rect 1570 -1001 1571 -999
rect 1573 -1001 1574 -999
rect 1570 -1007 1571 -1005
rect 1577 -1001 1578 -999
rect 1580 -1007 1581 -1005
rect 1584 -1001 1585 -999
rect 1584 -1007 1585 -1005
rect 1591 -1001 1592 -999
rect 1591 -1007 1592 -1005
rect 1598 -1001 1599 -999
rect 1598 -1007 1599 -1005
rect 1605 -1001 1606 -999
rect 1605 -1007 1606 -1005
rect 1612 -1001 1613 -999
rect 1612 -1007 1613 -1005
rect 1619 -1001 1620 -999
rect 1619 -1007 1620 -1005
rect 1626 -1001 1627 -999
rect 1626 -1007 1627 -1005
rect 1633 -1001 1634 -999
rect 1633 -1007 1634 -1005
rect 1640 -1001 1641 -999
rect 1640 -1007 1641 -1005
rect 1647 -1001 1648 -999
rect 1647 -1007 1648 -1005
rect 1654 -1001 1655 -999
rect 1654 -1007 1655 -1005
rect 1661 -1001 1662 -999
rect 1661 -1007 1662 -1005
rect 1668 -1001 1669 -999
rect 1668 -1007 1669 -1005
rect 1675 -1001 1676 -999
rect 1675 -1007 1676 -1005
rect 1682 -1001 1683 -999
rect 1682 -1007 1683 -1005
rect 1689 -1001 1690 -999
rect 1689 -1007 1690 -1005
rect 1696 -1001 1697 -999
rect 1696 -1007 1697 -1005
rect 1703 -1001 1704 -999
rect 1703 -1007 1704 -1005
rect 1710 -1001 1711 -999
rect 1710 -1007 1711 -1005
rect 1717 -1001 1718 -999
rect 1717 -1007 1718 -1005
rect 1724 -1001 1725 -999
rect 1724 -1007 1725 -1005
rect 1731 -1001 1732 -999
rect 1731 -1007 1732 -1005
rect 1738 -1001 1739 -999
rect 1738 -1007 1739 -1005
rect 1745 -1001 1746 -999
rect 1745 -1007 1746 -1005
rect 1752 -1001 1753 -999
rect 1752 -1007 1753 -1005
rect 1759 -1001 1760 -999
rect 1759 -1007 1760 -1005
rect 1766 -1001 1767 -999
rect 1766 -1007 1767 -1005
rect 1773 -1001 1774 -999
rect 1773 -1007 1774 -1005
rect 1780 -1001 1781 -999
rect 1780 -1007 1781 -1005
rect 1787 -1001 1788 -999
rect 1787 -1007 1788 -1005
rect 1794 -1001 1795 -999
rect 1794 -1007 1795 -1005
rect 1801 -1001 1802 -999
rect 1801 -1007 1802 -1005
rect 1808 -1001 1809 -999
rect 1808 -1007 1809 -1005
rect 1815 -1001 1816 -999
rect 1815 -1007 1816 -1005
rect 1822 -1001 1823 -999
rect 1822 -1007 1823 -1005
rect 1829 -1001 1830 -999
rect 1829 -1007 1830 -1005
rect 1836 -1001 1837 -999
rect 1836 -1007 1837 -1005
rect 1843 -1001 1844 -999
rect 1843 -1007 1844 -1005
rect 1850 -1001 1851 -999
rect 1850 -1007 1851 -1005
rect 1857 -1001 1858 -999
rect 1857 -1007 1858 -1005
rect 1864 -1001 1865 -999
rect 1864 -1007 1865 -1005
rect 1871 -1001 1872 -999
rect 1871 -1007 1872 -1005
rect 1878 -1001 1879 -999
rect 1878 -1007 1879 -1005
rect 1885 -1001 1886 -999
rect 1885 -1007 1886 -1005
rect 1892 -1001 1893 -999
rect 1892 -1007 1893 -1005
rect 1899 -1001 1900 -999
rect 1899 -1007 1900 -1005
rect 1906 -1001 1907 -999
rect 1906 -1007 1907 -1005
rect 1913 -1001 1914 -999
rect 1913 -1007 1914 -1005
rect 1920 -1001 1921 -999
rect 1920 -1007 1921 -1005
rect 1927 -1001 1928 -999
rect 1927 -1007 1928 -1005
rect 1934 -1001 1935 -999
rect 1934 -1007 1935 -1005
rect 1941 -1001 1942 -999
rect 1941 -1007 1942 -1005
rect 1948 -1001 1949 -999
rect 1948 -1007 1949 -1005
rect 1955 -1001 1956 -999
rect 1955 -1007 1956 -1005
rect 1962 -1001 1963 -999
rect 1962 -1007 1963 -1005
rect 1969 -1001 1970 -999
rect 1969 -1007 1970 -1005
rect 1976 -1001 1977 -999
rect 1976 -1007 1977 -1005
rect 1983 -1001 1984 -999
rect 1983 -1007 1984 -1005
rect 1990 -1001 1991 -999
rect 1990 -1007 1991 -1005
rect 1997 -1001 1998 -999
rect 1997 -1007 1998 -1005
rect 2004 -1001 2005 -999
rect 2004 -1007 2005 -1005
rect 2011 -1001 2012 -999
rect 2011 -1007 2012 -1005
rect 2018 -1001 2019 -999
rect 2018 -1007 2019 -1005
rect 2025 -1001 2026 -999
rect 2025 -1007 2026 -1005
rect 2032 -1001 2033 -999
rect 2032 -1007 2033 -1005
rect 2039 -1001 2040 -999
rect 2039 -1007 2040 -1005
rect 2046 -1001 2047 -999
rect 2046 -1007 2047 -1005
rect 2053 -1001 2054 -999
rect 2053 -1007 2054 -1005
rect 2060 -1001 2061 -999
rect 2060 -1007 2061 -1005
rect 2067 -1001 2068 -999
rect 2067 -1007 2068 -1005
rect 2074 -1001 2075 -999
rect 2074 -1007 2075 -1005
rect 2081 -1001 2082 -999
rect 2081 -1007 2082 -1005
rect 2088 -1001 2089 -999
rect 2088 -1007 2089 -1005
rect 2095 -1001 2096 -999
rect 2095 -1007 2096 -1005
rect 2102 -1001 2103 -999
rect 2102 -1007 2103 -1005
rect 2109 -1001 2110 -999
rect 2109 -1007 2110 -1005
rect 2116 -1001 2117 -999
rect 2116 -1007 2117 -1005
rect 2123 -1001 2124 -999
rect 2123 -1007 2124 -1005
rect 2130 -1001 2131 -999
rect 2130 -1007 2131 -1005
rect 2137 -1001 2138 -999
rect 2137 -1007 2138 -1005
rect 2144 -1001 2145 -999
rect 2144 -1007 2145 -1005
rect 2151 -1001 2152 -999
rect 2151 -1007 2152 -1005
rect 2158 -1001 2159 -999
rect 2158 -1007 2159 -1005
rect 2165 -1001 2166 -999
rect 2165 -1007 2166 -1005
rect 2172 -1001 2173 -999
rect 2172 -1007 2173 -1005
rect 2179 -1001 2180 -999
rect 2179 -1007 2180 -1005
rect 2186 -1001 2187 -999
rect 2186 -1007 2187 -1005
rect 2193 -1001 2194 -999
rect 2193 -1007 2194 -1005
rect 2200 -1001 2201 -999
rect 2200 -1007 2201 -1005
rect 2207 -1001 2208 -999
rect 2207 -1007 2208 -1005
rect 2214 -1001 2215 -999
rect 2214 -1007 2215 -1005
rect 2221 -1001 2222 -999
rect 2221 -1007 2222 -1005
rect 2228 -1001 2229 -999
rect 2228 -1007 2229 -1005
rect 2235 -1001 2236 -999
rect 2235 -1007 2236 -1005
rect 2242 -1001 2243 -999
rect 2242 -1007 2243 -1005
rect 2249 -1001 2250 -999
rect 2249 -1007 2250 -1005
rect 2256 -1001 2257 -999
rect 2256 -1007 2257 -1005
rect 2263 -1001 2264 -999
rect 2263 -1007 2264 -1005
rect 2270 -1001 2271 -999
rect 2270 -1007 2271 -1005
rect 2277 -1001 2278 -999
rect 2277 -1007 2278 -1005
rect 2284 -1001 2285 -999
rect 2284 -1007 2285 -1005
rect 2291 -1001 2292 -999
rect 2291 -1007 2292 -1005
rect 2298 -1001 2299 -999
rect 2298 -1007 2299 -1005
rect 2305 -1001 2306 -999
rect 2305 -1007 2306 -1005
rect 2312 -1001 2313 -999
rect 2312 -1007 2313 -1005
rect 2319 -1001 2320 -999
rect 2319 -1007 2320 -1005
rect 2326 -1001 2327 -999
rect 2326 -1007 2327 -1005
rect 2336 -1001 2337 -999
rect 2333 -1007 2334 -1005
rect 2336 -1007 2337 -1005
rect 2340 -1001 2341 -999
rect 2343 -1001 2344 -999
rect 2343 -1007 2344 -1005
rect 2347 -1001 2348 -999
rect 2350 -1001 2351 -999
rect 2347 -1007 2348 -1005
rect 2354 -1001 2355 -999
rect 2354 -1007 2355 -1005
rect 2361 -1001 2362 -999
rect 2361 -1007 2362 -1005
rect 2368 -1001 2369 -999
rect 2368 -1007 2369 -1005
rect 2375 -1001 2376 -999
rect 2375 -1007 2376 -1005
rect 2403 -1001 2404 -999
rect 2403 -1007 2404 -1005
rect 2417 -1001 2418 -999
rect 2417 -1007 2418 -1005
rect 9 -1168 10 -1166
rect 9 -1174 10 -1172
rect 16 -1168 17 -1166
rect 16 -1174 17 -1172
rect 23 -1168 24 -1166
rect 23 -1174 24 -1172
rect 30 -1168 31 -1166
rect 30 -1174 31 -1172
rect 37 -1168 38 -1166
rect 37 -1174 38 -1172
rect 44 -1168 45 -1166
rect 44 -1174 45 -1172
rect 51 -1168 52 -1166
rect 51 -1174 52 -1172
rect 58 -1168 59 -1166
rect 58 -1174 59 -1172
rect 65 -1168 66 -1166
rect 65 -1174 66 -1172
rect 72 -1168 73 -1166
rect 72 -1174 73 -1172
rect 79 -1168 80 -1166
rect 79 -1174 80 -1172
rect 86 -1168 87 -1166
rect 89 -1168 90 -1166
rect 86 -1174 87 -1172
rect 89 -1174 90 -1172
rect 93 -1168 94 -1166
rect 93 -1174 94 -1172
rect 100 -1168 101 -1166
rect 100 -1174 101 -1172
rect 107 -1168 108 -1166
rect 110 -1168 111 -1166
rect 110 -1174 111 -1172
rect 114 -1168 115 -1166
rect 117 -1168 118 -1166
rect 114 -1174 115 -1172
rect 121 -1168 122 -1166
rect 121 -1174 122 -1172
rect 128 -1168 129 -1166
rect 128 -1174 129 -1172
rect 135 -1168 136 -1166
rect 138 -1168 139 -1166
rect 135 -1174 136 -1172
rect 138 -1174 139 -1172
rect 142 -1168 143 -1166
rect 145 -1168 146 -1166
rect 142 -1174 143 -1172
rect 145 -1174 146 -1172
rect 149 -1168 150 -1166
rect 149 -1174 150 -1172
rect 156 -1168 157 -1166
rect 156 -1174 157 -1172
rect 163 -1168 164 -1166
rect 163 -1174 164 -1172
rect 170 -1168 171 -1166
rect 170 -1174 171 -1172
rect 177 -1168 178 -1166
rect 177 -1174 178 -1172
rect 184 -1168 185 -1166
rect 184 -1174 185 -1172
rect 191 -1168 192 -1166
rect 191 -1174 192 -1172
rect 198 -1168 199 -1166
rect 198 -1174 199 -1172
rect 205 -1168 206 -1166
rect 205 -1174 206 -1172
rect 212 -1168 213 -1166
rect 212 -1174 213 -1172
rect 219 -1168 220 -1166
rect 219 -1174 220 -1172
rect 226 -1168 227 -1166
rect 226 -1174 227 -1172
rect 233 -1168 234 -1166
rect 233 -1174 234 -1172
rect 240 -1168 241 -1166
rect 240 -1174 241 -1172
rect 243 -1174 244 -1172
rect 247 -1168 248 -1166
rect 247 -1174 248 -1172
rect 254 -1168 255 -1166
rect 254 -1174 255 -1172
rect 261 -1168 262 -1166
rect 261 -1174 262 -1172
rect 268 -1168 269 -1166
rect 268 -1174 269 -1172
rect 275 -1168 276 -1166
rect 275 -1174 276 -1172
rect 282 -1168 283 -1166
rect 282 -1174 283 -1172
rect 289 -1168 290 -1166
rect 289 -1174 290 -1172
rect 296 -1168 297 -1166
rect 296 -1174 297 -1172
rect 303 -1168 304 -1166
rect 303 -1174 304 -1172
rect 310 -1168 311 -1166
rect 310 -1174 311 -1172
rect 317 -1168 318 -1166
rect 317 -1174 318 -1172
rect 324 -1168 325 -1166
rect 324 -1174 325 -1172
rect 331 -1168 332 -1166
rect 331 -1174 332 -1172
rect 338 -1168 339 -1166
rect 338 -1174 339 -1172
rect 345 -1168 346 -1166
rect 345 -1174 346 -1172
rect 352 -1168 353 -1166
rect 352 -1174 353 -1172
rect 359 -1168 360 -1166
rect 359 -1174 360 -1172
rect 366 -1168 367 -1166
rect 366 -1174 367 -1172
rect 373 -1168 374 -1166
rect 373 -1174 374 -1172
rect 380 -1168 381 -1166
rect 380 -1174 381 -1172
rect 387 -1168 388 -1166
rect 387 -1174 388 -1172
rect 394 -1168 395 -1166
rect 394 -1174 395 -1172
rect 401 -1168 402 -1166
rect 401 -1174 402 -1172
rect 408 -1168 409 -1166
rect 408 -1174 409 -1172
rect 415 -1168 416 -1166
rect 415 -1174 416 -1172
rect 422 -1168 423 -1166
rect 425 -1168 426 -1166
rect 422 -1174 423 -1172
rect 429 -1168 430 -1166
rect 432 -1168 433 -1166
rect 432 -1174 433 -1172
rect 436 -1168 437 -1166
rect 436 -1174 437 -1172
rect 443 -1168 444 -1166
rect 443 -1174 444 -1172
rect 450 -1168 451 -1166
rect 450 -1174 451 -1172
rect 457 -1168 458 -1166
rect 457 -1174 458 -1172
rect 464 -1168 465 -1166
rect 464 -1174 465 -1172
rect 471 -1168 472 -1166
rect 471 -1174 472 -1172
rect 478 -1168 479 -1166
rect 478 -1174 479 -1172
rect 485 -1168 486 -1166
rect 485 -1174 486 -1172
rect 492 -1168 493 -1166
rect 492 -1174 493 -1172
rect 499 -1168 500 -1166
rect 499 -1174 500 -1172
rect 506 -1168 507 -1166
rect 506 -1174 507 -1172
rect 509 -1174 510 -1172
rect 513 -1168 514 -1166
rect 513 -1174 514 -1172
rect 520 -1168 521 -1166
rect 520 -1174 521 -1172
rect 527 -1168 528 -1166
rect 527 -1174 528 -1172
rect 534 -1168 535 -1166
rect 534 -1174 535 -1172
rect 541 -1168 542 -1166
rect 541 -1174 542 -1172
rect 548 -1168 549 -1166
rect 548 -1174 549 -1172
rect 555 -1168 556 -1166
rect 555 -1174 556 -1172
rect 562 -1168 563 -1166
rect 562 -1174 563 -1172
rect 569 -1168 570 -1166
rect 569 -1174 570 -1172
rect 576 -1168 577 -1166
rect 576 -1174 577 -1172
rect 583 -1168 584 -1166
rect 583 -1174 584 -1172
rect 590 -1168 591 -1166
rect 593 -1168 594 -1166
rect 590 -1174 591 -1172
rect 597 -1168 598 -1166
rect 597 -1174 598 -1172
rect 604 -1168 605 -1166
rect 607 -1168 608 -1166
rect 607 -1174 608 -1172
rect 611 -1168 612 -1166
rect 611 -1174 612 -1172
rect 618 -1168 619 -1166
rect 618 -1174 619 -1172
rect 625 -1168 626 -1166
rect 625 -1174 626 -1172
rect 632 -1168 633 -1166
rect 632 -1174 633 -1172
rect 639 -1168 640 -1166
rect 639 -1174 640 -1172
rect 646 -1168 647 -1166
rect 646 -1174 647 -1172
rect 656 -1168 657 -1166
rect 653 -1174 654 -1172
rect 656 -1174 657 -1172
rect 660 -1168 661 -1166
rect 660 -1174 661 -1172
rect 667 -1168 668 -1166
rect 667 -1174 668 -1172
rect 674 -1168 675 -1166
rect 674 -1174 675 -1172
rect 681 -1168 682 -1166
rect 681 -1174 682 -1172
rect 688 -1168 689 -1166
rect 688 -1174 689 -1172
rect 695 -1168 696 -1166
rect 695 -1174 696 -1172
rect 702 -1168 703 -1166
rect 702 -1174 703 -1172
rect 709 -1168 710 -1166
rect 709 -1174 710 -1172
rect 716 -1168 717 -1166
rect 716 -1174 717 -1172
rect 723 -1168 724 -1166
rect 723 -1174 724 -1172
rect 730 -1168 731 -1166
rect 733 -1168 734 -1166
rect 730 -1174 731 -1172
rect 737 -1168 738 -1166
rect 737 -1174 738 -1172
rect 744 -1168 745 -1166
rect 744 -1174 745 -1172
rect 751 -1168 752 -1166
rect 751 -1174 752 -1172
rect 761 -1168 762 -1166
rect 758 -1174 759 -1172
rect 761 -1174 762 -1172
rect 765 -1168 766 -1166
rect 765 -1174 766 -1172
rect 772 -1168 773 -1166
rect 775 -1168 776 -1166
rect 772 -1174 773 -1172
rect 779 -1168 780 -1166
rect 779 -1174 780 -1172
rect 786 -1168 787 -1166
rect 786 -1174 787 -1172
rect 793 -1168 794 -1166
rect 793 -1174 794 -1172
rect 800 -1168 801 -1166
rect 800 -1174 801 -1172
rect 807 -1168 808 -1166
rect 807 -1174 808 -1172
rect 814 -1168 815 -1166
rect 814 -1174 815 -1172
rect 821 -1168 822 -1166
rect 824 -1168 825 -1166
rect 821 -1174 822 -1172
rect 824 -1174 825 -1172
rect 828 -1168 829 -1166
rect 828 -1174 829 -1172
rect 835 -1168 836 -1166
rect 835 -1174 836 -1172
rect 842 -1168 843 -1166
rect 842 -1174 843 -1172
rect 849 -1168 850 -1166
rect 852 -1174 853 -1172
rect 856 -1168 857 -1166
rect 856 -1174 857 -1172
rect 863 -1168 864 -1166
rect 866 -1168 867 -1166
rect 866 -1174 867 -1172
rect 870 -1168 871 -1166
rect 877 -1168 878 -1166
rect 880 -1168 881 -1166
rect 877 -1174 878 -1172
rect 880 -1174 881 -1172
rect 884 -1168 885 -1166
rect 884 -1174 885 -1172
rect 891 -1168 892 -1166
rect 891 -1174 892 -1172
rect 898 -1168 899 -1166
rect 898 -1174 899 -1172
rect 905 -1168 906 -1166
rect 908 -1174 909 -1172
rect 912 -1168 913 -1166
rect 912 -1174 913 -1172
rect 919 -1168 920 -1166
rect 919 -1174 920 -1172
rect 926 -1168 927 -1166
rect 926 -1174 927 -1172
rect 933 -1168 934 -1166
rect 933 -1174 934 -1172
rect 940 -1168 941 -1166
rect 940 -1174 941 -1172
rect 947 -1168 948 -1166
rect 950 -1168 951 -1166
rect 947 -1174 948 -1172
rect 950 -1174 951 -1172
rect 957 -1168 958 -1166
rect 954 -1174 955 -1172
rect 961 -1168 962 -1166
rect 964 -1168 965 -1166
rect 961 -1174 962 -1172
rect 964 -1174 965 -1172
rect 968 -1168 969 -1166
rect 968 -1174 969 -1172
rect 975 -1168 976 -1166
rect 975 -1174 976 -1172
rect 982 -1168 983 -1166
rect 982 -1174 983 -1172
rect 989 -1168 990 -1166
rect 989 -1174 990 -1172
rect 996 -1168 997 -1166
rect 996 -1174 997 -1172
rect 1003 -1168 1004 -1166
rect 1006 -1168 1007 -1166
rect 1003 -1174 1004 -1172
rect 1006 -1174 1007 -1172
rect 1010 -1168 1011 -1166
rect 1010 -1174 1011 -1172
rect 1017 -1168 1018 -1166
rect 1017 -1174 1018 -1172
rect 1024 -1168 1025 -1166
rect 1024 -1174 1025 -1172
rect 1031 -1168 1032 -1166
rect 1031 -1174 1032 -1172
rect 1038 -1168 1039 -1166
rect 1038 -1174 1039 -1172
rect 1045 -1168 1046 -1166
rect 1045 -1174 1046 -1172
rect 1048 -1174 1049 -1172
rect 1052 -1168 1053 -1166
rect 1052 -1174 1053 -1172
rect 1059 -1168 1060 -1166
rect 1059 -1174 1060 -1172
rect 1066 -1168 1067 -1166
rect 1066 -1174 1067 -1172
rect 1073 -1168 1074 -1166
rect 1073 -1174 1074 -1172
rect 1080 -1168 1081 -1166
rect 1080 -1174 1081 -1172
rect 1087 -1168 1088 -1166
rect 1087 -1174 1088 -1172
rect 1094 -1168 1095 -1166
rect 1094 -1174 1095 -1172
rect 1101 -1168 1102 -1166
rect 1101 -1174 1102 -1172
rect 1108 -1168 1109 -1166
rect 1108 -1174 1109 -1172
rect 1115 -1168 1116 -1166
rect 1115 -1174 1116 -1172
rect 1122 -1168 1123 -1166
rect 1122 -1174 1123 -1172
rect 1129 -1168 1130 -1166
rect 1129 -1174 1130 -1172
rect 1136 -1168 1137 -1166
rect 1136 -1174 1137 -1172
rect 1143 -1168 1144 -1166
rect 1143 -1174 1144 -1172
rect 1150 -1168 1151 -1166
rect 1150 -1174 1151 -1172
rect 1157 -1168 1158 -1166
rect 1160 -1168 1161 -1166
rect 1157 -1174 1158 -1172
rect 1160 -1174 1161 -1172
rect 1164 -1168 1165 -1166
rect 1167 -1168 1168 -1166
rect 1164 -1174 1165 -1172
rect 1167 -1174 1168 -1172
rect 1171 -1168 1172 -1166
rect 1171 -1174 1172 -1172
rect 1178 -1168 1179 -1166
rect 1181 -1168 1182 -1166
rect 1178 -1174 1179 -1172
rect 1181 -1174 1182 -1172
rect 1185 -1168 1186 -1166
rect 1185 -1174 1186 -1172
rect 1192 -1168 1193 -1166
rect 1192 -1174 1193 -1172
rect 1199 -1168 1200 -1166
rect 1202 -1168 1203 -1166
rect 1199 -1174 1200 -1172
rect 1202 -1174 1203 -1172
rect 1206 -1168 1207 -1166
rect 1206 -1174 1207 -1172
rect 1213 -1168 1214 -1166
rect 1213 -1174 1214 -1172
rect 1220 -1168 1221 -1166
rect 1223 -1168 1224 -1166
rect 1220 -1174 1221 -1172
rect 1227 -1168 1228 -1166
rect 1227 -1174 1228 -1172
rect 1234 -1168 1235 -1166
rect 1237 -1168 1238 -1166
rect 1234 -1174 1235 -1172
rect 1237 -1174 1238 -1172
rect 1241 -1168 1242 -1166
rect 1241 -1174 1242 -1172
rect 1248 -1168 1249 -1166
rect 1248 -1174 1249 -1172
rect 1255 -1168 1256 -1166
rect 1255 -1174 1256 -1172
rect 1262 -1168 1263 -1166
rect 1262 -1174 1263 -1172
rect 1269 -1168 1270 -1166
rect 1269 -1174 1270 -1172
rect 1276 -1168 1277 -1166
rect 1276 -1174 1277 -1172
rect 1283 -1168 1284 -1166
rect 1283 -1174 1284 -1172
rect 1290 -1168 1291 -1166
rect 1290 -1174 1291 -1172
rect 1297 -1168 1298 -1166
rect 1297 -1174 1298 -1172
rect 1304 -1168 1305 -1166
rect 1307 -1168 1308 -1166
rect 1304 -1174 1305 -1172
rect 1307 -1174 1308 -1172
rect 1311 -1168 1312 -1166
rect 1311 -1174 1312 -1172
rect 1318 -1168 1319 -1166
rect 1318 -1174 1319 -1172
rect 1325 -1168 1326 -1166
rect 1325 -1174 1326 -1172
rect 1332 -1168 1333 -1166
rect 1335 -1168 1336 -1166
rect 1332 -1174 1333 -1172
rect 1335 -1174 1336 -1172
rect 1339 -1168 1340 -1166
rect 1339 -1174 1340 -1172
rect 1346 -1168 1347 -1166
rect 1346 -1174 1347 -1172
rect 1353 -1168 1354 -1166
rect 1353 -1174 1354 -1172
rect 1360 -1168 1361 -1166
rect 1360 -1174 1361 -1172
rect 1367 -1168 1368 -1166
rect 1367 -1174 1368 -1172
rect 1374 -1168 1375 -1166
rect 1374 -1174 1375 -1172
rect 1381 -1168 1382 -1166
rect 1381 -1174 1382 -1172
rect 1388 -1168 1389 -1166
rect 1388 -1174 1389 -1172
rect 1391 -1174 1392 -1172
rect 1395 -1168 1396 -1166
rect 1395 -1174 1396 -1172
rect 1402 -1168 1403 -1166
rect 1402 -1174 1403 -1172
rect 1409 -1168 1410 -1166
rect 1409 -1174 1410 -1172
rect 1416 -1168 1417 -1166
rect 1416 -1174 1417 -1172
rect 1423 -1168 1424 -1166
rect 1423 -1174 1424 -1172
rect 1430 -1168 1431 -1166
rect 1430 -1174 1431 -1172
rect 1437 -1168 1438 -1166
rect 1437 -1174 1438 -1172
rect 1447 -1168 1448 -1166
rect 1444 -1174 1445 -1172
rect 1447 -1174 1448 -1172
rect 1451 -1168 1452 -1166
rect 1451 -1174 1452 -1172
rect 1458 -1168 1459 -1166
rect 1458 -1174 1459 -1172
rect 1465 -1168 1466 -1166
rect 1465 -1174 1466 -1172
rect 1472 -1168 1473 -1166
rect 1472 -1174 1473 -1172
rect 1479 -1168 1480 -1166
rect 1479 -1174 1480 -1172
rect 1486 -1168 1487 -1166
rect 1486 -1174 1487 -1172
rect 1493 -1168 1494 -1166
rect 1493 -1174 1494 -1172
rect 1500 -1168 1501 -1166
rect 1500 -1174 1501 -1172
rect 1507 -1168 1508 -1166
rect 1507 -1174 1508 -1172
rect 1514 -1168 1515 -1166
rect 1514 -1174 1515 -1172
rect 1521 -1168 1522 -1166
rect 1521 -1174 1522 -1172
rect 1528 -1168 1529 -1166
rect 1528 -1174 1529 -1172
rect 1535 -1168 1536 -1166
rect 1535 -1174 1536 -1172
rect 1542 -1168 1543 -1166
rect 1542 -1174 1543 -1172
rect 1549 -1168 1550 -1166
rect 1549 -1174 1550 -1172
rect 1552 -1174 1553 -1172
rect 1556 -1168 1557 -1166
rect 1556 -1174 1557 -1172
rect 1563 -1168 1564 -1166
rect 1563 -1174 1564 -1172
rect 1570 -1168 1571 -1166
rect 1570 -1174 1571 -1172
rect 1577 -1168 1578 -1166
rect 1577 -1174 1578 -1172
rect 1584 -1168 1585 -1166
rect 1584 -1174 1585 -1172
rect 1591 -1168 1592 -1166
rect 1591 -1174 1592 -1172
rect 1598 -1168 1599 -1166
rect 1598 -1174 1599 -1172
rect 1605 -1168 1606 -1166
rect 1605 -1174 1606 -1172
rect 1612 -1168 1613 -1166
rect 1612 -1174 1613 -1172
rect 1619 -1168 1620 -1166
rect 1619 -1174 1620 -1172
rect 1626 -1168 1627 -1166
rect 1626 -1174 1627 -1172
rect 1633 -1168 1634 -1166
rect 1633 -1174 1634 -1172
rect 1640 -1168 1641 -1166
rect 1640 -1174 1641 -1172
rect 1647 -1168 1648 -1166
rect 1647 -1174 1648 -1172
rect 1654 -1168 1655 -1166
rect 1654 -1174 1655 -1172
rect 1661 -1168 1662 -1166
rect 1661 -1174 1662 -1172
rect 1668 -1168 1669 -1166
rect 1668 -1174 1669 -1172
rect 1675 -1168 1676 -1166
rect 1675 -1174 1676 -1172
rect 1682 -1168 1683 -1166
rect 1682 -1174 1683 -1172
rect 1689 -1168 1690 -1166
rect 1689 -1174 1690 -1172
rect 1696 -1168 1697 -1166
rect 1696 -1174 1697 -1172
rect 1703 -1168 1704 -1166
rect 1703 -1174 1704 -1172
rect 1710 -1168 1711 -1166
rect 1710 -1174 1711 -1172
rect 1717 -1168 1718 -1166
rect 1717 -1174 1718 -1172
rect 1724 -1168 1725 -1166
rect 1724 -1174 1725 -1172
rect 1731 -1168 1732 -1166
rect 1731 -1174 1732 -1172
rect 1741 -1168 1742 -1166
rect 1738 -1174 1739 -1172
rect 1741 -1174 1742 -1172
rect 1745 -1168 1746 -1166
rect 1745 -1174 1746 -1172
rect 1752 -1168 1753 -1166
rect 1752 -1174 1753 -1172
rect 1759 -1168 1760 -1166
rect 1759 -1174 1760 -1172
rect 1766 -1168 1767 -1166
rect 1766 -1174 1767 -1172
rect 1773 -1168 1774 -1166
rect 1773 -1174 1774 -1172
rect 1780 -1168 1781 -1166
rect 1780 -1174 1781 -1172
rect 1787 -1168 1788 -1166
rect 1787 -1174 1788 -1172
rect 1794 -1168 1795 -1166
rect 1794 -1174 1795 -1172
rect 1801 -1168 1802 -1166
rect 1801 -1174 1802 -1172
rect 1808 -1168 1809 -1166
rect 1808 -1174 1809 -1172
rect 1815 -1168 1816 -1166
rect 1815 -1174 1816 -1172
rect 1822 -1168 1823 -1166
rect 1822 -1174 1823 -1172
rect 1829 -1168 1830 -1166
rect 1829 -1174 1830 -1172
rect 1836 -1168 1837 -1166
rect 1836 -1174 1837 -1172
rect 1843 -1168 1844 -1166
rect 1843 -1174 1844 -1172
rect 1850 -1168 1851 -1166
rect 1850 -1174 1851 -1172
rect 1857 -1168 1858 -1166
rect 1857 -1174 1858 -1172
rect 1864 -1168 1865 -1166
rect 1864 -1174 1865 -1172
rect 1871 -1168 1872 -1166
rect 1871 -1174 1872 -1172
rect 1878 -1168 1879 -1166
rect 1878 -1174 1879 -1172
rect 1885 -1168 1886 -1166
rect 1885 -1174 1886 -1172
rect 1892 -1168 1893 -1166
rect 1892 -1174 1893 -1172
rect 1899 -1168 1900 -1166
rect 1899 -1174 1900 -1172
rect 1906 -1168 1907 -1166
rect 1906 -1174 1907 -1172
rect 1913 -1168 1914 -1166
rect 1913 -1174 1914 -1172
rect 1920 -1168 1921 -1166
rect 1920 -1174 1921 -1172
rect 1927 -1168 1928 -1166
rect 1927 -1174 1928 -1172
rect 1934 -1168 1935 -1166
rect 1934 -1174 1935 -1172
rect 1941 -1168 1942 -1166
rect 1941 -1174 1942 -1172
rect 1948 -1168 1949 -1166
rect 1948 -1174 1949 -1172
rect 1955 -1168 1956 -1166
rect 1955 -1174 1956 -1172
rect 1962 -1168 1963 -1166
rect 1962 -1174 1963 -1172
rect 1969 -1168 1970 -1166
rect 1969 -1174 1970 -1172
rect 1976 -1168 1977 -1166
rect 1976 -1174 1977 -1172
rect 1983 -1168 1984 -1166
rect 1983 -1174 1984 -1172
rect 1990 -1168 1991 -1166
rect 1990 -1174 1991 -1172
rect 1997 -1168 1998 -1166
rect 1997 -1174 1998 -1172
rect 2004 -1168 2005 -1166
rect 2004 -1174 2005 -1172
rect 2011 -1168 2012 -1166
rect 2011 -1174 2012 -1172
rect 2018 -1168 2019 -1166
rect 2018 -1174 2019 -1172
rect 2025 -1168 2026 -1166
rect 2025 -1174 2026 -1172
rect 2032 -1168 2033 -1166
rect 2032 -1174 2033 -1172
rect 2039 -1168 2040 -1166
rect 2039 -1174 2040 -1172
rect 2046 -1168 2047 -1166
rect 2046 -1174 2047 -1172
rect 2053 -1168 2054 -1166
rect 2053 -1174 2054 -1172
rect 2060 -1168 2061 -1166
rect 2060 -1174 2061 -1172
rect 2067 -1168 2068 -1166
rect 2067 -1174 2068 -1172
rect 2074 -1168 2075 -1166
rect 2074 -1174 2075 -1172
rect 2081 -1168 2082 -1166
rect 2081 -1174 2082 -1172
rect 2088 -1168 2089 -1166
rect 2088 -1174 2089 -1172
rect 2095 -1168 2096 -1166
rect 2095 -1174 2096 -1172
rect 2102 -1168 2103 -1166
rect 2102 -1174 2103 -1172
rect 2109 -1168 2110 -1166
rect 2109 -1174 2110 -1172
rect 2116 -1168 2117 -1166
rect 2116 -1174 2117 -1172
rect 2123 -1168 2124 -1166
rect 2123 -1174 2124 -1172
rect 2130 -1168 2131 -1166
rect 2130 -1174 2131 -1172
rect 2137 -1168 2138 -1166
rect 2137 -1174 2138 -1172
rect 2144 -1168 2145 -1166
rect 2144 -1174 2145 -1172
rect 2151 -1168 2152 -1166
rect 2151 -1174 2152 -1172
rect 2158 -1168 2159 -1166
rect 2158 -1174 2159 -1172
rect 2165 -1168 2166 -1166
rect 2165 -1174 2166 -1172
rect 2172 -1168 2173 -1166
rect 2172 -1174 2173 -1172
rect 2179 -1168 2180 -1166
rect 2179 -1174 2180 -1172
rect 2186 -1168 2187 -1166
rect 2186 -1174 2187 -1172
rect 2193 -1168 2194 -1166
rect 2193 -1174 2194 -1172
rect 2200 -1168 2201 -1166
rect 2200 -1174 2201 -1172
rect 2207 -1168 2208 -1166
rect 2207 -1174 2208 -1172
rect 2214 -1168 2215 -1166
rect 2214 -1174 2215 -1172
rect 2221 -1168 2222 -1166
rect 2221 -1174 2222 -1172
rect 2228 -1168 2229 -1166
rect 2228 -1174 2229 -1172
rect 2235 -1168 2236 -1166
rect 2235 -1174 2236 -1172
rect 2242 -1168 2243 -1166
rect 2242 -1174 2243 -1172
rect 2249 -1168 2250 -1166
rect 2249 -1174 2250 -1172
rect 2256 -1168 2257 -1166
rect 2256 -1174 2257 -1172
rect 2263 -1168 2264 -1166
rect 2263 -1174 2264 -1172
rect 2270 -1168 2271 -1166
rect 2270 -1174 2271 -1172
rect 2277 -1168 2278 -1166
rect 2277 -1174 2278 -1172
rect 2284 -1168 2285 -1166
rect 2284 -1174 2285 -1172
rect 2291 -1168 2292 -1166
rect 2291 -1174 2292 -1172
rect 2298 -1168 2299 -1166
rect 2298 -1174 2299 -1172
rect 2305 -1168 2306 -1166
rect 2305 -1174 2306 -1172
rect 2312 -1168 2313 -1166
rect 2312 -1174 2313 -1172
rect 2319 -1168 2320 -1166
rect 2319 -1174 2320 -1172
rect 2326 -1168 2327 -1166
rect 2326 -1174 2327 -1172
rect 2333 -1168 2334 -1166
rect 2333 -1174 2334 -1172
rect 2340 -1168 2341 -1166
rect 2340 -1174 2341 -1172
rect 2347 -1168 2348 -1166
rect 2347 -1174 2348 -1172
rect 2354 -1168 2355 -1166
rect 2354 -1174 2355 -1172
rect 2361 -1168 2362 -1166
rect 2361 -1174 2362 -1172
rect 2368 -1168 2369 -1166
rect 2368 -1174 2369 -1172
rect 2375 -1168 2376 -1166
rect 2375 -1174 2376 -1172
rect 2382 -1168 2383 -1166
rect 2382 -1174 2383 -1172
rect 2389 -1168 2390 -1166
rect 2392 -1168 2393 -1166
rect 2389 -1174 2390 -1172
rect 2392 -1174 2393 -1172
rect 2396 -1168 2397 -1166
rect 2399 -1168 2400 -1166
rect 2396 -1174 2397 -1172
rect 2403 -1168 2404 -1166
rect 2403 -1174 2404 -1172
rect 2424 -1168 2425 -1166
rect 2424 -1174 2425 -1172
rect 2431 -1168 2432 -1166
rect 2431 -1174 2432 -1172
rect 2438 -1168 2439 -1166
rect 2438 -1174 2439 -1172
rect 5 -1351 6 -1349
rect 2 -1357 3 -1355
rect 9 -1351 10 -1349
rect 9 -1357 10 -1355
rect 19 -1351 20 -1349
rect 16 -1357 17 -1355
rect 23 -1351 24 -1349
rect 23 -1357 24 -1355
rect 30 -1351 31 -1349
rect 30 -1357 31 -1355
rect 37 -1351 38 -1349
rect 37 -1357 38 -1355
rect 44 -1351 45 -1349
rect 44 -1357 45 -1355
rect 51 -1351 52 -1349
rect 51 -1357 52 -1355
rect 58 -1351 59 -1349
rect 58 -1357 59 -1355
rect 65 -1351 66 -1349
rect 72 -1351 73 -1349
rect 72 -1357 73 -1355
rect 79 -1351 80 -1349
rect 82 -1357 83 -1355
rect 86 -1351 87 -1349
rect 86 -1357 87 -1355
rect 93 -1351 94 -1349
rect 93 -1357 94 -1355
rect 100 -1351 101 -1349
rect 100 -1357 101 -1355
rect 107 -1351 108 -1349
rect 107 -1357 108 -1355
rect 114 -1351 115 -1349
rect 114 -1357 115 -1355
rect 121 -1351 122 -1349
rect 124 -1351 125 -1349
rect 121 -1357 122 -1355
rect 124 -1357 125 -1355
rect 128 -1351 129 -1349
rect 128 -1357 129 -1355
rect 135 -1351 136 -1349
rect 135 -1357 136 -1355
rect 142 -1351 143 -1349
rect 142 -1357 143 -1355
rect 149 -1351 150 -1349
rect 149 -1357 150 -1355
rect 156 -1351 157 -1349
rect 156 -1357 157 -1355
rect 163 -1351 164 -1349
rect 163 -1357 164 -1355
rect 170 -1351 171 -1349
rect 170 -1357 171 -1355
rect 177 -1351 178 -1349
rect 177 -1357 178 -1355
rect 184 -1351 185 -1349
rect 184 -1357 185 -1355
rect 191 -1351 192 -1349
rect 191 -1357 192 -1355
rect 198 -1351 199 -1349
rect 198 -1357 199 -1355
rect 205 -1351 206 -1349
rect 208 -1351 209 -1349
rect 205 -1357 206 -1355
rect 208 -1357 209 -1355
rect 212 -1351 213 -1349
rect 212 -1357 213 -1355
rect 219 -1351 220 -1349
rect 219 -1357 220 -1355
rect 229 -1351 230 -1349
rect 226 -1357 227 -1355
rect 229 -1357 230 -1355
rect 233 -1351 234 -1349
rect 233 -1357 234 -1355
rect 240 -1351 241 -1349
rect 240 -1357 241 -1355
rect 247 -1351 248 -1349
rect 247 -1357 248 -1355
rect 250 -1357 251 -1355
rect 254 -1357 255 -1355
rect 257 -1357 258 -1355
rect 261 -1351 262 -1349
rect 261 -1357 262 -1355
rect 268 -1351 269 -1349
rect 271 -1357 272 -1355
rect 275 -1351 276 -1349
rect 275 -1357 276 -1355
rect 282 -1351 283 -1349
rect 282 -1357 283 -1355
rect 289 -1351 290 -1349
rect 289 -1357 290 -1355
rect 296 -1351 297 -1349
rect 296 -1357 297 -1355
rect 303 -1351 304 -1349
rect 303 -1357 304 -1355
rect 310 -1351 311 -1349
rect 310 -1357 311 -1355
rect 317 -1351 318 -1349
rect 317 -1357 318 -1355
rect 324 -1351 325 -1349
rect 324 -1357 325 -1355
rect 331 -1351 332 -1349
rect 331 -1357 332 -1355
rect 338 -1351 339 -1349
rect 338 -1357 339 -1355
rect 345 -1351 346 -1349
rect 345 -1357 346 -1355
rect 352 -1351 353 -1349
rect 352 -1357 353 -1355
rect 359 -1351 360 -1349
rect 359 -1357 360 -1355
rect 366 -1351 367 -1349
rect 366 -1357 367 -1355
rect 373 -1351 374 -1349
rect 373 -1357 374 -1355
rect 380 -1351 381 -1349
rect 380 -1357 381 -1355
rect 387 -1351 388 -1349
rect 387 -1357 388 -1355
rect 394 -1351 395 -1349
rect 394 -1357 395 -1355
rect 401 -1351 402 -1349
rect 401 -1357 402 -1355
rect 408 -1351 409 -1349
rect 408 -1357 409 -1355
rect 415 -1351 416 -1349
rect 415 -1357 416 -1355
rect 422 -1351 423 -1349
rect 422 -1357 423 -1355
rect 429 -1351 430 -1349
rect 429 -1357 430 -1355
rect 436 -1351 437 -1349
rect 436 -1357 437 -1355
rect 443 -1351 444 -1349
rect 443 -1357 444 -1355
rect 450 -1351 451 -1349
rect 450 -1357 451 -1355
rect 457 -1351 458 -1349
rect 457 -1357 458 -1355
rect 464 -1351 465 -1349
rect 464 -1357 465 -1355
rect 471 -1351 472 -1349
rect 471 -1357 472 -1355
rect 478 -1351 479 -1349
rect 478 -1357 479 -1355
rect 485 -1351 486 -1349
rect 485 -1357 486 -1355
rect 492 -1351 493 -1349
rect 492 -1357 493 -1355
rect 499 -1351 500 -1349
rect 499 -1357 500 -1355
rect 506 -1351 507 -1349
rect 506 -1357 507 -1355
rect 513 -1351 514 -1349
rect 513 -1357 514 -1355
rect 520 -1351 521 -1349
rect 520 -1357 521 -1355
rect 527 -1351 528 -1349
rect 527 -1357 528 -1355
rect 534 -1351 535 -1349
rect 534 -1357 535 -1355
rect 541 -1351 542 -1349
rect 541 -1357 542 -1355
rect 548 -1351 549 -1349
rect 548 -1357 549 -1355
rect 555 -1351 556 -1349
rect 555 -1357 556 -1355
rect 562 -1351 563 -1349
rect 562 -1357 563 -1355
rect 569 -1351 570 -1349
rect 569 -1357 570 -1355
rect 576 -1351 577 -1349
rect 576 -1357 577 -1355
rect 583 -1351 584 -1349
rect 583 -1357 584 -1355
rect 590 -1351 591 -1349
rect 590 -1357 591 -1355
rect 597 -1351 598 -1349
rect 597 -1357 598 -1355
rect 604 -1351 605 -1349
rect 607 -1351 608 -1349
rect 604 -1357 605 -1355
rect 607 -1357 608 -1355
rect 611 -1351 612 -1349
rect 611 -1357 612 -1355
rect 618 -1351 619 -1349
rect 618 -1357 619 -1355
rect 625 -1351 626 -1349
rect 625 -1357 626 -1355
rect 632 -1351 633 -1349
rect 632 -1357 633 -1355
rect 639 -1351 640 -1349
rect 642 -1351 643 -1349
rect 639 -1357 640 -1355
rect 642 -1357 643 -1355
rect 646 -1351 647 -1349
rect 646 -1357 647 -1355
rect 653 -1351 654 -1349
rect 653 -1357 654 -1355
rect 660 -1351 661 -1349
rect 660 -1357 661 -1355
rect 667 -1351 668 -1349
rect 667 -1357 668 -1355
rect 674 -1351 675 -1349
rect 677 -1351 678 -1349
rect 674 -1357 675 -1355
rect 677 -1357 678 -1355
rect 681 -1351 682 -1349
rect 681 -1357 682 -1355
rect 688 -1351 689 -1349
rect 688 -1357 689 -1355
rect 695 -1351 696 -1349
rect 695 -1357 696 -1355
rect 702 -1351 703 -1349
rect 702 -1357 703 -1355
rect 709 -1351 710 -1349
rect 709 -1357 710 -1355
rect 716 -1351 717 -1349
rect 716 -1357 717 -1355
rect 723 -1351 724 -1349
rect 726 -1351 727 -1349
rect 726 -1357 727 -1355
rect 730 -1351 731 -1349
rect 730 -1357 731 -1355
rect 737 -1351 738 -1349
rect 737 -1357 738 -1355
rect 744 -1351 745 -1349
rect 744 -1357 745 -1355
rect 751 -1351 752 -1349
rect 751 -1357 752 -1355
rect 758 -1351 759 -1349
rect 758 -1357 759 -1355
rect 765 -1351 766 -1349
rect 765 -1357 766 -1355
rect 772 -1351 773 -1349
rect 772 -1357 773 -1355
rect 779 -1351 780 -1349
rect 782 -1351 783 -1349
rect 779 -1357 780 -1355
rect 782 -1357 783 -1355
rect 786 -1351 787 -1349
rect 789 -1351 790 -1349
rect 786 -1357 787 -1355
rect 789 -1357 790 -1355
rect 793 -1351 794 -1349
rect 796 -1351 797 -1349
rect 796 -1357 797 -1355
rect 800 -1351 801 -1349
rect 800 -1357 801 -1355
rect 807 -1351 808 -1349
rect 807 -1357 808 -1355
rect 814 -1351 815 -1349
rect 814 -1357 815 -1355
rect 821 -1351 822 -1349
rect 821 -1357 822 -1355
rect 828 -1351 829 -1349
rect 831 -1351 832 -1349
rect 828 -1357 829 -1355
rect 831 -1357 832 -1355
rect 835 -1351 836 -1349
rect 835 -1357 836 -1355
rect 838 -1357 839 -1355
rect 842 -1351 843 -1349
rect 842 -1357 843 -1355
rect 849 -1351 850 -1349
rect 849 -1357 850 -1355
rect 856 -1351 857 -1349
rect 856 -1357 857 -1355
rect 863 -1351 864 -1349
rect 866 -1351 867 -1349
rect 866 -1357 867 -1355
rect 870 -1357 871 -1355
rect 880 -1351 881 -1349
rect 877 -1357 878 -1355
rect 880 -1357 881 -1355
rect 884 -1351 885 -1349
rect 884 -1357 885 -1355
rect 891 -1351 892 -1349
rect 894 -1351 895 -1349
rect 891 -1357 892 -1355
rect 894 -1357 895 -1355
rect 898 -1351 899 -1349
rect 898 -1357 899 -1355
rect 905 -1351 906 -1349
rect 905 -1357 906 -1355
rect 912 -1351 913 -1349
rect 912 -1357 913 -1355
rect 919 -1351 920 -1349
rect 919 -1357 920 -1355
rect 926 -1351 927 -1349
rect 926 -1357 927 -1355
rect 933 -1351 934 -1349
rect 933 -1357 934 -1355
rect 940 -1351 941 -1349
rect 940 -1357 941 -1355
rect 947 -1351 948 -1349
rect 947 -1357 948 -1355
rect 954 -1351 955 -1349
rect 957 -1351 958 -1349
rect 954 -1357 955 -1355
rect 957 -1357 958 -1355
rect 961 -1351 962 -1349
rect 961 -1357 962 -1355
rect 968 -1351 969 -1349
rect 968 -1357 969 -1355
rect 975 -1351 976 -1349
rect 975 -1357 976 -1355
rect 985 -1351 986 -1349
rect 982 -1357 983 -1355
rect 985 -1357 986 -1355
rect 989 -1351 990 -1349
rect 992 -1351 993 -1349
rect 989 -1357 990 -1355
rect 992 -1357 993 -1355
rect 996 -1351 997 -1349
rect 999 -1351 1000 -1349
rect 996 -1357 997 -1355
rect 999 -1357 1000 -1355
rect 1003 -1351 1004 -1349
rect 1006 -1351 1007 -1349
rect 1003 -1357 1004 -1355
rect 1006 -1357 1007 -1355
rect 1010 -1351 1011 -1349
rect 1013 -1351 1014 -1349
rect 1010 -1357 1011 -1355
rect 1013 -1357 1014 -1355
rect 1017 -1351 1018 -1349
rect 1017 -1357 1018 -1355
rect 1024 -1351 1025 -1349
rect 1024 -1357 1025 -1355
rect 1031 -1351 1032 -1349
rect 1031 -1357 1032 -1355
rect 1038 -1351 1039 -1349
rect 1041 -1351 1042 -1349
rect 1038 -1357 1039 -1355
rect 1041 -1357 1042 -1355
rect 1045 -1351 1046 -1349
rect 1045 -1357 1046 -1355
rect 1052 -1351 1053 -1349
rect 1052 -1357 1053 -1355
rect 1059 -1351 1060 -1349
rect 1059 -1357 1060 -1355
rect 1066 -1351 1067 -1349
rect 1066 -1357 1067 -1355
rect 1073 -1351 1074 -1349
rect 1073 -1357 1074 -1355
rect 1080 -1351 1081 -1349
rect 1080 -1357 1081 -1355
rect 1087 -1351 1088 -1349
rect 1087 -1357 1088 -1355
rect 1094 -1351 1095 -1349
rect 1094 -1357 1095 -1355
rect 1101 -1351 1102 -1349
rect 1104 -1351 1105 -1349
rect 1101 -1357 1102 -1355
rect 1104 -1357 1105 -1355
rect 1108 -1351 1109 -1349
rect 1108 -1357 1109 -1355
rect 1115 -1351 1116 -1349
rect 1115 -1357 1116 -1355
rect 1122 -1351 1123 -1349
rect 1122 -1357 1123 -1355
rect 1129 -1351 1130 -1349
rect 1129 -1357 1130 -1355
rect 1136 -1351 1137 -1349
rect 1136 -1357 1137 -1355
rect 1143 -1351 1144 -1349
rect 1143 -1357 1144 -1355
rect 1150 -1351 1151 -1349
rect 1153 -1351 1154 -1349
rect 1150 -1357 1151 -1355
rect 1153 -1357 1154 -1355
rect 1157 -1351 1158 -1349
rect 1157 -1357 1158 -1355
rect 1164 -1351 1165 -1349
rect 1164 -1357 1165 -1355
rect 1171 -1351 1172 -1349
rect 1171 -1357 1172 -1355
rect 1178 -1351 1179 -1349
rect 1178 -1357 1179 -1355
rect 1185 -1351 1186 -1349
rect 1185 -1357 1186 -1355
rect 1192 -1351 1193 -1349
rect 1192 -1357 1193 -1355
rect 1199 -1351 1200 -1349
rect 1199 -1357 1200 -1355
rect 1206 -1351 1207 -1349
rect 1206 -1357 1207 -1355
rect 1213 -1351 1214 -1349
rect 1216 -1351 1217 -1349
rect 1213 -1357 1214 -1355
rect 1220 -1351 1221 -1349
rect 1220 -1357 1221 -1355
rect 1227 -1351 1228 -1349
rect 1227 -1357 1228 -1355
rect 1234 -1351 1235 -1349
rect 1234 -1357 1235 -1355
rect 1241 -1351 1242 -1349
rect 1241 -1357 1242 -1355
rect 1248 -1351 1249 -1349
rect 1248 -1357 1249 -1355
rect 1255 -1351 1256 -1349
rect 1255 -1357 1256 -1355
rect 1262 -1351 1263 -1349
rect 1262 -1357 1263 -1355
rect 1269 -1351 1270 -1349
rect 1269 -1357 1270 -1355
rect 1276 -1351 1277 -1349
rect 1276 -1357 1277 -1355
rect 1283 -1351 1284 -1349
rect 1283 -1357 1284 -1355
rect 1290 -1351 1291 -1349
rect 1290 -1357 1291 -1355
rect 1297 -1351 1298 -1349
rect 1297 -1357 1298 -1355
rect 1304 -1351 1305 -1349
rect 1304 -1357 1305 -1355
rect 1311 -1351 1312 -1349
rect 1311 -1357 1312 -1355
rect 1318 -1351 1319 -1349
rect 1318 -1357 1319 -1355
rect 1325 -1351 1326 -1349
rect 1325 -1357 1326 -1355
rect 1332 -1351 1333 -1349
rect 1332 -1357 1333 -1355
rect 1339 -1351 1340 -1349
rect 1339 -1357 1340 -1355
rect 1346 -1351 1347 -1349
rect 1346 -1357 1347 -1355
rect 1353 -1351 1354 -1349
rect 1353 -1357 1354 -1355
rect 1360 -1351 1361 -1349
rect 1360 -1357 1361 -1355
rect 1367 -1351 1368 -1349
rect 1370 -1351 1371 -1349
rect 1367 -1357 1368 -1355
rect 1370 -1357 1371 -1355
rect 1374 -1351 1375 -1349
rect 1374 -1357 1375 -1355
rect 1381 -1351 1382 -1349
rect 1384 -1351 1385 -1349
rect 1381 -1357 1382 -1355
rect 1384 -1357 1385 -1355
rect 1388 -1351 1389 -1349
rect 1391 -1351 1392 -1349
rect 1388 -1357 1389 -1355
rect 1395 -1351 1396 -1349
rect 1395 -1357 1396 -1355
rect 1402 -1351 1403 -1349
rect 1402 -1357 1403 -1355
rect 1409 -1351 1410 -1349
rect 1409 -1357 1410 -1355
rect 1416 -1351 1417 -1349
rect 1416 -1357 1417 -1355
rect 1419 -1357 1420 -1355
rect 1423 -1351 1424 -1349
rect 1423 -1357 1424 -1355
rect 1430 -1351 1431 -1349
rect 1433 -1351 1434 -1349
rect 1430 -1357 1431 -1355
rect 1433 -1357 1434 -1355
rect 1437 -1351 1438 -1349
rect 1437 -1357 1438 -1355
rect 1447 -1351 1448 -1349
rect 1444 -1357 1445 -1355
rect 1451 -1351 1452 -1349
rect 1451 -1357 1452 -1355
rect 1458 -1351 1459 -1349
rect 1458 -1357 1459 -1355
rect 1465 -1351 1466 -1349
rect 1465 -1357 1466 -1355
rect 1472 -1351 1473 -1349
rect 1472 -1357 1473 -1355
rect 1479 -1351 1480 -1349
rect 1479 -1357 1480 -1355
rect 1486 -1351 1487 -1349
rect 1486 -1357 1487 -1355
rect 1493 -1351 1494 -1349
rect 1493 -1357 1494 -1355
rect 1500 -1351 1501 -1349
rect 1500 -1357 1501 -1355
rect 1507 -1351 1508 -1349
rect 1510 -1351 1511 -1349
rect 1510 -1357 1511 -1355
rect 1514 -1351 1515 -1349
rect 1514 -1357 1515 -1355
rect 1521 -1351 1522 -1349
rect 1521 -1357 1522 -1355
rect 1528 -1351 1529 -1349
rect 1528 -1357 1529 -1355
rect 1535 -1351 1536 -1349
rect 1535 -1357 1536 -1355
rect 1542 -1351 1543 -1349
rect 1542 -1357 1543 -1355
rect 1549 -1351 1550 -1349
rect 1549 -1357 1550 -1355
rect 1556 -1351 1557 -1349
rect 1556 -1357 1557 -1355
rect 1563 -1351 1564 -1349
rect 1563 -1357 1564 -1355
rect 1570 -1351 1571 -1349
rect 1570 -1357 1571 -1355
rect 1577 -1351 1578 -1349
rect 1577 -1357 1578 -1355
rect 1584 -1351 1585 -1349
rect 1584 -1357 1585 -1355
rect 1591 -1351 1592 -1349
rect 1591 -1357 1592 -1355
rect 1598 -1351 1599 -1349
rect 1598 -1357 1599 -1355
rect 1605 -1351 1606 -1349
rect 1605 -1357 1606 -1355
rect 1612 -1351 1613 -1349
rect 1612 -1357 1613 -1355
rect 1619 -1351 1620 -1349
rect 1619 -1357 1620 -1355
rect 1626 -1351 1627 -1349
rect 1626 -1357 1627 -1355
rect 1633 -1351 1634 -1349
rect 1633 -1357 1634 -1355
rect 1640 -1351 1641 -1349
rect 1640 -1357 1641 -1355
rect 1647 -1351 1648 -1349
rect 1647 -1357 1648 -1355
rect 1654 -1351 1655 -1349
rect 1654 -1357 1655 -1355
rect 1661 -1351 1662 -1349
rect 1661 -1357 1662 -1355
rect 1668 -1351 1669 -1349
rect 1668 -1357 1669 -1355
rect 1675 -1351 1676 -1349
rect 1675 -1357 1676 -1355
rect 1678 -1357 1679 -1355
rect 1682 -1351 1683 -1349
rect 1682 -1357 1683 -1355
rect 1689 -1351 1690 -1349
rect 1689 -1357 1690 -1355
rect 1696 -1351 1697 -1349
rect 1696 -1357 1697 -1355
rect 1703 -1351 1704 -1349
rect 1703 -1357 1704 -1355
rect 1710 -1351 1711 -1349
rect 1710 -1357 1711 -1355
rect 1717 -1351 1718 -1349
rect 1717 -1357 1718 -1355
rect 1724 -1351 1725 -1349
rect 1724 -1357 1725 -1355
rect 1731 -1351 1732 -1349
rect 1731 -1357 1732 -1355
rect 1738 -1351 1739 -1349
rect 1738 -1357 1739 -1355
rect 1745 -1351 1746 -1349
rect 1745 -1357 1746 -1355
rect 1752 -1351 1753 -1349
rect 1752 -1357 1753 -1355
rect 1759 -1351 1760 -1349
rect 1759 -1357 1760 -1355
rect 1766 -1351 1767 -1349
rect 1766 -1357 1767 -1355
rect 1773 -1351 1774 -1349
rect 1773 -1357 1774 -1355
rect 1780 -1351 1781 -1349
rect 1780 -1357 1781 -1355
rect 1787 -1351 1788 -1349
rect 1787 -1357 1788 -1355
rect 1794 -1351 1795 -1349
rect 1794 -1357 1795 -1355
rect 1797 -1357 1798 -1355
rect 1801 -1351 1802 -1349
rect 1801 -1357 1802 -1355
rect 1808 -1351 1809 -1349
rect 1808 -1357 1809 -1355
rect 1815 -1351 1816 -1349
rect 1815 -1357 1816 -1355
rect 1822 -1351 1823 -1349
rect 1822 -1357 1823 -1355
rect 1829 -1351 1830 -1349
rect 1829 -1357 1830 -1355
rect 1836 -1351 1837 -1349
rect 1836 -1357 1837 -1355
rect 1843 -1351 1844 -1349
rect 1843 -1357 1844 -1355
rect 1850 -1351 1851 -1349
rect 1850 -1357 1851 -1355
rect 1857 -1351 1858 -1349
rect 1857 -1357 1858 -1355
rect 1864 -1351 1865 -1349
rect 1864 -1357 1865 -1355
rect 1871 -1351 1872 -1349
rect 1871 -1357 1872 -1355
rect 1878 -1351 1879 -1349
rect 1878 -1357 1879 -1355
rect 1885 -1351 1886 -1349
rect 1885 -1357 1886 -1355
rect 1892 -1351 1893 -1349
rect 1892 -1357 1893 -1355
rect 1899 -1351 1900 -1349
rect 1899 -1357 1900 -1355
rect 1906 -1351 1907 -1349
rect 1906 -1357 1907 -1355
rect 1913 -1351 1914 -1349
rect 1913 -1357 1914 -1355
rect 1920 -1351 1921 -1349
rect 1920 -1357 1921 -1355
rect 1927 -1351 1928 -1349
rect 1927 -1357 1928 -1355
rect 1934 -1351 1935 -1349
rect 1934 -1357 1935 -1355
rect 1941 -1351 1942 -1349
rect 1941 -1357 1942 -1355
rect 1948 -1351 1949 -1349
rect 1948 -1357 1949 -1355
rect 1955 -1351 1956 -1349
rect 1955 -1357 1956 -1355
rect 1962 -1351 1963 -1349
rect 1962 -1357 1963 -1355
rect 1969 -1351 1970 -1349
rect 1969 -1357 1970 -1355
rect 1976 -1351 1977 -1349
rect 1976 -1357 1977 -1355
rect 1983 -1351 1984 -1349
rect 1983 -1357 1984 -1355
rect 1990 -1351 1991 -1349
rect 1990 -1357 1991 -1355
rect 1997 -1351 1998 -1349
rect 1997 -1357 1998 -1355
rect 2004 -1351 2005 -1349
rect 2004 -1357 2005 -1355
rect 2011 -1351 2012 -1349
rect 2011 -1357 2012 -1355
rect 2018 -1351 2019 -1349
rect 2018 -1357 2019 -1355
rect 2025 -1351 2026 -1349
rect 2025 -1357 2026 -1355
rect 2032 -1351 2033 -1349
rect 2032 -1357 2033 -1355
rect 2039 -1351 2040 -1349
rect 2039 -1357 2040 -1355
rect 2046 -1351 2047 -1349
rect 2046 -1357 2047 -1355
rect 2053 -1351 2054 -1349
rect 2053 -1357 2054 -1355
rect 2060 -1351 2061 -1349
rect 2060 -1357 2061 -1355
rect 2067 -1351 2068 -1349
rect 2067 -1357 2068 -1355
rect 2074 -1351 2075 -1349
rect 2074 -1357 2075 -1355
rect 2081 -1351 2082 -1349
rect 2081 -1357 2082 -1355
rect 2088 -1351 2089 -1349
rect 2088 -1357 2089 -1355
rect 2095 -1351 2096 -1349
rect 2095 -1357 2096 -1355
rect 2102 -1351 2103 -1349
rect 2102 -1357 2103 -1355
rect 2109 -1351 2110 -1349
rect 2109 -1357 2110 -1355
rect 2116 -1351 2117 -1349
rect 2116 -1357 2117 -1355
rect 2123 -1351 2124 -1349
rect 2123 -1357 2124 -1355
rect 2130 -1351 2131 -1349
rect 2130 -1357 2131 -1355
rect 2137 -1351 2138 -1349
rect 2137 -1357 2138 -1355
rect 2144 -1351 2145 -1349
rect 2144 -1357 2145 -1355
rect 2151 -1351 2152 -1349
rect 2151 -1357 2152 -1355
rect 2158 -1351 2159 -1349
rect 2158 -1357 2159 -1355
rect 2165 -1351 2166 -1349
rect 2165 -1357 2166 -1355
rect 2172 -1351 2173 -1349
rect 2172 -1357 2173 -1355
rect 2179 -1351 2180 -1349
rect 2179 -1357 2180 -1355
rect 2186 -1351 2187 -1349
rect 2186 -1357 2187 -1355
rect 2193 -1351 2194 -1349
rect 2193 -1357 2194 -1355
rect 2200 -1351 2201 -1349
rect 2200 -1357 2201 -1355
rect 2207 -1351 2208 -1349
rect 2207 -1357 2208 -1355
rect 2214 -1351 2215 -1349
rect 2214 -1357 2215 -1355
rect 2221 -1351 2222 -1349
rect 2221 -1357 2222 -1355
rect 2228 -1351 2229 -1349
rect 2228 -1357 2229 -1355
rect 2235 -1351 2236 -1349
rect 2235 -1357 2236 -1355
rect 2242 -1351 2243 -1349
rect 2242 -1357 2243 -1355
rect 2249 -1351 2250 -1349
rect 2249 -1357 2250 -1355
rect 2256 -1351 2257 -1349
rect 2256 -1357 2257 -1355
rect 2263 -1351 2264 -1349
rect 2263 -1357 2264 -1355
rect 2270 -1351 2271 -1349
rect 2270 -1357 2271 -1355
rect 2277 -1351 2278 -1349
rect 2277 -1357 2278 -1355
rect 2284 -1351 2285 -1349
rect 2284 -1357 2285 -1355
rect 2291 -1351 2292 -1349
rect 2291 -1357 2292 -1355
rect 2298 -1351 2299 -1349
rect 2298 -1357 2299 -1355
rect 2305 -1351 2306 -1349
rect 2305 -1357 2306 -1355
rect 2312 -1351 2313 -1349
rect 2312 -1357 2313 -1355
rect 2319 -1351 2320 -1349
rect 2319 -1357 2320 -1355
rect 2326 -1351 2327 -1349
rect 2326 -1357 2327 -1355
rect 2333 -1351 2334 -1349
rect 2333 -1357 2334 -1355
rect 2340 -1351 2341 -1349
rect 2343 -1351 2344 -1349
rect 2340 -1357 2341 -1355
rect 2343 -1357 2344 -1355
rect 2347 -1351 2348 -1349
rect 2347 -1357 2348 -1355
rect 2354 -1351 2355 -1349
rect 2354 -1357 2355 -1355
rect 2361 -1351 2362 -1349
rect 2361 -1357 2362 -1355
rect 2368 -1351 2369 -1349
rect 2368 -1357 2369 -1355
rect 2375 -1351 2376 -1349
rect 2375 -1357 2376 -1355
rect 2382 -1351 2383 -1349
rect 2382 -1357 2383 -1355
rect 2389 -1351 2390 -1349
rect 2389 -1357 2390 -1355
rect 2396 -1351 2397 -1349
rect 2396 -1357 2397 -1355
rect 2403 -1351 2404 -1349
rect 2403 -1357 2404 -1355
rect 2410 -1351 2411 -1349
rect 2410 -1357 2411 -1355
rect 2417 -1351 2418 -1349
rect 2417 -1357 2418 -1355
rect 2424 -1351 2425 -1349
rect 2424 -1357 2425 -1355
rect 2431 -1351 2432 -1349
rect 2431 -1357 2432 -1355
rect 2438 -1351 2439 -1349
rect 2438 -1357 2439 -1355
rect 2445 -1351 2446 -1349
rect 2445 -1357 2446 -1355
rect 2452 -1351 2453 -1349
rect 2452 -1357 2453 -1355
rect 2459 -1351 2460 -1349
rect 2459 -1357 2460 -1355
rect 2466 -1351 2467 -1349
rect 2466 -1357 2467 -1355
rect 2473 -1351 2474 -1349
rect 2473 -1357 2474 -1355
rect 2480 -1351 2481 -1349
rect 2480 -1357 2481 -1355
rect 2487 -1351 2488 -1349
rect 2487 -1357 2488 -1355
rect 2494 -1351 2495 -1349
rect 2494 -1357 2495 -1355
rect 2501 -1351 2502 -1349
rect 2501 -1357 2502 -1355
rect 2508 -1351 2509 -1349
rect 2508 -1357 2509 -1355
rect 2515 -1351 2516 -1349
rect 2515 -1357 2516 -1355
rect 2522 -1351 2523 -1349
rect 2522 -1357 2523 -1355
rect 2529 -1351 2530 -1349
rect 2529 -1357 2530 -1355
rect 2536 -1351 2537 -1349
rect 2536 -1357 2537 -1355
rect 2543 -1351 2544 -1349
rect 2543 -1357 2544 -1355
rect 2550 -1351 2551 -1349
rect 2550 -1357 2551 -1355
rect 2557 -1351 2558 -1349
rect 2557 -1357 2558 -1355
rect 2564 -1351 2565 -1349
rect 2564 -1357 2565 -1355
rect 2571 -1351 2572 -1349
rect 2571 -1357 2572 -1355
rect 2578 -1351 2579 -1349
rect 2578 -1357 2579 -1355
rect 2 -1528 3 -1526
rect 2 -1534 3 -1532
rect 9 -1528 10 -1526
rect 9 -1534 10 -1532
rect 16 -1528 17 -1526
rect 19 -1528 20 -1526
rect 23 -1528 24 -1526
rect 26 -1528 27 -1526
rect 23 -1534 24 -1532
rect 30 -1528 31 -1526
rect 30 -1534 31 -1532
rect 37 -1528 38 -1526
rect 40 -1528 41 -1526
rect 37 -1534 38 -1532
rect 40 -1534 41 -1532
rect 44 -1528 45 -1526
rect 47 -1528 48 -1526
rect 44 -1534 45 -1532
rect 47 -1534 48 -1532
rect 51 -1528 52 -1526
rect 54 -1528 55 -1526
rect 51 -1534 52 -1532
rect 58 -1528 59 -1526
rect 58 -1534 59 -1532
rect 65 -1534 66 -1532
rect 72 -1528 73 -1526
rect 72 -1534 73 -1532
rect 79 -1528 80 -1526
rect 79 -1534 80 -1532
rect 86 -1528 87 -1526
rect 89 -1528 90 -1526
rect 86 -1534 87 -1532
rect 89 -1534 90 -1532
rect 93 -1528 94 -1526
rect 93 -1534 94 -1532
rect 100 -1528 101 -1526
rect 100 -1534 101 -1532
rect 107 -1528 108 -1526
rect 110 -1528 111 -1526
rect 110 -1534 111 -1532
rect 114 -1528 115 -1526
rect 117 -1528 118 -1526
rect 114 -1534 115 -1532
rect 117 -1534 118 -1532
rect 121 -1528 122 -1526
rect 121 -1534 122 -1532
rect 128 -1528 129 -1526
rect 128 -1534 129 -1532
rect 135 -1528 136 -1526
rect 135 -1534 136 -1532
rect 142 -1528 143 -1526
rect 142 -1534 143 -1532
rect 149 -1528 150 -1526
rect 149 -1534 150 -1532
rect 156 -1528 157 -1526
rect 156 -1534 157 -1532
rect 163 -1528 164 -1526
rect 163 -1534 164 -1532
rect 170 -1528 171 -1526
rect 170 -1534 171 -1532
rect 177 -1528 178 -1526
rect 177 -1534 178 -1532
rect 184 -1528 185 -1526
rect 184 -1534 185 -1532
rect 191 -1528 192 -1526
rect 191 -1534 192 -1532
rect 198 -1528 199 -1526
rect 201 -1528 202 -1526
rect 198 -1534 199 -1532
rect 201 -1534 202 -1532
rect 208 -1528 209 -1526
rect 205 -1534 206 -1532
rect 208 -1534 209 -1532
rect 212 -1528 213 -1526
rect 212 -1534 213 -1532
rect 219 -1528 220 -1526
rect 219 -1534 220 -1532
rect 226 -1528 227 -1526
rect 226 -1534 227 -1532
rect 233 -1528 234 -1526
rect 236 -1528 237 -1526
rect 233 -1534 234 -1532
rect 236 -1534 237 -1532
rect 240 -1528 241 -1526
rect 240 -1534 241 -1532
rect 247 -1528 248 -1526
rect 247 -1534 248 -1532
rect 254 -1528 255 -1526
rect 254 -1534 255 -1532
rect 261 -1528 262 -1526
rect 261 -1534 262 -1532
rect 268 -1528 269 -1526
rect 268 -1534 269 -1532
rect 275 -1528 276 -1526
rect 275 -1534 276 -1532
rect 282 -1528 283 -1526
rect 282 -1534 283 -1532
rect 289 -1528 290 -1526
rect 289 -1534 290 -1532
rect 296 -1528 297 -1526
rect 296 -1534 297 -1532
rect 303 -1528 304 -1526
rect 303 -1534 304 -1532
rect 310 -1528 311 -1526
rect 310 -1534 311 -1532
rect 317 -1528 318 -1526
rect 317 -1534 318 -1532
rect 324 -1528 325 -1526
rect 324 -1534 325 -1532
rect 331 -1528 332 -1526
rect 331 -1534 332 -1532
rect 338 -1528 339 -1526
rect 338 -1534 339 -1532
rect 345 -1528 346 -1526
rect 345 -1534 346 -1532
rect 352 -1528 353 -1526
rect 352 -1534 353 -1532
rect 359 -1528 360 -1526
rect 359 -1534 360 -1532
rect 366 -1528 367 -1526
rect 366 -1534 367 -1532
rect 373 -1528 374 -1526
rect 373 -1534 374 -1532
rect 380 -1528 381 -1526
rect 380 -1534 381 -1532
rect 387 -1528 388 -1526
rect 387 -1534 388 -1532
rect 394 -1528 395 -1526
rect 394 -1534 395 -1532
rect 401 -1528 402 -1526
rect 401 -1534 402 -1532
rect 408 -1528 409 -1526
rect 408 -1534 409 -1532
rect 415 -1528 416 -1526
rect 415 -1534 416 -1532
rect 422 -1528 423 -1526
rect 422 -1534 423 -1532
rect 429 -1528 430 -1526
rect 429 -1534 430 -1532
rect 436 -1528 437 -1526
rect 436 -1534 437 -1532
rect 443 -1528 444 -1526
rect 443 -1534 444 -1532
rect 450 -1528 451 -1526
rect 450 -1534 451 -1532
rect 457 -1528 458 -1526
rect 457 -1534 458 -1532
rect 464 -1528 465 -1526
rect 464 -1534 465 -1532
rect 471 -1528 472 -1526
rect 471 -1534 472 -1532
rect 478 -1528 479 -1526
rect 478 -1534 479 -1532
rect 485 -1528 486 -1526
rect 485 -1534 486 -1532
rect 492 -1528 493 -1526
rect 492 -1534 493 -1532
rect 499 -1528 500 -1526
rect 499 -1534 500 -1532
rect 506 -1528 507 -1526
rect 506 -1534 507 -1532
rect 513 -1528 514 -1526
rect 516 -1528 517 -1526
rect 513 -1534 514 -1532
rect 516 -1534 517 -1532
rect 520 -1528 521 -1526
rect 520 -1534 521 -1532
rect 527 -1528 528 -1526
rect 527 -1534 528 -1532
rect 534 -1528 535 -1526
rect 534 -1534 535 -1532
rect 541 -1528 542 -1526
rect 541 -1534 542 -1532
rect 548 -1528 549 -1526
rect 548 -1534 549 -1532
rect 555 -1528 556 -1526
rect 555 -1534 556 -1532
rect 562 -1528 563 -1526
rect 562 -1534 563 -1532
rect 569 -1528 570 -1526
rect 569 -1534 570 -1532
rect 576 -1528 577 -1526
rect 576 -1534 577 -1532
rect 583 -1528 584 -1526
rect 583 -1534 584 -1532
rect 593 -1528 594 -1526
rect 590 -1534 591 -1532
rect 593 -1534 594 -1532
rect 597 -1528 598 -1526
rect 597 -1534 598 -1532
rect 604 -1528 605 -1526
rect 604 -1534 605 -1532
rect 611 -1528 612 -1526
rect 611 -1534 612 -1532
rect 618 -1528 619 -1526
rect 618 -1534 619 -1532
rect 625 -1528 626 -1526
rect 628 -1528 629 -1526
rect 625 -1534 626 -1532
rect 628 -1534 629 -1532
rect 632 -1528 633 -1526
rect 632 -1534 633 -1532
rect 639 -1528 640 -1526
rect 642 -1528 643 -1526
rect 639 -1534 640 -1532
rect 642 -1534 643 -1532
rect 646 -1528 647 -1526
rect 646 -1534 647 -1532
rect 653 -1528 654 -1526
rect 653 -1534 654 -1532
rect 660 -1528 661 -1526
rect 660 -1534 661 -1532
rect 667 -1528 668 -1526
rect 667 -1534 668 -1532
rect 674 -1528 675 -1526
rect 674 -1534 675 -1532
rect 681 -1528 682 -1526
rect 681 -1534 682 -1532
rect 688 -1528 689 -1526
rect 691 -1528 692 -1526
rect 688 -1534 689 -1532
rect 691 -1534 692 -1532
rect 695 -1528 696 -1526
rect 695 -1534 696 -1532
rect 702 -1528 703 -1526
rect 702 -1534 703 -1532
rect 709 -1528 710 -1526
rect 709 -1534 710 -1532
rect 716 -1528 717 -1526
rect 716 -1534 717 -1532
rect 723 -1528 724 -1526
rect 723 -1534 724 -1532
rect 730 -1528 731 -1526
rect 730 -1534 731 -1532
rect 737 -1528 738 -1526
rect 740 -1528 741 -1526
rect 737 -1534 738 -1532
rect 744 -1528 745 -1526
rect 744 -1534 745 -1532
rect 751 -1528 752 -1526
rect 751 -1534 752 -1532
rect 758 -1528 759 -1526
rect 758 -1534 759 -1532
rect 765 -1528 766 -1526
rect 765 -1534 766 -1532
rect 772 -1528 773 -1526
rect 772 -1534 773 -1532
rect 779 -1528 780 -1526
rect 779 -1534 780 -1532
rect 786 -1528 787 -1526
rect 786 -1534 787 -1532
rect 793 -1528 794 -1526
rect 796 -1528 797 -1526
rect 793 -1534 794 -1532
rect 796 -1534 797 -1532
rect 800 -1528 801 -1526
rect 800 -1534 801 -1532
rect 807 -1528 808 -1526
rect 807 -1534 808 -1532
rect 810 -1534 811 -1532
rect 814 -1528 815 -1526
rect 814 -1534 815 -1532
rect 824 -1528 825 -1526
rect 821 -1534 822 -1532
rect 824 -1534 825 -1532
rect 828 -1528 829 -1526
rect 828 -1534 829 -1532
rect 835 -1528 836 -1526
rect 835 -1534 836 -1532
rect 842 -1528 843 -1526
rect 842 -1534 843 -1532
rect 849 -1528 850 -1526
rect 849 -1534 850 -1532
rect 856 -1528 857 -1526
rect 856 -1534 857 -1532
rect 863 -1528 864 -1526
rect 866 -1528 867 -1526
rect 863 -1534 864 -1532
rect 866 -1534 867 -1532
rect 870 -1528 871 -1526
rect 870 -1534 871 -1532
rect 877 -1528 878 -1526
rect 880 -1528 881 -1526
rect 880 -1534 881 -1532
rect 884 -1528 885 -1526
rect 887 -1528 888 -1526
rect 887 -1534 888 -1532
rect 891 -1528 892 -1526
rect 891 -1534 892 -1532
rect 898 -1528 899 -1526
rect 898 -1534 899 -1532
rect 905 -1528 906 -1526
rect 908 -1528 909 -1526
rect 905 -1534 906 -1532
rect 912 -1528 913 -1526
rect 912 -1534 913 -1532
rect 919 -1528 920 -1526
rect 919 -1534 920 -1532
rect 926 -1528 927 -1526
rect 926 -1534 927 -1532
rect 933 -1528 934 -1526
rect 933 -1534 934 -1532
rect 940 -1528 941 -1526
rect 943 -1528 944 -1526
rect 940 -1534 941 -1532
rect 943 -1534 944 -1532
rect 947 -1528 948 -1526
rect 947 -1534 948 -1532
rect 954 -1528 955 -1526
rect 954 -1534 955 -1532
rect 961 -1528 962 -1526
rect 961 -1534 962 -1532
rect 964 -1534 965 -1532
rect 968 -1528 969 -1526
rect 968 -1534 969 -1532
rect 975 -1528 976 -1526
rect 975 -1534 976 -1532
rect 982 -1528 983 -1526
rect 982 -1534 983 -1532
rect 989 -1528 990 -1526
rect 989 -1534 990 -1532
rect 996 -1528 997 -1526
rect 996 -1534 997 -1532
rect 1003 -1528 1004 -1526
rect 1003 -1534 1004 -1532
rect 1010 -1528 1011 -1526
rect 1010 -1534 1011 -1532
rect 1017 -1528 1018 -1526
rect 1017 -1534 1018 -1532
rect 1024 -1528 1025 -1526
rect 1024 -1534 1025 -1532
rect 1031 -1528 1032 -1526
rect 1031 -1534 1032 -1532
rect 1038 -1528 1039 -1526
rect 1038 -1534 1039 -1532
rect 1045 -1528 1046 -1526
rect 1045 -1534 1046 -1532
rect 1052 -1528 1053 -1526
rect 1052 -1534 1053 -1532
rect 1059 -1528 1060 -1526
rect 1059 -1534 1060 -1532
rect 1066 -1528 1067 -1526
rect 1066 -1534 1067 -1532
rect 1073 -1528 1074 -1526
rect 1073 -1534 1074 -1532
rect 1080 -1528 1081 -1526
rect 1080 -1534 1081 -1532
rect 1087 -1528 1088 -1526
rect 1090 -1528 1091 -1526
rect 1087 -1534 1088 -1532
rect 1090 -1534 1091 -1532
rect 1094 -1528 1095 -1526
rect 1094 -1534 1095 -1532
rect 1101 -1528 1102 -1526
rect 1101 -1534 1102 -1532
rect 1108 -1528 1109 -1526
rect 1108 -1534 1109 -1532
rect 1115 -1528 1116 -1526
rect 1115 -1534 1116 -1532
rect 1122 -1528 1123 -1526
rect 1122 -1534 1123 -1532
rect 1129 -1528 1130 -1526
rect 1129 -1534 1130 -1532
rect 1136 -1528 1137 -1526
rect 1136 -1534 1137 -1532
rect 1143 -1528 1144 -1526
rect 1143 -1534 1144 -1532
rect 1150 -1528 1151 -1526
rect 1153 -1528 1154 -1526
rect 1150 -1534 1151 -1532
rect 1153 -1534 1154 -1532
rect 1157 -1528 1158 -1526
rect 1160 -1528 1161 -1526
rect 1157 -1534 1158 -1532
rect 1160 -1534 1161 -1532
rect 1164 -1528 1165 -1526
rect 1164 -1534 1165 -1532
rect 1171 -1528 1172 -1526
rect 1171 -1534 1172 -1532
rect 1178 -1528 1179 -1526
rect 1178 -1534 1179 -1532
rect 1185 -1528 1186 -1526
rect 1185 -1534 1186 -1532
rect 1192 -1528 1193 -1526
rect 1192 -1534 1193 -1532
rect 1199 -1528 1200 -1526
rect 1199 -1534 1200 -1532
rect 1206 -1528 1207 -1526
rect 1206 -1534 1207 -1532
rect 1213 -1528 1214 -1526
rect 1213 -1534 1214 -1532
rect 1220 -1528 1221 -1526
rect 1220 -1534 1221 -1532
rect 1227 -1528 1228 -1526
rect 1227 -1534 1228 -1532
rect 1234 -1528 1235 -1526
rect 1234 -1534 1235 -1532
rect 1241 -1528 1242 -1526
rect 1241 -1534 1242 -1532
rect 1248 -1528 1249 -1526
rect 1251 -1528 1252 -1526
rect 1248 -1534 1249 -1532
rect 1251 -1534 1252 -1532
rect 1255 -1528 1256 -1526
rect 1258 -1528 1259 -1526
rect 1258 -1534 1259 -1532
rect 1262 -1528 1263 -1526
rect 1265 -1528 1266 -1526
rect 1262 -1534 1263 -1532
rect 1269 -1528 1270 -1526
rect 1269 -1534 1270 -1532
rect 1276 -1528 1277 -1526
rect 1276 -1534 1277 -1532
rect 1283 -1528 1284 -1526
rect 1286 -1528 1287 -1526
rect 1286 -1534 1287 -1532
rect 1290 -1528 1291 -1526
rect 1290 -1534 1291 -1532
rect 1297 -1528 1298 -1526
rect 1297 -1534 1298 -1532
rect 1304 -1528 1305 -1526
rect 1304 -1534 1305 -1532
rect 1311 -1528 1312 -1526
rect 1311 -1534 1312 -1532
rect 1318 -1528 1319 -1526
rect 1318 -1534 1319 -1532
rect 1325 -1528 1326 -1526
rect 1325 -1534 1326 -1532
rect 1332 -1528 1333 -1526
rect 1332 -1534 1333 -1532
rect 1339 -1528 1340 -1526
rect 1339 -1534 1340 -1532
rect 1346 -1528 1347 -1526
rect 1349 -1528 1350 -1526
rect 1346 -1534 1347 -1532
rect 1349 -1534 1350 -1532
rect 1353 -1528 1354 -1526
rect 1353 -1534 1354 -1532
rect 1360 -1528 1361 -1526
rect 1360 -1534 1361 -1532
rect 1367 -1528 1368 -1526
rect 1367 -1534 1368 -1532
rect 1374 -1528 1375 -1526
rect 1374 -1534 1375 -1532
rect 1381 -1528 1382 -1526
rect 1381 -1534 1382 -1532
rect 1388 -1528 1389 -1526
rect 1388 -1534 1389 -1532
rect 1395 -1528 1396 -1526
rect 1395 -1534 1396 -1532
rect 1402 -1528 1403 -1526
rect 1402 -1534 1403 -1532
rect 1409 -1528 1410 -1526
rect 1409 -1534 1410 -1532
rect 1416 -1528 1417 -1526
rect 1416 -1534 1417 -1532
rect 1426 -1528 1427 -1526
rect 1423 -1534 1424 -1532
rect 1430 -1528 1431 -1526
rect 1430 -1534 1431 -1532
rect 1437 -1528 1438 -1526
rect 1437 -1534 1438 -1532
rect 1444 -1528 1445 -1526
rect 1444 -1534 1445 -1532
rect 1451 -1528 1452 -1526
rect 1451 -1534 1452 -1532
rect 1458 -1528 1459 -1526
rect 1458 -1534 1459 -1532
rect 1465 -1528 1466 -1526
rect 1465 -1534 1466 -1532
rect 1472 -1528 1473 -1526
rect 1472 -1534 1473 -1532
rect 1479 -1528 1480 -1526
rect 1482 -1528 1483 -1526
rect 1479 -1534 1480 -1532
rect 1486 -1528 1487 -1526
rect 1489 -1528 1490 -1526
rect 1489 -1534 1490 -1532
rect 1493 -1528 1494 -1526
rect 1493 -1534 1494 -1532
rect 1500 -1528 1501 -1526
rect 1503 -1528 1504 -1526
rect 1500 -1534 1501 -1532
rect 1503 -1534 1504 -1532
rect 1507 -1528 1508 -1526
rect 1507 -1534 1508 -1532
rect 1514 -1528 1515 -1526
rect 1514 -1534 1515 -1532
rect 1521 -1528 1522 -1526
rect 1521 -1534 1522 -1532
rect 1528 -1528 1529 -1526
rect 1528 -1534 1529 -1532
rect 1535 -1528 1536 -1526
rect 1535 -1534 1536 -1532
rect 1542 -1528 1543 -1526
rect 1542 -1534 1543 -1532
rect 1549 -1528 1550 -1526
rect 1549 -1534 1550 -1532
rect 1556 -1528 1557 -1526
rect 1556 -1534 1557 -1532
rect 1563 -1528 1564 -1526
rect 1563 -1534 1564 -1532
rect 1570 -1528 1571 -1526
rect 1570 -1534 1571 -1532
rect 1577 -1528 1578 -1526
rect 1577 -1534 1578 -1532
rect 1584 -1528 1585 -1526
rect 1584 -1534 1585 -1532
rect 1591 -1528 1592 -1526
rect 1591 -1534 1592 -1532
rect 1598 -1528 1599 -1526
rect 1598 -1534 1599 -1532
rect 1605 -1528 1606 -1526
rect 1605 -1534 1606 -1532
rect 1612 -1528 1613 -1526
rect 1612 -1534 1613 -1532
rect 1619 -1528 1620 -1526
rect 1619 -1534 1620 -1532
rect 1626 -1528 1627 -1526
rect 1626 -1534 1627 -1532
rect 1633 -1528 1634 -1526
rect 1633 -1534 1634 -1532
rect 1640 -1528 1641 -1526
rect 1640 -1534 1641 -1532
rect 1647 -1528 1648 -1526
rect 1647 -1534 1648 -1532
rect 1654 -1528 1655 -1526
rect 1654 -1534 1655 -1532
rect 1661 -1528 1662 -1526
rect 1661 -1534 1662 -1532
rect 1668 -1528 1669 -1526
rect 1668 -1534 1669 -1532
rect 1675 -1528 1676 -1526
rect 1675 -1534 1676 -1532
rect 1682 -1528 1683 -1526
rect 1682 -1534 1683 -1532
rect 1689 -1528 1690 -1526
rect 1689 -1534 1690 -1532
rect 1696 -1528 1697 -1526
rect 1696 -1534 1697 -1532
rect 1703 -1528 1704 -1526
rect 1703 -1534 1704 -1532
rect 1710 -1528 1711 -1526
rect 1710 -1534 1711 -1532
rect 1717 -1528 1718 -1526
rect 1717 -1534 1718 -1532
rect 1724 -1528 1725 -1526
rect 1724 -1534 1725 -1532
rect 1731 -1528 1732 -1526
rect 1731 -1534 1732 -1532
rect 1738 -1528 1739 -1526
rect 1738 -1534 1739 -1532
rect 1745 -1528 1746 -1526
rect 1745 -1534 1746 -1532
rect 1752 -1528 1753 -1526
rect 1752 -1534 1753 -1532
rect 1759 -1528 1760 -1526
rect 1759 -1534 1760 -1532
rect 1766 -1528 1767 -1526
rect 1766 -1534 1767 -1532
rect 1773 -1528 1774 -1526
rect 1773 -1534 1774 -1532
rect 1780 -1528 1781 -1526
rect 1780 -1534 1781 -1532
rect 1787 -1528 1788 -1526
rect 1787 -1534 1788 -1532
rect 1794 -1528 1795 -1526
rect 1797 -1528 1798 -1526
rect 1794 -1534 1795 -1532
rect 1801 -1528 1802 -1526
rect 1801 -1534 1802 -1532
rect 1808 -1528 1809 -1526
rect 1808 -1534 1809 -1532
rect 1815 -1528 1816 -1526
rect 1815 -1534 1816 -1532
rect 1822 -1528 1823 -1526
rect 1822 -1534 1823 -1532
rect 1829 -1528 1830 -1526
rect 1829 -1534 1830 -1532
rect 1836 -1528 1837 -1526
rect 1836 -1534 1837 -1532
rect 1843 -1528 1844 -1526
rect 1843 -1534 1844 -1532
rect 1850 -1528 1851 -1526
rect 1850 -1534 1851 -1532
rect 1857 -1528 1858 -1526
rect 1857 -1534 1858 -1532
rect 1864 -1528 1865 -1526
rect 1864 -1534 1865 -1532
rect 1871 -1528 1872 -1526
rect 1871 -1534 1872 -1532
rect 1878 -1528 1879 -1526
rect 1878 -1534 1879 -1532
rect 1885 -1528 1886 -1526
rect 1885 -1534 1886 -1532
rect 1892 -1528 1893 -1526
rect 1892 -1534 1893 -1532
rect 1899 -1528 1900 -1526
rect 1899 -1534 1900 -1532
rect 1906 -1528 1907 -1526
rect 1906 -1534 1907 -1532
rect 1913 -1528 1914 -1526
rect 1913 -1534 1914 -1532
rect 1920 -1528 1921 -1526
rect 1920 -1534 1921 -1532
rect 1927 -1528 1928 -1526
rect 1927 -1534 1928 -1532
rect 1934 -1528 1935 -1526
rect 1934 -1534 1935 -1532
rect 1941 -1528 1942 -1526
rect 1941 -1534 1942 -1532
rect 1948 -1528 1949 -1526
rect 1948 -1534 1949 -1532
rect 1955 -1528 1956 -1526
rect 1955 -1534 1956 -1532
rect 1962 -1528 1963 -1526
rect 1962 -1534 1963 -1532
rect 1969 -1528 1970 -1526
rect 1969 -1534 1970 -1532
rect 1976 -1528 1977 -1526
rect 1976 -1534 1977 -1532
rect 1983 -1528 1984 -1526
rect 1983 -1534 1984 -1532
rect 1990 -1528 1991 -1526
rect 1990 -1534 1991 -1532
rect 1997 -1528 1998 -1526
rect 1997 -1534 1998 -1532
rect 2004 -1528 2005 -1526
rect 2004 -1534 2005 -1532
rect 2011 -1528 2012 -1526
rect 2011 -1534 2012 -1532
rect 2018 -1528 2019 -1526
rect 2018 -1534 2019 -1532
rect 2025 -1528 2026 -1526
rect 2025 -1534 2026 -1532
rect 2032 -1528 2033 -1526
rect 2032 -1534 2033 -1532
rect 2039 -1528 2040 -1526
rect 2039 -1534 2040 -1532
rect 2046 -1528 2047 -1526
rect 2046 -1534 2047 -1532
rect 2053 -1528 2054 -1526
rect 2053 -1534 2054 -1532
rect 2060 -1528 2061 -1526
rect 2060 -1534 2061 -1532
rect 2067 -1528 2068 -1526
rect 2067 -1534 2068 -1532
rect 2074 -1528 2075 -1526
rect 2074 -1534 2075 -1532
rect 2081 -1528 2082 -1526
rect 2081 -1534 2082 -1532
rect 2088 -1528 2089 -1526
rect 2088 -1534 2089 -1532
rect 2095 -1528 2096 -1526
rect 2095 -1534 2096 -1532
rect 2102 -1528 2103 -1526
rect 2102 -1534 2103 -1532
rect 2109 -1528 2110 -1526
rect 2109 -1534 2110 -1532
rect 2116 -1528 2117 -1526
rect 2116 -1534 2117 -1532
rect 2123 -1528 2124 -1526
rect 2123 -1534 2124 -1532
rect 2130 -1528 2131 -1526
rect 2130 -1534 2131 -1532
rect 2137 -1528 2138 -1526
rect 2137 -1534 2138 -1532
rect 2144 -1528 2145 -1526
rect 2144 -1534 2145 -1532
rect 2151 -1528 2152 -1526
rect 2151 -1534 2152 -1532
rect 2158 -1528 2159 -1526
rect 2158 -1534 2159 -1532
rect 2165 -1528 2166 -1526
rect 2165 -1534 2166 -1532
rect 2172 -1528 2173 -1526
rect 2172 -1534 2173 -1532
rect 2179 -1528 2180 -1526
rect 2179 -1534 2180 -1532
rect 2186 -1528 2187 -1526
rect 2186 -1534 2187 -1532
rect 2193 -1528 2194 -1526
rect 2193 -1534 2194 -1532
rect 2200 -1528 2201 -1526
rect 2200 -1534 2201 -1532
rect 2207 -1528 2208 -1526
rect 2207 -1534 2208 -1532
rect 2214 -1528 2215 -1526
rect 2214 -1534 2215 -1532
rect 2221 -1528 2222 -1526
rect 2221 -1534 2222 -1532
rect 2228 -1528 2229 -1526
rect 2228 -1534 2229 -1532
rect 2235 -1528 2236 -1526
rect 2235 -1534 2236 -1532
rect 2242 -1528 2243 -1526
rect 2242 -1534 2243 -1532
rect 2249 -1528 2250 -1526
rect 2249 -1534 2250 -1532
rect 2256 -1528 2257 -1526
rect 2256 -1534 2257 -1532
rect 2263 -1528 2264 -1526
rect 2263 -1534 2264 -1532
rect 2270 -1528 2271 -1526
rect 2270 -1534 2271 -1532
rect 2277 -1528 2278 -1526
rect 2277 -1534 2278 -1532
rect 2284 -1528 2285 -1526
rect 2284 -1534 2285 -1532
rect 2291 -1528 2292 -1526
rect 2291 -1534 2292 -1532
rect 2298 -1528 2299 -1526
rect 2298 -1534 2299 -1532
rect 2305 -1528 2306 -1526
rect 2305 -1534 2306 -1532
rect 2312 -1528 2313 -1526
rect 2312 -1534 2313 -1532
rect 2319 -1528 2320 -1526
rect 2319 -1534 2320 -1532
rect 2326 -1528 2327 -1526
rect 2326 -1534 2327 -1532
rect 2333 -1528 2334 -1526
rect 2333 -1534 2334 -1532
rect 2340 -1528 2341 -1526
rect 2340 -1534 2341 -1532
rect 2347 -1528 2348 -1526
rect 2347 -1534 2348 -1532
rect 2354 -1528 2355 -1526
rect 2354 -1534 2355 -1532
rect 2361 -1528 2362 -1526
rect 2361 -1534 2362 -1532
rect 2368 -1528 2369 -1526
rect 2368 -1534 2369 -1532
rect 2375 -1528 2376 -1526
rect 2375 -1534 2376 -1532
rect 2382 -1528 2383 -1526
rect 2382 -1534 2383 -1532
rect 2389 -1528 2390 -1526
rect 2389 -1534 2390 -1532
rect 2396 -1528 2397 -1526
rect 2396 -1534 2397 -1532
rect 2403 -1528 2404 -1526
rect 2403 -1534 2404 -1532
rect 2410 -1528 2411 -1526
rect 2410 -1534 2411 -1532
rect 2417 -1528 2418 -1526
rect 2417 -1534 2418 -1532
rect 2424 -1528 2425 -1526
rect 2424 -1534 2425 -1532
rect 2431 -1528 2432 -1526
rect 2431 -1534 2432 -1532
rect 2438 -1528 2439 -1526
rect 2438 -1534 2439 -1532
rect 2445 -1528 2446 -1526
rect 2445 -1534 2446 -1532
rect 2452 -1528 2453 -1526
rect 2452 -1534 2453 -1532
rect 2459 -1528 2460 -1526
rect 2459 -1534 2460 -1532
rect 2466 -1528 2467 -1526
rect 2466 -1534 2467 -1532
rect 2473 -1528 2474 -1526
rect 2473 -1534 2474 -1532
rect 2480 -1528 2481 -1526
rect 2480 -1534 2481 -1532
rect 2487 -1528 2488 -1526
rect 2487 -1534 2488 -1532
rect 2494 -1528 2495 -1526
rect 2494 -1534 2495 -1532
rect 2501 -1528 2502 -1526
rect 2501 -1534 2502 -1532
rect 2508 -1528 2509 -1526
rect 2508 -1534 2509 -1532
rect 2515 -1528 2516 -1526
rect 2515 -1534 2516 -1532
rect 2522 -1528 2523 -1526
rect 2522 -1534 2523 -1532
rect 2529 -1528 2530 -1526
rect 2529 -1534 2530 -1532
rect 2536 -1528 2537 -1526
rect 2536 -1534 2537 -1532
rect 2543 -1528 2544 -1526
rect 2543 -1534 2544 -1532
rect 2550 -1528 2551 -1526
rect 2550 -1534 2551 -1532
rect 2557 -1528 2558 -1526
rect 2557 -1534 2558 -1532
rect 16 -1701 17 -1699
rect 16 -1707 17 -1705
rect 23 -1701 24 -1699
rect 23 -1707 24 -1705
rect 30 -1701 31 -1699
rect 30 -1707 31 -1705
rect 37 -1701 38 -1699
rect 37 -1707 38 -1705
rect 44 -1701 45 -1699
rect 44 -1707 45 -1705
rect 51 -1701 52 -1699
rect 51 -1707 52 -1705
rect 58 -1701 59 -1699
rect 58 -1707 59 -1705
rect 65 -1701 66 -1699
rect 65 -1707 66 -1705
rect 72 -1701 73 -1699
rect 72 -1707 73 -1705
rect 79 -1701 80 -1699
rect 79 -1707 80 -1705
rect 86 -1701 87 -1699
rect 86 -1707 87 -1705
rect 93 -1701 94 -1699
rect 96 -1701 97 -1699
rect 93 -1707 94 -1705
rect 96 -1707 97 -1705
rect 100 -1701 101 -1699
rect 100 -1707 101 -1705
rect 107 -1701 108 -1699
rect 107 -1707 108 -1705
rect 114 -1701 115 -1699
rect 114 -1707 115 -1705
rect 121 -1701 122 -1699
rect 121 -1707 122 -1705
rect 128 -1701 129 -1699
rect 128 -1707 129 -1705
rect 135 -1701 136 -1699
rect 135 -1707 136 -1705
rect 142 -1701 143 -1699
rect 142 -1707 143 -1705
rect 149 -1701 150 -1699
rect 149 -1707 150 -1705
rect 156 -1701 157 -1699
rect 156 -1707 157 -1705
rect 163 -1701 164 -1699
rect 163 -1707 164 -1705
rect 170 -1701 171 -1699
rect 170 -1707 171 -1705
rect 180 -1701 181 -1699
rect 177 -1707 178 -1705
rect 180 -1707 181 -1705
rect 184 -1701 185 -1699
rect 184 -1707 185 -1705
rect 191 -1701 192 -1699
rect 194 -1701 195 -1699
rect 191 -1707 192 -1705
rect 194 -1707 195 -1705
rect 198 -1701 199 -1699
rect 198 -1707 199 -1705
rect 205 -1701 206 -1699
rect 205 -1707 206 -1705
rect 212 -1701 213 -1699
rect 212 -1707 213 -1705
rect 215 -1707 216 -1705
rect 219 -1701 220 -1699
rect 219 -1707 220 -1705
rect 226 -1701 227 -1699
rect 229 -1701 230 -1699
rect 229 -1707 230 -1705
rect 233 -1701 234 -1699
rect 233 -1707 234 -1705
rect 240 -1701 241 -1699
rect 240 -1707 241 -1705
rect 250 -1701 251 -1699
rect 247 -1707 248 -1705
rect 254 -1701 255 -1699
rect 254 -1707 255 -1705
rect 261 -1701 262 -1699
rect 261 -1707 262 -1705
rect 268 -1701 269 -1699
rect 268 -1707 269 -1705
rect 275 -1701 276 -1699
rect 275 -1707 276 -1705
rect 282 -1701 283 -1699
rect 282 -1707 283 -1705
rect 289 -1701 290 -1699
rect 289 -1707 290 -1705
rect 296 -1701 297 -1699
rect 296 -1707 297 -1705
rect 303 -1701 304 -1699
rect 303 -1707 304 -1705
rect 310 -1701 311 -1699
rect 310 -1707 311 -1705
rect 317 -1701 318 -1699
rect 317 -1707 318 -1705
rect 324 -1701 325 -1699
rect 324 -1707 325 -1705
rect 331 -1701 332 -1699
rect 331 -1707 332 -1705
rect 338 -1701 339 -1699
rect 338 -1707 339 -1705
rect 345 -1701 346 -1699
rect 345 -1707 346 -1705
rect 352 -1701 353 -1699
rect 352 -1707 353 -1705
rect 359 -1701 360 -1699
rect 359 -1707 360 -1705
rect 366 -1701 367 -1699
rect 366 -1707 367 -1705
rect 373 -1701 374 -1699
rect 373 -1707 374 -1705
rect 380 -1701 381 -1699
rect 380 -1707 381 -1705
rect 387 -1701 388 -1699
rect 387 -1707 388 -1705
rect 394 -1701 395 -1699
rect 394 -1707 395 -1705
rect 401 -1701 402 -1699
rect 401 -1707 402 -1705
rect 408 -1701 409 -1699
rect 408 -1707 409 -1705
rect 415 -1701 416 -1699
rect 415 -1707 416 -1705
rect 422 -1701 423 -1699
rect 422 -1707 423 -1705
rect 429 -1701 430 -1699
rect 429 -1707 430 -1705
rect 436 -1701 437 -1699
rect 436 -1707 437 -1705
rect 443 -1701 444 -1699
rect 443 -1707 444 -1705
rect 450 -1701 451 -1699
rect 453 -1701 454 -1699
rect 453 -1707 454 -1705
rect 457 -1701 458 -1699
rect 460 -1701 461 -1699
rect 460 -1707 461 -1705
rect 464 -1701 465 -1699
rect 464 -1707 465 -1705
rect 471 -1701 472 -1699
rect 471 -1707 472 -1705
rect 478 -1701 479 -1699
rect 481 -1701 482 -1699
rect 478 -1707 479 -1705
rect 481 -1707 482 -1705
rect 485 -1701 486 -1699
rect 485 -1707 486 -1705
rect 492 -1701 493 -1699
rect 492 -1707 493 -1705
rect 499 -1701 500 -1699
rect 499 -1707 500 -1705
rect 506 -1701 507 -1699
rect 506 -1707 507 -1705
rect 513 -1701 514 -1699
rect 513 -1707 514 -1705
rect 520 -1701 521 -1699
rect 520 -1707 521 -1705
rect 527 -1701 528 -1699
rect 527 -1707 528 -1705
rect 534 -1701 535 -1699
rect 534 -1707 535 -1705
rect 541 -1701 542 -1699
rect 541 -1707 542 -1705
rect 548 -1701 549 -1699
rect 548 -1707 549 -1705
rect 555 -1701 556 -1699
rect 555 -1707 556 -1705
rect 562 -1701 563 -1699
rect 562 -1707 563 -1705
rect 569 -1701 570 -1699
rect 569 -1707 570 -1705
rect 576 -1707 577 -1705
rect 579 -1707 580 -1705
rect 583 -1701 584 -1699
rect 583 -1707 584 -1705
rect 590 -1701 591 -1699
rect 590 -1707 591 -1705
rect 597 -1701 598 -1699
rect 597 -1707 598 -1705
rect 604 -1701 605 -1699
rect 604 -1707 605 -1705
rect 611 -1701 612 -1699
rect 611 -1707 612 -1705
rect 618 -1701 619 -1699
rect 618 -1707 619 -1705
rect 625 -1701 626 -1699
rect 625 -1707 626 -1705
rect 632 -1701 633 -1699
rect 632 -1707 633 -1705
rect 639 -1701 640 -1699
rect 642 -1701 643 -1699
rect 642 -1707 643 -1705
rect 646 -1701 647 -1699
rect 646 -1707 647 -1705
rect 653 -1701 654 -1699
rect 653 -1707 654 -1705
rect 660 -1701 661 -1699
rect 660 -1707 661 -1705
rect 667 -1701 668 -1699
rect 667 -1707 668 -1705
rect 674 -1701 675 -1699
rect 674 -1707 675 -1705
rect 681 -1701 682 -1699
rect 681 -1707 682 -1705
rect 688 -1701 689 -1699
rect 688 -1707 689 -1705
rect 695 -1701 696 -1699
rect 698 -1701 699 -1699
rect 695 -1707 696 -1705
rect 698 -1707 699 -1705
rect 702 -1701 703 -1699
rect 702 -1707 703 -1705
rect 709 -1701 710 -1699
rect 709 -1707 710 -1705
rect 716 -1701 717 -1699
rect 719 -1701 720 -1699
rect 716 -1707 717 -1705
rect 719 -1707 720 -1705
rect 723 -1701 724 -1699
rect 723 -1707 724 -1705
rect 730 -1701 731 -1699
rect 730 -1707 731 -1705
rect 737 -1701 738 -1699
rect 737 -1707 738 -1705
rect 744 -1701 745 -1699
rect 744 -1707 745 -1705
rect 751 -1701 752 -1699
rect 751 -1707 752 -1705
rect 758 -1701 759 -1699
rect 758 -1707 759 -1705
rect 765 -1701 766 -1699
rect 765 -1707 766 -1705
rect 772 -1701 773 -1699
rect 772 -1707 773 -1705
rect 779 -1701 780 -1699
rect 779 -1707 780 -1705
rect 786 -1701 787 -1699
rect 786 -1707 787 -1705
rect 793 -1701 794 -1699
rect 793 -1707 794 -1705
rect 800 -1701 801 -1699
rect 800 -1707 801 -1705
rect 807 -1701 808 -1699
rect 807 -1707 808 -1705
rect 814 -1701 815 -1699
rect 814 -1707 815 -1705
rect 821 -1701 822 -1699
rect 821 -1707 822 -1705
rect 828 -1701 829 -1699
rect 828 -1707 829 -1705
rect 835 -1701 836 -1699
rect 835 -1707 836 -1705
rect 842 -1701 843 -1699
rect 842 -1707 843 -1705
rect 849 -1701 850 -1699
rect 849 -1707 850 -1705
rect 856 -1701 857 -1699
rect 859 -1701 860 -1699
rect 856 -1707 857 -1705
rect 859 -1707 860 -1705
rect 863 -1701 864 -1699
rect 863 -1707 864 -1705
rect 870 -1701 871 -1699
rect 870 -1707 871 -1705
rect 877 -1701 878 -1699
rect 877 -1707 878 -1705
rect 884 -1701 885 -1699
rect 884 -1707 885 -1705
rect 891 -1701 892 -1699
rect 891 -1707 892 -1705
rect 898 -1701 899 -1699
rect 898 -1707 899 -1705
rect 905 -1701 906 -1699
rect 905 -1707 906 -1705
rect 912 -1701 913 -1699
rect 912 -1707 913 -1705
rect 919 -1701 920 -1699
rect 919 -1707 920 -1705
rect 926 -1701 927 -1699
rect 926 -1707 927 -1705
rect 933 -1701 934 -1699
rect 936 -1701 937 -1699
rect 933 -1707 934 -1705
rect 936 -1707 937 -1705
rect 940 -1701 941 -1699
rect 940 -1707 941 -1705
rect 947 -1701 948 -1699
rect 947 -1707 948 -1705
rect 954 -1701 955 -1699
rect 954 -1707 955 -1705
rect 961 -1701 962 -1699
rect 961 -1707 962 -1705
rect 968 -1701 969 -1699
rect 968 -1707 969 -1705
rect 971 -1707 972 -1705
rect 975 -1701 976 -1699
rect 975 -1707 976 -1705
rect 982 -1701 983 -1699
rect 982 -1707 983 -1705
rect 989 -1701 990 -1699
rect 989 -1707 990 -1705
rect 996 -1701 997 -1699
rect 996 -1707 997 -1705
rect 1003 -1701 1004 -1699
rect 1003 -1707 1004 -1705
rect 1010 -1701 1011 -1699
rect 1010 -1707 1011 -1705
rect 1017 -1701 1018 -1699
rect 1020 -1701 1021 -1699
rect 1017 -1707 1018 -1705
rect 1020 -1707 1021 -1705
rect 1024 -1701 1025 -1699
rect 1024 -1707 1025 -1705
rect 1034 -1701 1035 -1699
rect 1031 -1707 1032 -1705
rect 1038 -1701 1039 -1699
rect 1038 -1707 1039 -1705
rect 1045 -1701 1046 -1699
rect 1045 -1707 1046 -1705
rect 1052 -1701 1053 -1699
rect 1052 -1707 1053 -1705
rect 1059 -1701 1060 -1699
rect 1059 -1707 1060 -1705
rect 1066 -1701 1067 -1699
rect 1066 -1707 1067 -1705
rect 1073 -1701 1074 -1699
rect 1076 -1701 1077 -1699
rect 1073 -1707 1074 -1705
rect 1076 -1707 1077 -1705
rect 1080 -1701 1081 -1699
rect 1080 -1707 1081 -1705
rect 1087 -1701 1088 -1699
rect 1087 -1707 1088 -1705
rect 1094 -1701 1095 -1699
rect 1094 -1707 1095 -1705
rect 1101 -1701 1102 -1699
rect 1101 -1707 1102 -1705
rect 1108 -1701 1109 -1699
rect 1111 -1701 1112 -1699
rect 1108 -1707 1109 -1705
rect 1111 -1707 1112 -1705
rect 1115 -1701 1116 -1699
rect 1115 -1707 1116 -1705
rect 1122 -1701 1123 -1699
rect 1122 -1707 1123 -1705
rect 1129 -1701 1130 -1699
rect 1129 -1707 1130 -1705
rect 1136 -1701 1137 -1699
rect 1136 -1707 1137 -1705
rect 1143 -1701 1144 -1699
rect 1143 -1707 1144 -1705
rect 1153 -1701 1154 -1699
rect 1150 -1707 1151 -1705
rect 1153 -1707 1154 -1705
rect 1157 -1701 1158 -1699
rect 1157 -1707 1158 -1705
rect 1164 -1701 1165 -1699
rect 1164 -1707 1165 -1705
rect 1171 -1701 1172 -1699
rect 1171 -1707 1172 -1705
rect 1178 -1701 1179 -1699
rect 1178 -1707 1179 -1705
rect 1185 -1701 1186 -1699
rect 1185 -1707 1186 -1705
rect 1192 -1701 1193 -1699
rect 1192 -1707 1193 -1705
rect 1199 -1701 1200 -1699
rect 1199 -1707 1200 -1705
rect 1206 -1701 1207 -1699
rect 1206 -1707 1207 -1705
rect 1213 -1701 1214 -1699
rect 1213 -1707 1214 -1705
rect 1220 -1701 1221 -1699
rect 1220 -1707 1221 -1705
rect 1227 -1701 1228 -1699
rect 1227 -1707 1228 -1705
rect 1234 -1701 1235 -1699
rect 1234 -1707 1235 -1705
rect 1241 -1701 1242 -1699
rect 1241 -1707 1242 -1705
rect 1248 -1701 1249 -1699
rect 1248 -1707 1249 -1705
rect 1255 -1701 1256 -1699
rect 1255 -1707 1256 -1705
rect 1262 -1701 1263 -1699
rect 1265 -1701 1266 -1699
rect 1262 -1707 1263 -1705
rect 1265 -1707 1266 -1705
rect 1269 -1701 1270 -1699
rect 1269 -1707 1270 -1705
rect 1276 -1701 1277 -1699
rect 1276 -1707 1277 -1705
rect 1279 -1707 1280 -1705
rect 1283 -1701 1284 -1699
rect 1283 -1707 1284 -1705
rect 1290 -1701 1291 -1699
rect 1293 -1701 1294 -1699
rect 1290 -1707 1291 -1705
rect 1293 -1707 1294 -1705
rect 1297 -1701 1298 -1699
rect 1297 -1707 1298 -1705
rect 1304 -1701 1305 -1699
rect 1304 -1707 1305 -1705
rect 1311 -1701 1312 -1699
rect 1311 -1707 1312 -1705
rect 1318 -1701 1319 -1699
rect 1318 -1707 1319 -1705
rect 1325 -1701 1326 -1699
rect 1325 -1707 1326 -1705
rect 1332 -1701 1333 -1699
rect 1332 -1707 1333 -1705
rect 1339 -1701 1340 -1699
rect 1339 -1707 1340 -1705
rect 1346 -1701 1347 -1699
rect 1346 -1707 1347 -1705
rect 1353 -1701 1354 -1699
rect 1353 -1707 1354 -1705
rect 1360 -1701 1361 -1699
rect 1363 -1701 1364 -1699
rect 1360 -1707 1361 -1705
rect 1363 -1707 1364 -1705
rect 1367 -1701 1368 -1699
rect 1367 -1707 1368 -1705
rect 1374 -1701 1375 -1699
rect 1374 -1707 1375 -1705
rect 1381 -1701 1382 -1699
rect 1381 -1707 1382 -1705
rect 1388 -1701 1389 -1699
rect 1388 -1707 1389 -1705
rect 1395 -1701 1396 -1699
rect 1395 -1707 1396 -1705
rect 1402 -1701 1403 -1699
rect 1402 -1707 1403 -1705
rect 1409 -1701 1410 -1699
rect 1409 -1707 1410 -1705
rect 1416 -1701 1417 -1699
rect 1416 -1707 1417 -1705
rect 1423 -1701 1424 -1699
rect 1423 -1707 1424 -1705
rect 1430 -1701 1431 -1699
rect 1430 -1707 1431 -1705
rect 1437 -1701 1438 -1699
rect 1440 -1701 1441 -1699
rect 1437 -1707 1438 -1705
rect 1440 -1707 1441 -1705
rect 1444 -1701 1445 -1699
rect 1444 -1707 1445 -1705
rect 1451 -1701 1452 -1699
rect 1451 -1707 1452 -1705
rect 1458 -1701 1459 -1699
rect 1458 -1707 1459 -1705
rect 1465 -1701 1466 -1699
rect 1468 -1701 1469 -1699
rect 1465 -1707 1466 -1705
rect 1468 -1707 1469 -1705
rect 1472 -1701 1473 -1699
rect 1472 -1707 1473 -1705
rect 1479 -1701 1480 -1699
rect 1479 -1707 1480 -1705
rect 1486 -1701 1487 -1699
rect 1486 -1707 1487 -1705
rect 1493 -1701 1494 -1699
rect 1496 -1701 1497 -1699
rect 1493 -1707 1494 -1705
rect 1496 -1707 1497 -1705
rect 1500 -1701 1501 -1699
rect 1500 -1707 1501 -1705
rect 1507 -1701 1508 -1699
rect 1510 -1701 1511 -1699
rect 1507 -1707 1508 -1705
rect 1510 -1707 1511 -1705
rect 1514 -1701 1515 -1699
rect 1514 -1707 1515 -1705
rect 1521 -1701 1522 -1699
rect 1521 -1707 1522 -1705
rect 1528 -1701 1529 -1699
rect 1531 -1701 1532 -1699
rect 1528 -1707 1529 -1705
rect 1531 -1707 1532 -1705
rect 1535 -1701 1536 -1699
rect 1538 -1701 1539 -1699
rect 1535 -1707 1536 -1705
rect 1538 -1707 1539 -1705
rect 1542 -1701 1543 -1699
rect 1542 -1707 1543 -1705
rect 1549 -1701 1550 -1699
rect 1549 -1707 1550 -1705
rect 1556 -1701 1557 -1699
rect 1556 -1707 1557 -1705
rect 1563 -1701 1564 -1699
rect 1563 -1707 1564 -1705
rect 1570 -1701 1571 -1699
rect 1570 -1707 1571 -1705
rect 1577 -1701 1578 -1699
rect 1577 -1707 1578 -1705
rect 1584 -1701 1585 -1699
rect 1584 -1707 1585 -1705
rect 1591 -1701 1592 -1699
rect 1591 -1707 1592 -1705
rect 1598 -1701 1599 -1699
rect 1598 -1707 1599 -1705
rect 1605 -1701 1606 -1699
rect 1605 -1707 1606 -1705
rect 1612 -1701 1613 -1699
rect 1612 -1707 1613 -1705
rect 1619 -1701 1620 -1699
rect 1619 -1707 1620 -1705
rect 1626 -1701 1627 -1699
rect 1626 -1707 1627 -1705
rect 1633 -1701 1634 -1699
rect 1633 -1707 1634 -1705
rect 1640 -1701 1641 -1699
rect 1640 -1707 1641 -1705
rect 1647 -1701 1648 -1699
rect 1647 -1707 1648 -1705
rect 1654 -1701 1655 -1699
rect 1654 -1707 1655 -1705
rect 1661 -1701 1662 -1699
rect 1661 -1707 1662 -1705
rect 1668 -1701 1669 -1699
rect 1668 -1707 1669 -1705
rect 1675 -1701 1676 -1699
rect 1675 -1707 1676 -1705
rect 1682 -1701 1683 -1699
rect 1682 -1707 1683 -1705
rect 1689 -1701 1690 -1699
rect 1689 -1707 1690 -1705
rect 1696 -1701 1697 -1699
rect 1696 -1707 1697 -1705
rect 1703 -1701 1704 -1699
rect 1706 -1707 1707 -1705
rect 1710 -1701 1711 -1699
rect 1710 -1707 1711 -1705
rect 1717 -1701 1718 -1699
rect 1717 -1707 1718 -1705
rect 1724 -1701 1725 -1699
rect 1724 -1707 1725 -1705
rect 1731 -1701 1732 -1699
rect 1731 -1707 1732 -1705
rect 1738 -1701 1739 -1699
rect 1738 -1707 1739 -1705
rect 1745 -1701 1746 -1699
rect 1745 -1707 1746 -1705
rect 1752 -1701 1753 -1699
rect 1752 -1707 1753 -1705
rect 1759 -1701 1760 -1699
rect 1759 -1707 1760 -1705
rect 1766 -1701 1767 -1699
rect 1766 -1707 1767 -1705
rect 1773 -1701 1774 -1699
rect 1773 -1707 1774 -1705
rect 1780 -1701 1781 -1699
rect 1780 -1707 1781 -1705
rect 1787 -1701 1788 -1699
rect 1787 -1707 1788 -1705
rect 1794 -1701 1795 -1699
rect 1794 -1707 1795 -1705
rect 1801 -1701 1802 -1699
rect 1801 -1707 1802 -1705
rect 1808 -1701 1809 -1699
rect 1811 -1701 1812 -1699
rect 1808 -1707 1809 -1705
rect 1811 -1707 1812 -1705
rect 1815 -1701 1816 -1699
rect 1815 -1707 1816 -1705
rect 1822 -1701 1823 -1699
rect 1822 -1707 1823 -1705
rect 1829 -1701 1830 -1699
rect 1829 -1707 1830 -1705
rect 1836 -1701 1837 -1699
rect 1836 -1707 1837 -1705
rect 1843 -1701 1844 -1699
rect 1843 -1707 1844 -1705
rect 1850 -1701 1851 -1699
rect 1850 -1707 1851 -1705
rect 1857 -1701 1858 -1699
rect 1857 -1707 1858 -1705
rect 1864 -1701 1865 -1699
rect 1864 -1707 1865 -1705
rect 1871 -1701 1872 -1699
rect 1871 -1707 1872 -1705
rect 1878 -1701 1879 -1699
rect 1878 -1707 1879 -1705
rect 1885 -1701 1886 -1699
rect 1885 -1707 1886 -1705
rect 1892 -1701 1893 -1699
rect 1892 -1707 1893 -1705
rect 1899 -1701 1900 -1699
rect 1899 -1707 1900 -1705
rect 1906 -1701 1907 -1699
rect 1906 -1707 1907 -1705
rect 1913 -1701 1914 -1699
rect 1913 -1707 1914 -1705
rect 1920 -1701 1921 -1699
rect 1920 -1707 1921 -1705
rect 1927 -1701 1928 -1699
rect 1927 -1707 1928 -1705
rect 1934 -1701 1935 -1699
rect 1934 -1707 1935 -1705
rect 1941 -1701 1942 -1699
rect 1941 -1707 1942 -1705
rect 1948 -1701 1949 -1699
rect 1948 -1707 1949 -1705
rect 1955 -1701 1956 -1699
rect 1955 -1707 1956 -1705
rect 1962 -1701 1963 -1699
rect 1962 -1707 1963 -1705
rect 1969 -1701 1970 -1699
rect 1969 -1707 1970 -1705
rect 1976 -1701 1977 -1699
rect 1976 -1707 1977 -1705
rect 1983 -1701 1984 -1699
rect 1983 -1707 1984 -1705
rect 1990 -1701 1991 -1699
rect 1990 -1707 1991 -1705
rect 1997 -1701 1998 -1699
rect 1997 -1707 1998 -1705
rect 2004 -1701 2005 -1699
rect 2004 -1707 2005 -1705
rect 2011 -1701 2012 -1699
rect 2011 -1707 2012 -1705
rect 2018 -1701 2019 -1699
rect 2018 -1707 2019 -1705
rect 2025 -1701 2026 -1699
rect 2025 -1707 2026 -1705
rect 2032 -1701 2033 -1699
rect 2032 -1707 2033 -1705
rect 2039 -1701 2040 -1699
rect 2039 -1707 2040 -1705
rect 2042 -1707 2043 -1705
rect 2046 -1701 2047 -1699
rect 2046 -1707 2047 -1705
rect 2053 -1701 2054 -1699
rect 2053 -1707 2054 -1705
rect 2060 -1701 2061 -1699
rect 2060 -1707 2061 -1705
rect 2067 -1701 2068 -1699
rect 2067 -1707 2068 -1705
rect 2074 -1701 2075 -1699
rect 2074 -1707 2075 -1705
rect 2081 -1701 2082 -1699
rect 2081 -1707 2082 -1705
rect 2088 -1701 2089 -1699
rect 2088 -1707 2089 -1705
rect 2095 -1701 2096 -1699
rect 2095 -1707 2096 -1705
rect 2102 -1701 2103 -1699
rect 2102 -1707 2103 -1705
rect 2109 -1701 2110 -1699
rect 2109 -1707 2110 -1705
rect 2116 -1701 2117 -1699
rect 2116 -1707 2117 -1705
rect 2123 -1701 2124 -1699
rect 2123 -1707 2124 -1705
rect 2130 -1701 2131 -1699
rect 2130 -1707 2131 -1705
rect 2137 -1701 2138 -1699
rect 2137 -1707 2138 -1705
rect 2144 -1701 2145 -1699
rect 2144 -1707 2145 -1705
rect 2151 -1701 2152 -1699
rect 2151 -1707 2152 -1705
rect 2158 -1701 2159 -1699
rect 2158 -1707 2159 -1705
rect 2165 -1701 2166 -1699
rect 2165 -1707 2166 -1705
rect 2172 -1701 2173 -1699
rect 2172 -1707 2173 -1705
rect 2179 -1701 2180 -1699
rect 2179 -1707 2180 -1705
rect 2186 -1701 2187 -1699
rect 2186 -1707 2187 -1705
rect 2193 -1701 2194 -1699
rect 2193 -1707 2194 -1705
rect 2200 -1701 2201 -1699
rect 2200 -1707 2201 -1705
rect 2207 -1701 2208 -1699
rect 2207 -1707 2208 -1705
rect 2214 -1701 2215 -1699
rect 2214 -1707 2215 -1705
rect 2221 -1701 2222 -1699
rect 2221 -1707 2222 -1705
rect 2228 -1701 2229 -1699
rect 2228 -1707 2229 -1705
rect 2235 -1701 2236 -1699
rect 2235 -1707 2236 -1705
rect 2242 -1701 2243 -1699
rect 2242 -1707 2243 -1705
rect 2249 -1701 2250 -1699
rect 2249 -1707 2250 -1705
rect 2256 -1701 2257 -1699
rect 2256 -1707 2257 -1705
rect 2263 -1701 2264 -1699
rect 2263 -1707 2264 -1705
rect 2270 -1701 2271 -1699
rect 2270 -1707 2271 -1705
rect 2277 -1701 2278 -1699
rect 2277 -1707 2278 -1705
rect 2284 -1701 2285 -1699
rect 2284 -1707 2285 -1705
rect 2291 -1701 2292 -1699
rect 2291 -1707 2292 -1705
rect 2298 -1701 2299 -1699
rect 2298 -1707 2299 -1705
rect 2305 -1701 2306 -1699
rect 2305 -1707 2306 -1705
rect 2312 -1701 2313 -1699
rect 2312 -1707 2313 -1705
rect 2319 -1701 2320 -1699
rect 2319 -1707 2320 -1705
rect 2326 -1701 2327 -1699
rect 2326 -1707 2327 -1705
rect 2333 -1701 2334 -1699
rect 2333 -1707 2334 -1705
rect 2340 -1701 2341 -1699
rect 2340 -1707 2341 -1705
rect 2347 -1701 2348 -1699
rect 2347 -1707 2348 -1705
rect 2354 -1701 2355 -1699
rect 2354 -1707 2355 -1705
rect 2361 -1701 2362 -1699
rect 2361 -1707 2362 -1705
rect 2368 -1701 2369 -1699
rect 2368 -1707 2369 -1705
rect 2375 -1701 2376 -1699
rect 2375 -1707 2376 -1705
rect 2382 -1701 2383 -1699
rect 2382 -1707 2383 -1705
rect 2389 -1701 2390 -1699
rect 2389 -1707 2390 -1705
rect 2396 -1701 2397 -1699
rect 2396 -1707 2397 -1705
rect 2403 -1701 2404 -1699
rect 2403 -1707 2404 -1705
rect 2410 -1701 2411 -1699
rect 2410 -1707 2411 -1705
rect 2417 -1701 2418 -1699
rect 2417 -1707 2418 -1705
rect 2424 -1701 2425 -1699
rect 2427 -1701 2428 -1699
rect 2424 -1707 2425 -1705
rect 2427 -1707 2428 -1705
rect 2434 -1701 2435 -1699
rect 2431 -1707 2432 -1705
rect 2434 -1707 2435 -1705
rect 2438 -1701 2439 -1699
rect 2441 -1701 2442 -1699
rect 2441 -1707 2442 -1705
rect 2445 -1701 2446 -1699
rect 2445 -1707 2446 -1705
rect 2452 -1701 2453 -1699
rect 2452 -1707 2453 -1705
rect 2494 -1701 2495 -1699
rect 2494 -1707 2495 -1705
rect 2 -1852 3 -1850
rect 2 -1858 3 -1856
rect 9 -1852 10 -1850
rect 9 -1858 10 -1856
rect 16 -1852 17 -1850
rect 16 -1858 17 -1856
rect 23 -1852 24 -1850
rect 23 -1858 24 -1856
rect 30 -1852 31 -1850
rect 30 -1858 31 -1856
rect 37 -1852 38 -1850
rect 37 -1858 38 -1856
rect 47 -1852 48 -1850
rect 44 -1858 45 -1856
rect 47 -1858 48 -1856
rect 51 -1852 52 -1850
rect 51 -1858 52 -1856
rect 58 -1852 59 -1850
rect 58 -1858 59 -1856
rect 65 -1852 66 -1850
rect 65 -1858 66 -1856
rect 72 -1852 73 -1850
rect 72 -1858 73 -1856
rect 79 -1852 80 -1850
rect 79 -1858 80 -1856
rect 86 -1852 87 -1850
rect 86 -1858 87 -1856
rect 93 -1852 94 -1850
rect 93 -1858 94 -1856
rect 100 -1852 101 -1850
rect 100 -1858 101 -1856
rect 107 -1852 108 -1850
rect 107 -1858 108 -1856
rect 114 -1852 115 -1850
rect 114 -1858 115 -1856
rect 121 -1852 122 -1850
rect 124 -1852 125 -1850
rect 121 -1858 122 -1856
rect 124 -1858 125 -1856
rect 128 -1852 129 -1850
rect 128 -1858 129 -1856
rect 135 -1852 136 -1850
rect 135 -1858 136 -1856
rect 142 -1852 143 -1850
rect 142 -1858 143 -1856
rect 149 -1852 150 -1850
rect 149 -1858 150 -1856
rect 159 -1852 160 -1850
rect 159 -1858 160 -1856
rect 163 -1852 164 -1850
rect 163 -1858 164 -1856
rect 170 -1852 171 -1850
rect 170 -1858 171 -1856
rect 177 -1852 178 -1850
rect 177 -1858 178 -1856
rect 184 -1852 185 -1850
rect 187 -1852 188 -1850
rect 184 -1858 185 -1856
rect 187 -1858 188 -1856
rect 191 -1852 192 -1850
rect 191 -1858 192 -1856
rect 198 -1852 199 -1850
rect 201 -1852 202 -1850
rect 198 -1858 199 -1856
rect 205 -1852 206 -1850
rect 205 -1858 206 -1856
rect 212 -1852 213 -1850
rect 212 -1858 213 -1856
rect 219 -1852 220 -1850
rect 219 -1858 220 -1856
rect 226 -1852 227 -1850
rect 226 -1858 227 -1856
rect 229 -1858 230 -1856
rect 233 -1852 234 -1850
rect 236 -1852 237 -1850
rect 233 -1858 234 -1856
rect 240 -1852 241 -1850
rect 240 -1858 241 -1856
rect 250 -1852 251 -1850
rect 247 -1858 248 -1856
rect 250 -1858 251 -1856
rect 254 -1852 255 -1850
rect 254 -1858 255 -1856
rect 261 -1852 262 -1850
rect 261 -1858 262 -1856
rect 268 -1852 269 -1850
rect 268 -1858 269 -1856
rect 275 -1852 276 -1850
rect 275 -1858 276 -1856
rect 282 -1852 283 -1850
rect 282 -1858 283 -1856
rect 289 -1852 290 -1850
rect 289 -1858 290 -1856
rect 296 -1852 297 -1850
rect 296 -1858 297 -1856
rect 303 -1852 304 -1850
rect 303 -1858 304 -1856
rect 310 -1852 311 -1850
rect 310 -1858 311 -1856
rect 317 -1852 318 -1850
rect 317 -1858 318 -1856
rect 324 -1852 325 -1850
rect 324 -1858 325 -1856
rect 331 -1852 332 -1850
rect 331 -1858 332 -1856
rect 338 -1852 339 -1850
rect 338 -1858 339 -1856
rect 345 -1852 346 -1850
rect 345 -1858 346 -1856
rect 352 -1852 353 -1850
rect 352 -1858 353 -1856
rect 359 -1852 360 -1850
rect 359 -1858 360 -1856
rect 366 -1852 367 -1850
rect 366 -1858 367 -1856
rect 373 -1852 374 -1850
rect 373 -1858 374 -1856
rect 380 -1852 381 -1850
rect 380 -1858 381 -1856
rect 387 -1852 388 -1850
rect 387 -1858 388 -1856
rect 394 -1852 395 -1850
rect 394 -1858 395 -1856
rect 401 -1852 402 -1850
rect 401 -1858 402 -1856
rect 408 -1852 409 -1850
rect 408 -1858 409 -1856
rect 415 -1852 416 -1850
rect 415 -1858 416 -1856
rect 422 -1852 423 -1850
rect 422 -1858 423 -1856
rect 429 -1852 430 -1850
rect 429 -1858 430 -1856
rect 432 -1858 433 -1856
rect 436 -1852 437 -1850
rect 436 -1858 437 -1856
rect 443 -1852 444 -1850
rect 446 -1852 447 -1850
rect 443 -1858 444 -1856
rect 446 -1858 447 -1856
rect 450 -1858 451 -1856
rect 457 -1852 458 -1850
rect 457 -1858 458 -1856
rect 464 -1852 465 -1850
rect 464 -1858 465 -1856
rect 471 -1852 472 -1850
rect 471 -1858 472 -1856
rect 478 -1852 479 -1850
rect 478 -1858 479 -1856
rect 485 -1852 486 -1850
rect 485 -1858 486 -1856
rect 492 -1852 493 -1850
rect 492 -1858 493 -1856
rect 499 -1852 500 -1850
rect 499 -1858 500 -1856
rect 506 -1852 507 -1850
rect 506 -1858 507 -1856
rect 513 -1852 514 -1850
rect 516 -1852 517 -1850
rect 513 -1858 514 -1856
rect 516 -1858 517 -1856
rect 520 -1852 521 -1850
rect 520 -1858 521 -1856
rect 527 -1852 528 -1850
rect 527 -1858 528 -1856
rect 534 -1852 535 -1850
rect 534 -1858 535 -1856
rect 541 -1852 542 -1850
rect 541 -1858 542 -1856
rect 548 -1852 549 -1850
rect 548 -1858 549 -1856
rect 555 -1852 556 -1850
rect 555 -1858 556 -1856
rect 562 -1852 563 -1850
rect 565 -1852 566 -1850
rect 562 -1858 563 -1856
rect 565 -1858 566 -1856
rect 569 -1852 570 -1850
rect 569 -1858 570 -1856
rect 576 -1852 577 -1850
rect 576 -1858 577 -1856
rect 583 -1852 584 -1850
rect 583 -1858 584 -1856
rect 590 -1852 591 -1850
rect 590 -1858 591 -1856
rect 597 -1852 598 -1850
rect 597 -1858 598 -1856
rect 604 -1852 605 -1850
rect 604 -1858 605 -1856
rect 611 -1852 612 -1850
rect 614 -1852 615 -1850
rect 611 -1858 612 -1856
rect 614 -1858 615 -1856
rect 618 -1852 619 -1850
rect 618 -1858 619 -1856
rect 625 -1852 626 -1850
rect 625 -1858 626 -1856
rect 632 -1858 633 -1856
rect 635 -1858 636 -1856
rect 639 -1852 640 -1850
rect 639 -1858 640 -1856
rect 646 -1852 647 -1850
rect 649 -1852 650 -1850
rect 646 -1858 647 -1856
rect 649 -1858 650 -1856
rect 653 -1852 654 -1850
rect 653 -1858 654 -1856
rect 660 -1852 661 -1850
rect 660 -1858 661 -1856
rect 667 -1852 668 -1850
rect 667 -1858 668 -1856
rect 674 -1852 675 -1850
rect 674 -1858 675 -1856
rect 681 -1852 682 -1850
rect 681 -1858 682 -1856
rect 688 -1852 689 -1850
rect 688 -1858 689 -1856
rect 695 -1852 696 -1850
rect 695 -1858 696 -1856
rect 702 -1852 703 -1850
rect 702 -1858 703 -1856
rect 709 -1852 710 -1850
rect 709 -1858 710 -1856
rect 716 -1852 717 -1850
rect 716 -1858 717 -1856
rect 723 -1852 724 -1850
rect 723 -1858 724 -1856
rect 726 -1858 727 -1856
rect 730 -1852 731 -1850
rect 733 -1852 734 -1850
rect 730 -1858 731 -1856
rect 737 -1852 738 -1850
rect 740 -1852 741 -1850
rect 737 -1858 738 -1856
rect 740 -1858 741 -1856
rect 744 -1852 745 -1850
rect 744 -1858 745 -1856
rect 751 -1852 752 -1850
rect 751 -1858 752 -1856
rect 758 -1852 759 -1850
rect 758 -1858 759 -1856
rect 765 -1852 766 -1850
rect 765 -1858 766 -1856
rect 772 -1852 773 -1850
rect 772 -1858 773 -1856
rect 779 -1852 780 -1850
rect 779 -1858 780 -1856
rect 786 -1852 787 -1850
rect 786 -1858 787 -1856
rect 793 -1852 794 -1850
rect 793 -1858 794 -1856
rect 800 -1852 801 -1850
rect 803 -1852 804 -1850
rect 800 -1858 801 -1856
rect 803 -1858 804 -1856
rect 807 -1852 808 -1850
rect 807 -1858 808 -1856
rect 814 -1852 815 -1850
rect 814 -1858 815 -1856
rect 821 -1852 822 -1850
rect 821 -1858 822 -1856
rect 828 -1852 829 -1850
rect 828 -1858 829 -1856
rect 835 -1852 836 -1850
rect 835 -1858 836 -1856
rect 842 -1852 843 -1850
rect 842 -1858 843 -1856
rect 849 -1858 850 -1856
rect 852 -1858 853 -1856
rect 856 -1852 857 -1850
rect 856 -1858 857 -1856
rect 863 -1852 864 -1850
rect 863 -1858 864 -1856
rect 870 -1852 871 -1850
rect 870 -1858 871 -1856
rect 877 -1852 878 -1850
rect 877 -1858 878 -1856
rect 884 -1852 885 -1850
rect 884 -1858 885 -1856
rect 891 -1852 892 -1850
rect 894 -1852 895 -1850
rect 891 -1858 892 -1856
rect 894 -1858 895 -1856
rect 898 -1852 899 -1850
rect 898 -1858 899 -1856
rect 905 -1852 906 -1850
rect 908 -1852 909 -1850
rect 908 -1858 909 -1856
rect 912 -1852 913 -1850
rect 912 -1858 913 -1856
rect 919 -1852 920 -1850
rect 919 -1858 920 -1856
rect 926 -1852 927 -1850
rect 926 -1858 927 -1856
rect 933 -1852 934 -1850
rect 933 -1858 934 -1856
rect 940 -1852 941 -1850
rect 943 -1852 944 -1850
rect 940 -1858 941 -1856
rect 943 -1858 944 -1856
rect 947 -1852 948 -1850
rect 947 -1858 948 -1856
rect 954 -1852 955 -1850
rect 957 -1852 958 -1850
rect 954 -1858 955 -1856
rect 957 -1858 958 -1856
rect 961 -1852 962 -1850
rect 961 -1858 962 -1856
rect 968 -1852 969 -1850
rect 968 -1858 969 -1856
rect 975 -1852 976 -1850
rect 975 -1858 976 -1856
rect 982 -1852 983 -1850
rect 982 -1858 983 -1856
rect 989 -1852 990 -1850
rect 989 -1858 990 -1856
rect 996 -1852 997 -1850
rect 996 -1858 997 -1856
rect 1003 -1852 1004 -1850
rect 1003 -1858 1004 -1856
rect 1010 -1852 1011 -1850
rect 1010 -1858 1011 -1856
rect 1017 -1852 1018 -1850
rect 1017 -1858 1018 -1856
rect 1024 -1852 1025 -1850
rect 1024 -1858 1025 -1856
rect 1031 -1852 1032 -1850
rect 1031 -1858 1032 -1856
rect 1038 -1852 1039 -1850
rect 1038 -1858 1039 -1856
rect 1045 -1852 1046 -1850
rect 1045 -1858 1046 -1856
rect 1052 -1852 1053 -1850
rect 1052 -1858 1053 -1856
rect 1059 -1852 1060 -1850
rect 1059 -1858 1060 -1856
rect 1066 -1852 1067 -1850
rect 1066 -1858 1067 -1856
rect 1073 -1852 1074 -1850
rect 1073 -1858 1074 -1856
rect 1080 -1852 1081 -1850
rect 1080 -1858 1081 -1856
rect 1087 -1852 1088 -1850
rect 1087 -1858 1088 -1856
rect 1094 -1852 1095 -1850
rect 1094 -1858 1095 -1856
rect 1101 -1852 1102 -1850
rect 1101 -1858 1102 -1856
rect 1108 -1852 1109 -1850
rect 1108 -1858 1109 -1856
rect 1115 -1852 1116 -1850
rect 1115 -1858 1116 -1856
rect 1122 -1852 1123 -1850
rect 1122 -1858 1123 -1856
rect 1129 -1852 1130 -1850
rect 1129 -1858 1130 -1856
rect 1136 -1852 1137 -1850
rect 1136 -1858 1137 -1856
rect 1139 -1858 1140 -1856
rect 1143 -1852 1144 -1850
rect 1143 -1858 1144 -1856
rect 1150 -1852 1151 -1850
rect 1150 -1858 1151 -1856
rect 1157 -1852 1158 -1850
rect 1157 -1858 1158 -1856
rect 1164 -1852 1165 -1850
rect 1164 -1858 1165 -1856
rect 1171 -1852 1172 -1850
rect 1171 -1858 1172 -1856
rect 1178 -1852 1179 -1850
rect 1181 -1852 1182 -1850
rect 1178 -1858 1179 -1856
rect 1181 -1858 1182 -1856
rect 1185 -1852 1186 -1850
rect 1185 -1858 1186 -1856
rect 1192 -1852 1193 -1850
rect 1192 -1858 1193 -1856
rect 1199 -1852 1200 -1850
rect 1199 -1858 1200 -1856
rect 1209 -1852 1210 -1850
rect 1206 -1858 1207 -1856
rect 1209 -1858 1210 -1856
rect 1213 -1852 1214 -1850
rect 1213 -1858 1214 -1856
rect 1220 -1852 1221 -1850
rect 1220 -1858 1221 -1856
rect 1227 -1852 1228 -1850
rect 1227 -1858 1228 -1856
rect 1234 -1852 1235 -1850
rect 1234 -1858 1235 -1856
rect 1241 -1852 1242 -1850
rect 1241 -1858 1242 -1856
rect 1248 -1852 1249 -1850
rect 1248 -1858 1249 -1856
rect 1255 -1852 1256 -1850
rect 1255 -1858 1256 -1856
rect 1262 -1852 1263 -1850
rect 1262 -1858 1263 -1856
rect 1269 -1852 1270 -1850
rect 1269 -1858 1270 -1856
rect 1276 -1852 1277 -1850
rect 1279 -1852 1280 -1850
rect 1276 -1858 1277 -1856
rect 1279 -1858 1280 -1856
rect 1283 -1852 1284 -1850
rect 1283 -1858 1284 -1856
rect 1290 -1852 1291 -1850
rect 1293 -1852 1294 -1850
rect 1290 -1858 1291 -1856
rect 1297 -1852 1298 -1850
rect 1297 -1858 1298 -1856
rect 1304 -1852 1305 -1850
rect 1307 -1852 1308 -1850
rect 1304 -1858 1305 -1856
rect 1307 -1858 1308 -1856
rect 1311 -1852 1312 -1850
rect 1311 -1858 1312 -1856
rect 1318 -1852 1319 -1850
rect 1318 -1858 1319 -1856
rect 1325 -1852 1326 -1850
rect 1332 -1852 1333 -1850
rect 1332 -1858 1333 -1856
rect 1335 -1858 1336 -1856
rect 1339 -1852 1340 -1850
rect 1339 -1858 1340 -1856
rect 1346 -1852 1347 -1850
rect 1346 -1858 1347 -1856
rect 1353 -1852 1354 -1850
rect 1353 -1858 1354 -1856
rect 1360 -1852 1361 -1850
rect 1360 -1858 1361 -1856
rect 1367 -1852 1368 -1850
rect 1367 -1858 1368 -1856
rect 1374 -1852 1375 -1850
rect 1374 -1858 1375 -1856
rect 1381 -1852 1382 -1850
rect 1381 -1858 1382 -1856
rect 1388 -1852 1389 -1850
rect 1388 -1858 1389 -1856
rect 1395 -1852 1396 -1850
rect 1395 -1858 1396 -1856
rect 1402 -1852 1403 -1850
rect 1402 -1858 1403 -1856
rect 1409 -1852 1410 -1850
rect 1409 -1858 1410 -1856
rect 1416 -1852 1417 -1850
rect 1416 -1858 1417 -1856
rect 1423 -1852 1424 -1850
rect 1423 -1858 1424 -1856
rect 1430 -1852 1431 -1850
rect 1430 -1858 1431 -1856
rect 1437 -1852 1438 -1850
rect 1440 -1852 1441 -1850
rect 1437 -1858 1438 -1856
rect 1440 -1858 1441 -1856
rect 1444 -1852 1445 -1850
rect 1444 -1858 1445 -1856
rect 1451 -1852 1452 -1850
rect 1451 -1858 1452 -1856
rect 1458 -1852 1459 -1850
rect 1458 -1858 1459 -1856
rect 1465 -1852 1466 -1850
rect 1468 -1852 1469 -1850
rect 1465 -1858 1466 -1856
rect 1468 -1858 1469 -1856
rect 1472 -1852 1473 -1850
rect 1472 -1858 1473 -1856
rect 1479 -1852 1480 -1850
rect 1479 -1858 1480 -1856
rect 1486 -1852 1487 -1850
rect 1486 -1858 1487 -1856
rect 1493 -1852 1494 -1850
rect 1493 -1858 1494 -1856
rect 1500 -1852 1501 -1850
rect 1500 -1858 1501 -1856
rect 1507 -1852 1508 -1850
rect 1507 -1858 1508 -1856
rect 1510 -1858 1511 -1856
rect 1514 -1852 1515 -1850
rect 1514 -1858 1515 -1856
rect 1521 -1852 1522 -1850
rect 1521 -1858 1522 -1856
rect 1528 -1852 1529 -1850
rect 1528 -1858 1529 -1856
rect 1535 -1852 1536 -1850
rect 1535 -1858 1536 -1856
rect 1542 -1852 1543 -1850
rect 1542 -1858 1543 -1856
rect 1549 -1852 1550 -1850
rect 1549 -1858 1550 -1856
rect 1556 -1852 1557 -1850
rect 1556 -1858 1557 -1856
rect 1563 -1852 1564 -1850
rect 1563 -1858 1564 -1856
rect 1570 -1852 1571 -1850
rect 1570 -1858 1571 -1856
rect 1577 -1852 1578 -1850
rect 1577 -1858 1578 -1856
rect 1584 -1852 1585 -1850
rect 1584 -1858 1585 -1856
rect 1591 -1852 1592 -1850
rect 1591 -1858 1592 -1856
rect 1598 -1852 1599 -1850
rect 1598 -1858 1599 -1856
rect 1605 -1852 1606 -1850
rect 1605 -1858 1606 -1856
rect 1612 -1852 1613 -1850
rect 1612 -1858 1613 -1856
rect 1619 -1852 1620 -1850
rect 1619 -1858 1620 -1856
rect 1626 -1852 1627 -1850
rect 1629 -1852 1630 -1850
rect 1629 -1858 1630 -1856
rect 1633 -1852 1634 -1850
rect 1633 -1858 1634 -1856
rect 1640 -1852 1641 -1850
rect 1640 -1858 1641 -1856
rect 1647 -1852 1648 -1850
rect 1647 -1858 1648 -1856
rect 1654 -1852 1655 -1850
rect 1654 -1858 1655 -1856
rect 1664 -1852 1665 -1850
rect 1661 -1858 1662 -1856
rect 1664 -1858 1665 -1856
rect 1668 -1852 1669 -1850
rect 1668 -1858 1669 -1856
rect 1675 -1852 1676 -1850
rect 1675 -1858 1676 -1856
rect 1682 -1852 1683 -1850
rect 1682 -1858 1683 -1856
rect 1689 -1852 1690 -1850
rect 1689 -1858 1690 -1856
rect 1696 -1852 1697 -1850
rect 1696 -1858 1697 -1856
rect 1703 -1852 1704 -1850
rect 1703 -1858 1704 -1856
rect 1710 -1852 1711 -1850
rect 1710 -1858 1711 -1856
rect 1717 -1852 1718 -1850
rect 1717 -1858 1718 -1856
rect 1724 -1852 1725 -1850
rect 1724 -1858 1725 -1856
rect 1731 -1852 1732 -1850
rect 1731 -1858 1732 -1856
rect 1738 -1852 1739 -1850
rect 1738 -1858 1739 -1856
rect 1745 -1852 1746 -1850
rect 1745 -1858 1746 -1856
rect 1752 -1852 1753 -1850
rect 1752 -1858 1753 -1856
rect 1759 -1852 1760 -1850
rect 1759 -1858 1760 -1856
rect 1766 -1852 1767 -1850
rect 1766 -1858 1767 -1856
rect 1773 -1852 1774 -1850
rect 1773 -1858 1774 -1856
rect 1780 -1852 1781 -1850
rect 1780 -1858 1781 -1856
rect 1787 -1852 1788 -1850
rect 1787 -1858 1788 -1856
rect 1794 -1852 1795 -1850
rect 1794 -1858 1795 -1856
rect 1801 -1852 1802 -1850
rect 1801 -1858 1802 -1856
rect 1808 -1852 1809 -1850
rect 1808 -1858 1809 -1856
rect 1815 -1852 1816 -1850
rect 1815 -1858 1816 -1856
rect 1822 -1852 1823 -1850
rect 1822 -1858 1823 -1856
rect 1829 -1852 1830 -1850
rect 1829 -1858 1830 -1856
rect 1836 -1852 1837 -1850
rect 1836 -1858 1837 -1856
rect 1843 -1852 1844 -1850
rect 1843 -1858 1844 -1856
rect 1850 -1852 1851 -1850
rect 1853 -1852 1854 -1850
rect 1850 -1858 1851 -1856
rect 1853 -1858 1854 -1856
rect 1857 -1852 1858 -1850
rect 1857 -1858 1858 -1856
rect 1864 -1858 1865 -1856
rect 1867 -1858 1868 -1856
rect 1871 -1852 1872 -1850
rect 1871 -1858 1872 -1856
rect 1878 -1852 1879 -1850
rect 1878 -1858 1879 -1856
rect 1885 -1852 1886 -1850
rect 1885 -1858 1886 -1856
rect 1892 -1852 1893 -1850
rect 1892 -1858 1893 -1856
rect 1899 -1852 1900 -1850
rect 1899 -1858 1900 -1856
rect 1906 -1852 1907 -1850
rect 1906 -1858 1907 -1856
rect 1913 -1852 1914 -1850
rect 1913 -1858 1914 -1856
rect 1920 -1852 1921 -1850
rect 1920 -1858 1921 -1856
rect 1927 -1852 1928 -1850
rect 1927 -1858 1928 -1856
rect 1934 -1852 1935 -1850
rect 1934 -1858 1935 -1856
rect 1941 -1852 1942 -1850
rect 1941 -1858 1942 -1856
rect 1948 -1852 1949 -1850
rect 1948 -1858 1949 -1856
rect 1955 -1852 1956 -1850
rect 1955 -1858 1956 -1856
rect 1962 -1852 1963 -1850
rect 1962 -1858 1963 -1856
rect 1969 -1852 1970 -1850
rect 1969 -1858 1970 -1856
rect 1976 -1852 1977 -1850
rect 1976 -1858 1977 -1856
rect 1983 -1852 1984 -1850
rect 1983 -1858 1984 -1856
rect 1990 -1852 1991 -1850
rect 1990 -1858 1991 -1856
rect 1997 -1852 1998 -1850
rect 1997 -1858 1998 -1856
rect 2004 -1852 2005 -1850
rect 2004 -1858 2005 -1856
rect 2011 -1852 2012 -1850
rect 2011 -1858 2012 -1856
rect 2018 -1852 2019 -1850
rect 2018 -1858 2019 -1856
rect 2025 -1852 2026 -1850
rect 2025 -1858 2026 -1856
rect 2032 -1852 2033 -1850
rect 2032 -1858 2033 -1856
rect 2039 -1852 2040 -1850
rect 2042 -1852 2043 -1850
rect 2039 -1858 2040 -1856
rect 2046 -1852 2047 -1850
rect 2046 -1858 2047 -1856
rect 2053 -1852 2054 -1850
rect 2053 -1858 2054 -1856
rect 2060 -1852 2061 -1850
rect 2060 -1858 2061 -1856
rect 2067 -1852 2068 -1850
rect 2067 -1858 2068 -1856
rect 2074 -1852 2075 -1850
rect 2074 -1858 2075 -1856
rect 2081 -1852 2082 -1850
rect 2081 -1858 2082 -1856
rect 2088 -1852 2089 -1850
rect 2088 -1858 2089 -1856
rect 2095 -1852 2096 -1850
rect 2095 -1858 2096 -1856
rect 2102 -1852 2103 -1850
rect 2102 -1858 2103 -1856
rect 2109 -1852 2110 -1850
rect 2109 -1858 2110 -1856
rect 2116 -1852 2117 -1850
rect 2116 -1858 2117 -1856
rect 2123 -1852 2124 -1850
rect 2123 -1858 2124 -1856
rect 2130 -1852 2131 -1850
rect 2130 -1858 2131 -1856
rect 2137 -1852 2138 -1850
rect 2137 -1858 2138 -1856
rect 2144 -1852 2145 -1850
rect 2144 -1858 2145 -1856
rect 2151 -1852 2152 -1850
rect 2151 -1858 2152 -1856
rect 2158 -1852 2159 -1850
rect 2158 -1858 2159 -1856
rect 2165 -1852 2166 -1850
rect 2165 -1858 2166 -1856
rect 2172 -1852 2173 -1850
rect 2172 -1858 2173 -1856
rect 2179 -1852 2180 -1850
rect 2179 -1858 2180 -1856
rect 2186 -1852 2187 -1850
rect 2186 -1858 2187 -1856
rect 2193 -1852 2194 -1850
rect 2193 -1858 2194 -1856
rect 2200 -1852 2201 -1850
rect 2200 -1858 2201 -1856
rect 2207 -1852 2208 -1850
rect 2207 -1858 2208 -1856
rect 2214 -1852 2215 -1850
rect 2214 -1858 2215 -1856
rect 2221 -1852 2222 -1850
rect 2221 -1858 2222 -1856
rect 2228 -1852 2229 -1850
rect 2228 -1858 2229 -1856
rect 2235 -1852 2236 -1850
rect 2235 -1858 2236 -1856
rect 2242 -1852 2243 -1850
rect 2242 -1858 2243 -1856
rect 2249 -1852 2250 -1850
rect 2249 -1858 2250 -1856
rect 2256 -1852 2257 -1850
rect 2256 -1858 2257 -1856
rect 2263 -1852 2264 -1850
rect 2263 -1858 2264 -1856
rect 2270 -1852 2271 -1850
rect 2270 -1858 2271 -1856
rect 2277 -1852 2278 -1850
rect 2277 -1858 2278 -1856
rect 2284 -1852 2285 -1850
rect 2284 -1858 2285 -1856
rect 2291 -1852 2292 -1850
rect 2291 -1858 2292 -1856
rect 2298 -1852 2299 -1850
rect 2298 -1858 2299 -1856
rect 2305 -1852 2306 -1850
rect 2305 -1858 2306 -1856
rect 2312 -1852 2313 -1850
rect 2312 -1858 2313 -1856
rect 2319 -1852 2320 -1850
rect 2319 -1858 2320 -1856
rect 2326 -1852 2327 -1850
rect 2326 -1858 2327 -1856
rect 2333 -1852 2334 -1850
rect 2333 -1858 2334 -1856
rect 2340 -1852 2341 -1850
rect 2340 -1858 2341 -1856
rect 2347 -1852 2348 -1850
rect 2347 -1858 2348 -1856
rect 2354 -1852 2355 -1850
rect 2354 -1858 2355 -1856
rect 2361 -1852 2362 -1850
rect 2361 -1858 2362 -1856
rect 2368 -1852 2369 -1850
rect 2368 -1858 2369 -1856
rect 2375 -1852 2376 -1850
rect 2375 -1858 2376 -1856
rect 2382 -1852 2383 -1850
rect 2382 -1858 2383 -1856
rect 2389 -1852 2390 -1850
rect 2389 -1858 2390 -1856
rect 2396 -1852 2397 -1850
rect 2396 -1858 2397 -1856
rect 2403 -1852 2404 -1850
rect 2403 -1858 2404 -1856
rect 2410 -1852 2411 -1850
rect 2410 -1858 2411 -1856
rect 2417 -1852 2418 -1850
rect 2417 -1858 2418 -1856
rect 2424 -1852 2425 -1850
rect 2424 -1858 2425 -1856
rect 2431 -1852 2432 -1850
rect 2431 -1858 2432 -1856
rect 2438 -1852 2439 -1850
rect 2438 -1858 2439 -1856
rect 2445 -1852 2446 -1850
rect 2445 -1858 2446 -1856
rect 2452 -1852 2453 -1850
rect 2452 -1858 2453 -1856
rect 2459 -1852 2460 -1850
rect 2459 -1858 2460 -1856
rect 2466 -1852 2467 -1850
rect 2469 -1852 2470 -1850
rect 2466 -1858 2467 -1856
rect 2469 -1858 2470 -1856
rect 2473 -1852 2474 -1850
rect 2476 -1852 2477 -1850
rect 2473 -1858 2474 -1856
rect 2 -2027 3 -2025
rect 2 -2033 3 -2031
rect 9 -2027 10 -2025
rect 9 -2033 10 -2031
rect 16 -2027 17 -2025
rect 16 -2033 17 -2031
rect 23 -2027 24 -2025
rect 23 -2033 24 -2031
rect 30 -2027 31 -2025
rect 30 -2033 31 -2031
rect 37 -2027 38 -2025
rect 37 -2033 38 -2031
rect 44 -2027 45 -2025
rect 44 -2033 45 -2031
rect 51 -2027 52 -2025
rect 51 -2033 52 -2031
rect 54 -2033 55 -2031
rect 58 -2027 59 -2025
rect 58 -2033 59 -2031
rect 65 -2027 66 -2025
rect 65 -2033 66 -2031
rect 72 -2027 73 -2025
rect 72 -2033 73 -2031
rect 79 -2027 80 -2025
rect 79 -2033 80 -2031
rect 86 -2027 87 -2025
rect 89 -2027 90 -2025
rect 89 -2033 90 -2031
rect 93 -2027 94 -2025
rect 93 -2033 94 -2031
rect 100 -2027 101 -2025
rect 103 -2027 104 -2025
rect 100 -2033 101 -2031
rect 103 -2033 104 -2031
rect 107 -2027 108 -2025
rect 107 -2033 108 -2031
rect 114 -2027 115 -2025
rect 114 -2033 115 -2031
rect 121 -2027 122 -2025
rect 121 -2033 122 -2031
rect 128 -2027 129 -2025
rect 131 -2027 132 -2025
rect 131 -2033 132 -2031
rect 135 -2027 136 -2025
rect 135 -2033 136 -2031
rect 142 -2027 143 -2025
rect 142 -2033 143 -2031
rect 149 -2027 150 -2025
rect 149 -2033 150 -2031
rect 156 -2027 157 -2025
rect 159 -2027 160 -2025
rect 156 -2033 157 -2031
rect 159 -2033 160 -2031
rect 163 -2027 164 -2025
rect 163 -2033 164 -2031
rect 170 -2027 171 -2025
rect 173 -2027 174 -2025
rect 170 -2033 171 -2031
rect 173 -2033 174 -2031
rect 177 -2027 178 -2025
rect 177 -2033 178 -2031
rect 184 -2027 185 -2025
rect 184 -2033 185 -2031
rect 191 -2027 192 -2025
rect 194 -2027 195 -2025
rect 191 -2033 192 -2031
rect 194 -2033 195 -2031
rect 198 -2027 199 -2025
rect 198 -2033 199 -2031
rect 205 -2027 206 -2025
rect 205 -2033 206 -2031
rect 212 -2027 213 -2025
rect 215 -2027 216 -2025
rect 212 -2033 213 -2031
rect 215 -2033 216 -2031
rect 219 -2027 220 -2025
rect 219 -2033 220 -2031
rect 226 -2027 227 -2025
rect 226 -2033 227 -2031
rect 233 -2027 234 -2025
rect 233 -2033 234 -2031
rect 240 -2027 241 -2025
rect 240 -2033 241 -2031
rect 247 -2027 248 -2025
rect 247 -2033 248 -2031
rect 254 -2027 255 -2025
rect 254 -2033 255 -2031
rect 261 -2027 262 -2025
rect 261 -2033 262 -2031
rect 268 -2027 269 -2025
rect 268 -2033 269 -2031
rect 275 -2027 276 -2025
rect 275 -2033 276 -2031
rect 282 -2027 283 -2025
rect 282 -2033 283 -2031
rect 289 -2027 290 -2025
rect 289 -2033 290 -2031
rect 296 -2027 297 -2025
rect 296 -2033 297 -2031
rect 303 -2027 304 -2025
rect 303 -2033 304 -2031
rect 310 -2027 311 -2025
rect 310 -2033 311 -2031
rect 317 -2027 318 -2025
rect 317 -2033 318 -2031
rect 324 -2027 325 -2025
rect 324 -2033 325 -2031
rect 331 -2027 332 -2025
rect 331 -2033 332 -2031
rect 338 -2027 339 -2025
rect 338 -2033 339 -2031
rect 345 -2027 346 -2025
rect 345 -2033 346 -2031
rect 352 -2027 353 -2025
rect 352 -2033 353 -2031
rect 359 -2027 360 -2025
rect 359 -2033 360 -2031
rect 366 -2027 367 -2025
rect 366 -2033 367 -2031
rect 373 -2027 374 -2025
rect 373 -2033 374 -2031
rect 380 -2027 381 -2025
rect 380 -2033 381 -2031
rect 387 -2027 388 -2025
rect 387 -2033 388 -2031
rect 394 -2027 395 -2025
rect 394 -2033 395 -2031
rect 401 -2027 402 -2025
rect 401 -2033 402 -2031
rect 408 -2027 409 -2025
rect 408 -2033 409 -2031
rect 415 -2027 416 -2025
rect 415 -2033 416 -2031
rect 422 -2027 423 -2025
rect 422 -2033 423 -2031
rect 429 -2027 430 -2025
rect 429 -2033 430 -2031
rect 436 -2027 437 -2025
rect 436 -2033 437 -2031
rect 443 -2027 444 -2025
rect 443 -2033 444 -2031
rect 450 -2027 451 -2025
rect 450 -2033 451 -2031
rect 457 -2027 458 -2025
rect 457 -2033 458 -2031
rect 464 -2027 465 -2025
rect 464 -2033 465 -2031
rect 471 -2027 472 -2025
rect 471 -2033 472 -2031
rect 478 -2027 479 -2025
rect 478 -2033 479 -2031
rect 485 -2027 486 -2025
rect 485 -2033 486 -2031
rect 492 -2027 493 -2025
rect 492 -2033 493 -2031
rect 499 -2027 500 -2025
rect 499 -2033 500 -2031
rect 506 -2027 507 -2025
rect 506 -2033 507 -2031
rect 513 -2027 514 -2025
rect 513 -2033 514 -2031
rect 520 -2027 521 -2025
rect 520 -2033 521 -2031
rect 527 -2027 528 -2025
rect 527 -2033 528 -2031
rect 534 -2027 535 -2025
rect 534 -2033 535 -2031
rect 541 -2027 542 -2025
rect 544 -2027 545 -2025
rect 548 -2027 549 -2025
rect 548 -2033 549 -2031
rect 555 -2027 556 -2025
rect 555 -2033 556 -2031
rect 562 -2027 563 -2025
rect 562 -2033 563 -2031
rect 569 -2027 570 -2025
rect 569 -2033 570 -2031
rect 576 -2027 577 -2025
rect 576 -2033 577 -2031
rect 583 -2027 584 -2025
rect 586 -2027 587 -2025
rect 586 -2033 587 -2031
rect 590 -2027 591 -2025
rect 590 -2033 591 -2031
rect 597 -2027 598 -2025
rect 597 -2033 598 -2031
rect 604 -2027 605 -2025
rect 604 -2033 605 -2031
rect 611 -2027 612 -2025
rect 611 -2033 612 -2031
rect 618 -2027 619 -2025
rect 618 -2033 619 -2031
rect 625 -2027 626 -2025
rect 625 -2033 626 -2031
rect 632 -2027 633 -2025
rect 635 -2027 636 -2025
rect 632 -2033 633 -2031
rect 639 -2027 640 -2025
rect 639 -2033 640 -2031
rect 646 -2027 647 -2025
rect 646 -2033 647 -2031
rect 653 -2027 654 -2025
rect 653 -2033 654 -2031
rect 660 -2027 661 -2025
rect 660 -2033 661 -2031
rect 667 -2027 668 -2025
rect 667 -2033 668 -2031
rect 674 -2027 675 -2025
rect 674 -2033 675 -2031
rect 681 -2027 682 -2025
rect 681 -2033 682 -2031
rect 688 -2027 689 -2025
rect 688 -2033 689 -2031
rect 695 -2027 696 -2025
rect 695 -2033 696 -2031
rect 702 -2027 703 -2025
rect 702 -2033 703 -2031
rect 709 -2027 710 -2025
rect 709 -2033 710 -2031
rect 716 -2027 717 -2025
rect 716 -2033 717 -2031
rect 723 -2027 724 -2025
rect 723 -2033 724 -2031
rect 730 -2027 731 -2025
rect 730 -2033 731 -2031
rect 737 -2027 738 -2025
rect 740 -2027 741 -2025
rect 737 -2033 738 -2031
rect 740 -2033 741 -2031
rect 744 -2027 745 -2025
rect 744 -2033 745 -2031
rect 751 -2027 752 -2025
rect 751 -2033 752 -2031
rect 758 -2027 759 -2025
rect 758 -2033 759 -2031
rect 765 -2027 766 -2025
rect 765 -2033 766 -2031
rect 772 -2027 773 -2025
rect 772 -2033 773 -2031
rect 779 -2027 780 -2025
rect 782 -2027 783 -2025
rect 779 -2033 780 -2031
rect 786 -2027 787 -2025
rect 786 -2033 787 -2031
rect 793 -2027 794 -2025
rect 793 -2033 794 -2031
rect 800 -2033 801 -2031
rect 803 -2033 804 -2031
rect 807 -2027 808 -2025
rect 807 -2033 808 -2031
rect 814 -2027 815 -2025
rect 814 -2033 815 -2031
rect 821 -2027 822 -2025
rect 821 -2033 822 -2031
rect 828 -2027 829 -2025
rect 831 -2027 832 -2025
rect 828 -2033 829 -2031
rect 831 -2033 832 -2031
rect 835 -2027 836 -2025
rect 835 -2033 836 -2031
rect 842 -2027 843 -2025
rect 842 -2033 843 -2031
rect 849 -2027 850 -2025
rect 849 -2033 850 -2031
rect 856 -2027 857 -2025
rect 856 -2033 857 -2031
rect 863 -2027 864 -2025
rect 863 -2033 864 -2031
rect 870 -2027 871 -2025
rect 870 -2033 871 -2031
rect 877 -2027 878 -2025
rect 877 -2033 878 -2031
rect 884 -2027 885 -2025
rect 884 -2033 885 -2031
rect 891 -2027 892 -2025
rect 891 -2033 892 -2031
rect 898 -2027 899 -2025
rect 898 -2033 899 -2031
rect 905 -2027 906 -2025
rect 905 -2033 906 -2031
rect 912 -2027 913 -2025
rect 912 -2033 913 -2031
rect 919 -2027 920 -2025
rect 922 -2027 923 -2025
rect 919 -2033 920 -2031
rect 922 -2033 923 -2031
rect 926 -2027 927 -2025
rect 926 -2033 927 -2031
rect 933 -2027 934 -2025
rect 933 -2033 934 -2031
rect 940 -2027 941 -2025
rect 940 -2033 941 -2031
rect 947 -2027 948 -2025
rect 947 -2033 948 -2031
rect 954 -2027 955 -2025
rect 957 -2027 958 -2025
rect 954 -2033 955 -2031
rect 957 -2033 958 -2031
rect 961 -2027 962 -2025
rect 961 -2033 962 -2031
rect 968 -2027 969 -2025
rect 968 -2033 969 -2031
rect 975 -2027 976 -2025
rect 978 -2027 979 -2025
rect 978 -2033 979 -2031
rect 982 -2027 983 -2025
rect 982 -2033 983 -2031
rect 989 -2027 990 -2025
rect 989 -2033 990 -2031
rect 996 -2027 997 -2025
rect 996 -2033 997 -2031
rect 1003 -2027 1004 -2025
rect 1003 -2033 1004 -2031
rect 1010 -2027 1011 -2025
rect 1010 -2033 1011 -2031
rect 1017 -2027 1018 -2025
rect 1017 -2033 1018 -2031
rect 1024 -2027 1025 -2025
rect 1024 -2033 1025 -2031
rect 1031 -2027 1032 -2025
rect 1031 -2033 1032 -2031
rect 1038 -2027 1039 -2025
rect 1038 -2033 1039 -2031
rect 1045 -2027 1046 -2025
rect 1045 -2033 1046 -2031
rect 1052 -2027 1053 -2025
rect 1052 -2033 1053 -2031
rect 1059 -2027 1060 -2025
rect 1062 -2027 1063 -2025
rect 1059 -2033 1060 -2031
rect 1062 -2033 1063 -2031
rect 1066 -2027 1067 -2025
rect 1066 -2033 1067 -2031
rect 1073 -2027 1074 -2025
rect 1073 -2033 1074 -2031
rect 1080 -2027 1081 -2025
rect 1080 -2033 1081 -2031
rect 1087 -2027 1088 -2025
rect 1087 -2033 1088 -2031
rect 1094 -2027 1095 -2025
rect 1094 -2033 1095 -2031
rect 1101 -2027 1102 -2025
rect 1101 -2033 1102 -2031
rect 1108 -2027 1109 -2025
rect 1111 -2027 1112 -2025
rect 1108 -2033 1109 -2031
rect 1111 -2033 1112 -2031
rect 1115 -2027 1116 -2025
rect 1115 -2033 1116 -2031
rect 1125 -2027 1126 -2025
rect 1122 -2033 1123 -2031
rect 1125 -2033 1126 -2031
rect 1129 -2027 1130 -2025
rect 1129 -2033 1130 -2031
rect 1136 -2027 1137 -2025
rect 1136 -2033 1137 -2031
rect 1143 -2027 1144 -2025
rect 1143 -2033 1144 -2031
rect 1153 -2027 1154 -2025
rect 1153 -2033 1154 -2031
rect 1157 -2027 1158 -2025
rect 1157 -2033 1158 -2031
rect 1164 -2027 1165 -2025
rect 1167 -2027 1168 -2025
rect 1164 -2033 1165 -2031
rect 1167 -2033 1168 -2031
rect 1171 -2027 1172 -2025
rect 1171 -2033 1172 -2031
rect 1178 -2027 1179 -2025
rect 1178 -2033 1179 -2031
rect 1185 -2027 1186 -2025
rect 1185 -2033 1186 -2031
rect 1188 -2033 1189 -2031
rect 1192 -2027 1193 -2025
rect 1192 -2033 1193 -2031
rect 1199 -2027 1200 -2025
rect 1199 -2033 1200 -2031
rect 1206 -2027 1207 -2025
rect 1206 -2033 1207 -2031
rect 1213 -2027 1214 -2025
rect 1213 -2033 1214 -2031
rect 1220 -2027 1221 -2025
rect 1220 -2033 1221 -2031
rect 1227 -2027 1228 -2025
rect 1230 -2033 1231 -2031
rect 1234 -2027 1235 -2025
rect 1234 -2033 1235 -2031
rect 1241 -2027 1242 -2025
rect 1241 -2033 1242 -2031
rect 1248 -2027 1249 -2025
rect 1248 -2033 1249 -2031
rect 1255 -2027 1256 -2025
rect 1255 -2033 1256 -2031
rect 1262 -2027 1263 -2025
rect 1262 -2033 1263 -2031
rect 1269 -2027 1270 -2025
rect 1269 -2033 1270 -2031
rect 1276 -2027 1277 -2025
rect 1276 -2033 1277 -2031
rect 1283 -2027 1284 -2025
rect 1283 -2033 1284 -2031
rect 1290 -2027 1291 -2025
rect 1290 -2033 1291 -2031
rect 1297 -2027 1298 -2025
rect 1300 -2027 1301 -2025
rect 1297 -2033 1298 -2031
rect 1300 -2033 1301 -2031
rect 1304 -2027 1305 -2025
rect 1304 -2033 1305 -2031
rect 1311 -2027 1312 -2025
rect 1311 -2033 1312 -2031
rect 1318 -2027 1319 -2025
rect 1318 -2033 1319 -2031
rect 1325 -2033 1326 -2031
rect 1332 -2027 1333 -2025
rect 1335 -2027 1336 -2025
rect 1332 -2033 1333 -2031
rect 1339 -2027 1340 -2025
rect 1339 -2033 1340 -2031
rect 1346 -2027 1347 -2025
rect 1346 -2033 1347 -2031
rect 1353 -2027 1354 -2025
rect 1353 -2033 1354 -2031
rect 1360 -2027 1361 -2025
rect 1363 -2027 1364 -2025
rect 1360 -2033 1361 -2031
rect 1363 -2033 1364 -2031
rect 1367 -2027 1368 -2025
rect 1367 -2033 1368 -2031
rect 1374 -2027 1375 -2025
rect 1374 -2033 1375 -2031
rect 1381 -2027 1382 -2025
rect 1381 -2033 1382 -2031
rect 1388 -2027 1389 -2025
rect 1388 -2033 1389 -2031
rect 1395 -2027 1396 -2025
rect 1395 -2033 1396 -2031
rect 1402 -2027 1403 -2025
rect 1402 -2033 1403 -2031
rect 1409 -2027 1410 -2025
rect 1409 -2033 1410 -2031
rect 1416 -2027 1417 -2025
rect 1416 -2033 1417 -2031
rect 1423 -2027 1424 -2025
rect 1423 -2033 1424 -2031
rect 1430 -2027 1431 -2025
rect 1430 -2033 1431 -2031
rect 1437 -2027 1438 -2025
rect 1440 -2027 1441 -2025
rect 1437 -2033 1438 -2031
rect 1440 -2033 1441 -2031
rect 1444 -2027 1445 -2025
rect 1444 -2033 1445 -2031
rect 1451 -2027 1452 -2025
rect 1451 -2033 1452 -2031
rect 1458 -2027 1459 -2025
rect 1458 -2033 1459 -2031
rect 1465 -2027 1466 -2025
rect 1465 -2033 1466 -2031
rect 1472 -2027 1473 -2025
rect 1475 -2027 1476 -2025
rect 1475 -2033 1476 -2031
rect 1479 -2027 1480 -2025
rect 1479 -2033 1480 -2031
rect 1486 -2027 1487 -2025
rect 1489 -2027 1490 -2025
rect 1486 -2033 1487 -2031
rect 1489 -2033 1490 -2031
rect 1493 -2027 1494 -2025
rect 1496 -2027 1497 -2025
rect 1493 -2033 1494 -2031
rect 1496 -2033 1497 -2031
rect 1500 -2027 1501 -2025
rect 1500 -2033 1501 -2031
rect 1507 -2027 1508 -2025
rect 1507 -2033 1508 -2031
rect 1514 -2027 1515 -2025
rect 1514 -2033 1515 -2031
rect 1524 -2027 1525 -2025
rect 1521 -2033 1522 -2031
rect 1528 -2027 1529 -2025
rect 1528 -2033 1529 -2031
rect 1535 -2027 1536 -2025
rect 1535 -2033 1536 -2031
rect 1538 -2033 1539 -2031
rect 1542 -2027 1543 -2025
rect 1542 -2033 1543 -2031
rect 1549 -2027 1550 -2025
rect 1549 -2033 1550 -2031
rect 1552 -2033 1553 -2031
rect 1556 -2027 1557 -2025
rect 1556 -2033 1557 -2031
rect 1563 -2027 1564 -2025
rect 1563 -2033 1564 -2031
rect 1570 -2027 1571 -2025
rect 1570 -2033 1571 -2031
rect 1577 -2027 1578 -2025
rect 1577 -2033 1578 -2031
rect 1584 -2027 1585 -2025
rect 1584 -2033 1585 -2031
rect 1591 -2027 1592 -2025
rect 1591 -2033 1592 -2031
rect 1598 -2027 1599 -2025
rect 1598 -2033 1599 -2031
rect 1605 -2027 1606 -2025
rect 1605 -2033 1606 -2031
rect 1612 -2027 1613 -2025
rect 1612 -2033 1613 -2031
rect 1619 -2027 1620 -2025
rect 1622 -2027 1623 -2025
rect 1619 -2033 1620 -2031
rect 1622 -2033 1623 -2031
rect 1626 -2027 1627 -2025
rect 1626 -2033 1627 -2031
rect 1633 -2027 1634 -2025
rect 1636 -2027 1637 -2025
rect 1633 -2033 1634 -2031
rect 1636 -2033 1637 -2031
rect 1640 -2027 1641 -2025
rect 1640 -2033 1641 -2031
rect 1647 -2027 1648 -2025
rect 1647 -2033 1648 -2031
rect 1654 -2027 1655 -2025
rect 1654 -2033 1655 -2031
rect 1661 -2027 1662 -2025
rect 1664 -2027 1665 -2025
rect 1661 -2033 1662 -2031
rect 1664 -2033 1665 -2031
rect 1668 -2027 1669 -2025
rect 1668 -2033 1669 -2031
rect 1675 -2027 1676 -2025
rect 1675 -2033 1676 -2031
rect 1682 -2027 1683 -2025
rect 1682 -2033 1683 -2031
rect 1689 -2027 1690 -2025
rect 1689 -2033 1690 -2031
rect 1696 -2027 1697 -2025
rect 1696 -2033 1697 -2031
rect 1703 -2027 1704 -2025
rect 1703 -2033 1704 -2031
rect 1710 -2027 1711 -2025
rect 1710 -2033 1711 -2031
rect 1717 -2027 1718 -2025
rect 1717 -2033 1718 -2031
rect 1724 -2027 1725 -2025
rect 1724 -2033 1725 -2031
rect 1731 -2027 1732 -2025
rect 1734 -2027 1735 -2025
rect 1738 -2027 1739 -2025
rect 1738 -2033 1739 -2031
rect 1745 -2027 1746 -2025
rect 1745 -2033 1746 -2031
rect 1752 -2027 1753 -2025
rect 1752 -2033 1753 -2031
rect 1759 -2027 1760 -2025
rect 1759 -2033 1760 -2031
rect 1766 -2027 1767 -2025
rect 1766 -2033 1767 -2031
rect 1773 -2027 1774 -2025
rect 1773 -2033 1774 -2031
rect 1780 -2027 1781 -2025
rect 1780 -2033 1781 -2031
rect 1787 -2027 1788 -2025
rect 1787 -2033 1788 -2031
rect 1794 -2027 1795 -2025
rect 1794 -2033 1795 -2031
rect 1801 -2027 1802 -2025
rect 1801 -2033 1802 -2031
rect 1808 -2027 1809 -2025
rect 1808 -2033 1809 -2031
rect 1815 -2027 1816 -2025
rect 1815 -2033 1816 -2031
rect 1822 -2027 1823 -2025
rect 1822 -2033 1823 -2031
rect 1829 -2027 1830 -2025
rect 1829 -2033 1830 -2031
rect 1836 -2027 1837 -2025
rect 1836 -2033 1837 -2031
rect 1843 -2027 1844 -2025
rect 1843 -2033 1844 -2031
rect 1850 -2027 1851 -2025
rect 1850 -2033 1851 -2031
rect 1857 -2027 1858 -2025
rect 1857 -2033 1858 -2031
rect 1864 -2027 1865 -2025
rect 1864 -2033 1865 -2031
rect 1871 -2027 1872 -2025
rect 1871 -2033 1872 -2031
rect 1878 -2027 1879 -2025
rect 1878 -2033 1879 -2031
rect 1885 -2027 1886 -2025
rect 1885 -2033 1886 -2031
rect 1892 -2027 1893 -2025
rect 1892 -2033 1893 -2031
rect 1899 -2027 1900 -2025
rect 1899 -2033 1900 -2031
rect 1906 -2027 1907 -2025
rect 1906 -2033 1907 -2031
rect 1913 -2027 1914 -2025
rect 1913 -2033 1914 -2031
rect 1920 -2027 1921 -2025
rect 1920 -2033 1921 -2031
rect 1927 -2027 1928 -2025
rect 1927 -2033 1928 -2031
rect 1934 -2027 1935 -2025
rect 1934 -2033 1935 -2031
rect 1941 -2027 1942 -2025
rect 1941 -2033 1942 -2031
rect 1948 -2027 1949 -2025
rect 1948 -2033 1949 -2031
rect 1955 -2027 1956 -2025
rect 1955 -2033 1956 -2031
rect 1962 -2027 1963 -2025
rect 1962 -2033 1963 -2031
rect 1969 -2027 1970 -2025
rect 1969 -2033 1970 -2031
rect 1976 -2027 1977 -2025
rect 1976 -2033 1977 -2031
rect 1983 -2027 1984 -2025
rect 1983 -2033 1984 -2031
rect 1990 -2027 1991 -2025
rect 1990 -2033 1991 -2031
rect 1997 -2027 1998 -2025
rect 1997 -2033 1998 -2031
rect 2004 -2027 2005 -2025
rect 2004 -2033 2005 -2031
rect 2011 -2027 2012 -2025
rect 2011 -2033 2012 -2031
rect 2018 -2027 2019 -2025
rect 2018 -2033 2019 -2031
rect 2025 -2027 2026 -2025
rect 2025 -2033 2026 -2031
rect 2032 -2027 2033 -2025
rect 2032 -2033 2033 -2031
rect 2039 -2027 2040 -2025
rect 2039 -2033 2040 -2031
rect 2046 -2027 2047 -2025
rect 2046 -2033 2047 -2031
rect 2053 -2027 2054 -2025
rect 2053 -2033 2054 -2031
rect 2060 -2027 2061 -2025
rect 2060 -2033 2061 -2031
rect 2067 -2027 2068 -2025
rect 2067 -2033 2068 -2031
rect 2074 -2027 2075 -2025
rect 2074 -2033 2075 -2031
rect 2081 -2027 2082 -2025
rect 2081 -2033 2082 -2031
rect 2088 -2027 2089 -2025
rect 2088 -2033 2089 -2031
rect 2095 -2027 2096 -2025
rect 2095 -2033 2096 -2031
rect 2102 -2027 2103 -2025
rect 2102 -2033 2103 -2031
rect 2109 -2027 2110 -2025
rect 2109 -2033 2110 -2031
rect 2116 -2027 2117 -2025
rect 2116 -2033 2117 -2031
rect 2123 -2027 2124 -2025
rect 2123 -2033 2124 -2031
rect 2130 -2027 2131 -2025
rect 2130 -2033 2131 -2031
rect 2137 -2027 2138 -2025
rect 2137 -2033 2138 -2031
rect 2144 -2027 2145 -2025
rect 2144 -2033 2145 -2031
rect 2151 -2027 2152 -2025
rect 2151 -2033 2152 -2031
rect 2158 -2027 2159 -2025
rect 2158 -2033 2159 -2031
rect 2165 -2027 2166 -2025
rect 2165 -2033 2166 -2031
rect 2172 -2027 2173 -2025
rect 2172 -2033 2173 -2031
rect 2179 -2027 2180 -2025
rect 2179 -2033 2180 -2031
rect 2186 -2027 2187 -2025
rect 2186 -2033 2187 -2031
rect 2193 -2027 2194 -2025
rect 2193 -2033 2194 -2031
rect 2200 -2027 2201 -2025
rect 2200 -2033 2201 -2031
rect 2207 -2027 2208 -2025
rect 2207 -2033 2208 -2031
rect 2214 -2027 2215 -2025
rect 2214 -2033 2215 -2031
rect 2221 -2027 2222 -2025
rect 2221 -2033 2222 -2031
rect 2228 -2027 2229 -2025
rect 2228 -2033 2229 -2031
rect 2235 -2027 2236 -2025
rect 2235 -2033 2236 -2031
rect 2242 -2027 2243 -2025
rect 2242 -2033 2243 -2031
rect 2249 -2027 2250 -2025
rect 2249 -2033 2250 -2031
rect 2256 -2027 2257 -2025
rect 2256 -2033 2257 -2031
rect 2263 -2027 2264 -2025
rect 2263 -2033 2264 -2031
rect 2270 -2027 2271 -2025
rect 2270 -2033 2271 -2031
rect 2277 -2027 2278 -2025
rect 2277 -2033 2278 -2031
rect 2284 -2027 2285 -2025
rect 2284 -2033 2285 -2031
rect 2291 -2027 2292 -2025
rect 2291 -2033 2292 -2031
rect 2298 -2027 2299 -2025
rect 2298 -2033 2299 -2031
rect 2305 -2027 2306 -2025
rect 2305 -2033 2306 -2031
rect 2312 -2027 2313 -2025
rect 2312 -2033 2313 -2031
rect 2319 -2027 2320 -2025
rect 2319 -2033 2320 -2031
rect 2326 -2027 2327 -2025
rect 2326 -2033 2327 -2031
rect 2333 -2027 2334 -2025
rect 2333 -2033 2334 -2031
rect 2340 -2027 2341 -2025
rect 2340 -2033 2341 -2031
rect 2347 -2027 2348 -2025
rect 2347 -2033 2348 -2031
rect 2354 -2027 2355 -2025
rect 2354 -2033 2355 -2031
rect 2361 -2027 2362 -2025
rect 2361 -2033 2362 -2031
rect 2368 -2027 2369 -2025
rect 2368 -2033 2369 -2031
rect 2375 -2027 2376 -2025
rect 2375 -2033 2376 -2031
rect 2382 -2027 2383 -2025
rect 2382 -2033 2383 -2031
rect 2389 -2027 2390 -2025
rect 2389 -2033 2390 -2031
rect 2396 -2027 2397 -2025
rect 2396 -2033 2397 -2031
rect 2403 -2027 2404 -2025
rect 2403 -2033 2404 -2031
rect 2410 -2027 2411 -2025
rect 2410 -2033 2411 -2031
rect 2420 -2027 2421 -2025
rect 2424 -2027 2425 -2025
rect 2424 -2033 2425 -2031
rect 9 -2178 10 -2176
rect 9 -2184 10 -2182
rect 16 -2178 17 -2176
rect 16 -2184 17 -2182
rect 23 -2178 24 -2176
rect 23 -2184 24 -2182
rect 30 -2178 31 -2176
rect 30 -2184 31 -2182
rect 37 -2178 38 -2176
rect 40 -2184 41 -2182
rect 44 -2178 45 -2176
rect 44 -2184 45 -2182
rect 51 -2178 52 -2176
rect 51 -2184 52 -2182
rect 54 -2184 55 -2182
rect 58 -2178 59 -2176
rect 58 -2184 59 -2182
rect 65 -2178 66 -2176
rect 65 -2184 66 -2182
rect 72 -2178 73 -2176
rect 72 -2184 73 -2182
rect 79 -2178 80 -2176
rect 79 -2184 80 -2182
rect 86 -2178 87 -2176
rect 86 -2184 87 -2182
rect 93 -2178 94 -2176
rect 96 -2178 97 -2176
rect 93 -2184 94 -2182
rect 96 -2184 97 -2182
rect 100 -2178 101 -2176
rect 100 -2184 101 -2182
rect 107 -2178 108 -2176
rect 107 -2184 108 -2182
rect 114 -2178 115 -2176
rect 114 -2184 115 -2182
rect 121 -2178 122 -2176
rect 124 -2178 125 -2176
rect 121 -2184 122 -2182
rect 124 -2184 125 -2182
rect 131 -2178 132 -2176
rect 128 -2184 129 -2182
rect 131 -2184 132 -2182
rect 135 -2178 136 -2176
rect 138 -2178 139 -2176
rect 135 -2184 136 -2182
rect 138 -2184 139 -2182
rect 142 -2178 143 -2176
rect 142 -2184 143 -2182
rect 149 -2178 150 -2176
rect 149 -2184 150 -2182
rect 156 -2178 157 -2176
rect 156 -2184 157 -2182
rect 163 -2178 164 -2176
rect 163 -2184 164 -2182
rect 170 -2178 171 -2176
rect 170 -2184 171 -2182
rect 177 -2178 178 -2176
rect 177 -2184 178 -2182
rect 184 -2178 185 -2176
rect 184 -2184 185 -2182
rect 191 -2178 192 -2176
rect 191 -2184 192 -2182
rect 198 -2178 199 -2176
rect 198 -2184 199 -2182
rect 205 -2178 206 -2176
rect 205 -2184 206 -2182
rect 212 -2178 213 -2176
rect 212 -2184 213 -2182
rect 219 -2178 220 -2176
rect 219 -2184 220 -2182
rect 226 -2178 227 -2176
rect 226 -2184 227 -2182
rect 233 -2178 234 -2176
rect 236 -2178 237 -2176
rect 233 -2184 234 -2182
rect 236 -2184 237 -2182
rect 240 -2178 241 -2176
rect 243 -2178 244 -2176
rect 247 -2178 248 -2176
rect 247 -2184 248 -2182
rect 257 -2178 258 -2176
rect 257 -2184 258 -2182
rect 261 -2178 262 -2176
rect 261 -2184 262 -2182
rect 268 -2178 269 -2176
rect 268 -2184 269 -2182
rect 275 -2178 276 -2176
rect 275 -2184 276 -2182
rect 282 -2178 283 -2176
rect 282 -2184 283 -2182
rect 289 -2178 290 -2176
rect 289 -2184 290 -2182
rect 296 -2178 297 -2176
rect 296 -2184 297 -2182
rect 303 -2178 304 -2176
rect 303 -2184 304 -2182
rect 310 -2178 311 -2176
rect 310 -2184 311 -2182
rect 317 -2178 318 -2176
rect 317 -2184 318 -2182
rect 324 -2178 325 -2176
rect 324 -2184 325 -2182
rect 331 -2178 332 -2176
rect 331 -2184 332 -2182
rect 338 -2178 339 -2176
rect 338 -2184 339 -2182
rect 345 -2178 346 -2176
rect 345 -2184 346 -2182
rect 352 -2178 353 -2176
rect 352 -2184 353 -2182
rect 359 -2178 360 -2176
rect 359 -2184 360 -2182
rect 366 -2178 367 -2176
rect 366 -2184 367 -2182
rect 373 -2178 374 -2176
rect 373 -2184 374 -2182
rect 380 -2178 381 -2176
rect 380 -2184 381 -2182
rect 387 -2178 388 -2176
rect 387 -2184 388 -2182
rect 394 -2178 395 -2176
rect 394 -2184 395 -2182
rect 401 -2178 402 -2176
rect 404 -2178 405 -2176
rect 401 -2184 402 -2182
rect 408 -2178 409 -2176
rect 408 -2184 409 -2182
rect 415 -2178 416 -2176
rect 415 -2184 416 -2182
rect 422 -2178 423 -2176
rect 422 -2184 423 -2182
rect 429 -2178 430 -2176
rect 429 -2184 430 -2182
rect 436 -2178 437 -2176
rect 436 -2184 437 -2182
rect 443 -2178 444 -2176
rect 443 -2184 444 -2182
rect 450 -2178 451 -2176
rect 450 -2184 451 -2182
rect 457 -2178 458 -2176
rect 457 -2184 458 -2182
rect 464 -2178 465 -2176
rect 464 -2184 465 -2182
rect 471 -2178 472 -2176
rect 471 -2184 472 -2182
rect 478 -2178 479 -2176
rect 478 -2184 479 -2182
rect 485 -2178 486 -2176
rect 485 -2184 486 -2182
rect 492 -2178 493 -2176
rect 492 -2184 493 -2182
rect 495 -2184 496 -2182
rect 499 -2178 500 -2176
rect 499 -2184 500 -2182
rect 506 -2178 507 -2176
rect 506 -2184 507 -2182
rect 513 -2178 514 -2176
rect 516 -2178 517 -2176
rect 513 -2184 514 -2182
rect 516 -2184 517 -2182
rect 520 -2178 521 -2176
rect 520 -2184 521 -2182
rect 527 -2178 528 -2176
rect 527 -2184 528 -2182
rect 534 -2178 535 -2176
rect 534 -2184 535 -2182
rect 541 -2178 542 -2176
rect 541 -2184 542 -2182
rect 548 -2178 549 -2176
rect 548 -2184 549 -2182
rect 555 -2178 556 -2176
rect 555 -2184 556 -2182
rect 562 -2178 563 -2176
rect 562 -2184 563 -2182
rect 569 -2178 570 -2176
rect 569 -2184 570 -2182
rect 576 -2178 577 -2176
rect 576 -2184 577 -2182
rect 583 -2178 584 -2176
rect 583 -2184 584 -2182
rect 590 -2178 591 -2176
rect 590 -2184 591 -2182
rect 597 -2178 598 -2176
rect 597 -2184 598 -2182
rect 604 -2178 605 -2176
rect 604 -2184 605 -2182
rect 611 -2178 612 -2176
rect 611 -2184 612 -2182
rect 618 -2178 619 -2176
rect 618 -2184 619 -2182
rect 625 -2178 626 -2176
rect 625 -2184 626 -2182
rect 632 -2178 633 -2176
rect 632 -2184 633 -2182
rect 639 -2178 640 -2176
rect 639 -2184 640 -2182
rect 646 -2178 647 -2176
rect 646 -2184 647 -2182
rect 653 -2178 654 -2176
rect 656 -2178 657 -2176
rect 656 -2184 657 -2182
rect 660 -2178 661 -2176
rect 660 -2184 661 -2182
rect 667 -2178 668 -2176
rect 670 -2178 671 -2176
rect 670 -2184 671 -2182
rect 674 -2178 675 -2176
rect 674 -2184 675 -2182
rect 681 -2178 682 -2176
rect 681 -2184 682 -2182
rect 688 -2178 689 -2176
rect 688 -2184 689 -2182
rect 695 -2178 696 -2176
rect 695 -2184 696 -2182
rect 702 -2178 703 -2176
rect 702 -2184 703 -2182
rect 709 -2178 710 -2176
rect 709 -2184 710 -2182
rect 716 -2178 717 -2176
rect 716 -2184 717 -2182
rect 723 -2178 724 -2176
rect 723 -2184 724 -2182
rect 730 -2178 731 -2176
rect 730 -2184 731 -2182
rect 737 -2178 738 -2176
rect 737 -2184 738 -2182
rect 744 -2178 745 -2176
rect 747 -2178 748 -2176
rect 744 -2184 745 -2182
rect 747 -2184 748 -2182
rect 751 -2178 752 -2176
rect 751 -2184 752 -2182
rect 758 -2178 759 -2176
rect 761 -2178 762 -2176
rect 758 -2184 759 -2182
rect 765 -2178 766 -2176
rect 765 -2184 766 -2182
rect 772 -2178 773 -2176
rect 772 -2184 773 -2182
rect 779 -2178 780 -2176
rect 779 -2184 780 -2182
rect 786 -2178 787 -2176
rect 786 -2184 787 -2182
rect 789 -2184 790 -2182
rect 793 -2178 794 -2176
rect 793 -2184 794 -2182
rect 800 -2178 801 -2176
rect 800 -2184 801 -2182
rect 807 -2178 808 -2176
rect 807 -2184 808 -2182
rect 814 -2178 815 -2176
rect 814 -2184 815 -2182
rect 821 -2178 822 -2176
rect 821 -2184 822 -2182
rect 828 -2178 829 -2176
rect 828 -2184 829 -2182
rect 835 -2178 836 -2176
rect 835 -2184 836 -2182
rect 842 -2178 843 -2176
rect 842 -2184 843 -2182
rect 849 -2178 850 -2176
rect 849 -2184 850 -2182
rect 856 -2178 857 -2176
rect 856 -2184 857 -2182
rect 863 -2178 864 -2176
rect 863 -2184 864 -2182
rect 870 -2178 871 -2176
rect 870 -2184 871 -2182
rect 877 -2178 878 -2176
rect 877 -2184 878 -2182
rect 884 -2178 885 -2176
rect 884 -2184 885 -2182
rect 891 -2178 892 -2176
rect 891 -2184 892 -2182
rect 898 -2178 899 -2176
rect 898 -2184 899 -2182
rect 905 -2178 906 -2176
rect 905 -2184 906 -2182
rect 912 -2178 913 -2176
rect 912 -2184 913 -2182
rect 919 -2178 920 -2176
rect 919 -2184 920 -2182
rect 926 -2178 927 -2176
rect 926 -2184 927 -2182
rect 933 -2178 934 -2176
rect 933 -2184 934 -2182
rect 940 -2178 941 -2176
rect 940 -2184 941 -2182
rect 947 -2178 948 -2176
rect 947 -2184 948 -2182
rect 954 -2178 955 -2176
rect 954 -2184 955 -2182
rect 961 -2178 962 -2176
rect 961 -2184 962 -2182
rect 968 -2178 969 -2176
rect 968 -2184 969 -2182
rect 975 -2178 976 -2176
rect 978 -2178 979 -2176
rect 975 -2184 976 -2182
rect 978 -2184 979 -2182
rect 982 -2178 983 -2176
rect 982 -2184 983 -2182
rect 989 -2178 990 -2176
rect 989 -2184 990 -2182
rect 996 -2178 997 -2176
rect 996 -2184 997 -2182
rect 1003 -2178 1004 -2176
rect 1003 -2184 1004 -2182
rect 1010 -2178 1011 -2176
rect 1010 -2184 1011 -2182
rect 1017 -2178 1018 -2176
rect 1017 -2184 1018 -2182
rect 1024 -2178 1025 -2176
rect 1024 -2184 1025 -2182
rect 1031 -2178 1032 -2176
rect 1031 -2184 1032 -2182
rect 1038 -2178 1039 -2176
rect 1038 -2184 1039 -2182
rect 1045 -2178 1046 -2176
rect 1045 -2184 1046 -2182
rect 1052 -2178 1053 -2176
rect 1055 -2178 1056 -2176
rect 1052 -2184 1053 -2182
rect 1055 -2184 1056 -2182
rect 1059 -2178 1060 -2176
rect 1059 -2184 1060 -2182
rect 1066 -2178 1067 -2176
rect 1066 -2184 1067 -2182
rect 1073 -2178 1074 -2176
rect 1073 -2184 1074 -2182
rect 1080 -2178 1081 -2176
rect 1080 -2184 1081 -2182
rect 1087 -2178 1088 -2176
rect 1087 -2184 1088 -2182
rect 1094 -2178 1095 -2176
rect 1094 -2184 1095 -2182
rect 1101 -2178 1102 -2176
rect 1101 -2184 1102 -2182
rect 1108 -2178 1109 -2176
rect 1108 -2184 1109 -2182
rect 1115 -2178 1116 -2176
rect 1115 -2184 1116 -2182
rect 1122 -2178 1123 -2176
rect 1122 -2184 1123 -2182
rect 1129 -2178 1130 -2176
rect 1129 -2184 1130 -2182
rect 1136 -2178 1137 -2176
rect 1136 -2184 1137 -2182
rect 1143 -2178 1144 -2176
rect 1143 -2184 1144 -2182
rect 1150 -2178 1151 -2176
rect 1153 -2178 1154 -2176
rect 1157 -2178 1158 -2176
rect 1157 -2184 1158 -2182
rect 1164 -2178 1165 -2176
rect 1164 -2184 1165 -2182
rect 1171 -2178 1172 -2176
rect 1171 -2184 1172 -2182
rect 1178 -2178 1179 -2176
rect 1178 -2184 1179 -2182
rect 1185 -2178 1186 -2176
rect 1188 -2178 1189 -2176
rect 1185 -2184 1186 -2182
rect 1188 -2184 1189 -2182
rect 1192 -2178 1193 -2176
rect 1192 -2184 1193 -2182
rect 1199 -2178 1200 -2176
rect 1202 -2178 1203 -2176
rect 1199 -2184 1200 -2182
rect 1202 -2184 1203 -2182
rect 1206 -2178 1207 -2176
rect 1206 -2184 1207 -2182
rect 1213 -2178 1214 -2176
rect 1213 -2184 1214 -2182
rect 1220 -2178 1221 -2176
rect 1223 -2178 1224 -2176
rect 1220 -2184 1221 -2182
rect 1223 -2184 1224 -2182
rect 1230 -2178 1231 -2176
rect 1227 -2184 1228 -2182
rect 1230 -2184 1231 -2182
rect 1234 -2178 1235 -2176
rect 1234 -2184 1235 -2182
rect 1241 -2178 1242 -2176
rect 1241 -2184 1242 -2182
rect 1248 -2178 1249 -2176
rect 1248 -2184 1249 -2182
rect 1255 -2178 1256 -2176
rect 1258 -2178 1259 -2176
rect 1255 -2184 1256 -2182
rect 1258 -2184 1259 -2182
rect 1262 -2178 1263 -2176
rect 1262 -2184 1263 -2182
rect 1269 -2178 1270 -2176
rect 1269 -2184 1270 -2182
rect 1276 -2178 1277 -2176
rect 1276 -2184 1277 -2182
rect 1283 -2178 1284 -2176
rect 1283 -2184 1284 -2182
rect 1290 -2178 1291 -2176
rect 1290 -2184 1291 -2182
rect 1297 -2178 1298 -2176
rect 1297 -2184 1298 -2182
rect 1304 -2178 1305 -2176
rect 1307 -2178 1308 -2176
rect 1304 -2184 1305 -2182
rect 1307 -2184 1308 -2182
rect 1311 -2178 1312 -2176
rect 1311 -2184 1312 -2182
rect 1318 -2178 1319 -2176
rect 1318 -2184 1319 -2182
rect 1325 -2178 1326 -2176
rect 1325 -2184 1326 -2182
rect 1332 -2178 1333 -2176
rect 1335 -2178 1336 -2176
rect 1332 -2184 1333 -2182
rect 1335 -2184 1336 -2182
rect 1339 -2178 1340 -2176
rect 1342 -2178 1343 -2176
rect 1339 -2184 1340 -2182
rect 1342 -2184 1343 -2182
rect 1346 -2178 1347 -2176
rect 1346 -2184 1347 -2182
rect 1353 -2178 1354 -2176
rect 1353 -2184 1354 -2182
rect 1360 -2178 1361 -2176
rect 1360 -2184 1361 -2182
rect 1367 -2178 1368 -2176
rect 1367 -2184 1368 -2182
rect 1370 -2184 1371 -2182
rect 1374 -2178 1375 -2176
rect 1374 -2184 1375 -2182
rect 1381 -2178 1382 -2176
rect 1384 -2178 1385 -2176
rect 1381 -2184 1382 -2182
rect 1384 -2184 1385 -2182
rect 1388 -2178 1389 -2176
rect 1388 -2184 1389 -2182
rect 1395 -2178 1396 -2176
rect 1395 -2184 1396 -2182
rect 1402 -2178 1403 -2176
rect 1405 -2178 1406 -2176
rect 1402 -2184 1403 -2182
rect 1405 -2184 1406 -2182
rect 1409 -2178 1410 -2176
rect 1409 -2184 1410 -2182
rect 1416 -2178 1417 -2176
rect 1416 -2184 1417 -2182
rect 1423 -2178 1424 -2176
rect 1423 -2184 1424 -2182
rect 1430 -2178 1431 -2176
rect 1430 -2184 1431 -2182
rect 1437 -2178 1438 -2176
rect 1437 -2184 1438 -2182
rect 1444 -2178 1445 -2176
rect 1444 -2184 1445 -2182
rect 1451 -2178 1452 -2176
rect 1451 -2184 1452 -2182
rect 1458 -2178 1459 -2176
rect 1458 -2184 1459 -2182
rect 1465 -2178 1466 -2176
rect 1465 -2184 1466 -2182
rect 1472 -2178 1473 -2176
rect 1472 -2184 1473 -2182
rect 1479 -2178 1480 -2176
rect 1479 -2184 1480 -2182
rect 1486 -2178 1487 -2176
rect 1489 -2178 1490 -2176
rect 1486 -2184 1487 -2182
rect 1489 -2184 1490 -2182
rect 1493 -2178 1494 -2176
rect 1493 -2184 1494 -2182
rect 1500 -2178 1501 -2176
rect 1500 -2184 1501 -2182
rect 1507 -2178 1508 -2176
rect 1507 -2184 1508 -2182
rect 1514 -2178 1515 -2176
rect 1514 -2184 1515 -2182
rect 1521 -2178 1522 -2176
rect 1521 -2184 1522 -2182
rect 1528 -2178 1529 -2176
rect 1528 -2184 1529 -2182
rect 1535 -2178 1536 -2176
rect 1535 -2184 1536 -2182
rect 1542 -2178 1543 -2176
rect 1542 -2184 1543 -2182
rect 1549 -2178 1550 -2176
rect 1549 -2184 1550 -2182
rect 1556 -2178 1557 -2176
rect 1556 -2184 1557 -2182
rect 1563 -2178 1564 -2176
rect 1563 -2184 1564 -2182
rect 1570 -2178 1571 -2176
rect 1570 -2184 1571 -2182
rect 1577 -2178 1578 -2176
rect 1580 -2178 1581 -2176
rect 1580 -2184 1581 -2182
rect 1584 -2178 1585 -2176
rect 1584 -2184 1585 -2182
rect 1591 -2178 1592 -2176
rect 1591 -2184 1592 -2182
rect 1598 -2178 1599 -2176
rect 1598 -2184 1599 -2182
rect 1605 -2178 1606 -2176
rect 1605 -2184 1606 -2182
rect 1612 -2178 1613 -2176
rect 1612 -2184 1613 -2182
rect 1619 -2178 1620 -2176
rect 1619 -2184 1620 -2182
rect 1626 -2178 1627 -2176
rect 1626 -2184 1627 -2182
rect 1633 -2178 1634 -2176
rect 1633 -2184 1634 -2182
rect 1640 -2178 1641 -2176
rect 1640 -2184 1641 -2182
rect 1647 -2178 1648 -2176
rect 1650 -2178 1651 -2176
rect 1647 -2184 1648 -2182
rect 1650 -2184 1651 -2182
rect 1654 -2178 1655 -2176
rect 1654 -2184 1655 -2182
rect 1661 -2178 1662 -2176
rect 1661 -2184 1662 -2182
rect 1668 -2178 1669 -2176
rect 1668 -2184 1669 -2182
rect 1675 -2178 1676 -2176
rect 1675 -2184 1676 -2182
rect 1682 -2178 1683 -2176
rect 1682 -2184 1683 -2182
rect 1689 -2178 1690 -2176
rect 1689 -2184 1690 -2182
rect 1696 -2178 1697 -2176
rect 1696 -2184 1697 -2182
rect 1703 -2178 1704 -2176
rect 1703 -2184 1704 -2182
rect 1713 -2178 1714 -2176
rect 1717 -2178 1718 -2176
rect 1717 -2184 1718 -2182
rect 1724 -2178 1725 -2176
rect 1724 -2184 1725 -2182
rect 1731 -2178 1732 -2176
rect 1731 -2184 1732 -2182
rect 1738 -2178 1739 -2176
rect 1738 -2184 1739 -2182
rect 1745 -2178 1746 -2176
rect 1745 -2184 1746 -2182
rect 1752 -2178 1753 -2176
rect 1752 -2184 1753 -2182
rect 1759 -2178 1760 -2176
rect 1759 -2184 1760 -2182
rect 1766 -2178 1767 -2176
rect 1766 -2184 1767 -2182
rect 1773 -2178 1774 -2176
rect 1773 -2184 1774 -2182
rect 1780 -2178 1781 -2176
rect 1780 -2184 1781 -2182
rect 1787 -2178 1788 -2176
rect 1787 -2184 1788 -2182
rect 1794 -2178 1795 -2176
rect 1794 -2184 1795 -2182
rect 1801 -2178 1802 -2176
rect 1801 -2184 1802 -2182
rect 1808 -2178 1809 -2176
rect 1808 -2184 1809 -2182
rect 1815 -2178 1816 -2176
rect 1815 -2184 1816 -2182
rect 1822 -2178 1823 -2176
rect 1822 -2184 1823 -2182
rect 1829 -2178 1830 -2176
rect 1829 -2184 1830 -2182
rect 1836 -2178 1837 -2176
rect 1843 -2178 1844 -2176
rect 1843 -2184 1844 -2182
rect 1850 -2178 1851 -2176
rect 1850 -2184 1851 -2182
rect 1857 -2178 1858 -2176
rect 1857 -2184 1858 -2182
rect 1860 -2184 1861 -2182
rect 1864 -2178 1865 -2176
rect 1864 -2184 1865 -2182
rect 1871 -2178 1872 -2176
rect 1871 -2184 1872 -2182
rect 1878 -2178 1879 -2176
rect 1878 -2184 1879 -2182
rect 1885 -2178 1886 -2176
rect 1885 -2184 1886 -2182
rect 1892 -2178 1893 -2176
rect 1892 -2184 1893 -2182
rect 1899 -2178 1900 -2176
rect 1899 -2184 1900 -2182
rect 1906 -2178 1907 -2176
rect 1906 -2184 1907 -2182
rect 1913 -2178 1914 -2176
rect 1913 -2184 1914 -2182
rect 1920 -2178 1921 -2176
rect 1920 -2184 1921 -2182
rect 1927 -2178 1928 -2176
rect 1927 -2184 1928 -2182
rect 1934 -2178 1935 -2176
rect 1934 -2184 1935 -2182
rect 1941 -2178 1942 -2176
rect 1941 -2184 1942 -2182
rect 1948 -2178 1949 -2176
rect 1948 -2184 1949 -2182
rect 1955 -2178 1956 -2176
rect 1955 -2184 1956 -2182
rect 1962 -2178 1963 -2176
rect 1962 -2184 1963 -2182
rect 1969 -2178 1970 -2176
rect 1969 -2184 1970 -2182
rect 1976 -2178 1977 -2176
rect 1976 -2184 1977 -2182
rect 1983 -2178 1984 -2176
rect 1983 -2184 1984 -2182
rect 1990 -2178 1991 -2176
rect 1990 -2184 1991 -2182
rect 1997 -2178 1998 -2176
rect 1997 -2184 1998 -2182
rect 2004 -2178 2005 -2176
rect 2004 -2184 2005 -2182
rect 2011 -2178 2012 -2176
rect 2011 -2184 2012 -2182
rect 2018 -2178 2019 -2176
rect 2018 -2184 2019 -2182
rect 2025 -2178 2026 -2176
rect 2025 -2184 2026 -2182
rect 2032 -2178 2033 -2176
rect 2032 -2184 2033 -2182
rect 2039 -2178 2040 -2176
rect 2039 -2184 2040 -2182
rect 2046 -2178 2047 -2176
rect 2046 -2184 2047 -2182
rect 2053 -2178 2054 -2176
rect 2053 -2184 2054 -2182
rect 2060 -2178 2061 -2176
rect 2060 -2184 2061 -2182
rect 2067 -2178 2068 -2176
rect 2067 -2184 2068 -2182
rect 2074 -2178 2075 -2176
rect 2074 -2184 2075 -2182
rect 2081 -2178 2082 -2176
rect 2081 -2184 2082 -2182
rect 2088 -2178 2089 -2176
rect 2088 -2184 2089 -2182
rect 2095 -2178 2096 -2176
rect 2095 -2184 2096 -2182
rect 2102 -2178 2103 -2176
rect 2102 -2184 2103 -2182
rect 2109 -2178 2110 -2176
rect 2109 -2184 2110 -2182
rect 2116 -2178 2117 -2176
rect 2116 -2184 2117 -2182
rect 2123 -2178 2124 -2176
rect 2123 -2184 2124 -2182
rect 2130 -2178 2131 -2176
rect 2130 -2184 2131 -2182
rect 2137 -2178 2138 -2176
rect 2137 -2184 2138 -2182
rect 2144 -2178 2145 -2176
rect 2144 -2184 2145 -2182
rect 2151 -2178 2152 -2176
rect 2151 -2184 2152 -2182
rect 2158 -2178 2159 -2176
rect 2158 -2184 2159 -2182
rect 2165 -2178 2166 -2176
rect 2165 -2184 2166 -2182
rect 2172 -2178 2173 -2176
rect 2172 -2184 2173 -2182
rect 2179 -2178 2180 -2176
rect 2179 -2184 2180 -2182
rect 2186 -2178 2187 -2176
rect 2186 -2184 2187 -2182
rect 2193 -2178 2194 -2176
rect 2193 -2184 2194 -2182
rect 2200 -2178 2201 -2176
rect 2200 -2184 2201 -2182
rect 2207 -2178 2208 -2176
rect 2207 -2184 2208 -2182
rect 2214 -2178 2215 -2176
rect 2214 -2184 2215 -2182
rect 2221 -2178 2222 -2176
rect 2221 -2184 2222 -2182
rect 2228 -2178 2229 -2176
rect 2228 -2184 2229 -2182
rect 2235 -2178 2236 -2176
rect 2235 -2184 2236 -2182
rect 2242 -2178 2243 -2176
rect 2242 -2184 2243 -2182
rect 2249 -2178 2250 -2176
rect 2249 -2184 2250 -2182
rect 2256 -2178 2257 -2176
rect 2256 -2184 2257 -2182
rect 2263 -2178 2264 -2176
rect 2263 -2184 2264 -2182
rect 2270 -2178 2271 -2176
rect 2270 -2184 2271 -2182
rect 2277 -2178 2278 -2176
rect 2277 -2184 2278 -2182
rect 2284 -2178 2285 -2176
rect 2284 -2184 2285 -2182
rect 2291 -2178 2292 -2176
rect 2291 -2184 2292 -2182
rect 2298 -2178 2299 -2176
rect 2298 -2184 2299 -2182
rect 2305 -2178 2306 -2176
rect 2305 -2184 2306 -2182
rect 2312 -2178 2313 -2176
rect 2312 -2184 2313 -2182
rect 2319 -2178 2320 -2176
rect 2319 -2184 2320 -2182
rect 2326 -2178 2327 -2176
rect 2326 -2184 2327 -2182
rect 2333 -2178 2334 -2176
rect 2333 -2184 2334 -2182
rect 2340 -2178 2341 -2176
rect 2340 -2184 2341 -2182
rect 2347 -2178 2348 -2176
rect 2347 -2184 2348 -2182
rect 2354 -2178 2355 -2176
rect 2354 -2184 2355 -2182
rect 2361 -2178 2362 -2176
rect 2361 -2184 2362 -2182
rect 2368 -2178 2369 -2176
rect 2368 -2184 2369 -2182
rect 2375 -2178 2376 -2176
rect 2375 -2184 2376 -2182
rect 2382 -2178 2383 -2176
rect 2382 -2184 2383 -2182
rect 2389 -2178 2390 -2176
rect 2389 -2184 2390 -2182
rect 2396 -2178 2397 -2176
rect 2396 -2184 2397 -2182
rect 2403 -2178 2404 -2176
rect 2403 -2184 2404 -2182
rect 2410 -2178 2411 -2176
rect 2410 -2184 2411 -2182
rect 2417 -2178 2418 -2176
rect 2417 -2184 2418 -2182
rect 2424 -2178 2425 -2176
rect 2424 -2184 2425 -2182
rect 2 -2327 3 -2325
rect 2 -2333 3 -2331
rect 16 -2327 17 -2325
rect 16 -2333 17 -2331
rect 23 -2327 24 -2325
rect 23 -2333 24 -2331
rect 33 -2327 34 -2325
rect 30 -2333 31 -2331
rect 33 -2333 34 -2331
rect 37 -2327 38 -2325
rect 37 -2333 38 -2331
rect 44 -2327 45 -2325
rect 44 -2333 45 -2331
rect 51 -2327 52 -2325
rect 51 -2333 52 -2331
rect 58 -2327 59 -2325
rect 58 -2333 59 -2331
rect 65 -2327 66 -2325
rect 65 -2333 66 -2331
rect 72 -2327 73 -2325
rect 72 -2333 73 -2331
rect 79 -2327 80 -2325
rect 79 -2333 80 -2331
rect 86 -2327 87 -2325
rect 86 -2333 87 -2331
rect 93 -2327 94 -2325
rect 93 -2333 94 -2331
rect 96 -2333 97 -2331
rect 100 -2327 101 -2325
rect 100 -2333 101 -2331
rect 107 -2327 108 -2325
rect 107 -2333 108 -2331
rect 114 -2327 115 -2325
rect 114 -2333 115 -2331
rect 121 -2327 122 -2325
rect 121 -2333 122 -2331
rect 128 -2327 129 -2325
rect 128 -2333 129 -2331
rect 135 -2327 136 -2325
rect 135 -2333 136 -2331
rect 142 -2327 143 -2325
rect 145 -2327 146 -2325
rect 142 -2333 143 -2331
rect 145 -2333 146 -2331
rect 149 -2327 150 -2325
rect 149 -2333 150 -2331
rect 156 -2327 157 -2325
rect 156 -2333 157 -2331
rect 163 -2327 164 -2325
rect 166 -2327 167 -2325
rect 163 -2333 164 -2331
rect 166 -2333 167 -2331
rect 170 -2327 171 -2325
rect 170 -2333 171 -2331
rect 177 -2327 178 -2325
rect 184 -2327 185 -2325
rect 184 -2333 185 -2331
rect 191 -2327 192 -2325
rect 191 -2333 192 -2331
rect 198 -2327 199 -2325
rect 198 -2333 199 -2331
rect 205 -2327 206 -2325
rect 205 -2333 206 -2331
rect 212 -2327 213 -2325
rect 212 -2333 213 -2331
rect 219 -2327 220 -2325
rect 219 -2333 220 -2331
rect 226 -2327 227 -2325
rect 226 -2333 227 -2331
rect 233 -2327 234 -2325
rect 233 -2333 234 -2331
rect 243 -2327 244 -2325
rect 243 -2333 244 -2331
rect 247 -2327 248 -2325
rect 250 -2327 251 -2325
rect 247 -2333 248 -2331
rect 254 -2327 255 -2325
rect 254 -2333 255 -2331
rect 261 -2327 262 -2325
rect 261 -2333 262 -2331
rect 268 -2327 269 -2325
rect 268 -2333 269 -2331
rect 275 -2327 276 -2325
rect 275 -2333 276 -2331
rect 282 -2327 283 -2325
rect 282 -2333 283 -2331
rect 289 -2327 290 -2325
rect 289 -2333 290 -2331
rect 296 -2327 297 -2325
rect 296 -2333 297 -2331
rect 303 -2327 304 -2325
rect 303 -2333 304 -2331
rect 310 -2327 311 -2325
rect 310 -2333 311 -2331
rect 317 -2327 318 -2325
rect 317 -2333 318 -2331
rect 324 -2327 325 -2325
rect 324 -2333 325 -2331
rect 331 -2327 332 -2325
rect 331 -2333 332 -2331
rect 338 -2327 339 -2325
rect 338 -2333 339 -2331
rect 345 -2327 346 -2325
rect 345 -2333 346 -2331
rect 352 -2327 353 -2325
rect 352 -2333 353 -2331
rect 359 -2327 360 -2325
rect 359 -2333 360 -2331
rect 366 -2327 367 -2325
rect 366 -2333 367 -2331
rect 373 -2327 374 -2325
rect 373 -2333 374 -2331
rect 380 -2327 381 -2325
rect 380 -2333 381 -2331
rect 387 -2327 388 -2325
rect 387 -2333 388 -2331
rect 394 -2327 395 -2325
rect 394 -2333 395 -2331
rect 401 -2327 402 -2325
rect 401 -2333 402 -2331
rect 408 -2327 409 -2325
rect 408 -2333 409 -2331
rect 415 -2327 416 -2325
rect 415 -2333 416 -2331
rect 422 -2327 423 -2325
rect 422 -2333 423 -2331
rect 429 -2327 430 -2325
rect 436 -2327 437 -2325
rect 436 -2333 437 -2331
rect 443 -2327 444 -2325
rect 443 -2333 444 -2331
rect 450 -2327 451 -2325
rect 450 -2333 451 -2331
rect 457 -2327 458 -2325
rect 457 -2333 458 -2331
rect 464 -2327 465 -2325
rect 464 -2333 465 -2331
rect 471 -2327 472 -2325
rect 471 -2333 472 -2331
rect 478 -2327 479 -2325
rect 478 -2333 479 -2331
rect 485 -2327 486 -2325
rect 485 -2333 486 -2331
rect 492 -2327 493 -2325
rect 492 -2333 493 -2331
rect 499 -2327 500 -2325
rect 499 -2333 500 -2331
rect 506 -2327 507 -2325
rect 506 -2333 507 -2331
rect 513 -2327 514 -2325
rect 513 -2333 514 -2331
rect 520 -2327 521 -2325
rect 520 -2333 521 -2331
rect 527 -2327 528 -2325
rect 527 -2333 528 -2331
rect 534 -2327 535 -2325
rect 534 -2333 535 -2331
rect 541 -2327 542 -2325
rect 541 -2333 542 -2331
rect 548 -2327 549 -2325
rect 548 -2333 549 -2331
rect 555 -2327 556 -2325
rect 555 -2333 556 -2331
rect 562 -2327 563 -2325
rect 562 -2333 563 -2331
rect 569 -2327 570 -2325
rect 569 -2333 570 -2331
rect 576 -2327 577 -2325
rect 576 -2333 577 -2331
rect 583 -2327 584 -2325
rect 583 -2333 584 -2331
rect 590 -2327 591 -2325
rect 593 -2327 594 -2325
rect 593 -2333 594 -2331
rect 597 -2327 598 -2325
rect 597 -2333 598 -2331
rect 604 -2327 605 -2325
rect 604 -2333 605 -2331
rect 611 -2327 612 -2325
rect 611 -2333 612 -2331
rect 618 -2327 619 -2325
rect 621 -2327 622 -2325
rect 618 -2333 619 -2331
rect 621 -2333 622 -2331
rect 625 -2327 626 -2325
rect 628 -2333 629 -2331
rect 632 -2327 633 -2325
rect 632 -2333 633 -2331
rect 639 -2327 640 -2325
rect 639 -2333 640 -2331
rect 646 -2327 647 -2325
rect 646 -2333 647 -2331
rect 653 -2327 654 -2325
rect 653 -2333 654 -2331
rect 660 -2327 661 -2325
rect 663 -2327 664 -2325
rect 660 -2333 661 -2331
rect 667 -2327 668 -2325
rect 670 -2327 671 -2325
rect 667 -2333 668 -2331
rect 670 -2333 671 -2331
rect 674 -2327 675 -2325
rect 674 -2333 675 -2331
rect 681 -2327 682 -2325
rect 681 -2333 682 -2331
rect 688 -2327 689 -2325
rect 688 -2333 689 -2331
rect 695 -2327 696 -2325
rect 695 -2333 696 -2331
rect 702 -2327 703 -2325
rect 705 -2327 706 -2325
rect 702 -2333 703 -2331
rect 709 -2327 710 -2325
rect 709 -2333 710 -2331
rect 716 -2327 717 -2325
rect 716 -2333 717 -2331
rect 723 -2327 724 -2325
rect 726 -2327 727 -2325
rect 723 -2333 724 -2331
rect 726 -2333 727 -2331
rect 730 -2327 731 -2325
rect 730 -2333 731 -2331
rect 737 -2327 738 -2325
rect 737 -2333 738 -2331
rect 744 -2327 745 -2325
rect 744 -2333 745 -2331
rect 751 -2327 752 -2325
rect 751 -2333 752 -2331
rect 758 -2327 759 -2325
rect 758 -2333 759 -2331
rect 765 -2327 766 -2325
rect 768 -2333 769 -2331
rect 772 -2327 773 -2325
rect 772 -2333 773 -2331
rect 779 -2327 780 -2325
rect 782 -2327 783 -2325
rect 782 -2333 783 -2331
rect 786 -2327 787 -2325
rect 786 -2333 787 -2331
rect 793 -2327 794 -2325
rect 793 -2333 794 -2331
rect 800 -2327 801 -2325
rect 800 -2333 801 -2331
rect 807 -2327 808 -2325
rect 807 -2333 808 -2331
rect 814 -2327 815 -2325
rect 814 -2333 815 -2331
rect 821 -2327 822 -2325
rect 821 -2333 822 -2331
rect 828 -2327 829 -2325
rect 828 -2333 829 -2331
rect 835 -2327 836 -2325
rect 835 -2333 836 -2331
rect 842 -2327 843 -2325
rect 842 -2333 843 -2331
rect 849 -2327 850 -2325
rect 849 -2333 850 -2331
rect 856 -2327 857 -2325
rect 859 -2327 860 -2325
rect 856 -2333 857 -2331
rect 859 -2333 860 -2331
rect 863 -2327 864 -2325
rect 863 -2333 864 -2331
rect 870 -2327 871 -2325
rect 870 -2333 871 -2331
rect 877 -2327 878 -2325
rect 877 -2333 878 -2331
rect 884 -2327 885 -2325
rect 884 -2333 885 -2331
rect 891 -2327 892 -2325
rect 891 -2333 892 -2331
rect 898 -2327 899 -2325
rect 898 -2333 899 -2331
rect 905 -2327 906 -2325
rect 905 -2333 906 -2331
rect 912 -2327 913 -2325
rect 912 -2333 913 -2331
rect 919 -2327 920 -2325
rect 919 -2333 920 -2331
rect 922 -2333 923 -2331
rect 926 -2327 927 -2325
rect 926 -2333 927 -2331
rect 936 -2327 937 -2325
rect 933 -2333 934 -2331
rect 936 -2333 937 -2331
rect 940 -2327 941 -2325
rect 940 -2333 941 -2331
rect 947 -2327 948 -2325
rect 947 -2333 948 -2331
rect 954 -2327 955 -2325
rect 954 -2333 955 -2331
rect 961 -2327 962 -2325
rect 961 -2333 962 -2331
rect 968 -2327 969 -2325
rect 968 -2333 969 -2331
rect 975 -2327 976 -2325
rect 978 -2327 979 -2325
rect 975 -2333 976 -2331
rect 978 -2333 979 -2331
rect 982 -2327 983 -2325
rect 982 -2333 983 -2331
rect 989 -2327 990 -2325
rect 992 -2327 993 -2325
rect 989 -2333 990 -2331
rect 992 -2333 993 -2331
rect 996 -2327 997 -2325
rect 996 -2333 997 -2331
rect 1003 -2327 1004 -2325
rect 1003 -2333 1004 -2331
rect 1010 -2327 1011 -2325
rect 1010 -2333 1011 -2331
rect 1017 -2327 1018 -2325
rect 1017 -2333 1018 -2331
rect 1024 -2327 1025 -2325
rect 1024 -2333 1025 -2331
rect 1031 -2327 1032 -2325
rect 1031 -2333 1032 -2331
rect 1041 -2327 1042 -2325
rect 1038 -2333 1039 -2331
rect 1041 -2333 1042 -2331
rect 1045 -2327 1046 -2325
rect 1045 -2333 1046 -2331
rect 1052 -2327 1053 -2325
rect 1052 -2333 1053 -2331
rect 1059 -2327 1060 -2325
rect 1059 -2333 1060 -2331
rect 1066 -2327 1067 -2325
rect 1066 -2333 1067 -2331
rect 1073 -2327 1074 -2325
rect 1073 -2333 1074 -2331
rect 1080 -2327 1081 -2325
rect 1080 -2333 1081 -2331
rect 1087 -2327 1088 -2325
rect 1087 -2333 1088 -2331
rect 1094 -2327 1095 -2325
rect 1094 -2333 1095 -2331
rect 1101 -2327 1102 -2325
rect 1101 -2333 1102 -2331
rect 1108 -2327 1109 -2325
rect 1108 -2333 1109 -2331
rect 1115 -2327 1116 -2325
rect 1115 -2333 1116 -2331
rect 1122 -2327 1123 -2325
rect 1122 -2333 1123 -2331
rect 1129 -2327 1130 -2325
rect 1129 -2333 1130 -2331
rect 1136 -2327 1137 -2325
rect 1139 -2327 1140 -2325
rect 1136 -2333 1137 -2331
rect 1139 -2333 1140 -2331
rect 1143 -2327 1144 -2325
rect 1143 -2333 1144 -2331
rect 1150 -2327 1151 -2325
rect 1150 -2333 1151 -2331
rect 1157 -2327 1158 -2325
rect 1157 -2333 1158 -2331
rect 1164 -2327 1165 -2325
rect 1164 -2333 1165 -2331
rect 1171 -2327 1172 -2325
rect 1171 -2333 1172 -2331
rect 1178 -2327 1179 -2325
rect 1178 -2333 1179 -2331
rect 1185 -2327 1186 -2325
rect 1185 -2333 1186 -2331
rect 1192 -2327 1193 -2325
rect 1192 -2333 1193 -2331
rect 1199 -2327 1200 -2325
rect 1199 -2333 1200 -2331
rect 1206 -2327 1207 -2325
rect 1206 -2333 1207 -2331
rect 1213 -2327 1214 -2325
rect 1213 -2333 1214 -2331
rect 1220 -2327 1221 -2325
rect 1220 -2333 1221 -2331
rect 1227 -2327 1228 -2325
rect 1227 -2333 1228 -2331
rect 1234 -2327 1235 -2325
rect 1234 -2333 1235 -2331
rect 1241 -2327 1242 -2325
rect 1241 -2333 1242 -2331
rect 1248 -2327 1249 -2325
rect 1248 -2333 1249 -2331
rect 1251 -2333 1252 -2331
rect 1255 -2327 1256 -2325
rect 1255 -2333 1256 -2331
rect 1262 -2327 1263 -2325
rect 1262 -2333 1263 -2331
rect 1269 -2327 1270 -2325
rect 1269 -2333 1270 -2331
rect 1276 -2327 1277 -2325
rect 1276 -2333 1277 -2331
rect 1283 -2327 1284 -2325
rect 1283 -2333 1284 -2331
rect 1290 -2327 1291 -2325
rect 1293 -2327 1294 -2325
rect 1290 -2333 1291 -2331
rect 1293 -2333 1294 -2331
rect 1297 -2327 1298 -2325
rect 1297 -2333 1298 -2331
rect 1304 -2327 1305 -2325
rect 1304 -2333 1305 -2331
rect 1311 -2327 1312 -2325
rect 1311 -2333 1312 -2331
rect 1318 -2327 1319 -2325
rect 1321 -2327 1322 -2325
rect 1318 -2333 1319 -2331
rect 1321 -2333 1322 -2331
rect 1325 -2327 1326 -2325
rect 1325 -2333 1326 -2331
rect 1332 -2327 1333 -2325
rect 1332 -2333 1333 -2331
rect 1339 -2327 1340 -2325
rect 1339 -2333 1340 -2331
rect 1346 -2327 1347 -2325
rect 1346 -2333 1347 -2331
rect 1353 -2327 1354 -2325
rect 1353 -2333 1354 -2331
rect 1360 -2327 1361 -2325
rect 1360 -2333 1361 -2331
rect 1367 -2327 1368 -2325
rect 1367 -2333 1368 -2331
rect 1374 -2327 1375 -2325
rect 1374 -2333 1375 -2331
rect 1381 -2327 1382 -2325
rect 1381 -2333 1382 -2331
rect 1388 -2327 1389 -2325
rect 1388 -2333 1389 -2331
rect 1395 -2327 1396 -2325
rect 1398 -2327 1399 -2325
rect 1398 -2333 1399 -2331
rect 1402 -2327 1403 -2325
rect 1402 -2333 1403 -2331
rect 1409 -2327 1410 -2325
rect 1409 -2333 1410 -2331
rect 1416 -2327 1417 -2325
rect 1416 -2333 1417 -2331
rect 1423 -2327 1424 -2325
rect 1423 -2333 1424 -2331
rect 1430 -2327 1431 -2325
rect 1430 -2333 1431 -2331
rect 1437 -2327 1438 -2325
rect 1437 -2333 1438 -2331
rect 1444 -2327 1445 -2325
rect 1444 -2333 1445 -2331
rect 1451 -2327 1452 -2325
rect 1451 -2333 1452 -2331
rect 1458 -2327 1459 -2325
rect 1458 -2333 1459 -2331
rect 1465 -2327 1466 -2325
rect 1465 -2333 1466 -2331
rect 1472 -2327 1473 -2325
rect 1472 -2333 1473 -2331
rect 1479 -2327 1480 -2325
rect 1479 -2333 1480 -2331
rect 1486 -2327 1487 -2325
rect 1486 -2333 1487 -2331
rect 1493 -2327 1494 -2325
rect 1496 -2327 1497 -2325
rect 1493 -2333 1494 -2331
rect 1496 -2333 1497 -2331
rect 1500 -2327 1501 -2325
rect 1503 -2327 1504 -2325
rect 1500 -2333 1501 -2331
rect 1507 -2327 1508 -2325
rect 1507 -2333 1508 -2331
rect 1514 -2327 1515 -2325
rect 1517 -2327 1518 -2325
rect 1517 -2333 1518 -2331
rect 1521 -2327 1522 -2325
rect 1521 -2333 1522 -2331
rect 1528 -2327 1529 -2325
rect 1528 -2333 1529 -2331
rect 1535 -2327 1536 -2325
rect 1535 -2333 1536 -2331
rect 1542 -2327 1543 -2325
rect 1545 -2327 1546 -2325
rect 1542 -2333 1543 -2331
rect 1545 -2333 1546 -2331
rect 1549 -2327 1550 -2325
rect 1549 -2333 1550 -2331
rect 1556 -2327 1557 -2325
rect 1556 -2333 1557 -2331
rect 1563 -2327 1564 -2325
rect 1563 -2333 1564 -2331
rect 1570 -2327 1571 -2325
rect 1570 -2333 1571 -2331
rect 1577 -2327 1578 -2325
rect 1577 -2333 1578 -2331
rect 1584 -2327 1585 -2325
rect 1584 -2333 1585 -2331
rect 1591 -2327 1592 -2325
rect 1591 -2333 1592 -2331
rect 1598 -2327 1599 -2325
rect 1598 -2333 1599 -2331
rect 1605 -2327 1606 -2325
rect 1605 -2333 1606 -2331
rect 1612 -2327 1613 -2325
rect 1612 -2333 1613 -2331
rect 1619 -2327 1620 -2325
rect 1619 -2333 1620 -2331
rect 1626 -2327 1627 -2325
rect 1629 -2327 1630 -2325
rect 1626 -2333 1627 -2331
rect 1629 -2333 1630 -2331
rect 1633 -2327 1634 -2325
rect 1633 -2333 1634 -2331
rect 1640 -2327 1641 -2325
rect 1640 -2333 1641 -2331
rect 1647 -2327 1648 -2325
rect 1647 -2333 1648 -2331
rect 1654 -2327 1655 -2325
rect 1654 -2333 1655 -2331
rect 1661 -2327 1662 -2325
rect 1661 -2333 1662 -2331
rect 1668 -2327 1669 -2325
rect 1668 -2333 1669 -2331
rect 1675 -2327 1676 -2325
rect 1675 -2333 1676 -2331
rect 1685 -2327 1686 -2325
rect 1682 -2333 1683 -2331
rect 1685 -2333 1686 -2331
rect 1689 -2327 1690 -2325
rect 1689 -2333 1690 -2331
rect 1696 -2327 1697 -2325
rect 1696 -2333 1697 -2331
rect 1703 -2327 1704 -2325
rect 1703 -2333 1704 -2331
rect 1710 -2327 1711 -2325
rect 1710 -2333 1711 -2331
rect 1717 -2327 1718 -2325
rect 1717 -2333 1718 -2331
rect 1724 -2327 1725 -2325
rect 1724 -2333 1725 -2331
rect 1731 -2327 1732 -2325
rect 1731 -2333 1732 -2331
rect 1738 -2327 1739 -2325
rect 1738 -2333 1739 -2331
rect 1745 -2327 1746 -2325
rect 1745 -2333 1746 -2331
rect 1752 -2327 1753 -2325
rect 1752 -2333 1753 -2331
rect 1759 -2327 1760 -2325
rect 1759 -2333 1760 -2331
rect 1766 -2327 1767 -2325
rect 1766 -2333 1767 -2331
rect 1773 -2327 1774 -2325
rect 1773 -2333 1774 -2331
rect 1780 -2327 1781 -2325
rect 1780 -2333 1781 -2331
rect 1787 -2327 1788 -2325
rect 1787 -2333 1788 -2331
rect 1794 -2327 1795 -2325
rect 1794 -2333 1795 -2331
rect 1801 -2327 1802 -2325
rect 1801 -2333 1802 -2331
rect 1808 -2327 1809 -2325
rect 1808 -2333 1809 -2331
rect 1815 -2327 1816 -2325
rect 1815 -2333 1816 -2331
rect 1822 -2327 1823 -2325
rect 1822 -2333 1823 -2331
rect 1829 -2327 1830 -2325
rect 1829 -2333 1830 -2331
rect 1836 -2327 1837 -2325
rect 1836 -2333 1837 -2331
rect 1843 -2327 1844 -2325
rect 1843 -2333 1844 -2331
rect 1850 -2327 1851 -2325
rect 1850 -2333 1851 -2331
rect 1853 -2333 1854 -2331
rect 1857 -2327 1858 -2325
rect 1857 -2333 1858 -2331
rect 1864 -2327 1865 -2325
rect 1864 -2333 1865 -2331
rect 1871 -2327 1872 -2325
rect 1871 -2333 1872 -2331
rect 1878 -2327 1879 -2325
rect 1878 -2333 1879 -2331
rect 1885 -2327 1886 -2325
rect 1885 -2333 1886 -2331
rect 1895 -2327 1896 -2325
rect 1895 -2333 1896 -2331
rect 1899 -2327 1900 -2325
rect 1899 -2333 1900 -2331
rect 1906 -2327 1907 -2325
rect 1906 -2333 1907 -2331
rect 1913 -2327 1914 -2325
rect 1913 -2333 1914 -2331
rect 1920 -2327 1921 -2325
rect 1920 -2333 1921 -2331
rect 1927 -2327 1928 -2325
rect 1927 -2333 1928 -2331
rect 1934 -2327 1935 -2325
rect 1937 -2327 1938 -2325
rect 1934 -2333 1935 -2331
rect 1937 -2333 1938 -2331
rect 1941 -2327 1942 -2325
rect 1941 -2333 1942 -2331
rect 1948 -2327 1949 -2325
rect 1948 -2333 1949 -2331
rect 1955 -2327 1956 -2325
rect 1955 -2333 1956 -2331
rect 1962 -2327 1963 -2325
rect 1962 -2333 1963 -2331
rect 1969 -2327 1970 -2325
rect 1969 -2333 1970 -2331
rect 1976 -2327 1977 -2325
rect 1979 -2327 1980 -2325
rect 1979 -2333 1980 -2331
rect 1983 -2327 1984 -2325
rect 1983 -2333 1984 -2331
rect 1990 -2327 1991 -2325
rect 1990 -2333 1991 -2331
rect 1997 -2327 1998 -2325
rect 1997 -2333 1998 -2331
rect 2004 -2327 2005 -2325
rect 2004 -2333 2005 -2331
rect 2011 -2327 2012 -2325
rect 2011 -2333 2012 -2331
rect 2018 -2327 2019 -2325
rect 2018 -2333 2019 -2331
rect 2025 -2327 2026 -2325
rect 2025 -2333 2026 -2331
rect 2032 -2327 2033 -2325
rect 2032 -2333 2033 -2331
rect 2039 -2327 2040 -2325
rect 2039 -2333 2040 -2331
rect 2046 -2327 2047 -2325
rect 2046 -2333 2047 -2331
rect 2053 -2327 2054 -2325
rect 2053 -2333 2054 -2331
rect 2060 -2327 2061 -2325
rect 2060 -2333 2061 -2331
rect 2067 -2327 2068 -2325
rect 2067 -2333 2068 -2331
rect 2074 -2327 2075 -2325
rect 2074 -2333 2075 -2331
rect 2081 -2327 2082 -2325
rect 2081 -2333 2082 -2331
rect 2088 -2327 2089 -2325
rect 2088 -2333 2089 -2331
rect 2095 -2327 2096 -2325
rect 2095 -2333 2096 -2331
rect 2102 -2327 2103 -2325
rect 2102 -2333 2103 -2331
rect 2109 -2327 2110 -2325
rect 2109 -2333 2110 -2331
rect 2116 -2327 2117 -2325
rect 2116 -2333 2117 -2331
rect 2123 -2327 2124 -2325
rect 2123 -2333 2124 -2331
rect 2130 -2327 2131 -2325
rect 2130 -2333 2131 -2331
rect 2137 -2327 2138 -2325
rect 2137 -2333 2138 -2331
rect 2144 -2327 2145 -2325
rect 2144 -2333 2145 -2331
rect 2151 -2327 2152 -2325
rect 2151 -2333 2152 -2331
rect 2158 -2327 2159 -2325
rect 2158 -2333 2159 -2331
rect 2165 -2327 2166 -2325
rect 2165 -2333 2166 -2331
rect 2172 -2327 2173 -2325
rect 2172 -2333 2173 -2331
rect 2179 -2327 2180 -2325
rect 2179 -2333 2180 -2331
rect 2186 -2327 2187 -2325
rect 2186 -2333 2187 -2331
rect 2193 -2327 2194 -2325
rect 2193 -2333 2194 -2331
rect 2200 -2327 2201 -2325
rect 2200 -2333 2201 -2331
rect 2207 -2327 2208 -2325
rect 2207 -2333 2208 -2331
rect 2214 -2327 2215 -2325
rect 2214 -2333 2215 -2331
rect 2221 -2327 2222 -2325
rect 2221 -2333 2222 -2331
rect 2228 -2327 2229 -2325
rect 2228 -2333 2229 -2331
rect 2235 -2327 2236 -2325
rect 2235 -2333 2236 -2331
rect 2242 -2327 2243 -2325
rect 2242 -2333 2243 -2331
rect 2249 -2327 2250 -2325
rect 2249 -2333 2250 -2331
rect 2256 -2327 2257 -2325
rect 2256 -2333 2257 -2331
rect 2263 -2327 2264 -2325
rect 2263 -2333 2264 -2331
rect 2270 -2327 2271 -2325
rect 2270 -2333 2271 -2331
rect 2277 -2327 2278 -2325
rect 2277 -2333 2278 -2331
rect 2284 -2327 2285 -2325
rect 2284 -2333 2285 -2331
rect 2291 -2327 2292 -2325
rect 2291 -2333 2292 -2331
rect 2298 -2327 2299 -2325
rect 2298 -2333 2299 -2331
rect 2305 -2327 2306 -2325
rect 2305 -2333 2306 -2331
rect 2312 -2327 2313 -2325
rect 2312 -2333 2313 -2331
rect 2319 -2327 2320 -2325
rect 2319 -2333 2320 -2331
rect 2326 -2327 2327 -2325
rect 2326 -2333 2327 -2331
rect 2333 -2327 2334 -2325
rect 2336 -2327 2337 -2325
rect 2333 -2333 2334 -2331
rect 2336 -2333 2337 -2331
rect 2343 -2327 2344 -2325
rect 2343 -2333 2344 -2331
rect 2347 -2327 2348 -2325
rect 2347 -2333 2348 -2331
rect 2 -2500 3 -2498
rect 5 -2500 6 -2498
rect 5 -2506 6 -2504
rect 9 -2500 10 -2498
rect 9 -2506 10 -2504
rect 16 -2500 17 -2498
rect 19 -2506 20 -2504
rect 23 -2500 24 -2498
rect 23 -2506 24 -2504
rect 30 -2506 31 -2504
rect 33 -2506 34 -2504
rect 37 -2500 38 -2498
rect 37 -2506 38 -2504
rect 40 -2506 41 -2504
rect 44 -2500 45 -2498
rect 44 -2506 45 -2504
rect 51 -2500 52 -2498
rect 51 -2506 52 -2504
rect 58 -2500 59 -2498
rect 58 -2506 59 -2504
rect 61 -2506 62 -2504
rect 65 -2500 66 -2498
rect 65 -2506 66 -2504
rect 72 -2500 73 -2498
rect 72 -2506 73 -2504
rect 79 -2500 80 -2498
rect 79 -2506 80 -2504
rect 86 -2500 87 -2498
rect 86 -2506 87 -2504
rect 93 -2500 94 -2498
rect 96 -2500 97 -2498
rect 93 -2506 94 -2504
rect 96 -2506 97 -2504
rect 100 -2500 101 -2498
rect 100 -2506 101 -2504
rect 107 -2500 108 -2498
rect 110 -2500 111 -2498
rect 110 -2506 111 -2504
rect 114 -2500 115 -2498
rect 114 -2506 115 -2504
rect 121 -2500 122 -2498
rect 121 -2506 122 -2504
rect 128 -2500 129 -2498
rect 128 -2506 129 -2504
rect 135 -2500 136 -2498
rect 135 -2506 136 -2504
rect 142 -2500 143 -2498
rect 142 -2506 143 -2504
rect 149 -2500 150 -2498
rect 149 -2506 150 -2504
rect 156 -2500 157 -2498
rect 156 -2506 157 -2504
rect 163 -2500 164 -2498
rect 163 -2506 164 -2504
rect 166 -2506 167 -2504
rect 170 -2500 171 -2498
rect 170 -2506 171 -2504
rect 177 -2506 178 -2504
rect 184 -2500 185 -2498
rect 184 -2506 185 -2504
rect 191 -2500 192 -2498
rect 191 -2506 192 -2504
rect 198 -2500 199 -2498
rect 198 -2506 199 -2504
rect 205 -2500 206 -2498
rect 205 -2506 206 -2504
rect 212 -2500 213 -2498
rect 212 -2506 213 -2504
rect 219 -2500 220 -2498
rect 219 -2506 220 -2504
rect 226 -2500 227 -2498
rect 226 -2506 227 -2504
rect 233 -2500 234 -2498
rect 233 -2506 234 -2504
rect 240 -2500 241 -2498
rect 240 -2506 241 -2504
rect 247 -2500 248 -2498
rect 247 -2506 248 -2504
rect 254 -2500 255 -2498
rect 254 -2506 255 -2504
rect 261 -2500 262 -2498
rect 261 -2506 262 -2504
rect 268 -2500 269 -2498
rect 268 -2506 269 -2504
rect 275 -2500 276 -2498
rect 275 -2506 276 -2504
rect 282 -2500 283 -2498
rect 282 -2506 283 -2504
rect 289 -2500 290 -2498
rect 289 -2506 290 -2504
rect 296 -2500 297 -2498
rect 296 -2506 297 -2504
rect 303 -2500 304 -2498
rect 303 -2506 304 -2504
rect 310 -2500 311 -2498
rect 310 -2506 311 -2504
rect 317 -2500 318 -2498
rect 317 -2506 318 -2504
rect 324 -2500 325 -2498
rect 324 -2506 325 -2504
rect 331 -2500 332 -2498
rect 331 -2506 332 -2504
rect 338 -2500 339 -2498
rect 338 -2506 339 -2504
rect 345 -2500 346 -2498
rect 345 -2506 346 -2504
rect 352 -2500 353 -2498
rect 352 -2506 353 -2504
rect 359 -2500 360 -2498
rect 359 -2506 360 -2504
rect 366 -2500 367 -2498
rect 366 -2506 367 -2504
rect 373 -2500 374 -2498
rect 373 -2506 374 -2504
rect 380 -2500 381 -2498
rect 380 -2506 381 -2504
rect 387 -2500 388 -2498
rect 387 -2506 388 -2504
rect 394 -2500 395 -2498
rect 394 -2506 395 -2504
rect 401 -2500 402 -2498
rect 401 -2506 402 -2504
rect 408 -2500 409 -2498
rect 408 -2506 409 -2504
rect 415 -2500 416 -2498
rect 415 -2506 416 -2504
rect 422 -2500 423 -2498
rect 422 -2506 423 -2504
rect 429 -2500 430 -2498
rect 429 -2506 430 -2504
rect 436 -2500 437 -2498
rect 436 -2506 437 -2504
rect 443 -2500 444 -2498
rect 443 -2506 444 -2504
rect 450 -2500 451 -2498
rect 450 -2506 451 -2504
rect 457 -2500 458 -2498
rect 457 -2506 458 -2504
rect 464 -2500 465 -2498
rect 464 -2506 465 -2504
rect 471 -2500 472 -2498
rect 471 -2506 472 -2504
rect 478 -2500 479 -2498
rect 481 -2500 482 -2498
rect 478 -2506 479 -2504
rect 481 -2506 482 -2504
rect 485 -2500 486 -2498
rect 485 -2506 486 -2504
rect 492 -2500 493 -2498
rect 492 -2506 493 -2504
rect 499 -2500 500 -2498
rect 499 -2506 500 -2504
rect 506 -2500 507 -2498
rect 506 -2506 507 -2504
rect 513 -2500 514 -2498
rect 513 -2506 514 -2504
rect 520 -2500 521 -2498
rect 520 -2506 521 -2504
rect 527 -2500 528 -2498
rect 527 -2506 528 -2504
rect 534 -2500 535 -2498
rect 534 -2506 535 -2504
rect 541 -2500 542 -2498
rect 541 -2506 542 -2504
rect 548 -2500 549 -2498
rect 548 -2506 549 -2504
rect 555 -2500 556 -2498
rect 555 -2506 556 -2504
rect 562 -2500 563 -2498
rect 562 -2506 563 -2504
rect 569 -2500 570 -2498
rect 569 -2506 570 -2504
rect 576 -2500 577 -2498
rect 576 -2506 577 -2504
rect 583 -2500 584 -2498
rect 583 -2506 584 -2504
rect 590 -2500 591 -2498
rect 590 -2506 591 -2504
rect 597 -2500 598 -2498
rect 597 -2506 598 -2504
rect 604 -2500 605 -2498
rect 607 -2500 608 -2498
rect 607 -2506 608 -2504
rect 611 -2500 612 -2498
rect 611 -2506 612 -2504
rect 618 -2500 619 -2498
rect 618 -2506 619 -2504
rect 625 -2500 626 -2498
rect 625 -2506 626 -2504
rect 632 -2500 633 -2498
rect 632 -2506 633 -2504
rect 639 -2500 640 -2498
rect 639 -2506 640 -2504
rect 646 -2500 647 -2498
rect 646 -2506 647 -2504
rect 653 -2500 654 -2498
rect 653 -2506 654 -2504
rect 660 -2500 661 -2498
rect 660 -2506 661 -2504
rect 667 -2500 668 -2498
rect 670 -2500 671 -2498
rect 667 -2506 668 -2504
rect 670 -2506 671 -2504
rect 674 -2500 675 -2498
rect 674 -2506 675 -2504
rect 681 -2500 682 -2498
rect 681 -2506 682 -2504
rect 688 -2500 689 -2498
rect 688 -2506 689 -2504
rect 695 -2500 696 -2498
rect 695 -2506 696 -2504
rect 702 -2500 703 -2498
rect 702 -2506 703 -2504
rect 709 -2500 710 -2498
rect 709 -2506 710 -2504
rect 716 -2500 717 -2498
rect 716 -2506 717 -2504
rect 723 -2500 724 -2498
rect 723 -2506 724 -2504
rect 730 -2500 731 -2498
rect 730 -2506 731 -2504
rect 737 -2500 738 -2498
rect 740 -2500 741 -2498
rect 737 -2506 738 -2504
rect 740 -2506 741 -2504
rect 744 -2500 745 -2498
rect 744 -2506 745 -2504
rect 751 -2500 752 -2498
rect 751 -2506 752 -2504
rect 758 -2500 759 -2498
rect 758 -2506 759 -2504
rect 765 -2500 766 -2498
rect 765 -2506 766 -2504
rect 772 -2500 773 -2498
rect 775 -2500 776 -2498
rect 775 -2506 776 -2504
rect 779 -2500 780 -2498
rect 779 -2506 780 -2504
rect 786 -2500 787 -2498
rect 786 -2506 787 -2504
rect 793 -2500 794 -2498
rect 796 -2500 797 -2498
rect 793 -2506 794 -2504
rect 796 -2506 797 -2504
rect 800 -2500 801 -2498
rect 800 -2506 801 -2504
rect 807 -2500 808 -2498
rect 807 -2506 808 -2504
rect 814 -2500 815 -2498
rect 814 -2506 815 -2504
rect 821 -2500 822 -2498
rect 821 -2506 822 -2504
rect 828 -2500 829 -2498
rect 828 -2506 829 -2504
rect 835 -2500 836 -2498
rect 835 -2506 836 -2504
rect 842 -2500 843 -2498
rect 842 -2506 843 -2504
rect 849 -2500 850 -2498
rect 849 -2506 850 -2504
rect 856 -2500 857 -2498
rect 859 -2500 860 -2498
rect 856 -2506 857 -2504
rect 859 -2506 860 -2504
rect 863 -2500 864 -2498
rect 863 -2506 864 -2504
rect 870 -2500 871 -2498
rect 873 -2500 874 -2498
rect 873 -2506 874 -2504
rect 877 -2500 878 -2498
rect 877 -2506 878 -2504
rect 884 -2500 885 -2498
rect 884 -2506 885 -2504
rect 891 -2500 892 -2498
rect 891 -2506 892 -2504
rect 898 -2500 899 -2498
rect 898 -2506 899 -2504
rect 905 -2500 906 -2498
rect 905 -2506 906 -2504
rect 912 -2500 913 -2498
rect 912 -2506 913 -2504
rect 919 -2500 920 -2498
rect 922 -2500 923 -2498
rect 919 -2506 920 -2504
rect 922 -2506 923 -2504
rect 926 -2500 927 -2498
rect 926 -2506 927 -2504
rect 933 -2500 934 -2498
rect 933 -2506 934 -2504
rect 940 -2500 941 -2498
rect 940 -2506 941 -2504
rect 947 -2500 948 -2498
rect 947 -2506 948 -2504
rect 954 -2500 955 -2498
rect 957 -2500 958 -2498
rect 954 -2506 955 -2504
rect 957 -2506 958 -2504
rect 961 -2500 962 -2498
rect 961 -2506 962 -2504
rect 968 -2500 969 -2498
rect 968 -2506 969 -2504
rect 975 -2500 976 -2498
rect 978 -2500 979 -2498
rect 975 -2506 976 -2504
rect 978 -2506 979 -2504
rect 982 -2500 983 -2498
rect 982 -2506 983 -2504
rect 992 -2500 993 -2498
rect 989 -2506 990 -2504
rect 992 -2506 993 -2504
rect 996 -2500 997 -2498
rect 996 -2506 997 -2504
rect 1003 -2500 1004 -2498
rect 1003 -2506 1004 -2504
rect 1010 -2500 1011 -2498
rect 1013 -2500 1014 -2498
rect 1010 -2506 1011 -2504
rect 1013 -2506 1014 -2504
rect 1017 -2500 1018 -2498
rect 1017 -2506 1018 -2504
rect 1024 -2500 1025 -2498
rect 1024 -2506 1025 -2504
rect 1031 -2500 1032 -2498
rect 1031 -2506 1032 -2504
rect 1038 -2500 1039 -2498
rect 1038 -2506 1039 -2504
rect 1045 -2500 1046 -2498
rect 1045 -2506 1046 -2504
rect 1052 -2500 1053 -2498
rect 1055 -2500 1056 -2498
rect 1052 -2506 1053 -2504
rect 1055 -2506 1056 -2504
rect 1059 -2500 1060 -2498
rect 1059 -2506 1060 -2504
rect 1066 -2500 1067 -2498
rect 1066 -2506 1067 -2504
rect 1073 -2500 1074 -2498
rect 1076 -2500 1077 -2498
rect 1073 -2506 1074 -2504
rect 1080 -2500 1081 -2498
rect 1083 -2500 1084 -2498
rect 1080 -2506 1081 -2504
rect 1083 -2506 1084 -2504
rect 1087 -2500 1088 -2498
rect 1087 -2506 1088 -2504
rect 1094 -2500 1095 -2498
rect 1094 -2506 1095 -2504
rect 1101 -2500 1102 -2498
rect 1101 -2506 1102 -2504
rect 1108 -2500 1109 -2498
rect 1108 -2506 1109 -2504
rect 1115 -2500 1116 -2498
rect 1115 -2506 1116 -2504
rect 1122 -2500 1123 -2498
rect 1122 -2506 1123 -2504
rect 1129 -2500 1130 -2498
rect 1129 -2506 1130 -2504
rect 1136 -2500 1137 -2498
rect 1136 -2506 1137 -2504
rect 1143 -2500 1144 -2498
rect 1143 -2506 1144 -2504
rect 1150 -2500 1151 -2498
rect 1150 -2506 1151 -2504
rect 1157 -2500 1158 -2498
rect 1157 -2506 1158 -2504
rect 1164 -2500 1165 -2498
rect 1164 -2506 1165 -2504
rect 1171 -2500 1172 -2498
rect 1174 -2500 1175 -2498
rect 1171 -2506 1172 -2504
rect 1174 -2506 1175 -2504
rect 1178 -2500 1179 -2498
rect 1178 -2506 1179 -2504
rect 1185 -2500 1186 -2498
rect 1185 -2506 1186 -2504
rect 1192 -2500 1193 -2498
rect 1192 -2506 1193 -2504
rect 1199 -2500 1200 -2498
rect 1199 -2506 1200 -2504
rect 1206 -2500 1207 -2498
rect 1206 -2506 1207 -2504
rect 1213 -2500 1214 -2498
rect 1213 -2506 1214 -2504
rect 1216 -2506 1217 -2504
rect 1220 -2500 1221 -2498
rect 1220 -2506 1221 -2504
rect 1227 -2500 1228 -2498
rect 1227 -2506 1228 -2504
rect 1234 -2500 1235 -2498
rect 1234 -2506 1235 -2504
rect 1241 -2500 1242 -2498
rect 1241 -2506 1242 -2504
rect 1248 -2500 1249 -2498
rect 1248 -2506 1249 -2504
rect 1255 -2500 1256 -2498
rect 1255 -2506 1256 -2504
rect 1262 -2500 1263 -2498
rect 1262 -2506 1263 -2504
rect 1269 -2500 1270 -2498
rect 1272 -2500 1273 -2498
rect 1269 -2506 1270 -2504
rect 1272 -2506 1273 -2504
rect 1276 -2500 1277 -2498
rect 1276 -2506 1277 -2504
rect 1283 -2500 1284 -2498
rect 1283 -2506 1284 -2504
rect 1290 -2506 1291 -2504
rect 1297 -2500 1298 -2498
rect 1297 -2506 1298 -2504
rect 1304 -2500 1305 -2498
rect 1304 -2506 1305 -2504
rect 1311 -2500 1312 -2498
rect 1311 -2506 1312 -2504
rect 1318 -2500 1319 -2498
rect 1318 -2506 1319 -2504
rect 1325 -2500 1326 -2498
rect 1325 -2506 1326 -2504
rect 1332 -2500 1333 -2498
rect 1335 -2500 1336 -2498
rect 1332 -2506 1333 -2504
rect 1335 -2506 1336 -2504
rect 1339 -2500 1340 -2498
rect 1339 -2506 1340 -2504
rect 1346 -2500 1347 -2498
rect 1346 -2506 1347 -2504
rect 1353 -2500 1354 -2498
rect 1356 -2500 1357 -2498
rect 1353 -2506 1354 -2504
rect 1356 -2506 1357 -2504
rect 1363 -2500 1364 -2498
rect 1360 -2506 1361 -2504
rect 1363 -2506 1364 -2504
rect 1367 -2500 1368 -2498
rect 1367 -2506 1368 -2504
rect 1374 -2500 1375 -2498
rect 1377 -2500 1378 -2498
rect 1374 -2506 1375 -2504
rect 1377 -2506 1378 -2504
rect 1381 -2500 1382 -2498
rect 1381 -2506 1382 -2504
rect 1388 -2500 1389 -2498
rect 1388 -2506 1389 -2504
rect 1395 -2500 1396 -2498
rect 1395 -2506 1396 -2504
rect 1402 -2500 1403 -2498
rect 1402 -2506 1403 -2504
rect 1409 -2500 1410 -2498
rect 1409 -2506 1410 -2504
rect 1416 -2500 1417 -2498
rect 1416 -2506 1417 -2504
rect 1423 -2500 1424 -2498
rect 1423 -2506 1424 -2504
rect 1430 -2500 1431 -2498
rect 1430 -2506 1431 -2504
rect 1437 -2500 1438 -2498
rect 1437 -2506 1438 -2504
rect 1444 -2500 1445 -2498
rect 1444 -2506 1445 -2504
rect 1451 -2500 1452 -2498
rect 1451 -2506 1452 -2504
rect 1458 -2500 1459 -2498
rect 1458 -2506 1459 -2504
rect 1465 -2500 1466 -2498
rect 1465 -2506 1466 -2504
rect 1472 -2500 1473 -2498
rect 1472 -2506 1473 -2504
rect 1479 -2500 1480 -2498
rect 1479 -2506 1480 -2504
rect 1486 -2500 1487 -2498
rect 1486 -2506 1487 -2504
rect 1493 -2500 1494 -2498
rect 1493 -2506 1494 -2504
rect 1500 -2500 1501 -2498
rect 1500 -2506 1501 -2504
rect 1507 -2500 1508 -2498
rect 1507 -2506 1508 -2504
rect 1514 -2500 1515 -2498
rect 1514 -2506 1515 -2504
rect 1521 -2500 1522 -2498
rect 1521 -2506 1522 -2504
rect 1528 -2500 1529 -2498
rect 1528 -2506 1529 -2504
rect 1535 -2500 1536 -2498
rect 1535 -2506 1536 -2504
rect 1542 -2500 1543 -2498
rect 1542 -2506 1543 -2504
rect 1549 -2500 1550 -2498
rect 1549 -2506 1550 -2504
rect 1556 -2500 1557 -2498
rect 1556 -2506 1557 -2504
rect 1563 -2500 1564 -2498
rect 1563 -2506 1564 -2504
rect 1570 -2500 1571 -2498
rect 1570 -2506 1571 -2504
rect 1577 -2500 1578 -2498
rect 1580 -2500 1581 -2498
rect 1577 -2506 1578 -2504
rect 1580 -2506 1581 -2504
rect 1584 -2500 1585 -2498
rect 1584 -2506 1585 -2504
rect 1591 -2500 1592 -2498
rect 1591 -2506 1592 -2504
rect 1598 -2500 1599 -2498
rect 1601 -2500 1602 -2498
rect 1598 -2506 1599 -2504
rect 1601 -2506 1602 -2504
rect 1605 -2500 1606 -2498
rect 1605 -2506 1606 -2504
rect 1612 -2500 1613 -2498
rect 1612 -2506 1613 -2504
rect 1619 -2500 1620 -2498
rect 1619 -2506 1620 -2504
rect 1626 -2500 1627 -2498
rect 1626 -2506 1627 -2504
rect 1633 -2500 1634 -2498
rect 1633 -2506 1634 -2504
rect 1640 -2500 1641 -2498
rect 1640 -2506 1641 -2504
rect 1647 -2500 1648 -2498
rect 1647 -2506 1648 -2504
rect 1654 -2500 1655 -2498
rect 1654 -2506 1655 -2504
rect 1661 -2500 1662 -2498
rect 1661 -2506 1662 -2504
rect 1668 -2500 1669 -2498
rect 1668 -2506 1669 -2504
rect 1678 -2500 1679 -2498
rect 1678 -2506 1679 -2504
rect 1682 -2500 1683 -2498
rect 1682 -2506 1683 -2504
rect 1689 -2500 1690 -2498
rect 1689 -2506 1690 -2504
rect 1696 -2500 1697 -2498
rect 1696 -2506 1697 -2504
rect 1703 -2500 1704 -2498
rect 1703 -2506 1704 -2504
rect 1710 -2500 1711 -2498
rect 1710 -2506 1711 -2504
rect 1717 -2500 1718 -2498
rect 1717 -2506 1718 -2504
rect 1724 -2500 1725 -2498
rect 1724 -2506 1725 -2504
rect 1731 -2500 1732 -2498
rect 1731 -2506 1732 -2504
rect 1738 -2500 1739 -2498
rect 1738 -2506 1739 -2504
rect 1745 -2500 1746 -2498
rect 1745 -2506 1746 -2504
rect 1752 -2500 1753 -2498
rect 1752 -2506 1753 -2504
rect 1759 -2500 1760 -2498
rect 1759 -2506 1760 -2504
rect 1766 -2500 1767 -2498
rect 1766 -2506 1767 -2504
rect 1773 -2500 1774 -2498
rect 1773 -2506 1774 -2504
rect 1780 -2500 1781 -2498
rect 1780 -2506 1781 -2504
rect 1787 -2500 1788 -2498
rect 1787 -2506 1788 -2504
rect 1794 -2500 1795 -2498
rect 1794 -2506 1795 -2504
rect 1801 -2500 1802 -2498
rect 1804 -2500 1805 -2498
rect 1804 -2506 1805 -2504
rect 1808 -2500 1809 -2498
rect 1808 -2506 1809 -2504
rect 1815 -2500 1816 -2498
rect 1815 -2506 1816 -2504
rect 1822 -2500 1823 -2498
rect 1822 -2506 1823 -2504
rect 1829 -2500 1830 -2498
rect 1829 -2506 1830 -2504
rect 1836 -2500 1837 -2498
rect 1836 -2506 1837 -2504
rect 1843 -2500 1844 -2498
rect 1843 -2506 1844 -2504
rect 1850 -2500 1851 -2498
rect 1853 -2500 1854 -2498
rect 1850 -2506 1851 -2504
rect 1857 -2500 1858 -2498
rect 1857 -2506 1858 -2504
rect 1864 -2500 1865 -2498
rect 1864 -2506 1865 -2504
rect 1871 -2500 1872 -2498
rect 1871 -2506 1872 -2504
rect 1878 -2500 1879 -2498
rect 1878 -2506 1879 -2504
rect 1885 -2500 1886 -2498
rect 1885 -2506 1886 -2504
rect 1892 -2500 1893 -2498
rect 1892 -2506 1893 -2504
rect 1899 -2500 1900 -2498
rect 1899 -2506 1900 -2504
rect 1906 -2500 1907 -2498
rect 1906 -2506 1907 -2504
rect 1913 -2500 1914 -2498
rect 1913 -2506 1914 -2504
rect 1920 -2500 1921 -2498
rect 1920 -2506 1921 -2504
rect 1927 -2500 1928 -2498
rect 1927 -2506 1928 -2504
rect 1934 -2500 1935 -2498
rect 1934 -2506 1935 -2504
rect 1941 -2500 1942 -2498
rect 1941 -2506 1942 -2504
rect 1948 -2500 1949 -2498
rect 1948 -2506 1949 -2504
rect 1955 -2500 1956 -2498
rect 1955 -2506 1956 -2504
rect 1962 -2500 1963 -2498
rect 1962 -2506 1963 -2504
rect 1969 -2500 1970 -2498
rect 1969 -2506 1970 -2504
rect 1976 -2500 1977 -2498
rect 1976 -2506 1977 -2504
rect 1983 -2500 1984 -2498
rect 1983 -2506 1984 -2504
rect 1990 -2500 1991 -2498
rect 1990 -2506 1991 -2504
rect 1997 -2500 1998 -2498
rect 1997 -2506 1998 -2504
rect 2004 -2500 2005 -2498
rect 2004 -2506 2005 -2504
rect 2011 -2500 2012 -2498
rect 2011 -2506 2012 -2504
rect 2018 -2500 2019 -2498
rect 2018 -2506 2019 -2504
rect 2025 -2500 2026 -2498
rect 2025 -2506 2026 -2504
rect 2032 -2500 2033 -2498
rect 2032 -2506 2033 -2504
rect 2039 -2500 2040 -2498
rect 2039 -2506 2040 -2504
rect 2046 -2500 2047 -2498
rect 2046 -2506 2047 -2504
rect 2053 -2500 2054 -2498
rect 2053 -2506 2054 -2504
rect 2060 -2500 2061 -2498
rect 2060 -2506 2061 -2504
rect 2067 -2500 2068 -2498
rect 2067 -2506 2068 -2504
rect 2074 -2500 2075 -2498
rect 2074 -2506 2075 -2504
rect 2081 -2500 2082 -2498
rect 2081 -2506 2082 -2504
rect 2088 -2500 2089 -2498
rect 2088 -2506 2089 -2504
rect 2095 -2500 2096 -2498
rect 2095 -2506 2096 -2504
rect 2102 -2500 2103 -2498
rect 2102 -2506 2103 -2504
rect 2109 -2500 2110 -2498
rect 2109 -2506 2110 -2504
rect 2116 -2500 2117 -2498
rect 2116 -2506 2117 -2504
rect 2123 -2500 2124 -2498
rect 2123 -2506 2124 -2504
rect 2130 -2500 2131 -2498
rect 2130 -2506 2131 -2504
rect 2137 -2500 2138 -2498
rect 2137 -2506 2138 -2504
rect 2144 -2500 2145 -2498
rect 2144 -2506 2145 -2504
rect 2151 -2500 2152 -2498
rect 2151 -2506 2152 -2504
rect 2158 -2500 2159 -2498
rect 2158 -2506 2159 -2504
rect 2165 -2500 2166 -2498
rect 2165 -2506 2166 -2504
rect 2172 -2500 2173 -2498
rect 2172 -2506 2173 -2504
rect 2179 -2500 2180 -2498
rect 2179 -2506 2180 -2504
rect 2186 -2500 2187 -2498
rect 2186 -2506 2187 -2504
rect 2193 -2500 2194 -2498
rect 2193 -2506 2194 -2504
rect 2200 -2500 2201 -2498
rect 2200 -2506 2201 -2504
rect 2207 -2500 2208 -2498
rect 2207 -2506 2208 -2504
rect 2214 -2500 2215 -2498
rect 2214 -2506 2215 -2504
rect 2221 -2500 2222 -2498
rect 2221 -2506 2222 -2504
rect 2228 -2500 2229 -2498
rect 2228 -2506 2229 -2504
rect 2235 -2500 2236 -2498
rect 2235 -2506 2236 -2504
rect 2242 -2500 2243 -2498
rect 2242 -2506 2243 -2504
rect 2249 -2500 2250 -2498
rect 2249 -2506 2250 -2504
rect 2256 -2500 2257 -2498
rect 2256 -2506 2257 -2504
rect 2263 -2500 2264 -2498
rect 2263 -2506 2264 -2504
rect 2270 -2500 2271 -2498
rect 2270 -2506 2271 -2504
rect 2280 -2500 2281 -2498
rect 2280 -2506 2281 -2504
rect 2284 -2500 2285 -2498
rect 2284 -2506 2285 -2504
rect 2291 -2500 2292 -2498
rect 2291 -2506 2292 -2504
rect 2298 -2500 2299 -2498
rect 2298 -2506 2299 -2504
rect 2305 -2500 2306 -2498
rect 2305 -2506 2306 -2504
rect 2312 -2500 2313 -2498
rect 2312 -2506 2313 -2504
rect 9 -2673 10 -2671
rect 9 -2679 10 -2677
rect 16 -2673 17 -2671
rect 16 -2679 17 -2677
rect 26 -2673 27 -2671
rect 23 -2679 24 -2677
rect 26 -2679 27 -2677
rect 30 -2673 31 -2671
rect 30 -2679 31 -2677
rect 37 -2673 38 -2671
rect 37 -2679 38 -2677
rect 44 -2673 45 -2671
rect 44 -2679 45 -2677
rect 51 -2673 52 -2671
rect 54 -2673 55 -2671
rect 51 -2679 52 -2677
rect 54 -2679 55 -2677
rect 58 -2673 59 -2671
rect 58 -2679 59 -2677
rect 65 -2673 66 -2671
rect 68 -2673 69 -2671
rect 65 -2679 66 -2677
rect 68 -2679 69 -2677
rect 72 -2673 73 -2671
rect 75 -2673 76 -2671
rect 72 -2679 73 -2677
rect 75 -2679 76 -2677
rect 79 -2673 80 -2671
rect 79 -2679 80 -2677
rect 86 -2673 87 -2671
rect 86 -2679 87 -2677
rect 93 -2673 94 -2671
rect 93 -2679 94 -2677
rect 100 -2673 101 -2671
rect 103 -2673 104 -2671
rect 100 -2679 101 -2677
rect 103 -2679 104 -2677
rect 107 -2673 108 -2671
rect 107 -2679 108 -2677
rect 114 -2673 115 -2671
rect 114 -2679 115 -2677
rect 121 -2673 122 -2671
rect 121 -2679 122 -2677
rect 128 -2673 129 -2671
rect 131 -2673 132 -2671
rect 128 -2679 129 -2677
rect 131 -2679 132 -2677
rect 135 -2673 136 -2671
rect 135 -2679 136 -2677
rect 142 -2673 143 -2671
rect 142 -2679 143 -2677
rect 149 -2673 150 -2671
rect 149 -2679 150 -2677
rect 156 -2673 157 -2671
rect 156 -2679 157 -2677
rect 163 -2673 164 -2671
rect 163 -2679 164 -2677
rect 170 -2673 171 -2671
rect 170 -2679 171 -2677
rect 177 -2673 178 -2671
rect 177 -2679 178 -2677
rect 184 -2673 185 -2671
rect 184 -2679 185 -2677
rect 191 -2673 192 -2671
rect 191 -2679 192 -2677
rect 198 -2673 199 -2671
rect 201 -2673 202 -2671
rect 198 -2679 199 -2677
rect 205 -2673 206 -2671
rect 205 -2679 206 -2677
rect 212 -2673 213 -2671
rect 212 -2679 213 -2677
rect 219 -2673 220 -2671
rect 219 -2679 220 -2677
rect 226 -2673 227 -2671
rect 226 -2679 227 -2677
rect 233 -2673 234 -2671
rect 233 -2679 234 -2677
rect 240 -2673 241 -2671
rect 240 -2679 241 -2677
rect 243 -2679 244 -2677
rect 247 -2673 248 -2671
rect 247 -2679 248 -2677
rect 254 -2673 255 -2671
rect 254 -2679 255 -2677
rect 261 -2673 262 -2671
rect 261 -2679 262 -2677
rect 268 -2673 269 -2671
rect 268 -2679 269 -2677
rect 275 -2673 276 -2671
rect 275 -2679 276 -2677
rect 282 -2673 283 -2671
rect 282 -2679 283 -2677
rect 289 -2673 290 -2671
rect 289 -2679 290 -2677
rect 296 -2673 297 -2671
rect 296 -2679 297 -2677
rect 303 -2673 304 -2671
rect 303 -2679 304 -2677
rect 310 -2673 311 -2671
rect 310 -2679 311 -2677
rect 317 -2673 318 -2671
rect 317 -2679 318 -2677
rect 324 -2673 325 -2671
rect 324 -2679 325 -2677
rect 331 -2673 332 -2671
rect 331 -2679 332 -2677
rect 338 -2673 339 -2671
rect 338 -2679 339 -2677
rect 345 -2673 346 -2671
rect 345 -2679 346 -2677
rect 352 -2673 353 -2671
rect 352 -2679 353 -2677
rect 359 -2673 360 -2671
rect 359 -2679 360 -2677
rect 366 -2673 367 -2671
rect 366 -2679 367 -2677
rect 373 -2673 374 -2671
rect 373 -2679 374 -2677
rect 380 -2673 381 -2671
rect 380 -2679 381 -2677
rect 387 -2673 388 -2671
rect 387 -2679 388 -2677
rect 394 -2673 395 -2671
rect 394 -2679 395 -2677
rect 401 -2673 402 -2671
rect 401 -2679 402 -2677
rect 408 -2673 409 -2671
rect 411 -2673 412 -2671
rect 408 -2679 409 -2677
rect 411 -2679 412 -2677
rect 415 -2673 416 -2671
rect 415 -2679 416 -2677
rect 422 -2673 423 -2671
rect 422 -2679 423 -2677
rect 429 -2673 430 -2671
rect 429 -2679 430 -2677
rect 436 -2673 437 -2671
rect 436 -2679 437 -2677
rect 443 -2673 444 -2671
rect 443 -2679 444 -2677
rect 450 -2673 451 -2671
rect 450 -2679 451 -2677
rect 457 -2673 458 -2671
rect 457 -2679 458 -2677
rect 464 -2673 465 -2671
rect 464 -2679 465 -2677
rect 471 -2673 472 -2671
rect 471 -2679 472 -2677
rect 478 -2673 479 -2671
rect 478 -2679 479 -2677
rect 485 -2673 486 -2671
rect 485 -2679 486 -2677
rect 492 -2673 493 -2671
rect 492 -2679 493 -2677
rect 499 -2673 500 -2671
rect 499 -2679 500 -2677
rect 506 -2673 507 -2671
rect 506 -2679 507 -2677
rect 513 -2673 514 -2671
rect 513 -2679 514 -2677
rect 520 -2673 521 -2671
rect 520 -2679 521 -2677
rect 527 -2673 528 -2671
rect 527 -2679 528 -2677
rect 534 -2673 535 -2671
rect 534 -2679 535 -2677
rect 541 -2673 542 -2671
rect 541 -2679 542 -2677
rect 548 -2673 549 -2671
rect 548 -2679 549 -2677
rect 555 -2673 556 -2671
rect 558 -2673 559 -2671
rect 555 -2679 556 -2677
rect 558 -2679 559 -2677
rect 562 -2673 563 -2671
rect 562 -2679 563 -2677
rect 569 -2673 570 -2671
rect 569 -2679 570 -2677
rect 576 -2673 577 -2671
rect 576 -2679 577 -2677
rect 583 -2673 584 -2671
rect 583 -2679 584 -2677
rect 590 -2673 591 -2671
rect 590 -2679 591 -2677
rect 597 -2673 598 -2671
rect 597 -2679 598 -2677
rect 604 -2673 605 -2671
rect 604 -2679 605 -2677
rect 611 -2673 612 -2671
rect 611 -2679 612 -2677
rect 618 -2673 619 -2671
rect 618 -2679 619 -2677
rect 625 -2673 626 -2671
rect 625 -2679 626 -2677
rect 632 -2673 633 -2671
rect 632 -2679 633 -2677
rect 639 -2673 640 -2671
rect 639 -2679 640 -2677
rect 646 -2673 647 -2671
rect 646 -2679 647 -2677
rect 653 -2673 654 -2671
rect 653 -2679 654 -2677
rect 660 -2673 661 -2671
rect 660 -2679 661 -2677
rect 667 -2673 668 -2671
rect 667 -2679 668 -2677
rect 674 -2673 675 -2671
rect 674 -2679 675 -2677
rect 681 -2673 682 -2671
rect 681 -2679 682 -2677
rect 688 -2673 689 -2671
rect 688 -2679 689 -2677
rect 695 -2673 696 -2671
rect 695 -2679 696 -2677
rect 702 -2673 703 -2671
rect 702 -2679 703 -2677
rect 709 -2673 710 -2671
rect 709 -2679 710 -2677
rect 716 -2673 717 -2671
rect 716 -2679 717 -2677
rect 726 -2673 727 -2671
rect 726 -2679 727 -2677
rect 730 -2673 731 -2671
rect 730 -2679 731 -2677
rect 737 -2673 738 -2671
rect 737 -2679 738 -2677
rect 744 -2673 745 -2671
rect 744 -2679 745 -2677
rect 751 -2673 752 -2671
rect 751 -2679 752 -2677
rect 758 -2673 759 -2671
rect 758 -2679 759 -2677
rect 765 -2673 766 -2671
rect 765 -2679 766 -2677
rect 772 -2673 773 -2671
rect 772 -2679 773 -2677
rect 779 -2673 780 -2671
rect 779 -2679 780 -2677
rect 786 -2673 787 -2671
rect 789 -2673 790 -2671
rect 786 -2679 787 -2677
rect 789 -2679 790 -2677
rect 793 -2673 794 -2671
rect 793 -2679 794 -2677
rect 800 -2673 801 -2671
rect 800 -2679 801 -2677
rect 810 -2673 811 -2671
rect 807 -2679 808 -2677
rect 810 -2679 811 -2677
rect 814 -2673 815 -2671
rect 817 -2673 818 -2671
rect 814 -2679 815 -2677
rect 817 -2679 818 -2677
rect 821 -2673 822 -2671
rect 824 -2673 825 -2671
rect 821 -2679 822 -2677
rect 824 -2679 825 -2677
rect 828 -2673 829 -2671
rect 828 -2679 829 -2677
rect 835 -2673 836 -2671
rect 835 -2679 836 -2677
rect 842 -2673 843 -2671
rect 842 -2679 843 -2677
rect 849 -2673 850 -2671
rect 849 -2679 850 -2677
rect 856 -2673 857 -2671
rect 856 -2679 857 -2677
rect 863 -2673 864 -2671
rect 863 -2679 864 -2677
rect 870 -2673 871 -2671
rect 870 -2679 871 -2677
rect 877 -2673 878 -2671
rect 877 -2679 878 -2677
rect 884 -2673 885 -2671
rect 884 -2679 885 -2677
rect 891 -2673 892 -2671
rect 894 -2673 895 -2671
rect 894 -2679 895 -2677
rect 898 -2673 899 -2671
rect 898 -2679 899 -2677
rect 905 -2673 906 -2671
rect 905 -2679 906 -2677
rect 912 -2673 913 -2671
rect 912 -2679 913 -2677
rect 919 -2679 920 -2677
rect 922 -2679 923 -2677
rect 926 -2673 927 -2671
rect 926 -2679 927 -2677
rect 933 -2673 934 -2671
rect 933 -2679 934 -2677
rect 940 -2673 941 -2671
rect 940 -2679 941 -2677
rect 947 -2673 948 -2671
rect 950 -2673 951 -2671
rect 947 -2679 948 -2677
rect 950 -2679 951 -2677
rect 954 -2673 955 -2671
rect 954 -2679 955 -2677
rect 957 -2679 958 -2677
rect 961 -2673 962 -2671
rect 961 -2679 962 -2677
rect 968 -2673 969 -2671
rect 968 -2679 969 -2677
rect 975 -2673 976 -2671
rect 975 -2679 976 -2677
rect 982 -2673 983 -2671
rect 982 -2679 983 -2677
rect 989 -2673 990 -2671
rect 989 -2679 990 -2677
rect 996 -2673 997 -2671
rect 996 -2679 997 -2677
rect 1003 -2673 1004 -2671
rect 1006 -2673 1007 -2671
rect 1003 -2679 1004 -2677
rect 1010 -2673 1011 -2671
rect 1013 -2673 1014 -2671
rect 1010 -2679 1011 -2677
rect 1013 -2679 1014 -2677
rect 1017 -2673 1018 -2671
rect 1017 -2679 1018 -2677
rect 1024 -2673 1025 -2671
rect 1024 -2679 1025 -2677
rect 1031 -2673 1032 -2671
rect 1031 -2679 1032 -2677
rect 1038 -2673 1039 -2671
rect 1038 -2679 1039 -2677
rect 1041 -2679 1042 -2677
rect 1045 -2673 1046 -2671
rect 1045 -2679 1046 -2677
rect 1052 -2673 1053 -2671
rect 1052 -2679 1053 -2677
rect 1059 -2673 1060 -2671
rect 1059 -2679 1060 -2677
rect 1066 -2673 1067 -2671
rect 1066 -2679 1067 -2677
rect 1073 -2673 1074 -2671
rect 1073 -2679 1074 -2677
rect 1080 -2673 1081 -2671
rect 1080 -2679 1081 -2677
rect 1087 -2673 1088 -2671
rect 1087 -2679 1088 -2677
rect 1094 -2673 1095 -2671
rect 1094 -2679 1095 -2677
rect 1101 -2673 1102 -2671
rect 1101 -2679 1102 -2677
rect 1108 -2673 1109 -2671
rect 1108 -2679 1109 -2677
rect 1115 -2673 1116 -2671
rect 1115 -2679 1116 -2677
rect 1122 -2673 1123 -2671
rect 1125 -2673 1126 -2671
rect 1122 -2679 1123 -2677
rect 1125 -2679 1126 -2677
rect 1129 -2673 1130 -2671
rect 1129 -2679 1130 -2677
rect 1136 -2673 1137 -2671
rect 1139 -2679 1140 -2677
rect 1143 -2673 1144 -2671
rect 1143 -2679 1144 -2677
rect 1150 -2673 1151 -2671
rect 1150 -2679 1151 -2677
rect 1157 -2673 1158 -2671
rect 1157 -2679 1158 -2677
rect 1164 -2673 1165 -2671
rect 1164 -2679 1165 -2677
rect 1171 -2673 1172 -2671
rect 1171 -2679 1172 -2677
rect 1178 -2673 1179 -2671
rect 1178 -2679 1179 -2677
rect 1185 -2673 1186 -2671
rect 1188 -2673 1189 -2671
rect 1185 -2679 1186 -2677
rect 1192 -2673 1193 -2671
rect 1195 -2673 1196 -2671
rect 1192 -2679 1193 -2677
rect 1195 -2679 1196 -2677
rect 1199 -2673 1200 -2671
rect 1199 -2679 1200 -2677
rect 1206 -2673 1207 -2671
rect 1206 -2679 1207 -2677
rect 1213 -2673 1214 -2671
rect 1213 -2679 1214 -2677
rect 1220 -2673 1221 -2671
rect 1220 -2679 1221 -2677
rect 1227 -2673 1228 -2671
rect 1227 -2679 1228 -2677
rect 1234 -2673 1235 -2671
rect 1237 -2673 1238 -2671
rect 1234 -2679 1235 -2677
rect 1241 -2673 1242 -2671
rect 1241 -2679 1242 -2677
rect 1244 -2679 1245 -2677
rect 1248 -2673 1249 -2671
rect 1248 -2679 1249 -2677
rect 1255 -2673 1256 -2671
rect 1255 -2679 1256 -2677
rect 1262 -2673 1263 -2671
rect 1262 -2679 1263 -2677
rect 1269 -2673 1270 -2671
rect 1269 -2679 1270 -2677
rect 1276 -2673 1277 -2671
rect 1276 -2679 1277 -2677
rect 1283 -2673 1284 -2671
rect 1283 -2679 1284 -2677
rect 1290 -2673 1291 -2671
rect 1290 -2679 1291 -2677
rect 1297 -2673 1298 -2671
rect 1297 -2679 1298 -2677
rect 1304 -2673 1305 -2671
rect 1304 -2679 1305 -2677
rect 1311 -2673 1312 -2671
rect 1314 -2673 1315 -2671
rect 1311 -2679 1312 -2677
rect 1314 -2679 1315 -2677
rect 1318 -2673 1319 -2671
rect 1318 -2679 1319 -2677
rect 1325 -2679 1326 -2677
rect 1328 -2679 1329 -2677
rect 1332 -2673 1333 -2671
rect 1332 -2679 1333 -2677
rect 1339 -2673 1340 -2671
rect 1339 -2679 1340 -2677
rect 1346 -2673 1347 -2671
rect 1346 -2679 1347 -2677
rect 1353 -2673 1354 -2671
rect 1353 -2679 1354 -2677
rect 1360 -2673 1361 -2671
rect 1360 -2679 1361 -2677
rect 1367 -2673 1368 -2671
rect 1367 -2679 1368 -2677
rect 1374 -2673 1375 -2671
rect 1374 -2679 1375 -2677
rect 1381 -2673 1382 -2671
rect 1381 -2679 1382 -2677
rect 1388 -2673 1389 -2671
rect 1388 -2679 1389 -2677
rect 1395 -2673 1396 -2671
rect 1398 -2673 1399 -2671
rect 1395 -2679 1396 -2677
rect 1398 -2679 1399 -2677
rect 1402 -2673 1403 -2671
rect 1402 -2679 1403 -2677
rect 1409 -2673 1410 -2671
rect 1412 -2673 1413 -2671
rect 1409 -2679 1410 -2677
rect 1416 -2673 1417 -2671
rect 1416 -2679 1417 -2677
rect 1423 -2673 1424 -2671
rect 1423 -2679 1424 -2677
rect 1430 -2673 1431 -2671
rect 1430 -2679 1431 -2677
rect 1433 -2679 1434 -2677
rect 1437 -2673 1438 -2671
rect 1440 -2673 1441 -2671
rect 1437 -2679 1438 -2677
rect 1440 -2679 1441 -2677
rect 1444 -2673 1445 -2671
rect 1447 -2673 1448 -2671
rect 1444 -2679 1445 -2677
rect 1451 -2673 1452 -2671
rect 1451 -2679 1452 -2677
rect 1458 -2673 1459 -2671
rect 1458 -2679 1459 -2677
rect 1465 -2673 1466 -2671
rect 1465 -2679 1466 -2677
rect 1472 -2673 1473 -2671
rect 1472 -2679 1473 -2677
rect 1479 -2673 1480 -2671
rect 1479 -2679 1480 -2677
rect 1486 -2673 1487 -2671
rect 1486 -2679 1487 -2677
rect 1493 -2673 1494 -2671
rect 1493 -2679 1494 -2677
rect 1500 -2673 1501 -2671
rect 1500 -2679 1501 -2677
rect 1507 -2673 1508 -2671
rect 1510 -2673 1511 -2671
rect 1507 -2679 1508 -2677
rect 1510 -2679 1511 -2677
rect 1514 -2673 1515 -2671
rect 1514 -2679 1515 -2677
rect 1521 -2673 1522 -2671
rect 1521 -2679 1522 -2677
rect 1528 -2673 1529 -2671
rect 1528 -2679 1529 -2677
rect 1535 -2673 1536 -2671
rect 1535 -2679 1536 -2677
rect 1542 -2673 1543 -2671
rect 1542 -2679 1543 -2677
rect 1549 -2673 1550 -2671
rect 1549 -2679 1550 -2677
rect 1556 -2673 1557 -2671
rect 1556 -2679 1557 -2677
rect 1563 -2673 1564 -2671
rect 1563 -2679 1564 -2677
rect 1570 -2673 1571 -2671
rect 1570 -2679 1571 -2677
rect 1577 -2673 1578 -2671
rect 1580 -2673 1581 -2671
rect 1577 -2679 1578 -2677
rect 1580 -2679 1581 -2677
rect 1584 -2673 1585 -2671
rect 1584 -2679 1585 -2677
rect 1591 -2673 1592 -2671
rect 1591 -2679 1592 -2677
rect 1598 -2673 1599 -2671
rect 1598 -2679 1599 -2677
rect 1605 -2673 1606 -2671
rect 1605 -2679 1606 -2677
rect 1612 -2673 1613 -2671
rect 1612 -2679 1613 -2677
rect 1619 -2673 1620 -2671
rect 1619 -2679 1620 -2677
rect 1626 -2673 1627 -2671
rect 1626 -2679 1627 -2677
rect 1633 -2673 1634 -2671
rect 1633 -2679 1634 -2677
rect 1640 -2673 1641 -2671
rect 1640 -2679 1641 -2677
rect 1647 -2673 1648 -2671
rect 1647 -2679 1648 -2677
rect 1654 -2673 1655 -2671
rect 1654 -2679 1655 -2677
rect 1661 -2673 1662 -2671
rect 1661 -2679 1662 -2677
rect 1668 -2673 1669 -2671
rect 1668 -2679 1669 -2677
rect 1675 -2673 1676 -2671
rect 1675 -2679 1676 -2677
rect 1682 -2673 1683 -2671
rect 1682 -2679 1683 -2677
rect 1689 -2673 1690 -2671
rect 1689 -2679 1690 -2677
rect 1696 -2673 1697 -2671
rect 1696 -2679 1697 -2677
rect 1703 -2673 1704 -2671
rect 1703 -2679 1704 -2677
rect 1710 -2673 1711 -2671
rect 1710 -2679 1711 -2677
rect 1717 -2673 1718 -2671
rect 1717 -2679 1718 -2677
rect 1724 -2673 1725 -2671
rect 1724 -2679 1725 -2677
rect 1731 -2673 1732 -2671
rect 1731 -2679 1732 -2677
rect 1738 -2673 1739 -2671
rect 1738 -2679 1739 -2677
rect 1745 -2673 1746 -2671
rect 1745 -2679 1746 -2677
rect 1752 -2673 1753 -2671
rect 1755 -2673 1756 -2671
rect 1752 -2679 1753 -2677
rect 1755 -2679 1756 -2677
rect 1759 -2673 1760 -2671
rect 1759 -2679 1760 -2677
rect 1766 -2673 1767 -2671
rect 1766 -2679 1767 -2677
rect 1773 -2673 1774 -2671
rect 1773 -2679 1774 -2677
rect 1780 -2673 1781 -2671
rect 1780 -2679 1781 -2677
rect 1787 -2673 1788 -2671
rect 1787 -2679 1788 -2677
rect 1794 -2673 1795 -2671
rect 1794 -2679 1795 -2677
rect 1801 -2673 1802 -2671
rect 1801 -2679 1802 -2677
rect 1808 -2673 1809 -2671
rect 1808 -2679 1809 -2677
rect 1815 -2673 1816 -2671
rect 1815 -2679 1816 -2677
rect 1822 -2673 1823 -2671
rect 1822 -2679 1823 -2677
rect 1829 -2673 1830 -2671
rect 1829 -2679 1830 -2677
rect 1836 -2673 1837 -2671
rect 1836 -2679 1837 -2677
rect 1843 -2673 1844 -2671
rect 1843 -2679 1844 -2677
rect 1850 -2673 1851 -2671
rect 1850 -2679 1851 -2677
rect 1857 -2673 1858 -2671
rect 1857 -2679 1858 -2677
rect 1864 -2673 1865 -2671
rect 1864 -2679 1865 -2677
rect 1871 -2673 1872 -2671
rect 1871 -2679 1872 -2677
rect 1878 -2673 1879 -2671
rect 1878 -2679 1879 -2677
rect 1885 -2673 1886 -2671
rect 1885 -2679 1886 -2677
rect 1892 -2673 1893 -2671
rect 1892 -2679 1893 -2677
rect 1899 -2673 1900 -2671
rect 1899 -2679 1900 -2677
rect 1906 -2673 1907 -2671
rect 1906 -2679 1907 -2677
rect 1913 -2673 1914 -2671
rect 1913 -2679 1914 -2677
rect 1920 -2673 1921 -2671
rect 1920 -2679 1921 -2677
rect 1927 -2673 1928 -2671
rect 1927 -2679 1928 -2677
rect 1934 -2673 1935 -2671
rect 1934 -2679 1935 -2677
rect 1941 -2673 1942 -2671
rect 1941 -2679 1942 -2677
rect 1948 -2673 1949 -2671
rect 1948 -2679 1949 -2677
rect 1955 -2673 1956 -2671
rect 1955 -2679 1956 -2677
rect 1962 -2673 1963 -2671
rect 1962 -2679 1963 -2677
rect 1969 -2673 1970 -2671
rect 1969 -2679 1970 -2677
rect 1976 -2673 1977 -2671
rect 1976 -2679 1977 -2677
rect 1983 -2673 1984 -2671
rect 1983 -2679 1984 -2677
rect 1990 -2673 1991 -2671
rect 1990 -2679 1991 -2677
rect 1997 -2673 1998 -2671
rect 1997 -2679 1998 -2677
rect 2004 -2673 2005 -2671
rect 2004 -2679 2005 -2677
rect 2011 -2673 2012 -2671
rect 2011 -2679 2012 -2677
rect 2018 -2673 2019 -2671
rect 2018 -2679 2019 -2677
rect 2025 -2673 2026 -2671
rect 2025 -2679 2026 -2677
rect 2032 -2673 2033 -2671
rect 2032 -2679 2033 -2677
rect 2039 -2673 2040 -2671
rect 2039 -2679 2040 -2677
rect 2046 -2673 2047 -2671
rect 2046 -2679 2047 -2677
rect 2053 -2673 2054 -2671
rect 2053 -2679 2054 -2677
rect 2060 -2673 2061 -2671
rect 2060 -2679 2061 -2677
rect 2067 -2673 2068 -2671
rect 2067 -2679 2068 -2677
rect 2074 -2673 2075 -2671
rect 2074 -2679 2075 -2677
rect 2081 -2673 2082 -2671
rect 2081 -2679 2082 -2677
rect 2088 -2673 2089 -2671
rect 2088 -2679 2089 -2677
rect 2095 -2673 2096 -2671
rect 2095 -2679 2096 -2677
rect 2102 -2673 2103 -2671
rect 2102 -2679 2103 -2677
rect 2109 -2673 2110 -2671
rect 2109 -2679 2110 -2677
rect 2116 -2673 2117 -2671
rect 2116 -2679 2117 -2677
rect 2123 -2673 2124 -2671
rect 2123 -2679 2124 -2677
rect 2130 -2673 2131 -2671
rect 2130 -2679 2131 -2677
rect 2137 -2673 2138 -2671
rect 2137 -2679 2138 -2677
rect 2144 -2673 2145 -2671
rect 2144 -2679 2145 -2677
rect 2151 -2673 2152 -2671
rect 2151 -2679 2152 -2677
rect 2158 -2673 2159 -2671
rect 2158 -2679 2159 -2677
rect 2165 -2673 2166 -2671
rect 2165 -2679 2166 -2677
rect 2172 -2673 2173 -2671
rect 2172 -2679 2173 -2677
rect 2179 -2673 2180 -2671
rect 2179 -2679 2180 -2677
rect 2186 -2673 2187 -2671
rect 2186 -2679 2187 -2677
rect 2193 -2673 2194 -2671
rect 2193 -2679 2194 -2677
rect 2200 -2673 2201 -2671
rect 2200 -2679 2201 -2677
rect 2207 -2673 2208 -2671
rect 2207 -2679 2208 -2677
rect 2214 -2673 2215 -2671
rect 2214 -2679 2215 -2677
rect 2221 -2673 2222 -2671
rect 2221 -2679 2222 -2677
rect 2228 -2673 2229 -2671
rect 2228 -2679 2229 -2677
rect 2235 -2673 2236 -2671
rect 2235 -2679 2236 -2677
rect 2242 -2673 2243 -2671
rect 2242 -2679 2243 -2677
rect 2263 -2673 2264 -2671
rect 2263 -2679 2264 -2677
rect 2270 -2673 2271 -2671
rect 2270 -2679 2271 -2677
rect 2 -2836 3 -2834
rect 2 -2842 3 -2840
rect 9 -2836 10 -2834
rect 9 -2842 10 -2840
rect 16 -2836 17 -2834
rect 16 -2842 17 -2840
rect 23 -2836 24 -2834
rect 23 -2842 24 -2840
rect 30 -2836 31 -2834
rect 30 -2842 31 -2840
rect 37 -2836 38 -2834
rect 37 -2842 38 -2840
rect 44 -2836 45 -2834
rect 44 -2842 45 -2840
rect 51 -2836 52 -2834
rect 54 -2836 55 -2834
rect 51 -2842 52 -2840
rect 58 -2836 59 -2834
rect 58 -2842 59 -2840
rect 65 -2836 66 -2834
rect 65 -2842 66 -2840
rect 72 -2836 73 -2834
rect 72 -2842 73 -2840
rect 79 -2836 80 -2834
rect 82 -2836 83 -2834
rect 79 -2842 80 -2840
rect 82 -2842 83 -2840
rect 86 -2836 87 -2834
rect 86 -2842 87 -2840
rect 93 -2836 94 -2834
rect 93 -2842 94 -2840
rect 100 -2836 101 -2834
rect 100 -2842 101 -2840
rect 110 -2836 111 -2834
rect 107 -2842 108 -2840
rect 114 -2836 115 -2834
rect 114 -2842 115 -2840
rect 121 -2836 122 -2834
rect 121 -2842 122 -2840
rect 128 -2836 129 -2834
rect 128 -2842 129 -2840
rect 135 -2836 136 -2834
rect 135 -2842 136 -2840
rect 142 -2836 143 -2834
rect 142 -2842 143 -2840
rect 149 -2836 150 -2834
rect 149 -2842 150 -2840
rect 156 -2836 157 -2834
rect 156 -2842 157 -2840
rect 163 -2836 164 -2834
rect 163 -2842 164 -2840
rect 170 -2836 171 -2834
rect 170 -2842 171 -2840
rect 177 -2836 178 -2834
rect 177 -2842 178 -2840
rect 184 -2836 185 -2834
rect 184 -2842 185 -2840
rect 191 -2836 192 -2834
rect 191 -2842 192 -2840
rect 198 -2836 199 -2834
rect 198 -2842 199 -2840
rect 205 -2836 206 -2834
rect 205 -2842 206 -2840
rect 212 -2836 213 -2834
rect 212 -2842 213 -2840
rect 219 -2836 220 -2834
rect 222 -2836 223 -2834
rect 219 -2842 220 -2840
rect 222 -2842 223 -2840
rect 226 -2836 227 -2834
rect 226 -2842 227 -2840
rect 236 -2836 237 -2834
rect 233 -2842 234 -2840
rect 236 -2842 237 -2840
rect 240 -2836 241 -2834
rect 240 -2842 241 -2840
rect 247 -2836 248 -2834
rect 250 -2836 251 -2834
rect 247 -2842 248 -2840
rect 250 -2842 251 -2840
rect 254 -2836 255 -2834
rect 254 -2842 255 -2840
rect 261 -2836 262 -2834
rect 261 -2842 262 -2840
rect 268 -2836 269 -2834
rect 268 -2842 269 -2840
rect 275 -2836 276 -2834
rect 275 -2842 276 -2840
rect 282 -2836 283 -2834
rect 282 -2842 283 -2840
rect 289 -2836 290 -2834
rect 289 -2842 290 -2840
rect 296 -2836 297 -2834
rect 296 -2842 297 -2840
rect 303 -2836 304 -2834
rect 303 -2842 304 -2840
rect 310 -2836 311 -2834
rect 310 -2842 311 -2840
rect 317 -2836 318 -2834
rect 317 -2842 318 -2840
rect 324 -2836 325 -2834
rect 324 -2842 325 -2840
rect 331 -2836 332 -2834
rect 331 -2842 332 -2840
rect 338 -2836 339 -2834
rect 338 -2842 339 -2840
rect 345 -2836 346 -2834
rect 345 -2842 346 -2840
rect 352 -2836 353 -2834
rect 352 -2842 353 -2840
rect 359 -2836 360 -2834
rect 359 -2842 360 -2840
rect 366 -2836 367 -2834
rect 366 -2842 367 -2840
rect 373 -2836 374 -2834
rect 373 -2842 374 -2840
rect 380 -2836 381 -2834
rect 380 -2842 381 -2840
rect 387 -2836 388 -2834
rect 387 -2842 388 -2840
rect 394 -2836 395 -2834
rect 394 -2842 395 -2840
rect 401 -2836 402 -2834
rect 401 -2842 402 -2840
rect 408 -2836 409 -2834
rect 408 -2842 409 -2840
rect 415 -2836 416 -2834
rect 415 -2842 416 -2840
rect 422 -2836 423 -2834
rect 422 -2842 423 -2840
rect 432 -2836 433 -2834
rect 429 -2842 430 -2840
rect 436 -2836 437 -2834
rect 436 -2842 437 -2840
rect 443 -2836 444 -2834
rect 443 -2842 444 -2840
rect 450 -2836 451 -2834
rect 450 -2842 451 -2840
rect 457 -2836 458 -2834
rect 460 -2836 461 -2834
rect 460 -2842 461 -2840
rect 464 -2836 465 -2834
rect 464 -2842 465 -2840
rect 471 -2836 472 -2834
rect 471 -2842 472 -2840
rect 478 -2836 479 -2834
rect 478 -2842 479 -2840
rect 485 -2836 486 -2834
rect 485 -2842 486 -2840
rect 492 -2836 493 -2834
rect 492 -2842 493 -2840
rect 499 -2836 500 -2834
rect 499 -2842 500 -2840
rect 506 -2836 507 -2834
rect 506 -2842 507 -2840
rect 513 -2836 514 -2834
rect 513 -2842 514 -2840
rect 520 -2836 521 -2834
rect 520 -2842 521 -2840
rect 527 -2836 528 -2834
rect 527 -2842 528 -2840
rect 534 -2836 535 -2834
rect 534 -2842 535 -2840
rect 541 -2836 542 -2834
rect 544 -2836 545 -2834
rect 544 -2842 545 -2840
rect 548 -2836 549 -2834
rect 548 -2842 549 -2840
rect 555 -2836 556 -2834
rect 555 -2842 556 -2840
rect 562 -2836 563 -2834
rect 562 -2842 563 -2840
rect 569 -2836 570 -2834
rect 569 -2842 570 -2840
rect 576 -2836 577 -2834
rect 576 -2842 577 -2840
rect 583 -2836 584 -2834
rect 583 -2842 584 -2840
rect 590 -2836 591 -2834
rect 590 -2842 591 -2840
rect 597 -2836 598 -2834
rect 597 -2842 598 -2840
rect 604 -2836 605 -2834
rect 604 -2842 605 -2840
rect 611 -2836 612 -2834
rect 611 -2842 612 -2840
rect 618 -2836 619 -2834
rect 621 -2836 622 -2834
rect 618 -2842 619 -2840
rect 621 -2842 622 -2840
rect 625 -2836 626 -2834
rect 625 -2842 626 -2840
rect 632 -2836 633 -2834
rect 632 -2842 633 -2840
rect 639 -2836 640 -2834
rect 639 -2842 640 -2840
rect 646 -2836 647 -2834
rect 646 -2842 647 -2840
rect 653 -2836 654 -2834
rect 653 -2842 654 -2840
rect 660 -2836 661 -2834
rect 663 -2836 664 -2834
rect 660 -2842 661 -2840
rect 663 -2842 664 -2840
rect 667 -2836 668 -2834
rect 667 -2842 668 -2840
rect 674 -2836 675 -2834
rect 674 -2842 675 -2840
rect 681 -2836 682 -2834
rect 681 -2842 682 -2840
rect 688 -2836 689 -2834
rect 688 -2842 689 -2840
rect 695 -2836 696 -2834
rect 695 -2842 696 -2840
rect 702 -2836 703 -2834
rect 705 -2836 706 -2834
rect 702 -2842 703 -2840
rect 705 -2842 706 -2840
rect 709 -2836 710 -2834
rect 709 -2842 710 -2840
rect 716 -2836 717 -2834
rect 716 -2842 717 -2840
rect 723 -2836 724 -2834
rect 723 -2842 724 -2840
rect 730 -2836 731 -2834
rect 733 -2836 734 -2834
rect 730 -2842 731 -2840
rect 733 -2842 734 -2840
rect 737 -2836 738 -2834
rect 737 -2842 738 -2840
rect 744 -2836 745 -2834
rect 744 -2842 745 -2840
rect 747 -2842 748 -2840
rect 751 -2836 752 -2834
rect 751 -2842 752 -2840
rect 758 -2836 759 -2834
rect 758 -2842 759 -2840
rect 765 -2836 766 -2834
rect 765 -2842 766 -2840
rect 772 -2836 773 -2834
rect 772 -2842 773 -2840
rect 779 -2836 780 -2834
rect 779 -2842 780 -2840
rect 786 -2836 787 -2834
rect 789 -2836 790 -2834
rect 789 -2842 790 -2840
rect 793 -2836 794 -2834
rect 793 -2842 794 -2840
rect 800 -2836 801 -2834
rect 800 -2842 801 -2840
rect 807 -2836 808 -2834
rect 807 -2842 808 -2840
rect 814 -2836 815 -2834
rect 814 -2842 815 -2840
rect 821 -2836 822 -2834
rect 821 -2842 822 -2840
rect 828 -2836 829 -2834
rect 828 -2842 829 -2840
rect 835 -2836 836 -2834
rect 838 -2836 839 -2834
rect 842 -2836 843 -2834
rect 842 -2842 843 -2840
rect 849 -2836 850 -2834
rect 849 -2842 850 -2840
rect 856 -2836 857 -2834
rect 856 -2842 857 -2840
rect 863 -2836 864 -2834
rect 866 -2836 867 -2834
rect 863 -2842 864 -2840
rect 866 -2842 867 -2840
rect 870 -2836 871 -2834
rect 870 -2842 871 -2840
rect 877 -2836 878 -2834
rect 877 -2842 878 -2840
rect 884 -2836 885 -2834
rect 884 -2842 885 -2840
rect 891 -2836 892 -2834
rect 891 -2842 892 -2840
rect 898 -2836 899 -2834
rect 898 -2842 899 -2840
rect 905 -2836 906 -2834
rect 905 -2842 906 -2840
rect 912 -2836 913 -2834
rect 915 -2836 916 -2834
rect 912 -2842 913 -2840
rect 919 -2836 920 -2834
rect 919 -2842 920 -2840
rect 926 -2836 927 -2834
rect 926 -2842 927 -2840
rect 933 -2836 934 -2834
rect 933 -2842 934 -2840
rect 940 -2836 941 -2834
rect 943 -2836 944 -2834
rect 940 -2842 941 -2840
rect 943 -2842 944 -2840
rect 947 -2836 948 -2834
rect 947 -2842 948 -2840
rect 954 -2836 955 -2834
rect 954 -2842 955 -2840
rect 961 -2836 962 -2834
rect 964 -2836 965 -2834
rect 961 -2842 962 -2840
rect 968 -2836 969 -2834
rect 968 -2842 969 -2840
rect 975 -2836 976 -2834
rect 978 -2836 979 -2834
rect 978 -2842 979 -2840
rect 982 -2836 983 -2834
rect 982 -2842 983 -2840
rect 989 -2836 990 -2834
rect 989 -2842 990 -2840
rect 996 -2836 997 -2834
rect 996 -2842 997 -2840
rect 1003 -2836 1004 -2834
rect 1003 -2842 1004 -2840
rect 1010 -2836 1011 -2834
rect 1010 -2842 1011 -2840
rect 1017 -2836 1018 -2834
rect 1017 -2842 1018 -2840
rect 1024 -2836 1025 -2834
rect 1024 -2842 1025 -2840
rect 1031 -2836 1032 -2834
rect 1031 -2842 1032 -2840
rect 1038 -2836 1039 -2834
rect 1038 -2842 1039 -2840
rect 1045 -2836 1046 -2834
rect 1045 -2842 1046 -2840
rect 1052 -2836 1053 -2834
rect 1055 -2836 1056 -2834
rect 1052 -2842 1053 -2840
rect 1055 -2842 1056 -2840
rect 1059 -2836 1060 -2834
rect 1062 -2836 1063 -2834
rect 1059 -2842 1060 -2840
rect 1066 -2836 1067 -2834
rect 1066 -2842 1067 -2840
rect 1073 -2836 1074 -2834
rect 1073 -2842 1074 -2840
rect 1080 -2836 1081 -2834
rect 1080 -2842 1081 -2840
rect 1087 -2836 1088 -2834
rect 1087 -2842 1088 -2840
rect 1094 -2836 1095 -2834
rect 1097 -2836 1098 -2834
rect 1094 -2842 1095 -2840
rect 1097 -2842 1098 -2840
rect 1101 -2836 1102 -2834
rect 1101 -2842 1102 -2840
rect 1108 -2836 1109 -2834
rect 1108 -2842 1109 -2840
rect 1115 -2836 1116 -2834
rect 1115 -2842 1116 -2840
rect 1122 -2836 1123 -2834
rect 1122 -2842 1123 -2840
rect 1129 -2836 1130 -2834
rect 1129 -2842 1130 -2840
rect 1136 -2836 1137 -2834
rect 1136 -2842 1137 -2840
rect 1143 -2836 1144 -2834
rect 1143 -2842 1144 -2840
rect 1150 -2836 1151 -2834
rect 1150 -2842 1151 -2840
rect 1157 -2836 1158 -2834
rect 1157 -2842 1158 -2840
rect 1164 -2836 1165 -2834
rect 1164 -2842 1165 -2840
rect 1171 -2836 1172 -2834
rect 1171 -2842 1172 -2840
rect 1178 -2836 1179 -2834
rect 1178 -2842 1179 -2840
rect 1185 -2836 1186 -2834
rect 1185 -2842 1186 -2840
rect 1192 -2836 1193 -2834
rect 1192 -2842 1193 -2840
rect 1199 -2836 1200 -2834
rect 1199 -2842 1200 -2840
rect 1206 -2836 1207 -2834
rect 1206 -2842 1207 -2840
rect 1213 -2836 1214 -2834
rect 1213 -2842 1214 -2840
rect 1220 -2836 1221 -2834
rect 1220 -2842 1221 -2840
rect 1227 -2836 1228 -2834
rect 1227 -2842 1228 -2840
rect 1234 -2836 1235 -2834
rect 1234 -2842 1235 -2840
rect 1241 -2836 1242 -2834
rect 1241 -2842 1242 -2840
rect 1248 -2836 1249 -2834
rect 1248 -2842 1249 -2840
rect 1255 -2836 1256 -2834
rect 1258 -2836 1259 -2834
rect 1258 -2842 1259 -2840
rect 1262 -2836 1263 -2834
rect 1262 -2842 1263 -2840
rect 1269 -2836 1270 -2834
rect 1269 -2842 1270 -2840
rect 1276 -2836 1277 -2834
rect 1276 -2842 1277 -2840
rect 1283 -2836 1284 -2834
rect 1286 -2836 1287 -2834
rect 1286 -2842 1287 -2840
rect 1290 -2836 1291 -2834
rect 1290 -2842 1291 -2840
rect 1297 -2836 1298 -2834
rect 1297 -2842 1298 -2840
rect 1304 -2836 1305 -2834
rect 1304 -2842 1305 -2840
rect 1311 -2836 1312 -2834
rect 1314 -2836 1315 -2834
rect 1311 -2842 1312 -2840
rect 1314 -2842 1315 -2840
rect 1318 -2836 1319 -2834
rect 1318 -2842 1319 -2840
rect 1325 -2836 1326 -2834
rect 1325 -2842 1326 -2840
rect 1332 -2836 1333 -2834
rect 1332 -2842 1333 -2840
rect 1339 -2836 1340 -2834
rect 1339 -2842 1340 -2840
rect 1346 -2836 1347 -2834
rect 1346 -2842 1347 -2840
rect 1349 -2842 1350 -2840
rect 1353 -2836 1354 -2834
rect 1353 -2842 1354 -2840
rect 1360 -2836 1361 -2834
rect 1360 -2842 1361 -2840
rect 1367 -2836 1368 -2834
rect 1367 -2842 1368 -2840
rect 1374 -2836 1375 -2834
rect 1374 -2842 1375 -2840
rect 1381 -2836 1382 -2834
rect 1381 -2842 1382 -2840
rect 1391 -2836 1392 -2834
rect 1388 -2842 1389 -2840
rect 1391 -2842 1392 -2840
rect 1395 -2836 1396 -2834
rect 1395 -2842 1396 -2840
rect 1402 -2836 1403 -2834
rect 1402 -2842 1403 -2840
rect 1409 -2836 1410 -2834
rect 1409 -2842 1410 -2840
rect 1416 -2836 1417 -2834
rect 1416 -2842 1417 -2840
rect 1423 -2836 1424 -2834
rect 1423 -2842 1424 -2840
rect 1433 -2836 1434 -2834
rect 1430 -2842 1431 -2840
rect 1433 -2842 1434 -2840
rect 1437 -2836 1438 -2834
rect 1437 -2842 1438 -2840
rect 1444 -2836 1445 -2834
rect 1444 -2842 1445 -2840
rect 1451 -2836 1452 -2834
rect 1451 -2842 1452 -2840
rect 1458 -2836 1459 -2834
rect 1458 -2842 1459 -2840
rect 1465 -2836 1466 -2834
rect 1465 -2842 1466 -2840
rect 1472 -2836 1473 -2834
rect 1472 -2842 1473 -2840
rect 1479 -2836 1480 -2834
rect 1479 -2842 1480 -2840
rect 1489 -2836 1490 -2834
rect 1486 -2842 1487 -2840
rect 1489 -2842 1490 -2840
rect 1493 -2836 1494 -2834
rect 1496 -2836 1497 -2834
rect 1493 -2842 1494 -2840
rect 1496 -2842 1497 -2840
rect 1500 -2836 1501 -2834
rect 1500 -2842 1501 -2840
rect 1507 -2836 1508 -2834
rect 1507 -2842 1508 -2840
rect 1514 -2836 1515 -2834
rect 1514 -2842 1515 -2840
rect 1521 -2836 1522 -2834
rect 1521 -2842 1522 -2840
rect 1528 -2836 1529 -2834
rect 1528 -2842 1529 -2840
rect 1535 -2836 1536 -2834
rect 1535 -2842 1536 -2840
rect 1542 -2836 1543 -2834
rect 1542 -2842 1543 -2840
rect 1549 -2836 1550 -2834
rect 1549 -2842 1550 -2840
rect 1556 -2836 1557 -2834
rect 1556 -2842 1557 -2840
rect 1563 -2842 1564 -2840
rect 1566 -2842 1567 -2840
rect 1570 -2836 1571 -2834
rect 1570 -2842 1571 -2840
rect 1577 -2836 1578 -2834
rect 1577 -2842 1578 -2840
rect 1584 -2836 1585 -2834
rect 1584 -2842 1585 -2840
rect 1591 -2836 1592 -2834
rect 1591 -2842 1592 -2840
rect 1598 -2836 1599 -2834
rect 1598 -2842 1599 -2840
rect 1605 -2836 1606 -2834
rect 1605 -2842 1606 -2840
rect 1612 -2836 1613 -2834
rect 1612 -2842 1613 -2840
rect 1619 -2836 1620 -2834
rect 1619 -2842 1620 -2840
rect 1626 -2836 1627 -2834
rect 1626 -2842 1627 -2840
rect 1633 -2836 1634 -2834
rect 1633 -2842 1634 -2840
rect 1640 -2836 1641 -2834
rect 1640 -2842 1641 -2840
rect 1647 -2836 1648 -2834
rect 1647 -2842 1648 -2840
rect 1654 -2836 1655 -2834
rect 1654 -2842 1655 -2840
rect 1661 -2836 1662 -2834
rect 1661 -2842 1662 -2840
rect 1668 -2836 1669 -2834
rect 1668 -2842 1669 -2840
rect 1675 -2836 1676 -2834
rect 1675 -2842 1676 -2840
rect 1685 -2836 1686 -2834
rect 1682 -2842 1683 -2840
rect 1685 -2842 1686 -2840
rect 1689 -2836 1690 -2834
rect 1689 -2842 1690 -2840
rect 1696 -2836 1697 -2834
rect 1696 -2842 1697 -2840
rect 1706 -2836 1707 -2834
rect 1703 -2842 1704 -2840
rect 1706 -2842 1707 -2840
rect 1710 -2836 1711 -2834
rect 1710 -2842 1711 -2840
rect 1717 -2836 1718 -2834
rect 1717 -2842 1718 -2840
rect 1724 -2836 1725 -2834
rect 1724 -2842 1725 -2840
rect 1731 -2836 1732 -2834
rect 1731 -2842 1732 -2840
rect 1738 -2836 1739 -2834
rect 1738 -2842 1739 -2840
rect 1745 -2836 1746 -2834
rect 1745 -2842 1746 -2840
rect 1755 -2836 1756 -2834
rect 1752 -2842 1753 -2840
rect 1755 -2842 1756 -2840
rect 1759 -2836 1760 -2834
rect 1759 -2842 1760 -2840
rect 1766 -2836 1767 -2834
rect 1766 -2842 1767 -2840
rect 1773 -2836 1774 -2834
rect 1773 -2842 1774 -2840
rect 1780 -2836 1781 -2834
rect 1780 -2842 1781 -2840
rect 1787 -2836 1788 -2834
rect 1787 -2842 1788 -2840
rect 1794 -2836 1795 -2834
rect 1794 -2842 1795 -2840
rect 1801 -2836 1802 -2834
rect 1801 -2842 1802 -2840
rect 1808 -2836 1809 -2834
rect 1808 -2842 1809 -2840
rect 1815 -2836 1816 -2834
rect 1815 -2842 1816 -2840
rect 1822 -2836 1823 -2834
rect 1822 -2842 1823 -2840
rect 1829 -2836 1830 -2834
rect 1829 -2842 1830 -2840
rect 1836 -2836 1837 -2834
rect 1836 -2842 1837 -2840
rect 1843 -2836 1844 -2834
rect 1843 -2842 1844 -2840
rect 1850 -2836 1851 -2834
rect 1850 -2842 1851 -2840
rect 1857 -2836 1858 -2834
rect 1857 -2842 1858 -2840
rect 1864 -2836 1865 -2834
rect 1864 -2842 1865 -2840
rect 1871 -2836 1872 -2834
rect 1871 -2842 1872 -2840
rect 1878 -2836 1879 -2834
rect 1878 -2842 1879 -2840
rect 1885 -2836 1886 -2834
rect 1885 -2842 1886 -2840
rect 1892 -2836 1893 -2834
rect 1892 -2842 1893 -2840
rect 1899 -2836 1900 -2834
rect 1899 -2842 1900 -2840
rect 1906 -2836 1907 -2834
rect 1906 -2842 1907 -2840
rect 1913 -2836 1914 -2834
rect 1913 -2842 1914 -2840
rect 1920 -2836 1921 -2834
rect 1920 -2842 1921 -2840
rect 1927 -2836 1928 -2834
rect 1927 -2842 1928 -2840
rect 1934 -2836 1935 -2834
rect 1934 -2842 1935 -2840
rect 1941 -2836 1942 -2834
rect 1941 -2842 1942 -2840
rect 1948 -2836 1949 -2834
rect 1948 -2842 1949 -2840
rect 1955 -2836 1956 -2834
rect 1955 -2842 1956 -2840
rect 1962 -2836 1963 -2834
rect 1962 -2842 1963 -2840
rect 1969 -2836 1970 -2834
rect 1969 -2842 1970 -2840
rect 1976 -2836 1977 -2834
rect 1976 -2842 1977 -2840
rect 1983 -2836 1984 -2834
rect 1983 -2842 1984 -2840
rect 1990 -2836 1991 -2834
rect 1990 -2842 1991 -2840
rect 1997 -2836 1998 -2834
rect 1997 -2842 1998 -2840
rect 2004 -2836 2005 -2834
rect 2004 -2842 2005 -2840
rect 2011 -2836 2012 -2834
rect 2011 -2842 2012 -2840
rect 2018 -2836 2019 -2834
rect 2018 -2842 2019 -2840
rect 2025 -2836 2026 -2834
rect 2025 -2842 2026 -2840
rect 2032 -2836 2033 -2834
rect 2032 -2842 2033 -2840
rect 2039 -2836 2040 -2834
rect 2039 -2842 2040 -2840
rect 2046 -2836 2047 -2834
rect 2046 -2842 2047 -2840
rect 2053 -2836 2054 -2834
rect 2053 -2842 2054 -2840
rect 2060 -2836 2061 -2834
rect 2060 -2842 2061 -2840
rect 2067 -2836 2068 -2834
rect 2067 -2842 2068 -2840
rect 2074 -2836 2075 -2834
rect 2074 -2842 2075 -2840
rect 2081 -2836 2082 -2834
rect 2081 -2842 2082 -2840
rect 2088 -2836 2089 -2834
rect 2088 -2842 2089 -2840
rect 2095 -2836 2096 -2834
rect 2095 -2842 2096 -2840
rect 2102 -2836 2103 -2834
rect 2102 -2842 2103 -2840
rect 2109 -2836 2110 -2834
rect 2109 -2842 2110 -2840
rect 2116 -2836 2117 -2834
rect 2116 -2842 2117 -2840
rect 2123 -2836 2124 -2834
rect 2123 -2842 2124 -2840
rect 2130 -2836 2131 -2834
rect 2130 -2842 2131 -2840
rect 2137 -2836 2138 -2834
rect 2137 -2842 2138 -2840
rect 2144 -2836 2145 -2834
rect 2144 -2842 2145 -2840
rect 2151 -2836 2152 -2834
rect 2151 -2842 2152 -2840
rect 2158 -2836 2159 -2834
rect 2158 -2842 2159 -2840
rect 2165 -2836 2166 -2834
rect 2165 -2842 2166 -2840
rect 2172 -2836 2173 -2834
rect 2172 -2842 2173 -2840
rect 2179 -2836 2180 -2834
rect 2179 -2842 2180 -2840
rect 2186 -2836 2187 -2834
rect 2186 -2842 2187 -2840
rect 2193 -2836 2194 -2834
rect 2193 -2842 2194 -2840
rect 2200 -2836 2201 -2834
rect 2200 -2842 2201 -2840
rect 2207 -2836 2208 -2834
rect 2207 -2842 2208 -2840
rect 2214 -2836 2215 -2834
rect 2214 -2842 2215 -2840
rect 2221 -2836 2222 -2834
rect 2224 -2836 2225 -2834
rect 2221 -2842 2222 -2840
rect 2224 -2842 2225 -2840
rect 2228 -2836 2229 -2834
rect 2228 -2842 2229 -2840
rect 2235 -2836 2236 -2834
rect 2235 -2842 2236 -2840
rect 2242 -2836 2243 -2834
rect 2242 -2842 2243 -2840
rect 2249 -2836 2250 -2834
rect 2249 -2842 2250 -2840
rect 2259 -2836 2260 -2834
rect 2256 -2842 2257 -2840
rect 2259 -2842 2260 -2840
rect 2263 -2836 2264 -2834
rect 2263 -2842 2264 -2840
rect 2270 -2836 2271 -2834
rect 2270 -2842 2271 -2840
rect 16 -2981 17 -2979
rect 16 -2987 17 -2985
rect 23 -2981 24 -2979
rect 23 -2987 24 -2985
rect 30 -2981 31 -2979
rect 30 -2987 31 -2985
rect 37 -2981 38 -2979
rect 37 -2987 38 -2985
rect 44 -2981 45 -2979
rect 44 -2987 45 -2985
rect 54 -2981 55 -2979
rect 51 -2987 52 -2985
rect 58 -2981 59 -2979
rect 58 -2987 59 -2985
rect 65 -2981 66 -2979
rect 65 -2987 66 -2985
rect 72 -2981 73 -2979
rect 72 -2987 73 -2985
rect 79 -2981 80 -2979
rect 79 -2987 80 -2985
rect 86 -2981 87 -2979
rect 86 -2987 87 -2985
rect 93 -2981 94 -2979
rect 93 -2987 94 -2985
rect 100 -2981 101 -2979
rect 103 -2981 104 -2979
rect 100 -2987 101 -2985
rect 103 -2987 104 -2985
rect 110 -2981 111 -2979
rect 110 -2987 111 -2985
rect 114 -2981 115 -2979
rect 117 -2981 118 -2979
rect 117 -2987 118 -2985
rect 121 -2981 122 -2979
rect 124 -2981 125 -2979
rect 121 -2987 122 -2985
rect 124 -2987 125 -2985
rect 128 -2981 129 -2979
rect 128 -2987 129 -2985
rect 135 -2981 136 -2979
rect 135 -2987 136 -2985
rect 142 -2981 143 -2979
rect 142 -2987 143 -2985
rect 149 -2981 150 -2979
rect 149 -2987 150 -2985
rect 159 -2981 160 -2979
rect 156 -2987 157 -2985
rect 159 -2987 160 -2985
rect 163 -2981 164 -2979
rect 163 -2987 164 -2985
rect 170 -2981 171 -2979
rect 170 -2987 171 -2985
rect 177 -2981 178 -2979
rect 177 -2987 178 -2985
rect 184 -2981 185 -2979
rect 184 -2987 185 -2985
rect 191 -2981 192 -2979
rect 191 -2987 192 -2985
rect 198 -2981 199 -2979
rect 198 -2987 199 -2985
rect 205 -2981 206 -2979
rect 205 -2987 206 -2985
rect 212 -2981 213 -2979
rect 215 -2981 216 -2979
rect 212 -2987 213 -2985
rect 215 -2987 216 -2985
rect 219 -2981 220 -2979
rect 219 -2987 220 -2985
rect 226 -2981 227 -2979
rect 226 -2987 227 -2985
rect 233 -2981 234 -2979
rect 233 -2987 234 -2985
rect 240 -2981 241 -2979
rect 240 -2987 241 -2985
rect 247 -2981 248 -2979
rect 247 -2987 248 -2985
rect 254 -2981 255 -2979
rect 257 -2981 258 -2979
rect 254 -2987 255 -2985
rect 261 -2981 262 -2979
rect 261 -2987 262 -2985
rect 268 -2981 269 -2979
rect 268 -2987 269 -2985
rect 275 -2981 276 -2979
rect 275 -2987 276 -2985
rect 282 -2981 283 -2979
rect 282 -2987 283 -2985
rect 289 -2981 290 -2979
rect 289 -2987 290 -2985
rect 296 -2981 297 -2979
rect 296 -2987 297 -2985
rect 303 -2981 304 -2979
rect 303 -2987 304 -2985
rect 310 -2981 311 -2979
rect 310 -2987 311 -2985
rect 317 -2981 318 -2979
rect 317 -2987 318 -2985
rect 324 -2981 325 -2979
rect 324 -2987 325 -2985
rect 331 -2981 332 -2979
rect 331 -2987 332 -2985
rect 338 -2981 339 -2979
rect 338 -2987 339 -2985
rect 345 -2981 346 -2979
rect 345 -2987 346 -2985
rect 352 -2981 353 -2979
rect 352 -2987 353 -2985
rect 359 -2981 360 -2979
rect 359 -2987 360 -2985
rect 366 -2981 367 -2979
rect 366 -2987 367 -2985
rect 373 -2981 374 -2979
rect 373 -2987 374 -2985
rect 380 -2981 381 -2979
rect 380 -2987 381 -2985
rect 387 -2981 388 -2979
rect 387 -2987 388 -2985
rect 394 -2981 395 -2979
rect 394 -2987 395 -2985
rect 401 -2981 402 -2979
rect 401 -2987 402 -2985
rect 408 -2981 409 -2979
rect 408 -2987 409 -2985
rect 415 -2981 416 -2979
rect 415 -2987 416 -2985
rect 422 -2981 423 -2979
rect 422 -2987 423 -2985
rect 429 -2981 430 -2979
rect 429 -2987 430 -2985
rect 436 -2981 437 -2979
rect 436 -2987 437 -2985
rect 443 -2981 444 -2979
rect 443 -2987 444 -2985
rect 450 -2981 451 -2979
rect 450 -2987 451 -2985
rect 457 -2981 458 -2979
rect 457 -2987 458 -2985
rect 464 -2981 465 -2979
rect 467 -2981 468 -2979
rect 471 -2981 472 -2979
rect 471 -2987 472 -2985
rect 478 -2981 479 -2979
rect 478 -2987 479 -2985
rect 485 -2981 486 -2979
rect 485 -2987 486 -2985
rect 492 -2981 493 -2979
rect 492 -2987 493 -2985
rect 499 -2981 500 -2979
rect 499 -2987 500 -2985
rect 506 -2981 507 -2979
rect 506 -2987 507 -2985
rect 513 -2981 514 -2979
rect 513 -2987 514 -2985
rect 520 -2981 521 -2979
rect 520 -2987 521 -2985
rect 527 -2981 528 -2979
rect 527 -2987 528 -2985
rect 534 -2981 535 -2979
rect 534 -2987 535 -2985
rect 541 -2981 542 -2979
rect 544 -2981 545 -2979
rect 541 -2987 542 -2985
rect 544 -2987 545 -2985
rect 548 -2981 549 -2979
rect 548 -2987 549 -2985
rect 555 -2981 556 -2979
rect 555 -2987 556 -2985
rect 562 -2981 563 -2979
rect 565 -2981 566 -2979
rect 565 -2987 566 -2985
rect 569 -2981 570 -2979
rect 569 -2987 570 -2985
rect 572 -2987 573 -2985
rect 576 -2981 577 -2979
rect 576 -2987 577 -2985
rect 583 -2981 584 -2979
rect 583 -2987 584 -2985
rect 590 -2981 591 -2979
rect 590 -2987 591 -2985
rect 597 -2981 598 -2979
rect 597 -2987 598 -2985
rect 604 -2981 605 -2979
rect 604 -2987 605 -2985
rect 611 -2981 612 -2979
rect 611 -2987 612 -2985
rect 618 -2981 619 -2979
rect 618 -2987 619 -2985
rect 625 -2981 626 -2979
rect 625 -2987 626 -2985
rect 632 -2981 633 -2979
rect 632 -2987 633 -2985
rect 639 -2981 640 -2979
rect 642 -2981 643 -2979
rect 642 -2987 643 -2985
rect 646 -2981 647 -2979
rect 646 -2987 647 -2985
rect 653 -2981 654 -2979
rect 653 -2987 654 -2985
rect 660 -2981 661 -2979
rect 663 -2981 664 -2979
rect 660 -2987 661 -2985
rect 663 -2987 664 -2985
rect 667 -2981 668 -2979
rect 667 -2987 668 -2985
rect 674 -2981 675 -2979
rect 674 -2987 675 -2985
rect 681 -2981 682 -2979
rect 681 -2987 682 -2985
rect 688 -2981 689 -2979
rect 688 -2987 689 -2985
rect 695 -2981 696 -2979
rect 695 -2987 696 -2985
rect 702 -2981 703 -2979
rect 702 -2987 703 -2985
rect 709 -2981 710 -2979
rect 709 -2987 710 -2985
rect 716 -2981 717 -2979
rect 716 -2987 717 -2985
rect 723 -2981 724 -2979
rect 723 -2987 724 -2985
rect 730 -2981 731 -2979
rect 730 -2987 731 -2985
rect 737 -2981 738 -2979
rect 740 -2981 741 -2979
rect 737 -2987 738 -2985
rect 740 -2987 741 -2985
rect 744 -2981 745 -2979
rect 744 -2987 745 -2985
rect 751 -2981 752 -2979
rect 751 -2987 752 -2985
rect 758 -2981 759 -2979
rect 758 -2987 759 -2985
rect 765 -2981 766 -2979
rect 765 -2987 766 -2985
rect 772 -2981 773 -2979
rect 772 -2987 773 -2985
rect 779 -2981 780 -2979
rect 779 -2987 780 -2985
rect 786 -2981 787 -2979
rect 786 -2987 787 -2985
rect 793 -2981 794 -2979
rect 793 -2987 794 -2985
rect 800 -2981 801 -2979
rect 807 -2981 808 -2979
rect 807 -2987 808 -2985
rect 814 -2981 815 -2979
rect 814 -2987 815 -2985
rect 821 -2981 822 -2979
rect 821 -2987 822 -2985
rect 828 -2981 829 -2979
rect 828 -2987 829 -2985
rect 835 -2981 836 -2979
rect 835 -2987 836 -2985
rect 842 -2981 843 -2979
rect 842 -2987 843 -2985
rect 849 -2981 850 -2979
rect 849 -2987 850 -2985
rect 856 -2981 857 -2979
rect 856 -2987 857 -2985
rect 863 -2981 864 -2979
rect 863 -2987 864 -2985
rect 870 -2981 871 -2979
rect 870 -2987 871 -2985
rect 880 -2981 881 -2979
rect 880 -2987 881 -2985
rect 884 -2981 885 -2979
rect 884 -2987 885 -2985
rect 891 -2981 892 -2979
rect 891 -2987 892 -2985
rect 898 -2981 899 -2979
rect 898 -2987 899 -2985
rect 905 -2981 906 -2979
rect 905 -2987 906 -2985
rect 912 -2981 913 -2979
rect 912 -2987 913 -2985
rect 922 -2981 923 -2979
rect 919 -2987 920 -2985
rect 922 -2987 923 -2985
rect 926 -2981 927 -2979
rect 926 -2987 927 -2985
rect 933 -2981 934 -2979
rect 933 -2987 934 -2985
rect 940 -2981 941 -2979
rect 940 -2987 941 -2985
rect 947 -2981 948 -2979
rect 947 -2987 948 -2985
rect 954 -2981 955 -2979
rect 954 -2987 955 -2985
rect 961 -2981 962 -2979
rect 964 -2981 965 -2979
rect 961 -2987 962 -2985
rect 964 -2987 965 -2985
rect 968 -2981 969 -2979
rect 968 -2987 969 -2985
rect 975 -2981 976 -2979
rect 975 -2987 976 -2985
rect 982 -2981 983 -2979
rect 985 -2981 986 -2979
rect 982 -2987 983 -2985
rect 985 -2987 986 -2985
rect 989 -2981 990 -2979
rect 989 -2987 990 -2985
rect 996 -2981 997 -2979
rect 996 -2987 997 -2985
rect 1003 -2981 1004 -2979
rect 1003 -2987 1004 -2985
rect 1010 -2981 1011 -2979
rect 1010 -2987 1011 -2985
rect 1017 -2981 1018 -2979
rect 1017 -2987 1018 -2985
rect 1024 -2981 1025 -2979
rect 1024 -2987 1025 -2985
rect 1031 -2981 1032 -2979
rect 1031 -2987 1032 -2985
rect 1034 -2987 1035 -2985
rect 1038 -2981 1039 -2979
rect 1041 -2981 1042 -2979
rect 1038 -2987 1039 -2985
rect 1041 -2987 1042 -2985
rect 1045 -2981 1046 -2979
rect 1045 -2987 1046 -2985
rect 1055 -2981 1056 -2979
rect 1052 -2987 1053 -2985
rect 1055 -2987 1056 -2985
rect 1059 -2981 1060 -2979
rect 1062 -2981 1063 -2979
rect 1059 -2987 1060 -2985
rect 1062 -2987 1063 -2985
rect 1066 -2981 1067 -2979
rect 1069 -2981 1070 -2979
rect 1066 -2987 1067 -2985
rect 1069 -2987 1070 -2985
rect 1073 -2981 1074 -2979
rect 1073 -2987 1074 -2985
rect 1080 -2981 1081 -2979
rect 1080 -2987 1081 -2985
rect 1087 -2981 1088 -2979
rect 1087 -2987 1088 -2985
rect 1094 -2981 1095 -2979
rect 1097 -2981 1098 -2979
rect 1097 -2987 1098 -2985
rect 1101 -2981 1102 -2979
rect 1101 -2987 1102 -2985
rect 1108 -2981 1109 -2979
rect 1108 -2987 1109 -2985
rect 1115 -2981 1116 -2979
rect 1115 -2987 1116 -2985
rect 1122 -2981 1123 -2979
rect 1125 -2981 1126 -2979
rect 1125 -2987 1126 -2985
rect 1129 -2981 1130 -2979
rect 1129 -2987 1130 -2985
rect 1136 -2981 1137 -2979
rect 1139 -2981 1140 -2979
rect 1136 -2987 1137 -2985
rect 1139 -2987 1140 -2985
rect 1143 -2981 1144 -2979
rect 1143 -2987 1144 -2985
rect 1150 -2981 1151 -2979
rect 1150 -2987 1151 -2985
rect 1157 -2981 1158 -2979
rect 1160 -2981 1161 -2979
rect 1157 -2987 1158 -2985
rect 1160 -2987 1161 -2985
rect 1164 -2981 1165 -2979
rect 1164 -2987 1165 -2985
rect 1171 -2981 1172 -2979
rect 1171 -2987 1172 -2985
rect 1178 -2981 1179 -2979
rect 1178 -2987 1179 -2985
rect 1185 -2981 1186 -2979
rect 1185 -2987 1186 -2985
rect 1192 -2981 1193 -2979
rect 1192 -2987 1193 -2985
rect 1199 -2981 1200 -2979
rect 1202 -2981 1203 -2979
rect 1199 -2987 1200 -2985
rect 1202 -2987 1203 -2985
rect 1206 -2981 1207 -2979
rect 1209 -2981 1210 -2979
rect 1209 -2987 1210 -2985
rect 1213 -2981 1214 -2979
rect 1213 -2987 1214 -2985
rect 1220 -2981 1221 -2979
rect 1220 -2987 1221 -2985
rect 1227 -2981 1228 -2979
rect 1227 -2987 1228 -2985
rect 1234 -2981 1235 -2979
rect 1234 -2987 1235 -2985
rect 1241 -2981 1242 -2979
rect 1241 -2987 1242 -2985
rect 1248 -2981 1249 -2979
rect 1248 -2987 1249 -2985
rect 1255 -2981 1256 -2979
rect 1255 -2987 1256 -2985
rect 1262 -2981 1263 -2979
rect 1262 -2987 1263 -2985
rect 1269 -2981 1270 -2979
rect 1269 -2987 1270 -2985
rect 1276 -2981 1277 -2979
rect 1276 -2987 1277 -2985
rect 1283 -2981 1284 -2979
rect 1283 -2987 1284 -2985
rect 1290 -2981 1291 -2979
rect 1290 -2987 1291 -2985
rect 1297 -2981 1298 -2979
rect 1297 -2987 1298 -2985
rect 1304 -2981 1305 -2979
rect 1304 -2987 1305 -2985
rect 1314 -2981 1315 -2979
rect 1311 -2987 1312 -2985
rect 1314 -2987 1315 -2985
rect 1318 -2981 1319 -2979
rect 1318 -2987 1319 -2985
rect 1325 -2981 1326 -2979
rect 1325 -2987 1326 -2985
rect 1332 -2981 1333 -2979
rect 1332 -2987 1333 -2985
rect 1339 -2981 1340 -2979
rect 1339 -2987 1340 -2985
rect 1346 -2981 1347 -2979
rect 1346 -2987 1347 -2985
rect 1353 -2981 1354 -2979
rect 1353 -2987 1354 -2985
rect 1360 -2981 1361 -2979
rect 1363 -2981 1364 -2979
rect 1363 -2987 1364 -2985
rect 1367 -2981 1368 -2979
rect 1367 -2987 1368 -2985
rect 1374 -2981 1375 -2979
rect 1374 -2987 1375 -2985
rect 1381 -2981 1382 -2979
rect 1381 -2987 1382 -2985
rect 1388 -2981 1389 -2979
rect 1388 -2987 1389 -2985
rect 1395 -2981 1396 -2979
rect 1395 -2987 1396 -2985
rect 1402 -2981 1403 -2979
rect 1402 -2987 1403 -2985
rect 1409 -2981 1410 -2979
rect 1409 -2987 1410 -2985
rect 1419 -2981 1420 -2979
rect 1416 -2987 1417 -2985
rect 1419 -2987 1420 -2985
rect 1423 -2981 1424 -2979
rect 1423 -2987 1424 -2985
rect 1430 -2981 1431 -2979
rect 1430 -2987 1431 -2985
rect 1437 -2981 1438 -2979
rect 1437 -2987 1438 -2985
rect 1444 -2981 1445 -2979
rect 1444 -2987 1445 -2985
rect 1451 -2981 1452 -2979
rect 1451 -2987 1452 -2985
rect 1458 -2981 1459 -2979
rect 1458 -2987 1459 -2985
rect 1465 -2981 1466 -2979
rect 1465 -2987 1466 -2985
rect 1472 -2981 1473 -2979
rect 1472 -2987 1473 -2985
rect 1479 -2981 1480 -2979
rect 1479 -2987 1480 -2985
rect 1486 -2981 1487 -2979
rect 1486 -2987 1487 -2985
rect 1493 -2981 1494 -2979
rect 1493 -2987 1494 -2985
rect 1500 -2981 1501 -2979
rect 1500 -2987 1501 -2985
rect 1507 -2981 1508 -2979
rect 1507 -2987 1508 -2985
rect 1514 -2981 1515 -2979
rect 1514 -2987 1515 -2985
rect 1521 -2981 1522 -2979
rect 1521 -2987 1522 -2985
rect 1528 -2981 1529 -2979
rect 1528 -2987 1529 -2985
rect 1535 -2981 1536 -2979
rect 1535 -2987 1536 -2985
rect 1542 -2981 1543 -2979
rect 1542 -2987 1543 -2985
rect 1549 -2981 1550 -2979
rect 1549 -2987 1550 -2985
rect 1556 -2981 1557 -2979
rect 1556 -2987 1557 -2985
rect 1563 -2981 1564 -2979
rect 1563 -2987 1564 -2985
rect 1570 -2981 1571 -2979
rect 1570 -2987 1571 -2985
rect 1573 -2987 1574 -2985
rect 1577 -2981 1578 -2979
rect 1577 -2987 1578 -2985
rect 1584 -2981 1585 -2979
rect 1584 -2987 1585 -2985
rect 1591 -2981 1592 -2979
rect 1591 -2987 1592 -2985
rect 1598 -2981 1599 -2979
rect 1598 -2987 1599 -2985
rect 1605 -2981 1606 -2979
rect 1605 -2987 1606 -2985
rect 1612 -2981 1613 -2979
rect 1612 -2987 1613 -2985
rect 1619 -2981 1620 -2979
rect 1619 -2987 1620 -2985
rect 1626 -2981 1627 -2979
rect 1626 -2987 1627 -2985
rect 1633 -2981 1634 -2979
rect 1633 -2987 1634 -2985
rect 1640 -2981 1641 -2979
rect 1640 -2987 1641 -2985
rect 1647 -2981 1648 -2979
rect 1647 -2987 1648 -2985
rect 1654 -2981 1655 -2979
rect 1654 -2987 1655 -2985
rect 1661 -2981 1662 -2979
rect 1661 -2987 1662 -2985
rect 1668 -2981 1669 -2979
rect 1668 -2987 1669 -2985
rect 1675 -2981 1676 -2979
rect 1675 -2987 1676 -2985
rect 1682 -2981 1683 -2979
rect 1682 -2987 1683 -2985
rect 1689 -2981 1690 -2979
rect 1689 -2987 1690 -2985
rect 1696 -2981 1697 -2979
rect 1696 -2987 1697 -2985
rect 1703 -2981 1704 -2979
rect 1703 -2987 1704 -2985
rect 1710 -2981 1711 -2979
rect 1710 -2987 1711 -2985
rect 1717 -2981 1718 -2979
rect 1717 -2987 1718 -2985
rect 1724 -2981 1725 -2979
rect 1724 -2987 1725 -2985
rect 1731 -2981 1732 -2979
rect 1731 -2987 1732 -2985
rect 1738 -2981 1739 -2979
rect 1738 -2987 1739 -2985
rect 1745 -2981 1746 -2979
rect 1745 -2987 1746 -2985
rect 1752 -2981 1753 -2979
rect 1752 -2987 1753 -2985
rect 1759 -2981 1760 -2979
rect 1759 -2987 1760 -2985
rect 1766 -2987 1767 -2985
rect 1769 -2987 1770 -2985
rect 1773 -2981 1774 -2979
rect 1773 -2987 1774 -2985
rect 1780 -2981 1781 -2979
rect 1780 -2987 1781 -2985
rect 1787 -2981 1788 -2979
rect 1787 -2987 1788 -2985
rect 1794 -2981 1795 -2979
rect 1794 -2987 1795 -2985
rect 1801 -2981 1802 -2979
rect 1801 -2987 1802 -2985
rect 1808 -2981 1809 -2979
rect 1808 -2987 1809 -2985
rect 1815 -2981 1816 -2979
rect 1815 -2987 1816 -2985
rect 1822 -2981 1823 -2979
rect 1822 -2987 1823 -2985
rect 1829 -2981 1830 -2979
rect 1829 -2987 1830 -2985
rect 1836 -2981 1837 -2979
rect 1836 -2987 1837 -2985
rect 1843 -2981 1844 -2979
rect 1843 -2987 1844 -2985
rect 1850 -2981 1851 -2979
rect 1850 -2987 1851 -2985
rect 1857 -2981 1858 -2979
rect 1857 -2987 1858 -2985
rect 1864 -2981 1865 -2979
rect 1864 -2987 1865 -2985
rect 1871 -2981 1872 -2979
rect 1871 -2987 1872 -2985
rect 1874 -2987 1875 -2985
rect 1878 -2981 1879 -2979
rect 1878 -2987 1879 -2985
rect 1885 -2981 1886 -2979
rect 1885 -2987 1886 -2985
rect 1892 -2981 1893 -2979
rect 1892 -2987 1893 -2985
rect 1899 -2981 1900 -2979
rect 1899 -2987 1900 -2985
rect 1906 -2981 1907 -2979
rect 1906 -2987 1907 -2985
rect 1913 -2981 1914 -2979
rect 1913 -2987 1914 -2985
rect 1920 -2981 1921 -2979
rect 1920 -2987 1921 -2985
rect 1927 -2981 1928 -2979
rect 1927 -2987 1928 -2985
rect 1934 -2981 1935 -2979
rect 1934 -2987 1935 -2985
rect 1941 -2981 1942 -2979
rect 1941 -2987 1942 -2985
rect 1948 -2981 1949 -2979
rect 1948 -2987 1949 -2985
rect 1955 -2981 1956 -2979
rect 1955 -2987 1956 -2985
rect 1962 -2981 1963 -2979
rect 1962 -2987 1963 -2985
rect 1969 -2981 1970 -2979
rect 1969 -2987 1970 -2985
rect 1976 -2981 1977 -2979
rect 1976 -2987 1977 -2985
rect 1983 -2981 1984 -2979
rect 1983 -2987 1984 -2985
rect 1990 -2981 1991 -2979
rect 1990 -2987 1991 -2985
rect 1997 -2981 1998 -2979
rect 1997 -2987 1998 -2985
rect 2004 -2981 2005 -2979
rect 2004 -2987 2005 -2985
rect 2011 -2981 2012 -2979
rect 2011 -2987 2012 -2985
rect 2018 -2981 2019 -2979
rect 2018 -2987 2019 -2985
rect 2025 -2981 2026 -2979
rect 2025 -2987 2026 -2985
rect 2032 -2981 2033 -2979
rect 2032 -2987 2033 -2985
rect 2039 -2981 2040 -2979
rect 2039 -2987 2040 -2985
rect 2046 -2981 2047 -2979
rect 2046 -2987 2047 -2985
rect 2053 -2981 2054 -2979
rect 2053 -2987 2054 -2985
rect 2060 -2981 2061 -2979
rect 2060 -2987 2061 -2985
rect 2067 -2981 2068 -2979
rect 2067 -2987 2068 -2985
rect 2074 -2981 2075 -2979
rect 2074 -2987 2075 -2985
rect 2081 -2981 2082 -2979
rect 2081 -2987 2082 -2985
rect 2088 -2981 2089 -2979
rect 2088 -2987 2089 -2985
rect 2095 -2981 2096 -2979
rect 2098 -2981 2099 -2979
rect 2095 -2987 2096 -2985
rect 2098 -2987 2099 -2985
rect 2102 -2981 2103 -2979
rect 2102 -2987 2103 -2985
rect 2109 -2981 2110 -2979
rect 2109 -2987 2110 -2985
rect 2116 -2981 2117 -2979
rect 2116 -2987 2117 -2985
rect 2123 -2981 2124 -2979
rect 2123 -2987 2124 -2985
rect 2130 -2981 2131 -2979
rect 2130 -2987 2131 -2985
rect 2137 -2981 2138 -2979
rect 2137 -2987 2138 -2985
rect 2144 -2981 2145 -2979
rect 2144 -2987 2145 -2985
rect 2151 -2981 2152 -2979
rect 2151 -2987 2152 -2985
rect 23 -3096 24 -3094
rect 23 -3102 24 -3100
rect 30 -3096 31 -3094
rect 30 -3102 31 -3100
rect 37 -3096 38 -3094
rect 37 -3102 38 -3100
rect 58 -3096 59 -3094
rect 58 -3102 59 -3100
rect 65 -3096 66 -3094
rect 65 -3102 66 -3100
rect 72 -3096 73 -3094
rect 72 -3102 73 -3100
rect 79 -3102 80 -3100
rect 82 -3102 83 -3100
rect 86 -3096 87 -3094
rect 86 -3102 87 -3100
rect 93 -3096 94 -3094
rect 100 -3096 101 -3094
rect 100 -3102 101 -3100
rect 107 -3096 108 -3094
rect 107 -3102 108 -3100
rect 114 -3096 115 -3094
rect 114 -3102 115 -3100
rect 121 -3096 122 -3094
rect 121 -3102 122 -3100
rect 131 -3096 132 -3094
rect 128 -3102 129 -3100
rect 131 -3102 132 -3100
rect 138 -3096 139 -3094
rect 135 -3102 136 -3100
rect 138 -3102 139 -3100
rect 142 -3096 143 -3094
rect 142 -3102 143 -3100
rect 149 -3096 150 -3094
rect 149 -3102 150 -3100
rect 156 -3096 157 -3094
rect 156 -3102 157 -3100
rect 166 -3096 167 -3094
rect 163 -3102 164 -3100
rect 166 -3102 167 -3100
rect 173 -3096 174 -3094
rect 170 -3102 171 -3100
rect 173 -3102 174 -3100
rect 177 -3096 178 -3094
rect 177 -3102 178 -3100
rect 184 -3096 185 -3094
rect 184 -3102 185 -3100
rect 191 -3096 192 -3094
rect 191 -3102 192 -3100
rect 198 -3096 199 -3094
rect 198 -3102 199 -3100
rect 205 -3096 206 -3094
rect 208 -3096 209 -3094
rect 205 -3102 206 -3100
rect 208 -3102 209 -3100
rect 212 -3096 213 -3094
rect 212 -3102 213 -3100
rect 219 -3096 220 -3094
rect 219 -3102 220 -3100
rect 226 -3096 227 -3094
rect 226 -3102 227 -3100
rect 236 -3096 237 -3094
rect 236 -3102 237 -3100
rect 240 -3096 241 -3094
rect 240 -3102 241 -3100
rect 247 -3096 248 -3094
rect 247 -3102 248 -3100
rect 254 -3096 255 -3094
rect 254 -3102 255 -3100
rect 261 -3096 262 -3094
rect 261 -3102 262 -3100
rect 268 -3096 269 -3094
rect 268 -3102 269 -3100
rect 275 -3096 276 -3094
rect 275 -3102 276 -3100
rect 282 -3096 283 -3094
rect 282 -3102 283 -3100
rect 289 -3096 290 -3094
rect 289 -3102 290 -3100
rect 296 -3096 297 -3094
rect 296 -3102 297 -3100
rect 303 -3096 304 -3094
rect 303 -3102 304 -3100
rect 310 -3096 311 -3094
rect 310 -3102 311 -3100
rect 317 -3096 318 -3094
rect 317 -3102 318 -3100
rect 324 -3096 325 -3094
rect 324 -3102 325 -3100
rect 331 -3096 332 -3094
rect 331 -3102 332 -3100
rect 338 -3096 339 -3094
rect 338 -3102 339 -3100
rect 345 -3096 346 -3094
rect 345 -3102 346 -3100
rect 352 -3096 353 -3094
rect 352 -3102 353 -3100
rect 359 -3096 360 -3094
rect 359 -3102 360 -3100
rect 366 -3096 367 -3094
rect 366 -3102 367 -3100
rect 373 -3096 374 -3094
rect 373 -3102 374 -3100
rect 380 -3096 381 -3094
rect 380 -3102 381 -3100
rect 387 -3096 388 -3094
rect 387 -3102 388 -3100
rect 394 -3096 395 -3094
rect 394 -3102 395 -3100
rect 401 -3096 402 -3094
rect 401 -3102 402 -3100
rect 408 -3096 409 -3094
rect 408 -3102 409 -3100
rect 415 -3096 416 -3094
rect 415 -3102 416 -3100
rect 422 -3096 423 -3094
rect 422 -3102 423 -3100
rect 429 -3096 430 -3094
rect 429 -3102 430 -3100
rect 436 -3096 437 -3094
rect 436 -3102 437 -3100
rect 443 -3096 444 -3094
rect 443 -3102 444 -3100
rect 450 -3096 451 -3094
rect 450 -3102 451 -3100
rect 457 -3096 458 -3094
rect 460 -3096 461 -3094
rect 457 -3102 458 -3100
rect 460 -3102 461 -3100
rect 464 -3096 465 -3094
rect 464 -3102 465 -3100
rect 471 -3096 472 -3094
rect 471 -3102 472 -3100
rect 478 -3096 479 -3094
rect 478 -3102 479 -3100
rect 485 -3096 486 -3094
rect 485 -3102 486 -3100
rect 492 -3096 493 -3094
rect 492 -3102 493 -3100
rect 499 -3096 500 -3094
rect 499 -3102 500 -3100
rect 506 -3096 507 -3094
rect 506 -3102 507 -3100
rect 513 -3096 514 -3094
rect 513 -3102 514 -3100
rect 520 -3096 521 -3094
rect 520 -3102 521 -3100
rect 527 -3102 528 -3100
rect 530 -3102 531 -3100
rect 534 -3096 535 -3094
rect 534 -3102 535 -3100
rect 541 -3096 542 -3094
rect 541 -3102 542 -3100
rect 548 -3096 549 -3094
rect 548 -3102 549 -3100
rect 555 -3096 556 -3094
rect 555 -3102 556 -3100
rect 562 -3096 563 -3094
rect 562 -3102 563 -3100
rect 569 -3096 570 -3094
rect 569 -3102 570 -3100
rect 576 -3096 577 -3094
rect 576 -3102 577 -3100
rect 583 -3096 584 -3094
rect 583 -3102 584 -3100
rect 590 -3096 591 -3094
rect 590 -3102 591 -3100
rect 597 -3096 598 -3094
rect 597 -3102 598 -3100
rect 604 -3096 605 -3094
rect 604 -3102 605 -3100
rect 611 -3096 612 -3094
rect 614 -3096 615 -3094
rect 611 -3102 612 -3100
rect 614 -3102 615 -3100
rect 618 -3096 619 -3094
rect 618 -3102 619 -3100
rect 625 -3096 626 -3094
rect 625 -3102 626 -3100
rect 632 -3096 633 -3094
rect 632 -3102 633 -3100
rect 639 -3096 640 -3094
rect 639 -3102 640 -3100
rect 646 -3096 647 -3094
rect 646 -3102 647 -3100
rect 653 -3096 654 -3094
rect 653 -3102 654 -3100
rect 660 -3096 661 -3094
rect 660 -3102 661 -3100
rect 667 -3096 668 -3094
rect 667 -3102 668 -3100
rect 674 -3096 675 -3094
rect 674 -3102 675 -3100
rect 681 -3096 682 -3094
rect 681 -3102 682 -3100
rect 688 -3096 689 -3094
rect 688 -3102 689 -3100
rect 695 -3096 696 -3094
rect 695 -3102 696 -3100
rect 702 -3096 703 -3094
rect 702 -3102 703 -3100
rect 709 -3096 710 -3094
rect 709 -3102 710 -3100
rect 716 -3096 717 -3094
rect 716 -3102 717 -3100
rect 723 -3096 724 -3094
rect 723 -3102 724 -3100
rect 730 -3096 731 -3094
rect 730 -3102 731 -3100
rect 737 -3096 738 -3094
rect 737 -3102 738 -3100
rect 744 -3096 745 -3094
rect 744 -3102 745 -3100
rect 751 -3096 752 -3094
rect 751 -3102 752 -3100
rect 758 -3096 759 -3094
rect 758 -3102 759 -3100
rect 765 -3096 766 -3094
rect 765 -3102 766 -3100
rect 772 -3096 773 -3094
rect 772 -3102 773 -3100
rect 779 -3096 780 -3094
rect 779 -3102 780 -3100
rect 786 -3096 787 -3094
rect 786 -3102 787 -3100
rect 793 -3096 794 -3094
rect 793 -3102 794 -3100
rect 800 -3102 801 -3100
rect 807 -3096 808 -3094
rect 807 -3102 808 -3100
rect 817 -3096 818 -3094
rect 814 -3102 815 -3100
rect 817 -3102 818 -3100
rect 821 -3096 822 -3094
rect 821 -3102 822 -3100
rect 828 -3096 829 -3094
rect 828 -3102 829 -3100
rect 835 -3096 836 -3094
rect 835 -3102 836 -3100
rect 842 -3096 843 -3094
rect 842 -3102 843 -3100
rect 849 -3096 850 -3094
rect 849 -3102 850 -3100
rect 856 -3096 857 -3094
rect 856 -3102 857 -3100
rect 863 -3096 864 -3094
rect 866 -3102 867 -3100
rect 870 -3096 871 -3094
rect 870 -3102 871 -3100
rect 877 -3096 878 -3094
rect 880 -3096 881 -3094
rect 877 -3102 878 -3100
rect 880 -3102 881 -3100
rect 884 -3096 885 -3094
rect 884 -3102 885 -3100
rect 894 -3096 895 -3094
rect 891 -3102 892 -3100
rect 898 -3096 899 -3094
rect 898 -3102 899 -3100
rect 905 -3096 906 -3094
rect 905 -3102 906 -3100
rect 912 -3096 913 -3094
rect 915 -3096 916 -3094
rect 912 -3102 913 -3100
rect 919 -3096 920 -3094
rect 919 -3102 920 -3100
rect 926 -3096 927 -3094
rect 926 -3102 927 -3100
rect 933 -3096 934 -3094
rect 933 -3102 934 -3100
rect 940 -3096 941 -3094
rect 940 -3102 941 -3100
rect 947 -3096 948 -3094
rect 947 -3102 948 -3100
rect 954 -3096 955 -3094
rect 954 -3102 955 -3100
rect 961 -3096 962 -3094
rect 961 -3102 962 -3100
rect 968 -3096 969 -3094
rect 968 -3102 969 -3100
rect 975 -3096 976 -3094
rect 975 -3102 976 -3100
rect 982 -3096 983 -3094
rect 982 -3102 983 -3100
rect 989 -3096 990 -3094
rect 989 -3102 990 -3100
rect 996 -3096 997 -3094
rect 996 -3102 997 -3100
rect 1003 -3096 1004 -3094
rect 1003 -3102 1004 -3100
rect 1010 -3096 1011 -3094
rect 1010 -3102 1011 -3100
rect 1017 -3096 1018 -3094
rect 1017 -3102 1018 -3100
rect 1024 -3096 1025 -3094
rect 1024 -3102 1025 -3100
rect 1031 -3096 1032 -3094
rect 1031 -3102 1032 -3100
rect 1038 -3096 1039 -3094
rect 1038 -3102 1039 -3100
rect 1045 -3096 1046 -3094
rect 1045 -3102 1046 -3100
rect 1055 -3096 1056 -3094
rect 1055 -3102 1056 -3100
rect 1059 -3096 1060 -3094
rect 1059 -3102 1060 -3100
rect 1066 -3096 1067 -3094
rect 1066 -3102 1067 -3100
rect 1073 -3096 1074 -3094
rect 1076 -3096 1077 -3094
rect 1073 -3102 1074 -3100
rect 1076 -3102 1077 -3100
rect 1083 -3096 1084 -3094
rect 1080 -3102 1081 -3100
rect 1083 -3102 1084 -3100
rect 1087 -3096 1088 -3094
rect 1087 -3102 1088 -3100
rect 1094 -3096 1095 -3094
rect 1094 -3102 1095 -3100
rect 1101 -3096 1102 -3094
rect 1101 -3102 1102 -3100
rect 1108 -3096 1109 -3094
rect 1108 -3102 1109 -3100
rect 1115 -3096 1116 -3094
rect 1115 -3102 1116 -3100
rect 1122 -3096 1123 -3094
rect 1122 -3102 1123 -3100
rect 1125 -3102 1126 -3100
rect 1129 -3096 1130 -3094
rect 1129 -3102 1130 -3100
rect 1136 -3096 1137 -3094
rect 1136 -3102 1137 -3100
rect 1143 -3096 1144 -3094
rect 1143 -3102 1144 -3100
rect 1150 -3096 1151 -3094
rect 1150 -3102 1151 -3100
rect 1157 -3096 1158 -3094
rect 1160 -3096 1161 -3094
rect 1157 -3102 1158 -3100
rect 1160 -3102 1161 -3100
rect 1164 -3096 1165 -3094
rect 1164 -3102 1165 -3100
rect 1171 -3096 1172 -3094
rect 1171 -3102 1172 -3100
rect 1178 -3096 1179 -3094
rect 1178 -3102 1179 -3100
rect 1185 -3096 1186 -3094
rect 1185 -3102 1186 -3100
rect 1192 -3096 1193 -3094
rect 1192 -3102 1193 -3100
rect 1199 -3096 1200 -3094
rect 1199 -3102 1200 -3100
rect 1206 -3096 1207 -3094
rect 1206 -3102 1207 -3100
rect 1213 -3096 1214 -3094
rect 1216 -3096 1217 -3094
rect 1213 -3102 1214 -3100
rect 1216 -3102 1217 -3100
rect 1220 -3096 1221 -3094
rect 1220 -3102 1221 -3100
rect 1227 -3096 1228 -3094
rect 1227 -3102 1228 -3100
rect 1234 -3096 1235 -3094
rect 1237 -3096 1238 -3094
rect 1234 -3102 1235 -3100
rect 1237 -3102 1238 -3100
rect 1241 -3096 1242 -3094
rect 1241 -3102 1242 -3100
rect 1248 -3102 1249 -3100
rect 1255 -3096 1256 -3094
rect 1255 -3102 1256 -3100
rect 1262 -3096 1263 -3094
rect 1262 -3102 1263 -3100
rect 1269 -3096 1270 -3094
rect 1269 -3102 1270 -3100
rect 1276 -3102 1277 -3100
rect 1283 -3096 1284 -3094
rect 1283 -3102 1284 -3100
rect 1290 -3096 1291 -3094
rect 1290 -3102 1291 -3100
rect 1297 -3096 1298 -3094
rect 1297 -3102 1298 -3100
rect 1304 -3096 1305 -3094
rect 1304 -3102 1305 -3100
rect 1311 -3096 1312 -3094
rect 1311 -3102 1312 -3100
rect 1314 -3102 1315 -3100
rect 1318 -3096 1319 -3094
rect 1318 -3102 1319 -3100
rect 1325 -3096 1326 -3094
rect 1325 -3102 1326 -3100
rect 1332 -3096 1333 -3094
rect 1332 -3102 1333 -3100
rect 1339 -3096 1340 -3094
rect 1339 -3102 1340 -3100
rect 1346 -3096 1347 -3094
rect 1346 -3102 1347 -3100
rect 1353 -3096 1354 -3094
rect 1353 -3102 1354 -3100
rect 1360 -3096 1361 -3094
rect 1360 -3102 1361 -3100
rect 1367 -3096 1368 -3094
rect 1367 -3102 1368 -3100
rect 1374 -3096 1375 -3094
rect 1374 -3102 1375 -3100
rect 1381 -3096 1382 -3094
rect 1381 -3102 1382 -3100
rect 1388 -3096 1389 -3094
rect 1388 -3102 1389 -3100
rect 1398 -3096 1399 -3094
rect 1395 -3102 1396 -3100
rect 1398 -3102 1399 -3100
rect 1402 -3096 1403 -3094
rect 1405 -3096 1406 -3094
rect 1402 -3102 1403 -3100
rect 1409 -3096 1410 -3094
rect 1409 -3102 1410 -3100
rect 1416 -3096 1417 -3094
rect 1416 -3102 1417 -3100
rect 1423 -3096 1424 -3094
rect 1423 -3102 1424 -3100
rect 1430 -3096 1431 -3094
rect 1430 -3102 1431 -3100
rect 1437 -3096 1438 -3094
rect 1437 -3102 1438 -3100
rect 1444 -3102 1445 -3100
rect 1447 -3102 1448 -3100
rect 1451 -3096 1452 -3094
rect 1451 -3102 1452 -3100
rect 1458 -3096 1459 -3094
rect 1458 -3102 1459 -3100
rect 1465 -3096 1466 -3094
rect 1465 -3102 1466 -3100
rect 1472 -3096 1473 -3094
rect 1472 -3102 1473 -3100
rect 1479 -3096 1480 -3094
rect 1479 -3102 1480 -3100
rect 1486 -3096 1487 -3094
rect 1486 -3102 1487 -3100
rect 1493 -3096 1494 -3094
rect 1493 -3102 1494 -3100
rect 1500 -3096 1501 -3094
rect 1500 -3102 1501 -3100
rect 1507 -3096 1508 -3094
rect 1507 -3102 1508 -3100
rect 1514 -3096 1515 -3094
rect 1514 -3102 1515 -3100
rect 1521 -3096 1522 -3094
rect 1521 -3102 1522 -3100
rect 1528 -3096 1529 -3094
rect 1528 -3102 1529 -3100
rect 1535 -3096 1536 -3094
rect 1535 -3102 1536 -3100
rect 1542 -3096 1543 -3094
rect 1542 -3102 1543 -3100
rect 1549 -3096 1550 -3094
rect 1549 -3102 1550 -3100
rect 1556 -3096 1557 -3094
rect 1559 -3096 1560 -3094
rect 1556 -3102 1557 -3100
rect 1559 -3102 1560 -3100
rect 1566 -3096 1567 -3094
rect 1563 -3102 1564 -3100
rect 1566 -3102 1567 -3100
rect 1570 -3096 1571 -3094
rect 1570 -3102 1571 -3100
rect 1577 -3096 1578 -3094
rect 1577 -3102 1578 -3100
rect 1584 -3096 1585 -3094
rect 1584 -3102 1585 -3100
rect 1591 -3096 1592 -3094
rect 1591 -3102 1592 -3100
rect 1598 -3096 1599 -3094
rect 1598 -3102 1599 -3100
rect 1605 -3096 1606 -3094
rect 1605 -3102 1606 -3100
rect 1612 -3096 1613 -3094
rect 1612 -3102 1613 -3100
rect 1619 -3096 1620 -3094
rect 1619 -3102 1620 -3100
rect 1626 -3096 1627 -3094
rect 1626 -3102 1627 -3100
rect 1633 -3096 1634 -3094
rect 1633 -3102 1634 -3100
rect 1640 -3096 1641 -3094
rect 1640 -3102 1641 -3100
rect 1647 -3096 1648 -3094
rect 1647 -3102 1648 -3100
rect 1654 -3096 1655 -3094
rect 1654 -3102 1655 -3100
rect 1661 -3096 1662 -3094
rect 1661 -3102 1662 -3100
rect 1668 -3096 1669 -3094
rect 1668 -3102 1669 -3100
rect 1675 -3096 1676 -3094
rect 1675 -3102 1676 -3100
rect 1682 -3096 1683 -3094
rect 1685 -3096 1686 -3094
rect 1685 -3102 1686 -3100
rect 1689 -3096 1690 -3094
rect 1689 -3102 1690 -3100
rect 1696 -3096 1697 -3094
rect 1696 -3102 1697 -3100
rect 1703 -3096 1704 -3094
rect 1703 -3102 1704 -3100
rect 1710 -3096 1711 -3094
rect 1710 -3102 1711 -3100
rect 1717 -3096 1718 -3094
rect 1717 -3102 1718 -3100
rect 1724 -3096 1725 -3094
rect 1724 -3102 1725 -3100
rect 1731 -3096 1732 -3094
rect 1731 -3102 1732 -3100
rect 1738 -3096 1739 -3094
rect 1738 -3102 1739 -3100
rect 1745 -3096 1746 -3094
rect 1745 -3102 1746 -3100
rect 1752 -3096 1753 -3094
rect 1752 -3102 1753 -3100
rect 1759 -3096 1760 -3094
rect 1759 -3102 1760 -3100
rect 1766 -3096 1767 -3094
rect 1766 -3102 1767 -3100
rect 1773 -3096 1774 -3094
rect 1773 -3102 1774 -3100
rect 1780 -3096 1781 -3094
rect 1780 -3102 1781 -3100
rect 1787 -3096 1788 -3094
rect 1787 -3102 1788 -3100
rect 1794 -3096 1795 -3094
rect 1794 -3102 1795 -3100
rect 1801 -3096 1802 -3094
rect 1801 -3102 1802 -3100
rect 1808 -3096 1809 -3094
rect 1808 -3102 1809 -3100
rect 1815 -3096 1816 -3094
rect 1815 -3102 1816 -3100
rect 1822 -3096 1823 -3094
rect 1822 -3102 1823 -3100
rect 1829 -3096 1830 -3094
rect 1829 -3102 1830 -3100
rect 1836 -3096 1837 -3094
rect 1836 -3102 1837 -3100
rect 1843 -3096 1844 -3094
rect 1843 -3102 1844 -3100
rect 1850 -3096 1851 -3094
rect 1850 -3102 1851 -3100
rect 1857 -3096 1858 -3094
rect 1857 -3102 1858 -3100
rect 1864 -3096 1865 -3094
rect 1864 -3102 1865 -3100
rect 1871 -3096 1872 -3094
rect 1874 -3096 1875 -3094
rect 1871 -3102 1872 -3100
rect 1881 -3096 1882 -3094
rect 1878 -3102 1879 -3100
rect 1881 -3102 1882 -3100
rect 1885 -3096 1886 -3094
rect 1885 -3102 1886 -3100
rect 1892 -3096 1893 -3094
rect 1892 -3102 1893 -3100
rect 1899 -3096 1900 -3094
rect 1899 -3102 1900 -3100
rect 1906 -3096 1907 -3094
rect 1906 -3102 1907 -3100
rect 1913 -3096 1914 -3094
rect 1913 -3102 1914 -3100
rect 1920 -3096 1921 -3094
rect 1920 -3102 1921 -3100
rect 1927 -3096 1928 -3094
rect 1927 -3102 1928 -3100
rect 1934 -3096 1935 -3094
rect 1934 -3102 1935 -3100
rect 1941 -3096 1942 -3094
rect 1941 -3102 1942 -3100
rect 1948 -3096 1949 -3094
rect 1948 -3102 1949 -3100
rect 1955 -3096 1956 -3094
rect 1955 -3102 1956 -3100
rect 1962 -3096 1963 -3094
rect 1965 -3096 1966 -3094
rect 1962 -3102 1963 -3100
rect 1965 -3102 1966 -3100
rect 1969 -3096 1970 -3094
rect 1969 -3102 1970 -3100
rect 1976 -3096 1977 -3094
rect 1976 -3102 1977 -3100
rect 1983 -3096 1984 -3094
rect 1983 -3102 1984 -3100
rect 1990 -3096 1991 -3094
rect 1990 -3102 1991 -3100
rect 1997 -3096 1998 -3094
rect 1997 -3102 1998 -3100
rect 2004 -3096 2005 -3094
rect 2004 -3102 2005 -3100
rect 2032 -3096 2033 -3094
rect 2032 -3102 2033 -3100
rect 2046 -3096 2047 -3094
rect 2046 -3102 2047 -3100
rect 2074 -3096 2075 -3094
rect 2074 -3102 2075 -3100
rect 93 -3227 94 -3225
rect 93 -3233 94 -3231
rect 100 -3227 101 -3225
rect 100 -3233 101 -3231
rect 107 -3227 108 -3225
rect 107 -3233 108 -3231
rect 114 -3227 115 -3225
rect 117 -3233 118 -3231
rect 121 -3227 122 -3225
rect 121 -3233 122 -3231
rect 128 -3227 129 -3225
rect 128 -3233 129 -3231
rect 135 -3227 136 -3225
rect 135 -3233 136 -3231
rect 142 -3227 143 -3225
rect 142 -3233 143 -3231
rect 149 -3227 150 -3225
rect 149 -3233 150 -3231
rect 156 -3227 157 -3225
rect 156 -3233 157 -3231
rect 163 -3227 164 -3225
rect 163 -3233 164 -3231
rect 170 -3227 171 -3225
rect 173 -3233 174 -3231
rect 177 -3227 178 -3225
rect 177 -3233 178 -3231
rect 187 -3227 188 -3225
rect 187 -3233 188 -3231
rect 191 -3227 192 -3225
rect 194 -3227 195 -3225
rect 191 -3233 192 -3231
rect 198 -3227 199 -3225
rect 198 -3233 199 -3231
rect 205 -3227 206 -3225
rect 208 -3227 209 -3225
rect 205 -3233 206 -3231
rect 208 -3233 209 -3231
rect 212 -3227 213 -3225
rect 212 -3233 213 -3231
rect 219 -3227 220 -3225
rect 219 -3233 220 -3231
rect 226 -3227 227 -3225
rect 226 -3233 227 -3231
rect 233 -3227 234 -3225
rect 233 -3233 234 -3231
rect 240 -3227 241 -3225
rect 240 -3233 241 -3231
rect 247 -3227 248 -3225
rect 247 -3233 248 -3231
rect 254 -3227 255 -3225
rect 254 -3233 255 -3231
rect 261 -3227 262 -3225
rect 261 -3233 262 -3231
rect 268 -3227 269 -3225
rect 268 -3233 269 -3231
rect 275 -3227 276 -3225
rect 275 -3233 276 -3231
rect 282 -3227 283 -3225
rect 282 -3233 283 -3231
rect 289 -3227 290 -3225
rect 289 -3233 290 -3231
rect 296 -3227 297 -3225
rect 296 -3233 297 -3231
rect 303 -3227 304 -3225
rect 303 -3233 304 -3231
rect 310 -3227 311 -3225
rect 310 -3233 311 -3231
rect 317 -3227 318 -3225
rect 317 -3233 318 -3231
rect 324 -3227 325 -3225
rect 324 -3233 325 -3231
rect 331 -3227 332 -3225
rect 331 -3233 332 -3231
rect 338 -3227 339 -3225
rect 338 -3233 339 -3231
rect 345 -3227 346 -3225
rect 345 -3233 346 -3231
rect 352 -3227 353 -3225
rect 352 -3233 353 -3231
rect 359 -3227 360 -3225
rect 359 -3233 360 -3231
rect 366 -3227 367 -3225
rect 366 -3233 367 -3231
rect 373 -3227 374 -3225
rect 373 -3233 374 -3231
rect 380 -3227 381 -3225
rect 380 -3233 381 -3231
rect 387 -3227 388 -3225
rect 387 -3233 388 -3231
rect 394 -3227 395 -3225
rect 394 -3233 395 -3231
rect 401 -3227 402 -3225
rect 404 -3227 405 -3225
rect 401 -3233 402 -3231
rect 404 -3233 405 -3231
rect 408 -3227 409 -3225
rect 408 -3233 409 -3231
rect 415 -3227 416 -3225
rect 418 -3227 419 -3225
rect 415 -3233 416 -3231
rect 418 -3233 419 -3231
rect 425 -3227 426 -3225
rect 422 -3233 423 -3231
rect 429 -3227 430 -3225
rect 429 -3233 430 -3231
rect 436 -3227 437 -3225
rect 436 -3233 437 -3231
rect 443 -3227 444 -3225
rect 443 -3233 444 -3231
rect 450 -3227 451 -3225
rect 450 -3233 451 -3231
rect 457 -3227 458 -3225
rect 457 -3233 458 -3231
rect 464 -3227 465 -3225
rect 464 -3233 465 -3231
rect 471 -3227 472 -3225
rect 471 -3233 472 -3231
rect 478 -3227 479 -3225
rect 478 -3233 479 -3231
rect 485 -3227 486 -3225
rect 485 -3233 486 -3231
rect 492 -3227 493 -3225
rect 495 -3233 496 -3231
rect 499 -3227 500 -3225
rect 499 -3233 500 -3231
rect 506 -3227 507 -3225
rect 506 -3233 507 -3231
rect 513 -3227 514 -3225
rect 513 -3233 514 -3231
rect 520 -3227 521 -3225
rect 520 -3233 521 -3231
rect 527 -3227 528 -3225
rect 527 -3233 528 -3231
rect 534 -3227 535 -3225
rect 534 -3233 535 -3231
rect 541 -3227 542 -3225
rect 541 -3233 542 -3231
rect 548 -3227 549 -3225
rect 548 -3233 549 -3231
rect 555 -3227 556 -3225
rect 555 -3233 556 -3231
rect 562 -3227 563 -3225
rect 562 -3233 563 -3231
rect 569 -3227 570 -3225
rect 569 -3233 570 -3231
rect 576 -3227 577 -3225
rect 579 -3227 580 -3225
rect 576 -3233 577 -3231
rect 579 -3233 580 -3231
rect 583 -3227 584 -3225
rect 583 -3233 584 -3231
rect 590 -3227 591 -3225
rect 590 -3233 591 -3231
rect 597 -3227 598 -3225
rect 597 -3233 598 -3231
rect 604 -3227 605 -3225
rect 604 -3233 605 -3231
rect 611 -3227 612 -3225
rect 614 -3227 615 -3225
rect 611 -3233 612 -3231
rect 614 -3233 615 -3231
rect 618 -3227 619 -3225
rect 618 -3233 619 -3231
rect 625 -3227 626 -3225
rect 625 -3233 626 -3231
rect 632 -3227 633 -3225
rect 632 -3233 633 -3231
rect 639 -3227 640 -3225
rect 639 -3233 640 -3231
rect 646 -3227 647 -3225
rect 646 -3233 647 -3231
rect 653 -3227 654 -3225
rect 653 -3233 654 -3231
rect 660 -3227 661 -3225
rect 660 -3233 661 -3231
rect 667 -3227 668 -3225
rect 667 -3233 668 -3231
rect 674 -3227 675 -3225
rect 677 -3233 678 -3231
rect 681 -3227 682 -3225
rect 681 -3233 682 -3231
rect 688 -3227 689 -3225
rect 688 -3233 689 -3231
rect 695 -3227 696 -3225
rect 695 -3233 696 -3231
rect 702 -3227 703 -3225
rect 702 -3233 703 -3231
rect 709 -3227 710 -3225
rect 709 -3233 710 -3231
rect 716 -3227 717 -3225
rect 716 -3233 717 -3231
rect 719 -3233 720 -3231
rect 723 -3227 724 -3225
rect 723 -3233 724 -3231
rect 730 -3227 731 -3225
rect 730 -3233 731 -3231
rect 737 -3227 738 -3225
rect 737 -3233 738 -3231
rect 744 -3227 745 -3225
rect 747 -3227 748 -3225
rect 751 -3227 752 -3225
rect 751 -3233 752 -3231
rect 758 -3227 759 -3225
rect 758 -3233 759 -3231
rect 765 -3227 766 -3225
rect 768 -3227 769 -3225
rect 765 -3233 766 -3231
rect 768 -3233 769 -3231
rect 772 -3227 773 -3225
rect 772 -3233 773 -3231
rect 779 -3227 780 -3225
rect 779 -3233 780 -3231
rect 786 -3227 787 -3225
rect 786 -3233 787 -3231
rect 793 -3227 794 -3225
rect 793 -3233 794 -3231
rect 800 -3227 801 -3225
rect 800 -3233 801 -3231
rect 803 -3233 804 -3231
rect 807 -3227 808 -3225
rect 807 -3233 808 -3231
rect 814 -3227 815 -3225
rect 817 -3227 818 -3225
rect 817 -3233 818 -3231
rect 821 -3227 822 -3225
rect 821 -3233 822 -3231
rect 828 -3227 829 -3225
rect 828 -3233 829 -3231
rect 835 -3227 836 -3225
rect 835 -3233 836 -3231
rect 842 -3227 843 -3225
rect 842 -3233 843 -3231
rect 849 -3227 850 -3225
rect 849 -3233 850 -3231
rect 856 -3227 857 -3225
rect 856 -3233 857 -3231
rect 863 -3227 864 -3225
rect 863 -3233 864 -3231
rect 873 -3227 874 -3225
rect 870 -3233 871 -3231
rect 873 -3233 874 -3231
rect 877 -3227 878 -3225
rect 877 -3233 878 -3231
rect 884 -3227 885 -3225
rect 884 -3233 885 -3231
rect 891 -3227 892 -3225
rect 891 -3233 892 -3231
rect 898 -3227 899 -3225
rect 898 -3233 899 -3231
rect 905 -3227 906 -3225
rect 905 -3233 906 -3231
rect 912 -3227 913 -3225
rect 912 -3233 913 -3231
rect 919 -3227 920 -3225
rect 919 -3233 920 -3231
rect 926 -3227 927 -3225
rect 926 -3233 927 -3231
rect 933 -3227 934 -3225
rect 933 -3233 934 -3231
rect 940 -3227 941 -3225
rect 943 -3227 944 -3225
rect 940 -3233 941 -3231
rect 943 -3233 944 -3231
rect 947 -3227 948 -3225
rect 947 -3233 948 -3231
rect 954 -3227 955 -3225
rect 954 -3233 955 -3231
rect 957 -3233 958 -3231
rect 961 -3227 962 -3225
rect 961 -3233 962 -3231
rect 968 -3227 969 -3225
rect 968 -3233 969 -3231
rect 975 -3227 976 -3225
rect 975 -3233 976 -3231
rect 985 -3227 986 -3225
rect 985 -3233 986 -3231
rect 989 -3227 990 -3225
rect 989 -3233 990 -3231
rect 996 -3227 997 -3225
rect 996 -3233 997 -3231
rect 1003 -3227 1004 -3225
rect 1003 -3233 1004 -3231
rect 1010 -3227 1011 -3225
rect 1010 -3233 1011 -3231
rect 1017 -3227 1018 -3225
rect 1017 -3233 1018 -3231
rect 1024 -3227 1025 -3225
rect 1024 -3233 1025 -3231
rect 1031 -3227 1032 -3225
rect 1031 -3233 1032 -3231
rect 1038 -3227 1039 -3225
rect 1038 -3233 1039 -3231
rect 1045 -3227 1046 -3225
rect 1045 -3233 1046 -3231
rect 1052 -3227 1053 -3225
rect 1052 -3233 1053 -3231
rect 1059 -3227 1060 -3225
rect 1059 -3233 1060 -3231
rect 1066 -3227 1067 -3225
rect 1066 -3233 1067 -3231
rect 1073 -3227 1074 -3225
rect 1073 -3233 1074 -3231
rect 1080 -3227 1081 -3225
rect 1080 -3233 1081 -3231
rect 1087 -3227 1088 -3225
rect 1087 -3233 1088 -3231
rect 1094 -3227 1095 -3225
rect 1094 -3233 1095 -3231
rect 1101 -3227 1102 -3225
rect 1101 -3233 1102 -3231
rect 1108 -3227 1109 -3225
rect 1111 -3227 1112 -3225
rect 1108 -3233 1109 -3231
rect 1115 -3227 1116 -3225
rect 1115 -3233 1116 -3231
rect 1122 -3227 1123 -3225
rect 1122 -3233 1123 -3231
rect 1129 -3227 1130 -3225
rect 1129 -3233 1130 -3231
rect 1136 -3227 1137 -3225
rect 1136 -3233 1137 -3231
rect 1143 -3227 1144 -3225
rect 1143 -3233 1144 -3231
rect 1150 -3227 1151 -3225
rect 1150 -3233 1151 -3231
rect 1157 -3227 1158 -3225
rect 1157 -3233 1158 -3231
rect 1164 -3227 1165 -3225
rect 1167 -3227 1168 -3225
rect 1164 -3233 1165 -3231
rect 1167 -3233 1168 -3231
rect 1171 -3227 1172 -3225
rect 1171 -3233 1172 -3231
rect 1178 -3227 1179 -3225
rect 1178 -3233 1179 -3231
rect 1185 -3227 1186 -3225
rect 1185 -3233 1186 -3231
rect 1192 -3227 1193 -3225
rect 1192 -3233 1193 -3231
rect 1199 -3227 1200 -3225
rect 1199 -3233 1200 -3231
rect 1206 -3227 1207 -3225
rect 1206 -3233 1207 -3231
rect 1213 -3227 1214 -3225
rect 1216 -3227 1217 -3225
rect 1213 -3233 1214 -3231
rect 1216 -3233 1217 -3231
rect 1220 -3227 1221 -3225
rect 1220 -3233 1221 -3231
rect 1227 -3227 1228 -3225
rect 1227 -3233 1228 -3231
rect 1234 -3233 1235 -3231
rect 1237 -3233 1238 -3231
rect 1241 -3227 1242 -3225
rect 1241 -3233 1242 -3231
rect 1248 -3227 1249 -3225
rect 1248 -3233 1249 -3231
rect 1255 -3227 1256 -3225
rect 1258 -3227 1259 -3225
rect 1255 -3233 1256 -3231
rect 1262 -3227 1263 -3225
rect 1262 -3233 1263 -3231
rect 1269 -3227 1270 -3225
rect 1269 -3233 1270 -3231
rect 1276 -3227 1277 -3225
rect 1276 -3233 1277 -3231
rect 1283 -3227 1284 -3225
rect 1283 -3233 1284 -3231
rect 1290 -3227 1291 -3225
rect 1290 -3233 1291 -3231
rect 1297 -3227 1298 -3225
rect 1297 -3233 1298 -3231
rect 1304 -3227 1305 -3225
rect 1304 -3233 1305 -3231
rect 1311 -3227 1312 -3225
rect 1311 -3233 1312 -3231
rect 1318 -3227 1319 -3225
rect 1318 -3233 1319 -3231
rect 1325 -3227 1326 -3225
rect 1325 -3233 1326 -3231
rect 1332 -3227 1333 -3225
rect 1332 -3233 1333 -3231
rect 1339 -3227 1340 -3225
rect 1339 -3233 1340 -3231
rect 1346 -3227 1347 -3225
rect 1346 -3233 1347 -3231
rect 1353 -3227 1354 -3225
rect 1356 -3227 1357 -3225
rect 1353 -3233 1354 -3231
rect 1360 -3227 1361 -3225
rect 1360 -3233 1361 -3231
rect 1367 -3227 1368 -3225
rect 1367 -3233 1368 -3231
rect 1374 -3227 1375 -3225
rect 1374 -3233 1375 -3231
rect 1381 -3227 1382 -3225
rect 1381 -3233 1382 -3231
rect 1388 -3227 1389 -3225
rect 1388 -3233 1389 -3231
rect 1395 -3227 1396 -3225
rect 1395 -3233 1396 -3231
rect 1402 -3227 1403 -3225
rect 1402 -3233 1403 -3231
rect 1409 -3227 1410 -3225
rect 1409 -3233 1410 -3231
rect 1416 -3227 1417 -3225
rect 1416 -3233 1417 -3231
rect 1423 -3227 1424 -3225
rect 1423 -3233 1424 -3231
rect 1430 -3227 1431 -3225
rect 1430 -3233 1431 -3231
rect 1437 -3227 1438 -3225
rect 1437 -3233 1438 -3231
rect 1444 -3227 1445 -3225
rect 1444 -3233 1445 -3231
rect 1451 -3227 1452 -3225
rect 1451 -3233 1452 -3231
rect 1458 -3227 1459 -3225
rect 1461 -3227 1462 -3225
rect 1458 -3233 1459 -3231
rect 1465 -3227 1466 -3225
rect 1465 -3233 1466 -3231
rect 1472 -3227 1473 -3225
rect 1472 -3233 1473 -3231
rect 1479 -3227 1480 -3225
rect 1479 -3233 1480 -3231
rect 1486 -3227 1487 -3225
rect 1486 -3233 1487 -3231
rect 1493 -3227 1494 -3225
rect 1493 -3233 1494 -3231
rect 1500 -3227 1501 -3225
rect 1500 -3233 1501 -3231
rect 1507 -3227 1508 -3225
rect 1507 -3233 1508 -3231
rect 1514 -3227 1515 -3225
rect 1514 -3233 1515 -3231
rect 1521 -3227 1522 -3225
rect 1521 -3233 1522 -3231
rect 1528 -3227 1529 -3225
rect 1528 -3233 1529 -3231
rect 1535 -3227 1536 -3225
rect 1535 -3233 1536 -3231
rect 1542 -3227 1543 -3225
rect 1542 -3233 1543 -3231
rect 1549 -3227 1550 -3225
rect 1549 -3233 1550 -3231
rect 1556 -3227 1557 -3225
rect 1556 -3233 1557 -3231
rect 1563 -3227 1564 -3225
rect 1563 -3233 1564 -3231
rect 1570 -3227 1571 -3225
rect 1570 -3233 1571 -3231
rect 1577 -3227 1578 -3225
rect 1580 -3233 1581 -3231
rect 1584 -3227 1585 -3225
rect 1584 -3233 1585 -3231
rect 1591 -3227 1592 -3225
rect 1591 -3233 1592 -3231
rect 1598 -3227 1599 -3225
rect 1598 -3233 1599 -3231
rect 1605 -3227 1606 -3225
rect 1605 -3233 1606 -3231
rect 1612 -3227 1613 -3225
rect 1612 -3233 1613 -3231
rect 1619 -3227 1620 -3225
rect 1619 -3233 1620 -3231
rect 1626 -3227 1627 -3225
rect 1626 -3233 1627 -3231
rect 1633 -3227 1634 -3225
rect 1633 -3233 1634 -3231
rect 1640 -3227 1641 -3225
rect 1643 -3227 1644 -3225
rect 1640 -3233 1641 -3231
rect 1643 -3233 1644 -3231
rect 1647 -3227 1648 -3225
rect 1650 -3227 1651 -3225
rect 1647 -3233 1648 -3231
rect 1650 -3233 1651 -3231
rect 1654 -3227 1655 -3225
rect 1657 -3227 1658 -3225
rect 1654 -3233 1655 -3231
rect 1661 -3227 1662 -3225
rect 1661 -3233 1662 -3231
rect 1671 -3227 1672 -3225
rect 1671 -3233 1672 -3231
rect 1675 -3227 1676 -3225
rect 1675 -3233 1676 -3231
rect 1682 -3227 1683 -3225
rect 1685 -3227 1686 -3225
rect 1682 -3233 1683 -3231
rect 1685 -3233 1686 -3231
rect 1689 -3227 1690 -3225
rect 1689 -3233 1690 -3231
rect 1696 -3227 1697 -3225
rect 1696 -3233 1697 -3231
rect 1703 -3227 1704 -3225
rect 1703 -3233 1704 -3231
rect 1710 -3227 1711 -3225
rect 1710 -3233 1711 -3231
rect 1717 -3227 1718 -3225
rect 1717 -3233 1718 -3231
rect 1724 -3227 1725 -3225
rect 1724 -3233 1725 -3231
rect 1731 -3227 1732 -3225
rect 1731 -3233 1732 -3231
rect 1738 -3227 1739 -3225
rect 1738 -3233 1739 -3231
rect 1745 -3227 1746 -3225
rect 1745 -3233 1746 -3231
rect 1752 -3227 1753 -3225
rect 1752 -3233 1753 -3231
rect 1759 -3227 1760 -3225
rect 1759 -3233 1760 -3231
rect 1766 -3227 1767 -3225
rect 1766 -3233 1767 -3231
rect 1773 -3227 1774 -3225
rect 1773 -3233 1774 -3231
rect 1780 -3227 1781 -3225
rect 1780 -3233 1781 -3231
rect 1808 -3227 1809 -3225
rect 1808 -3233 1809 -3231
rect 1815 -3227 1816 -3225
rect 1815 -3233 1816 -3231
rect 1822 -3227 1823 -3225
rect 1822 -3233 1823 -3231
rect 1850 -3227 1851 -3225
rect 1853 -3227 1854 -3225
rect 1850 -3233 1851 -3231
rect 1853 -3233 1854 -3231
rect 1857 -3227 1858 -3225
rect 1857 -3233 1858 -3231
rect 1864 -3227 1865 -3225
rect 1864 -3233 1865 -3231
rect 1878 -3227 1879 -3225
rect 1878 -3233 1879 -3231
rect 1885 -3227 1886 -3225
rect 1885 -3233 1886 -3231
rect 1892 -3227 1893 -3225
rect 1892 -3233 1893 -3231
rect 1906 -3227 1907 -3225
rect 1906 -3233 1907 -3231
rect 1920 -3227 1921 -3225
rect 1920 -3233 1921 -3231
rect 1962 -3227 1963 -3225
rect 1965 -3227 1966 -3225
rect 1962 -3233 1963 -3231
rect 1965 -3233 1966 -3231
rect 1969 -3227 1970 -3225
rect 1969 -3233 1970 -3231
rect 1976 -3227 1977 -3225
rect 1976 -3233 1977 -3231
rect 1983 -3227 1984 -3225
rect 1983 -3233 1984 -3231
rect 2018 -3227 2019 -3225
rect 2018 -3233 2019 -3231
rect 2046 -3227 2047 -3225
rect 2046 -3233 2047 -3231
rect 142 -3330 143 -3328
rect 142 -3336 143 -3334
rect 163 -3330 164 -3328
rect 163 -3336 164 -3334
rect 170 -3330 171 -3328
rect 170 -3336 171 -3334
rect 177 -3330 178 -3328
rect 177 -3336 178 -3334
rect 184 -3330 185 -3328
rect 184 -3336 185 -3334
rect 191 -3330 192 -3328
rect 191 -3336 192 -3334
rect 198 -3330 199 -3328
rect 198 -3336 199 -3334
rect 205 -3330 206 -3328
rect 205 -3336 206 -3334
rect 215 -3330 216 -3328
rect 212 -3336 213 -3334
rect 215 -3336 216 -3334
rect 219 -3330 220 -3328
rect 219 -3336 220 -3334
rect 226 -3330 227 -3328
rect 229 -3330 230 -3328
rect 236 -3336 237 -3334
rect 240 -3330 241 -3328
rect 240 -3336 241 -3334
rect 247 -3330 248 -3328
rect 247 -3336 248 -3334
rect 254 -3330 255 -3328
rect 257 -3330 258 -3328
rect 257 -3336 258 -3334
rect 261 -3330 262 -3328
rect 261 -3336 262 -3334
rect 268 -3330 269 -3328
rect 268 -3336 269 -3334
rect 275 -3330 276 -3328
rect 275 -3336 276 -3334
rect 282 -3330 283 -3328
rect 282 -3336 283 -3334
rect 289 -3330 290 -3328
rect 289 -3336 290 -3334
rect 296 -3330 297 -3328
rect 296 -3336 297 -3334
rect 303 -3330 304 -3328
rect 303 -3336 304 -3334
rect 310 -3330 311 -3328
rect 310 -3336 311 -3334
rect 317 -3330 318 -3328
rect 317 -3336 318 -3334
rect 324 -3330 325 -3328
rect 324 -3336 325 -3334
rect 331 -3330 332 -3328
rect 331 -3336 332 -3334
rect 338 -3330 339 -3328
rect 338 -3336 339 -3334
rect 345 -3330 346 -3328
rect 345 -3336 346 -3334
rect 352 -3330 353 -3328
rect 352 -3336 353 -3334
rect 359 -3330 360 -3328
rect 359 -3336 360 -3334
rect 366 -3330 367 -3328
rect 366 -3336 367 -3334
rect 373 -3330 374 -3328
rect 373 -3336 374 -3334
rect 380 -3330 381 -3328
rect 383 -3330 384 -3328
rect 380 -3336 381 -3334
rect 383 -3336 384 -3334
rect 387 -3330 388 -3328
rect 387 -3336 388 -3334
rect 394 -3330 395 -3328
rect 394 -3336 395 -3334
rect 401 -3330 402 -3328
rect 401 -3336 402 -3334
rect 408 -3330 409 -3328
rect 408 -3336 409 -3334
rect 415 -3330 416 -3328
rect 415 -3336 416 -3334
rect 418 -3336 419 -3334
rect 422 -3330 423 -3328
rect 422 -3336 423 -3334
rect 429 -3330 430 -3328
rect 429 -3336 430 -3334
rect 436 -3330 437 -3328
rect 436 -3336 437 -3334
rect 443 -3330 444 -3328
rect 443 -3336 444 -3334
rect 450 -3330 451 -3328
rect 450 -3336 451 -3334
rect 457 -3330 458 -3328
rect 457 -3336 458 -3334
rect 464 -3330 465 -3328
rect 464 -3336 465 -3334
rect 471 -3330 472 -3328
rect 471 -3336 472 -3334
rect 478 -3330 479 -3328
rect 478 -3336 479 -3334
rect 485 -3330 486 -3328
rect 485 -3336 486 -3334
rect 492 -3330 493 -3328
rect 492 -3336 493 -3334
rect 499 -3330 500 -3328
rect 499 -3336 500 -3334
rect 506 -3330 507 -3328
rect 506 -3336 507 -3334
rect 513 -3330 514 -3328
rect 513 -3336 514 -3334
rect 520 -3330 521 -3328
rect 520 -3336 521 -3334
rect 527 -3330 528 -3328
rect 527 -3336 528 -3334
rect 534 -3330 535 -3328
rect 537 -3330 538 -3328
rect 534 -3336 535 -3334
rect 537 -3336 538 -3334
rect 541 -3330 542 -3328
rect 541 -3336 542 -3334
rect 548 -3330 549 -3328
rect 548 -3336 549 -3334
rect 555 -3330 556 -3328
rect 555 -3336 556 -3334
rect 562 -3330 563 -3328
rect 562 -3336 563 -3334
rect 569 -3330 570 -3328
rect 569 -3336 570 -3334
rect 576 -3330 577 -3328
rect 583 -3330 584 -3328
rect 583 -3336 584 -3334
rect 590 -3330 591 -3328
rect 590 -3336 591 -3334
rect 597 -3330 598 -3328
rect 600 -3330 601 -3328
rect 597 -3336 598 -3334
rect 600 -3336 601 -3334
rect 604 -3330 605 -3328
rect 604 -3336 605 -3334
rect 611 -3330 612 -3328
rect 611 -3336 612 -3334
rect 618 -3330 619 -3328
rect 618 -3336 619 -3334
rect 625 -3330 626 -3328
rect 625 -3336 626 -3334
rect 632 -3330 633 -3328
rect 632 -3336 633 -3334
rect 639 -3330 640 -3328
rect 642 -3330 643 -3328
rect 646 -3330 647 -3328
rect 646 -3336 647 -3334
rect 653 -3330 654 -3328
rect 653 -3336 654 -3334
rect 660 -3330 661 -3328
rect 660 -3336 661 -3334
rect 667 -3330 668 -3328
rect 667 -3336 668 -3334
rect 674 -3330 675 -3328
rect 674 -3336 675 -3334
rect 681 -3330 682 -3328
rect 681 -3336 682 -3334
rect 688 -3330 689 -3328
rect 688 -3336 689 -3334
rect 695 -3330 696 -3328
rect 695 -3336 696 -3334
rect 702 -3330 703 -3328
rect 702 -3336 703 -3334
rect 709 -3330 710 -3328
rect 709 -3336 710 -3334
rect 716 -3330 717 -3328
rect 716 -3336 717 -3334
rect 726 -3330 727 -3328
rect 723 -3336 724 -3334
rect 733 -3330 734 -3328
rect 730 -3336 731 -3334
rect 737 -3330 738 -3328
rect 737 -3336 738 -3334
rect 744 -3330 745 -3328
rect 744 -3336 745 -3334
rect 751 -3330 752 -3328
rect 751 -3336 752 -3334
rect 758 -3330 759 -3328
rect 758 -3336 759 -3334
rect 765 -3330 766 -3328
rect 765 -3336 766 -3334
rect 772 -3330 773 -3328
rect 772 -3336 773 -3334
rect 779 -3330 780 -3328
rect 782 -3330 783 -3328
rect 779 -3336 780 -3334
rect 786 -3330 787 -3328
rect 786 -3336 787 -3334
rect 793 -3330 794 -3328
rect 793 -3336 794 -3334
rect 800 -3330 801 -3328
rect 800 -3336 801 -3334
rect 807 -3330 808 -3328
rect 807 -3336 808 -3334
rect 814 -3330 815 -3328
rect 814 -3336 815 -3334
rect 821 -3330 822 -3328
rect 821 -3336 822 -3334
rect 828 -3330 829 -3328
rect 828 -3336 829 -3334
rect 835 -3330 836 -3328
rect 835 -3336 836 -3334
rect 842 -3330 843 -3328
rect 842 -3336 843 -3334
rect 849 -3330 850 -3328
rect 849 -3336 850 -3334
rect 852 -3336 853 -3334
rect 856 -3330 857 -3328
rect 856 -3336 857 -3334
rect 863 -3330 864 -3328
rect 863 -3336 864 -3334
rect 870 -3330 871 -3328
rect 870 -3336 871 -3334
rect 877 -3330 878 -3328
rect 877 -3336 878 -3334
rect 884 -3330 885 -3328
rect 884 -3336 885 -3334
rect 891 -3330 892 -3328
rect 891 -3336 892 -3334
rect 898 -3330 899 -3328
rect 898 -3336 899 -3334
rect 905 -3330 906 -3328
rect 905 -3336 906 -3334
rect 912 -3330 913 -3328
rect 912 -3336 913 -3334
rect 919 -3330 920 -3328
rect 919 -3336 920 -3334
rect 926 -3330 927 -3328
rect 929 -3330 930 -3328
rect 926 -3336 927 -3334
rect 933 -3330 934 -3328
rect 933 -3336 934 -3334
rect 940 -3330 941 -3328
rect 940 -3336 941 -3334
rect 947 -3330 948 -3328
rect 947 -3336 948 -3334
rect 957 -3330 958 -3328
rect 954 -3336 955 -3334
rect 957 -3336 958 -3334
rect 961 -3330 962 -3328
rect 961 -3336 962 -3334
rect 968 -3330 969 -3328
rect 968 -3336 969 -3334
rect 971 -3336 972 -3334
rect 978 -3330 979 -3328
rect 975 -3336 976 -3334
rect 978 -3336 979 -3334
rect 982 -3330 983 -3328
rect 982 -3336 983 -3334
rect 989 -3330 990 -3328
rect 992 -3330 993 -3328
rect 989 -3336 990 -3334
rect 996 -3330 997 -3328
rect 996 -3336 997 -3334
rect 1003 -3330 1004 -3328
rect 1003 -3336 1004 -3334
rect 1010 -3330 1011 -3328
rect 1010 -3336 1011 -3334
rect 1017 -3330 1018 -3328
rect 1017 -3336 1018 -3334
rect 1024 -3330 1025 -3328
rect 1024 -3336 1025 -3334
rect 1031 -3330 1032 -3328
rect 1031 -3336 1032 -3334
rect 1038 -3330 1039 -3328
rect 1038 -3336 1039 -3334
rect 1045 -3330 1046 -3328
rect 1045 -3336 1046 -3334
rect 1052 -3330 1053 -3328
rect 1052 -3336 1053 -3334
rect 1059 -3330 1060 -3328
rect 1059 -3336 1060 -3334
rect 1066 -3330 1067 -3328
rect 1069 -3330 1070 -3328
rect 1066 -3336 1067 -3334
rect 1073 -3330 1074 -3328
rect 1073 -3336 1074 -3334
rect 1080 -3330 1081 -3328
rect 1080 -3336 1081 -3334
rect 1083 -3336 1084 -3334
rect 1087 -3330 1088 -3328
rect 1087 -3336 1088 -3334
rect 1094 -3330 1095 -3328
rect 1094 -3336 1095 -3334
rect 1097 -3336 1098 -3334
rect 1104 -3330 1105 -3328
rect 1104 -3336 1105 -3334
rect 1108 -3330 1109 -3328
rect 1108 -3336 1109 -3334
rect 1115 -3330 1116 -3328
rect 1115 -3336 1116 -3334
rect 1122 -3330 1123 -3328
rect 1122 -3336 1123 -3334
rect 1129 -3330 1130 -3328
rect 1129 -3336 1130 -3334
rect 1136 -3330 1137 -3328
rect 1136 -3336 1137 -3334
rect 1143 -3330 1144 -3328
rect 1143 -3336 1144 -3334
rect 1150 -3330 1151 -3328
rect 1150 -3336 1151 -3334
rect 1157 -3330 1158 -3328
rect 1157 -3336 1158 -3334
rect 1164 -3330 1165 -3328
rect 1164 -3336 1165 -3334
rect 1171 -3330 1172 -3328
rect 1171 -3336 1172 -3334
rect 1178 -3330 1179 -3328
rect 1178 -3336 1179 -3334
rect 1185 -3330 1186 -3328
rect 1185 -3336 1186 -3334
rect 1192 -3330 1193 -3328
rect 1192 -3336 1193 -3334
rect 1199 -3330 1200 -3328
rect 1199 -3336 1200 -3334
rect 1206 -3330 1207 -3328
rect 1206 -3336 1207 -3334
rect 1216 -3330 1217 -3328
rect 1213 -3336 1214 -3334
rect 1216 -3336 1217 -3334
rect 1220 -3330 1221 -3328
rect 1220 -3336 1221 -3334
rect 1227 -3330 1228 -3328
rect 1227 -3336 1228 -3334
rect 1234 -3330 1235 -3328
rect 1237 -3330 1238 -3328
rect 1234 -3336 1235 -3334
rect 1237 -3336 1238 -3334
rect 1241 -3330 1242 -3328
rect 1241 -3336 1242 -3334
rect 1248 -3330 1249 -3328
rect 1248 -3336 1249 -3334
rect 1255 -3330 1256 -3328
rect 1255 -3336 1256 -3334
rect 1262 -3330 1263 -3328
rect 1262 -3336 1263 -3334
rect 1269 -3330 1270 -3328
rect 1269 -3336 1270 -3334
rect 1272 -3336 1273 -3334
rect 1276 -3330 1277 -3328
rect 1276 -3336 1277 -3334
rect 1283 -3330 1284 -3328
rect 1283 -3336 1284 -3334
rect 1290 -3330 1291 -3328
rect 1290 -3336 1291 -3334
rect 1297 -3330 1298 -3328
rect 1297 -3336 1298 -3334
rect 1304 -3330 1305 -3328
rect 1304 -3336 1305 -3334
rect 1311 -3330 1312 -3328
rect 1311 -3336 1312 -3334
rect 1318 -3330 1319 -3328
rect 1318 -3336 1319 -3334
rect 1325 -3330 1326 -3328
rect 1325 -3336 1326 -3334
rect 1332 -3330 1333 -3328
rect 1332 -3336 1333 -3334
rect 1339 -3330 1340 -3328
rect 1339 -3336 1340 -3334
rect 1346 -3330 1347 -3328
rect 1346 -3336 1347 -3334
rect 1353 -3330 1354 -3328
rect 1353 -3336 1354 -3334
rect 1360 -3330 1361 -3328
rect 1360 -3336 1361 -3334
rect 1367 -3330 1368 -3328
rect 1370 -3336 1371 -3334
rect 1374 -3330 1375 -3328
rect 1374 -3336 1375 -3334
rect 1381 -3336 1382 -3334
rect 1384 -3336 1385 -3334
rect 1388 -3330 1389 -3328
rect 1388 -3336 1389 -3334
rect 1395 -3330 1396 -3328
rect 1395 -3336 1396 -3334
rect 1402 -3330 1403 -3328
rect 1402 -3336 1403 -3334
rect 1409 -3330 1410 -3328
rect 1409 -3336 1410 -3334
rect 1416 -3336 1417 -3334
rect 1419 -3336 1420 -3334
rect 1423 -3330 1424 -3328
rect 1423 -3336 1424 -3334
rect 1430 -3330 1431 -3328
rect 1430 -3336 1431 -3334
rect 1437 -3330 1438 -3328
rect 1437 -3336 1438 -3334
rect 1444 -3330 1445 -3328
rect 1444 -3336 1445 -3334
rect 1451 -3330 1452 -3328
rect 1451 -3336 1452 -3334
rect 1458 -3330 1459 -3328
rect 1458 -3336 1459 -3334
rect 1465 -3330 1466 -3328
rect 1465 -3336 1466 -3334
rect 1472 -3330 1473 -3328
rect 1472 -3336 1473 -3334
rect 1479 -3330 1480 -3328
rect 1479 -3336 1480 -3334
rect 1486 -3330 1487 -3328
rect 1486 -3336 1487 -3334
rect 1493 -3330 1494 -3328
rect 1493 -3336 1494 -3334
rect 1500 -3330 1501 -3328
rect 1500 -3336 1501 -3334
rect 1507 -3330 1508 -3328
rect 1507 -3336 1508 -3334
rect 1514 -3330 1515 -3328
rect 1514 -3336 1515 -3334
rect 1521 -3330 1522 -3328
rect 1521 -3336 1522 -3334
rect 1528 -3330 1529 -3328
rect 1528 -3336 1529 -3334
rect 1556 -3330 1557 -3328
rect 1556 -3336 1557 -3334
rect 1563 -3330 1564 -3328
rect 1563 -3336 1564 -3334
rect 1591 -3330 1592 -3328
rect 1591 -3336 1592 -3334
rect 1598 -3330 1599 -3328
rect 1598 -3336 1599 -3334
rect 1605 -3330 1606 -3328
rect 1605 -3336 1606 -3334
rect 1608 -3336 1609 -3334
rect 1626 -3330 1627 -3328
rect 1626 -3336 1627 -3334
rect 1654 -3330 1655 -3328
rect 1654 -3336 1655 -3334
rect 1661 -3330 1662 -3328
rect 1661 -3336 1662 -3334
rect 1668 -3330 1669 -3328
rect 1668 -3336 1669 -3334
rect 1717 -3330 1718 -3328
rect 1717 -3336 1718 -3334
rect 1724 -3330 1725 -3328
rect 1727 -3330 1728 -3328
rect 1727 -3336 1728 -3334
rect 1731 -3330 1732 -3328
rect 1731 -3336 1732 -3334
rect 1738 -3330 1739 -3328
rect 1738 -3336 1739 -3334
rect 1745 -3330 1746 -3328
rect 1745 -3336 1746 -3334
rect 1752 -3330 1753 -3328
rect 1752 -3336 1753 -3334
rect 1766 -3330 1767 -3328
rect 1766 -3336 1767 -3334
rect 1780 -3330 1781 -3328
rect 1780 -3336 1781 -3334
rect 1787 -3330 1788 -3328
rect 1787 -3336 1788 -3334
rect 1794 -3330 1795 -3328
rect 1794 -3336 1795 -3334
rect 1801 -3330 1802 -3328
rect 1801 -3336 1802 -3334
rect 1815 -3330 1816 -3328
rect 1815 -3336 1816 -3334
rect 1836 -3330 1837 -3328
rect 1836 -3336 1837 -3334
rect 1843 -3330 1844 -3328
rect 1843 -3336 1844 -3334
rect 1850 -3330 1851 -3328
rect 1853 -3330 1854 -3328
rect 1850 -3336 1851 -3334
rect 1853 -3336 1854 -3334
rect 1857 -3330 1858 -3328
rect 1857 -3336 1858 -3334
rect 1864 -3330 1865 -3328
rect 1864 -3336 1865 -3334
rect 1871 -3330 1872 -3328
rect 1871 -3336 1872 -3334
rect 1878 -3330 1879 -3328
rect 1878 -3336 1879 -3334
rect 1885 -3336 1886 -3334
rect 1888 -3336 1889 -3334
rect 1892 -3330 1893 -3328
rect 1892 -3336 1893 -3334
rect 1906 -3330 1907 -3328
rect 1906 -3336 1907 -3334
rect 1962 -3330 1963 -3328
rect 1962 -3336 1963 -3334
rect 1969 -3330 1970 -3328
rect 1969 -3336 1970 -3334
rect 2025 -3330 2026 -3328
rect 2025 -3336 2026 -3334
rect 2028 -3336 2029 -3334
rect 2032 -3330 2033 -3328
rect 2032 -3336 2033 -3334
rect 173 -3417 174 -3415
rect 170 -3423 171 -3421
rect 173 -3423 174 -3421
rect 180 -3417 181 -3415
rect 296 -3417 297 -3415
rect 296 -3423 297 -3421
rect 310 -3417 311 -3415
rect 310 -3423 311 -3421
rect 317 -3423 318 -3421
rect 331 -3417 332 -3415
rect 331 -3423 332 -3421
rect 338 -3417 339 -3415
rect 338 -3423 339 -3421
rect 345 -3417 346 -3415
rect 345 -3423 346 -3421
rect 359 -3417 360 -3415
rect 359 -3423 360 -3421
rect 373 -3417 374 -3415
rect 373 -3423 374 -3421
rect 380 -3417 381 -3415
rect 380 -3423 381 -3421
rect 387 -3417 388 -3415
rect 390 -3417 391 -3415
rect 390 -3423 391 -3421
rect 394 -3417 395 -3415
rect 394 -3423 395 -3421
rect 401 -3417 402 -3415
rect 401 -3423 402 -3421
rect 404 -3423 405 -3421
rect 408 -3417 409 -3415
rect 408 -3423 409 -3421
rect 422 -3417 423 -3415
rect 422 -3423 423 -3421
rect 429 -3417 430 -3415
rect 429 -3423 430 -3421
rect 436 -3417 437 -3415
rect 436 -3423 437 -3421
rect 439 -3423 440 -3421
rect 443 -3417 444 -3415
rect 443 -3423 444 -3421
rect 450 -3417 451 -3415
rect 450 -3423 451 -3421
rect 457 -3417 458 -3415
rect 457 -3423 458 -3421
rect 464 -3417 465 -3415
rect 464 -3423 465 -3421
rect 474 -3417 475 -3415
rect 471 -3423 472 -3421
rect 474 -3423 475 -3421
rect 478 -3417 479 -3415
rect 478 -3423 479 -3421
rect 488 -3417 489 -3415
rect 488 -3423 489 -3421
rect 492 -3417 493 -3415
rect 492 -3423 493 -3421
rect 499 -3417 500 -3415
rect 499 -3423 500 -3421
rect 506 -3417 507 -3415
rect 506 -3423 507 -3421
rect 513 -3417 514 -3415
rect 513 -3423 514 -3421
rect 520 -3417 521 -3415
rect 520 -3423 521 -3421
rect 527 -3417 528 -3415
rect 527 -3423 528 -3421
rect 534 -3417 535 -3415
rect 534 -3423 535 -3421
rect 541 -3417 542 -3415
rect 541 -3423 542 -3421
rect 548 -3417 549 -3415
rect 548 -3423 549 -3421
rect 555 -3417 556 -3415
rect 555 -3423 556 -3421
rect 558 -3423 559 -3421
rect 562 -3417 563 -3415
rect 562 -3423 563 -3421
rect 569 -3417 570 -3415
rect 569 -3423 570 -3421
rect 576 -3423 577 -3421
rect 583 -3417 584 -3415
rect 583 -3423 584 -3421
rect 590 -3417 591 -3415
rect 590 -3423 591 -3421
rect 597 -3417 598 -3415
rect 597 -3423 598 -3421
rect 604 -3417 605 -3415
rect 604 -3423 605 -3421
rect 611 -3417 612 -3415
rect 611 -3423 612 -3421
rect 618 -3417 619 -3415
rect 618 -3423 619 -3421
rect 625 -3417 626 -3415
rect 625 -3423 626 -3421
rect 632 -3417 633 -3415
rect 632 -3423 633 -3421
rect 639 -3417 640 -3415
rect 639 -3423 640 -3421
rect 646 -3417 647 -3415
rect 646 -3423 647 -3421
rect 653 -3417 654 -3415
rect 653 -3423 654 -3421
rect 660 -3417 661 -3415
rect 660 -3423 661 -3421
rect 667 -3417 668 -3415
rect 674 -3417 675 -3415
rect 674 -3423 675 -3421
rect 681 -3417 682 -3415
rect 681 -3423 682 -3421
rect 688 -3417 689 -3415
rect 695 -3417 696 -3415
rect 695 -3423 696 -3421
rect 702 -3417 703 -3415
rect 702 -3423 703 -3421
rect 709 -3417 710 -3415
rect 709 -3423 710 -3421
rect 716 -3417 717 -3415
rect 716 -3423 717 -3421
rect 723 -3417 724 -3415
rect 726 -3417 727 -3415
rect 723 -3423 724 -3421
rect 726 -3423 727 -3421
rect 730 -3417 731 -3415
rect 730 -3423 731 -3421
rect 737 -3417 738 -3415
rect 737 -3423 738 -3421
rect 744 -3417 745 -3415
rect 744 -3423 745 -3421
rect 751 -3417 752 -3415
rect 751 -3423 752 -3421
rect 758 -3417 759 -3415
rect 758 -3423 759 -3421
rect 765 -3417 766 -3415
rect 765 -3423 766 -3421
rect 772 -3417 773 -3415
rect 772 -3423 773 -3421
rect 779 -3417 780 -3415
rect 779 -3423 780 -3421
rect 786 -3417 787 -3415
rect 786 -3423 787 -3421
rect 793 -3417 794 -3415
rect 793 -3423 794 -3421
rect 800 -3417 801 -3415
rect 803 -3417 804 -3415
rect 807 -3417 808 -3415
rect 807 -3423 808 -3421
rect 814 -3417 815 -3415
rect 814 -3423 815 -3421
rect 821 -3417 822 -3415
rect 821 -3423 822 -3421
rect 828 -3417 829 -3415
rect 828 -3423 829 -3421
rect 835 -3417 836 -3415
rect 835 -3423 836 -3421
rect 842 -3417 843 -3415
rect 842 -3423 843 -3421
rect 845 -3423 846 -3421
rect 849 -3417 850 -3415
rect 849 -3423 850 -3421
rect 859 -3417 860 -3415
rect 859 -3423 860 -3421
rect 863 -3417 864 -3415
rect 863 -3423 864 -3421
rect 870 -3417 871 -3415
rect 870 -3423 871 -3421
rect 877 -3417 878 -3415
rect 877 -3423 878 -3421
rect 884 -3417 885 -3415
rect 884 -3423 885 -3421
rect 891 -3417 892 -3415
rect 891 -3423 892 -3421
rect 901 -3417 902 -3415
rect 898 -3423 899 -3421
rect 901 -3423 902 -3421
rect 905 -3417 906 -3415
rect 905 -3423 906 -3421
rect 912 -3417 913 -3415
rect 912 -3423 913 -3421
rect 919 -3417 920 -3415
rect 919 -3423 920 -3421
rect 922 -3423 923 -3421
rect 926 -3417 927 -3415
rect 926 -3423 927 -3421
rect 933 -3417 934 -3415
rect 936 -3417 937 -3415
rect 940 -3417 941 -3415
rect 940 -3423 941 -3421
rect 947 -3417 948 -3415
rect 947 -3423 948 -3421
rect 954 -3417 955 -3415
rect 954 -3423 955 -3421
rect 961 -3417 962 -3415
rect 961 -3423 962 -3421
rect 968 -3417 969 -3415
rect 968 -3423 969 -3421
rect 975 -3417 976 -3415
rect 975 -3423 976 -3421
rect 982 -3417 983 -3415
rect 982 -3423 983 -3421
rect 989 -3417 990 -3415
rect 992 -3417 993 -3415
rect 989 -3423 990 -3421
rect 992 -3423 993 -3421
rect 996 -3417 997 -3415
rect 996 -3423 997 -3421
rect 1003 -3417 1004 -3415
rect 1003 -3423 1004 -3421
rect 1010 -3417 1011 -3415
rect 1010 -3423 1011 -3421
rect 1017 -3417 1018 -3415
rect 1017 -3423 1018 -3421
rect 1024 -3417 1025 -3415
rect 1027 -3417 1028 -3415
rect 1031 -3417 1032 -3415
rect 1034 -3417 1035 -3415
rect 1031 -3423 1032 -3421
rect 1034 -3423 1035 -3421
rect 1038 -3417 1039 -3415
rect 1038 -3423 1039 -3421
rect 1045 -3417 1046 -3415
rect 1045 -3423 1046 -3421
rect 1052 -3417 1053 -3415
rect 1052 -3423 1053 -3421
rect 1059 -3417 1060 -3415
rect 1059 -3423 1060 -3421
rect 1066 -3417 1067 -3415
rect 1066 -3423 1067 -3421
rect 1069 -3423 1070 -3421
rect 1073 -3417 1074 -3415
rect 1073 -3423 1074 -3421
rect 1080 -3417 1081 -3415
rect 1080 -3423 1081 -3421
rect 1087 -3417 1088 -3415
rect 1087 -3423 1088 -3421
rect 1094 -3417 1095 -3415
rect 1094 -3423 1095 -3421
rect 1101 -3417 1102 -3415
rect 1101 -3423 1102 -3421
rect 1108 -3417 1109 -3415
rect 1108 -3423 1109 -3421
rect 1115 -3417 1116 -3415
rect 1115 -3423 1116 -3421
rect 1122 -3417 1123 -3415
rect 1125 -3417 1126 -3415
rect 1122 -3423 1123 -3421
rect 1125 -3423 1126 -3421
rect 1136 -3417 1137 -3415
rect 1136 -3423 1137 -3421
rect 1143 -3417 1144 -3415
rect 1143 -3423 1144 -3421
rect 1160 -3417 1161 -3415
rect 1157 -3423 1158 -3421
rect 1171 -3417 1172 -3415
rect 1171 -3423 1172 -3421
rect 1178 -3417 1179 -3415
rect 1178 -3423 1179 -3421
rect 1185 -3417 1186 -3415
rect 1185 -3423 1186 -3421
rect 1192 -3417 1193 -3415
rect 1192 -3423 1193 -3421
rect 1199 -3417 1200 -3415
rect 1199 -3423 1200 -3421
rect 1206 -3417 1207 -3415
rect 1209 -3417 1210 -3415
rect 1206 -3423 1207 -3421
rect 1213 -3417 1214 -3415
rect 1213 -3423 1214 -3421
rect 1220 -3417 1221 -3415
rect 1220 -3423 1221 -3421
rect 1227 -3417 1228 -3415
rect 1227 -3423 1228 -3421
rect 1234 -3417 1235 -3415
rect 1234 -3423 1235 -3421
rect 1241 -3417 1242 -3415
rect 1241 -3423 1242 -3421
rect 1248 -3417 1249 -3415
rect 1248 -3423 1249 -3421
rect 1255 -3417 1256 -3415
rect 1255 -3423 1256 -3421
rect 1262 -3417 1263 -3415
rect 1262 -3423 1263 -3421
rect 1269 -3417 1270 -3415
rect 1269 -3423 1270 -3421
rect 1276 -3423 1277 -3421
rect 1283 -3417 1284 -3415
rect 1283 -3423 1284 -3421
rect 1290 -3417 1291 -3415
rect 1290 -3423 1291 -3421
rect 1297 -3417 1298 -3415
rect 1297 -3423 1298 -3421
rect 1304 -3417 1305 -3415
rect 1307 -3423 1308 -3421
rect 1332 -3417 1333 -3415
rect 1332 -3423 1333 -3421
rect 1346 -3417 1347 -3415
rect 1346 -3423 1347 -3421
rect 1360 -3417 1361 -3415
rect 1360 -3423 1361 -3421
rect 1367 -3417 1368 -3415
rect 1367 -3423 1368 -3421
rect 1374 -3417 1375 -3415
rect 1377 -3417 1378 -3415
rect 1374 -3423 1375 -3421
rect 1381 -3417 1382 -3415
rect 1381 -3423 1382 -3421
rect 1451 -3417 1452 -3415
rect 1451 -3423 1452 -3421
rect 1458 -3417 1459 -3415
rect 1458 -3423 1459 -3421
rect 1465 -3417 1466 -3415
rect 1465 -3423 1466 -3421
rect 1472 -3417 1473 -3415
rect 1472 -3423 1473 -3421
rect 1500 -3417 1501 -3415
rect 1500 -3423 1501 -3421
rect 1521 -3417 1522 -3415
rect 1521 -3423 1522 -3421
rect 1528 -3417 1529 -3415
rect 1528 -3423 1529 -3421
rect 1549 -3417 1550 -3415
rect 1552 -3417 1553 -3415
rect 1584 -3417 1585 -3415
rect 1587 -3417 1588 -3415
rect 1584 -3423 1585 -3421
rect 1612 -3417 1613 -3415
rect 1612 -3423 1613 -3421
rect 1647 -3417 1648 -3415
rect 1647 -3423 1648 -3421
rect 1654 -3417 1655 -3415
rect 1654 -3423 1655 -3421
rect 1724 -3417 1725 -3415
rect 1724 -3423 1725 -3421
rect 1731 -3417 1732 -3415
rect 1731 -3423 1732 -3421
rect 1738 -3417 1739 -3415
rect 1738 -3423 1739 -3421
rect 1759 -3417 1760 -3415
rect 1759 -3423 1760 -3421
rect 1769 -3417 1770 -3415
rect 1766 -3423 1767 -3421
rect 1780 -3417 1781 -3415
rect 1780 -3423 1781 -3421
rect 1787 -3417 1788 -3415
rect 1787 -3423 1788 -3421
rect 1801 -3417 1802 -3415
rect 1801 -3423 1802 -3421
rect 1808 -3417 1809 -3415
rect 1811 -3417 1812 -3415
rect 1808 -3423 1809 -3421
rect 1822 -3417 1823 -3415
rect 1822 -3423 1823 -3421
rect 1829 -3417 1830 -3415
rect 1829 -3423 1830 -3421
rect 1836 -3417 1837 -3415
rect 1836 -3423 1837 -3421
rect 1843 -3417 1844 -3415
rect 1843 -3423 1844 -3421
rect 1850 -3417 1851 -3415
rect 1850 -3423 1851 -3421
rect 1857 -3417 1858 -3415
rect 1857 -3423 1858 -3421
rect 1864 -3417 1865 -3415
rect 1864 -3423 1865 -3421
rect 1867 -3423 1868 -3421
rect 1871 -3417 1872 -3415
rect 1871 -3423 1872 -3421
rect 1955 -3417 1956 -3415
rect 1955 -3423 1956 -3421
rect 1962 -3417 1963 -3415
rect 1962 -3423 1963 -3421
rect 2025 -3417 2026 -3415
rect 2028 -3417 2029 -3415
rect 2025 -3423 2026 -3421
rect 2032 -3417 2033 -3415
rect 2032 -3423 2033 -3421
rect 173 -3462 174 -3460
rect 268 -3462 269 -3460
rect 271 -3468 272 -3466
rect 324 -3462 325 -3460
rect 324 -3468 325 -3466
rect 380 -3462 381 -3460
rect 380 -3468 381 -3466
rect 415 -3462 416 -3460
rect 415 -3468 416 -3466
rect 422 -3462 423 -3460
rect 422 -3468 423 -3466
rect 439 -3468 440 -3466
rect 443 -3462 444 -3460
rect 443 -3468 444 -3466
rect 457 -3462 458 -3460
rect 457 -3468 458 -3466
rect 464 -3462 465 -3460
rect 467 -3462 468 -3460
rect 467 -3468 468 -3466
rect 485 -3462 486 -3460
rect 485 -3468 486 -3466
rect 492 -3462 493 -3460
rect 492 -3468 493 -3466
rect 499 -3462 500 -3460
rect 499 -3468 500 -3466
rect 506 -3462 507 -3460
rect 506 -3468 507 -3466
rect 513 -3462 514 -3460
rect 513 -3468 514 -3466
rect 520 -3462 521 -3460
rect 520 -3468 521 -3466
rect 523 -3468 524 -3466
rect 534 -3462 535 -3460
rect 534 -3468 535 -3466
rect 541 -3462 542 -3460
rect 541 -3468 542 -3466
rect 551 -3468 552 -3466
rect 555 -3462 556 -3460
rect 555 -3468 556 -3466
rect 562 -3462 563 -3460
rect 562 -3468 563 -3466
rect 569 -3462 570 -3460
rect 569 -3468 570 -3466
rect 576 -3462 577 -3460
rect 579 -3462 580 -3460
rect 579 -3468 580 -3466
rect 583 -3462 584 -3460
rect 583 -3468 584 -3466
rect 590 -3462 591 -3460
rect 593 -3462 594 -3460
rect 590 -3468 591 -3466
rect 597 -3462 598 -3460
rect 597 -3468 598 -3466
rect 604 -3462 605 -3460
rect 604 -3468 605 -3466
rect 611 -3462 612 -3460
rect 611 -3468 612 -3466
rect 621 -3462 622 -3460
rect 625 -3462 626 -3460
rect 628 -3462 629 -3460
rect 628 -3468 629 -3466
rect 632 -3462 633 -3460
rect 632 -3468 633 -3466
rect 639 -3462 640 -3460
rect 639 -3468 640 -3466
rect 642 -3468 643 -3466
rect 646 -3462 647 -3460
rect 646 -3468 647 -3466
rect 653 -3462 654 -3460
rect 653 -3468 654 -3466
rect 660 -3462 661 -3460
rect 660 -3468 661 -3466
rect 667 -3462 668 -3460
rect 667 -3468 668 -3466
rect 674 -3462 675 -3460
rect 674 -3468 675 -3466
rect 681 -3462 682 -3460
rect 684 -3462 685 -3460
rect 681 -3468 682 -3466
rect 688 -3468 689 -3466
rect 695 -3462 696 -3460
rect 695 -3468 696 -3466
rect 702 -3462 703 -3460
rect 705 -3462 706 -3460
rect 702 -3468 703 -3466
rect 705 -3468 706 -3466
rect 709 -3462 710 -3460
rect 709 -3468 710 -3466
rect 716 -3462 717 -3460
rect 716 -3468 717 -3466
rect 723 -3462 724 -3460
rect 723 -3468 724 -3466
rect 730 -3462 731 -3460
rect 730 -3468 731 -3466
rect 737 -3462 738 -3460
rect 737 -3468 738 -3466
rect 744 -3462 745 -3460
rect 744 -3468 745 -3466
rect 751 -3462 752 -3460
rect 751 -3468 752 -3466
rect 758 -3462 759 -3460
rect 758 -3468 759 -3466
rect 779 -3462 780 -3460
rect 779 -3468 780 -3466
rect 793 -3462 794 -3460
rect 793 -3468 794 -3466
rect 800 -3462 801 -3460
rect 800 -3468 801 -3466
rect 807 -3462 808 -3460
rect 807 -3468 808 -3466
rect 814 -3462 815 -3460
rect 814 -3468 815 -3466
rect 821 -3462 822 -3460
rect 821 -3468 822 -3466
rect 828 -3462 829 -3460
rect 828 -3468 829 -3466
rect 835 -3462 836 -3460
rect 835 -3468 836 -3466
rect 842 -3462 843 -3460
rect 842 -3468 843 -3466
rect 849 -3462 850 -3460
rect 849 -3468 850 -3466
rect 877 -3462 878 -3460
rect 877 -3468 878 -3466
rect 884 -3462 885 -3460
rect 884 -3468 885 -3466
rect 915 -3462 916 -3460
rect 912 -3468 913 -3466
rect 915 -3468 916 -3466
rect 922 -3462 923 -3460
rect 919 -3468 920 -3466
rect 922 -3468 923 -3466
rect 954 -3462 955 -3460
rect 954 -3468 955 -3466
rect 975 -3462 976 -3460
rect 975 -3468 976 -3466
rect 996 -3462 997 -3460
rect 1003 -3462 1004 -3460
rect 1003 -3468 1004 -3466
rect 1010 -3462 1011 -3460
rect 1010 -3468 1011 -3466
rect 1017 -3462 1018 -3460
rect 1017 -3468 1018 -3466
rect 1024 -3462 1025 -3460
rect 1024 -3468 1025 -3466
rect 1031 -3462 1032 -3460
rect 1031 -3468 1032 -3466
rect 1038 -3462 1039 -3460
rect 1038 -3468 1039 -3466
rect 1045 -3462 1046 -3460
rect 1045 -3468 1046 -3466
rect 1052 -3462 1053 -3460
rect 1052 -3468 1053 -3466
rect 1059 -3462 1060 -3460
rect 1059 -3468 1060 -3466
rect 1062 -3468 1063 -3466
rect 1066 -3462 1067 -3460
rect 1066 -3468 1067 -3466
rect 1073 -3462 1074 -3460
rect 1073 -3468 1074 -3466
rect 1080 -3462 1081 -3460
rect 1083 -3462 1084 -3460
rect 1083 -3468 1084 -3466
rect 1087 -3462 1088 -3460
rect 1087 -3468 1088 -3466
rect 1094 -3462 1095 -3460
rect 1094 -3468 1095 -3466
rect 1101 -3462 1102 -3460
rect 1101 -3468 1102 -3466
rect 1108 -3462 1109 -3460
rect 1108 -3468 1109 -3466
rect 1125 -3462 1126 -3460
rect 1122 -3468 1123 -3466
rect 1125 -3468 1126 -3466
rect 1129 -3462 1130 -3460
rect 1129 -3468 1130 -3466
rect 1157 -3462 1158 -3460
rect 1157 -3468 1158 -3466
rect 1164 -3462 1165 -3460
rect 1164 -3468 1165 -3466
rect 1171 -3462 1172 -3460
rect 1171 -3468 1172 -3466
rect 1178 -3462 1179 -3460
rect 1181 -3462 1182 -3460
rect 1178 -3468 1179 -3466
rect 1185 -3462 1186 -3460
rect 1185 -3468 1186 -3466
rect 1192 -3462 1193 -3460
rect 1192 -3468 1193 -3466
rect 1199 -3462 1200 -3460
rect 1199 -3468 1200 -3466
rect 1206 -3462 1207 -3460
rect 1206 -3468 1207 -3466
rect 1213 -3462 1214 -3460
rect 1213 -3468 1214 -3466
rect 1220 -3462 1221 -3460
rect 1220 -3468 1221 -3466
rect 1227 -3462 1228 -3460
rect 1227 -3468 1228 -3466
rect 1234 -3462 1235 -3460
rect 1234 -3468 1235 -3466
rect 1241 -3462 1242 -3460
rect 1241 -3468 1242 -3466
rect 1248 -3462 1249 -3460
rect 1248 -3468 1249 -3466
rect 1286 -3462 1287 -3460
rect 1283 -3468 1284 -3466
rect 1290 -3462 1291 -3460
rect 1290 -3468 1291 -3466
rect 1304 -3462 1305 -3460
rect 1307 -3462 1308 -3460
rect 1304 -3468 1305 -3466
rect 1307 -3468 1308 -3466
rect 1311 -3462 1312 -3460
rect 1311 -3468 1312 -3466
rect 1318 -3462 1319 -3460
rect 1321 -3462 1322 -3460
rect 1318 -3468 1319 -3466
rect 1325 -3462 1326 -3460
rect 1325 -3468 1326 -3466
rect 1332 -3462 1333 -3460
rect 1332 -3468 1333 -3466
rect 1360 -3462 1361 -3460
rect 1360 -3468 1361 -3466
rect 1437 -3462 1438 -3460
rect 1437 -3468 1438 -3466
rect 1444 -3462 1445 -3460
rect 1444 -3468 1445 -3466
rect 1451 -3462 1452 -3460
rect 1451 -3468 1452 -3466
rect 1458 -3462 1459 -3460
rect 1461 -3462 1462 -3460
rect 1458 -3468 1459 -3466
rect 1465 -3462 1466 -3460
rect 1465 -3468 1466 -3466
rect 1493 -3462 1494 -3460
rect 1493 -3468 1494 -3466
rect 1500 -3462 1501 -3460
rect 1500 -3468 1501 -3466
rect 1514 -3462 1515 -3460
rect 1514 -3468 1515 -3466
rect 1521 -3462 1522 -3460
rect 1521 -3468 1522 -3466
rect 1626 -3462 1627 -3460
rect 1629 -3462 1630 -3460
rect 1640 -3462 1641 -3460
rect 1640 -3468 1641 -3466
rect 1724 -3462 1725 -3460
rect 1724 -3468 1725 -3466
rect 1731 -3462 1732 -3460
rect 1731 -3468 1732 -3466
rect 1748 -3462 1749 -3460
rect 1745 -3468 1746 -3466
rect 1766 -3462 1767 -3460
rect 1766 -3468 1767 -3466
rect 1780 -3462 1781 -3460
rect 1780 -3468 1781 -3466
rect 1794 -3462 1795 -3460
rect 1794 -3468 1795 -3466
rect 1822 -3462 1823 -3460
rect 1822 -3468 1823 -3466
rect 1829 -3462 1830 -3460
rect 1829 -3468 1830 -3466
rect 1836 -3468 1837 -3466
rect 1839 -3468 1840 -3466
rect 1843 -3462 1844 -3460
rect 1843 -3468 1844 -3466
rect 1850 -3462 1851 -3460
rect 1850 -3468 1851 -3466
rect 1857 -3462 1858 -3460
rect 1860 -3462 1861 -3460
rect 1860 -3468 1861 -3466
rect 1864 -3462 1865 -3460
rect 1867 -3462 1868 -3460
rect 1864 -3468 1865 -3466
rect 1871 -3462 1872 -3460
rect 1871 -3468 1872 -3466
rect 1955 -3462 1956 -3460
rect 1955 -3468 1956 -3466
rect 1962 -3462 1963 -3460
rect 1962 -3468 1963 -3466
rect 2025 -3462 2026 -3460
rect 2025 -3468 2026 -3466
rect 2028 -3468 2029 -3466
rect 2032 -3462 2033 -3460
rect 2032 -3468 2033 -3466
rect 331 -3491 332 -3489
rect 331 -3497 332 -3495
rect 366 -3491 367 -3489
rect 369 -3491 370 -3489
rect 387 -3491 388 -3489
rect 387 -3497 388 -3495
rect 394 -3491 395 -3489
rect 394 -3497 395 -3495
rect 429 -3491 430 -3489
rect 429 -3497 430 -3495
rect 432 -3497 433 -3495
rect 464 -3491 465 -3489
rect 464 -3497 465 -3495
rect 471 -3491 472 -3489
rect 471 -3497 472 -3495
rect 478 -3491 479 -3489
rect 478 -3497 479 -3495
rect 485 -3491 486 -3489
rect 485 -3497 486 -3495
rect 523 -3491 524 -3489
rect 523 -3497 524 -3495
rect 534 -3491 535 -3489
rect 534 -3497 535 -3495
rect 541 -3491 542 -3489
rect 541 -3497 542 -3495
rect 569 -3491 570 -3489
rect 569 -3497 570 -3495
rect 583 -3491 584 -3489
rect 583 -3497 584 -3495
rect 590 -3491 591 -3489
rect 590 -3497 591 -3495
rect 604 -3491 605 -3489
rect 604 -3497 605 -3495
rect 611 -3491 612 -3489
rect 611 -3497 612 -3495
rect 618 -3491 619 -3489
rect 618 -3497 619 -3495
rect 632 -3491 633 -3489
rect 632 -3497 633 -3495
rect 639 -3491 640 -3489
rect 639 -3497 640 -3495
rect 646 -3491 647 -3489
rect 646 -3497 647 -3495
rect 653 -3491 654 -3489
rect 653 -3497 654 -3495
rect 656 -3497 657 -3495
rect 681 -3491 682 -3489
rect 681 -3497 682 -3495
rect 716 -3491 717 -3489
rect 716 -3497 717 -3495
rect 737 -3491 738 -3489
rect 737 -3497 738 -3495
rect 744 -3491 745 -3489
rect 744 -3497 745 -3495
rect 751 -3491 752 -3489
rect 751 -3497 752 -3495
rect 758 -3491 759 -3489
rect 758 -3497 759 -3495
rect 765 -3491 766 -3489
rect 765 -3497 766 -3495
rect 772 -3491 773 -3489
rect 772 -3497 773 -3495
rect 779 -3491 780 -3489
rect 779 -3497 780 -3495
rect 786 -3491 787 -3489
rect 789 -3491 790 -3489
rect 793 -3491 794 -3489
rect 793 -3497 794 -3495
rect 814 -3491 815 -3489
rect 814 -3497 815 -3495
rect 828 -3491 829 -3489
rect 828 -3497 829 -3495
rect 842 -3491 843 -3489
rect 842 -3497 843 -3495
rect 866 -3491 867 -3489
rect 863 -3497 864 -3495
rect 866 -3497 867 -3495
rect 870 -3491 871 -3489
rect 870 -3497 871 -3495
rect 887 -3491 888 -3489
rect 884 -3497 885 -3495
rect 898 -3491 899 -3489
rect 898 -3497 899 -3495
rect 975 -3491 976 -3489
rect 975 -3497 976 -3495
rect 996 -3497 997 -3495
rect 1010 -3491 1011 -3489
rect 1010 -3497 1011 -3495
rect 1017 -3491 1018 -3489
rect 1017 -3497 1018 -3495
rect 1024 -3491 1025 -3489
rect 1024 -3497 1025 -3495
rect 1031 -3491 1032 -3489
rect 1031 -3497 1032 -3495
rect 1038 -3491 1039 -3489
rect 1038 -3497 1039 -3495
rect 1045 -3491 1046 -3489
rect 1045 -3497 1046 -3495
rect 1052 -3491 1053 -3489
rect 1052 -3497 1053 -3495
rect 1059 -3491 1060 -3489
rect 1059 -3497 1060 -3495
rect 1066 -3491 1067 -3489
rect 1066 -3497 1067 -3495
rect 1080 -3491 1081 -3489
rect 1080 -3497 1081 -3495
rect 1143 -3491 1144 -3489
rect 1143 -3497 1144 -3495
rect 1178 -3491 1179 -3489
rect 1178 -3497 1179 -3495
rect 1192 -3491 1193 -3489
rect 1192 -3497 1193 -3495
rect 1234 -3491 1235 -3489
rect 1234 -3497 1235 -3495
rect 1241 -3491 1242 -3489
rect 1241 -3497 1242 -3495
rect 1248 -3491 1249 -3489
rect 1248 -3497 1249 -3495
rect 1251 -3497 1252 -3495
rect 1255 -3491 1256 -3489
rect 1255 -3497 1256 -3495
rect 1262 -3491 1263 -3489
rect 1262 -3497 1263 -3495
rect 1269 -3491 1270 -3489
rect 1272 -3491 1273 -3489
rect 1276 -3491 1277 -3489
rect 1276 -3497 1277 -3495
rect 1286 -3491 1287 -3489
rect 1283 -3497 1284 -3495
rect 1290 -3491 1291 -3489
rect 1290 -3497 1291 -3495
rect 1304 -3491 1305 -3489
rect 1304 -3497 1305 -3495
rect 1311 -3491 1312 -3489
rect 1311 -3497 1312 -3495
rect 1360 -3491 1361 -3489
rect 1360 -3497 1361 -3495
rect 1430 -3491 1431 -3489
rect 1433 -3491 1434 -3489
rect 1430 -3497 1431 -3495
rect 1437 -3491 1438 -3489
rect 1437 -3497 1438 -3495
rect 1493 -3491 1494 -3489
rect 1493 -3497 1494 -3495
rect 1500 -3491 1501 -3489
rect 1503 -3491 1504 -3489
rect 1500 -3497 1501 -3495
rect 1507 -3491 1508 -3489
rect 1507 -3497 1508 -3495
rect 1514 -3491 1515 -3489
rect 1514 -3497 1515 -3495
rect 1521 -3491 1522 -3489
rect 1521 -3497 1522 -3495
rect 1570 -3491 1571 -3489
rect 1570 -3497 1571 -3495
rect 1640 -3491 1641 -3489
rect 1640 -3497 1641 -3495
rect 1724 -3491 1725 -3489
rect 1727 -3491 1728 -3489
rect 1724 -3497 1725 -3495
rect 1731 -3491 1732 -3489
rect 1731 -3497 1732 -3495
rect 1780 -3491 1781 -3489
rect 1780 -3497 1781 -3495
rect 1790 -3491 1791 -3489
rect 1790 -3497 1791 -3495
rect 1843 -3491 1844 -3489
rect 1843 -3497 1844 -3495
rect 1850 -3491 1851 -3489
rect 1850 -3497 1851 -3495
rect 1864 -3491 1865 -3489
rect 1864 -3497 1865 -3495
rect 1955 -3491 1956 -3489
rect 1958 -3491 1959 -3489
rect 2025 -3491 2026 -3489
rect 2028 -3491 2029 -3489
rect 2025 -3497 2026 -3495
rect 2032 -3491 2033 -3489
rect 2032 -3497 2033 -3495
rect 338 -3514 339 -3512
rect 394 -3514 395 -3512
rect 394 -3520 395 -3518
rect 429 -3514 430 -3512
rect 429 -3520 430 -3518
rect 464 -3514 465 -3512
rect 464 -3520 465 -3518
rect 478 -3514 479 -3512
rect 478 -3520 479 -3518
rect 541 -3514 542 -3512
rect 541 -3520 542 -3518
rect 548 -3514 549 -3512
rect 548 -3520 549 -3518
rect 576 -3514 577 -3512
rect 576 -3520 577 -3518
rect 583 -3514 584 -3512
rect 583 -3520 584 -3518
rect 604 -3514 605 -3512
rect 604 -3520 605 -3518
rect 611 -3514 612 -3512
rect 611 -3520 612 -3518
rect 618 -3514 619 -3512
rect 618 -3520 619 -3518
rect 625 -3514 626 -3512
rect 625 -3520 626 -3518
rect 632 -3514 633 -3512
rect 632 -3520 633 -3518
rect 639 -3514 640 -3512
rect 639 -3520 640 -3518
rect 709 -3514 710 -3512
rect 709 -3520 710 -3518
rect 730 -3514 731 -3512
rect 730 -3520 731 -3518
rect 737 -3514 738 -3512
rect 737 -3520 738 -3518
rect 744 -3514 745 -3512
rect 744 -3520 745 -3518
rect 751 -3514 752 -3512
rect 751 -3520 752 -3518
rect 758 -3514 759 -3512
rect 758 -3520 759 -3518
rect 765 -3514 766 -3512
rect 765 -3520 766 -3518
rect 775 -3514 776 -3512
rect 772 -3520 773 -3518
rect 775 -3520 776 -3518
rect 779 -3514 780 -3512
rect 779 -3520 780 -3518
rect 789 -3514 790 -3512
rect 786 -3520 787 -3518
rect 789 -3520 790 -3518
rect 793 -3514 794 -3512
rect 793 -3520 794 -3518
rect 800 -3514 801 -3512
rect 800 -3520 801 -3518
rect 810 -3514 811 -3512
rect 810 -3520 811 -3518
rect 891 -3514 892 -3512
rect 891 -3520 892 -3518
rect 968 -3514 969 -3512
rect 968 -3520 969 -3518
rect 1003 -3514 1004 -3512
rect 1003 -3520 1004 -3518
rect 1010 -3514 1011 -3512
rect 1010 -3520 1011 -3518
rect 1017 -3514 1018 -3512
rect 1017 -3520 1018 -3518
rect 1024 -3514 1025 -3512
rect 1024 -3520 1025 -3518
rect 1031 -3514 1032 -3512
rect 1031 -3520 1032 -3518
rect 1038 -3514 1039 -3512
rect 1038 -3520 1039 -3518
rect 1045 -3514 1046 -3512
rect 1052 -3514 1053 -3512
rect 1052 -3520 1053 -3518
rect 1059 -3514 1060 -3512
rect 1062 -3514 1063 -3512
rect 1059 -3520 1060 -3518
rect 1066 -3514 1067 -3512
rect 1066 -3520 1067 -3518
rect 1122 -3514 1123 -3512
rect 1122 -3520 1123 -3518
rect 1150 -3514 1151 -3512
rect 1150 -3520 1151 -3518
rect 1160 -3514 1161 -3512
rect 1157 -3520 1158 -3518
rect 1160 -3520 1161 -3518
rect 1206 -3514 1207 -3512
rect 1206 -3520 1207 -3518
rect 1234 -3514 1235 -3512
rect 1234 -3520 1235 -3518
rect 1360 -3514 1361 -3512
rect 1360 -3520 1361 -3518
rect 1367 -3514 1368 -3512
rect 1367 -3520 1368 -3518
rect 1507 -3514 1508 -3512
rect 1507 -3520 1508 -3518
rect 1510 -3520 1511 -3518
rect 1514 -3514 1515 -3512
rect 1514 -3520 1515 -3518
rect 1521 -3514 1522 -3512
rect 1521 -3520 1522 -3518
rect 1612 -3514 1613 -3512
rect 1612 -3520 1613 -3518
rect 1640 -3514 1641 -3512
rect 1640 -3520 1641 -3518
rect 1850 -3514 1851 -3512
rect 1850 -3520 1851 -3518
rect 1857 -3514 1858 -3512
rect 1860 -3514 1861 -3512
rect 1857 -3520 1858 -3518
rect 2025 -3514 2026 -3512
rect 2025 -3520 2026 -3518
rect 2032 -3514 2033 -3512
rect 2032 -3520 2033 -3518
rect 394 -3533 395 -3531
rect 394 -3539 395 -3537
rect 408 -3533 409 -3531
rect 408 -3539 409 -3537
rect 464 -3533 465 -3531
rect 464 -3539 465 -3537
rect 471 -3539 472 -3537
rect 474 -3539 475 -3537
rect 478 -3533 479 -3531
rect 478 -3539 479 -3537
rect 541 -3533 542 -3531
rect 541 -3539 542 -3537
rect 548 -3533 549 -3531
rect 548 -3539 549 -3537
rect 576 -3533 577 -3531
rect 576 -3539 577 -3537
rect 583 -3533 584 -3531
rect 583 -3539 584 -3537
rect 604 -3533 605 -3531
rect 604 -3539 605 -3537
rect 611 -3533 612 -3531
rect 611 -3539 612 -3537
rect 618 -3533 619 -3531
rect 618 -3539 619 -3537
rect 625 -3533 626 -3531
rect 632 -3533 633 -3531
rect 635 -3533 636 -3531
rect 635 -3539 636 -3537
rect 639 -3533 640 -3531
rect 639 -3539 640 -3537
rect 646 -3533 647 -3531
rect 646 -3539 647 -3537
rect 709 -3533 710 -3531
rect 709 -3539 710 -3537
rect 716 -3533 717 -3531
rect 716 -3539 717 -3537
rect 723 -3533 724 -3531
rect 723 -3539 724 -3537
rect 730 -3533 731 -3531
rect 730 -3539 731 -3537
rect 740 -3533 741 -3531
rect 740 -3539 741 -3537
rect 744 -3533 745 -3531
rect 744 -3539 745 -3537
rect 765 -3533 766 -3531
rect 765 -3539 766 -3537
rect 786 -3533 787 -3531
rect 786 -3539 787 -3537
rect 793 -3533 794 -3531
rect 793 -3539 794 -3537
rect 926 -3533 927 -3531
rect 926 -3539 927 -3537
rect 971 -3533 972 -3531
rect 968 -3539 969 -3537
rect 1010 -3533 1011 -3531
rect 1010 -3539 1011 -3537
rect 1024 -3533 1025 -3531
rect 1027 -3533 1028 -3531
rect 1027 -3539 1028 -3537
rect 1031 -3533 1032 -3531
rect 1031 -3539 1032 -3537
rect 1038 -3533 1039 -3531
rect 1038 -3539 1039 -3537
rect 1045 -3539 1046 -3537
rect 1059 -3533 1060 -3531
rect 1059 -3539 1060 -3537
rect 1066 -3533 1067 -3531
rect 1066 -3539 1067 -3537
rect 1213 -3533 1214 -3531
rect 1213 -3539 1214 -3537
rect 1223 -3533 1224 -3531
rect 1223 -3539 1224 -3537
rect 1507 -3533 1508 -3531
rect 1510 -3533 1511 -3531
rect 1507 -3539 1508 -3537
rect 1514 -3533 1515 -3531
rect 1514 -3539 1515 -3537
rect 1521 -3533 1522 -3531
rect 1521 -3539 1522 -3537
rect 1633 -3533 1634 -3531
rect 1633 -3539 1634 -3537
rect 1640 -3533 1641 -3531
rect 1640 -3539 1641 -3537
rect 2025 -3533 2026 -3531
rect 2025 -3539 2026 -3537
rect 2032 -3533 2033 -3531
rect 2032 -3539 2033 -3537
rect 401 -3548 402 -3546
rect 401 -3554 402 -3552
rect 408 -3548 409 -3546
rect 541 -3548 542 -3546
rect 541 -3554 542 -3552
rect 548 -3554 549 -3552
rect 551 -3554 552 -3552
rect 555 -3548 556 -3546
rect 555 -3554 556 -3552
rect 583 -3548 584 -3546
rect 586 -3554 587 -3552
rect 590 -3548 591 -3546
rect 590 -3554 591 -3552
rect 604 -3548 605 -3546
rect 604 -3554 605 -3552
rect 607 -3554 608 -3552
rect 611 -3548 612 -3546
rect 611 -3554 612 -3552
rect 618 -3548 619 -3546
rect 618 -3554 619 -3552
rect 646 -3548 647 -3546
rect 646 -3554 647 -3552
rect 702 -3548 703 -3546
rect 702 -3554 703 -3552
rect 716 -3548 717 -3546
rect 716 -3554 717 -3552
rect 723 -3548 724 -3546
rect 723 -3554 724 -3552
rect 730 -3548 731 -3546
rect 730 -3554 731 -3552
rect 758 -3548 759 -3546
rect 758 -3554 759 -3552
rect 789 -3548 790 -3546
rect 789 -3554 790 -3552
rect 793 -3548 794 -3546
rect 793 -3554 794 -3552
rect 1020 -3548 1021 -3546
rect 1017 -3554 1018 -3552
rect 1038 -3548 1039 -3546
rect 1038 -3554 1039 -3552
rect 1059 -3548 1060 -3546
rect 1059 -3554 1060 -3552
rect 1507 -3548 1508 -3546
rect 1507 -3554 1508 -3552
rect 1514 -3548 1515 -3546
rect 1514 -3554 1515 -3552
rect 1521 -3548 1522 -3546
rect 1521 -3554 1522 -3552
rect 1640 -3548 1641 -3546
rect 1640 -3554 1641 -3552
rect 1647 -3548 1648 -3546
rect 1647 -3554 1648 -3552
rect 2025 -3548 2026 -3546
rect 2025 -3554 2026 -3552
rect 2032 -3548 2033 -3546
rect 2032 -3554 2033 -3552
rect 401 -3563 402 -3561
rect 401 -3569 402 -3567
rect 408 -3569 409 -3567
rect 604 -3563 605 -3561
rect 607 -3563 608 -3561
rect 604 -3569 605 -3567
rect 611 -3563 612 -3561
rect 611 -3569 612 -3567
rect 618 -3563 619 -3561
rect 618 -3569 619 -3567
rect 649 -3563 650 -3561
rect 702 -3563 703 -3561
rect 702 -3569 703 -3567
rect 716 -3563 717 -3561
rect 716 -3569 717 -3567
rect 723 -3563 724 -3561
rect 723 -3569 724 -3567
rect 730 -3563 731 -3561
rect 730 -3569 731 -3567
rect 758 -3563 759 -3561
rect 758 -3569 759 -3567
rect 1062 -3569 1063 -3567
rect 1066 -3563 1067 -3561
rect 1066 -3569 1067 -3567
rect 1514 -3563 1515 -3561
rect 1517 -3563 1518 -3561
rect 1514 -3569 1515 -3567
rect 1521 -3563 1522 -3561
rect 1521 -3569 1522 -3567
rect 1640 -3563 1641 -3561
rect 1640 -3569 1641 -3567
rect 1647 -3563 1648 -3561
rect 1647 -3569 1648 -3567
rect 2025 -3563 2026 -3561
rect 2028 -3563 2029 -3561
rect 401 -3578 402 -3576
rect 401 -3584 402 -3582
rect 408 -3578 409 -3576
rect 408 -3584 409 -3582
rect 604 -3578 605 -3576
rect 604 -3584 605 -3582
rect 611 -3578 612 -3576
rect 611 -3584 612 -3582
rect 618 -3578 619 -3576
rect 618 -3584 619 -3582
rect 702 -3578 703 -3576
rect 702 -3584 703 -3582
rect 716 -3578 717 -3576
rect 716 -3584 717 -3582
rect 723 -3578 724 -3576
rect 723 -3584 724 -3582
rect 730 -3578 731 -3576
rect 730 -3584 731 -3582
rect 758 -3578 759 -3576
rect 758 -3584 759 -3582
rect 1640 -3578 1641 -3576
rect 1640 -3584 1641 -3582
rect 1647 -3578 1648 -3576
rect 1647 -3584 1648 -3582
rect 394 -3591 395 -3589
rect 394 -3597 395 -3595
rect 401 -3591 402 -3589
rect 401 -3597 402 -3595
rect 604 -3591 605 -3589
rect 604 -3597 605 -3595
rect 611 -3591 612 -3589
rect 611 -3597 612 -3595
rect 621 -3591 622 -3589
rect 702 -3591 703 -3589
rect 702 -3597 703 -3595
rect 723 -3591 724 -3589
rect 726 -3591 727 -3589
rect 723 -3597 724 -3595
rect 730 -3591 731 -3589
rect 730 -3597 731 -3595
rect 758 -3591 759 -3589
rect 758 -3597 759 -3595
rect 1640 -3591 1641 -3589
rect 1640 -3597 1641 -3595
rect 1647 -3591 1648 -3589
rect 1647 -3597 1648 -3595
rect 394 -3602 395 -3600
rect 394 -3608 395 -3606
rect 401 -3602 402 -3600
rect 401 -3608 402 -3606
rect 604 -3602 605 -3600
rect 604 -3608 605 -3606
rect 611 -3602 612 -3600
rect 611 -3608 612 -3606
rect 702 -3602 703 -3600
rect 705 -3608 706 -3606
rect 758 -3602 759 -3600
rect 758 -3608 759 -3606
rect 1640 -3602 1641 -3600
rect 1640 -3608 1641 -3606
rect 1647 -3602 1648 -3600
rect 1647 -3608 1648 -3606
rect 394 -3613 395 -3611
rect 394 -3619 395 -3617
rect 401 -3613 402 -3611
rect 401 -3619 402 -3617
rect 604 -3613 605 -3611
rect 604 -3619 605 -3617
rect 611 -3613 612 -3611
rect 611 -3619 612 -3617
rect 695 -3613 696 -3611
rect 695 -3619 696 -3617
rect 758 -3613 759 -3611
rect 758 -3619 759 -3617
rect 1643 -3613 1644 -3611
rect 1640 -3619 1641 -3617
rect 1647 -3613 1648 -3611
rect 1647 -3619 1648 -3617
rect 394 -3624 395 -3622
rect 394 -3630 395 -3628
rect 401 -3624 402 -3622
rect 401 -3630 402 -3628
rect 604 -3624 605 -3622
rect 604 -3630 605 -3628
rect 611 -3624 612 -3622
rect 611 -3630 612 -3628
rect 695 -3624 696 -3622
rect 695 -3630 696 -3628
rect 761 -3630 762 -3628
rect 765 -3624 766 -3622
rect 765 -3630 766 -3628
rect 394 -3635 395 -3633
rect 394 -3641 395 -3639
rect 401 -3635 402 -3633
rect 401 -3641 402 -3639
rect 604 -3635 605 -3633
rect 604 -3641 605 -3639
rect 611 -3635 612 -3633
rect 611 -3641 612 -3639
rect 695 -3635 696 -3633
rect 695 -3641 696 -3639
rect 394 -3646 395 -3644
rect 394 -3652 395 -3650
rect 401 -3646 402 -3644
rect 401 -3652 402 -3650
rect 604 -3646 605 -3644
rect 604 -3652 605 -3650
rect 611 -3646 612 -3644
rect 611 -3652 612 -3650
rect 695 -3646 696 -3644
rect 695 -3652 696 -3650
rect 394 -3661 395 -3659
rect 397 -3667 398 -3665
rect 401 -3661 402 -3659
rect 401 -3667 402 -3665
rect 604 -3661 605 -3659
rect 604 -3667 605 -3665
rect 611 -3661 612 -3659
rect 611 -3667 612 -3665
rect 698 -3661 699 -3659
<< metal1 >>
rect 254 0 433 1
rect 485 0 633 1
rect 635 0 773 1
rect 796 0 815 1
rect 824 0 962 1
rect 968 0 1207 1
rect 352 -2 573 -1
rect 576 -2 682 -1
rect 688 -2 766 -1
rect 800 -2 892 -1
rect 978 -2 983 -1
rect 1038 -2 1438 -1
rect 397 -4 549 -3
rect 555 -4 584 -3
rect 604 -4 843 -3
rect 863 -4 920 -3
rect 1073 -4 1130 -3
rect 415 -6 423 -5
rect 611 -6 626 -5
rect 639 -6 846 -5
rect 884 -6 1088 -5
rect 1094 -6 1126 -5
rect 618 -8 853 -7
rect 646 -10 706 -9
rect 709 -10 916 -9
rect 663 -12 990 -11
rect 716 -14 822 -13
rect 828 -14 888 -13
rect 730 -16 804 -15
rect 810 -16 871 -15
rect 835 -18 860 -17
rect 184 -29 213 -28
rect 240 -29 398 -28
rect 404 -29 479 -28
rect 492 -29 619 -28
rect 646 -29 724 -28
rect 737 -29 759 -28
rect 765 -29 829 -28
rect 842 -29 1221 -28
rect 1234 -29 1361 -28
rect 1437 -29 1487 -28
rect 1629 -29 1634 -28
rect 198 -31 255 -30
rect 275 -31 314 -30
rect 317 -31 661 -30
rect 667 -31 741 -30
rect 744 -31 864 -30
rect 870 -31 885 -30
rect 908 -31 948 -30
rect 961 -31 1046 -30
rect 1066 -31 1102 -30
rect 1108 -31 1151 -30
rect 1206 -31 1291 -30
rect 1321 -31 1333 -30
rect 1440 -31 1760 -30
rect 296 -33 353 -32
rect 355 -33 465 -32
rect 471 -33 612 -32
rect 618 -33 626 -32
rect 660 -33 696 -32
rect 702 -33 822 -32
rect 828 -33 1039 -32
rect 1087 -33 1179 -32
rect 394 -35 486 -34
rect 499 -35 640 -34
rect 677 -35 976 -34
rect 978 -35 1004 -34
rect 1010 -35 1095 -34
rect 1132 -35 1214 -34
rect 415 -37 423 -36
rect 432 -37 591 -36
rect 611 -37 657 -36
rect 702 -37 717 -36
rect 751 -37 888 -36
rect 912 -37 1018 -36
rect 1073 -37 1088 -36
rect 1094 -37 1116 -36
rect 422 -39 447 -38
rect 485 -39 605 -38
rect 639 -39 654 -38
rect 716 -39 808 -38
rect 842 -39 899 -38
rect 926 -39 1126 -38
rect 506 -41 853 -40
rect 856 -41 1039 -40
rect 520 -43 577 -42
rect 583 -43 647 -42
rect 653 -43 962 -42
rect 982 -43 1032 -42
rect 534 -45 689 -44
rect 768 -45 864 -44
rect 870 -45 920 -44
rect 982 -45 1070 -44
rect 548 -47 598 -46
rect 604 -47 902 -46
rect 989 -47 1060 -46
rect 548 -49 573 -48
rect 583 -49 934 -48
rect 1024 -49 1074 -48
rect 569 -51 780 -50
rect 793 -51 836 -50
rect 849 -51 1081 -50
rect 569 -53 675 -52
rect 688 -53 710 -52
rect 772 -53 836 -52
rect 849 -53 913 -52
rect 709 -55 731 -54
rect 772 -55 811 -54
rect 877 -55 941 -54
rect 730 -57 969 -56
rect 800 -59 920 -58
rect 807 -61 815 -60
rect 887 -61 1053 -60
rect 681 -63 815 -62
rect 891 -63 990 -62
rect 565 -65 682 -64
rect 803 -65 892 -64
rect 915 -65 969 -64
rect 58 -76 524 -75
rect 530 -76 1242 -75
rect 1290 -76 1298 -75
rect 1332 -76 1375 -75
rect 1486 -76 1515 -75
rect 1633 -76 1641 -75
rect 1759 -76 1886 -75
rect 65 -78 227 -77
rect 233 -78 850 -77
rect 852 -78 1137 -77
rect 1157 -78 1168 -77
rect 1171 -78 1270 -77
rect 1360 -78 1424 -77
rect 72 -80 402 -79
rect 404 -80 437 -79
rect 450 -80 521 -79
rect 555 -80 661 -79
rect 674 -80 710 -79
rect 740 -80 1326 -79
rect 79 -82 353 -81
rect 359 -82 423 -81
rect 429 -82 605 -81
rect 625 -82 829 -81
rect 835 -82 906 -81
rect 919 -82 941 -81
rect 943 -82 1291 -81
rect 1321 -82 1361 -81
rect 86 -84 265 -83
rect 282 -84 500 -83
rect 513 -84 542 -83
rect 562 -84 633 -83
rect 653 -84 766 -83
rect 786 -84 822 -83
rect 856 -84 1123 -83
rect 1125 -84 1319 -83
rect 93 -86 472 -85
rect 499 -86 528 -85
rect 541 -86 612 -85
rect 660 -86 752 -85
rect 779 -86 822 -85
rect 856 -86 1011 -85
rect 1038 -86 1109 -85
rect 1115 -86 1151 -85
rect 1178 -86 1256 -85
rect 100 -88 601 -87
rect 604 -88 619 -87
rect 702 -88 829 -87
rect 863 -88 885 -87
rect 919 -88 969 -87
rect 975 -88 1284 -87
rect 107 -90 185 -89
rect 191 -90 241 -89
rect 247 -90 444 -89
rect 471 -90 976 -89
rect 989 -90 1193 -89
rect 1213 -90 1305 -89
rect 114 -92 237 -91
rect 240 -92 276 -91
rect 296 -92 332 -91
rect 338 -92 650 -91
rect 702 -92 871 -91
rect 898 -92 1214 -91
rect 1220 -92 1354 -91
rect 124 -94 304 -93
rect 310 -94 325 -93
rect 345 -94 545 -93
rect 576 -94 640 -93
rect 709 -94 717 -93
rect 751 -94 1235 -93
rect 1237 -94 1508 -93
rect 128 -96 584 -95
rect 590 -96 612 -95
rect 618 -96 958 -95
rect 961 -96 1151 -95
rect 1227 -96 1312 -95
rect 135 -98 507 -97
rect 583 -98 598 -97
rect 639 -98 836 -97
rect 863 -98 878 -97
rect 954 -98 990 -97
rect 999 -98 1095 -97
rect 1101 -98 1277 -97
rect 149 -100 353 -99
rect 366 -100 570 -99
rect 758 -100 899 -99
rect 933 -100 1102 -99
rect 1118 -100 1186 -99
rect 152 -102 290 -101
rect 310 -102 860 -101
rect 870 -102 983 -101
rect 996 -102 1095 -101
rect 156 -104 318 -103
rect 380 -104 493 -103
rect 730 -104 759 -103
rect 779 -104 909 -103
rect 912 -104 983 -103
rect 1003 -104 1165 -103
rect 163 -106 699 -105
rect 789 -106 801 -105
rect 803 -106 955 -105
rect 968 -106 1018 -105
rect 1027 -106 1235 -105
rect 170 -108 409 -107
rect 411 -108 416 -107
rect 422 -108 549 -107
rect 807 -108 1004 -107
rect 1010 -108 1144 -107
rect 177 -110 535 -109
rect 548 -110 745 -109
rect 807 -110 927 -109
rect 933 -110 1200 -109
rect 184 -112 657 -111
rect 744 -112 843 -111
rect 947 -112 997 -111
rect 1017 -112 1060 -111
rect 1073 -112 1221 -111
rect 198 -114 220 -113
rect 229 -114 318 -113
rect 373 -114 731 -113
rect 814 -114 878 -113
rect 912 -114 948 -113
rect 1024 -114 1060 -113
rect 1080 -114 1179 -113
rect 198 -116 475 -115
rect 492 -116 766 -115
rect 891 -116 1081 -115
rect 1087 -116 1207 -115
rect 205 -118 468 -117
rect 534 -118 1077 -117
rect 1087 -118 1249 -117
rect 212 -120 388 -119
rect 390 -120 570 -119
rect 597 -120 892 -119
rect 1038 -120 1112 -119
rect 261 -122 678 -121
rect 681 -122 1025 -121
rect 1045 -122 1130 -121
rect 275 -124 395 -123
rect 401 -124 486 -123
rect 646 -124 843 -123
rect 1052 -124 1067 -123
rect 296 -126 682 -125
rect 688 -126 815 -125
rect 142 -128 689 -127
rect 723 -128 1053 -127
rect 394 -130 738 -129
rect 408 -132 566 -131
rect 723 -132 794 -131
rect 121 -134 794 -133
rect 415 -136 465 -135
rect 485 -136 668 -135
rect 446 -138 591 -137
rect 667 -138 773 -137
rect 457 -140 507 -139
rect 565 -140 717 -139
rect 772 -140 1046 -139
rect 460 -142 1228 -141
rect 16 -153 262 -152
rect 282 -153 388 -152
rect 408 -153 696 -152
rect 768 -153 1347 -152
rect 1353 -153 1368 -152
rect 1374 -153 1501 -152
rect 1507 -153 1627 -152
rect 1640 -153 1669 -152
rect 1885 -153 1942 -152
rect 23 -155 108 -154
rect 114 -155 227 -154
rect 240 -155 269 -154
rect 282 -155 332 -154
rect 345 -155 531 -154
rect 541 -155 601 -154
rect 611 -155 738 -154
rect 803 -155 941 -154
rect 950 -155 1403 -154
rect 1423 -155 1494 -154
rect 1514 -155 1557 -154
rect 1566 -155 1585 -154
rect 1615 -155 1634 -154
rect 37 -157 258 -156
rect 331 -157 416 -156
rect 422 -157 444 -156
rect 450 -157 538 -156
rect 541 -157 556 -156
rect 590 -157 682 -156
rect 684 -157 927 -156
rect 1013 -157 1431 -156
rect 1542 -157 1816 -156
rect 44 -159 73 -158
rect 86 -159 766 -158
rect 814 -159 941 -158
rect 1076 -159 1249 -158
rect 1276 -159 1571 -158
rect 51 -161 80 -160
rect 93 -161 647 -160
rect 649 -161 1081 -160
rect 1090 -161 1466 -160
rect 72 -163 367 -162
rect 380 -163 409 -162
rect 429 -163 458 -162
rect 467 -163 1025 -162
rect 1073 -163 1249 -162
rect 1283 -163 1578 -162
rect 79 -165 94 -164
rect 100 -165 125 -164
rect 128 -165 153 -164
rect 163 -165 234 -164
rect 240 -165 1508 -164
rect 100 -167 566 -166
rect 618 -167 696 -166
rect 737 -167 1011 -166
rect 1073 -167 1109 -166
rect 1129 -167 1452 -166
rect 107 -169 570 -168
rect 621 -169 731 -168
rect 814 -169 839 -168
rect 849 -169 948 -168
rect 975 -169 1277 -168
rect 1290 -169 1375 -168
rect 117 -171 612 -170
rect 849 -171 878 -170
rect 884 -171 1109 -170
rect 1122 -171 1291 -170
rect 1304 -171 1445 -170
rect 121 -173 202 -172
rect 226 -173 773 -172
rect 856 -173 878 -172
rect 887 -173 1228 -172
rect 1311 -173 1473 -172
rect 128 -175 255 -174
rect 275 -175 430 -174
rect 450 -175 479 -174
rect 492 -175 598 -174
rect 667 -175 773 -174
rect 870 -175 1025 -174
rect 1059 -175 1130 -174
rect 1136 -175 1396 -174
rect 65 -177 255 -176
rect 275 -177 360 -176
rect 366 -177 895 -176
rect 905 -177 976 -176
rect 989 -177 1137 -176
rect 1150 -177 1284 -176
rect 1318 -177 1438 -176
rect 135 -179 262 -178
rect 338 -179 479 -178
rect 513 -179 563 -178
rect 569 -179 930 -178
rect 961 -179 1305 -178
rect 1325 -179 1592 -178
rect 142 -181 213 -180
rect 243 -181 272 -180
rect 296 -181 339 -180
rect 345 -181 486 -180
rect 513 -181 594 -180
rect 705 -181 1228 -180
rect 1325 -181 1333 -180
rect 1360 -181 1459 -180
rect 145 -183 157 -182
rect 163 -183 391 -182
rect 401 -183 416 -182
rect 471 -183 1011 -182
rect 1017 -183 1123 -182
rect 1164 -183 1424 -182
rect 149 -185 717 -184
rect 786 -185 906 -184
rect 919 -185 1060 -184
rect 1080 -185 1116 -184
rect 1171 -185 1389 -184
rect 156 -187 1515 -186
rect 170 -189 493 -188
rect 520 -189 990 -188
rect 1003 -189 1361 -188
rect 177 -191 360 -190
rect 373 -191 668 -190
rect 709 -191 857 -190
rect 912 -191 920 -190
rect 954 -191 1165 -190
rect 1171 -191 1266 -190
rect 177 -193 437 -192
rect 520 -193 948 -192
rect 968 -193 1116 -192
rect 1174 -193 1242 -192
rect 58 -195 437 -194
rect 527 -195 1053 -194
rect 1094 -195 1522 -194
rect 58 -197 160 -196
rect 184 -197 297 -196
rect 310 -197 486 -196
rect 506 -197 528 -196
rect 534 -197 717 -196
rect 758 -197 787 -196
rect 793 -197 962 -196
rect 1017 -197 1151 -196
rect 1178 -197 1354 -196
rect 170 -199 311 -198
rect 317 -199 374 -198
rect 394 -199 507 -198
rect 555 -199 780 -198
rect 821 -199 871 -198
rect 1038 -199 1053 -198
rect 1094 -199 1144 -198
rect 1185 -199 1410 -198
rect 184 -201 461 -200
rect 674 -201 969 -200
rect 1038 -201 1550 -200
rect 194 -203 934 -202
rect 1101 -203 1417 -202
rect 198 -205 423 -204
rect 660 -205 675 -204
rect 688 -205 955 -204
rect 1066 -205 1102 -204
rect 1143 -205 1270 -204
rect 30 -207 199 -206
rect 212 -207 822 -206
rect 898 -207 1186 -206
rect 1192 -207 1529 -206
rect 219 -209 318 -208
rect 324 -209 395 -208
rect 401 -209 640 -208
rect 698 -209 1193 -208
rect 1199 -209 1487 -208
rect 219 -211 500 -210
rect 548 -211 661 -210
rect 709 -211 1235 -210
rect 1241 -211 1298 -210
rect 247 -213 1000 -212
rect 1031 -213 1067 -212
rect 1157 -213 1235 -212
rect 1255 -213 1298 -212
rect 89 -215 248 -214
rect 324 -215 1263 -214
rect 1269 -215 1613 -214
rect 352 -217 381 -216
rect 499 -217 752 -216
rect 758 -217 1088 -216
rect 1199 -217 1382 -216
rect 352 -219 524 -218
rect 548 -219 916 -218
rect 996 -219 1088 -218
rect 1202 -219 1340 -218
rect 523 -221 843 -220
rect 863 -221 1032 -220
rect 1045 -221 1158 -220
rect 1206 -221 1480 -220
rect 583 -223 752 -222
rect 765 -223 1179 -222
rect 1213 -223 1312 -222
rect 576 -225 584 -224
rect 604 -225 689 -224
rect 702 -225 864 -224
rect 891 -225 1263 -224
rect 303 -227 605 -226
rect 632 -227 843 -226
rect 982 -227 1046 -226
rect 1216 -227 1319 -226
rect 205 -229 304 -228
rect 576 -229 734 -228
rect 744 -229 794 -228
rect 807 -229 899 -228
rect 936 -229 983 -228
rect 1003 -229 1214 -228
rect 1220 -229 1536 -228
rect 439 -231 1221 -230
rect 1255 -231 1329 -230
rect 625 -233 633 -232
rect 639 -233 713 -232
rect 779 -233 1147 -232
rect 191 -235 626 -234
rect 653 -235 745 -234
rect 807 -235 885 -234
rect 135 -237 654 -236
rect 835 -237 1207 -236
rect 800 -239 836 -238
rect 800 -241 829 -240
rect 723 -243 829 -242
rect 534 -245 724 -244
rect 16 -256 195 -255
rect 198 -256 339 -255
rect 366 -256 748 -255
rect 761 -256 916 -255
rect 992 -256 1599 -255
rect 1612 -256 1970 -255
rect 16 -258 150 -257
rect 156 -258 538 -257
rect 618 -258 801 -257
rect 810 -258 1802 -257
rect 1815 -258 1928 -257
rect 1941 -258 1984 -257
rect 44 -260 209 -259
rect 240 -260 314 -259
rect 338 -260 409 -259
rect 432 -260 797 -259
rect 828 -260 846 -259
rect 880 -260 1529 -259
rect 1542 -260 1606 -259
rect 1615 -260 1662 -259
rect 1668 -260 1732 -259
rect 1962 -260 2194 -259
rect 23 -262 241 -261
rect 247 -262 437 -261
rect 439 -262 591 -261
rect 653 -262 885 -261
rect 891 -262 1641 -261
rect 23 -264 38 -263
rect 54 -264 1508 -263
rect 1514 -264 1844 -263
rect 37 -266 416 -265
rect 422 -266 591 -265
rect 709 -266 1032 -265
rect 1083 -266 1690 -265
rect 65 -268 129 -267
rect 149 -268 171 -267
rect 187 -268 255 -267
rect 268 -268 304 -267
rect 310 -268 983 -267
rect 996 -268 1830 -267
rect 86 -270 94 -269
rect 114 -270 143 -269
rect 156 -270 633 -269
rect 709 -270 815 -269
rect 828 -270 850 -269
rect 856 -270 997 -269
rect 1010 -270 1781 -269
rect 58 -272 143 -271
rect 233 -272 409 -271
rect 422 -272 458 -271
rect 506 -272 521 -271
rect 534 -272 941 -271
rect 954 -272 1032 -271
rect 1094 -272 1550 -271
rect 1552 -272 1767 -271
rect 58 -274 745 -273
rect 772 -274 815 -273
rect 856 -274 990 -273
rect 1010 -274 1018 -273
rect 1020 -274 1452 -273
rect 1465 -274 1795 -273
rect 93 -276 101 -275
rect 128 -276 262 -275
rect 268 -276 472 -275
rect 506 -276 780 -275
rect 863 -276 941 -275
rect 954 -276 1004 -275
rect 1101 -276 1200 -275
rect 1227 -276 1648 -275
rect 100 -278 178 -277
rect 205 -278 780 -277
rect 842 -278 864 -277
rect 894 -278 1536 -277
rect 1556 -278 1655 -277
rect 72 -280 178 -279
rect 191 -280 206 -279
rect 219 -280 535 -279
rect 555 -280 619 -279
rect 628 -280 1004 -279
rect 1153 -280 1711 -279
rect 72 -282 836 -281
rect 926 -282 1095 -281
rect 1178 -282 1515 -281
rect 1591 -282 1816 -281
rect 107 -284 262 -283
rect 275 -284 465 -283
rect 471 -284 486 -283
rect 513 -284 654 -283
rect 667 -284 850 -283
rect 947 -284 1228 -283
rect 1262 -284 1753 -283
rect 107 -286 213 -285
rect 219 -286 227 -285
rect 233 -286 895 -285
rect 947 -286 1546 -285
rect 1626 -286 1718 -285
rect 135 -288 304 -287
rect 310 -288 451 -287
rect 548 -288 556 -287
rect 569 -288 927 -287
rect 968 -288 983 -287
rect 1213 -288 1536 -287
rect 1633 -288 1746 -287
rect 30 -290 451 -289
rect 548 -290 913 -289
rect 1122 -290 1214 -289
rect 1276 -290 1508 -289
rect 30 -292 52 -291
rect 138 -292 171 -291
rect 226 -292 353 -291
rect 394 -292 458 -291
rect 611 -292 969 -291
rect 975 -292 1123 -291
rect 1136 -292 1277 -291
rect 1297 -292 1529 -291
rect 47 -294 52 -293
rect 138 -294 367 -293
rect 394 -294 482 -293
rect 611 -294 682 -293
rect 702 -294 1263 -293
rect 1318 -294 1557 -293
rect 89 -296 682 -295
rect 688 -296 703 -295
rect 723 -296 913 -295
rect 919 -296 1319 -295
rect 1328 -296 2005 -295
rect 243 -298 416 -297
rect 429 -298 465 -297
rect 576 -298 920 -297
rect 1108 -298 1298 -297
rect 1353 -298 1627 -297
rect 247 -300 405 -299
rect 576 -300 839 -299
rect 1024 -300 1109 -299
rect 1360 -300 1739 -299
rect 254 -302 272 -301
rect 275 -302 325 -301
rect 345 -302 570 -301
rect 597 -302 689 -301
rect 723 -302 759 -301
rect 772 -302 1592 -301
rect 282 -304 437 -303
rect 660 -304 668 -303
rect 730 -304 843 -303
rect 1171 -304 1361 -303
rect 1374 -304 1823 -303
rect 135 -306 283 -305
rect 289 -306 486 -305
rect 660 -306 1326 -305
rect 1381 -306 1466 -305
rect 1472 -306 1788 -305
rect 289 -308 388 -307
rect 401 -308 514 -307
rect 716 -308 731 -307
rect 786 -308 1137 -307
rect 1185 -308 1375 -307
rect 1388 -308 1620 -307
rect 296 -310 500 -309
rect 646 -310 717 -309
rect 786 -310 1028 -309
rect 1073 -310 1172 -309
rect 1185 -310 1333 -309
rect 1395 -310 1683 -309
rect 212 -312 647 -311
rect 1073 -312 1270 -311
rect 1402 -312 1669 -311
rect 299 -314 808 -313
rect 1076 -314 1396 -313
rect 1409 -314 1676 -313
rect 324 -316 542 -315
rect 1157 -316 1270 -315
rect 1311 -316 1403 -315
rect 1416 -316 1697 -315
rect 331 -318 500 -317
rect 933 -318 1417 -317
rect 1423 -318 1760 -317
rect 331 -320 801 -319
rect 870 -320 934 -319
rect 1104 -320 1312 -319
rect 1430 -320 1725 -319
rect 345 -322 528 -321
rect 632 -322 871 -321
rect 1157 -322 1256 -321
rect 1437 -322 1704 -321
rect 79 -324 528 -323
rect 712 -324 1256 -323
rect 1444 -324 1774 -323
rect 79 -326 164 -325
rect 352 -326 622 -325
rect 1164 -326 1333 -325
rect 1451 -326 1613 -325
rect 163 -328 167 -327
rect 359 -328 598 -327
rect 1017 -328 1165 -327
rect 1192 -328 1389 -327
rect 1472 -328 1585 -327
rect 359 -330 524 -329
rect 1066 -330 1193 -329
rect 1206 -330 1424 -329
rect 1486 -330 1837 -329
rect 117 -332 1067 -331
rect 1087 -332 1207 -331
rect 1220 -332 1431 -331
rect 1493 -332 1634 -331
rect 380 -334 388 -333
rect 443 -334 542 -333
rect 961 -334 1088 -333
rect 1234 -334 1410 -333
rect 1500 -334 1809 -333
rect 373 -336 381 -335
rect 443 -336 479 -335
rect 765 -336 962 -335
rect 1038 -336 1221 -335
rect 1248 -336 1438 -335
rect 1479 -336 1501 -335
rect 1563 -336 1585 -335
rect 373 -338 706 -337
rect 1038 -338 1151 -337
rect 1248 -338 1578 -337
rect 478 -340 1543 -339
rect 639 -342 766 -341
rect 1129 -342 1235 -341
rect 1283 -342 1494 -341
rect 639 -344 696 -343
rect 1045 -344 1284 -343
rect 1290 -344 1445 -343
rect 695 -346 738 -345
rect 877 -346 1046 -345
rect 1052 -346 1130 -345
rect 1150 -346 1571 -345
rect 604 -348 738 -347
rect 877 -348 1382 -347
rect 1458 -348 1571 -347
rect 317 -350 605 -349
rect 625 -350 1459 -349
rect 121 -352 318 -351
rect 401 -352 626 -351
rect 898 -352 1053 -351
rect 1304 -352 1480 -351
rect 121 -354 584 -353
rect 898 -354 1144 -353
rect 1339 -354 1564 -353
rect 492 -356 584 -355
rect 1024 -356 1291 -355
rect 1346 -356 1578 -355
rect 492 -358 563 -357
rect 821 -358 1347 -357
rect 1367 -358 1487 -357
rect 184 -360 563 -359
rect 751 -360 822 -359
rect 1059 -360 1144 -359
rect 1181 -360 1368 -359
rect 674 -362 752 -361
rect 905 -362 1060 -361
rect 1115 -362 1305 -361
rect 467 -364 675 -363
rect 793 -364 906 -363
rect 1080 -364 1116 -363
rect 1241 -364 1340 -363
rect 793 -366 1522 -365
rect 835 -368 1522 -367
rect 887 -370 1242 -369
rect 16 -381 622 -380
rect 625 -381 703 -380
rect 758 -381 1298 -380
rect 1353 -381 1949 -380
rect 1958 -381 2117 -380
rect 2193 -381 2285 -380
rect 23 -383 748 -382
rect 751 -383 759 -382
rect 761 -383 801 -382
rect 810 -383 829 -382
rect 845 -383 1753 -382
rect 1766 -383 1963 -382
rect 1969 -383 2089 -382
rect 23 -385 45 -384
rect 51 -385 80 -384
rect 96 -385 1179 -384
rect 1185 -385 1298 -384
rect 1353 -385 1473 -384
rect 1591 -385 1753 -384
rect 1773 -385 1900 -384
rect 1927 -385 1998 -384
rect 2004 -385 2264 -384
rect 37 -387 482 -386
rect 495 -387 563 -386
rect 600 -387 1137 -386
rect 1167 -387 1683 -386
rect 1710 -387 1851 -386
rect 1976 -387 1991 -386
rect 2011 -387 2145 -386
rect 44 -389 447 -388
rect 478 -389 857 -388
rect 971 -389 1760 -388
rect 1794 -389 1907 -388
rect 1983 -389 2040 -388
rect 61 -391 248 -390
rect 345 -391 479 -390
rect 513 -391 563 -390
rect 625 -391 885 -390
rect 978 -391 1347 -390
rect 1356 -391 1431 -390
rect 1440 -391 1984 -390
rect 72 -393 136 -392
rect 163 -393 1802 -392
rect 1808 -393 1914 -392
rect 16 -395 164 -394
rect 170 -395 216 -394
rect 222 -395 591 -394
rect 635 -395 1592 -394
rect 1612 -395 1942 -394
rect 72 -397 87 -396
rect 173 -397 206 -396
rect 233 -397 752 -396
rect 765 -397 892 -396
rect 978 -397 1088 -396
rect 1125 -397 1858 -396
rect 30 -399 234 -398
rect 247 -399 374 -398
rect 401 -399 507 -398
rect 513 -399 689 -398
rect 702 -399 1007 -398
rect 1017 -399 1781 -398
rect 1815 -399 1921 -398
rect 79 -401 612 -400
rect 646 -401 913 -400
rect 982 -401 1105 -400
rect 1136 -401 1249 -400
rect 1262 -401 1347 -400
rect 1360 -401 1431 -400
rect 1493 -401 1613 -400
rect 1633 -401 1760 -400
rect 1787 -401 1816 -400
rect 1836 -401 1935 -400
rect 86 -403 416 -402
rect 443 -403 507 -402
rect 527 -403 983 -402
rect 1020 -403 1326 -402
rect 1360 -403 1543 -402
rect 1549 -403 1634 -402
rect 1654 -403 1865 -402
rect 121 -405 206 -404
rect 212 -405 444 -404
rect 527 -405 549 -404
rect 667 -405 773 -404
rect 793 -405 1739 -404
rect 1745 -405 1893 -404
rect 114 -407 122 -406
rect 156 -407 766 -406
rect 849 -407 892 -406
rect 1024 -407 1774 -406
rect 1843 -407 1970 -406
rect 156 -409 192 -408
rect 219 -409 668 -408
rect 674 -409 829 -408
rect 852 -409 1123 -408
rect 1129 -409 1249 -408
rect 1388 -409 1473 -408
rect 1500 -409 1844 -408
rect 149 -411 192 -410
rect 226 -411 612 -410
rect 674 -411 710 -410
rect 716 -411 773 -410
rect 856 -411 986 -410
rect 1027 -411 1963 -410
rect 149 -413 433 -412
rect 541 -413 591 -412
rect 653 -413 710 -412
rect 730 -413 794 -412
rect 863 -413 913 -412
rect 1031 -413 1088 -412
rect 1164 -413 1543 -412
rect 1563 -413 1655 -412
rect 1661 -413 1781 -412
rect 187 -415 1767 -414
rect 226 -417 241 -416
rect 345 -417 465 -416
rect 541 -417 650 -416
rect 653 -417 1480 -416
rect 1507 -417 1550 -416
rect 1570 -417 1802 -416
rect 240 -419 269 -418
rect 359 -419 430 -418
rect 548 -419 570 -418
rect 681 -419 1018 -418
rect 1059 -419 1130 -418
rect 1178 -419 1291 -418
rect 1311 -419 1389 -418
rect 1402 -419 1494 -418
rect 1584 -419 1711 -418
rect 1724 -419 1879 -418
rect 166 -421 360 -420
rect 373 -421 437 -420
rect 471 -421 682 -420
rect 688 -421 958 -420
rect 968 -421 1032 -420
rect 1073 -421 1872 -420
rect 100 -423 437 -422
rect 457 -423 472 -422
rect 730 -423 808 -422
rect 1076 -423 1648 -422
rect 1668 -423 1788 -422
rect 100 -425 521 -424
rect 744 -425 1263 -424
rect 1328 -425 1669 -424
rect 1675 -425 1795 -424
rect 166 -427 332 -426
rect 401 -427 486 -426
rect 737 -427 745 -426
rect 779 -427 1074 -426
rect 1080 -427 1228 -426
rect 1332 -427 1403 -426
rect 1409 -427 1501 -426
rect 1556 -427 1676 -426
rect 1682 -427 1830 -426
rect 212 -429 1060 -428
rect 1083 -429 1662 -428
rect 1689 -429 1809 -428
rect 268 -431 906 -430
rect 968 -431 1648 -430
rect 1703 -431 1837 -430
rect 296 -433 780 -432
rect 803 -433 1333 -432
rect 1367 -433 1480 -432
rect 1486 -433 1585 -432
rect 1619 -433 1739 -432
rect 296 -435 787 -434
rect 807 -435 1123 -434
rect 1192 -435 1291 -434
rect 1437 -435 1508 -434
rect 1514 -435 1620 -434
rect 1626 -435 1746 -434
rect 303 -437 486 -436
rect 632 -437 787 -436
rect 842 -437 1410 -436
rect 1423 -437 1515 -436
rect 1521 -437 1627 -436
rect 1640 -437 1725 -436
rect 1731 -437 1886 -436
rect 177 -439 304 -438
rect 310 -439 570 -438
rect 632 -439 878 -438
rect 887 -439 1641 -438
rect 1717 -439 1830 -438
rect 177 -441 339 -440
rect 408 -441 521 -440
rect 719 -441 1424 -440
rect 1444 -441 1522 -440
rect 1577 -441 1690 -440
rect 107 -443 409 -442
rect 415 -443 640 -442
rect 775 -443 1445 -442
rect 1451 -443 1578 -442
rect 1598 -443 1718 -442
rect 107 -445 276 -444
rect 310 -445 367 -444
rect 429 -445 619 -444
rect 814 -445 843 -444
rect 870 -445 1228 -444
rect 1241 -445 1557 -444
rect 1605 -445 1732 -444
rect 2 -447 619 -446
rect 821 -447 878 -446
rect 905 -447 941 -446
rect 1010 -447 1242 -446
rect 1255 -447 1452 -446
rect 1458 -447 1606 -446
rect 58 -449 815 -448
rect 870 -449 1081 -448
rect 1083 -449 1396 -448
rect 1465 -449 1571 -448
rect 128 -451 367 -450
rect 450 -451 1704 -450
rect 128 -453 143 -452
rect 198 -453 640 -452
rect 695 -453 822 -452
rect 940 -453 1151 -452
rect 1181 -453 1459 -452
rect 1486 -453 1823 -452
rect 142 -455 927 -454
rect 1010 -455 1039 -454
rect 1066 -455 1193 -454
rect 1220 -455 1312 -454
rect 1318 -455 1466 -454
rect 1696 -455 1823 -454
rect 184 -457 696 -456
rect 726 -457 1256 -456
rect 1269 -457 1396 -456
rect 1535 -457 1697 -456
rect 184 -459 577 -458
rect 1038 -459 1053 -458
rect 1066 -459 1956 -458
rect 198 -461 353 -460
rect 450 -461 724 -460
rect 898 -461 1053 -460
rect 1101 -461 1599 -460
rect 219 -463 927 -462
rect 1045 -463 1102 -462
rect 1108 -463 1151 -462
rect 1199 -463 1270 -462
rect 1283 -463 1368 -462
rect 1416 -463 1536 -462
rect 275 -465 388 -464
rect 576 -465 605 -464
rect 723 -465 1375 -464
rect 289 -467 388 -466
rect 583 -467 605 -466
rect 849 -467 1284 -466
rect 1339 -467 1417 -466
rect 282 -469 290 -468
rect 317 -469 458 -468
rect 583 -469 797 -468
rect 898 -469 955 -468
rect 961 -469 1109 -468
rect 1115 -469 1221 -468
rect 1276 -469 1340 -468
rect 1374 -469 1382 -468
rect 254 -471 283 -470
rect 317 -471 717 -470
rect 740 -471 1116 -470
rect 1171 -471 1200 -470
rect 1206 -471 1319 -470
rect 254 -473 598 -472
rect 863 -473 955 -472
rect 992 -473 1172 -472
rect 1213 -473 1277 -472
rect 1304 -473 1382 -472
rect 324 -475 738 -474
rect 919 -475 1046 -474
rect 1143 -475 1207 -474
rect 1234 -475 1305 -474
rect 324 -477 423 -476
rect 464 -477 598 -476
rect 919 -477 990 -476
rect 1094 -477 1144 -476
rect 1157 -477 1235 -476
rect 331 -479 381 -478
rect 422 -479 535 -478
rect 947 -479 962 -478
rect 975 -479 1214 -478
rect 93 -481 381 -480
rect 933 -481 948 -480
rect 989 -481 1928 -480
rect 93 -483 535 -482
rect 933 -483 1564 -482
rect 338 -485 395 -484
rect 996 -485 1095 -484
rect 261 -487 395 -486
rect 835 -487 997 -486
rect 1003 -487 1158 -486
rect 261 -489 661 -488
rect 54 -491 661 -490
rect 352 -493 1028 -492
rect 555 -495 836 -494
rect 492 -497 556 -496
rect 492 -499 1186 -498
rect 30 -510 73 -509
rect 93 -510 174 -509
rect 205 -510 734 -509
rect 737 -510 1634 -509
rect 1682 -510 2152 -509
rect 2214 -510 2292 -509
rect 37 -512 647 -511
rect 656 -512 696 -511
rect 723 -512 773 -511
rect 824 -512 1130 -511
rect 1146 -512 1375 -511
rect 1535 -512 2033 -511
rect 2039 -512 2173 -511
rect 2263 -512 2362 -511
rect 44 -514 213 -513
rect 215 -514 1767 -513
rect 1836 -514 2005 -513
rect 2014 -514 2180 -513
rect 2284 -514 2327 -513
rect 44 -516 167 -515
rect 170 -516 451 -515
rect 541 -516 633 -515
rect 635 -516 773 -515
rect 842 -516 885 -515
rect 898 -516 969 -515
rect 982 -516 1753 -515
rect 1864 -516 2047 -515
rect 2088 -516 2211 -515
rect 135 -518 738 -517
rect 751 -518 755 -517
rect 786 -518 843 -517
rect 849 -518 920 -517
rect 975 -518 1753 -517
rect 1864 -518 1980 -517
rect 1983 -518 2159 -517
rect 75 -520 920 -519
rect 985 -520 1767 -519
rect 1794 -520 1984 -519
rect 1990 -520 2008 -519
rect 2116 -520 2194 -519
rect 114 -522 976 -521
rect 992 -522 1214 -521
rect 1269 -522 1375 -521
rect 1472 -522 1536 -521
rect 1612 -522 1795 -521
rect 1808 -522 1991 -521
rect 2116 -522 2225 -521
rect 114 -524 332 -523
rect 380 -524 990 -523
rect 996 -524 1126 -523
rect 1164 -524 2138 -523
rect 2144 -524 2201 -523
rect 138 -526 899 -525
rect 940 -526 997 -525
rect 1003 -526 1844 -525
rect 1871 -526 2054 -525
rect 163 -528 717 -527
rect 723 -528 1109 -527
rect 1167 -528 1361 -527
rect 1395 -528 1473 -527
rect 1619 -528 1809 -527
rect 1878 -528 2061 -527
rect 205 -530 1263 -529
rect 1290 -530 1396 -529
rect 1479 -530 1620 -529
rect 1633 -530 2208 -529
rect 219 -532 2082 -531
rect 219 -534 654 -533
rect 660 -534 1007 -533
rect 1017 -534 1109 -533
rect 1192 -534 1270 -533
rect 1290 -534 1368 -533
rect 1479 -534 2022 -533
rect 79 -536 654 -535
rect 702 -536 1004 -535
rect 1024 -536 1347 -535
rect 1367 -536 1487 -535
rect 1640 -536 1837 -535
rect 1885 -536 2068 -535
rect 222 -538 283 -537
rect 310 -538 664 -537
rect 716 -538 727 -537
rect 730 -538 990 -537
rect 1031 -538 1123 -537
rect 1136 -538 1193 -537
rect 1227 -538 1347 -537
rect 1493 -538 1641 -537
rect 1661 -538 2040 -537
rect 103 -540 1494 -539
rect 1710 -540 1872 -539
rect 1899 -540 2075 -539
rect 226 -542 237 -541
rect 240 -542 311 -541
rect 324 -542 493 -541
rect 534 -542 1214 -541
rect 1255 -542 1361 -541
rect 1717 -542 1879 -541
rect 1906 -542 2110 -541
rect 65 -544 227 -543
rect 233 -544 1718 -543
rect 1731 -544 2103 -543
rect 9 -546 66 -545
rect 72 -546 241 -545
rect 254 -546 598 -545
rect 600 -546 1438 -545
rect 1570 -546 1732 -545
rect 1738 -546 1900 -545
rect 1913 -546 2131 -545
rect 9 -548 199 -547
rect 233 -548 430 -547
rect 450 -548 514 -547
rect 541 -548 741 -547
rect 751 -548 906 -547
rect 947 -548 1018 -547
rect 1034 -548 1935 -547
rect 1941 -548 2096 -547
rect 107 -550 199 -549
rect 282 -550 388 -549
rect 394 -550 1014 -549
rect 1062 -550 2026 -549
rect 16 -552 108 -551
rect 177 -552 255 -551
rect 317 -552 325 -551
rect 331 -552 538 -551
rect 565 -552 1242 -551
rect 1262 -552 1956 -551
rect 1962 -552 2124 -551
rect 16 -554 157 -553
rect 177 -554 888 -553
rect 891 -554 969 -553
rect 978 -554 1739 -553
rect 1759 -554 1942 -553
rect 1948 -554 2166 -553
rect 93 -556 538 -555
rect 569 -556 594 -555
rect 611 -556 703 -555
rect 786 -556 1613 -555
rect 1675 -556 1907 -555
rect 1920 -556 1956 -555
rect 1969 -556 2145 -555
rect 121 -558 157 -557
rect 303 -558 318 -557
rect 345 -558 430 -557
rect 492 -558 563 -557
rect 569 -558 745 -557
rect 835 -558 892 -557
rect 905 -558 962 -557
rect 1031 -558 1242 -557
rect 1283 -558 1571 -557
rect 1591 -558 1760 -557
rect 1773 -558 1949 -557
rect 1976 -558 1998 -557
rect 121 -560 549 -559
rect 604 -560 612 -559
rect 621 -560 871 -559
rect 877 -560 1228 -559
rect 1297 -560 1592 -559
rect 1696 -560 1935 -559
rect 100 -562 549 -561
rect 649 -562 1844 -561
rect 1927 -562 2089 -561
rect 100 -564 640 -563
rect 688 -564 731 -563
rect 754 -564 962 -563
rect 985 -564 1697 -563
rect 1703 -564 1928 -563
rect 61 -566 689 -565
rect 793 -566 871 -565
rect 1073 -566 1130 -565
rect 1150 -566 1256 -565
rect 1297 -566 1802 -565
rect 1829 -566 1886 -565
rect 2 -568 62 -567
rect 303 -568 528 -567
rect 639 -568 710 -567
rect 793 -568 829 -567
rect 852 -568 1039 -567
rect 1080 -568 1711 -567
rect 1724 -568 1963 -567
rect 250 -570 1039 -569
rect 1083 -570 1788 -569
rect 338 -572 346 -571
rect 366 -572 381 -571
rect 387 -572 433 -571
rect 436 -572 605 -571
rect 709 -572 759 -571
rect 765 -572 829 -571
rect 863 -572 948 -571
rect 971 -572 1725 -571
rect 1745 -572 1921 -571
rect 142 -574 766 -573
rect 821 -574 836 -573
rect 863 -574 1648 -573
rect 1703 -574 1823 -573
rect 142 -576 402 -575
rect 408 -576 514 -575
rect 527 -576 556 -575
rect 695 -576 822 -575
rect 954 -576 1746 -575
rect 1780 -576 1970 -575
rect 117 -578 402 -577
rect 415 -578 811 -577
rect 856 -578 955 -577
rect 1010 -578 1074 -577
rect 1094 -578 1165 -577
rect 1216 -578 1998 -577
rect 275 -580 409 -579
rect 422 -580 437 -579
rect 495 -580 745 -579
rect 758 -580 780 -579
rect 800 -580 857 -579
rect 1010 -580 1977 -579
rect 86 -582 801 -581
rect 1094 -582 1683 -581
rect 86 -584 353 -583
rect 359 -584 423 -583
rect 506 -584 563 -583
rect 586 -584 1781 -583
rect 58 -586 353 -585
rect 359 -586 479 -585
rect 555 -586 682 -585
rect 1101 -586 1137 -585
rect 1220 -586 1284 -585
rect 1325 -586 1662 -585
rect 23 -588 1326 -587
rect 1332 -588 2012 -587
rect 23 -590 52 -589
rect 275 -590 458 -589
rect 471 -590 507 -589
rect 674 -590 780 -589
rect 1080 -590 1102 -589
rect 1199 -590 1221 -589
rect 1234 -590 1333 -589
rect 1353 -590 1438 -589
rect 1465 -590 1914 -589
rect 51 -592 626 -591
rect 667 -592 675 -591
rect 681 -592 1151 -591
rect 1248 -592 1354 -591
rect 1416 -592 1774 -591
rect 1850 -592 2012 -591
rect 135 -594 458 -593
rect 464 -594 626 -593
rect 1157 -594 1249 -593
rect 1318 -594 1466 -593
rect 1500 -594 1648 -593
rect 184 -596 465 -595
rect 576 -596 668 -595
rect 1087 -596 1158 -595
rect 1311 -596 1319 -595
rect 1402 -596 1501 -595
rect 1521 -596 1676 -595
rect 184 -598 262 -597
rect 289 -598 472 -597
rect 576 -598 591 -597
rect 618 -598 1235 -597
rect 1304 -598 1403 -597
rect 1416 -598 2019 -597
rect 149 -600 262 -599
rect 289 -600 934 -599
rect 1206 -600 1312 -599
rect 1430 -600 1522 -599
rect 1528 -600 1830 -599
rect 1857 -600 2019 -599
rect 149 -602 248 -601
rect 338 -602 941 -601
rect 1115 -602 1207 -601
rect 1440 -602 1851 -601
rect 79 -604 248 -603
rect 366 -604 850 -603
rect 912 -604 1305 -603
rect 1528 -604 1578 -603
rect 1598 -604 1788 -603
rect 373 -606 479 -605
rect 590 -606 878 -605
rect 929 -606 1088 -605
rect 1178 -606 1431 -605
rect 1458 -606 1599 -605
rect 1605 -606 1823 -605
rect 191 -608 374 -607
rect 394 -608 500 -607
rect 807 -608 913 -607
rect 933 -608 937 -607
rect 1045 -608 1116 -607
rect 1143 -608 1179 -607
rect 1388 -608 1459 -607
rect 1507 -608 1578 -607
rect 1668 -608 1858 -607
rect 173 -610 192 -609
rect 443 -610 619 -609
rect 926 -610 1046 -609
rect 1143 -610 1816 -609
rect 443 -612 521 -611
rect 926 -612 1543 -611
rect 1549 -612 1802 -611
rect 485 -614 521 -613
rect 1202 -614 1543 -613
rect 1626 -614 1816 -613
rect 485 -616 584 -615
rect 1276 -616 1389 -615
rect 1423 -616 1606 -615
rect 1668 -616 1690 -615
rect 499 -618 661 -617
rect 1185 -618 1277 -617
rect 1339 -618 1424 -617
rect 1444 -618 1550 -617
rect 1556 -618 1690 -617
rect 583 -620 1655 -619
rect 1059 -622 1186 -621
rect 1381 -622 1445 -621
rect 1451 -622 1627 -621
rect 1059 -624 2187 -623
rect 1066 -626 1452 -625
rect 1507 -626 1515 -625
rect 1556 -626 1564 -625
rect 1584 -626 1655 -625
rect 1052 -628 1067 -627
rect 1171 -628 1340 -627
rect 1409 -628 1515 -627
rect 1563 -628 2222 -627
rect 268 -630 1053 -629
rect 1199 -630 1382 -629
rect 1409 -630 1959 -629
rect 268 -632 416 -631
rect 915 -632 1172 -631
rect 1489 -632 1585 -631
rect 2 -643 122 -642
rect 131 -643 2138 -642
rect 2144 -643 2320 -642
rect 2326 -643 2348 -642
rect 2361 -643 2404 -642
rect 44 -645 1224 -644
rect 1300 -645 2131 -644
rect 2137 -645 2173 -644
rect 2193 -645 2208 -644
rect 2214 -645 2278 -644
rect 2291 -645 2327 -644
rect 47 -647 66 -646
rect 68 -647 755 -646
rect 807 -647 1123 -646
rect 1143 -647 1592 -646
rect 1703 -647 2236 -646
rect 12 -649 66 -648
rect 72 -649 1781 -648
rect 1843 -649 2222 -648
rect 51 -651 927 -650
rect 940 -651 1907 -650
rect 1955 -651 2257 -650
rect 51 -653 682 -652
rect 698 -653 983 -652
rect 1010 -653 2152 -652
rect 2158 -653 2313 -652
rect 58 -655 1683 -654
rect 1885 -655 2131 -654
rect 2200 -655 2225 -654
rect 72 -657 1004 -656
rect 1059 -657 1627 -656
rect 1885 -657 1970 -656
rect 2004 -657 2145 -656
rect 82 -659 1032 -658
rect 1059 -659 1074 -658
rect 1083 -659 1466 -658
rect 1486 -659 2166 -658
rect 16 -661 1074 -660
rect 1094 -661 2187 -660
rect 93 -663 563 -662
rect 618 -663 941 -662
rect 957 -663 1053 -662
rect 1062 -663 2180 -662
rect 93 -665 143 -664
rect 145 -665 944 -664
rect 1052 -665 1109 -664
rect 1150 -665 2187 -664
rect 75 -667 1109 -666
rect 1136 -667 1151 -666
rect 1174 -667 2306 -666
rect 135 -669 1823 -668
rect 1857 -669 2005 -668
rect 2011 -669 2152 -668
rect 170 -671 311 -670
rect 401 -671 1032 -670
rect 1101 -671 1123 -670
rect 1178 -671 1214 -670
rect 1216 -671 2110 -670
rect 2116 -671 2299 -670
rect 173 -673 1928 -672
rect 1983 -673 2110 -672
rect 2123 -673 2292 -672
rect 187 -675 703 -674
rect 733 -675 2180 -674
rect 205 -677 1452 -676
rect 1493 -677 1627 -676
rect 1717 -677 1823 -676
rect 1864 -677 2012 -676
rect 2018 -677 2159 -676
rect 212 -679 748 -678
rect 765 -679 1004 -678
rect 1101 -679 1112 -678
rect 1199 -679 1984 -678
rect 1990 -679 2124 -678
rect 191 -681 213 -680
rect 236 -681 1179 -680
rect 1213 -681 1410 -680
rect 1430 -681 1592 -680
rect 1605 -681 1718 -680
rect 1738 -681 1858 -680
rect 1990 -681 2068 -680
rect 2074 -681 2243 -680
rect 149 -683 192 -682
rect 247 -683 318 -682
rect 366 -683 766 -682
rect 800 -683 808 -682
rect 824 -683 2285 -682
rect 30 -685 318 -684
rect 366 -685 773 -684
rect 849 -685 864 -684
rect 891 -685 927 -684
rect 929 -685 1956 -684
rect 1962 -685 2068 -684
rect 2081 -685 2250 -684
rect 9 -687 864 -686
rect 877 -687 892 -686
rect 1080 -687 1739 -686
rect 1752 -687 2075 -686
rect 2088 -687 2264 -686
rect 19 -689 2082 -688
rect 2095 -689 2271 -688
rect 30 -691 38 -690
rect 149 -691 986 -690
rect 1080 -691 1088 -690
rect 1129 -691 1200 -690
rect 1360 -691 1452 -690
rect 1549 -691 1683 -690
rect 1759 -691 2096 -690
rect 37 -693 724 -692
rect 730 -693 1494 -692
rect 1556 -693 1970 -692
rect 1976 -693 2089 -692
rect 261 -695 363 -694
rect 401 -695 556 -694
rect 562 -695 668 -694
rect 681 -695 1711 -694
rect 1794 -695 1928 -694
rect 1997 -695 2117 -694
rect 156 -697 262 -696
rect 282 -697 584 -696
rect 590 -697 668 -696
rect 702 -697 1305 -696
rect 1360 -697 1774 -696
rect 1829 -697 1963 -696
rect 2025 -697 2166 -696
rect 128 -699 157 -698
rect 240 -699 283 -698
rect 310 -699 507 -698
rect 523 -699 1487 -698
rect 1507 -699 1795 -698
rect 1829 -699 1942 -698
rect 2039 -699 2218 -698
rect 114 -701 241 -700
rect 324 -701 507 -700
rect 548 -701 566 -700
rect 569 -701 801 -700
rect 814 -701 850 -700
rect 852 -701 1746 -700
rect 1808 -701 1942 -700
rect 2046 -701 2173 -700
rect 86 -703 115 -702
rect 324 -703 465 -702
rect 492 -703 685 -702
rect 744 -703 2208 -702
rect 5 -705 87 -704
rect 415 -705 465 -704
rect 492 -705 696 -704
rect 747 -705 2103 -704
rect 408 -707 416 -706
rect 429 -707 556 -706
rect 590 -707 1466 -706
rect 1584 -707 1704 -706
rect 1836 -707 1977 -706
rect 2053 -707 2201 -706
rect 303 -709 409 -708
rect 422 -709 430 -708
rect 432 -709 626 -708
rect 639 -709 1781 -708
rect 1850 -709 1998 -708
rect 2060 -709 2194 -708
rect 100 -711 640 -710
rect 646 -711 1228 -710
rect 1248 -711 1760 -710
rect 1871 -711 2026 -710
rect 100 -713 199 -712
rect 219 -713 304 -712
rect 422 -713 1203 -712
rect 1248 -713 1459 -712
rect 1528 -713 1872 -712
rect 1878 -713 2047 -712
rect 163 -715 199 -714
rect 443 -715 549 -714
rect 604 -715 619 -714
rect 653 -715 790 -714
rect 814 -715 871 -714
rect 947 -715 1130 -714
rect 1136 -715 1746 -714
rect 1899 -715 2040 -714
rect 163 -717 486 -716
rect 534 -717 570 -716
rect 576 -717 605 -716
rect 611 -717 626 -716
rect 660 -717 2229 -716
rect 23 -719 486 -718
rect 583 -719 948 -718
rect 996 -719 1088 -718
rect 1097 -719 1529 -718
rect 1598 -719 1711 -718
rect 1724 -719 1837 -718
rect 1920 -719 2061 -718
rect 23 -721 745 -720
rect 772 -721 780 -720
rect 793 -721 871 -720
rect 989 -721 997 -720
rect 1045 -721 1557 -720
rect 1598 -721 1676 -720
rect 1689 -721 1809 -720
rect 1920 -721 1949 -720
rect 289 -723 654 -722
rect 663 -723 710 -722
rect 758 -723 794 -722
rect 1045 -723 1067 -722
rect 1143 -723 2103 -722
rect 184 -725 759 -724
rect 779 -725 1116 -724
rect 1192 -725 1228 -724
rect 1255 -725 1305 -724
rect 1367 -725 1431 -724
rect 1437 -725 1550 -724
rect 1570 -725 1690 -724
rect 1731 -725 1851 -724
rect 1934 -725 2054 -724
rect 184 -727 717 -726
rect 898 -727 1067 -726
rect 1171 -727 1438 -726
rect 1577 -727 1676 -726
rect 1766 -727 1900 -726
rect 177 -729 717 -728
rect 898 -729 1147 -728
rect 1171 -729 1410 -728
rect 1423 -729 1571 -728
rect 1605 -729 1641 -728
rect 1647 -729 1774 -728
rect 1801 -729 1935 -728
rect 58 -731 1147 -730
rect 1234 -731 1256 -730
rect 1290 -731 1585 -730
rect 1612 -731 1725 -730
rect 1815 -731 1949 -730
rect 177 -733 1270 -732
rect 1339 -733 1424 -732
rect 1444 -733 1802 -732
rect 219 -735 1613 -734
rect 1619 -735 1753 -734
rect 250 -737 1193 -736
rect 1206 -737 1270 -736
rect 1353 -737 1445 -736
rect 1472 -737 1620 -736
rect 1633 -737 1732 -736
rect 142 -739 1473 -738
rect 1500 -739 1641 -738
rect 1654 -739 1879 -738
rect 205 -741 1501 -740
rect 1514 -741 1655 -740
rect 1668 -741 2019 -740
rect 289 -743 500 -742
rect 537 -743 990 -742
rect 1024 -743 1578 -742
rect 1696 -743 1816 -742
rect 373 -745 1697 -744
rect 352 -747 374 -746
rect 380 -747 577 -746
rect 611 -747 689 -746
rect 726 -747 1354 -746
rect 1370 -747 1844 -746
rect 254 -749 381 -748
rect 394 -749 535 -748
rect 632 -749 661 -748
rect 674 -749 710 -748
rect 1017 -749 1025 -748
rect 1038 -749 1116 -748
rect 1185 -749 1235 -748
rect 1241 -749 1291 -748
rect 1374 -749 1459 -748
rect 1514 -749 1522 -748
rect 1535 -749 1634 -748
rect 254 -751 521 -750
rect 597 -751 675 -750
rect 688 -751 1165 -750
rect 1185 -751 1564 -750
rect 331 -753 353 -752
rect 387 -753 598 -752
rect 968 -753 1018 -752
rect 1094 -753 1340 -752
rect 1346 -753 1522 -752
rect 1535 -753 1865 -752
rect 275 -755 332 -754
rect 387 -755 479 -754
rect 499 -755 514 -754
rect 933 -755 969 -754
rect 975 -755 1039 -754
rect 1139 -755 1375 -754
rect 1381 -755 1648 -754
rect 275 -757 297 -756
rect 359 -757 479 -756
rect 513 -757 920 -756
rect 954 -757 976 -756
rect 1153 -757 1242 -756
rect 1283 -757 1347 -756
rect 1395 -757 1508 -756
rect 1538 -757 1767 -756
rect 208 -759 920 -758
rect 1157 -759 1165 -758
rect 1206 -759 1221 -758
rect 1311 -759 1382 -758
rect 1395 -759 1403 -758
rect 1542 -759 1669 -758
rect 44 -761 1543 -760
rect 135 -763 209 -762
rect 296 -763 542 -762
rect 786 -763 955 -762
rect 961 -763 1312 -762
rect 1318 -763 1564 -762
rect 345 -765 360 -764
rect 443 -765 528 -764
rect 810 -765 1284 -764
rect 79 -767 528 -766
rect 884 -767 934 -766
rect 1157 -767 2033 -766
rect 79 -769 633 -768
rect 905 -769 962 -768
rect 1209 -769 2033 -768
rect 107 -771 885 -770
rect 1220 -771 2215 -770
rect 107 -773 822 -772
rect 1262 -773 1403 -772
rect 268 -775 906 -774
rect 268 -777 339 -776
rect 345 -777 650 -776
rect 821 -777 836 -776
rect 880 -777 1263 -776
rect 338 -779 752 -778
rect 828 -779 836 -778
rect 450 -781 731 -780
rect 751 -781 1417 -780
rect 128 -783 1417 -782
rect 233 -785 451 -784
rect 457 -785 542 -784
rect 828 -785 1914 -784
rect 233 -787 395 -786
rect 457 -787 843 -786
rect 1787 -787 1914 -786
rect 471 -789 647 -788
rect 842 -789 913 -788
rect 1661 -789 1788 -788
rect 471 -791 1011 -790
rect 1276 -791 1662 -790
rect 520 -793 1319 -792
rect 912 -795 1298 -794
rect 1276 -797 1480 -796
rect 1297 -799 1333 -798
rect 1388 -799 1480 -798
rect 1325 -801 1389 -800
rect 226 -803 1326 -802
rect 1332 -803 1907 -802
rect 226 -805 587 -804
rect 436 -807 587 -806
rect 222 -809 437 -808
rect 9 -820 1627 -819
rect 1661 -820 2362 -819
rect 2403 -820 2418 -819
rect 9 -822 94 -821
rect 103 -822 353 -821
rect 457 -822 591 -821
rect 614 -822 654 -821
rect 674 -822 748 -821
rect 782 -822 850 -821
rect 947 -822 1315 -821
rect 1332 -822 1424 -821
rect 1538 -822 2096 -821
rect 2326 -822 2337 -821
rect 2343 -822 2404 -821
rect 16 -824 192 -823
rect 222 -824 2250 -823
rect 2277 -824 2327 -823
rect 2347 -824 2376 -823
rect 16 -826 1326 -825
rect 1335 -826 1522 -825
rect 1598 -826 1602 -825
rect 1626 -826 1655 -825
rect 1661 -826 1816 -825
rect 2095 -826 2152 -825
rect 2277 -826 2341 -825
rect 2347 -826 2369 -825
rect 44 -828 1697 -827
rect 1815 -828 1879 -827
rect 2151 -828 2180 -827
rect 44 -830 941 -829
rect 947 -830 969 -829
rect 989 -830 1424 -829
rect 1598 -830 1718 -829
rect 1878 -830 1942 -829
rect 1990 -830 2180 -829
rect 58 -832 755 -831
rect 817 -832 1410 -831
rect 1601 -832 1718 -831
rect 1899 -832 1991 -831
rect 58 -834 136 -833
rect 142 -834 223 -833
rect 254 -834 591 -833
rect 635 -834 927 -833
rect 989 -834 1133 -833
rect 1136 -834 1802 -833
rect 1941 -834 1984 -833
rect 79 -836 262 -835
rect 282 -836 363 -835
rect 422 -836 850 -835
rect 870 -836 941 -835
rect 996 -836 1245 -835
rect 1248 -836 1522 -835
rect 1605 -836 1697 -835
rect 1983 -836 2026 -835
rect 72 -838 997 -837
rect 1020 -838 1557 -837
rect 1573 -838 2026 -837
rect 72 -840 668 -839
rect 681 -840 717 -839
rect 821 -840 871 -839
rect 926 -840 1193 -839
rect 1195 -840 2110 -839
rect 79 -842 325 -841
rect 352 -842 500 -841
rect 506 -842 724 -841
rect 772 -842 822 -841
rect 1010 -842 2110 -841
rect 121 -844 269 -843
rect 282 -844 1161 -843
rect 1174 -844 1774 -843
rect 47 -846 1774 -845
rect 128 -848 563 -847
rect 646 -848 832 -847
rect 1010 -848 1088 -847
rect 1094 -848 1123 -847
rect 1129 -848 2236 -847
rect 128 -850 1042 -849
rect 1045 -850 1088 -849
rect 1094 -850 1102 -849
rect 1111 -850 2047 -849
rect 2235 -850 2285 -849
rect 145 -852 801 -851
rect 828 -852 1130 -851
rect 1136 -852 1228 -851
rect 1248 -852 1389 -851
rect 1402 -852 1410 -851
rect 1430 -852 2047 -851
rect 170 -854 192 -853
rect 205 -854 1802 -853
rect 170 -856 272 -855
rect 296 -856 584 -855
rect 646 -856 1256 -855
rect 1272 -856 1970 -855
rect 184 -858 290 -857
rect 310 -858 377 -857
rect 422 -858 1109 -857
rect 1139 -858 1242 -857
rect 1255 -858 1354 -857
rect 1360 -858 2320 -857
rect 184 -860 759 -859
rect 775 -860 1109 -859
rect 1143 -860 2075 -859
rect 198 -862 290 -861
rect 310 -862 451 -861
rect 457 -862 549 -861
rect 562 -862 570 -861
rect 653 -862 1025 -861
rect 1045 -862 1060 -861
rect 1101 -862 1186 -861
rect 1206 -862 1760 -861
rect 1969 -862 2005 -861
rect 2074 -862 2131 -861
rect 156 -864 199 -863
rect 205 -864 234 -863
rect 254 -864 521 -863
rect 527 -864 1207 -863
rect 1209 -864 2124 -863
rect 2130 -864 2166 -863
rect 156 -866 444 -865
rect 478 -866 521 -865
rect 527 -866 808 -865
rect 828 -866 1781 -865
rect 2004 -866 2054 -865
rect 2123 -866 2138 -865
rect 163 -868 451 -867
rect 478 -868 773 -867
rect 807 -868 1081 -867
rect 1143 -868 1217 -867
rect 1220 -868 2061 -867
rect 2102 -868 2138 -867
rect 163 -870 332 -869
rect 359 -870 570 -869
rect 667 -870 2351 -869
rect 187 -872 1781 -871
rect 1787 -872 2061 -871
rect 2102 -872 2159 -871
rect 219 -874 801 -873
rect 957 -874 1403 -873
rect 1556 -874 1648 -873
rect 1654 -874 1746 -873
rect 1787 -874 1830 -873
rect 2053 -874 2089 -873
rect 233 -876 304 -875
rect 324 -876 374 -875
rect 387 -876 444 -875
rect 492 -876 969 -875
rect 1024 -876 1529 -875
rect 1605 -876 1676 -875
rect 1682 -876 1760 -875
rect 1829 -876 1914 -875
rect 100 -878 388 -877
rect 408 -878 549 -877
rect 688 -878 727 -877
rect 737 -878 759 -877
rect 1055 -878 2082 -877
rect 100 -880 937 -879
rect 1080 -880 1165 -879
rect 1185 -880 1767 -879
rect 1871 -880 2089 -879
rect 121 -882 374 -881
rect 408 -882 416 -881
rect 436 -882 507 -881
rect 513 -882 720 -881
rect 723 -882 1032 -881
rect 1146 -882 1518 -881
rect 1647 -882 1739 -881
rect 1745 -882 1844 -881
rect 1913 -882 1963 -881
rect 2081 -882 2145 -881
rect 2 -884 416 -883
rect 492 -884 766 -883
rect 1031 -884 1067 -883
rect 1157 -884 2299 -883
rect 2 -886 178 -885
rect 247 -886 304 -885
rect 359 -886 381 -885
rect 499 -886 531 -885
rect 534 -886 584 -885
rect 688 -886 710 -885
rect 737 -886 885 -885
rect 954 -886 2299 -885
rect 65 -888 1963 -887
rect 2144 -888 2173 -887
rect 65 -890 395 -889
rect 464 -890 535 -889
rect 541 -890 675 -889
rect 698 -890 920 -889
rect 1052 -890 1067 -889
rect 1157 -890 1200 -889
rect 1213 -890 2243 -889
rect 86 -892 395 -891
rect 401 -892 465 -891
rect 513 -892 598 -891
rect 702 -892 1172 -891
rect 1199 -892 1277 -891
rect 1286 -892 1529 -891
rect 1682 -892 1704 -891
rect 1738 -892 1865 -891
rect 2172 -892 2194 -891
rect 2207 -892 2243 -891
rect 86 -894 367 -893
rect 380 -894 612 -893
rect 702 -894 836 -893
rect 905 -894 1053 -893
rect 1125 -894 1865 -893
rect 2193 -894 2229 -893
rect 107 -896 906 -895
rect 919 -896 1116 -895
rect 1164 -896 1270 -895
rect 1290 -896 1389 -895
rect 1395 -896 1431 -895
rect 1766 -896 2313 -895
rect 107 -898 241 -897
rect 247 -898 1018 -897
rect 1038 -898 1116 -897
rect 1171 -898 2201 -897
rect 2207 -898 2264 -897
rect 51 -900 241 -899
rect 261 -900 633 -899
rect 765 -900 815 -899
rect 1192 -900 1277 -899
rect 1290 -900 1347 -899
rect 1353 -900 1585 -899
rect 1794 -900 1872 -899
rect 1892 -900 2264 -899
rect 51 -902 629 -901
rect 639 -902 1893 -901
rect 2018 -902 2313 -901
rect 124 -904 1676 -903
rect 1794 -904 1907 -903
rect 2018 -904 2068 -903
rect 2186 -904 2229 -903
rect 149 -906 437 -905
rect 541 -906 612 -905
rect 618 -906 633 -905
rect 786 -906 836 -905
rect 1213 -906 1270 -905
rect 1304 -906 2355 -905
rect 30 -908 787 -907
rect 796 -908 885 -907
rect 1220 -908 1235 -907
rect 1241 -908 1809 -907
rect 1843 -908 2040 -907
rect 2067 -908 2117 -907
rect 2200 -908 2257 -907
rect 30 -910 178 -909
rect 180 -910 710 -909
rect 716 -910 1809 -909
rect 1906 -910 1956 -909
rect 2039 -910 2292 -909
rect 135 -912 2117 -911
rect 2214 -912 2257 -911
rect 149 -914 1175 -913
rect 1223 -914 1704 -913
rect 1955 -914 1998 -913
rect 2214 -914 2271 -913
rect 226 -916 640 -915
rect 814 -916 1312 -915
rect 1325 -916 1417 -915
rect 1535 -916 2187 -915
rect 2270 -916 2306 -915
rect 226 -918 878 -917
rect 1178 -918 1417 -917
rect 1493 -918 2306 -917
rect 23 -920 878 -919
rect 1122 -920 1179 -919
rect 1227 -920 1263 -919
rect 1304 -920 1445 -919
rect 1493 -920 1550 -919
rect 1584 -920 1634 -919
rect 1997 -920 2033 -919
rect 23 -922 115 -921
rect 268 -922 2292 -921
rect 114 -924 486 -923
rect 593 -924 955 -923
rect 1234 -924 1438 -923
rect 1535 -924 1613 -923
rect 1633 -924 1711 -923
rect 1857 -924 2033 -923
rect 275 -926 297 -925
rect 345 -926 619 -925
rect 1262 -926 1298 -925
rect 1311 -926 2285 -925
rect 275 -928 430 -927
rect 485 -928 556 -927
rect 597 -928 605 -927
rect 684 -928 1298 -927
rect 1339 -928 1445 -927
rect 1549 -928 1564 -927
rect 1612 -928 1620 -927
rect 1710 -928 1823 -927
rect 1857 -928 1886 -927
rect 345 -930 661 -929
rect 1283 -930 1438 -929
rect 1563 -930 1669 -929
rect 1822 -930 1837 -929
rect 1885 -930 1949 -929
rect 19 -932 1837 -931
rect 331 -934 1284 -933
rect 1339 -934 1452 -933
rect 1500 -934 1669 -933
rect 366 -936 1399 -935
rect 1500 -936 1578 -935
rect 1619 -936 1725 -935
rect 401 -938 696 -937
rect 1059 -938 1949 -937
rect 187 -940 696 -939
rect 1318 -940 1452 -939
rect 1577 -940 1900 -939
rect 429 -942 1014 -941
rect 1318 -942 1508 -941
rect 1724 -942 1851 -941
rect 604 -944 843 -943
rect 1346 -944 1396 -943
rect 1507 -944 1592 -943
rect 1850 -944 1928 -943
rect 660 -946 913 -945
rect 1360 -946 1382 -945
rect 1591 -946 1690 -945
rect 1927 -946 1977 -945
rect 744 -948 1690 -947
rect 1976 -948 2012 -947
rect 744 -950 794 -949
rect 842 -950 934 -949
rect 1363 -950 2159 -949
rect 555 -952 934 -951
rect 1367 -952 1753 -951
rect 1920 -952 2012 -951
rect 793 -954 962 -953
rect 1017 -954 1753 -953
rect 856 -956 913 -955
rect 961 -956 983 -955
rect 1367 -956 1459 -955
rect 856 -958 892 -957
rect 982 -958 1004 -957
rect 1370 -958 2166 -957
rect 471 -960 892 -959
rect 1374 -960 1921 -959
rect 471 -962 577 -961
rect 586 -962 1004 -961
rect 1374 -962 1480 -961
rect 576 -964 626 -963
rect 1381 -964 1487 -963
rect 625 -966 2320 -965
rect 1458 -968 1543 -967
rect 1479 -970 1571 -969
rect 1486 -972 1732 -971
rect 1465 -974 1732 -973
rect 1465 -976 1473 -975
rect 1542 -976 1641 -975
rect 1073 -978 1473 -977
rect 1514 -978 1641 -977
rect 779 -980 1074 -979
rect 1514 -980 2250 -979
rect 1570 -982 2222 -981
rect 751 -984 2222 -983
rect 37 -986 752 -985
rect 37 -988 976 -987
rect 975 -990 1151 -989
rect 730 -992 1151 -991
rect 730 -994 864 -993
rect 338 -996 864 -995
rect 338 -998 391 -997
rect 9 -1009 762 -1008
rect 772 -1009 2138 -1008
rect 2284 -1009 2341 -1008
rect 2375 -1009 2432 -1008
rect 9 -1011 59 -1010
rect 93 -1011 2257 -1010
rect 2298 -1011 2376 -1010
rect 2382 -1011 2393 -1010
rect 2403 -1011 2439 -1010
rect 16 -1013 59 -1012
rect 93 -1013 843 -1012
rect 884 -1013 934 -1012
rect 936 -1013 1389 -1012
rect 1507 -1013 1578 -1012
rect 1703 -1013 2299 -1012
rect 2368 -1013 2404 -1012
rect 2417 -1013 2425 -1012
rect 16 -1015 332 -1014
rect 345 -1015 1007 -1014
rect 1020 -1015 2229 -1014
rect 103 -1017 1151 -1016
rect 1174 -1017 1872 -1016
rect 2123 -1017 2369 -1016
rect 110 -1019 318 -1018
rect 324 -1019 332 -1018
rect 345 -1019 444 -1018
rect 590 -1019 629 -1018
rect 646 -1019 955 -1018
rect 964 -1019 2243 -1018
rect 117 -1021 1452 -1020
rect 1514 -1021 1683 -1020
rect 1689 -1021 1704 -1020
rect 1787 -1021 2124 -1020
rect 2165 -1021 2229 -1020
rect 128 -1023 783 -1022
rect 793 -1023 1109 -1022
rect 1122 -1023 1361 -1022
rect 1514 -1023 1536 -1022
rect 1710 -1023 1788 -1022
rect 1801 -1023 2390 -1022
rect 128 -1025 262 -1024
rect 268 -1025 479 -1024
rect 590 -1025 668 -1024
rect 733 -1025 2292 -1024
rect 86 -1027 668 -1026
rect 779 -1027 1991 -1026
rect 2102 -1027 2292 -1026
rect 86 -1029 136 -1028
rect 138 -1029 1893 -1028
rect 1962 -1029 1991 -1028
rect 2172 -1029 2243 -1028
rect 135 -1031 1823 -1030
rect 1836 -1031 1893 -1030
rect 1962 -1031 2019 -1030
rect 2130 -1031 2173 -1030
rect 177 -1033 2320 -1032
rect 23 -1035 178 -1034
rect 180 -1035 465 -1034
rect 478 -1035 486 -1034
rect 611 -1035 2222 -1034
rect 23 -1037 45 -1036
rect 100 -1037 2320 -1036
rect 44 -1039 241 -1038
rect 261 -1039 276 -1038
rect 310 -1039 881 -1038
rect 940 -1039 1018 -1038
rect 1024 -1039 1508 -1038
rect 1517 -1039 2264 -1038
rect 184 -1041 255 -1040
rect 271 -1041 780 -1040
rect 793 -1041 857 -1040
rect 863 -1041 885 -1040
rect 891 -1041 941 -1040
rect 975 -1041 1109 -1040
rect 1125 -1041 2089 -1040
rect 2158 -1041 2222 -1040
rect 138 -1043 2159 -1042
rect 187 -1045 2278 -1044
rect 191 -1047 311 -1046
rect 324 -1047 682 -1046
rect 723 -1047 976 -1046
rect 989 -1047 1039 -1046
rect 1041 -1047 2019 -1046
rect 2067 -1047 2131 -1046
rect 2200 -1047 2278 -1046
rect 170 -1049 192 -1048
rect 205 -1049 318 -1048
rect 366 -1049 612 -1048
rect 625 -1049 1732 -1048
rect 1738 -1049 1823 -1048
rect 1843 -1049 2103 -1048
rect 2200 -1049 2250 -1048
rect 121 -1051 206 -1050
rect 219 -1051 654 -1050
rect 660 -1051 717 -1050
rect 730 -1051 857 -1050
rect 863 -1051 1690 -1050
rect 1710 -1051 2362 -1050
rect 121 -1053 360 -1052
rect 366 -1053 1172 -1052
rect 1181 -1053 1627 -1052
rect 1745 -1053 1802 -1052
rect 1843 -1053 1851 -1052
rect 1864 -1053 2138 -1052
rect 2186 -1053 2250 -1052
rect 145 -1055 731 -1054
rect 796 -1055 913 -1054
rect 996 -1055 1203 -1054
rect 1234 -1055 1389 -1054
rect 1437 -1055 1732 -1054
rect 1815 -1055 1851 -1054
rect 1871 -1055 1907 -1054
rect 1983 -1055 2264 -1054
rect 170 -1057 377 -1056
rect 380 -1057 776 -1056
rect 817 -1057 1669 -1056
rect 1675 -1057 1907 -1056
rect 1955 -1057 1984 -1056
rect 2004 -1057 2068 -1056
rect 2186 -1057 2400 -1056
rect 79 -1059 381 -1058
rect 387 -1059 815 -1058
rect 831 -1059 2033 -1058
rect 2039 -1059 2362 -1058
rect 79 -1061 115 -1060
rect 222 -1061 619 -1060
rect 639 -1061 724 -1060
rect 775 -1061 969 -1060
rect 982 -1061 997 -1060
rect 1003 -1061 1172 -1060
rect 1192 -1061 2047 -1060
rect 30 -1063 619 -1062
rect 646 -1063 710 -1062
rect 835 -1063 1123 -1062
rect 1136 -1063 1151 -1062
rect 1157 -1063 1193 -1062
rect 1234 -1063 1837 -1062
rect 1878 -1063 2166 -1062
rect 30 -1065 720 -1064
rect 835 -1065 948 -1064
rect 968 -1065 1074 -1064
rect 1129 -1065 1158 -1064
rect 1237 -1065 1291 -1064
rect 1307 -1065 2005 -1064
rect 2011 -1065 2089 -1064
rect 65 -1067 640 -1066
rect 660 -1067 759 -1066
rect 842 -1067 871 -1066
rect 877 -1067 913 -1066
rect 947 -1067 2257 -1066
rect 65 -1069 472 -1068
rect 485 -1069 535 -1068
rect 597 -1069 626 -1068
rect 635 -1069 1074 -1068
rect 1087 -1069 1130 -1068
rect 1136 -1069 1473 -1068
rect 1479 -1069 1536 -1068
rect 1542 -1069 1627 -1068
rect 1633 -1069 1676 -1068
rect 1815 -1069 2397 -1068
rect 226 -1071 465 -1070
rect 513 -1071 815 -1070
rect 891 -1071 899 -1070
rect 1003 -1071 1025 -1070
rect 1045 -1071 1088 -1070
rect 1241 -1071 2061 -1070
rect 51 -1073 514 -1072
rect 534 -1073 1270 -1072
rect 1272 -1073 2033 -1072
rect 2039 -1073 2348 -1072
rect 51 -1075 143 -1074
rect 212 -1075 227 -1074
rect 240 -1075 528 -1074
rect 597 -1075 1063 -1074
rect 1223 -1075 1242 -1074
rect 1244 -1075 2285 -1074
rect 142 -1077 990 -1076
rect 1010 -1077 1039 -1076
rect 1055 -1077 1550 -1076
rect 1598 -1077 1669 -1076
rect 1829 -1077 1865 -1076
rect 1878 -1077 1928 -1076
rect 1941 -1077 1956 -1076
rect 1969 -1077 2012 -1076
rect 2207 -1077 2348 -1076
rect 198 -1079 213 -1078
rect 254 -1079 542 -1078
rect 681 -1079 951 -1078
rect 1017 -1079 1116 -1078
rect 1248 -1079 1361 -1078
rect 1374 -1079 1438 -1078
rect 1486 -1079 1830 -1078
rect 1927 -1079 2194 -1078
rect 198 -1081 808 -1080
rect 877 -1081 1270 -1080
rect 1283 -1081 2313 -1080
rect 275 -1083 416 -1082
rect 429 -1083 1448 -1082
rect 1500 -1083 1543 -1082
rect 1580 -1083 1942 -1082
rect 1997 -1083 2047 -1082
rect 2109 -1083 2208 -1082
rect 2235 -1083 2313 -1082
rect 359 -1085 433 -1084
rect 443 -1085 500 -1084
rect 541 -1085 605 -1084
rect 607 -1085 2194 -1084
rect 114 -1087 500 -1086
rect 604 -1087 1046 -1086
rect 1059 -1087 1144 -1086
rect 1227 -1087 1249 -1086
rect 1286 -1087 1760 -1086
rect 1808 -1087 1970 -1086
rect 2151 -1087 2236 -1086
rect 401 -1089 405 -1088
rect 415 -1089 507 -1088
rect 695 -1089 983 -1088
rect 1080 -1089 1144 -1088
rect 1213 -1089 1228 -1088
rect 1314 -1089 1641 -1088
rect 1654 -1089 1746 -1088
rect 1857 -1089 2110 -1088
rect 401 -1091 409 -1090
rect 429 -1091 1774 -1090
rect 1794 -1091 1858 -1090
rect 2095 -1091 2152 -1090
rect 408 -1093 577 -1092
rect 688 -1093 696 -1092
rect 702 -1093 808 -1092
rect 898 -1093 1095 -1092
rect 1101 -1093 1116 -1092
rect 1213 -1093 2344 -1092
rect 2 -1095 689 -1094
rect 709 -1095 927 -1094
rect 1031 -1095 1102 -1094
rect 1318 -1095 1452 -1094
rect 1556 -1095 1641 -1094
rect 1696 -1095 1760 -1094
rect 2025 -1095 2096 -1094
rect 72 -1097 703 -1096
rect 737 -1097 1291 -1096
rect 1325 -1097 1375 -1096
rect 1381 -1097 1473 -1096
rect 1598 -1097 1606 -1096
rect 1717 -1097 1774 -1096
rect 1899 -1097 2026 -1096
rect 37 -1099 73 -1098
rect 89 -1099 1095 -1098
rect 1185 -1099 1697 -1098
rect 1717 -1099 1753 -1098
rect 1899 -1099 2334 -1098
rect 37 -1101 594 -1100
rect 751 -1101 871 -1100
rect 905 -1101 1032 -1100
rect 1066 -1101 1081 -1100
rect 1185 -1101 1200 -1100
rect 1206 -1101 1319 -1100
rect 1335 -1101 2306 -1100
rect 247 -1103 927 -1102
rect 961 -1103 1067 -1102
rect 1178 -1103 1207 -1102
rect 1255 -1103 1326 -1102
rect 1367 -1103 1382 -1102
rect 1395 -1103 1753 -1102
rect 2214 -1103 2306 -1102
rect 163 -1105 248 -1104
rect 373 -1105 1179 -1104
rect 1195 -1105 1557 -1104
rect 1724 -1105 1809 -1104
rect 2116 -1105 2215 -1104
rect 2270 -1105 2334 -1104
rect 163 -1107 339 -1106
rect 352 -1107 374 -1106
rect 390 -1107 738 -1106
rect 772 -1107 1634 -1106
rect 2053 -1107 2117 -1106
rect 233 -1109 962 -1108
rect 1052 -1109 1725 -1108
rect 2053 -1109 2337 -1108
rect 233 -1111 395 -1110
rect 450 -1111 472 -1110
rect 506 -1111 1795 -1110
rect 107 -1113 395 -1112
rect 450 -1113 493 -1112
rect 548 -1113 577 -1112
rect 674 -1113 752 -1112
rect 786 -1113 1011 -1112
rect 1199 -1113 1767 -1112
rect 107 -1115 2327 -1114
rect 338 -1117 521 -1116
rect 569 -1117 1053 -1116
rect 1220 -1117 1256 -1116
rect 1262 -1117 1368 -1116
rect 1402 -1117 2061 -1116
rect 352 -1119 867 -1118
rect 905 -1119 1683 -1118
rect 1766 -1119 1781 -1118
rect 422 -1121 570 -1120
rect 674 -1121 1168 -1120
rect 1220 -1121 2271 -1120
rect 100 -1123 423 -1122
rect 436 -1123 493 -1122
rect 520 -1123 584 -1122
rect 744 -1123 787 -1122
rect 800 -1123 1284 -1122
rect 1297 -1123 1396 -1122
rect 1423 -1123 1480 -1122
rect 1549 -1123 1606 -1122
rect 1661 -1123 1781 -1122
rect 289 -1125 584 -1124
rect 800 -1125 822 -1124
rect 1164 -1125 1263 -1124
rect 1297 -1125 2355 -1124
rect 289 -1127 297 -1126
rect 436 -1127 657 -1126
rect 821 -1127 1998 -1126
rect 296 -1129 304 -1128
rect 457 -1129 549 -1128
rect 555 -1129 745 -1128
rect 1164 -1129 1613 -1128
rect 1619 -1129 1662 -1128
rect 282 -1131 304 -1130
rect 404 -1131 458 -1130
rect 555 -1131 563 -1130
rect 1304 -1131 1403 -1130
rect 1416 -1131 1424 -1130
rect 1430 -1131 1487 -1130
rect 1584 -1131 1613 -1130
rect 149 -1133 283 -1132
rect 1304 -1133 1935 -1132
rect 149 -1135 426 -1134
rect 1311 -1135 2327 -1134
rect 156 -1137 563 -1136
rect 1311 -1137 1340 -1136
rect 1398 -1137 2355 -1136
rect 96 -1139 157 -1138
rect 824 -1139 1340 -1138
rect 1430 -1139 1522 -1138
rect 1528 -1139 1585 -1138
rect 1591 -1139 1620 -1138
rect 1934 -1139 2082 -1138
rect 632 -1141 1592 -1140
rect 2081 -1141 2180 -1140
rect 632 -1143 1161 -1142
rect 1444 -1143 1501 -1142
rect 2144 -1143 2180 -1142
rect 1458 -1145 1522 -1144
rect 2074 -1145 2145 -1144
rect 1276 -1147 1459 -1146
rect 1493 -1147 1529 -1146
rect 1976 -1147 2075 -1146
rect 828 -1149 1277 -1148
rect 1465 -1149 1494 -1148
rect 1948 -1149 1977 -1148
rect 765 -1151 829 -1150
rect 1465 -1151 1648 -1150
rect 1920 -1151 1949 -1150
rect 765 -1153 850 -1152
rect 1563 -1153 1648 -1152
rect 1913 -1153 1921 -1152
rect 849 -1155 1417 -1154
rect 1885 -1155 1914 -1154
rect 1353 -1157 1564 -1156
rect 1741 -1157 1886 -1156
rect 1346 -1159 1354 -1158
rect 1332 -1161 1347 -1160
rect 957 -1163 1333 -1162
rect 957 -1165 1655 -1164
rect 5 -1176 433 -1175
rect 485 -1176 654 -1175
rect 656 -1176 1515 -1175
rect 1549 -1176 2292 -1175
rect 2298 -1176 2495 -1175
rect 19 -1178 31 -1177
rect 89 -1178 857 -1177
rect 866 -1178 1032 -1177
rect 1041 -1178 2474 -1177
rect 23 -1180 822 -1179
rect 842 -1180 857 -1179
rect 880 -1180 1746 -1179
rect 1906 -1180 2453 -1179
rect 23 -1182 612 -1181
rect 667 -1182 850 -1181
rect 905 -1182 927 -1181
rect 947 -1182 1434 -1181
rect 1447 -1182 2362 -1181
rect 2368 -1182 2565 -1181
rect 30 -1184 678 -1183
rect 751 -1184 843 -1183
rect 912 -1184 1032 -1183
rect 1048 -1184 1123 -1183
rect 1157 -1184 2264 -1183
rect 2277 -1184 2467 -1183
rect 100 -1186 909 -1185
rect 947 -1186 1095 -1185
rect 1104 -1186 2544 -1185
rect 100 -1188 248 -1187
rect 254 -1188 913 -1187
rect 950 -1188 1452 -1187
rect 1458 -1188 1550 -1187
rect 1552 -1188 1599 -1187
rect 1605 -1188 1907 -1187
rect 1927 -1188 2460 -1187
rect 121 -1190 510 -1189
rect 513 -1190 612 -1189
rect 667 -1190 1270 -1189
rect 1307 -1190 2397 -1189
rect 2431 -1190 2579 -1189
rect 124 -1192 1291 -1191
rect 1335 -1192 2348 -1191
rect 2354 -1192 2558 -1191
rect 128 -1194 1928 -1193
rect 1969 -1194 2390 -1193
rect 2438 -1194 2481 -1193
rect 128 -1196 269 -1195
rect 275 -1196 783 -1195
rect 796 -1196 969 -1195
rect 982 -1196 1095 -1195
rect 1115 -1196 1270 -1195
rect 1339 -1196 1459 -1195
rect 1500 -1196 1599 -1195
rect 1605 -1196 1613 -1195
rect 1745 -1196 1802 -1195
rect 2060 -1196 2264 -1195
rect 2284 -1196 2488 -1195
rect 138 -1198 584 -1197
rect 590 -1198 1816 -1197
rect 1857 -1198 2061 -1197
rect 2095 -1198 2292 -1197
rect 2305 -1198 2502 -1197
rect 208 -1200 731 -1199
rect 751 -1200 885 -1199
rect 992 -1200 2432 -1199
rect 37 -1202 885 -1201
rect 1003 -1202 1830 -1201
rect 1962 -1202 2285 -1201
rect 2312 -1202 2509 -1201
rect 37 -1204 703 -1203
rect 758 -1204 1515 -1203
rect 1521 -1204 1613 -1203
rect 1668 -1204 1830 -1203
rect 2109 -1204 2299 -1203
rect 2319 -1204 2516 -1203
rect 268 -1206 2376 -1205
rect 2424 -1206 2439 -1205
rect 275 -1208 2344 -1207
rect 310 -1210 969 -1209
rect 1003 -1210 2271 -1209
rect 2333 -1210 2537 -1209
rect 72 -1212 311 -1211
rect 380 -1212 430 -1211
rect 436 -1212 514 -1211
rect 527 -1212 584 -1211
rect 604 -1212 822 -1211
rect 828 -1212 927 -1211
rect 1010 -1212 1116 -1211
rect 1164 -1212 2383 -1211
rect 72 -1214 444 -1213
rect 485 -1214 549 -1213
rect 555 -1214 591 -1213
rect 642 -1214 1858 -1213
rect 1920 -1214 2110 -1213
rect 2116 -1214 2306 -1213
rect 2340 -1214 2551 -1213
rect 9 -1216 556 -1215
rect 569 -1216 654 -1215
rect 702 -1216 958 -1215
rect 1038 -1216 1158 -1215
rect 1167 -1216 2572 -1215
rect 9 -1218 136 -1217
rect 219 -1218 1165 -1217
rect 1178 -1218 1844 -1217
rect 1934 -1218 2320 -1217
rect 16 -1220 444 -1219
rect 499 -1220 731 -1219
rect 758 -1220 787 -1219
rect 800 -1220 895 -1219
rect 1045 -1220 1123 -1219
rect 1185 -1220 1340 -1219
rect 1370 -1220 2103 -1219
rect 2116 -1220 2257 -1219
rect 65 -1222 570 -1221
rect 800 -1222 1039 -1221
rect 1045 -1222 1102 -1221
rect 1192 -1222 1291 -1221
rect 1311 -1222 1501 -1221
rect 1563 -1222 2530 -1221
rect 65 -1224 80 -1223
rect 114 -1224 2103 -1223
rect 2144 -1224 2313 -1223
rect 114 -1226 647 -1225
rect 807 -1226 811 -1225
rect 852 -1226 1802 -1225
rect 1815 -1226 1893 -1225
rect 1948 -1226 2145 -1225
rect 2151 -1226 2334 -1225
rect 135 -1228 682 -1227
rect 789 -1228 1949 -1227
rect 1955 -1228 2152 -1227
rect 2158 -1228 2348 -1227
rect 191 -1230 220 -1229
rect 373 -1230 500 -1229
rect 506 -1230 2446 -1229
rect 191 -1232 388 -1231
rect 408 -1232 608 -1231
rect 646 -1232 1088 -1231
rect 1192 -1232 1263 -1231
rect 1283 -1232 1564 -1231
rect 1570 -1232 1669 -1231
rect 1731 -1232 1893 -1231
rect 1955 -1232 2068 -1231
rect 2088 -1232 2257 -1231
rect 198 -1234 1088 -1233
rect 1234 -1234 2411 -1233
rect 149 -1236 1235 -1235
rect 1255 -1236 1263 -1235
rect 1283 -1236 1354 -1235
rect 1381 -1236 1392 -1235
rect 1416 -1236 1522 -1235
rect 1591 -1236 1732 -1235
rect 1738 -1236 2271 -1235
rect 145 -1238 150 -1237
rect 198 -1238 1361 -1237
rect 1381 -1238 1620 -1237
rect 1633 -1238 1739 -1237
rect 1741 -1238 2068 -1237
rect 2172 -1238 2355 -1237
rect 233 -1240 409 -1239
rect 422 -1240 1795 -1239
rect 1885 -1240 2089 -1239
rect 2179 -1240 2362 -1239
rect 226 -1242 234 -1241
rect 261 -1242 423 -1241
rect 436 -1242 675 -1241
rect 681 -1242 745 -1241
rect 807 -1242 1305 -1241
rect 1332 -1242 1963 -1241
rect 1983 -1242 2159 -1241
rect 2186 -1242 2369 -1241
rect 261 -1244 1011 -1243
rect 1059 -1244 1221 -1243
rect 1241 -1244 1354 -1243
rect 1384 -1244 2208 -1243
rect 2221 -1244 2383 -1243
rect 303 -1246 374 -1245
rect 380 -1246 458 -1245
rect 506 -1246 724 -1245
rect 744 -1246 955 -1245
rect 961 -1246 1634 -1245
rect 1654 -1246 1795 -1245
rect 1990 -1246 2180 -1245
rect 2193 -1246 2376 -1245
rect 229 -1248 458 -1247
rect 527 -1248 832 -1247
rect 877 -1248 2096 -1247
rect 2200 -1248 2523 -1247
rect 303 -1250 535 -1249
rect 548 -1250 1182 -1249
rect 1206 -1250 1305 -1249
rect 1325 -1250 1333 -1249
rect 1416 -1250 2124 -1249
rect 2137 -1250 2201 -1249
rect 2228 -1250 2390 -1249
rect 331 -1252 388 -1251
rect 520 -1252 535 -1251
rect 562 -1252 787 -1251
rect 891 -1252 962 -1251
rect 975 -1252 1060 -1251
rect 1073 -1252 1179 -1251
rect 1241 -1252 1249 -1251
rect 1255 -1252 1389 -1251
rect 1423 -1252 1571 -1251
rect 1591 -1252 1725 -1251
rect 1759 -1252 1921 -1251
rect 2004 -1252 2187 -1251
rect 2242 -1252 2397 -1251
rect 205 -1254 521 -1253
rect 562 -1254 640 -1253
rect 660 -1254 1221 -1253
rect 1276 -1254 1389 -1253
rect 1447 -1254 2166 -1253
rect 2249 -1254 2425 -1253
rect 205 -1256 2075 -1255
rect 282 -1258 332 -1257
rect 607 -1258 815 -1257
rect 863 -1258 2243 -1257
rect 282 -1260 465 -1259
rect 541 -1260 815 -1259
rect 898 -1260 976 -1259
rect 985 -1260 1984 -1259
rect 2004 -1260 2131 -1259
rect 93 -1262 899 -1261
rect 919 -1262 1186 -1261
rect 1276 -1262 1298 -1261
rect 1367 -1262 1424 -1261
rect 1451 -1262 1697 -1261
rect 1703 -1262 1886 -1261
rect 1913 -1262 2124 -1261
rect 86 -1264 94 -1263
rect 110 -1264 1704 -1263
rect 1752 -1264 1914 -1263
rect 2018 -1264 2194 -1263
rect 86 -1266 598 -1265
rect 632 -1266 675 -1265
rect 709 -1266 920 -1265
rect 954 -1266 965 -1265
rect 1073 -1266 1217 -1265
rect 1325 -1266 1368 -1265
rect 1402 -1266 2166 -1265
rect 44 -1268 710 -1267
rect 723 -1268 1942 -1267
rect 2032 -1268 2229 -1267
rect 44 -1270 325 -1269
rect 464 -1270 836 -1269
rect 1080 -1270 1207 -1269
rect 1402 -1270 1410 -1269
rect 1507 -1270 1753 -1269
rect 1766 -1270 2019 -1269
rect 2039 -1270 2222 -1269
rect 243 -1272 325 -1271
rect 541 -1272 619 -1271
rect 625 -1272 633 -1271
rect 639 -1272 2418 -1271
rect 597 -1274 881 -1273
rect 989 -1274 1081 -1273
rect 1143 -1274 1361 -1273
rect 1528 -1274 1620 -1273
rect 1626 -1274 1760 -1273
rect 1773 -1274 1942 -1273
rect 2046 -1274 2250 -1273
rect 142 -1276 2047 -1275
rect 2053 -1276 2208 -1275
rect 142 -1278 825 -1277
rect 870 -1278 990 -1277
rect 1136 -1278 1627 -1277
rect 1640 -1278 1767 -1277
rect 1780 -1278 1935 -1277
rect 2011 -1278 2054 -1277
rect 618 -1280 1200 -1279
rect 1227 -1280 1410 -1279
rect 1535 -1280 1641 -1279
rect 1647 -1280 1774 -1279
rect 1780 -1280 1977 -1279
rect 625 -1282 780 -1281
rect 996 -1282 1137 -1281
rect 1143 -1282 1161 -1281
rect 1171 -1282 1228 -1281
rect 1237 -1282 1648 -1281
rect 1661 -1282 1844 -1281
rect 1850 -1282 2040 -1281
rect 660 -1284 892 -1283
rect 996 -1284 2173 -1283
rect 688 -1286 836 -1285
rect 999 -1286 1200 -1285
rect 1311 -1286 1508 -1285
rect 1542 -1286 1655 -1285
rect 1717 -1286 2012 -1285
rect 688 -1288 867 -1287
rect 1052 -1288 1172 -1287
rect 1391 -1288 1529 -1287
rect 1556 -1288 1662 -1287
rect 1787 -1288 2278 -1287
rect 765 -1290 1249 -1289
rect 1430 -1290 1718 -1289
rect 1808 -1290 1991 -1289
rect 695 -1292 766 -1291
rect 1024 -1292 1053 -1291
rect 1150 -1292 1298 -1291
rect 1430 -1292 1970 -1291
rect 695 -1294 941 -1293
rect 1024 -1294 1067 -1293
rect 1108 -1294 1151 -1293
rect 1213 -1294 1788 -1293
rect 1836 -1294 2033 -1293
rect 51 -1296 941 -1295
rect 1108 -1296 1130 -1295
rect 1153 -1296 1837 -1295
rect 1850 -1296 2393 -1295
rect 51 -1298 59 -1297
rect 450 -1298 1067 -1297
rect 1213 -1298 2215 -1297
rect 58 -1300 80 -1299
rect 450 -1300 577 -1299
rect 1017 -1300 1130 -1299
rect 1444 -1300 1536 -1299
rect 1556 -1300 2404 -1299
rect 352 -1302 577 -1301
rect 933 -1302 1018 -1301
rect 1479 -1302 1977 -1301
rect 2025 -1302 2215 -1301
rect 352 -1304 402 -1303
rect 793 -1304 934 -1303
rect 1013 -1304 2026 -1303
rect 2081 -1304 2404 -1303
rect 394 -1306 402 -1305
rect 761 -1306 2082 -1305
rect 212 -1308 395 -1307
rect 793 -1308 1998 -1307
rect 212 -1310 416 -1309
rect 1395 -1310 1480 -1309
rect 1493 -1310 1543 -1309
rect 1577 -1310 1697 -1309
rect 1864 -1310 2075 -1309
rect 170 -1312 416 -1311
rect 1006 -1312 1865 -1311
rect 1871 -1312 2131 -1311
rect 107 -1314 1007 -1313
rect 1346 -1314 1494 -1313
rect 1584 -1314 1725 -1313
rect 1878 -1314 2138 -1313
rect 170 -1316 738 -1315
rect 1395 -1316 1438 -1315
rect 1465 -1316 1879 -1315
rect 247 -1318 1347 -1317
rect 1472 -1318 1578 -1317
rect 1675 -1318 1809 -1317
rect 716 -1320 738 -1319
rect 779 -1320 1466 -1319
rect 1472 -1320 1711 -1319
rect 359 -1322 717 -1321
rect 1318 -1322 1438 -1321
rect 1486 -1322 1585 -1321
rect 1675 -1322 2236 -1321
rect 163 -1324 360 -1323
rect 1202 -1324 1319 -1323
rect 1374 -1324 1487 -1323
rect 1510 -1324 2236 -1323
rect 156 -1326 164 -1325
rect 177 -1326 1375 -1325
rect 1682 -1326 1872 -1325
rect 156 -1328 241 -1327
rect 1682 -1328 2327 -1327
rect 177 -1330 185 -1329
rect 240 -1330 297 -1329
rect 1689 -1330 1998 -1329
rect 184 -1332 290 -1331
rect 296 -1332 479 -1331
rect 1101 -1332 1690 -1331
rect 1710 -1332 1900 -1331
rect 289 -1334 472 -1333
rect 1822 -1334 2327 -1333
rect 317 -1336 479 -1335
rect 828 -1336 1823 -1335
rect 1899 -1336 2341 -1335
rect 317 -1338 727 -1337
rect 366 -1340 472 -1339
rect 345 -1342 367 -1341
rect 345 -1344 493 -1343
rect 338 -1346 493 -1345
rect 121 -1348 339 -1347
rect 2 -1359 839 -1358
rect 880 -1359 1137 -1358
rect 1150 -1359 2264 -1358
rect 2343 -1359 2579 -1358
rect 26 -1361 1578 -1360
rect 1794 -1361 1798 -1360
rect 2263 -1361 2362 -1360
rect 37 -1363 990 -1362
rect 996 -1363 1718 -1362
rect 1794 -1363 1851 -1362
rect 2361 -1363 2425 -1362
rect 40 -1365 1984 -1364
rect 44 -1367 202 -1366
rect 208 -1367 437 -1366
rect 464 -1367 909 -1366
rect 943 -1367 1977 -1366
rect 1983 -1367 2369 -1366
rect 44 -1369 87 -1368
rect 89 -1369 969 -1368
rect 989 -1369 1116 -1368
rect 1136 -1369 1193 -1368
rect 1213 -1369 1557 -1368
rect 1577 -1369 1606 -1368
rect 1717 -1369 1767 -1368
rect 1850 -1369 1914 -1368
rect 1976 -1369 2040 -1368
rect 2368 -1369 2432 -1368
rect 54 -1371 87 -1370
rect 93 -1371 125 -1370
rect 170 -1371 269 -1370
rect 317 -1371 465 -1370
rect 499 -1371 629 -1370
rect 642 -1371 969 -1370
rect 996 -1371 1501 -1370
rect 1507 -1371 1774 -1370
rect 1913 -1371 1963 -1370
rect 2431 -1371 2481 -1370
rect 58 -1373 62 -1372
rect 72 -1373 825 -1372
rect 831 -1373 906 -1372
rect 957 -1373 1424 -1372
rect 1426 -1373 1865 -1372
rect 1962 -1373 2033 -1372
rect 58 -1375 66 -1374
rect 79 -1375 157 -1374
rect 170 -1375 237 -1374
rect 240 -1375 640 -1374
rect 646 -1375 955 -1374
rect 982 -1375 2481 -1374
rect 82 -1377 1753 -1376
rect 1766 -1377 2110 -1376
rect 93 -1379 297 -1378
rect 317 -1379 888 -1378
rect 891 -1379 2530 -1378
rect 107 -1381 605 -1380
rect 646 -1381 654 -1380
rect 681 -1381 1000 -1380
rect 1006 -1381 1434 -1380
rect 1472 -1381 1753 -1380
rect 1773 -1381 1823 -1380
rect 1864 -1381 1921 -1380
rect 2109 -1381 2194 -1380
rect 2529 -1381 2558 -1380
rect 110 -1383 1788 -1382
rect 1797 -1383 2033 -1382
rect 2193 -1383 2292 -1382
rect 2340 -1383 2558 -1382
rect 117 -1385 209 -1384
rect 226 -1385 1375 -1384
rect 1430 -1385 1872 -1384
rect 2200 -1385 2341 -1384
rect 121 -1387 1235 -1386
rect 1251 -1387 2327 -1386
rect 107 -1389 122 -1388
rect 128 -1389 654 -1388
rect 681 -1389 738 -1388
rect 772 -1389 783 -1388
rect 796 -1389 913 -1388
rect 954 -1389 976 -1388
rect 982 -1389 1074 -1388
rect 1087 -1389 1193 -1388
rect 1213 -1389 1228 -1388
rect 1234 -1389 1305 -1388
rect 1332 -1389 1431 -1388
rect 1472 -1389 1487 -1388
rect 1500 -1389 2271 -1388
rect 128 -1391 993 -1390
rect 1013 -1391 1760 -1390
rect 1787 -1391 1837 -1390
rect 1871 -1391 1935 -1390
rect 2200 -1391 2509 -1390
rect 226 -1393 486 -1392
rect 516 -1393 570 -1392
rect 723 -1393 1091 -1392
rect 1104 -1393 1676 -1392
rect 1759 -1393 1816 -1392
rect 1822 -1393 1893 -1392
rect 1934 -1393 1998 -1392
rect 2270 -1393 2383 -1392
rect 2508 -1393 2523 -1392
rect 229 -1395 1921 -1394
rect 1997 -1395 2075 -1394
rect 2116 -1395 2383 -1394
rect 2522 -1395 2544 -1394
rect 240 -1397 752 -1396
rect 772 -1397 843 -1396
rect 880 -1397 920 -1396
rect 1038 -1397 1361 -1396
rect 1370 -1397 2425 -1396
rect 2543 -1397 2572 -1396
rect 254 -1399 689 -1398
rect 726 -1399 867 -1398
rect 891 -1399 962 -1398
rect 1031 -1399 1039 -1398
rect 1041 -1399 2166 -1398
rect 254 -1401 619 -1400
rect 688 -1401 759 -1400
rect 779 -1401 1879 -1400
rect 2165 -1401 2257 -1400
rect 296 -1403 895 -1402
rect 898 -1403 976 -1402
rect 1066 -1403 1102 -1402
rect 1115 -1403 1298 -1402
rect 1304 -1403 1452 -1402
rect 1482 -1403 2124 -1402
rect 2256 -1403 2355 -1402
rect 16 -1405 1452 -1404
rect 1510 -1405 2278 -1404
rect 16 -1407 2117 -1406
rect 2123 -1407 2208 -1406
rect 2277 -1407 2411 -1406
rect 310 -1409 605 -1408
rect 618 -1409 703 -1408
rect 730 -1409 741 -1408
rect 758 -1409 871 -1408
rect 905 -1409 2040 -1408
rect 2207 -1409 2446 -1408
rect 184 -1411 311 -1410
rect 408 -1411 864 -1410
rect 866 -1411 2131 -1410
rect 2410 -1411 2460 -1410
rect 184 -1413 276 -1412
rect 366 -1413 409 -1412
rect 415 -1413 608 -1412
rect 642 -1413 2355 -1412
rect 2445 -1413 2495 -1412
rect 257 -1415 416 -1414
rect 422 -1415 594 -1414
rect 702 -1415 1179 -1414
rect 1227 -1415 1249 -1414
rect 1258 -1415 2173 -1414
rect 219 -1417 423 -1416
rect 429 -1417 570 -1416
rect 730 -1417 1350 -1416
rect 1384 -1417 1676 -1416
rect 1682 -1417 2495 -1416
rect 19 -1419 430 -1418
rect 436 -1419 1312 -1418
rect 1332 -1419 1354 -1418
rect 1556 -1419 1585 -1418
rect 1591 -1419 1893 -1418
rect 2172 -1419 2243 -1418
rect 149 -1421 220 -1420
rect 247 -1421 1683 -1420
rect 1780 -1421 2075 -1420
rect 2242 -1421 2334 -1420
rect 149 -1423 766 -1422
rect 789 -1423 2460 -1422
rect 247 -1425 353 -1424
rect 366 -1425 493 -1424
rect 506 -1425 752 -1424
rect 765 -1425 1172 -1424
rect 1178 -1425 1291 -1424
rect 1297 -1425 1326 -1424
rect 1353 -1425 1494 -1424
rect 1584 -1425 1886 -1424
rect 142 -1427 1291 -1426
rect 1311 -1427 1340 -1426
rect 1591 -1427 1634 -1426
rect 1780 -1427 1830 -1426
rect 1836 -1427 1900 -1426
rect 142 -1429 986 -1428
rect 1003 -1429 1326 -1428
rect 1605 -1429 1648 -1428
rect 1815 -1429 1858 -1428
rect 1878 -1429 1956 -1428
rect 275 -1431 360 -1430
rect 471 -1431 507 -1430
rect 541 -1431 1011 -1430
rect 1024 -1431 1102 -1430
rect 1150 -1431 1186 -1430
rect 1241 -1431 1340 -1430
rect 1619 -1431 1830 -1430
rect 1857 -1431 1928 -1430
rect 1955 -1431 2026 -1430
rect 289 -1433 493 -1432
rect 541 -1433 1420 -1432
rect 1489 -1433 1620 -1432
rect 1633 -1433 1669 -1432
rect 1885 -1433 1949 -1432
rect 2025 -1433 2096 -1432
rect 289 -1435 549 -1434
rect 555 -1435 780 -1434
rect 814 -1435 1088 -1434
rect 1153 -1435 2292 -1434
rect 135 -1437 549 -1436
rect 716 -1437 1004 -1436
rect 1010 -1437 1053 -1436
rect 1059 -1437 1067 -1436
rect 1185 -1437 1207 -1436
rect 1241 -1437 1263 -1436
rect 1283 -1437 1361 -1436
rect 1647 -1437 1690 -1436
rect 1899 -1437 2180 -1436
rect 135 -1439 668 -1438
rect 716 -1439 829 -1438
rect 835 -1439 1074 -1438
rect 1206 -1439 1221 -1438
rect 1248 -1439 2327 -1438
rect 250 -1441 1221 -1440
rect 1255 -1441 1494 -1440
rect 1668 -1441 1725 -1440
rect 1927 -1441 2005 -1440
rect 2067 -1441 2180 -1440
rect 261 -1443 556 -1442
rect 677 -1443 1256 -1442
rect 1262 -1443 1270 -1442
rect 1283 -1443 1942 -1442
rect 1948 -1443 2019 -1442
rect 261 -1445 521 -1444
rect 674 -1445 1270 -1444
rect 1381 -1445 1690 -1444
rect 1941 -1445 2012 -1444
rect 2018 -1445 2089 -1444
rect 9 -1447 521 -1446
rect 674 -1447 692 -1446
rect 737 -1447 2131 -1446
rect 9 -1449 1266 -1448
rect 1381 -1449 1389 -1448
rect 1503 -1449 1725 -1448
rect 1969 -1449 2096 -1448
rect 303 -1451 360 -1450
rect 450 -1451 668 -1450
rect 744 -1451 1053 -1450
rect 1388 -1451 1403 -1450
rect 1514 -1451 2068 -1450
rect 2088 -1451 2187 -1450
rect 177 -1453 304 -1452
rect 352 -1453 374 -1452
rect 450 -1453 598 -1452
rect 709 -1453 745 -1452
rect 786 -1453 2187 -1452
rect 177 -1455 192 -1454
rect 271 -1455 710 -1454
rect 786 -1455 948 -1454
rect 1024 -1455 1165 -1454
rect 1276 -1455 1403 -1454
rect 1969 -1455 2061 -1454
rect 191 -1457 346 -1456
rect 373 -1457 402 -1456
rect 443 -1457 598 -1456
rect 660 -1457 948 -1456
rect 1031 -1457 1154 -1456
rect 1157 -1457 1515 -1456
rect 2004 -1457 2250 -1456
rect 331 -1459 346 -1458
rect 401 -1459 1287 -1458
rect 2011 -1459 2082 -1458
rect 2249 -1459 2348 -1458
rect 331 -1461 591 -1460
rect 632 -1461 661 -1460
rect 814 -1461 927 -1460
rect 940 -1461 1060 -1460
rect 1122 -1461 1277 -1460
rect 2060 -1461 2152 -1460
rect 2347 -1461 2418 -1460
rect 114 -1463 633 -1462
rect 828 -1463 1613 -1462
rect 2081 -1463 2159 -1462
rect 2417 -1463 2474 -1462
rect 51 -1465 115 -1464
rect 443 -1465 797 -1464
rect 835 -1465 850 -1464
rect 856 -1465 899 -1464
rect 912 -1465 1445 -1464
rect 1612 -1465 1655 -1464
rect 2151 -1465 2229 -1464
rect 2473 -1465 2516 -1464
rect 51 -1467 843 -1466
rect 870 -1467 885 -1466
rect 919 -1467 1018 -1466
rect 1122 -1467 1144 -1466
rect 1157 -1467 2453 -1466
rect 2515 -1467 2537 -1466
rect 471 -1469 801 -1468
rect 884 -1469 1564 -1468
rect 1654 -1469 1697 -1468
rect 2158 -1469 2236 -1468
rect 2452 -1469 2502 -1468
rect 2536 -1469 2551 -1468
rect 338 -1471 801 -1470
rect 926 -1471 934 -1470
rect 940 -1471 2334 -1470
rect 2375 -1471 2551 -1470
rect 205 -1473 934 -1472
rect 1017 -1473 2145 -1472
rect 2228 -1473 2313 -1472
rect 338 -1475 458 -1474
rect 478 -1475 500 -1474
rect 562 -1475 857 -1474
rect 877 -1475 2376 -1474
rect 23 -1477 563 -1476
rect 625 -1477 850 -1476
rect 1143 -1477 1522 -1476
rect 1563 -1477 1599 -1476
rect 1696 -1477 1732 -1476
rect 1990 -1477 2236 -1476
rect 2312 -1477 2397 -1476
rect 2 -1479 626 -1478
rect 793 -1479 1732 -1478
rect 1990 -1479 2299 -1478
rect 2396 -1479 2467 -1478
rect 23 -1481 2103 -1480
rect 2144 -1481 2222 -1480
rect 2284 -1481 2467 -1480
rect 156 -1483 878 -1482
rect 1160 -1483 1445 -1482
rect 1486 -1483 2502 -1482
rect 380 -1485 458 -1484
rect 485 -1485 514 -1484
rect 1164 -1485 1200 -1484
rect 1521 -1485 1543 -1484
rect 1598 -1485 1641 -1484
rect 2046 -1485 2222 -1484
rect 2284 -1485 2565 -1484
rect 47 -1487 514 -1486
rect 1080 -1487 1200 -1486
rect 1367 -1487 1641 -1486
rect 2046 -1487 2138 -1486
rect 2298 -1487 2390 -1486
rect 212 -1489 381 -1488
rect 394 -1489 479 -1488
rect 821 -1489 1368 -1488
rect 1542 -1489 1550 -1488
rect 2053 -1489 2103 -1488
rect 2137 -1489 2215 -1488
rect 2389 -1489 2439 -1488
rect 212 -1491 808 -1490
rect 1080 -1491 1095 -1490
rect 1549 -1491 1571 -1490
rect 1801 -1491 2054 -1490
rect 2214 -1491 2306 -1490
rect 2438 -1491 2488 -1490
rect 37 -1493 2488 -1492
rect 394 -1495 535 -1494
rect 807 -1495 1375 -1494
rect 1535 -1495 2306 -1494
rect 324 -1497 535 -1496
rect 1094 -1497 1109 -1496
rect 1395 -1497 1536 -1496
rect 1570 -1497 1627 -1496
rect 1801 -1497 1844 -1496
rect 324 -1499 612 -1498
rect 1045 -1499 1109 -1498
rect 1395 -1499 1410 -1498
rect 1626 -1499 1662 -1498
rect 1843 -1499 1907 -1498
rect 583 -1501 612 -1500
rect 695 -1501 1046 -1500
rect 1409 -1501 1529 -1500
rect 1661 -1501 1704 -1500
rect 1745 -1501 1907 -1500
rect 30 -1503 584 -1502
rect 639 -1503 1529 -1502
rect 1703 -1503 1739 -1502
rect 1745 -1503 1809 -1502
rect 30 -1505 528 -1504
rect 1416 -1505 1809 -1504
rect 100 -1507 528 -1506
rect 1416 -1507 1438 -1506
rect 1710 -1507 1739 -1506
rect 100 -1509 199 -1508
rect 233 -1509 696 -1508
rect 1437 -1509 1459 -1508
rect 72 -1511 234 -1510
rect 576 -1511 1711 -1510
rect 198 -1513 1172 -1512
rect 1458 -1513 1466 -1512
rect 576 -1515 962 -1514
rect 1465 -1515 1480 -1514
rect 1318 -1517 1480 -1516
rect 1318 -1519 1347 -1518
rect 1346 -1521 2320 -1520
rect 2319 -1523 2404 -1522
rect 1678 -1525 2404 -1524
rect 16 -1536 90 -1535
rect 93 -1536 209 -1535
rect 229 -1536 1711 -1535
rect 2389 -1536 2428 -1535
rect 2431 -1536 2435 -1535
rect 23 -1538 500 -1537
rect 583 -1538 794 -1537
rect 807 -1538 1333 -1537
rect 1360 -1538 1441 -1537
rect 1479 -1538 1977 -1537
rect 2284 -1538 2390 -1537
rect 23 -1540 629 -1539
rect 642 -1540 710 -1539
rect 719 -1540 2306 -1539
rect 40 -1542 829 -1541
rect 859 -1542 1494 -1541
rect 1496 -1542 2537 -1541
rect 44 -1544 55 -1543
rect 72 -1544 937 -1543
rect 943 -1544 1641 -1543
rect 1710 -1544 1823 -1543
rect 1976 -1544 2089 -1543
rect 2284 -1544 2418 -1543
rect 44 -1546 101 -1545
rect 107 -1546 811 -1545
rect 821 -1546 2033 -1545
rect 2305 -1546 2439 -1545
rect 47 -1548 423 -1547
rect 481 -1548 528 -1547
rect 583 -1548 661 -1547
rect 691 -1548 815 -1547
rect 821 -1548 1144 -1547
rect 1150 -1548 1585 -1547
rect 1822 -1548 1907 -1547
rect 1990 -1548 2089 -1547
rect 2340 -1548 2439 -1547
rect 30 -1550 423 -1549
rect 527 -1550 780 -1549
rect 793 -1550 990 -1549
rect 1076 -1550 2404 -1549
rect 30 -1552 283 -1551
rect 366 -1552 500 -1551
rect 590 -1552 605 -1551
rect 625 -1552 2054 -1551
rect 2403 -1552 2516 -1551
rect 51 -1554 304 -1553
rect 366 -1554 409 -1553
rect 590 -1554 619 -1553
rect 625 -1554 850 -1553
rect 880 -1554 1515 -1553
rect 1538 -1554 2124 -1553
rect 51 -1556 66 -1555
rect 72 -1556 262 -1555
rect 268 -1556 797 -1555
rect 814 -1556 1039 -1555
rect 1090 -1556 2411 -1555
rect 2 -1558 262 -1557
rect 268 -1558 724 -1557
rect 730 -1558 1021 -1557
rect 1038 -1558 1221 -1557
rect 1248 -1558 2348 -1557
rect 65 -1560 430 -1559
rect 604 -1560 1207 -1559
rect 1220 -1560 1312 -1559
rect 1332 -1560 1606 -1559
rect 1878 -1560 2054 -1559
rect 2123 -1560 2243 -1559
rect 2347 -1560 2474 -1559
rect 79 -1562 710 -1561
rect 723 -1562 1067 -1561
rect 1129 -1562 1207 -1561
rect 1248 -1562 1396 -1561
rect 1402 -1562 2418 -1561
rect 79 -1564 227 -1563
rect 233 -1564 521 -1563
rect 646 -1564 661 -1563
rect 698 -1564 2341 -1563
rect 100 -1566 472 -1565
rect 520 -1566 682 -1565
rect 702 -1566 885 -1565
rect 887 -1566 1025 -1565
rect 1066 -1566 1172 -1565
rect 1192 -1566 1252 -1565
rect 1255 -1566 1298 -1565
rect 1311 -1566 1459 -1565
rect 1479 -1566 1522 -1565
rect 1584 -1566 1676 -1565
rect 1878 -1566 1970 -1565
rect 1990 -1566 2061 -1565
rect 2095 -1566 2243 -1565
rect 37 -1568 1025 -1567
rect 1111 -1568 1676 -1567
rect 1906 -1568 2019 -1567
rect 2032 -1568 2145 -1567
rect 37 -1570 1613 -1569
rect 1955 -1570 2019 -1569
rect 2095 -1570 2215 -1569
rect 121 -1572 461 -1571
rect 471 -1572 507 -1571
rect 534 -1572 682 -1571
rect 702 -1572 752 -1571
rect 779 -1572 871 -1571
rect 898 -1572 941 -1571
rect 961 -1572 2173 -1571
rect 2214 -1572 2327 -1571
rect 114 -1574 752 -1573
rect 824 -1574 878 -1573
rect 898 -1574 1011 -1573
rect 1129 -1574 1235 -1573
rect 1283 -1574 1305 -1573
rect 1360 -1574 1865 -1573
rect 1955 -1574 2068 -1573
rect 2172 -1574 2292 -1573
rect 2326 -1574 2446 -1573
rect 114 -1576 202 -1575
rect 212 -1576 647 -1575
rect 737 -1576 1270 -1575
rect 1297 -1576 1354 -1575
rect 1395 -1576 1830 -1575
rect 1864 -1576 1942 -1575
rect 1969 -1576 2082 -1575
rect 2291 -1576 2362 -1575
rect 2445 -1576 2544 -1575
rect 121 -1578 913 -1577
rect 964 -1578 1403 -1577
rect 1423 -1578 1802 -1577
rect 1829 -1578 1963 -1577
rect 2067 -1578 2159 -1577
rect 2361 -1578 2488 -1577
rect 128 -1580 132 -1579
rect 198 -1580 2495 -1579
rect 128 -1582 675 -1581
rect 849 -1582 920 -1581
rect 989 -1582 1123 -1581
rect 1143 -1582 1179 -1581
rect 1192 -1582 1326 -1581
rect 1353 -1582 1550 -1581
rect 1605 -1582 1634 -1581
rect 1766 -1582 1942 -1581
rect 1962 -1582 2075 -1581
rect 2081 -1582 2194 -1581
rect 2494 -1582 2523 -1581
rect 184 -1584 199 -1583
rect 212 -1584 577 -1583
rect 593 -1584 2145 -1583
rect 2193 -1584 2299 -1583
rect 177 -1586 185 -1585
rect 219 -1586 962 -1585
rect 1122 -1586 1812 -1585
rect 2074 -1586 2166 -1585
rect 2298 -1586 2425 -1585
rect 135 -1588 220 -1587
rect 226 -1588 1011 -1587
rect 1153 -1588 1270 -1587
rect 1286 -1588 1802 -1587
rect 2165 -1588 2271 -1587
rect 135 -1590 1053 -1589
rect 1157 -1590 2222 -1589
rect 2270 -1590 2313 -1589
rect 233 -1592 696 -1591
rect 800 -1592 2425 -1591
rect 236 -1594 479 -1593
rect 506 -1594 542 -1593
rect 667 -1594 801 -1593
rect 870 -1594 1046 -1593
rect 1157 -1594 1375 -1593
rect 1423 -1594 1620 -1593
rect 1633 -1594 1739 -1593
rect 1766 -1594 1921 -1593
rect 2221 -1594 2278 -1593
rect 2312 -1594 2383 -1593
rect 240 -1596 1018 -1595
rect 1045 -1596 1109 -1595
rect 1160 -1596 1291 -1595
rect 1304 -1596 1438 -1595
rect 1458 -1596 1774 -1595
rect 2277 -1596 2397 -1595
rect 156 -1598 241 -1597
rect 247 -1598 409 -1597
rect 415 -1598 738 -1597
rect 828 -1598 1109 -1597
rect 1171 -1598 1417 -1597
rect 1486 -1598 1564 -1597
rect 1612 -1598 1795 -1597
rect 2382 -1598 2509 -1597
rect 156 -1600 171 -1599
rect 275 -1600 454 -1599
rect 464 -1600 535 -1599
rect 667 -1600 934 -1599
rect 954 -1600 1291 -1599
rect 1325 -1600 1445 -1599
rect 1489 -1600 2236 -1599
rect 2396 -1600 2481 -1599
rect 117 -1602 465 -1601
rect 478 -1602 493 -1601
rect 516 -1602 1053 -1601
rect 1178 -1602 1214 -1601
rect 1265 -1602 1774 -1601
rect 1794 -1602 1893 -1601
rect 2235 -1602 2355 -1601
rect 149 -1604 493 -1603
rect 674 -1604 892 -1603
rect 905 -1604 1452 -1603
rect 1493 -1604 1620 -1603
rect 1738 -1604 1788 -1603
rect 1892 -1604 1998 -1603
rect 2207 -1604 2355 -1603
rect 86 -1606 150 -1605
rect 170 -1606 255 -1605
rect 275 -1606 297 -1605
rect 303 -1606 402 -1605
rect 429 -1606 444 -1605
rect 695 -1606 773 -1605
rect 891 -1606 976 -1605
rect 982 -1606 1018 -1605
rect 1213 -1606 1753 -1605
rect 1759 -1606 1921 -1605
rect 1983 -1606 2208 -1605
rect 86 -1608 143 -1607
rect 250 -1608 1452 -1607
rect 1503 -1608 2467 -1607
rect 142 -1610 643 -1609
rect 772 -1610 843 -1609
rect 905 -1610 1382 -1609
rect 1416 -1610 1466 -1609
rect 1507 -1610 1641 -1609
rect 1752 -1610 1872 -1609
rect 1997 -1610 2103 -1609
rect 110 -1612 1466 -1611
rect 1514 -1612 1683 -1611
rect 1759 -1612 1900 -1611
rect 2102 -1612 2320 -1611
rect 205 -1614 1382 -1613
rect 1444 -1614 1599 -1613
rect 1787 -1614 2110 -1613
rect 2319 -1614 2530 -1613
rect 205 -1616 654 -1615
rect 842 -1616 927 -1615
rect 933 -1616 1116 -1615
rect 1234 -1616 1508 -1615
rect 1531 -1616 2159 -1615
rect 254 -1618 1154 -1617
rect 1276 -1618 1438 -1617
rect 1549 -1618 1669 -1617
rect 1815 -1618 1984 -1617
rect 282 -1620 374 -1619
rect 387 -1620 808 -1619
rect 912 -1620 1571 -1619
rect 1668 -1620 1781 -1619
rect 1871 -1620 1949 -1619
rect 96 -1622 1571 -1621
rect 1899 -1622 2012 -1621
rect 296 -1624 612 -1623
rect 919 -1624 1032 -1623
rect 1034 -1624 1599 -1623
rect 1927 -1624 2110 -1623
rect 338 -1626 402 -1625
rect 436 -1626 941 -1625
rect 954 -1626 1060 -1625
rect 1115 -1626 1137 -1625
rect 1258 -1626 1816 -1625
rect 1927 -1626 2026 -1625
rect 338 -1628 346 -1627
rect 352 -1628 416 -1627
rect 436 -1628 1501 -1627
rect 1563 -1628 1697 -1627
rect 1948 -1628 2047 -1627
rect 289 -1630 353 -1629
rect 373 -1630 458 -1629
rect 562 -1630 612 -1629
rect 926 -1630 1074 -1629
rect 1136 -1630 1319 -1629
rect 1349 -1630 1683 -1629
rect 1689 -1630 1697 -1629
rect 2004 -1630 2012 -1629
rect 2025 -1630 2131 -1629
rect 191 -1632 290 -1631
rect 317 -1632 346 -1631
rect 387 -1632 1004 -1631
rect 1059 -1632 1102 -1631
rect 1262 -1632 1781 -1631
rect 2004 -1632 2117 -1631
rect 2130 -1632 2250 -1631
rect 191 -1634 619 -1633
rect 975 -1634 1081 -1633
rect 1101 -1634 1228 -1633
rect 1276 -1634 1522 -1633
rect 1689 -1634 1809 -1633
rect 2046 -1634 2138 -1633
rect 2249 -1634 2460 -1633
rect 194 -1636 1263 -1635
rect 1318 -1636 1655 -1635
rect 1808 -1636 2180 -1635
rect 317 -1638 360 -1637
rect 394 -1638 640 -1637
rect 968 -1638 1228 -1637
rect 1293 -1638 1655 -1637
rect 2116 -1638 2229 -1637
rect 324 -1640 458 -1639
rect 548 -1640 563 -1639
rect 639 -1640 2551 -1639
rect 324 -1642 556 -1641
rect 856 -1642 969 -1641
rect 982 -1642 1165 -1641
rect 1374 -1642 1536 -1641
rect 2137 -1642 2376 -1641
rect 331 -1644 360 -1643
rect 394 -1644 633 -1643
rect 653 -1644 857 -1643
rect 1003 -1644 1186 -1643
rect 1500 -1644 1627 -1643
rect 2200 -1644 2376 -1643
rect 331 -1646 486 -1645
rect 548 -1646 759 -1645
rect 1073 -1646 2187 -1645
rect 2200 -1646 2264 -1645
rect 180 -1648 2187 -1647
rect 2228 -1648 2334 -1647
rect 443 -1650 1347 -1649
rect 1468 -1650 2264 -1649
rect 2333 -1650 2453 -1649
rect 450 -1652 633 -1651
rect 758 -1652 836 -1651
rect 996 -1652 1347 -1651
rect 1430 -1652 2453 -1651
rect 450 -1654 731 -1653
rect 765 -1654 836 -1653
rect 1080 -1654 1200 -1653
rect 1430 -1654 1557 -1653
rect 1626 -1654 1732 -1653
rect 485 -1656 717 -1655
rect 765 -1656 1088 -1655
rect 1164 -1656 1368 -1655
rect 1528 -1656 2180 -1655
rect 513 -1658 997 -1657
rect 1087 -1658 1364 -1657
rect 1367 -1658 1473 -1657
rect 1535 -1658 2061 -1657
rect 513 -1660 689 -1659
rect 786 -1660 1200 -1659
rect 1388 -1660 1529 -1659
rect 1556 -1660 1725 -1659
rect 131 -1662 787 -1661
rect 866 -1662 1732 -1661
rect 555 -1664 2442 -1663
rect 569 -1666 717 -1665
rect 1185 -1666 1242 -1665
rect 1388 -1666 1543 -1665
rect 1724 -1666 1851 -1665
rect 569 -1668 864 -1667
rect 1241 -1668 1340 -1667
rect 1472 -1668 1662 -1667
rect 1850 -1668 1935 -1667
rect 688 -1670 745 -1669
rect 863 -1670 948 -1669
rect 1339 -1670 1410 -1669
rect 1542 -1670 1648 -1669
rect 1661 -1670 1746 -1669
rect 1934 -1670 2040 -1669
rect 9 -1672 745 -1671
rect 947 -1672 2558 -1671
rect 93 -1674 2040 -1673
rect 1409 -1676 1592 -1675
rect 1745 -1676 1858 -1675
rect 1510 -1678 1858 -1677
rect 1577 -1680 1648 -1679
rect 1577 -1682 1704 -1681
rect 1591 -1684 1718 -1683
rect 1703 -1686 2411 -1685
rect 1717 -1688 1844 -1687
rect 1843 -1690 1914 -1689
rect 1913 -1692 2152 -1691
rect 2151 -1694 2257 -1693
rect 2256 -1696 2369 -1695
rect 2368 -1698 2502 -1697
rect 2 -1709 388 -1708
rect 429 -1709 1539 -1708
rect 1629 -1709 2047 -1708
rect 2389 -1709 2439 -1708
rect 2445 -1709 2460 -1708
rect 2469 -1709 2495 -1708
rect 9 -1711 108 -1710
rect 142 -1711 146 -1710
rect 187 -1711 1266 -1710
rect 1276 -1711 2411 -1710
rect 16 -1713 615 -1712
rect 649 -1713 944 -1712
rect 1017 -1713 1606 -1712
rect 1664 -1713 2313 -1712
rect 2347 -1713 2411 -1712
rect 16 -1715 1004 -1714
rect 1020 -1715 1193 -1714
rect 1206 -1715 1291 -1714
rect 1293 -1715 2271 -1714
rect 2389 -1715 2474 -1714
rect 30 -1717 895 -1716
rect 989 -1717 1018 -1716
rect 1031 -1717 1403 -1716
rect 1437 -1717 1739 -1716
rect 1801 -1717 2477 -1716
rect 30 -1719 332 -1718
rect 446 -1719 808 -1718
rect 821 -1719 1074 -1718
rect 1108 -1719 2418 -1718
rect 37 -1721 97 -1720
rect 107 -1721 374 -1720
rect 394 -1721 808 -1720
rect 821 -1721 1364 -1720
rect 1367 -1721 1403 -1720
rect 1440 -1721 2292 -1720
rect 2361 -1721 2418 -1720
rect 37 -1723 444 -1722
rect 457 -1723 829 -1722
rect 835 -1723 909 -1722
rect 961 -1723 1032 -1722
rect 1059 -1723 1063 -1722
rect 1111 -1723 1886 -1722
rect 1997 -1723 2047 -1722
rect 2228 -1723 2292 -1722
rect 2305 -1723 2362 -1722
rect 47 -1725 52 -1724
rect 65 -1725 181 -1724
rect 194 -1725 1102 -1724
rect 1153 -1725 1697 -1724
rect 1706 -1725 2376 -1724
rect 51 -1727 241 -1726
rect 247 -1727 535 -1726
rect 548 -1727 857 -1726
rect 870 -1727 962 -1726
rect 989 -1727 1011 -1726
rect 1059 -1727 1410 -1726
rect 1440 -1727 1704 -1726
rect 1836 -1727 2435 -1726
rect 58 -1729 66 -1728
rect 86 -1729 160 -1728
rect 198 -1729 1151 -1728
rect 1192 -1729 1284 -1728
rect 1293 -1729 1445 -1728
rect 1458 -1729 1998 -1728
rect 2039 -1729 2043 -1728
rect 2228 -1729 2320 -1728
rect 58 -1731 899 -1730
rect 957 -1731 1445 -1730
rect 1468 -1731 2397 -1730
rect 86 -1733 136 -1732
rect 142 -1733 451 -1732
rect 460 -1733 633 -1732
rect 653 -1733 829 -1732
rect 870 -1733 892 -1732
rect 1003 -1733 1095 -1732
rect 1143 -1733 1151 -1732
rect 1209 -1733 1375 -1732
rect 1388 -1733 1459 -1732
rect 1468 -1733 2320 -1732
rect 44 -1735 1375 -1734
rect 1493 -1735 1648 -1734
rect 1696 -1735 1942 -1734
rect 2039 -1735 2138 -1734
rect 2235 -1735 2306 -1734
rect 93 -1737 927 -1736
rect 1143 -1737 1182 -1736
rect 1213 -1737 1308 -1736
rect 1325 -1737 1368 -1736
rect 1493 -1737 1592 -1736
rect 1647 -1737 1809 -1736
rect 1815 -1737 1837 -1736
rect 1850 -1737 1886 -1736
rect 1941 -1737 2159 -1736
rect 2179 -1737 2236 -1736
rect 2242 -1737 2271 -1736
rect 2284 -1737 2376 -1736
rect 93 -1739 381 -1738
rect 429 -1739 927 -1738
rect 1171 -1739 1326 -1738
rect 1360 -1739 2208 -1738
rect 2221 -1739 2285 -1738
rect 135 -1741 206 -1740
rect 212 -1741 864 -1740
rect 884 -1741 1074 -1740
rect 1164 -1741 1172 -1740
rect 1213 -1741 1242 -1740
rect 1262 -1741 2019 -1740
rect 2081 -1741 2138 -1740
rect 2151 -1741 2222 -1740
rect 2263 -1741 2348 -1740
rect 100 -1743 206 -1742
rect 212 -1743 759 -1742
rect 793 -1743 1011 -1742
rect 1227 -1743 1389 -1742
rect 1510 -1743 2201 -1742
rect 198 -1745 367 -1744
rect 373 -1745 566 -1744
rect 579 -1745 1739 -1744
rect 1745 -1745 2243 -1744
rect 226 -1747 913 -1746
rect 940 -1747 1165 -1746
rect 1185 -1747 1228 -1746
rect 1241 -1747 1312 -1746
rect 1353 -1747 1361 -1746
rect 1528 -1747 2404 -1746
rect 229 -1749 1095 -1748
rect 1248 -1749 1263 -1748
rect 1283 -1749 1522 -1748
rect 1528 -1749 1543 -1748
rect 1556 -1749 1606 -1748
rect 1724 -1749 1746 -1748
rect 1759 -1749 2019 -1748
rect 2102 -1749 2264 -1748
rect 2333 -1749 2404 -1748
rect 124 -1751 1522 -1750
rect 1531 -1751 2313 -1750
rect 236 -1753 955 -1752
rect 1052 -1753 1186 -1752
rect 1297 -1753 1410 -1752
rect 1535 -1753 2089 -1752
rect 2130 -1753 2208 -1752
rect 240 -1755 1077 -1754
rect 1234 -1755 1298 -1754
rect 1304 -1755 1354 -1754
rect 1535 -1755 1613 -1754
rect 1619 -1755 1760 -1754
rect 1773 -1755 1816 -1754
rect 1850 -1755 2355 -1754
rect 289 -1757 699 -1756
rect 716 -1757 2159 -1756
rect 2165 -1757 2201 -1756
rect 2298 -1757 2355 -1756
rect 289 -1759 325 -1758
rect 331 -1759 514 -1758
rect 520 -1759 640 -1758
rect 653 -1759 738 -1758
rect 744 -1759 1053 -1758
rect 1157 -1759 1235 -1758
rect 1290 -1759 2166 -1758
rect 2179 -1759 2383 -1758
rect 324 -1761 591 -1760
rect 618 -1761 1109 -1760
rect 1115 -1761 1158 -1760
rect 1304 -1761 1802 -1760
rect 1808 -1761 1914 -1760
rect 2053 -1761 2103 -1760
rect 2151 -1761 2425 -1760
rect 121 -1763 619 -1762
rect 660 -1763 738 -1762
rect 744 -1763 906 -1762
rect 912 -1763 1046 -1762
rect 1496 -1763 2299 -1762
rect 2340 -1763 2383 -1762
rect 79 -1765 122 -1764
rect 345 -1765 367 -1764
rect 387 -1765 514 -1764
rect 520 -1765 612 -1764
rect 667 -1765 836 -1764
rect 849 -1765 885 -1764
rect 891 -1765 1984 -1764
rect 2004 -1765 2341 -1764
rect 79 -1767 269 -1766
rect 275 -1767 346 -1766
rect 352 -1767 381 -1766
rect 436 -1767 535 -1766
rect 548 -1767 948 -1766
rect 954 -1767 1280 -1766
rect 1556 -1767 1627 -1766
rect 1724 -1767 1872 -1766
rect 1934 -1767 1984 -1766
rect 2025 -1767 2054 -1766
rect 2249 -1767 2425 -1766
rect 149 -1769 437 -1768
rect 443 -1769 1543 -1768
rect 1563 -1769 1592 -1768
rect 1598 -1769 1613 -1768
rect 1619 -1769 1718 -1768
rect 1773 -1769 1900 -1768
rect 1955 -1769 2005 -1768
rect 2042 -1769 2082 -1768
rect 149 -1771 185 -1770
rect 268 -1771 339 -1770
rect 352 -1771 409 -1770
rect 481 -1771 1312 -1770
rect 1465 -1771 1935 -1770
rect 1969 -1771 2250 -1770
rect 114 -1773 339 -1772
rect 359 -1773 395 -1772
rect 408 -1773 416 -1772
rect 492 -1773 661 -1772
rect 667 -1773 682 -1772
rect 695 -1773 2446 -1772
rect 114 -1775 1424 -1774
rect 1465 -1775 1732 -1774
rect 1787 -1775 2334 -1774
rect 275 -1777 283 -1776
rect 317 -1777 360 -1776
rect 415 -1777 598 -1776
rect 646 -1777 948 -1776
rect 968 -1777 1914 -1776
rect 1927 -1777 1970 -1776
rect 1976 -1777 2026 -1776
rect 282 -1779 570 -1778
rect 590 -1779 689 -1778
rect 695 -1779 731 -1778
rect 733 -1779 997 -1778
rect 1045 -1779 1067 -1778
rect 1269 -1779 1424 -1778
rect 1479 -1779 1788 -1778
rect 1843 -1779 1872 -1778
rect 1878 -1779 1956 -1778
rect 1976 -1779 2173 -1778
rect 219 -1781 1270 -1780
rect 1276 -1781 1879 -1780
rect 2123 -1781 2173 -1780
rect 191 -1783 220 -1782
rect 296 -1783 598 -1782
rect 674 -1783 857 -1782
rect 863 -1783 1508 -1782
rect 1563 -1783 1795 -1782
rect 1857 -1783 1900 -1782
rect 2074 -1783 2124 -1782
rect 191 -1785 486 -1784
rect 492 -1785 507 -1784
rect 516 -1785 1067 -1784
rect 1472 -1785 1844 -1784
rect 2074 -1785 2327 -1784
rect 261 -1787 297 -1786
rect 310 -1787 318 -1786
rect 453 -1787 689 -1786
rect 716 -1787 752 -1786
rect 758 -1787 983 -1786
rect 1430 -1787 1473 -1786
rect 1479 -1787 1487 -1786
rect 1507 -1787 1991 -1786
rect 2116 -1787 2327 -1786
rect 250 -1789 262 -1788
rect 310 -1789 528 -1788
rect 562 -1789 577 -1788
rect 625 -1789 752 -1788
rect 779 -1789 794 -1788
rect 877 -1789 969 -1788
rect 971 -1789 2131 -1788
rect 100 -1791 563 -1790
rect 576 -1791 741 -1790
rect 803 -1791 878 -1790
rect 898 -1791 1280 -1790
rect 1332 -1791 1487 -1790
rect 1570 -1791 1599 -1790
rect 1675 -1791 1928 -1790
rect 1948 -1791 1991 -1790
rect 2060 -1791 2117 -1790
rect 128 -1793 528 -1792
rect 625 -1793 647 -1792
rect 674 -1793 710 -1792
rect 719 -1793 1249 -1792
rect 1346 -1793 1431 -1792
rect 1451 -1793 1571 -1792
rect 1661 -1793 1676 -1792
rect 1717 -1793 1854 -1792
rect 1920 -1793 1949 -1792
rect 2032 -1793 2061 -1792
rect 128 -1795 234 -1794
rect 464 -1795 682 -1794
rect 723 -1795 1102 -1794
rect 1199 -1795 1333 -1794
rect 1346 -1795 1578 -1794
rect 1752 -1795 1795 -1794
rect 1822 -1795 1858 -1794
rect 1892 -1795 1921 -1794
rect 2032 -1795 2442 -1794
rect 177 -1797 710 -1796
rect 730 -1797 1732 -1796
rect 1892 -1797 2096 -1796
rect 170 -1799 178 -1798
rect 201 -1799 780 -1798
rect 905 -1799 2397 -1798
rect 156 -1801 171 -1800
rect 215 -1801 1753 -1800
rect 2011 -1801 2096 -1800
rect 233 -1803 486 -1802
rect 499 -1803 570 -1802
rect 604 -1803 724 -1802
rect 933 -1803 2089 -1802
rect 464 -1805 472 -1804
rect 478 -1805 605 -1804
rect 611 -1805 1452 -1804
rect 1577 -1805 1585 -1804
rect 1962 -1805 2012 -1804
rect 72 -1807 472 -1806
rect 499 -1807 556 -1806
rect 936 -1807 997 -1806
rect 1024 -1807 1200 -1806
rect 1514 -1807 1585 -1806
rect 1710 -1807 1963 -1806
rect 72 -1809 402 -1808
rect 506 -1809 815 -1808
rect 940 -1809 2187 -1808
rect 184 -1811 479 -1810
rect 541 -1811 934 -1810
rect 975 -1811 983 -1810
rect 1024 -1811 1319 -1810
rect 1381 -1811 1515 -1810
rect 1689 -1811 1711 -1810
rect 2186 -1811 2467 -1810
rect 401 -1813 584 -1812
rect 814 -1813 843 -1812
rect 975 -1813 1039 -1812
rect 1136 -1813 1382 -1812
rect 1437 -1813 1690 -1812
rect 541 -1815 773 -1814
rect 786 -1815 843 -1814
rect 859 -1815 1039 -1814
rect 1136 -1815 1179 -1814
rect 1318 -1815 1340 -1814
rect 555 -1817 2428 -1816
rect 583 -1819 643 -1818
rect 772 -1819 801 -1818
rect 1178 -1819 1823 -1818
rect 786 -1821 1088 -1820
rect 1339 -1821 2453 -1820
rect 800 -1823 2068 -1822
rect 2193 -1823 2453 -1822
rect 1087 -1825 1123 -1824
rect 2067 -1825 2257 -1824
rect 1080 -1827 1123 -1826
rect 2144 -1827 2194 -1826
rect 2256 -1827 2432 -1826
rect 1080 -1829 1812 -1828
rect 2109 -1829 2145 -1828
rect 2368 -1829 2432 -1828
rect 1682 -1831 2110 -1830
rect 2277 -1831 2369 -1830
rect 1668 -1833 1683 -1832
rect 2214 -1833 2278 -1832
rect 1654 -1835 1669 -1834
rect 1906 -1835 2215 -1834
rect 1633 -1837 1655 -1836
rect 1864 -1837 1907 -1836
rect 1633 -1839 1767 -1838
rect 1766 -1841 1830 -1840
rect 1780 -1843 1830 -1842
rect 1395 -1845 1781 -1844
rect 1395 -1847 1417 -1846
rect 1416 -1849 1627 -1848
rect 30 -1860 612 -1859
rect 618 -1860 1182 -1859
rect 1206 -1860 1627 -1859
rect 1636 -1860 2369 -1859
rect 30 -1862 150 -1861
rect 184 -1862 1928 -1861
rect 2270 -1862 2470 -1861
rect 37 -1864 619 -1863
rect 632 -1864 1291 -1863
rect 1307 -1864 1648 -1863
rect 1664 -1864 2110 -1863
rect 2319 -1864 2421 -1863
rect 37 -1866 192 -1865
rect 194 -1866 615 -1865
rect 635 -1866 1200 -1865
rect 1206 -1866 1221 -1865
rect 1241 -1866 1245 -1865
rect 1276 -1866 1963 -1865
rect 2109 -1866 2278 -1865
rect 2319 -1866 2418 -1865
rect 47 -1868 2243 -1867
rect 2368 -1868 2411 -1867
rect 72 -1870 801 -1869
rect 852 -1870 1382 -1869
rect 1437 -1870 2222 -1869
rect 2410 -1870 2460 -1869
rect 72 -1872 129 -1871
rect 131 -1872 2271 -1871
rect 89 -1874 1732 -1873
rect 1734 -1874 2453 -1873
rect 100 -1876 188 -1875
rect 215 -1876 1301 -1875
rect 1332 -1876 1336 -1875
rect 1363 -1876 1935 -1875
rect 1962 -1876 1991 -1875
rect 2067 -1876 2278 -1875
rect 100 -1878 1424 -1877
rect 1468 -1878 2208 -1877
rect 2221 -1878 2285 -1877
rect 107 -1880 517 -1879
rect 548 -1880 1441 -1879
rect 1475 -1880 2250 -1879
rect 2256 -1880 2285 -1879
rect 107 -1882 136 -1881
rect 142 -1882 1154 -1881
rect 1164 -1882 1221 -1881
rect 1241 -1882 1326 -1881
rect 1332 -1882 1340 -1881
rect 1353 -1882 1424 -1881
rect 1489 -1882 1578 -1881
rect 1622 -1882 1956 -1881
rect 2067 -1882 2124 -1881
rect 2249 -1882 2292 -1881
rect 103 -1884 136 -1883
rect 142 -1884 381 -1883
rect 401 -1884 650 -1883
rect 688 -1884 731 -1883
rect 737 -1884 1025 -1883
rect 1059 -1884 1070 -1883
rect 1094 -1884 1732 -1883
rect 1773 -1884 1991 -1883
rect 2256 -1884 2306 -1883
rect 16 -1886 1095 -1885
rect 1136 -1886 2089 -1885
rect 16 -1888 353 -1887
rect 373 -1888 587 -1887
rect 611 -1888 682 -1887
rect 688 -1888 787 -1887
rect 894 -1888 1998 -1887
rect 124 -1890 1102 -1889
rect 1129 -1890 1137 -1889
rect 1150 -1890 1200 -1889
rect 1209 -1890 2446 -1889
rect 128 -1892 1074 -1891
rect 1080 -1892 1102 -1891
rect 1129 -1892 1140 -1891
rect 1164 -1892 1459 -1891
rect 1507 -1892 2390 -1891
rect 184 -1894 220 -1893
rect 233 -1894 2124 -1893
rect 2228 -1894 2390 -1893
rect 177 -1896 234 -1895
rect 250 -1896 1431 -1895
rect 1440 -1896 2292 -1895
rect 177 -1898 262 -1897
rect 275 -1898 430 -1897
rect 446 -1898 465 -1897
rect 478 -1898 783 -1897
rect 905 -1898 1613 -1897
rect 1633 -1898 1998 -1897
rect 2032 -1898 2229 -1897
rect 205 -1900 381 -1899
rect 401 -1900 633 -1899
rect 646 -1900 1270 -1899
rect 1290 -1900 1298 -1899
rect 1304 -1900 2208 -1899
rect 205 -1902 283 -1901
rect 303 -1902 353 -1901
rect 373 -1902 822 -1901
rect 908 -1902 948 -1901
rect 957 -1902 1844 -1901
rect 1853 -1902 2425 -1901
rect 51 -1904 283 -1903
rect 303 -1904 451 -1903
rect 464 -1904 528 -1903
rect 541 -1904 731 -1903
rect 744 -1904 1277 -1903
rect 1339 -1904 1368 -1903
rect 1381 -1904 1417 -1903
rect 1430 -1904 1452 -1903
rect 1458 -1904 1473 -1903
rect 1507 -1904 1585 -1903
rect 1605 -1904 1613 -1903
rect 1647 -1904 1851 -1903
rect 1864 -1904 2404 -1903
rect 51 -1906 1606 -1905
rect 1664 -1906 2376 -1905
rect 2403 -1906 2439 -1905
rect 219 -1908 1522 -1907
rect 1577 -1908 1592 -1907
rect 1773 -1908 1823 -1907
rect 1843 -1908 2082 -1907
rect 226 -1910 2376 -1909
rect 170 -1912 227 -1911
rect 261 -1912 269 -1911
rect 275 -1912 542 -1911
rect 562 -1912 1109 -1911
rect 1167 -1912 2306 -1911
rect 156 -1914 269 -1913
rect 394 -1914 528 -1913
rect 565 -1914 1053 -1913
rect 1059 -1914 1347 -1913
rect 1353 -1914 1403 -1913
rect 1416 -1914 1501 -1913
rect 1584 -1914 1620 -1913
rect 1822 -1914 1837 -1913
rect 1850 -1914 1879 -1913
rect 1934 -1914 1970 -1913
rect 2032 -1914 2145 -1913
rect 170 -1916 2159 -1915
rect 173 -1918 2159 -1917
rect 229 -1920 1837 -1919
rect 1864 -1920 1900 -1919
rect 1941 -1920 2145 -1919
rect 240 -1922 395 -1921
rect 422 -1922 549 -1921
rect 569 -1922 741 -1921
rect 744 -1922 808 -1921
rect 821 -1922 941 -1921
rect 943 -1922 1186 -1921
rect 1227 -1922 1270 -1921
rect 1346 -1922 1571 -1921
rect 1591 -1922 1781 -1921
rect 1878 -1922 1914 -1921
rect 1941 -1922 1984 -1921
rect 2081 -1922 2138 -1921
rect 2 -1924 241 -1923
rect 422 -1924 545 -1923
rect 646 -1924 864 -1923
rect 919 -1924 948 -1923
rect 957 -1924 2243 -1923
rect 2 -1926 738 -1925
rect 807 -1926 1011 -1925
rect 1024 -1926 1438 -1925
rect 1444 -1926 1571 -1925
rect 1780 -1926 1830 -1925
rect 1899 -1926 2467 -1925
rect 159 -1928 1011 -1927
rect 1038 -1928 1081 -1927
rect 1178 -1928 2334 -1927
rect 9 -1930 160 -1929
rect 429 -1930 500 -1929
rect 506 -1930 741 -1929
rect 863 -1930 976 -1929
rect 978 -1930 1511 -1929
rect 1913 -1930 1949 -1929
rect 1955 -1930 2012 -1929
rect 2074 -1930 2334 -1929
rect 9 -1932 199 -1931
rect 324 -1932 500 -1931
rect 506 -1932 878 -1931
rect 919 -1932 1123 -1931
rect 1178 -1932 1630 -1931
rect 1696 -1932 1949 -1931
rect 1969 -1932 2005 -1931
rect 2011 -1932 2061 -1931
rect 2074 -1932 2131 -1931
rect 2137 -1932 2194 -1931
rect 58 -1934 1039 -1933
rect 1062 -1934 2299 -1933
rect 23 -1936 59 -1935
rect 198 -1936 1004 -1935
rect 1066 -1936 1620 -1935
rect 1696 -1936 1704 -1935
rect 1983 -1936 2026 -1935
rect 2060 -1936 2117 -1935
rect 2130 -1936 2173 -1935
rect 2298 -1936 2313 -1935
rect 23 -1938 115 -1937
rect 324 -1938 1466 -1937
rect 1472 -1938 2425 -1937
rect 114 -1940 759 -1939
rect 828 -1940 878 -1939
rect 926 -1940 1305 -1939
rect 1367 -1940 1410 -1939
rect 1444 -1940 1480 -1939
rect 1486 -1940 1501 -1939
rect 1703 -1940 1886 -1939
rect 1892 -1940 2117 -1939
rect 2312 -1940 2348 -1939
rect 432 -1942 570 -1941
rect 674 -1942 682 -1941
rect 695 -1942 1004 -1941
rect 1066 -1942 1116 -1941
rect 1185 -1942 1319 -1941
rect 1335 -1942 1410 -1941
rect 1451 -1942 1599 -1941
rect 1724 -1942 2026 -1941
rect 2347 -1942 2383 -1941
rect 191 -1944 675 -1943
rect 702 -1944 955 -1943
rect 975 -1944 1753 -1943
rect 1766 -1944 1886 -1943
rect 1892 -1944 2166 -1943
rect 2179 -1944 2383 -1943
rect 450 -1946 591 -1945
rect 660 -1946 696 -1945
rect 702 -1946 997 -1945
rect 1073 -1946 1868 -1945
rect 1976 -1946 2173 -1945
rect 2179 -1946 2236 -1945
rect 121 -1948 661 -1947
rect 709 -1948 941 -1947
rect 982 -1948 997 -1947
rect 1087 -1948 1116 -1947
rect 1125 -1948 1977 -1947
rect 2004 -1948 2054 -1947
rect 86 -1950 983 -1949
rect 1111 -1950 2194 -1949
rect 121 -1952 297 -1951
rect 443 -1952 1088 -1951
rect 1227 -1952 2236 -1951
rect 296 -1954 360 -1953
rect 443 -1954 556 -1953
rect 590 -1954 727 -1953
rect 772 -1954 955 -1953
rect 1248 -1954 1830 -1953
rect 2053 -1954 2103 -1953
rect 289 -1956 556 -1955
rect 653 -1956 710 -1955
rect 723 -1956 759 -1955
rect 772 -1956 923 -1955
rect 926 -1956 1046 -1955
rect 1213 -1956 1249 -1955
rect 1395 -1956 1403 -1955
rect 1465 -1956 1634 -1955
rect 1654 -1956 1725 -1955
rect 1752 -1956 1760 -1955
rect 1766 -1956 1816 -1955
rect 2102 -1956 2152 -1955
rect 289 -1958 850 -1957
rect 933 -1958 1319 -1957
rect 1360 -1958 1396 -1957
rect 1486 -1958 1928 -1957
rect 2151 -1958 2201 -1957
rect 359 -1960 437 -1959
rect 478 -1960 605 -1959
rect 653 -1960 843 -1959
rect 849 -1960 899 -1959
rect 933 -1960 2474 -1959
rect 436 -1962 598 -1961
rect 604 -1962 752 -1961
rect 842 -1962 857 -1961
rect 1017 -1962 1046 -1961
rect 1213 -1962 1235 -1961
rect 1279 -1962 1816 -1961
rect 310 -1964 1018 -1963
rect 1234 -1964 1312 -1963
rect 1360 -1964 2089 -1963
rect 310 -1966 318 -1965
rect 485 -1966 563 -1965
rect 576 -1966 857 -1965
rect 1297 -1966 2201 -1965
rect 212 -1968 318 -1967
rect 485 -1968 493 -1967
rect 513 -1968 804 -1967
rect 1311 -1968 1662 -1967
rect 1675 -1968 1760 -1967
rect 1801 -1968 2166 -1967
rect 149 -1970 213 -1969
rect 247 -1970 493 -1969
rect 534 -1970 598 -1969
rect 625 -1970 899 -1969
rect 1549 -1970 1599 -1969
rect 1654 -1970 1746 -1969
rect 1801 -1970 1858 -1969
rect 86 -1972 248 -1971
rect 387 -1972 514 -1971
rect 576 -1972 794 -1971
rect 1524 -1972 1746 -1971
rect 93 -1974 535 -1973
rect 716 -1974 724 -1973
rect 751 -1974 892 -1973
rect 1535 -1974 1858 -1973
rect 93 -1976 339 -1975
rect 387 -1976 416 -1975
rect 457 -1976 626 -1975
rect 639 -1976 717 -1975
rect 793 -1976 1109 -1975
rect 1549 -1976 2341 -1975
rect 79 -1978 640 -1977
rect 828 -1978 2341 -1977
rect 79 -1980 832 -1979
rect 870 -1980 892 -1979
rect 1052 -1980 1536 -1979
rect 1661 -1980 2327 -1979
rect 254 -1982 458 -1981
rect 870 -1982 913 -1981
rect 1675 -1982 1683 -1981
rect 2326 -1982 2362 -1981
rect 44 -1984 255 -1983
rect 331 -1984 339 -1983
rect 345 -1984 416 -1983
rect 583 -1984 913 -1983
rect 1682 -1984 1690 -1983
rect 2361 -1984 2397 -1983
rect 44 -1986 66 -1985
rect 331 -1986 1263 -1985
rect 1689 -1986 1711 -1985
rect 1787 -1986 2397 -1985
rect 65 -1988 1375 -1987
rect 1563 -1988 1788 -1987
rect 345 -1990 367 -1989
rect 583 -1990 787 -1989
rect 1255 -1990 1263 -1989
rect 1283 -1990 1564 -1989
rect 1710 -1990 1739 -1989
rect 366 -1992 409 -1991
rect 1171 -1992 1256 -1991
rect 1374 -1992 1389 -1991
rect 1640 -1992 1739 -1991
rect 408 -1994 472 -1993
rect 765 -1994 1172 -1993
rect 1192 -1994 1284 -1993
rect 1388 -1994 1497 -1993
rect 1556 -1994 1641 -1993
rect 471 -1996 521 -1995
rect 765 -1996 1032 -1995
rect 1157 -1996 1193 -1995
rect 1514 -1996 1557 -1995
rect 520 -1998 668 -1997
rect 989 -1998 1032 -1997
rect 1143 -1998 1158 -1997
rect 1514 -1998 1543 -1997
rect 635 -2000 668 -1999
rect 779 -2000 1144 -1999
rect 1493 -2000 1543 -1999
rect 968 -2002 990 -2001
rect 1493 -2002 2215 -2001
rect 884 -2004 969 -2003
rect 2214 -2004 2264 -2003
rect 884 -2006 1669 -2005
rect 2039 -2006 2264 -2005
rect 1668 -2008 1795 -2007
rect 2039 -2008 2096 -2007
rect 1794 -2010 2019 -2009
rect 2095 -2010 2355 -2009
rect 1808 -2012 2019 -2011
rect 2354 -2012 2432 -2011
rect 1808 -2014 1872 -2013
rect 1871 -2016 1907 -2015
rect 1906 -2018 1921 -2017
rect 1920 -2020 2047 -2019
rect 1717 -2022 2047 -2021
rect 779 -2024 1718 -2023
rect 9 -2035 762 -2034
rect 800 -2035 850 -2034
rect 898 -2035 1109 -2034
rect 1111 -2035 1207 -2034
rect 1230 -2035 1301 -2034
rect 1335 -2035 1977 -2034
rect 2403 -2035 2418 -2034
rect 9 -2037 45 -2036
rect 51 -2037 66 -2036
rect 86 -2037 136 -2036
rect 138 -2037 1018 -2036
rect 1024 -2037 1109 -2036
rect 1122 -2037 1424 -2036
rect 1437 -2037 2425 -2036
rect 37 -2039 832 -2038
rect 898 -2039 1305 -2038
rect 1360 -2039 1641 -2038
rect 1713 -2039 1970 -2038
rect 37 -2041 241 -2040
rect 296 -2041 1063 -2040
rect 1073 -2041 1207 -2040
rect 1297 -2041 1858 -2040
rect 1934 -2041 2404 -2040
rect 30 -2043 241 -2042
rect 296 -2043 472 -2042
rect 492 -2043 1018 -2042
rect 1024 -2043 1431 -2042
rect 1437 -2043 1445 -2042
rect 1472 -2043 1879 -2042
rect 1969 -2043 2376 -2042
rect 16 -2045 472 -2044
rect 499 -2045 542 -2044
rect 569 -2045 1123 -2044
rect 1150 -2045 2292 -2044
rect 2340 -2045 2376 -2044
rect 16 -2047 808 -2046
rect 828 -2047 1410 -2046
rect 1430 -2047 1984 -2046
rect 2249 -2047 2292 -2046
rect 2298 -2047 2341 -2046
rect 30 -2049 73 -2048
rect 89 -2049 885 -2048
rect 919 -2049 927 -2048
rect 954 -2049 2355 -2048
rect 44 -2051 696 -2050
rect 751 -2051 850 -2050
rect 922 -2051 1032 -2050
rect 1153 -2051 1396 -2050
rect 1402 -2051 1424 -2050
rect 1440 -2051 2117 -2050
rect 2214 -2051 2250 -2050
rect 2 -2053 1154 -2052
rect 1171 -2053 1343 -2052
rect 1363 -2053 2229 -2052
rect 51 -2055 1697 -2054
rect 1766 -2055 2425 -2054
rect 58 -2057 1361 -2056
rect 1384 -2057 1599 -2056
rect 1605 -2057 1697 -2056
rect 1808 -2057 1879 -2056
rect 2095 -2057 2355 -2056
rect 58 -2059 97 -2058
rect 100 -2059 108 -2058
rect 156 -2059 2306 -2058
rect 65 -2061 703 -2060
rect 758 -2061 804 -2060
rect 807 -2061 1319 -2060
rect 1402 -2061 2026 -2060
rect 2095 -2061 2187 -2060
rect 2228 -2061 2285 -2060
rect 2305 -2061 2313 -2060
rect 72 -2063 962 -2062
rect 1031 -2063 1130 -2062
rect 1178 -2063 1641 -2062
rect 1654 -2063 1809 -2062
rect 1815 -2063 1977 -2062
rect 2046 -2063 2313 -2062
rect 100 -2065 1406 -2064
rect 1409 -2065 1886 -2064
rect 1920 -2065 2047 -2064
rect 2116 -2065 2131 -2064
rect 2172 -2065 2215 -2064
rect 2256 -2065 2285 -2064
rect 107 -2067 1168 -2066
rect 1178 -2067 1193 -2066
rect 1220 -2067 1319 -2066
rect 1486 -2067 1991 -2066
rect 2074 -2067 2131 -2066
rect 2137 -2067 2173 -2066
rect 2186 -2067 2348 -2066
rect 156 -2069 458 -2068
rect 516 -2069 1004 -2068
rect 1038 -2069 1130 -2068
rect 1192 -2069 1291 -2068
rect 1297 -2069 1308 -2068
rect 1486 -2069 1725 -2068
rect 1745 -2069 1816 -2068
rect 1871 -2069 1921 -2068
rect 1948 -2069 1991 -2068
rect 2018 -2069 2075 -2068
rect 2081 -2069 2138 -2068
rect 2207 -2069 2257 -2068
rect 2333 -2069 2348 -2068
rect 159 -2071 906 -2070
rect 1003 -2071 1256 -2070
rect 1269 -2071 1984 -2070
rect 173 -2073 1242 -2072
rect 1276 -2073 1396 -2072
rect 1489 -2073 2299 -2072
rect 191 -2075 507 -2074
rect 569 -2075 979 -2074
rect 1038 -2075 1067 -2074
rect 1080 -2075 1172 -2074
rect 1234 -2075 1445 -2074
rect 1521 -2075 1760 -2074
rect 1843 -2075 2082 -2074
rect 191 -2077 587 -2076
rect 590 -2077 657 -2076
rect 670 -2077 745 -2076
rect 758 -2077 885 -2076
rect 891 -2077 906 -2076
rect 978 -2077 1823 -2076
rect 1871 -2077 1942 -2076
rect 1955 -2077 2019 -2076
rect 170 -2079 591 -2078
rect 604 -2079 780 -2078
rect 786 -2079 801 -2078
rect 828 -2079 969 -2078
rect 989 -2079 1235 -2078
rect 1283 -2079 1291 -2078
rect 1304 -2079 1417 -2078
rect 1521 -2079 1613 -2078
rect 1622 -2079 2033 -2078
rect 170 -2081 731 -2080
rect 740 -2081 2026 -2080
rect 194 -2083 1725 -2082
rect 1752 -2083 1823 -2082
rect 1899 -2083 1942 -2082
rect 1955 -2083 2390 -2082
rect 212 -2085 318 -2084
rect 331 -2085 962 -2084
rect 1059 -2085 2334 -2084
rect 2361 -2085 2390 -2084
rect 93 -2087 332 -2086
rect 338 -2087 458 -2086
rect 464 -2087 605 -2086
rect 618 -2087 752 -2086
rect 793 -2087 927 -2086
rect 940 -2087 990 -2086
rect 1066 -2087 1665 -2086
rect 1689 -2087 1767 -2086
rect 1773 -2087 1844 -2086
rect 1850 -2087 1900 -2086
rect 1906 -2087 1949 -2086
rect 2326 -2087 2362 -2086
rect 93 -2089 1466 -2088
rect 1479 -2089 1753 -2088
rect 1780 -2089 1851 -2088
rect 2004 -2089 2327 -2088
rect 103 -2091 1774 -2090
rect 1780 -2091 1914 -2090
rect 114 -2093 794 -2092
rect 835 -2093 920 -2092
rect 940 -2093 983 -2092
rect 1080 -2093 1095 -2092
rect 1143 -2093 1242 -2092
rect 1311 -2093 1417 -2092
rect 1451 -2093 1690 -2092
rect 1703 -2093 1907 -2092
rect 114 -2095 353 -2094
rect 366 -2095 465 -2094
rect 562 -2095 619 -2094
rect 653 -2095 955 -2094
rect 1094 -2095 1102 -2094
rect 1136 -2095 1312 -2094
rect 1332 -2095 1466 -2094
rect 1500 -2095 1613 -2094
rect 1626 -2095 1746 -2094
rect 1794 -2095 2033 -2094
rect 205 -2097 353 -2096
rect 404 -2097 969 -2096
rect 1010 -2097 1102 -2096
rect 1136 -2097 1214 -2096
rect 1325 -2097 1501 -2096
rect 1528 -2097 1655 -2096
rect 1703 -2097 1865 -2096
rect 177 -2099 206 -2098
rect 215 -2099 1732 -2098
rect 1801 -2099 1865 -2098
rect 163 -2101 178 -2100
rect 219 -2101 1060 -2100
rect 1143 -2101 1224 -2100
rect 1262 -2101 1326 -2100
rect 1332 -2101 2271 -2100
rect 124 -2103 164 -2102
rect 219 -2103 1651 -2102
rect 2221 -2103 2271 -2102
rect 236 -2105 682 -2104
rect 688 -2105 1277 -2104
rect 1353 -2105 1529 -2104
rect 1535 -2105 1963 -2104
rect 2179 -2105 2222 -2104
rect 247 -2107 1760 -2106
rect 1927 -2107 1963 -2106
rect 2165 -2107 2180 -2106
rect 247 -2109 290 -2108
rect 303 -2109 507 -2108
rect 583 -2109 612 -2108
rect 625 -2109 682 -2108
rect 695 -2109 958 -2108
rect 1010 -2109 1046 -2108
rect 1164 -2109 2005 -2108
rect 2123 -2109 2166 -2108
rect 261 -2111 318 -2110
rect 338 -2111 1553 -2110
rect 1563 -2111 1935 -2110
rect 2067 -2111 2124 -2110
rect 142 -2113 262 -2112
rect 275 -2113 689 -2112
rect 702 -2113 1259 -2112
rect 1262 -2113 1476 -2112
rect 1538 -2113 1928 -2112
rect 2011 -2113 2068 -2112
rect 142 -2115 1581 -2114
rect 1584 -2115 1795 -2114
rect 275 -2117 549 -2116
rect 597 -2117 612 -2116
rect 625 -2117 857 -2116
rect 863 -2117 1270 -2116
rect 1367 -2117 1536 -2116
rect 1542 -2117 1914 -2116
rect 289 -2119 388 -2118
rect 422 -2119 1074 -2118
rect 1164 -2119 1200 -2118
rect 1213 -2119 1494 -2118
rect 1549 -2119 2110 -2118
rect 226 -2121 388 -2120
rect 436 -2121 598 -2120
rect 653 -2121 2208 -2120
rect 226 -2123 647 -2122
rect 660 -2123 1627 -2122
rect 1636 -2123 2012 -2122
rect 2060 -2123 2110 -2122
rect 233 -2125 423 -2124
rect 443 -2125 647 -2124
rect 660 -2125 976 -2124
rect 1188 -2125 1284 -2124
rect 1339 -2125 1494 -2124
rect 1549 -2125 1634 -2124
rect 2060 -2125 2264 -2124
rect 303 -2127 556 -2126
rect 576 -2127 864 -2126
rect 891 -2127 1620 -2126
rect 1633 -2127 1711 -2126
rect 2235 -2127 2264 -2126
rect 23 -2129 1620 -2128
rect 2193 -2129 2236 -2128
rect 23 -2131 132 -2130
rect 345 -2131 367 -2130
rect 373 -2131 549 -2130
rect 555 -2131 871 -2130
rect 933 -2131 1046 -2130
rect 1188 -2131 1998 -2130
rect 2151 -2131 2194 -2130
rect 131 -2133 213 -2132
rect 345 -2133 402 -2132
rect 443 -2133 997 -2132
rect 1199 -2133 2320 -2132
rect 149 -2135 871 -2134
rect 947 -2135 983 -2134
rect 1248 -2135 1354 -2134
rect 1381 -2135 1543 -2134
rect 1563 -2135 1788 -2134
rect 2151 -2135 2383 -2134
rect 54 -2137 150 -2136
rect 373 -2137 1203 -2136
rect 1381 -2137 1998 -2136
rect 2144 -2137 2383 -2136
rect 394 -2139 437 -2138
rect 450 -2139 633 -2138
rect 639 -2139 997 -2138
rect 1157 -2139 1249 -2138
rect 1570 -2139 1802 -2138
rect 2088 -2139 2145 -2138
rect 79 -2141 395 -2140
rect 401 -2141 409 -2140
rect 492 -2141 563 -2140
rect 632 -2141 1056 -2140
rect 1125 -2141 1158 -2140
rect 1458 -2141 1571 -2140
rect 1577 -2141 1886 -2140
rect 2039 -2141 2089 -2140
rect 79 -2143 535 -2142
rect 674 -2143 857 -2142
rect 1052 -2143 1459 -2142
rect 1584 -2143 1592 -2142
rect 1598 -2143 1683 -2142
rect 1787 -2143 2397 -2142
rect 121 -2145 451 -2144
rect 527 -2145 577 -2144
rect 709 -2145 780 -2144
rect 821 -2145 1452 -2144
rect 1556 -2145 1592 -2144
rect 1605 -2145 1676 -2144
rect 1682 -2145 1830 -2144
rect 2396 -2145 2411 -2144
rect 135 -2147 528 -2146
rect 534 -2147 1340 -2146
rect 1507 -2147 1676 -2146
rect 2102 -2147 2411 -2146
rect 254 -2149 675 -2148
rect 716 -2149 787 -2148
rect 842 -2149 948 -2148
rect 1052 -2149 1739 -2148
rect 2053 -2149 2103 -2148
rect 257 -2151 822 -2150
rect 1185 -2151 2040 -2150
rect 268 -2153 640 -2152
rect 723 -2153 836 -2152
rect 1185 -2153 2243 -2152
rect 268 -2155 1368 -2154
rect 1374 -2155 1508 -2154
rect 1556 -2155 1718 -2154
rect 2200 -2155 2243 -2154
rect 408 -2157 416 -2156
rect 478 -2157 710 -2156
rect 730 -2157 878 -2156
rect 1230 -2157 1739 -2156
rect 2158 -2157 2201 -2156
rect 233 -2159 479 -2158
rect 513 -2159 724 -2158
rect 747 -2159 934 -2158
rect 1255 -2159 1375 -2158
rect 1647 -2159 2054 -2158
rect 282 -2161 514 -2160
rect 520 -2161 717 -2160
rect 765 -2161 1480 -2160
rect 1647 -2161 2278 -2160
rect 282 -2163 325 -2162
rect 359 -2163 521 -2162
rect 765 -2163 773 -2162
rect 814 -2163 843 -2162
rect 877 -2163 1662 -2162
rect 1668 -2163 1830 -2162
rect 1892 -2163 2159 -2162
rect 324 -2165 430 -2164
rect 667 -2165 815 -2164
rect 1346 -2165 1669 -2164
rect 1717 -2165 1858 -2164
rect 359 -2167 486 -2166
rect 499 -2167 668 -2166
rect 772 -2167 913 -2166
rect 1346 -2167 1389 -2166
rect 1496 -2167 2278 -2166
rect 198 -2169 486 -2168
rect 737 -2169 1389 -2168
rect 1514 -2169 1662 -2168
rect 1836 -2169 1893 -2168
rect 184 -2171 199 -2170
rect 380 -2171 416 -2170
rect 429 -2171 745 -2170
rect 912 -2171 1578 -2170
rect 1836 -2171 2320 -2170
rect 121 -2173 381 -2172
rect 737 -2173 1490 -2172
rect 184 -2175 244 -2174
rect 1220 -2175 1515 -2174
rect 2 -2186 675 -2185
rect 744 -2186 1235 -2185
rect 1258 -2186 2313 -2185
rect 2343 -2186 2397 -2185
rect 9 -2188 52 -2187
rect 54 -2188 1389 -2187
rect 1398 -2188 1886 -2187
rect 1937 -2188 2299 -2187
rect 37 -2190 997 -2189
rect 1038 -2190 1224 -2189
rect 1227 -2190 2306 -2189
rect 51 -2192 1032 -2191
rect 1080 -2192 1151 -2191
rect 1157 -2192 1389 -2191
rect 1405 -2192 1438 -2191
rect 1489 -2192 2404 -2191
rect 65 -2194 1042 -2193
rect 1080 -2194 1102 -2193
rect 1115 -2194 1140 -2193
rect 1143 -2194 1235 -2193
rect 1293 -2194 1984 -2193
rect 2151 -2194 2306 -2193
rect 65 -2196 1277 -2195
rect 1304 -2196 1928 -2195
rect 1969 -2196 2299 -2195
rect 93 -2198 1480 -2197
rect 1496 -2198 1753 -2197
rect 1780 -2198 1784 -2197
rect 1836 -2198 1872 -2197
rect 1885 -2198 1963 -2197
rect 1969 -2198 2033 -2197
rect 2151 -2198 2271 -2197
rect 93 -2200 1361 -2199
rect 1367 -2200 2173 -2199
rect 2228 -2200 2337 -2199
rect 96 -2202 927 -2201
rect 936 -2202 1011 -2201
rect 1031 -2202 1046 -2201
rect 1094 -2202 1158 -2201
rect 1192 -2202 1256 -2201
rect 1304 -2202 1417 -2201
rect 1437 -2202 1515 -2201
rect 1521 -2202 1753 -2201
rect 1780 -2202 1844 -2201
rect 1860 -2202 2369 -2201
rect 107 -2204 129 -2203
rect 131 -2204 258 -2203
rect 296 -2204 657 -2203
rect 674 -2204 1896 -2203
rect 1927 -2204 1991 -2203
rect 2032 -2204 2103 -2203
rect 107 -2206 507 -2205
rect 527 -2206 1385 -2205
rect 1416 -2206 1494 -2205
rect 1521 -2206 1627 -2205
rect 1629 -2206 2250 -2205
rect 121 -2208 1711 -2207
rect 1843 -2208 1907 -2207
rect 1962 -2208 2026 -2207
rect 2060 -2208 2229 -2207
rect 16 -2210 122 -2209
rect 124 -2210 388 -2209
rect 450 -2210 496 -2209
rect 506 -2210 780 -2209
rect 782 -2210 993 -2209
rect 996 -2210 1942 -2209
rect 1983 -2210 2047 -2209
rect 2060 -2210 2131 -2209
rect 16 -2212 87 -2211
rect 128 -2212 1189 -2211
rect 1192 -2212 1270 -2211
rect 1332 -2212 1347 -2211
rect 1367 -2212 1536 -2211
rect 1545 -2212 2348 -2211
rect 86 -2214 626 -2213
rect 681 -2214 745 -2213
rect 800 -2214 1186 -2213
rect 1202 -2214 1277 -2213
rect 1283 -2214 1347 -2213
rect 1381 -2214 1550 -2213
rect 1580 -2214 2117 -2213
rect 2130 -2214 2257 -2213
rect 138 -2216 2264 -2215
rect 145 -2218 857 -2217
rect 877 -2218 1504 -2217
rect 1517 -2218 2348 -2217
rect 166 -2220 2208 -2219
rect 2256 -2220 2355 -2219
rect 236 -2222 941 -2221
rect 975 -2222 1760 -2221
rect 1783 -2222 1907 -2221
rect 1941 -2222 1998 -2221
rect 2025 -2222 2089 -2221
rect 2102 -2222 2201 -2221
rect 2207 -2222 2341 -2221
rect 243 -2224 885 -2223
rect 912 -2224 1011 -2223
rect 1094 -2224 1172 -2223
rect 1185 -2224 1263 -2223
rect 1269 -2224 1291 -2223
rect 1342 -2224 1431 -2223
rect 1479 -2224 1788 -2223
rect 1871 -2224 1949 -2223
rect 1990 -2224 2054 -2223
rect 2088 -2224 2166 -2223
rect 2200 -2224 2334 -2223
rect 156 -2226 1172 -2225
rect 1220 -2226 2285 -2225
rect 40 -2228 157 -2227
rect 250 -2228 1221 -2227
rect 1227 -2228 1452 -2227
rect 1535 -2228 1669 -2227
rect 1759 -2228 1816 -2227
rect 1934 -2228 2166 -2227
rect 2186 -2228 2285 -2227
rect 289 -2230 780 -2229
rect 821 -2230 927 -2229
rect 940 -2230 955 -2229
rect 975 -2230 1980 -2229
rect 1997 -2230 2068 -2229
rect 2116 -2230 2222 -2229
rect 289 -2232 353 -2231
rect 359 -2232 1056 -2231
rect 1101 -2232 1130 -2231
rect 1136 -2232 1333 -2231
rect 1381 -2232 1466 -2231
rect 1549 -2232 1592 -2231
rect 1647 -2232 2264 -2231
rect 261 -2234 360 -2233
rect 457 -2234 517 -2233
rect 527 -2234 584 -2233
rect 590 -2234 955 -2233
rect 978 -2234 2313 -2233
rect 100 -2236 262 -2235
rect 296 -2236 605 -2235
rect 618 -2236 668 -2235
rect 681 -2236 710 -2235
rect 726 -2236 2173 -2235
rect 2186 -2236 2418 -2235
rect 100 -2238 1018 -2237
rect 1115 -2238 1697 -2237
rect 1787 -2238 1851 -2237
rect 1934 -2238 2180 -2237
rect 2221 -2238 2320 -2237
rect 170 -2240 458 -2239
rect 492 -2240 1074 -2239
rect 1129 -2240 1165 -2239
rect 1248 -2240 1361 -2239
rect 1423 -2240 1452 -2239
rect 1465 -2240 1571 -2239
rect 1591 -2240 1690 -2239
rect 1703 -2240 1851 -2239
rect 1948 -2240 2005 -2239
rect 2046 -2240 2334 -2239
rect 79 -2242 493 -2241
rect 555 -2242 1231 -2241
rect 1248 -2242 2271 -2241
rect 79 -2244 640 -2243
rect 653 -2244 1137 -2243
rect 1143 -2244 1207 -2243
rect 1255 -2244 1375 -2243
rect 1423 -2244 1515 -2243
rect 1570 -2244 1662 -2243
rect 1682 -2244 1816 -2243
rect 1857 -2244 2005 -2243
rect 2053 -2244 2124 -2243
rect 2179 -2244 2292 -2243
rect 170 -2246 178 -2245
rect 338 -2246 451 -2245
rect 576 -2246 619 -2245
rect 621 -2246 1578 -2245
rect 1605 -2246 1690 -2245
rect 1703 -2246 1767 -2245
rect 1857 -2246 1921 -2245
rect 2067 -2246 2138 -2245
rect 177 -2248 1686 -2247
rect 1766 -2248 1823 -2247
rect 2123 -2248 2236 -2247
rect 317 -2250 339 -2249
rect 352 -2250 367 -2249
rect 394 -2250 556 -2249
rect 583 -2250 598 -2249
rect 604 -2250 696 -2249
rect 709 -2250 920 -2249
rect 978 -2250 2292 -2249
rect 275 -2252 598 -2251
rect 639 -2252 892 -2251
rect 912 -2252 990 -2251
rect 1073 -2252 1123 -2251
rect 1164 -2252 1242 -2251
rect 1262 -2252 1396 -2251
rect 1430 -2252 1501 -2251
rect 1605 -2252 1641 -2251
rect 1647 -2252 1809 -2251
rect 2074 -2252 2236 -2251
rect 275 -2254 626 -2253
rect 688 -2254 822 -2253
rect 828 -2254 885 -2253
rect 982 -2254 1046 -2253
rect 1087 -2254 1123 -2253
rect 1178 -2254 1242 -2253
rect 1283 -2254 1319 -2253
rect 1339 -2254 1823 -2253
rect 2018 -2254 2075 -2253
rect 310 -2256 318 -2255
rect 324 -2256 395 -2255
rect 443 -2256 892 -2255
rect 961 -2256 1088 -2255
rect 1178 -2256 1445 -2255
rect 1486 -2256 1921 -2255
rect 2018 -2256 2362 -2255
rect 114 -2258 325 -2257
rect 366 -2258 664 -2257
rect 695 -2258 1308 -2257
rect 1318 -2258 2411 -2257
rect 114 -2260 227 -2259
rect 310 -2260 542 -2259
rect 590 -2260 871 -2259
rect 933 -2260 962 -2259
rect 989 -2260 2425 -2259
rect 163 -2262 227 -2261
rect 380 -2262 689 -2261
rect 751 -2262 1018 -2261
rect 1206 -2262 1298 -2261
rect 1339 -2262 1459 -2261
rect 1472 -2262 1487 -2261
rect 1500 -2262 2383 -2261
rect 163 -2264 2250 -2263
rect 380 -2266 836 -2265
rect 856 -2266 1977 -2265
rect 443 -2268 472 -2267
rect 478 -2268 577 -2267
rect 593 -2268 2040 -2267
rect 142 -2270 472 -2269
rect 478 -2270 920 -2269
rect 1290 -2270 1914 -2269
rect 2039 -2270 2110 -2269
rect 142 -2272 255 -2271
rect 513 -2272 871 -2271
rect 1297 -2272 1354 -2271
rect 1370 -2272 1459 -2271
rect 1472 -2272 1956 -2271
rect 2109 -2272 2215 -2271
rect 513 -2274 535 -2273
rect 541 -2274 549 -2273
rect 737 -2274 752 -2273
rect 758 -2274 1669 -2273
rect 1808 -2274 2012 -2273
rect 2095 -2274 2215 -2273
rect 422 -2276 535 -2275
rect 548 -2276 717 -2275
rect 758 -2276 864 -2275
rect 1353 -2276 1529 -2275
rect 1563 -2276 1956 -2275
rect 2011 -2276 2082 -2275
rect 2095 -2276 2194 -2275
rect 184 -2278 717 -2277
rect 765 -2278 878 -2277
rect 1059 -2278 1529 -2277
rect 1563 -2278 1655 -2277
rect 1661 -2278 1739 -2277
rect 1892 -2278 1914 -2277
rect 2081 -2278 2159 -2277
rect 149 -2280 185 -2279
rect 219 -2280 423 -2279
rect 485 -2280 738 -2279
rect 772 -2280 801 -2279
rect 814 -2280 864 -2279
rect 1059 -2280 1336 -2279
rect 1374 -2280 1543 -2279
rect 1619 -2280 1697 -2279
rect 1738 -2280 1795 -2279
rect 135 -2282 150 -2281
rect 191 -2282 220 -2281
rect 373 -2282 766 -2281
rect 786 -2282 2320 -2281
rect 135 -2284 570 -2283
rect 611 -2284 815 -2283
rect 828 -2284 843 -2283
rect 859 -2284 2138 -2283
rect 191 -2286 1067 -2285
rect 1321 -2286 2194 -2285
rect 373 -2288 521 -2287
rect 569 -2288 724 -2287
rect 786 -2288 1004 -2287
rect 1066 -2288 1109 -2287
rect 1395 -2288 1977 -2287
rect 415 -2290 521 -2289
rect 646 -2290 773 -2289
rect 807 -2290 843 -2289
rect 968 -2290 1543 -2289
rect 1619 -2290 1718 -2289
rect 1794 -2290 1865 -2289
rect 331 -2292 416 -2291
rect 436 -2292 486 -2291
rect 499 -2292 612 -2291
rect 646 -2292 661 -2291
rect 723 -2292 983 -2291
rect 1052 -2292 1109 -2291
rect 1402 -2292 2159 -2291
rect 233 -2294 500 -2293
rect 562 -2294 1403 -2293
rect 1409 -2294 1865 -2293
rect 233 -2296 706 -2295
rect 730 -2296 1053 -2295
rect 1409 -2296 1627 -2295
rect 1633 -2296 1718 -2295
rect 268 -2298 437 -2297
rect 730 -2298 899 -2297
rect 905 -2298 969 -2297
rect 1444 -2298 1585 -2297
rect 1633 -2298 1725 -2297
rect 205 -2300 899 -2299
rect 905 -2300 1326 -2299
rect 1584 -2300 1676 -2299
rect 44 -2302 206 -2301
rect 212 -2302 269 -2301
rect 331 -2302 346 -2301
rect 429 -2302 563 -2301
rect 747 -2302 1004 -2301
rect 1024 -2302 1725 -2301
rect 44 -2304 59 -2303
rect 72 -2304 1025 -2303
rect 1325 -2304 1613 -2303
rect 1640 -2304 1732 -2303
rect 23 -2306 59 -2305
rect 72 -2306 402 -2305
rect 807 -2306 850 -2305
rect 1507 -2306 1613 -2305
rect 1650 -2306 2327 -2305
rect 23 -2308 199 -2307
rect 212 -2308 248 -2307
rect 282 -2308 346 -2307
rect 401 -2308 465 -2307
rect 835 -2308 1214 -2307
rect 1507 -2308 1557 -2307
rect 1675 -2308 1746 -2307
rect 2277 -2308 2327 -2307
rect 198 -2310 671 -2309
rect 793 -2310 1214 -2309
rect 1556 -2310 1599 -2309
rect 1731 -2310 2145 -2309
rect 2277 -2310 2390 -2309
rect 247 -2312 430 -2311
rect 464 -2312 633 -2311
rect 789 -2312 1599 -2311
rect 1745 -2312 1802 -2311
rect 2144 -2312 2243 -2311
rect 282 -2314 304 -2313
rect 387 -2314 671 -2313
rect 793 -2314 1494 -2313
rect 1801 -2314 1879 -2313
rect 2242 -2314 2376 -2313
rect 303 -2316 409 -2315
rect 632 -2316 703 -2315
rect 849 -2316 1312 -2315
rect 1773 -2316 1879 -2315
rect 30 -2318 409 -2317
rect 660 -2318 1312 -2317
rect 1773 -2318 1830 -2317
rect 702 -2320 1655 -2319
rect 1829 -2320 1900 -2319
rect 1199 -2322 1900 -2321
rect 33 -2324 1200 -2323
rect 5 -2335 66 -2334
rect 163 -2335 1025 -2334
rect 1038 -2335 1361 -2334
rect 1363 -2335 2222 -2334
rect 2326 -2335 2344 -2334
rect 9 -2337 874 -2336
rect 905 -2337 1249 -2336
rect 1272 -2337 2075 -2336
rect 2165 -2337 2334 -2336
rect 23 -2339 146 -2338
rect 170 -2339 174 -2338
rect 226 -2339 594 -2338
rect 597 -2339 727 -2338
rect 782 -2339 1536 -2338
rect 1542 -2339 1879 -2338
rect 1892 -2339 1949 -2338
rect 1976 -2339 2040 -2338
rect 2165 -2339 2194 -2338
rect 2221 -2339 2243 -2338
rect 16 -2341 227 -2340
rect 240 -2341 608 -2340
rect 618 -2341 1319 -2340
rect 1374 -2341 1396 -2340
rect 1398 -2341 1410 -2340
rect 1493 -2341 2236 -2340
rect 2242 -2341 2292 -2340
rect 16 -2343 38 -2342
rect 51 -2343 1025 -2342
rect 1041 -2343 1494 -2342
rect 1517 -2343 1907 -2342
rect 1934 -2343 2285 -2342
rect 30 -2345 1081 -2344
rect 1108 -2345 1980 -2344
rect 2039 -2345 2089 -2344
rect 2186 -2345 2292 -2344
rect 33 -2347 45 -2346
rect 51 -2347 1578 -2346
rect 1580 -2347 2257 -2346
rect 44 -2349 115 -2348
rect 170 -2349 178 -2348
rect 243 -2349 507 -2348
rect 569 -2349 619 -2348
rect 625 -2349 892 -2348
rect 905 -2349 941 -2348
rect 954 -2349 1322 -2348
rect 1377 -2349 1452 -2348
rect 1542 -2349 1599 -2348
rect 1682 -2349 2229 -2348
rect 2235 -2349 2278 -2348
rect 65 -2351 276 -2350
rect 282 -2351 1077 -2350
rect 1080 -2351 1613 -2350
rect 1682 -2351 1746 -2350
rect 1850 -2351 1854 -2350
rect 1878 -2351 2103 -2350
rect 2179 -2351 2187 -2350
rect 2193 -2351 2208 -2350
rect 2228 -2351 2264 -2350
rect 114 -2353 262 -2352
rect 275 -2353 388 -2352
rect 408 -2353 766 -2352
rect 775 -2353 941 -2352
rect 978 -2353 1214 -2352
rect 1248 -2353 1263 -2352
rect 1276 -2353 1357 -2352
rect 1451 -2353 1529 -2352
rect 1685 -2353 2159 -2352
rect 2207 -2353 2281 -2352
rect 166 -2355 2180 -2354
rect 2256 -2355 2313 -2354
rect 247 -2357 843 -2356
rect 859 -2357 1613 -2356
rect 1745 -2357 1774 -2356
rect 1850 -2357 1886 -2356
rect 1895 -2357 2215 -2356
rect 2263 -2357 2320 -2356
rect 247 -2359 479 -2358
rect 481 -2359 1630 -2358
rect 1773 -2359 1788 -2358
rect 1885 -2359 1942 -2358
rect 1948 -2359 2117 -2358
rect 261 -2361 402 -2360
rect 408 -2361 486 -2360
rect 492 -2361 507 -2360
rect 527 -2361 570 -2360
rect 576 -2361 780 -2360
rect 786 -2361 955 -2360
rect 982 -2361 1039 -2360
rect 1055 -2361 1487 -2360
rect 1528 -2361 1592 -2360
rect 1787 -2361 1844 -2360
rect 1853 -2361 1942 -2360
rect 2011 -2361 2117 -2360
rect 282 -2363 836 -2362
rect 842 -2363 913 -2362
rect 919 -2363 1697 -2362
rect 1843 -2363 1858 -2362
rect 1906 -2363 1928 -2362
rect 1934 -2363 1998 -2362
rect 2011 -2363 2068 -2362
rect 2088 -2363 2306 -2362
rect 296 -2365 724 -2364
rect 730 -2365 1410 -2364
rect 1486 -2365 1571 -2364
rect 1591 -2365 1823 -2364
rect 1836 -2365 1858 -2364
rect 1927 -2365 1991 -2364
rect 1997 -2365 2061 -2364
rect 2102 -2365 2131 -2364
rect 2305 -2365 2348 -2364
rect 191 -2367 724 -2366
rect 730 -2367 794 -2366
rect 796 -2367 1669 -2366
rect 1678 -2367 1697 -2366
rect 1836 -2367 1984 -2366
rect 1990 -2367 2124 -2366
rect 72 -2369 192 -2368
rect 296 -2369 1053 -2368
rect 1108 -2369 1151 -2368
rect 1262 -2369 1305 -2368
rect 1318 -2369 1382 -2368
rect 1668 -2369 1739 -2368
rect 1983 -2369 2054 -2368
rect 2060 -2369 2110 -2368
rect 2123 -2369 2138 -2368
rect 310 -2371 430 -2370
rect 457 -2371 857 -2370
rect 859 -2371 1333 -2370
rect 1381 -2371 1438 -2370
rect 1738 -2371 1767 -2370
rect 1969 -2371 2110 -2370
rect 2137 -2371 2152 -2370
rect 268 -2373 311 -2372
rect 387 -2373 857 -2372
rect 863 -2373 983 -2372
rect 1052 -2373 2075 -2372
rect 2151 -2373 2173 -2372
rect 401 -2375 682 -2374
rect 716 -2375 2068 -2374
rect 2172 -2375 2201 -2374
rect 37 -2377 2201 -2376
rect 100 -2379 717 -2378
rect 786 -2379 1165 -2378
rect 1227 -2379 1305 -2378
rect 1437 -2379 1445 -2378
rect 1766 -2379 1830 -2378
rect 2018 -2379 2215 -2378
rect 100 -2381 962 -2380
rect 1087 -2381 1165 -2380
rect 1227 -2381 1256 -2380
rect 1276 -2381 1546 -2380
rect 1647 -2381 1830 -2380
rect 2046 -2381 2285 -2380
rect 422 -2383 769 -2382
rect 821 -2383 979 -2382
rect 1087 -2383 1130 -2382
rect 1136 -2383 1298 -2382
rect 1444 -2383 1480 -2382
rect 1549 -2383 1648 -2382
rect 1801 -2383 1970 -2382
rect 2053 -2383 2096 -2382
rect 110 -2385 1137 -2384
rect 1150 -2385 1186 -2384
rect 1293 -2385 1753 -2384
rect 1899 -2385 2096 -2384
rect 324 -2387 423 -2386
rect 457 -2387 647 -2386
rect 660 -2387 759 -2386
rect 821 -2387 878 -2386
rect 884 -2387 892 -2386
rect 912 -2387 1336 -2386
rect 1479 -2387 1704 -2386
rect 1752 -2387 1781 -2386
rect 1801 -2387 1900 -2386
rect 324 -2389 395 -2388
rect 464 -2389 486 -2388
rect 492 -2389 1312 -2388
rect 1465 -2389 1781 -2388
rect 303 -2391 395 -2390
rect 464 -2391 1018 -2390
rect 1115 -2391 1536 -2390
rect 1703 -2391 1718 -2390
rect 303 -2393 332 -2392
rect 520 -2393 682 -2392
rect 702 -2393 1186 -2392
rect 1311 -2393 1340 -2392
rect 1710 -2393 1718 -2392
rect 331 -2395 353 -2394
rect 380 -2395 521 -2394
rect 527 -2395 1252 -2394
rect 1339 -2395 1389 -2394
rect 1598 -2395 1711 -2394
rect 345 -2397 353 -2396
rect 380 -2397 437 -2396
rect 499 -2397 703 -2396
rect 758 -2397 1060 -2396
rect 1115 -2397 1193 -2396
rect 1367 -2397 1389 -2396
rect 219 -2399 346 -2398
rect 436 -2399 472 -2398
rect 499 -2399 535 -2398
rect 576 -2399 741 -2398
rect 814 -2399 1060 -2398
rect 1129 -2399 1403 -2398
rect 149 -2401 220 -2400
rect 233 -2401 535 -2400
rect 590 -2401 612 -2400
rect 621 -2401 2131 -2400
rect 149 -2403 164 -2402
rect 233 -2403 451 -2402
rect 597 -2403 1032 -2402
rect 1171 -2403 1466 -2402
rect 359 -2405 451 -2404
rect 611 -2405 633 -2404
rect 646 -2405 738 -2404
rect 814 -2405 871 -2404
rect 884 -2405 1375 -2404
rect 198 -2407 360 -2406
rect 443 -2407 472 -2406
rect 478 -2407 871 -2406
rect 919 -2407 2250 -2406
rect 184 -2409 199 -2408
rect 443 -2409 605 -2408
rect 628 -2409 801 -2408
rect 828 -2409 878 -2408
rect 922 -2409 2313 -2408
rect 135 -2411 605 -2410
rect 632 -2411 710 -2410
rect 737 -2411 1515 -2410
rect 135 -2413 416 -2412
rect 660 -2413 990 -2412
rect 1013 -2413 1403 -2412
rect 184 -2415 640 -2414
rect 670 -2415 2271 -2414
rect 268 -2417 671 -2416
rect 800 -2417 808 -2416
rect 828 -2417 899 -2416
rect 922 -2417 1725 -2416
rect 2270 -2417 2299 -2416
rect 366 -2419 710 -2418
rect 835 -2419 1004 -2418
rect 1017 -2419 1158 -2418
rect 1171 -2419 1914 -2418
rect 121 -2421 1004 -2420
rect 1031 -2421 1732 -2420
rect 1808 -2421 1914 -2420
rect 121 -2423 668 -2422
rect 863 -2423 948 -2422
rect 957 -2423 1158 -2422
rect 1174 -2423 1298 -2422
rect 1332 -2423 2299 -2422
rect 107 -2425 668 -2424
rect 898 -2425 969 -2424
rect 975 -2425 1550 -2424
rect 1633 -2425 1809 -2424
rect 107 -2427 129 -2426
rect 156 -2427 367 -2426
rect 415 -2427 514 -2426
rect 555 -2427 808 -2426
rect 933 -2427 2159 -2426
rect 79 -2429 556 -2428
rect 639 -2429 745 -2428
rect 936 -2429 1627 -2428
rect 1724 -2429 1938 -2428
rect 2 -2431 80 -2430
rect 86 -2431 934 -2430
rect 947 -2431 1067 -2430
rect 1139 -2431 2250 -2430
rect 2 -2433 73 -2432
rect 86 -2433 1501 -2432
rect 1507 -2433 1634 -2432
rect 1731 -2433 1865 -2432
rect 128 -2435 549 -2434
rect 695 -2435 745 -2434
rect 961 -2435 1123 -2434
rect 1178 -2435 1256 -2434
rect 1346 -2435 1865 -2434
rect 96 -2437 1179 -2436
rect 1192 -2437 1326 -2436
rect 1346 -2437 1424 -2436
rect 1500 -2437 1585 -2436
rect 1605 -2437 1627 -2436
rect 58 -2439 97 -2438
rect 156 -2439 213 -2438
rect 513 -2439 563 -2438
rect 688 -2439 696 -2438
rect 968 -2439 1011 -2438
rect 1066 -2439 1144 -2438
rect 1213 -2439 1606 -2438
rect 58 -2441 997 -2440
rect 1010 -2441 1102 -2440
rect 1122 -2441 1207 -2440
rect 1325 -2441 1497 -2440
rect 1507 -2441 1557 -2440
rect 1584 -2441 1655 -2440
rect 142 -2443 563 -2442
rect 793 -2443 1102 -2442
rect 1143 -2443 1522 -2442
rect 1556 -2443 1620 -2442
rect 93 -2445 143 -2444
rect 205 -2445 689 -2444
rect 975 -2445 2019 -2444
rect 93 -2447 1823 -2446
rect 205 -2449 675 -2448
rect 996 -2449 1046 -2448
rect 1206 -2449 1235 -2448
rect 1353 -2449 1424 -2448
rect 1458 -2449 1620 -2448
rect 212 -2451 290 -2450
rect 548 -2451 1805 -2450
rect 289 -2453 339 -2452
rect 674 -2453 993 -2452
rect 1045 -2453 1095 -2452
rect 1234 -2453 2337 -2452
rect 338 -2455 542 -2454
rect 926 -2455 1095 -2454
rect 1353 -2455 2145 -2454
rect 541 -2457 850 -2456
rect 992 -2457 2047 -2456
rect 772 -2459 927 -2458
rect 1199 -2459 2145 -2458
rect 23 -2461 773 -2460
rect 849 -2461 1291 -2460
rect 1367 -2461 1431 -2460
rect 1458 -2461 1578 -2460
rect 1199 -2463 1284 -2462
rect 1430 -2463 1641 -2462
rect 1283 -2465 1417 -2464
rect 1521 -2465 1662 -2464
rect 373 -2467 1662 -2466
rect 373 -2469 584 -2468
rect 1416 -2469 1473 -2468
rect 1563 -2469 1655 -2468
rect 583 -2471 654 -2470
rect 1472 -2471 1602 -2470
rect 1640 -2471 1816 -2470
rect 653 -2473 752 -2472
rect 1563 -2473 1690 -2472
rect 1815 -2473 1872 -2472
rect 751 -2475 1074 -2474
rect 1689 -2475 1760 -2474
rect 1871 -2475 1921 -2474
rect 1073 -2477 1956 -2476
rect 1759 -2479 1795 -2478
rect 1920 -2479 1963 -2478
rect 1675 -2481 1795 -2480
rect 1955 -2481 2005 -2480
rect 1962 -2483 2026 -2482
rect 1083 -2485 2026 -2484
rect 2004 -2487 2033 -2486
rect 2032 -2489 2082 -2488
rect 1220 -2491 2082 -2490
rect 1220 -2493 1242 -2492
rect 1241 -2495 1270 -2494
rect 1269 -2497 1571 -2496
rect 5 -2508 416 -2507
rect 464 -2508 990 -2507
rect 992 -2508 1074 -2507
rect 1080 -2508 1795 -2507
rect 1801 -2508 1935 -2507
rect 2088 -2508 2092 -2507
rect 9 -2510 1410 -2509
rect 1510 -2510 2054 -2509
rect 2088 -2510 2159 -2509
rect 9 -2512 52 -2511
rect 54 -2512 766 -2511
rect 775 -2512 878 -2511
rect 926 -2512 1084 -2511
rect 1188 -2512 1697 -2511
rect 1794 -2512 1886 -2511
rect 1934 -2512 2026 -2511
rect 2053 -2512 2131 -2511
rect 16 -2514 38 -2513
rect 40 -2514 1249 -2513
rect 1290 -2514 1809 -2513
rect 1885 -2514 1998 -2513
rect 2025 -2514 2103 -2513
rect 2130 -2514 2194 -2513
rect 33 -2516 934 -2515
rect 950 -2516 1291 -2515
rect 1335 -2516 2110 -2515
rect 37 -2518 52 -2517
rect 58 -2518 1466 -2517
rect 1580 -2518 1648 -2517
rect 1678 -2518 1970 -2517
rect 1997 -2518 2061 -2517
rect 2102 -2518 2243 -2517
rect 44 -2520 76 -2519
rect 93 -2520 1151 -2519
rect 1195 -2520 1907 -2519
rect 1969 -2520 2033 -2519
rect 2109 -2520 2173 -2519
rect 2242 -2520 2292 -2519
rect 44 -2522 528 -2521
rect 541 -2522 979 -2521
rect 989 -2522 1175 -2521
rect 1199 -2522 1333 -2521
rect 1356 -2522 1697 -2521
rect 1804 -2522 2187 -2521
rect 58 -2524 62 -2523
rect 72 -2524 1238 -2523
rect 1332 -2524 1417 -2523
rect 1458 -2524 2033 -2523
rect 2172 -2524 2236 -2523
rect 72 -2526 367 -2525
rect 373 -2526 790 -2525
rect 817 -2526 2061 -2525
rect 2186 -2526 2257 -2525
rect 93 -2528 115 -2527
rect 128 -2528 811 -2527
rect 859 -2528 1676 -2527
rect 1808 -2528 1872 -2527
rect 2235 -2528 2285 -2527
rect 107 -2530 262 -2529
rect 268 -2530 871 -2529
rect 877 -2530 1312 -2529
rect 1360 -2530 2117 -2529
rect 110 -2532 1361 -2531
rect 1374 -2532 1942 -2531
rect 2116 -2532 2124 -2531
rect 131 -2534 969 -2533
rect 1006 -2534 1032 -2533
rect 1038 -2534 1151 -2533
rect 1216 -2534 2271 -2533
rect 19 -2536 1032 -2535
rect 1038 -2536 1158 -2535
rect 1311 -2536 1844 -2535
rect 1871 -2536 1928 -2535
rect 1941 -2536 2166 -2535
rect 2270 -2536 2313 -2535
rect 149 -2538 269 -2537
rect 275 -2538 794 -2537
rect 898 -2538 934 -2537
rect 940 -2538 1200 -2537
rect 1377 -2538 1655 -2537
rect 1843 -2538 1900 -2537
rect 2123 -2538 2180 -2537
rect 103 -2540 899 -2539
rect 919 -2540 969 -2539
rect 1010 -2540 1123 -2539
rect 1402 -2540 1406 -2539
rect 1416 -2540 1438 -2539
rect 1458 -2540 1515 -2539
rect 1580 -2540 2005 -2539
rect 2165 -2540 2229 -2539
rect 128 -2542 941 -2541
rect 1013 -2542 1375 -2541
rect 1402 -2542 1445 -2541
rect 1465 -2542 1543 -2541
rect 1601 -2542 2096 -2541
rect 2179 -2542 2250 -2541
rect 149 -2544 430 -2543
rect 478 -2544 1662 -2543
rect 1766 -2544 2229 -2543
rect 163 -2546 178 -2545
rect 191 -2546 262 -2545
rect 303 -2546 412 -2545
rect 429 -2546 1441 -2545
rect 1444 -2546 1620 -2545
rect 1647 -2546 1711 -2545
rect 1899 -2546 1963 -2545
rect 163 -2548 1354 -2547
rect 1437 -2548 1704 -2547
rect 1710 -2548 1921 -2547
rect 96 -2550 1354 -2549
rect 1500 -2550 1515 -2549
rect 1542 -2550 1564 -2549
rect 1612 -2550 1928 -2549
rect 177 -2552 584 -2551
rect 604 -2552 892 -2551
rect 894 -2552 1767 -2551
rect 1920 -2552 2012 -2551
rect 191 -2554 1578 -2553
rect 1619 -2554 1977 -2553
rect 201 -2556 608 -2555
rect 632 -2556 1214 -2555
rect 1272 -2556 1704 -2555
rect 1948 -2556 2012 -2555
rect 205 -2558 276 -2557
rect 310 -2558 1270 -2557
rect 1314 -2558 2096 -2557
rect 198 -2560 206 -2559
rect 240 -2560 542 -2559
rect 555 -2560 741 -2559
rect 751 -2560 773 -2559
rect 926 -2560 1298 -2559
rect 1451 -2560 1613 -2559
rect 1654 -2560 1756 -2559
rect 1948 -2560 2040 -2559
rect 198 -2562 612 -2561
rect 709 -2562 1053 -2561
rect 1066 -2562 1410 -2561
rect 1451 -2562 1571 -2561
rect 1661 -2562 1739 -2561
rect 1976 -2562 2047 -2561
rect 240 -2564 416 -2563
rect 457 -2564 612 -2563
rect 709 -2564 731 -2563
rect 737 -2564 2005 -2563
rect 2046 -2564 2208 -2563
rect 254 -2566 304 -2565
rect 310 -2566 423 -2565
rect 457 -2566 559 -2565
rect 562 -2566 766 -2565
rect 873 -2566 2040 -2565
rect 2091 -2566 2159 -2565
rect 135 -2568 255 -2567
rect 352 -2568 1011 -2567
rect 1017 -2568 2194 -2567
rect 135 -2570 248 -2569
rect 352 -2570 451 -2569
rect 492 -2570 1158 -2569
rect 1185 -2570 1963 -2569
rect 184 -2572 493 -2571
rect 562 -2572 864 -2571
rect 1017 -2572 1109 -2571
rect 1122 -2572 1424 -2571
rect 1479 -2572 1564 -2571
rect 1570 -2572 1606 -2571
rect 1738 -2572 1788 -2571
rect 142 -2574 864 -2573
rect 1052 -2574 1116 -2573
rect 1213 -2574 1326 -2573
rect 1423 -2574 1529 -2573
rect 1605 -2574 1683 -2573
rect 1787 -2574 1865 -2573
rect 142 -2576 892 -2575
rect 1066 -2576 1319 -2575
rect 1479 -2576 1487 -2575
rect 1500 -2576 1585 -2575
rect 1682 -2576 1760 -2575
rect 1850 -2576 1865 -2575
rect 184 -2578 976 -2577
rect 1073 -2578 1095 -2577
rect 1269 -2578 1389 -2577
rect 1486 -2578 1550 -2577
rect 1584 -2578 1627 -2577
rect 1731 -2578 1760 -2577
rect 1850 -2578 1956 -2577
rect 219 -2580 423 -2579
rect 450 -2580 829 -2579
rect 842 -2580 976 -2579
rect 1080 -2580 1088 -2579
rect 1094 -2580 1144 -2579
rect 1297 -2580 1396 -2579
rect 1528 -2580 1634 -2579
rect 1955 -2580 2019 -2579
rect 86 -2582 843 -2581
rect 1087 -2582 1382 -2581
rect 1388 -2582 1494 -2581
rect 1549 -2582 1746 -2581
rect 1990 -2582 2019 -2581
rect 86 -2584 923 -2583
rect 1143 -2584 1221 -2583
rect 1234 -2584 1382 -2583
rect 1395 -2584 1830 -2583
rect 1878 -2584 1991 -2583
rect 26 -2586 1879 -2585
rect 219 -2588 318 -2587
rect 359 -2588 1364 -2587
rect 1430 -2588 1494 -2587
rect 1591 -2588 1732 -2587
rect 1745 -2588 1816 -2587
rect 1829 -2588 1837 -2587
rect 212 -2590 318 -2589
rect 331 -2590 360 -2589
rect 366 -2590 507 -2589
rect 569 -2590 633 -2589
rect 646 -2590 1186 -2589
rect 1220 -2590 1340 -2589
rect 1430 -2590 1599 -2589
rect 1626 -2590 1690 -2589
rect 1815 -2590 1858 -2589
rect 212 -2592 598 -2591
rect 646 -2592 689 -2591
rect 716 -2592 794 -2591
rect 828 -2592 1305 -2591
rect 1318 -2592 1536 -2591
rect 1591 -2592 1774 -2591
rect 1836 -2592 1893 -2591
rect 68 -2594 689 -2593
rect 716 -2594 1207 -2593
rect 1234 -2594 1263 -2593
rect 1339 -2594 1399 -2593
rect 1472 -2594 1536 -2593
rect 1598 -2594 1669 -2593
rect 1773 -2594 1823 -2593
rect 1857 -2594 2075 -2593
rect 226 -2596 248 -2595
rect 282 -2596 1116 -2595
rect 1171 -2596 1893 -2595
rect 2074 -2596 2145 -2595
rect 170 -2598 227 -2597
rect 282 -2598 671 -2597
rect 723 -2598 738 -2597
rect 751 -2598 1126 -2597
rect 1171 -2598 1256 -2597
rect 1262 -2598 1347 -2597
rect 1412 -2598 1473 -2597
rect 1633 -2598 2281 -2597
rect 166 -2600 171 -2599
rect 331 -2600 346 -2599
rect 373 -2600 395 -2599
rect 401 -2600 857 -2599
rect 954 -2600 1347 -2599
rect 1640 -2600 1690 -2599
rect 1822 -2600 1914 -2599
rect 2144 -2600 2215 -2599
rect 30 -2602 346 -2601
rect 380 -2602 528 -2601
rect 569 -2602 815 -2601
rect 824 -2602 1305 -2601
rect 1640 -2602 1725 -2601
rect 1913 -2602 1984 -2601
rect 2214 -2602 2264 -2601
rect 30 -2604 486 -2603
rect 506 -2604 850 -2603
rect 1178 -2604 1984 -2603
rect 2263 -2604 2306 -2603
rect 79 -2606 857 -2605
rect 1003 -2606 1179 -2605
rect 1206 -2606 1284 -2605
rect 1447 -2606 1725 -2605
rect 79 -2608 549 -2607
rect 583 -2608 801 -2607
rect 807 -2608 1004 -2607
rect 1255 -2608 1578 -2607
rect 1668 -2608 1753 -2607
rect 156 -2610 402 -2609
rect 408 -2610 465 -2609
rect 485 -2610 640 -2609
rect 726 -2610 2082 -2609
rect 156 -2612 556 -2611
rect 597 -2612 958 -2611
rect 1752 -2612 2299 -2611
rect 289 -2614 409 -2613
rect 520 -2614 955 -2613
rect 2081 -2614 2152 -2613
rect 65 -2616 290 -2615
rect 380 -2616 661 -2615
rect 730 -2616 983 -2615
rect 2151 -2616 2222 -2615
rect 65 -2618 2068 -2617
rect 387 -2620 479 -2619
rect 513 -2620 661 -2619
rect 758 -2620 1109 -2619
rect 2067 -2620 2138 -2619
rect 338 -2622 388 -2621
rect 394 -2622 1056 -2621
rect 2137 -2622 2201 -2621
rect 338 -2624 500 -2623
rect 513 -2624 696 -2623
rect 786 -2624 1284 -2623
rect 443 -2626 500 -2625
rect 520 -2626 577 -2625
rect 590 -2626 759 -2625
rect 800 -2626 1557 -2625
rect 233 -2628 444 -2627
rect 534 -2628 591 -2627
rect 618 -2628 815 -2627
rect 849 -2628 1102 -2627
rect 1507 -2628 1557 -2627
rect 233 -2630 675 -2629
rect 695 -2630 997 -2629
rect 1101 -2630 1137 -2629
rect 1248 -2630 1508 -2629
rect 324 -2632 535 -2631
rect 548 -2632 836 -2631
rect 982 -2632 1060 -2631
rect 1136 -2632 2222 -2631
rect 324 -2634 472 -2633
rect 576 -2634 787 -2633
rect 796 -2634 1060 -2633
rect 23 -2636 472 -2635
rect 618 -2636 885 -2635
rect 996 -2636 1046 -2635
rect 639 -2638 682 -2637
rect 779 -2638 836 -2637
rect 884 -2638 906 -2637
rect 1045 -2638 1277 -2637
rect 121 -2640 780 -2639
rect 1241 -2640 1277 -2639
rect 481 -2642 906 -2641
rect 1241 -2642 1781 -2641
rect 625 -2644 682 -2643
rect 1013 -2644 1781 -2643
rect 625 -2646 913 -2645
rect 667 -2648 2201 -2647
rect 667 -2650 703 -2649
rect 912 -2650 1130 -2649
rect 674 -2652 822 -2651
rect 1129 -2652 1165 -2651
rect 114 -2654 822 -2653
rect 1164 -2654 1228 -2653
rect 702 -2656 745 -2655
rect 1227 -2656 1368 -2655
rect 744 -2658 962 -2657
rect 1192 -2658 1368 -2657
rect 947 -2660 962 -2659
rect 1192 -2660 1907 -2659
rect 296 -2662 948 -2661
rect 296 -2664 437 -2663
rect 436 -2666 654 -2665
rect 100 -2668 654 -2667
rect 100 -2670 122 -2669
rect 2 -2681 69 -2680
rect 103 -2681 339 -2680
rect 432 -2681 465 -2680
rect 506 -2681 734 -2680
rect 758 -2681 839 -2680
rect 915 -2681 2047 -2680
rect 2224 -2681 2271 -2680
rect 16 -2683 251 -2682
rect 338 -2683 346 -2682
rect 506 -2683 780 -2682
rect 786 -2683 1151 -2682
rect 1185 -2683 1886 -2682
rect 1927 -2683 2260 -2682
rect 16 -2685 696 -2684
rect 709 -2685 958 -2684
rect 978 -2685 1284 -2684
rect 1286 -2685 1459 -2684
rect 1489 -2685 1592 -2684
rect 1619 -2685 1886 -2684
rect 23 -2687 136 -2686
rect 156 -2687 1056 -2686
rect 1062 -2687 1137 -2686
rect 1139 -2687 1480 -2686
rect 1577 -2687 2250 -2686
rect 23 -2689 521 -2688
rect 548 -2689 818 -2688
rect 821 -2689 934 -2688
rect 954 -2689 1144 -2688
rect 1185 -2689 1207 -2688
rect 1234 -2689 2005 -2688
rect 26 -2691 843 -2690
rect 919 -2691 1956 -2690
rect 65 -2693 87 -2692
rect 110 -2693 283 -2692
rect 345 -2693 360 -2692
rect 387 -2693 521 -2692
rect 555 -2693 633 -2692
rect 681 -2693 724 -2692
rect 765 -2693 951 -2692
rect 954 -2693 976 -2692
rect 1013 -2693 2103 -2692
rect 65 -2695 997 -2694
rect 1041 -2695 1872 -2694
rect 1955 -2695 1977 -2694
rect 2102 -2695 2138 -2694
rect 82 -2697 633 -2696
rect 681 -2697 717 -2696
rect 765 -2697 1221 -2696
rect 1234 -2697 1396 -2696
rect 1423 -2697 1459 -2696
rect 1479 -2697 1557 -2696
rect 1584 -2697 1686 -2696
rect 1755 -2697 2159 -2696
rect 86 -2699 1259 -2698
rect 1318 -2699 2271 -2698
rect 107 -2701 556 -2700
rect 558 -2701 661 -2700
rect 695 -2701 738 -2700
rect 772 -2701 892 -2700
rect 919 -2701 962 -2700
rect 975 -2701 1928 -2700
rect 1976 -2701 2019 -2700
rect 2130 -2701 2138 -2700
rect 2158 -2701 2173 -2700
rect 121 -2703 129 -2702
rect 163 -2703 549 -2702
rect 562 -2703 1039 -2702
rect 1066 -2703 1144 -2702
rect 1195 -2703 1445 -2702
rect 1556 -2703 1788 -2702
rect 1871 -2703 1907 -2702
rect 2011 -2703 2019 -2702
rect 2130 -2703 2145 -2702
rect 51 -2705 1445 -2704
rect 1584 -2705 1697 -2704
rect 1759 -2705 2005 -2704
rect 2144 -2705 2152 -2704
rect 51 -2707 983 -2706
rect 996 -2707 1214 -2706
rect 1220 -2707 1263 -2706
rect 1360 -2707 1592 -2706
rect 1619 -2707 1634 -2706
rect 1647 -2707 1707 -2706
rect 1759 -2707 1767 -2706
rect 1899 -2707 1907 -2706
rect 2151 -2707 2166 -2706
rect 121 -2709 668 -2708
rect 730 -2709 1039 -2708
rect 1066 -2709 1130 -2708
rect 1206 -2709 1228 -2708
rect 1241 -2709 1893 -2708
rect 1899 -2709 1914 -2708
rect 2165 -2709 2180 -2708
rect 128 -2711 437 -2710
rect 457 -2711 563 -2710
rect 576 -2711 710 -2710
rect 730 -2711 2180 -2710
rect 93 -2713 437 -2712
rect 513 -2713 738 -2712
rect 772 -2713 1172 -2712
rect 1213 -2713 1270 -2712
rect 1276 -2713 1361 -2712
rect 1374 -2713 1508 -2712
rect 1598 -2713 1634 -2712
rect 1647 -2713 1655 -2712
rect 1668 -2713 1697 -2712
rect 1766 -2713 2054 -2712
rect 93 -2715 115 -2714
rect 163 -2715 353 -2714
rect 366 -2715 661 -2714
rect 663 -2715 1277 -2714
rect 1388 -2715 1424 -2714
rect 1430 -2715 1984 -2714
rect 2053 -2715 2082 -2714
rect 114 -2717 479 -2716
rect 513 -2717 1032 -2716
rect 1073 -2717 1284 -2716
rect 1395 -2717 2222 -2716
rect 184 -2719 1392 -2718
rect 1398 -2719 2012 -2718
rect 2060 -2719 2082 -2718
rect 2221 -2719 2264 -2718
rect 75 -2721 185 -2720
rect 226 -2721 388 -2720
rect 478 -2721 857 -2720
rect 877 -2721 1130 -2720
rect 1227 -2721 1315 -2720
rect 1433 -2721 2229 -2720
rect 44 -2723 857 -2722
rect 877 -2723 1088 -2722
rect 1097 -2723 2033 -2722
rect 2060 -2723 2089 -2722
rect 2214 -2723 2229 -2722
rect 44 -2725 472 -2724
rect 576 -2725 647 -2724
rect 667 -2725 703 -2724
rect 779 -2725 850 -2724
rect 912 -2725 1172 -2724
rect 1262 -2725 1291 -2724
rect 1437 -2725 1865 -2724
rect 1962 -2725 1984 -2724
rect 2088 -2725 2096 -2724
rect 135 -2727 913 -2726
rect 933 -2727 1004 -2726
rect 1010 -2727 1242 -2726
rect 1244 -2727 1865 -2726
rect 2095 -2727 2110 -2726
rect 142 -2729 647 -2728
rect 688 -2729 1893 -2728
rect 142 -2731 171 -2730
rect 226 -2731 332 -2730
rect 352 -2731 542 -2730
rect 604 -2731 1193 -2730
rect 1269 -2731 1298 -2730
rect 1437 -2731 1487 -2730
rect 1500 -2731 1508 -2730
rect 1528 -2731 1599 -2730
rect 1626 -2731 1655 -2730
rect 1668 -2731 1683 -2730
rect 1780 -2731 2033 -2730
rect 79 -2733 605 -2732
rect 625 -2733 759 -2732
rect 786 -2733 2173 -2732
rect 9 -2735 80 -2734
rect 149 -2735 332 -2734
rect 415 -2735 1011 -2734
rect 1073 -2735 1158 -2734
rect 1192 -2735 1354 -2734
rect 1440 -2735 2215 -2734
rect 9 -2737 864 -2736
rect 870 -2737 1158 -2736
rect 1290 -2737 1333 -2736
rect 1353 -2737 1368 -2736
rect 1472 -2737 2264 -2736
rect 30 -2739 416 -2738
rect 471 -2739 493 -2738
rect 527 -2739 864 -2738
rect 870 -2739 1046 -2738
rect 1087 -2739 1102 -2738
rect 1108 -2739 1151 -2738
rect 1332 -2739 2208 -2738
rect 30 -2741 255 -2740
rect 261 -2741 360 -2740
rect 408 -2741 1109 -2740
rect 1115 -2741 1312 -2740
rect 1314 -2741 2208 -2740
rect 54 -2743 1046 -2742
rect 1101 -2743 1326 -2742
rect 1367 -2743 1403 -2742
rect 1451 -2743 1473 -2742
rect 1521 -2743 1529 -2742
rect 1580 -2743 1963 -2742
rect 37 -2745 1403 -2744
rect 1521 -2745 1550 -2744
rect 1626 -2745 1641 -2744
rect 1850 -2745 2110 -2744
rect 37 -2747 451 -2746
rect 492 -2747 727 -2746
rect 793 -2747 843 -2746
rect 849 -2747 1256 -2746
rect 1549 -2747 1571 -2746
rect 1689 -2747 1851 -2746
rect 54 -2749 1914 -2748
rect 131 -2751 150 -2750
rect 156 -2751 1434 -2750
rect 1570 -2751 1662 -2750
rect 1689 -2751 1718 -2750
rect 170 -2753 318 -2752
rect 408 -2753 423 -2752
rect 450 -2753 598 -2752
rect 625 -2753 965 -2752
rect 968 -2753 1375 -2752
rect 1542 -2753 1718 -2752
rect 205 -2755 255 -2754
rect 282 -2755 311 -2754
rect 317 -2755 444 -2754
rect 527 -2755 752 -2754
rect 793 -2755 1511 -2754
rect 1542 -2755 1564 -2754
rect 1661 -2755 1676 -2754
rect 205 -2757 1753 -2756
rect 233 -2759 262 -2758
rect 289 -2759 367 -2758
rect 411 -2759 1326 -2758
rect 1675 -2759 1732 -2758
rect 240 -2761 1179 -2760
rect 1255 -2761 1515 -2760
rect 1731 -2761 1858 -2760
rect 243 -2763 402 -2762
rect 443 -2763 706 -2762
rect 744 -2763 969 -2762
rect 982 -2763 1018 -2762
rect 1059 -2763 1179 -2762
rect 1514 -2763 1725 -2762
rect 1857 -2763 1879 -2762
rect 212 -2765 402 -2764
rect 464 -2765 1060 -2764
rect 1115 -2765 1165 -2764
rect 1724 -2765 1739 -2764
rect 1878 -2765 2124 -2764
rect 212 -2767 304 -2766
rect 310 -2767 591 -2766
rect 597 -2767 1466 -2766
rect 1738 -2767 1746 -2766
rect 177 -2769 591 -2768
rect 621 -2769 752 -2768
rect 789 -2769 2124 -2768
rect 177 -2771 899 -2770
rect 943 -2771 1788 -2770
rect 247 -2773 304 -2772
rect 324 -2773 423 -2772
rect 541 -2773 1319 -2772
rect 1465 -2773 1494 -2772
rect 1496 -2773 1746 -2772
rect 289 -2775 570 -2774
rect 639 -2775 717 -2774
rect 744 -2775 1578 -2774
rect 296 -2777 325 -2776
rect 569 -2777 675 -2776
rect 688 -2777 941 -2776
rect 947 -2777 1032 -2776
rect 1122 -2777 1298 -2776
rect 1493 -2777 1711 -2776
rect 72 -2779 297 -2778
rect 460 -2779 1123 -2778
rect 1125 -2779 1844 -2778
rect 72 -2781 237 -2780
rect 268 -2781 675 -2780
rect 702 -2781 1501 -2780
rect 1710 -2781 1802 -2780
rect 198 -2783 948 -2782
rect 961 -2783 2040 -2782
rect 198 -2785 1452 -2784
rect 1794 -2785 1802 -2784
rect 2039 -2785 2075 -2784
rect 219 -2787 269 -2786
rect 611 -2787 640 -2786
rect 789 -2787 1641 -2786
rect 1794 -2787 1809 -2786
rect 2074 -2787 2117 -2786
rect 100 -2789 612 -2788
rect 800 -2789 1329 -2788
rect 1703 -2789 1809 -2788
rect 100 -2791 248 -2790
rect 380 -2791 801 -2790
rect 807 -2791 2047 -2790
rect 219 -2793 899 -2792
rect 940 -2793 1844 -2792
rect 380 -2795 619 -2794
rect 807 -2795 829 -2794
rect 835 -2795 923 -2794
rect 1003 -2795 1025 -2794
rect 1164 -2795 1200 -2794
rect 810 -2797 2194 -2796
rect 814 -2799 1382 -2798
rect 2186 -2799 2194 -2798
rect 544 -2801 2187 -2800
rect 814 -2803 885 -2802
rect 1017 -2803 1081 -2802
rect 1199 -2803 1340 -2802
rect 1381 -2803 1613 -2802
rect 394 -2805 885 -2804
rect 1024 -2805 1756 -2804
rect 394 -2807 458 -2806
rect 821 -2807 906 -2806
rect 1080 -2807 1249 -2806
rect 1339 -2807 1347 -2806
rect 1409 -2807 1613 -2806
rect 618 -2809 1249 -2808
rect 1346 -2809 1970 -2808
rect 824 -2811 1781 -2810
rect 1969 -2811 1991 -2810
rect 828 -2813 1053 -2812
rect 1409 -2813 1417 -2812
rect 1815 -2813 1991 -2812
rect 835 -2815 927 -2814
rect 1052 -2815 1837 -2814
rect 191 -2817 927 -2816
rect 1815 -2817 1823 -2816
rect 1836 -2817 1921 -2816
rect 191 -2819 535 -2818
rect 866 -2819 2117 -2818
rect 275 -2821 535 -2820
rect 894 -2821 1417 -2820
rect 1535 -2821 1921 -2820
rect 275 -2823 500 -2822
rect 905 -2823 1305 -2822
rect 1822 -2823 1830 -2822
rect 485 -2825 500 -2824
rect 989 -2825 1536 -2824
rect 1829 -2825 1998 -2824
rect 429 -2827 486 -2826
rect 989 -2827 1095 -2826
rect 1304 -2827 1312 -2826
rect 1997 -2827 2026 -2826
rect 240 -2829 1095 -2828
rect 2025 -2829 2068 -2828
rect 1941 -2831 2068 -2830
rect 222 -2833 1942 -2832
rect 23 -2844 468 -2843
rect 541 -2844 1497 -2843
rect 1500 -2844 2257 -2843
rect 23 -2846 185 -2845
rect 219 -2846 381 -2845
rect 429 -2846 493 -2845
rect 548 -2846 787 -2845
rect 814 -2846 941 -2845
rect 943 -2846 1333 -2845
rect 1346 -2846 1634 -2845
rect 1682 -2846 2138 -2845
rect 2221 -2846 2250 -2845
rect 30 -2848 545 -2847
rect 548 -2848 892 -2847
rect 919 -2848 1140 -2847
rect 1202 -2848 1210 -2847
rect 1255 -2848 1326 -2847
rect 1332 -2848 1620 -2847
rect 1682 -2848 2061 -2847
rect 2074 -2848 2138 -2847
rect 30 -2850 258 -2849
rect 317 -2850 790 -2849
rect 828 -2850 892 -2849
rect 922 -2850 1501 -2849
rect 1566 -2850 2005 -2849
rect 2060 -2850 2208 -2849
rect 51 -2852 479 -2851
rect 492 -2852 528 -2851
rect 544 -2852 913 -2851
rect 964 -2852 1235 -2851
rect 1258 -2852 1921 -2851
rect 2004 -2852 2103 -2851
rect 82 -2854 409 -2853
rect 457 -2854 500 -2853
rect 527 -2854 738 -2853
rect 744 -2854 843 -2853
rect 863 -2854 1984 -2853
rect 2074 -2854 2215 -2853
rect 103 -2856 353 -2855
rect 373 -2856 409 -2855
rect 460 -2856 556 -2855
rect 565 -2856 941 -2855
rect 968 -2856 972 -2855
rect 975 -2856 1375 -2855
rect 1391 -2856 1851 -2855
rect 1983 -2856 2089 -2855
rect 2098 -2856 2103 -2855
rect 107 -2858 388 -2857
rect 401 -2858 815 -2857
rect 835 -2858 927 -2857
rect 968 -2858 983 -2857
rect 1017 -2858 1060 -2857
rect 1062 -2858 1088 -2857
rect 1136 -2858 1620 -2857
rect 1703 -2858 2033 -2857
rect 2088 -2858 2236 -2857
rect 117 -2860 1893 -2859
rect 2032 -2860 2152 -2859
rect 124 -2862 857 -2861
rect 866 -2862 1098 -2861
rect 1234 -2862 1291 -2861
rect 1314 -2862 1557 -2861
rect 1703 -2862 1774 -2861
rect 1850 -2862 1998 -2861
rect 191 -2864 402 -2863
rect 485 -2864 556 -2863
rect 597 -2864 661 -2863
rect 674 -2864 927 -2863
rect 971 -2864 983 -2863
rect 1017 -2864 1137 -2863
rect 1283 -2864 1382 -2863
rect 1433 -2864 1718 -2863
rect 1731 -2864 1921 -2863
rect 128 -2866 598 -2865
rect 611 -2866 1126 -2865
rect 1286 -2866 1697 -2865
rect 1706 -2866 2019 -2865
rect 86 -2868 129 -2867
rect 191 -2868 213 -2867
rect 219 -2868 444 -2867
rect 485 -2868 521 -2867
rect 583 -2868 612 -2867
rect 621 -2868 801 -2867
rect 856 -2868 1242 -2867
rect 1290 -2868 1340 -2867
rect 1346 -2868 1473 -2867
rect 1486 -2868 2110 -2867
rect 86 -2870 248 -2869
rect 250 -2870 1403 -2869
rect 1419 -2870 1473 -2869
rect 1489 -2870 1634 -2869
rect 1696 -2870 1816 -2869
rect 1878 -2870 1998 -2869
rect 2018 -2870 2124 -2869
rect 72 -2872 248 -2871
rect 289 -2872 318 -2871
rect 324 -2872 430 -2871
rect 443 -2872 472 -2871
rect 499 -2872 605 -2871
rect 674 -2872 1312 -2871
rect 1314 -2872 2201 -2871
rect 58 -2874 73 -2873
rect 135 -2874 605 -2873
rect 681 -2874 913 -2873
rect 1038 -2874 1350 -2873
rect 1360 -2874 1364 -2873
rect 1374 -2874 1424 -2873
rect 1451 -2874 2194 -2873
rect 58 -2876 1249 -2875
rect 1339 -2876 1368 -2875
rect 1381 -2876 1438 -2875
rect 1493 -2876 1686 -2875
rect 1717 -2876 1858 -2875
rect 1892 -2876 1977 -2875
rect 2109 -2876 2243 -2875
rect 100 -2878 1368 -2877
rect 1402 -2878 1410 -2877
rect 1437 -2878 2271 -2877
rect 100 -2880 1732 -2879
rect 1752 -2880 1907 -2879
rect 1976 -2880 2180 -2879
rect 110 -2882 1410 -2881
rect 1493 -2882 1543 -2881
rect 1556 -2882 1641 -2881
rect 1752 -2882 1872 -2881
rect 1906 -2882 2012 -2881
rect 2123 -2882 2225 -2881
rect 135 -2884 577 -2883
rect 583 -2884 850 -2883
rect 880 -2884 1102 -2883
rect 1115 -2884 1424 -2883
rect 1444 -2884 1543 -2883
rect 1640 -2884 1760 -2883
rect 1773 -2884 1886 -2883
rect 2011 -2884 2117 -2883
rect 65 -2886 850 -2885
rect 961 -2886 2117 -2885
rect 205 -2888 479 -2887
rect 520 -2888 1053 -2887
rect 1059 -2888 1459 -2887
rect 1755 -2888 1991 -2887
rect 2 -2890 206 -2889
rect 212 -2890 633 -2889
rect 642 -2890 1452 -2889
rect 1759 -2890 1830 -2889
rect 1871 -2890 2260 -2889
rect 222 -2892 2047 -2891
rect 233 -2894 304 -2893
rect 310 -2894 353 -2893
rect 373 -2894 416 -2893
rect 576 -2894 1417 -2893
rect 1444 -2894 1480 -2893
rect 1801 -2894 1879 -2893
rect 1990 -2894 2096 -2893
rect 233 -2896 269 -2895
rect 289 -2896 535 -2895
rect 590 -2896 682 -2895
rect 688 -2896 829 -2895
rect 961 -2896 2152 -2895
rect 163 -2898 269 -2897
rect 275 -2898 535 -2897
rect 590 -2898 808 -2897
rect 978 -2898 1886 -2897
rect 2046 -2898 2166 -2897
rect 163 -2900 934 -2899
rect 1010 -2900 1459 -2899
rect 1479 -2900 1599 -2899
rect 1801 -2900 1942 -2899
rect 236 -2902 304 -2901
rect 310 -2902 423 -2901
rect 632 -2902 724 -2901
rect 730 -2902 1389 -2901
rect 1598 -2902 1613 -2901
rect 1815 -2902 1837 -2901
rect 1941 -2902 2040 -2901
rect 16 -2904 731 -2903
rect 744 -2904 1074 -2903
rect 1087 -2904 1123 -2903
rect 1199 -2904 1858 -2903
rect 2039 -2904 2159 -2903
rect 37 -2906 724 -2905
rect 747 -2906 948 -2905
rect 954 -2906 1123 -2905
rect 1241 -2906 1298 -2905
rect 1360 -2906 1522 -2905
rect 1612 -2906 1676 -2905
rect 1829 -2906 1949 -2905
rect 37 -2908 143 -2907
rect 275 -2908 367 -2907
rect 380 -2908 734 -2907
rect 737 -2908 1676 -2907
rect 1836 -2908 1914 -2907
rect 142 -2910 766 -2909
rect 772 -2910 864 -2909
rect 933 -2910 1095 -2909
rect 1101 -2910 1144 -2909
rect 1248 -2910 1277 -2909
rect 1297 -2910 1396 -2909
rect 1521 -2910 1627 -2909
rect 1913 -2910 2026 -2909
rect 324 -2912 395 -2911
rect 415 -2912 1056 -2911
rect 1066 -2912 1326 -2911
rect 1388 -2912 1466 -2911
rect 2025 -2912 2131 -2911
rect 44 -2914 1067 -2913
rect 1069 -2914 1655 -2913
rect 2130 -2914 2264 -2913
rect 44 -2916 619 -2915
rect 646 -2916 808 -2915
rect 842 -2916 1200 -2915
rect 1276 -2916 1354 -2915
rect 1395 -2916 1508 -2915
rect 1654 -2916 1690 -2915
rect 9 -2918 619 -2917
rect 660 -2918 1627 -2917
rect 1689 -2918 1746 -2917
rect 198 -2920 395 -2919
rect 422 -2920 465 -2919
rect 562 -2920 647 -2919
rect 663 -2920 948 -2919
rect 954 -2920 1039 -2919
rect 1045 -2920 1487 -2919
rect 1507 -2920 1592 -2919
rect 1745 -2920 1865 -2919
rect 65 -2922 465 -2921
rect 506 -2922 563 -2921
rect 663 -2922 1179 -2921
rect 1465 -2922 1578 -2921
rect 1710 -2922 1865 -2921
rect 121 -2924 507 -2923
rect 688 -2924 1172 -2923
rect 1178 -2924 1305 -2923
rect 1430 -2924 1578 -2923
rect 1710 -2924 1795 -2923
rect 121 -2926 185 -2925
rect 331 -2926 472 -2925
rect 702 -2926 1158 -2925
rect 1171 -2926 1214 -2925
rect 1304 -2926 1844 -2925
rect 149 -2928 199 -2927
rect 240 -2928 332 -2927
rect 345 -2928 367 -2927
rect 387 -2928 1056 -2927
rect 1073 -2928 1130 -2927
rect 1213 -2928 1263 -2927
rect 1430 -2928 1529 -2927
rect 1570 -2928 1592 -2927
rect 1794 -2928 1956 -2927
rect 149 -2930 1025 -2929
rect 1031 -2930 1046 -2929
rect 1080 -2930 1354 -2929
rect 1528 -2930 1585 -2929
rect 1843 -2930 1963 -2929
rect 156 -2932 241 -2931
rect 345 -2932 794 -2931
rect 989 -2932 1025 -2931
rect 1080 -2932 1662 -2931
rect 1955 -2932 2068 -2931
rect 513 -2934 1130 -2933
rect 1192 -2934 1263 -2933
rect 1514 -2934 1585 -2933
rect 1661 -2934 1739 -2933
rect 1962 -2934 2082 -2933
rect 296 -2936 514 -2935
rect 569 -2936 703 -2935
rect 705 -2936 885 -2935
rect 989 -2936 1032 -2935
rect 1094 -2936 1144 -2935
rect 1192 -2936 1270 -2935
rect 1514 -2936 1606 -2935
rect 1738 -2936 2096 -2935
rect 54 -2938 1270 -2937
rect 1605 -2938 1669 -2937
rect 2067 -2938 2187 -2937
rect 170 -2940 570 -2939
rect 709 -2940 885 -2939
rect 1010 -2940 1207 -2939
rect 1668 -2940 1788 -2939
rect 2081 -2940 2229 -2939
rect 170 -2942 262 -2941
rect 296 -2942 339 -2941
rect 695 -2942 710 -2941
rect 740 -2942 1949 -2941
rect 254 -2944 339 -2943
rect 667 -2944 696 -2943
rect 751 -2944 1564 -2943
rect 1787 -2944 1935 -2943
rect 16 -2946 255 -2945
rect 261 -2946 360 -2945
rect 667 -2946 1571 -2945
rect 177 -2948 752 -2947
rect 765 -2948 1151 -2947
rect 1157 -2948 1935 -2947
rect 177 -2950 216 -2949
rect 226 -2950 360 -2949
rect 772 -2950 1004 -2949
rect 1115 -2950 1165 -2949
rect 1206 -2950 1536 -2949
rect 1563 -2950 1648 -2949
rect 159 -2952 227 -2951
rect 779 -2952 801 -2951
rect 870 -2952 1004 -2951
rect 1150 -2952 1186 -2951
rect 1535 -2952 1725 -2951
rect 779 -2954 878 -2953
rect 905 -2954 1165 -2953
rect 1185 -2954 1221 -2953
rect 1647 -2954 1781 -2953
rect 93 -2956 906 -2955
rect 1097 -2956 1221 -2955
rect 1724 -2956 1823 -2955
rect 79 -2958 94 -2957
rect 793 -2958 822 -2957
rect 870 -2958 899 -2957
rect 1780 -2958 1928 -2957
rect 79 -2960 997 -2959
rect 1822 -2960 1970 -2959
rect 114 -2962 899 -2961
rect 996 -2962 1109 -2961
rect 1927 -2962 2054 -2961
rect 114 -2964 451 -2963
rect 758 -2964 822 -2963
rect 1108 -2964 1228 -2963
rect 1808 -2964 2054 -2963
rect 450 -2966 1042 -2965
rect 1227 -2966 1319 -2965
rect 1808 -2966 1900 -2965
rect 1969 -2966 2173 -2965
rect 653 -2968 759 -2967
rect 1318 -2968 1550 -2967
rect 1766 -2968 1900 -2967
rect 639 -2970 654 -2969
rect 1160 -2970 1550 -2969
rect 282 -2972 640 -2971
rect 282 -2974 626 -2973
rect 625 -2976 717 -2975
rect 716 -2978 986 -2977
rect 16 -2989 111 -2988
rect 114 -2989 388 -2988
rect 422 -2989 461 -2988
rect 471 -2989 563 -2988
rect 569 -2989 976 -2988
rect 1041 -2989 2061 -2988
rect 2095 -2989 2138 -2988
rect 51 -2991 73 -2990
rect 100 -2991 934 -2990
rect 961 -2991 969 -2990
rect 1052 -2991 1326 -2990
rect 1360 -2991 1410 -2990
rect 1416 -2991 1858 -2990
rect 1871 -2991 1875 -2990
rect 2098 -2991 2117 -2990
rect 37 -2993 73 -2992
rect 93 -2993 101 -2992
rect 107 -2993 780 -2992
rect 880 -2993 1690 -2992
rect 1769 -2993 1816 -2992
rect 1836 -2993 1858 -2992
rect 1871 -2993 1991 -2992
rect 30 -2995 94 -2994
rect 142 -2995 920 -2994
rect 964 -2995 1032 -2994
rect 1055 -2995 1837 -2994
rect 1892 -2995 1991 -2994
rect 30 -2997 59 -2996
rect 65 -2997 566 -2996
rect 572 -2997 962 -2996
rect 968 -2997 1088 -2996
rect 1125 -2997 1494 -2996
rect 1566 -2997 1886 -2996
rect 37 -2999 521 -2998
rect 541 -2999 815 -2998
rect 884 -2999 934 -2998
rect 1031 -2999 1186 -2998
rect 1199 -2999 1977 -2998
rect 44 -3001 66 -3000
rect 135 -3001 542 -3000
rect 590 -3001 916 -3000
rect 954 -3001 1186 -3000
rect 1199 -3001 1249 -3000
rect 1318 -3001 1417 -3000
rect 1419 -3001 1921 -3000
rect 1976 -3001 2103 -3000
rect 58 -3003 199 -3002
rect 208 -3003 444 -3002
rect 471 -3003 881 -3002
rect 894 -3003 1879 -3002
rect 1885 -3003 1984 -3002
rect 142 -3005 206 -3004
rect 212 -3005 339 -3004
rect 422 -3005 430 -3004
rect 443 -3005 1277 -3004
rect 1318 -3005 1340 -3004
rect 1398 -3005 1942 -3004
rect 86 -3007 213 -3006
rect 236 -3007 619 -3006
rect 642 -3007 759 -3006
rect 786 -3007 955 -3006
rect 1055 -3007 1704 -3006
rect 1808 -3007 1882 -3006
rect 1920 -3007 2026 -3006
rect 86 -3009 220 -3008
rect 240 -3009 430 -3008
rect 478 -3009 619 -3008
rect 688 -3009 1039 -3008
rect 1066 -3009 1095 -3008
rect 1139 -3009 1634 -3008
rect 1654 -3009 1942 -3008
rect 131 -3011 787 -3010
rect 905 -3011 920 -3010
rect 1038 -3011 1221 -3010
rect 1325 -3011 1560 -3010
rect 1570 -3011 1865 -3010
rect 149 -3013 465 -3012
rect 478 -3013 668 -3012
rect 688 -3013 1256 -3012
rect 1339 -3013 1431 -3012
rect 1486 -3013 1767 -3012
rect 1808 -3013 2054 -3012
rect 138 -3015 150 -3014
rect 156 -3015 664 -3014
rect 667 -3015 696 -3014
rect 716 -3015 720 -3014
rect 730 -3015 923 -3014
rect 1045 -3015 1067 -3014
rect 1069 -3015 1214 -3014
rect 1220 -3015 1228 -3014
rect 1255 -3015 1270 -3014
rect 1402 -3015 1406 -3014
rect 1430 -3015 1501 -3014
rect 1570 -3015 1606 -3014
rect 1633 -3015 1676 -3014
rect 1689 -3015 1774 -3014
rect 1815 -3015 1949 -3014
rect 156 -3017 192 -3016
rect 198 -3017 262 -3016
rect 282 -3017 570 -3016
rect 590 -3017 703 -3016
rect 716 -3017 801 -3016
rect 849 -3017 906 -3016
rect 1045 -3017 1144 -3016
rect 1160 -3017 1354 -3016
rect 1402 -3017 1529 -3016
rect 1549 -3017 1676 -3016
rect 1703 -3017 1781 -3016
rect 1864 -3017 2040 -3016
rect 128 -3019 1161 -3018
rect 1178 -3019 1207 -3018
rect 1213 -3019 1424 -3018
rect 1486 -3019 1564 -3018
rect 1573 -3019 2131 -3018
rect 159 -3021 1074 -3020
rect 1076 -3021 1438 -3020
rect 1493 -3021 1522 -3020
rect 1528 -3021 1683 -3020
rect 1759 -3021 1781 -3020
rect 1874 -3021 1893 -3020
rect 1948 -3021 2089 -3020
rect 163 -3023 521 -3022
rect 597 -3023 640 -3022
rect 695 -3023 710 -3022
rect 730 -3023 1081 -3022
rect 1083 -3023 1935 -3022
rect 166 -3025 927 -3024
rect 1087 -3025 1116 -3024
rect 1143 -3025 1305 -3024
rect 1353 -3025 1396 -3024
rect 1423 -3025 1480 -3024
rect 1500 -3025 1557 -3024
rect 1654 -3025 1746 -3024
rect 1759 -3025 1851 -3024
rect 1934 -3025 2012 -3024
rect 79 -3027 927 -3026
rect 985 -3027 1851 -3026
rect 170 -3029 262 -3028
rect 282 -3029 381 -3028
rect 457 -3029 598 -3028
rect 614 -3029 899 -3028
rect 1178 -3029 1242 -3028
rect 1269 -3029 1291 -3028
rect 1304 -3029 1473 -3028
rect 1549 -3029 1613 -3028
rect 1661 -3029 1686 -3028
rect 1745 -3029 1956 -3028
rect 173 -3031 605 -3030
rect 625 -3031 1116 -3030
rect 1192 -3031 1606 -3030
rect 1612 -3031 1641 -3030
rect 1661 -3031 1725 -3030
rect 1766 -3031 1844 -3030
rect 184 -3033 192 -3032
rect 219 -3033 374 -3032
rect 457 -3033 976 -3032
rect 1164 -3033 1193 -3032
rect 1202 -3033 1410 -3032
rect 1437 -3033 1515 -3032
rect 1598 -3033 1641 -3032
rect 1682 -3033 1984 -3032
rect 184 -3035 206 -3034
rect 215 -3035 374 -3034
rect 485 -3035 738 -3034
rect 740 -3035 871 -3034
rect 1136 -3035 1599 -3034
rect 1724 -3035 2075 -3034
rect 240 -3037 269 -3036
rect 296 -3037 661 -3036
rect 702 -3037 724 -3036
rect 737 -3037 913 -3036
rect 1136 -3037 1235 -3036
rect 1241 -3037 1389 -3036
rect 1451 -3037 1522 -3036
rect 1773 -3037 1823 -3036
rect 1843 -3037 2005 -3036
rect 2074 -3037 2152 -3036
rect 254 -3039 1368 -3038
rect 1388 -3039 1718 -3038
rect 1822 -3039 2019 -3038
rect 247 -3041 255 -3040
rect 268 -3041 1060 -3040
rect 1157 -3041 1368 -3040
rect 1451 -3041 1732 -3040
rect 2004 -3041 2082 -3040
rect 103 -3043 248 -3042
rect 296 -3043 402 -3042
rect 415 -3043 724 -3042
rect 758 -3043 818 -3042
rect 870 -3043 948 -3042
rect 1017 -3043 1732 -3042
rect 275 -3045 402 -3044
rect 415 -3045 507 -3044
rect 513 -3045 780 -3044
rect 835 -3045 948 -3044
rect 1003 -3045 1018 -3044
rect 1059 -3045 1102 -3044
rect 1164 -3045 1238 -3044
rect 1283 -3045 1291 -3044
rect 1332 -3045 1480 -3044
rect 1514 -3045 1543 -3044
rect 1717 -3045 1795 -3044
rect 275 -3047 325 -3046
rect 338 -3047 367 -3046
rect 485 -3047 556 -3046
rect 625 -3047 675 -3046
rect 709 -3047 1063 -3046
rect 1097 -3047 1333 -3046
rect 1465 -3047 1956 -3046
rect 289 -3049 556 -3048
rect 660 -3049 682 -3048
rect 765 -3049 850 -3048
rect 884 -3049 1235 -3048
rect 1283 -3049 1298 -3048
rect 1465 -3049 1739 -3048
rect 1794 -3049 1928 -3048
rect 289 -3051 633 -3050
rect 674 -3051 1130 -3050
rect 1227 -3051 1263 -3050
rect 1297 -3051 1312 -3050
rect 1472 -3051 1966 -3050
rect 310 -3053 388 -3052
rect 506 -3053 997 -3052
rect 1024 -3053 1263 -3052
rect 1311 -3053 1536 -3052
rect 1542 -3053 1585 -3052
rect 1738 -3053 1802 -3052
rect 1927 -3053 2068 -3052
rect 310 -3055 1074 -3054
rect 1101 -3055 1151 -3054
rect 1535 -3055 1592 -3054
rect 1801 -3055 1907 -3054
rect 324 -3057 500 -3056
rect 513 -3057 535 -3056
rect 548 -3057 1158 -3056
rect 1584 -3057 1620 -3056
rect 1906 -3057 2033 -3056
rect 226 -3059 535 -3058
rect 632 -3059 829 -3058
rect 835 -3059 1382 -3058
rect 1591 -3059 1627 -3058
rect 2032 -3059 2110 -3058
rect 121 -3061 227 -3060
rect 352 -3061 549 -3060
rect 681 -3061 843 -3060
rect 940 -3061 1004 -3060
rect 1024 -3061 1109 -3060
rect 1122 -3061 1151 -3060
rect 1381 -3061 1445 -3060
rect 1619 -3061 1648 -3060
rect 121 -3063 577 -3062
rect 765 -3063 857 -3062
rect 940 -3063 1375 -3062
rect 1626 -3063 1697 -3062
rect 124 -3065 353 -3064
rect 359 -3065 381 -3064
rect 450 -3065 829 -3064
rect 856 -3065 864 -3064
rect 996 -3065 1217 -3064
rect 1556 -3065 1697 -3064
rect 359 -3067 545 -3066
rect 576 -3067 654 -3066
rect 772 -3067 899 -3066
rect 1010 -3067 1109 -3066
rect 1129 -3067 1172 -3066
rect 1647 -3067 1711 -3066
rect 366 -3069 395 -3068
rect 450 -3069 493 -3068
rect 499 -3069 1364 -3068
rect 1710 -3069 1788 -3068
rect 317 -3071 395 -3070
rect 492 -3071 647 -3070
rect 653 -3071 892 -3070
rect 1034 -3071 1375 -3070
rect 1787 -3071 1900 -3070
rect 177 -3073 318 -3072
rect 527 -3073 605 -3072
rect 611 -3073 647 -3072
rect 744 -3073 1011 -3072
rect 1171 -3073 1315 -3072
rect 1899 -3073 1998 -3072
rect 23 -3075 612 -3074
rect 772 -3075 822 -3074
rect 863 -3075 1970 -3074
rect 23 -3077 983 -3076
rect 1507 -3077 1970 -3076
rect 177 -3079 304 -3078
rect 331 -3079 822 -3078
rect 982 -3079 990 -3078
rect 1507 -3079 1578 -3078
rect 1913 -3079 1998 -3078
rect 233 -3081 304 -3080
rect 331 -3081 346 -3080
rect 583 -3081 745 -3080
rect 807 -3081 843 -3080
rect 877 -3081 1578 -3080
rect 1913 -3081 2047 -3080
rect 345 -3083 409 -3082
rect 583 -3083 752 -3082
rect 793 -3083 808 -3082
rect 989 -3083 1459 -3082
rect 2046 -3083 2124 -3082
rect 117 -3085 409 -3084
rect 751 -3085 913 -3084
rect 1458 -3085 1669 -3084
rect 793 -3087 1210 -3086
rect 1668 -3087 1753 -3086
rect 1752 -3089 1830 -3088
rect 1829 -3091 1963 -3090
rect 1962 -3093 2145 -3092
rect 23 -3104 209 -3103
rect 212 -3104 234 -3103
rect 380 -3104 458 -3103
rect 520 -3104 818 -3103
rect 821 -3104 1312 -3103
rect 1381 -3104 1403 -3103
rect 1461 -3104 1865 -3103
rect 1962 -3104 2047 -3103
rect 30 -3106 206 -3105
rect 212 -3106 1168 -3105
rect 1199 -3106 1259 -3105
rect 1276 -3106 1452 -3105
rect 1465 -3106 1564 -3105
rect 1566 -3106 1683 -3105
rect 1853 -3106 1893 -3105
rect 1997 -3106 2019 -3105
rect 2046 -3106 2075 -3105
rect 58 -3108 132 -3107
rect 187 -3108 689 -3107
rect 737 -3108 1445 -3107
rect 1451 -3108 1536 -3107
rect 1640 -3108 1879 -3107
rect 1892 -3108 1949 -3107
rect 65 -3110 1112 -3109
rect 1199 -3110 1305 -3109
rect 1311 -3110 1704 -3109
rect 1864 -3110 1872 -3109
rect 1878 -3110 1900 -3109
rect 72 -3112 237 -3111
rect 289 -3112 822 -3111
rect 835 -3112 1123 -3111
rect 1216 -3112 1606 -3111
rect 1671 -3112 1858 -3111
rect 79 -3114 675 -3113
rect 681 -3114 1161 -3113
rect 1234 -3114 1347 -3113
rect 1381 -3114 1634 -3113
rect 1675 -3114 1963 -3113
rect 86 -3116 139 -3115
rect 194 -3116 283 -3115
rect 289 -3116 426 -3115
rect 506 -3116 738 -3115
rect 758 -3116 1644 -3115
rect 1857 -3116 1886 -3115
rect 93 -3118 143 -3117
rect 254 -3118 283 -3117
rect 352 -3118 1347 -3117
rect 1395 -3118 1473 -3117
rect 1486 -3118 1557 -3117
rect 1605 -3118 1851 -3117
rect 1885 -3118 1921 -3117
rect 107 -3120 881 -3119
rect 891 -3120 1116 -3119
rect 1122 -3120 1326 -3119
rect 1395 -3120 1711 -3119
rect 1920 -3120 1977 -3119
rect 107 -3122 178 -3121
rect 226 -3122 353 -3121
rect 380 -3122 580 -3121
rect 604 -3122 878 -3121
rect 898 -3122 1116 -3121
rect 1237 -3122 1410 -3121
rect 1437 -3122 1564 -3121
rect 1633 -3122 1788 -3121
rect 1976 -3122 2005 -3121
rect 114 -3124 167 -3123
rect 177 -3124 808 -3123
rect 828 -3124 892 -3123
rect 943 -3124 1725 -3123
rect 100 -3126 115 -3125
rect 121 -3126 209 -3125
rect 254 -3126 360 -3125
rect 401 -3126 531 -3125
rect 555 -3126 874 -3125
rect 877 -3126 1448 -3125
rect 1465 -3126 1613 -3125
rect 1647 -3126 1725 -3125
rect 100 -3128 311 -3127
rect 359 -3128 367 -3127
rect 373 -3128 556 -3127
rect 569 -3128 818 -3127
rect 828 -3128 1207 -3127
rect 1248 -3128 1270 -3127
rect 1276 -3128 1882 -3127
rect 121 -3130 157 -3129
rect 191 -3130 227 -3129
rect 275 -3130 402 -3129
rect 404 -3130 458 -3129
rect 471 -3130 605 -3129
rect 625 -3130 1084 -3129
rect 1094 -3130 1126 -3129
rect 1185 -3130 1270 -3129
rect 1297 -3130 1315 -3129
rect 1318 -3130 1641 -3129
rect 1647 -3130 1956 -3129
rect 135 -3132 276 -3131
rect 296 -3132 374 -3131
rect 471 -3132 535 -3131
rect 541 -3132 570 -3131
rect 625 -3132 710 -3131
rect 716 -3132 836 -3131
rect 863 -3132 920 -3131
rect 961 -3132 1704 -3131
rect 135 -3134 269 -3133
rect 310 -3134 318 -3133
rect 366 -3134 430 -3133
rect 443 -3134 710 -3133
rect 758 -3134 955 -3133
rect 961 -3134 1032 -3133
rect 1045 -3134 1711 -3133
rect 142 -3136 913 -3135
rect 968 -3136 1560 -3135
rect 1612 -3136 1823 -3135
rect 156 -3138 192 -3137
rect 219 -3138 297 -3137
rect 317 -3138 332 -3137
rect 429 -3138 598 -3137
rect 632 -3138 808 -3137
rect 856 -3138 920 -3137
rect 968 -3138 1228 -3137
rect 1248 -3138 1368 -3137
rect 1402 -3138 1550 -3137
rect 1556 -3138 1907 -3137
rect 173 -3140 1046 -3139
rect 1073 -3140 1305 -3139
rect 1318 -3140 1718 -3139
rect 1766 -3140 1823 -3139
rect 1906 -3140 1935 -3139
rect 205 -3142 633 -3141
rect 639 -3142 867 -3141
rect 912 -3142 1375 -3141
rect 1409 -3142 1543 -3141
rect 1549 -3142 1627 -3141
rect 1661 -3142 1767 -3141
rect 219 -3144 262 -3143
rect 268 -3144 346 -3143
rect 394 -3144 640 -3143
rect 681 -3144 703 -3143
rect 765 -3144 1032 -3143
rect 1073 -3144 1172 -3143
rect 1185 -3144 1361 -3143
rect 1367 -3144 1578 -3143
rect 1626 -3144 1928 -3143
rect 261 -3146 1158 -3145
rect 1171 -3146 1459 -3145
rect 1472 -3146 1669 -3145
rect 1675 -3146 1851 -3145
rect 331 -3148 584 -3147
rect 597 -3148 619 -3147
rect 688 -3148 794 -3147
rect 800 -3148 857 -3147
rect 1017 -3148 1053 -3147
rect 1076 -3148 1658 -3147
rect 1661 -3148 1844 -3147
rect 338 -3150 346 -3149
rect 394 -3150 661 -3149
rect 702 -3150 1025 -3149
rect 1094 -3150 1221 -3149
rect 1227 -3150 1333 -3149
rect 1360 -3150 1508 -3149
rect 1535 -3150 1592 -3149
rect 338 -3152 451 -3151
rect 485 -3152 542 -3151
rect 576 -3152 717 -3151
rect 768 -3152 1193 -3151
rect 1206 -3152 1217 -3151
rect 1220 -3152 1242 -3151
rect 1262 -3152 1445 -3151
rect 1486 -3152 1655 -3151
rect 37 -3154 577 -3153
rect 583 -3154 1056 -3153
rect 1101 -3154 1214 -3153
rect 1241 -3154 1417 -3153
rect 1437 -3154 1686 -3153
rect 418 -3156 451 -3155
rect 485 -3156 724 -3155
rect 793 -3156 843 -3155
rect 985 -3156 1508 -3155
rect 1542 -3156 1816 -3155
rect 443 -3158 1214 -3157
rect 1262 -3158 1494 -3157
rect 1570 -3158 1718 -3157
rect 1738 -3158 1816 -3157
rect 506 -3160 934 -3159
rect 989 -3160 1193 -3159
rect 1297 -3160 1966 -3159
rect 520 -3162 1399 -3161
rect 1416 -3162 1585 -3161
rect 1591 -3162 1802 -3161
rect 1965 -3162 2033 -3161
rect 527 -3164 885 -3163
rect 905 -3164 990 -3163
rect 1003 -3164 1018 -3163
rect 1024 -3164 1060 -3163
rect 1101 -3164 1137 -3163
rect 1157 -3164 1291 -3163
rect 1325 -3164 1515 -3163
rect 1521 -3164 1739 -3163
rect 324 -3166 1291 -3165
rect 1332 -3166 1480 -3165
rect 1493 -3166 1690 -3165
rect 324 -3168 388 -3167
rect 527 -3168 745 -3167
rect 786 -3168 885 -3167
rect 905 -3168 976 -3167
rect 1003 -3168 1067 -3167
rect 1143 -3168 1480 -3167
rect 1500 -3168 1571 -3167
rect 1577 -3168 1942 -3167
rect 387 -3170 514 -3169
rect 534 -3170 773 -3169
rect 800 -3170 1690 -3169
rect 464 -3172 745 -3171
rect 814 -3172 1375 -3171
rect 1500 -3172 1599 -3171
rect 1650 -3172 1686 -3171
rect 163 -3174 465 -3173
rect 492 -3174 976 -3173
rect 1059 -3174 1151 -3173
rect 1356 -3174 1522 -3173
rect 1584 -3174 1732 -3173
rect 163 -3176 766 -3175
rect 933 -3176 983 -3175
rect 1066 -3176 1109 -3175
rect 1143 -3176 1179 -3175
rect 1514 -3176 1697 -3175
rect 1731 -3176 1746 -3175
rect 415 -3178 493 -3177
rect 513 -3178 591 -3177
rect 611 -3178 787 -3177
rect 940 -3178 1137 -3177
rect 1150 -3178 1284 -3177
rect 1598 -3178 1837 -3177
rect 415 -3180 899 -3179
rect 954 -3180 1179 -3179
rect 1283 -3180 1340 -3179
rect 1654 -3180 1970 -3179
rect 184 -3182 1340 -3181
rect 1696 -3182 1809 -3181
rect 1969 -3182 1984 -3181
rect 590 -3184 696 -3183
rect 730 -3184 815 -3183
rect 1108 -3184 1354 -3183
rect 1745 -3184 1760 -3183
rect 1780 -3184 1809 -3183
rect 1983 -3184 1991 -3183
rect 82 -3186 731 -3185
rect 772 -3186 1354 -3185
rect 1752 -3186 1760 -3185
rect 1773 -3186 1781 -3185
rect 562 -3188 696 -3187
rect 1752 -3188 1795 -3187
rect 499 -3190 563 -3189
rect 611 -3190 668 -3189
rect 674 -3190 724 -3189
rect 1773 -3190 1830 -3189
rect 499 -3192 780 -3191
rect 614 -3194 941 -3193
rect 247 -3196 615 -3195
rect 618 -3196 647 -3195
rect 653 -3196 843 -3195
rect 240 -3198 248 -3197
rect 478 -3198 654 -3197
rect 660 -3198 1081 -3197
rect 170 -3200 241 -3199
rect 408 -3200 479 -3199
rect 548 -3200 647 -3199
rect 667 -3200 871 -3199
rect 170 -3202 752 -3201
rect 779 -3202 948 -3201
rect 128 -3204 752 -3203
rect 849 -3204 1081 -3203
rect 128 -3206 150 -3205
rect 408 -3206 423 -3205
rect 548 -3206 748 -3205
rect 849 -3206 1039 -3205
rect 149 -3208 461 -3207
rect 947 -3208 997 -3207
rect 1038 -3208 1088 -3207
rect 996 -3210 1011 -3209
rect 1087 -3210 1256 -3209
rect 1010 -3212 1459 -3211
rect 1255 -3214 1424 -3213
rect 1164 -3216 1424 -3215
rect 1164 -3218 1529 -3217
rect 1430 -3220 1529 -3219
rect 1430 -3222 1620 -3221
rect 1619 -3224 1914 -3223
rect 93 -3235 174 -3234
rect 184 -3235 538 -3234
rect 548 -3235 601 -3234
rect 642 -3235 773 -3234
rect 800 -3235 1445 -3234
rect 1563 -3235 1644 -3234
rect 1668 -3235 1728 -3234
rect 1738 -3235 1966 -3234
rect 2018 -3235 2026 -3234
rect 2032 -3235 2047 -3234
rect 107 -3237 678 -3236
rect 688 -3237 1165 -3236
rect 1213 -3237 1599 -3236
rect 1640 -3237 1746 -3236
rect 1766 -3237 1788 -3236
rect 1808 -3237 1851 -3236
rect 1871 -3237 1886 -3236
rect 1962 -3237 1984 -3236
rect 121 -3239 206 -3238
rect 208 -3239 227 -3238
rect 233 -3239 258 -3238
rect 275 -3239 783 -3238
rect 800 -3239 899 -3238
rect 929 -3239 1606 -3238
rect 1689 -3239 1795 -3238
rect 1815 -3239 1844 -3238
rect 1962 -3239 1977 -3238
rect 100 -3241 227 -3240
rect 247 -3241 276 -3240
rect 282 -3241 416 -3240
rect 464 -3241 871 -3240
rect 873 -3241 1466 -3240
rect 1528 -3241 1606 -3240
rect 1703 -3241 1802 -3240
rect 1815 -3241 1851 -3240
rect 128 -3243 188 -3242
rect 191 -3243 1585 -3242
rect 1598 -3243 1634 -3242
rect 1717 -3243 1739 -3242
rect 1745 -3243 1774 -3242
rect 1822 -3243 1837 -3242
rect 135 -3245 720 -3244
rect 751 -3245 944 -3244
rect 957 -3245 997 -3244
rect 1104 -3245 1221 -3244
rect 1237 -3245 1620 -3244
rect 1717 -3245 1732 -3244
rect 1759 -3245 1767 -3244
rect 156 -3247 171 -3246
rect 191 -3247 1648 -3246
rect 1731 -3247 1753 -3246
rect 205 -3249 213 -3248
rect 215 -3249 1070 -3248
rect 1108 -3249 1683 -3248
rect 1724 -3249 1753 -3248
rect 219 -3251 804 -3250
rect 814 -3251 1011 -3250
rect 1108 -3251 1130 -3250
rect 1216 -3251 1410 -3250
rect 1465 -3251 1655 -3250
rect 219 -3253 416 -3252
rect 464 -3253 507 -3252
rect 513 -3253 615 -3252
rect 632 -3253 1130 -3252
rect 1216 -3253 1347 -3252
rect 1353 -3253 1592 -3252
rect 1654 -3253 1697 -3252
rect 240 -3255 507 -3254
rect 576 -3255 1651 -3254
rect 240 -3257 640 -3256
rect 653 -3257 689 -3256
rect 716 -3257 1333 -3256
rect 1346 -3257 1487 -3256
rect 1549 -3257 1592 -3256
rect 247 -3259 262 -3258
rect 282 -3259 661 -3258
rect 674 -3259 703 -3258
rect 716 -3259 993 -3258
rect 1080 -3259 1354 -3258
rect 1374 -3259 1445 -3258
rect 1472 -3259 1529 -3258
rect 1563 -3259 1662 -3258
rect 254 -3261 262 -3260
rect 331 -3261 745 -3260
rect 751 -3261 808 -3260
rect 856 -3261 983 -3260
rect 985 -3261 1270 -3260
rect 1290 -3261 1459 -3260
rect 1486 -3261 1581 -3260
rect 1661 -3261 1676 -3260
rect 268 -3263 332 -3262
rect 338 -3263 727 -3262
rect 772 -3263 794 -3262
rect 807 -3263 948 -3262
rect 957 -3263 1165 -3262
rect 1167 -3263 1473 -3262
rect 268 -3265 290 -3264
rect 338 -3265 605 -3264
rect 653 -3265 696 -3264
rect 702 -3265 1256 -3264
rect 1269 -3265 1613 -3264
rect 289 -3267 346 -3266
rect 352 -3267 419 -3266
rect 485 -3267 514 -3266
rect 562 -3267 857 -3266
rect 863 -3267 871 -3266
rect 898 -3267 1095 -3266
rect 1115 -3267 1235 -3266
rect 1237 -3267 1686 -3266
rect 345 -3269 647 -3268
rect 660 -3269 668 -3268
rect 695 -3269 731 -3268
rect 793 -3269 1032 -3268
rect 1115 -3269 1193 -3268
rect 1220 -3269 1494 -3268
rect 352 -3271 444 -3270
rect 485 -3271 787 -3270
rect 912 -3271 1011 -3270
rect 1031 -3271 1151 -3270
rect 1171 -3271 1256 -3270
rect 1290 -3271 1312 -3270
rect 1332 -3271 1340 -3270
rect 1374 -3271 1515 -3270
rect 229 -3273 444 -3272
rect 495 -3273 580 -3272
rect 583 -3273 640 -3272
rect 646 -3273 682 -3272
rect 786 -3273 1060 -3272
rect 1066 -3273 1494 -3272
rect 1500 -3273 1515 -3272
rect 359 -3275 423 -3274
rect 499 -3275 734 -3274
rect 912 -3275 934 -3274
rect 947 -3275 1004 -3274
rect 1059 -3275 1179 -3274
rect 1192 -3275 1263 -3274
rect 1283 -3275 1501 -3274
rect 177 -3277 500 -3276
rect 527 -3277 682 -3276
rect 709 -3277 1004 -3276
rect 1066 -3277 1228 -3276
rect 1262 -3277 1557 -3276
rect 177 -3279 199 -3278
rect 359 -3279 437 -3278
rect 527 -3279 818 -3278
rect 919 -3279 934 -3278
rect 968 -3279 997 -3278
rect 1150 -3279 1298 -3278
rect 1311 -3279 1319 -3278
rect 1409 -3279 1854 -3278
rect 163 -3281 199 -3280
rect 366 -3281 423 -3280
rect 555 -3281 1340 -3280
rect 1458 -3281 1543 -3280
rect 1853 -3281 1865 -3280
rect 142 -3283 164 -3282
rect 324 -3283 367 -3282
rect 373 -3283 437 -3282
rect 478 -3283 556 -3282
rect 562 -3283 598 -3282
rect 604 -3283 738 -3282
rect 919 -3283 955 -3282
rect 968 -3283 1123 -3282
rect 1157 -3283 1228 -3282
rect 1283 -3283 1382 -3282
rect 1535 -3283 1557 -3282
rect 1864 -3283 1893 -3282
rect 117 -3285 143 -3284
rect 310 -3285 598 -3284
rect 667 -3285 780 -3284
rect 1122 -3285 1207 -3284
rect 1297 -3285 1368 -3284
rect 1892 -3285 1907 -3284
rect 310 -3287 318 -3286
rect 324 -3287 430 -3286
rect 576 -3287 941 -3286
rect 1143 -3287 1158 -3286
rect 1171 -3287 1389 -3286
rect 1906 -3287 1921 -3286
rect 317 -3289 626 -3288
rect 709 -3289 836 -3288
rect 940 -3289 1025 -3288
rect 1178 -3289 1417 -3288
rect 373 -3291 451 -3290
rect 583 -3291 612 -3290
rect 625 -3291 1095 -3290
rect 1206 -3291 1438 -3290
rect 149 -3293 612 -3292
rect 737 -3293 1018 -3292
rect 1024 -3293 1053 -3292
rect 1318 -3293 1431 -3292
rect 383 -3295 864 -3294
rect 961 -3295 1389 -3294
rect 1402 -3295 1438 -3294
rect 387 -3297 493 -3296
rect 590 -3297 633 -3296
rect 765 -3297 1018 -3296
rect 1038 -3297 1053 -3296
rect 1136 -3297 1403 -3296
rect 387 -3299 472 -3298
rect 590 -3299 1088 -3298
rect 1136 -3299 1200 -3298
rect 1325 -3299 1431 -3298
rect 394 -3301 549 -3300
rect 765 -3301 906 -3300
rect 961 -3301 990 -3300
rect 1038 -3301 1081 -3300
rect 1087 -3301 1186 -3300
rect 1199 -3301 1361 -3300
rect 1367 -3301 1571 -3300
rect 394 -3303 409 -3302
rect 429 -3303 535 -3302
rect 723 -3303 1186 -3302
rect 1325 -3303 1522 -3302
rect 380 -3305 409 -3304
rect 450 -3305 619 -3304
rect 779 -3305 1277 -3304
rect 1451 -3305 1522 -3304
rect 380 -3307 479 -3306
rect 534 -3307 1672 -3306
rect 401 -3309 619 -3308
rect 821 -3309 836 -3308
rect 884 -3309 1361 -3308
rect 1451 -3309 1508 -3308
rect 296 -3311 402 -3310
rect 404 -3311 458 -3310
rect 471 -3311 976 -3310
rect 978 -3311 1144 -3310
rect 1248 -3311 1277 -3310
rect 1423 -3311 1508 -3310
rect 296 -3313 769 -3312
rect 821 -3313 843 -3312
rect 849 -3313 885 -3312
rect 905 -3313 1235 -3312
rect 1248 -3313 1480 -3312
rect 457 -3315 521 -3314
rect 842 -3315 878 -3314
rect 989 -3315 1627 -3314
rect 520 -3317 759 -3316
rect 877 -3317 892 -3316
rect 1304 -3317 1424 -3316
rect 1479 -3317 1725 -3316
rect 758 -3319 850 -3318
rect 1304 -3319 1396 -3318
rect 1626 -3319 1711 -3318
rect 828 -3321 892 -3320
rect 1073 -3321 1396 -3320
rect 828 -3323 927 -3322
rect 1073 -3323 1242 -3322
rect 254 -3325 927 -3324
rect 1045 -3325 1242 -3324
rect 1045 -3327 1102 -3326
rect 142 -3338 174 -3337
rect 177 -3338 237 -3337
rect 257 -3338 374 -3337
rect 394 -3338 538 -3337
rect 541 -3338 545 -3337
rect 590 -3338 780 -3337
rect 814 -3338 1126 -3337
rect 1160 -3338 1228 -3337
rect 1234 -3338 1452 -3337
rect 1521 -3338 1585 -3337
rect 1591 -3338 1613 -3337
rect 1647 -3338 1662 -3337
rect 1717 -3338 1728 -3337
rect 1752 -3338 1760 -3337
rect 1766 -3338 1770 -3337
rect 1787 -3338 1812 -3337
rect 1829 -3338 1844 -3337
rect 1885 -3338 1907 -3337
rect 1955 -3338 1963 -3337
rect 2025 -3338 2029 -3337
rect 163 -3340 391 -3339
rect 415 -3340 486 -3339
rect 488 -3340 507 -3339
rect 513 -3340 993 -3339
rect 1034 -3340 1221 -3339
rect 1234 -3340 1284 -3339
rect 1339 -3340 1459 -3339
rect 1521 -3340 1529 -3339
rect 1549 -3340 1627 -3339
rect 1724 -3340 1746 -3339
rect 1787 -3340 1851 -3339
rect 1888 -3340 1893 -3339
rect 1962 -3340 1970 -3339
rect 2025 -3340 2033 -3339
rect 170 -3342 181 -3341
rect 212 -3342 409 -3341
rect 429 -3342 927 -3341
rect 968 -3342 1333 -3341
rect 1367 -3342 1494 -3341
rect 1528 -3342 1564 -3341
rect 1605 -3342 1655 -3341
rect 1794 -3342 1823 -3341
rect 1836 -3342 1844 -3341
rect 1850 -3342 1858 -3341
rect 215 -3344 804 -3343
rect 821 -3344 937 -3343
rect 968 -3344 1004 -3343
rect 1031 -3344 1221 -3343
rect 1237 -3344 1298 -3343
rect 1332 -3344 1375 -3343
rect 1381 -3344 1445 -3343
rect 1451 -3344 1487 -3343
rect 1552 -3344 1599 -3343
rect 1608 -3344 1669 -3343
rect 1801 -3344 1837 -3343
rect 1857 -3344 1872 -3343
rect 240 -3346 507 -3345
rect 541 -3346 577 -3345
rect 597 -3346 1084 -3345
rect 1097 -3346 1312 -3345
rect 1374 -3346 1459 -3345
rect 1556 -3346 1588 -3345
rect 1654 -3346 1854 -3345
rect 1864 -3346 1872 -3345
rect 275 -3348 374 -3347
rect 422 -3348 430 -3347
rect 474 -3348 1371 -3347
rect 1384 -3348 1424 -3347
rect 1801 -3348 1816 -3347
rect 1864 -3348 1879 -3347
rect 2028 -3348 2033 -3347
rect 205 -3350 423 -3349
rect 548 -3350 1032 -3349
rect 1066 -3350 1431 -3349
rect 282 -3352 860 -3351
rect 877 -3352 1004 -3351
rect 1080 -3352 1137 -3351
rect 1199 -3352 1228 -3351
rect 1269 -3352 1354 -3351
rect 1388 -3352 1420 -3351
rect 296 -3354 384 -3353
rect 492 -3354 549 -3353
rect 555 -3354 591 -3353
rect 597 -3354 647 -3353
rect 653 -3354 878 -3353
rect 891 -3354 955 -3353
rect 961 -3354 1081 -3353
rect 1101 -3354 1179 -3353
rect 1199 -3354 1326 -3353
rect 1416 -3354 1438 -3353
rect 268 -3356 297 -3355
rect 317 -3356 409 -3355
rect 450 -3356 493 -3355
rect 534 -3356 647 -3355
rect 674 -3356 1028 -3355
rect 1045 -3356 1179 -3355
rect 1213 -3356 1403 -3355
rect 359 -3358 514 -3357
rect 534 -3358 584 -3357
rect 618 -3358 640 -3357
rect 660 -3358 675 -3357
rect 681 -3358 1067 -3357
rect 1157 -3358 1214 -3357
rect 1269 -3358 1473 -3357
rect 303 -3360 360 -3359
rect 366 -3360 395 -3359
rect 478 -3360 556 -3359
rect 562 -3360 682 -3359
rect 723 -3360 1396 -3359
rect 1472 -3360 1515 -3359
rect 331 -3362 479 -3361
rect 562 -3362 727 -3361
rect 730 -3362 1809 -3361
rect 198 -3364 332 -3363
rect 345 -3364 661 -3363
rect 723 -3364 759 -3363
rect 772 -3364 815 -3363
rect 821 -3364 1060 -3363
rect 1272 -3364 1284 -3363
rect 1290 -3364 1298 -3363
rect 289 -3366 346 -3365
rect 387 -3366 451 -3365
rect 583 -3366 668 -3365
rect 737 -3366 962 -3365
rect 978 -3366 1025 -3365
rect 1045 -3366 1144 -3365
rect 1255 -3366 1291 -3365
rect 219 -3368 388 -3367
rect 443 -3368 731 -3367
rect 751 -3368 1095 -3367
rect 1192 -3368 1256 -3367
rect 352 -3370 668 -3369
rect 772 -3370 801 -3369
rect 835 -3370 850 -3369
rect 852 -3370 1011 -3369
rect 1024 -3370 1039 -3369
rect 1059 -3370 1074 -3369
rect 1094 -3370 1242 -3369
rect 401 -3372 444 -3371
rect 471 -3372 738 -3371
rect 779 -3372 976 -3371
rect 982 -3372 1105 -3371
rect 1192 -3372 1466 -3371
rect 401 -3374 752 -3373
rect 793 -3374 836 -3373
rect 842 -3374 958 -3373
rect 989 -3374 1361 -3373
rect 1465 -3374 1508 -3373
rect 600 -3376 1074 -3375
rect 1241 -3376 1305 -3375
rect 1346 -3376 1361 -3375
rect 604 -3378 759 -3377
rect 800 -3378 1378 -3377
rect 604 -3380 612 -3379
rect 618 -3380 710 -3379
rect 842 -3380 1207 -3379
rect 1318 -3380 1347 -3379
rect 520 -3382 710 -3381
rect 849 -3382 1151 -3381
rect 1185 -3382 1305 -3381
rect 418 -3384 521 -3383
rect 527 -3384 612 -3383
rect 625 -3384 654 -3383
rect 688 -3384 794 -3383
rect 856 -3384 983 -3383
rect 989 -3384 1249 -3383
rect 457 -3386 626 -3385
rect 688 -3386 787 -3385
rect 870 -3386 976 -3385
rect 1108 -3386 1207 -3385
rect 1209 -3386 1249 -3385
rect 310 -3388 458 -3387
rect 527 -3388 570 -3387
rect 786 -3388 885 -3387
rect 891 -3388 1123 -3387
rect 1185 -3388 1480 -3387
rect 184 -3390 570 -3389
rect 807 -3390 1109 -3389
rect 1122 -3390 1382 -3389
rect 261 -3392 311 -3391
rect 695 -3392 808 -3391
rect 863 -3392 885 -3391
rect 898 -3392 1039 -3391
rect 324 -3394 696 -3393
rect 744 -3394 864 -3393
rect 870 -3394 906 -3393
rect 919 -3394 1011 -3393
rect 702 -3396 745 -3395
rect 901 -3396 1277 -3395
rect 464 -3398 703 -3397
rect 905 -3398 1116 -3397
rect 436 -3400 465 -3399
rect 912 -3400 920 -3399
rect 926 -3400 1130 -3399
rect 380 -3402 437 -3401
rect 765 -3402 913 -3401
rect 940 -3402 1144 -3401
rect 247 -3404 381 -3403
rect 632 -3404 766 -3403
rect 940 -3404 1217 -3403
rect 499 -3406 633 -3405
rect 947 -3406 1137 -3405
rect 338 -3408 500 -3407
rect 828 -3408 948 -3407
rect 954 -3408 997 -3407
rect 1052 -3408 1116 -3407
rect 191 -3410 339 -3409
rect 828 -3410 934 -3409
rect 996 -3410 1172 -3409
rect 933 -3412 1018 -3411
rect 1052 -3412 1088 -3411
rect 1171 -3412 1263 -3411
rect 971 -3414 1018 -3413
rect 1087 -3414 1165 -3413
rect 1262 -3414 1410 -3413
rect 173 -3425 269 -3424
rect 296 -3425 318 -3424
rect 338 -3425 475 -3424
rect 478 -3425 594 -3424
rect 621 -3425 633 -3424
rect 639 -3425 724 -3424
rect 726 -3425 941 -3424
rect 961 -3425 1207 -3424
rect 1213 -3425 1287 -3424
rect 1297 -3425 1308 -3424
rect 1311 -3425 1333 -3424
rect 1346 -3425 1375 -3424
rect 1437 -3425 1452 -3424
rect 1458 -3425 1494 -3424
rect 1514 -3425 1529 -3424
rect 1584 -3425 1809 -3424
rect 1822 -3425 1861 -3424
rect 170 -3427 174 -3426
rect 310 -3427 325 -3426
rect 345 -3427 391 -3426
rect 394 -3427 402 -3426
rect 404 -3427 416 -3426
rect 429 -3427 468 -3426
rect 492 -3427 629 -3426
rect 646 -3427 724 -3426
rect 758 -3427 801 -3426
rect 807 -3427 843 -3426
rect 884 -3427 923 -3426
rect 975 -3427 1025 -3426
rect 1066 -3427 1200 -3426
rect 1206 -3427 1235 -3426
rect 1248 -3427 1308 -3426
rect 1321 -3427 1333 -3426
rect 1444 -3427 1466 -3426
rect 1612 -3427 1630 -3426
rect 1640 -3427 1648 -3426
rect 1724 -3427 1728 -3426
rect 1738 -3427 1749 -3426
rect 1759 -3427 1767 -3426
rect 1794 -3427 1802 -3426
rect 1822 -3427 1830 -3426
rect 1857 -3427 1868 -3426
rect 373 -3429 472 -3428
rect 492 -3429 563 -3428
rect 611 -3429 640 -3428
rect 653 -3429 657 -3428
rect 684 -3429 717 -3428
rect 744 -3429 759 -3428
rect 807 -3429 990 -3428
rect 992 -3429 1053 -3428
rect 1066 -3429 1102 -3428
rect 1108 -3429 1200 -3428
rect 1220 -3429 1459 -3428
rect 1461 -3429 1655 -3428
rect 1724 -3429 1732 -3428
rect 1766 -3429 1788 -3428
rect 1829 -3429 1844 -3428
rect 1857 -3429 1865 -3428
rect 408 -3431 489 -3430
rect 499 -3431 612 -3430
rect 625 -3431 668 -3430
rect 695 -3431 1032 -3430
rect 1052 -3431 1088 -3430
rect 1101 -3431 1186 -3430
rect 1255 -3431 1319 -3430
rect 1325 -3431 1368 -3430
rect 1381 -3431 1466 -3430
rect 1836 -3431 1844 -3430
rect 1864 -3431 1872 -3430
rect 450 -3433 486 -3432
rect 506 -3433 647 -3432
rect 653 -3433 689 -3432
rect 702 -3433 923 -3432
rect 1003 -3433 1032 -3432
rect 1069 -3433 1126 -3432
rect 1136 -3433 1221 -3432
rect 1276 -3433 1284 -3432
rect 1451 -3433 1473 -3432
rect 422 -3435 507 -3434
rect 548 -3435 580 -3434
rect 660 -3435 696 -3434
rect 702 -3435 787 -3434
rect 814 -3435 846 -3434
rect 863 -3435 885 -3434
rect 901 -3435 1095 -3434
rect 1108 -3435 1193 -3434
rect 1867 -3435 1872 -3434
rect 380 -3437 423 -3436
rect 464 -3437 500 -3436
rect 555 -3437 605 -3436
rect 660 -3437 706 -3436
rect 709 -3437 899 -3436
rect 912 -3437 976 -3436
rect 1010 -3437 1123 -3436
rect 1143 -3437 1235 -3436
rect 331 -3439 465 -3438
rect 541 -3439 556 -3438
rect 558 -3439 780 -3438
rect 814 -3439 829 -3438
rect 835 -3439 860 -3438
rect 915 -3439 969 -3438
rect 982 -3439 1011 -3438
rect 1034 -3439 1095 -3438
rect 1115 -3439 1182 -3438
rect 1185 -3439 1263 -3438
rect 359 -3441 381 -3440
rect 541 -3441 619 -3440
rect 674 -3441 710 -3440
rect 737 -3441 829 -3440
rect 835 -3441 871 -3440
rect 919 -3441 955 -3440
rect 1073 -3441 1249 -3440
rect 562 -3443 598 -3442
rect 604 -3443 626 -3442
rect 681 -3443 738 -3442
rect 744 -3443 822 -3442
rect 842 -3443 892 -3442
rect 947 -3443 1004 -3442
rect 1059 -3443 1074 -3442
rect 1080 -3443 1130 -3442
rect 1164 -3443 1627 -3442
rect 520 -3445 682 -3444
rect 751 -3445 1126 -3444
rect 1192 -3445 1242 -3444
rect 436 -3447 521 -3446
rect 569 -3447 717 -3446
rect 751 -3447 850 -3446
rect 877 -3447 1081 -3446
rect 1083 -3447 1172 -3446
rect 1227 -3447 1242 -3446
rect 527 -3449 570 -3448
rect 583 -3449 598 -3448
rect 632 -3449 1060 -3448
rect 1087 -3449 1305 -3448
rect 513 -3451 584 -3450
rect 590 -3451 675 -3450
rect 730 -3451 850 -3450
rect 877 -3451 906 -3450
rect 954 -3451 997 -3450
rect 1171 -3451 1270 -3450
rect 457 -3453 514 -3452
rect 730 -3453 927 -3452
rect 996 -3453 1046 -3452
rect 1178 -3453 1228 -3452
rect 443 -3455 458 -3454
rect 590 -3455 1046 -3454
rect 1178 -3455 1214 -3454
rect 439 -3457 444 -3456
rect 765 -3457 822 -3456
rect 772 -3459 780 -3458
rect 271 -3470 367 -3469
rect 369 -3470 395 -3469
rect 415 -3470 430 -3469
rect 439 -3470 444 -3469
rect 457 -3470 465 -3469
rect 478 -3470 493 -3469
rect 499 -3470 552 -3469
rect 569 -3470 640 -3469
rect 642 -3470 752 -3469
rect 765 -3470 808 -3469
rect 828 -3470 913 -3469
rect 919 -3470 955 -3469
rect 975 -3470 979 -3469
rect 1031 -3470 1063 -3469
rect 1080 -3470 1109 -3469
rect 1122 -3470 1186 -3469
rect 1199 -3470 1319 -3469
rect 1430 -3470 1445 -3469
rect 1458 -3470 1571 -3469
rect 1745 -3470 1767 -3469
rect 1790 -3470 1795 -3469
rect 1829 -3470 1837 -3469
rect 1839 -3470 1851 -3469
rect 1860 -3470 1865 -3469
rect 1958 -3470 1963 -3469
rect 2025 -3470 2029 -3469
rect 324 -3472 332 -3471
rect 380 -3472 388 -3471
rect 422 -3472 468 -3471
rect 485 -3472 524 -3471
rect 541 -3472 570 -3471
rect 579 -3472 605 -3471
rect 618 -3472 629 -3471
rect 639 -3472 654 -3471
rect 667 -3472 706 -3471
rect 730 -3472 738 -3471
rect 772 -3472 780 -3471
rect 789 -3472 815 -3471
rect 828 -3472 843 -3471
rect 849 -3472 923 -3471
rect 975 -3472 997 -3471
rect 1017 -3472 1032 -3471
rect 1059 -3472 1074 -3471
rect 1083 -3472 1172 -3471
rect 1178 -3472 1207 -3471
rect 1213 -3472 1273 -3471
rect 1276 -3472 1287 -3471
rect 1307 -3472 1312 -3471
rect 1433 -3472 1452 -3471
rect 1500 -3472 1504 -3471
rect 1507 -3472 1515 -3471
rect 1843 -3472 1851 -3471
rect 1864 -3472 1872 -3471
rect 2025 -3472 2033 -3471
rect 471 -3474 524 -3473
rect 562 -3474 605 -3473
rect 653 -3474 745 -3473
rect 800 -3474 888 -3473
rect 1010 -3474 1018 -3473
rect 1045 -3474 1501 -3473
rect 1822 -3474 1844 -3473
rect 2028 -3474 2033 -3473
rect 485 -3476 633 -3475
rect 674 -3476 703 -3475
rect 709 -3476 745 -3475
rect 814 -3476 836 -3475
rect 866 -3476 1088 -3475
rect 1094 -3476 1126 -3475
rect 1129 -3476 1144 -3475
rect 1178 -3476 1193 -3475
rect 1234 -3476 1263 -3475
rect 1269 -3476 1326 -3475
rect 1493 -3476 1515 -3475
rect 506 -3478 542 -3477
rect 590 -3478 598 -3477
rect 632 -3478 661 -3477
rect 681 -3478 752 -3477
rect 821 -3478 843 -3477
rect 870 -3478 878 -3477
rect 884 -3478 916 -3477
rect 1003 -3478 1011 -3477
rect 1038 -3478 1046 -3477
rect 1059 -3478 1102 -3477
rect 1157 -3478 1193 -3477
rect 1220 -3478 1235 -3477
rect 1255 -3478 1305 -3477
rect 1311 -3478 1333 -3477
rect 1465 -3478 1494 -3477
rect 520 -3480 899 -3479
rect 1024 -3480 1039 -3479
rect 1248 -3480 1305 -3479
rect 534 -3482 591 -3481
rect 611 -3482 682 -3481
rect 695 -3482 787 -3481
rect 1024 -3482 1165 -3481
rect 1241 -3482 1249 -3481
rect 1283 -3482 1291 -3481
rect 513 -3484 535 -3483
rect 555 -3484 612 -3483
rect 716 -3484 780 -3483
rect 1227 -3484 1242 -3483
rect 1290 -3484 1728 -3483
rect 688 -3486 717 -3485
rect 737 -3486 759 -3485
rect 723 -3488 759 -3487
rect 331 -3499 339 -3498
rect 394 -3499 430 -3498
rect 432 -3499 472 -3498
rect 523 -3499 654 -3498
rect 681 -3499 710 -3498
rect 716 -3499 731 -3498
rect 775 -3499 892 -3498
rect 968 -3499 976 -3498
rect 996 -3499 1004 -3498
rect 1038 -3499 1063 -3498
rect 1122 -3499 1291 -3498
rect 1304 -3499 1368 -3498
rect 1430 -3499 1438 -3498
rect 1500 -3499 1508 -3498
rect 1570 -3499 1613 -3498
rect 1724 -3499 1732 -3498
rect 1780 -3499 1791 -3498
rect 1850 -3499 1861 -3498
rect 387 -3501 395 -3500
rect 429 -3501 486 -3500
rect 534 -3501 549 -3500
rect 569 -3501 577 -3500
rect 625 -3501 633 -3500
rect 646 -3501 657 -3500
rect 779 -3501 801 -3500
rect 810 -3501 829 -3500
rect 842 -3501 867 -3500
rect 884 -3501 1025 -3500
rect 1038 -3501 1046 -3500
rect 1143 -3501 1151 -3500
rect 1160 -3501 1179 -3500
rect 1192 -3501 1207 -3500
rect 1234 -3501 1252 -3500
rect 1262 -3501 1277 -3500
rect 1283 -3501 1312 -3500
rect 1493 -3501 1508 -3500
rect 1843 -3501 1851 -3500
rect 1857 -3501 1865 -3500
rect 611 -3503 633 -3502
rect 751 -3503 780 -3502
rect 789 -3503 815 -3502
rect 863 -3503 871 -3502
rect 898 -3503 1025 -3502
rect 1031 -3503 1046 -3502
rect 1234 -3503 1256 -3502
rect 611 -3505 619 -3504
rect 751 -3505 759 -3504
rect 1031 -3505 1060 -3504
rect 1241 -3505 1249 -3504
rect 604 -3507 619 -3506
rect 744 -3507 759 -3506
rect 1059 -3507 1067 -3506
rect 590 -3509 605 -3508
rect 744 -3509 766 -3508
rect 1066 -3509 1081 -3508
rect 765 -3511 773 -3510
rect 408 -3522 430 -3521
rect 618 -3522 636 -3521
rect 709 -3522 717 -3521
rect 723 -3522 738 -3521
rect 751 -3522 787 -3521
rect 800 -3522 811 -3521
rect 891 -3522 927 -3521
rect 968 -3522 972 -3521
rect 1017 -3522 1028 -3521
rect 1038 -3522 1042 -3521
rect 1059 -3522 1067 -3521
rect 1150 -3522 1158 -3521
rect 1206 -3522 1214 -3521
rect 1223 -3522 1235 -3521
rect 1360 -3522 1368 -3521
rect 1507 -3522 1511 -3521
rect 1612 -3522 1634 -3521
rect 1850 -3522 1858 -3521
rect 611 -3524 619 -3523
rect 632 -3524 647 -3523
rect 709 -3524 741 -3523
rect 758 -3524 776 -3523
rect 779 -3524 787 -3523
rect 1024 -3524 1161 -3523
rect 1507 -3524 1515 -3523
rect 604 -3526 612 -3525
rect 765 -3526 790 -3525
rect 1010 -3526 1025 -3525
rect 1038 -3526 1046 -3525
rect 1052 -3526 1060 -3525
rect 1066 -3526 1123 -3525
rect 604 -3528 626 -3527
rect 765 -3528 773 -3527
rect 1003 -3528 1011 -3527
rect 1510 -3528 1515 -3527
rect 625 -3530 633 -3529
rect 394 -3541 402 -3540
rect 464 -3541 475 -3540
rect 548 -3541 556 -3540
rect 583 -3541 591 -3540
rect 635 -3541 640 -3540
rect 702 -3541 710 -3540
rect 730 -3541 741 -3540
rect 758 -3541 766 -3540
rect 786 -3541 790 -3540
rect 926 -3541 969 -3540
rect 1010 -3541 1021 -3540
rect 1027 -3541 1032 -3540
rect 1038 -3541 1046 -3540
rect 1213 -3541 1224 -3540
rect 1507 -3541 1511 -3540
rect 1640 -3541 1648 -3540
rect 471 -3543 479 -3542
rect 576 -3543 584 -3542
rect 730 -3543 745 -3542
rect 1038 -3543 1067 -3542
rect 1507 -3543 1522 -3542
rect 1633 -3543 1641 -3542
rect 1510 -3545 1522 -3544
rect 401 -3556 405 -3555
rect 541 -3556 549 -3555
rect 551 -3556 556 -3555
rect 586 -3556 591 -3555
rect 604 -3556 608 -3555
rect 646 -3556 650 -3555
rect 789 -3556 794 -3555
rect 1017 -3556 1039 -3555
rect 1059 -3556 1067 -3555
rect 1517 -3556 1522 -3555
rect 2028 -3556 2033 -3555
rect 401 -3558 409 -3557
rect 604 -3558 612 -3557
rect 1514 -3558 1522 -3557
rect 607 -3560 612 -3559
rect 1507 -3560 1515 -3559
rect 401 -3571 405 -3570
rect 1062 -3571 1067 -3570
rect 1514 -3571 1522 -3570
rect 401 -3573 409 -3572
rect 404 -3575 409 -3574
rect 394 -3586 402 -3585
rect 618 -3586 622 -3585
rect 723 -3586 727 -3585
rect 401 -3588 409 -3587
rect 716 -3588 724 -3587
rect 723 -3599 731 -3598
rect 695 -3610 706 -3609
rect 1640 -3610 1644 -3609
rect 758 -3621 766 -3620
rect 1640 -3621 1648 -3620
rect 761 -3632 766 -3631
rect 394 -3654 398 -3653
rect 695 -3654 699 -3653
rect 394 -3656 402 -3655
rect 397 -3658 402 -3657
rect 397 -3669 402 -3668
rect 604 -3669 612 -3668
<< m2contact >>
rect 254 0 255 1
rect 432 0 433 1
rect 485 0 486 1
rect 632 0 633 1
rect 635 0 636 1
rect 772 0 773 1
rect 796 0 797 1
rect 814 0 815 1
rect 824 0 825 1
rect 961 0 962 1
rect 968 0 969 1
rect 1206 0 1207 1
rect 352 -2 353 -1
rect 572 -2 573 -1
rect 576 -2 577 -1
rect 681 -2 682 -1
rect 688 -2 689 -1
rect 765 -2 766 -1
rect 800 -2 801 -1
rect 891 -2 892 -1
rect 978 -2 979 -1
rect 982 -2 983 -1
rect 1038 -2 1039 -1
rect 1437 -2 1438 -1
rect 397 -4 398 -3
rect 548 -4 549 -3
rect 555 -4 556 -3
rect 583 -4 584 -3
rect 604 -4 605 -3
rect 842 -4 843 -3
rect 863 -4 864 -3
rect 919 -4 920 -3
rect 1073 -4 1074 -3
rect 1129 -4 1130 -3
rect 415 -6 416 -5
rect 422 -6 423 -5
rect 611 -6 612 -5
rect 625 -6 626 -5
rect 639 -6 640 -5
rect 845 -6 846 -5
rect 884 -6 885 -5
rect 1087 -6 1088 -5
rect 1094 -6 1095 -5
rect 1125 -6 1126 -5
rect 618 -8 619 -7
rect 852 -8 853 -7
rect 646 -10 647 -9
rect 705 -10 706 -9
rect 709 -10 710 -9
rect 915 -10 916 -9
rect 663 -12 664 -11
rect 989 -12 990 -11
rect 716 -14 717 -13
rect 821 -14 822 -13
rect 828 -14 829 -13
rect 887 -14 888 -13
rect 730 -16 731 -15
rect 803 -16 804 -15
rect 810 -16 811 -15
rect 870 -16 871 -15
rect 835 -18 836 -17
rect 859 -18 860 -17
rect 184 -29 185 -28
rect 212 -29 213 -28
rect 240 -29 241 -28
rect 397 -29 398 -28
rect 404 -29 405 -28
rect 478 -29 479 -28
rect 492 -29 493 -28
rect 618 -29 619 -28
rect 646 -29 647 -28
rect 723 -29 724 -28
rect 737 -29 738 -28
rect 758 -29 759 -28
rect 765 -29 766 -28
rect 828 -29 829 -28
rect 842 -29 843 -28
rect 1220 -29 1221 -28
rect 1234 -29 1235 -28
rect 1360 -29 1361 -28
rect 1437 -29 1438 -28
rect 1486 -29 1487 -28
rect 1629 -29 1630 -28
rect 1633 -29 1634 -28
rect 198 -31 199 -30
rect 254 -31 255 -30
rect 275 -31 276 -30
rect 313 -31 314 -30
rect 317 -31 318 -30
rect 660 -31 661 -30
rect 667 -31 668 -30
rect 740 -31 741 -30
rect 744 -31 745 -30
rect 863 -31 864 -30
rect 870 -31 871 -30
rect 884 -31 885 -30
rect 908 -31 909 -30
rect 947 -31 948 -30
rect 961 -31 962 -30
rect 1045 -31 1046 -30
rect 1066 -31 1067 -30
rect 1101 -31 1102 -30
rect 1108 -31 1109 -30
rect 1150 -31 1151 -30
rect 1206 -31 1207 -30
rect 1290 -31 1291 -30
rect 1321 -31 1322 -30
rect 1332 -31 1333 -30
rect 1440 -31 1441 -30
rect 1759 -31 1760 -30
rect 296 -33 297 -32
rect 352 -33 353 -32
rect 355 -33 356 -32
rect 464 -33 465 -32
rect 471 -33 472 -32
rect 611 -33 612 -32
rect 618 -33 619 -32
rect 625 -33 626 -32
rect 660 -33 661 -32
rect 695 -33 696 -32
rect 702 -33 703 -32
rect 821 -33 822 -32
rect 828 -33 829 -32
rect 1038 -33 1039 -32
rect 1087 -33 1088 -32
rect 1178 -33 1179 -32
rect 394 -35 395 -34
rect 485 -35 486 -34
rect 499 -35 500 -34
rect 639 -35 640 -34
rect 677 -35 678 -34
rect 975 -35 976 -34
rect 978 -35 979 -34
rect 1003 -35 1004 -34
rect 1010 -35 1011 -34
rect 1094 -35 1095 -34
rect 1132 -35 1133 -34
rect 1213 -35 1214 -34
rect 415 -37 416 -36
rect 422 -37 423 -36
rect 432 -37 433 -36
rect 590 -37 591 -36
rect 611 -37 612 -36
rect 656 -37 657 -36
rect 702 -37 703 -36
rect 716 -37 717 -36
rect 751 -37 752 -36
rect 887 -37 888 -36
rect 912 -37 913 -36
rect 1017 -37 1018 -36
rect 1073 -37 1074 -36
rect 1087 -37 1088 -36
rect 1094 -37 1095 -36
rect 1115 -37 1116 -36
rect 422 -39 423 -38
rect 446 -39 447 -38
rect 485 -39 486 -38
rect 604 -39 605 -38
rect 639 -39 640 -38
rect 653 -39 654 -38
rect 716 -39 717 -38
rect 807 -39 808 -38
rect 842 -39 843 -38
rect 898 -39 899 -38
rect 926 -39 927 -38
rect 1125 -39 1126 -38
rect 506 -41 507 -40
rect 852 -41 853 -40
rect 856 -41 857 -40
rect 1038 -41 1039 -40
rect 520 -43 521 -42
rect 576 -43 577 -42
rect 583 -43 584 -42
rect 646 -43 647 -42
rect 653 -43 654 -42
rect 961 -43 962 -42
rect 982 -43 983 -42
rect 1031 -43 1032 -42
rect 534 -45 535 -44
rect 688 -45 689 -44
rect 768 -45 769 -44
rect 863 -45 864 -44
rect 870 -45 871 -44
rect 919 -45 920 -44
rect 982 -45 983 -44
rect 1069 -45 1070 -44
rect 548 -47 549 -46
rect 597 -47 598 -46
rect 604 -47 605 -46
rect 901 -47 902 -46
rect 989 -47 990 -46
rect 1059 -47 1060 -46
rect 548 -49 549 -48
rect 572 -49 573 -48
rect 583 -49 584 -48
rect 933 -49 934 -48
rect 1024 -49 1025 -48
rect 1073 -49 1074 -48
rect 569 -51 570 -50
rect 779 -51 780 -50
rect 793 -51 794 -50
rect 835 -51 836 -50
rect 849 -51 850 -50
rect 1080 -51 1081 -50
rect 569 -53 570 -52
rect 674 -53 675 -52
rect 688 -53 689 -52
rect 709 -53 710 -52
rect 772 -53 773 -52
rect 835 -53 836 -52
rect 849 -53 850 -52
rect 912 -53 913 -52
rect 709 -55 710 -54
rect 730 -55 731 -54
rect 772 -55 773 -54
rect 810 -55 811 -54
rect 877 -55 878 -54
rect 940 -55 941 -54
rect 730 -57 731 -56
rect 968 -57 969 -56
rect 800 -59 801 -58
rect 919 -59 920 -58
rect 807 -61 808 -60
rect 814 -61 815 -60
rect 887 -61 888 -60
rect 1052 -61 1053 -60
rect 681 -63 682 -62
rect 814 -63 815 -62
rect 891 -63 892 -62
rect 989 -63 990 -62
rect 565 -65 566 -64
rect 681 -65 682 -64
rect 803 -65 804 -64
rect 891 -65 892 -64
rect 915 -65 916 -64
rect 968 -65 969 -64
rect 58 -76 59 -75
rect 523 -76 524 -75
rect 530 -76 531 -75
rect 1241 -76 1242 -75
rect 1290 -76 1291 -75
rect 1297 -76 1298 -75
rect 1332 -76 1333 -75
rect 1374 -76 1375 -75
rect 1486 -76 1487 -75
rect 1514 -76 1515 -75
rect 1633 -76 1634 -75
rect 1640 -76 1641 -75
rect 1759 -76 1760 -75
rect 1885 -76 1886 -75
rect 65 -78 66 -77
rect 226 -78 227 -77
rect 233 -78 234 -77
rect 849 -78 850 -77
rect 852 -78 853 -77
rect 1136 -78 1137 -77
rect 1157 -78 1158 -77
rect 1167 -78 1168 -77
rect 1171 -78 1172 -77
rect 1269 -78 1270 -77
rect 1360 -78 1361 -77
rect 1423 -78 1424 -77
rect 72 -80 73 -79
rect 401 -80 402 -79
rect 404 -80 405 -79
rect 436 -80 437 -79
rect 450 -80 451 -79
rect 520 -80 521 -79
rect 555 -80 556 -79
rect 660 -80 661 -79
rect 674 -80 675 -79
rect 709 -80 710 -79
rect 740 -80 741 -79
rect 1325 -80 1326 -79
rect 79 -82 80 -81
rect 352 -82 353 -81
rect 359 -82 360 -81
rect 422 -82 423 -81
rect 429 -82 430 -81
rect 604 -82 605 -81
rect 625 -82 626 -81
rect 828 -82 829 -81
rect 835 -82 836 -81
rect 905 -82 906 -81
rect 919 -82 920 -81
rect 940 -82 941 -81
rect 943 -82 944 -81
rect 1290 -82 1291 -81
rect 1321 -82 1322 -81
rect 1360 -82 1361 -81
rect 86 -84 87 -83
rect 264 -84 265 -83
rect 282 -84 283 -83
rect 499 -84 500 -83
rect 513 -84 514 -83
rect 541 -84 542 -83
rect 562 -84 563 -83
rect 632 -84 633 -83
rect 653 -84 654 -83
rect 765 -84 766 -83
rect 786 -84 787 -83
rect 821 -84 822 -83
rect 856 -84 857 -83
rect 1122 -84 1123 -83
rect 1125 -84 1126 -83
rect 1318 -84 1319 -83
rect 93 -86 94 -85
rect 471 -86 472 -85
rect 499 -86 500 -85
rect 527 -86 528 -85
rect 541 -86 542 -85
rect 611 -86 612 -85
rect 660 -86 661 -85
rect 751 -86 752 -85
rect 779 -86 780 -85
rect 821 -86 822 -85
rect 856 -86 857 -85
rect 1010 -86 1011 -85
rect 1038 -86 1039 -85
rect 1108 -86 1109 -85
rect 1115 -86 1116 -85
rect 1150 -86 1151 -85
rect 1178 -86 1179 -85
rect 1255 -86 1256 -85
rect 100 -88 101 -87
rect 600 -88 601 -87
rect 604 -88 605 -87
rect 618 -88 619 -87
rect 702 -88 703 -87
rect 828 -88 829 -87
rect 863 -88 864 -87
rect 884 -88 885 -87
rect 919 -88 920 -87
rect 968 -88 969 -87
rect 975 -88 976 -87
rect 1283 -88 1284 -87
rect 107 -90 108 -89
rect 184 -90 185 -89
rect 191 -90 192 -89
rect 240 -90 241 -89
rect 247 -90 248 -89
rect 443 -90 444 -89
rect 471 -90 472 -89
rect 975 -90 976 -89
rect 989 -90 990 -89
rect 1192 -90 1193 -89
rect 1213 -90 1214 -89
rect 1304 -90 1305 -89
rect 114 -92 115 -91
rect 236 -92 237 -91
rect 240 -92 241 -91
rect 275 -92 276 -91
rect 296 -92 297 -91
rect 331 -92 332 -91
rect 338 -92 339 -91
rect 649 -92 650 -91
rect 702 -92 703 -91
rect 870 -92 871 -91
rect 898 -92 899 -91
rect 1213 -92 1214 -91
rect 1220 -92 1221 -91
rect 1353 -92 1354 -91
rect 124 -94 125 -93
rect 303 -94 304 -93
rect 310 -94 311 -93
rect 324 -94 325 -93
rect 345 -94 346 -93
rect 544 -94 545 -93
rect 576 -94 577 -93
rect 639 -94 640 -93
rect 709 -94 710 -93
rect 716 -94 717 -93
rect 751 -94 752 -93
rect 1234 -94 1235 -93
rect 1237 -94 1238 -93
rect 1507 -94 1508 -93
rect 128 -96 129 -95
rect 583 -96 584 -95
rect 590 -96 591 -95
rect 611 -96 612 -95
rect 618 -96 619 -95
rect 957 -96 958 -95
rect 961 -96 962 -95
rect 1150 -96 1151 -95
rect 1227 -96 1228 -95
rect 1311 -96 1312 -95
rect 135 -98 136 -97
rect 506 -98 507 -97
rect 583 -98 584 -97
rect 597 -98 598 -97
rect 639 -98 640 -97
rect 835 -98 836 -97
rect 863 -98 864 -97
rect 877 -98 878 -97
rect 954 -98 955 -97
rect 989 -98 990 -97
rect 999 -98 1000 -97
rect 1094 -98 1095 -97
rect 1101 -98 1102 -97
rect 1276 -98 1277 -97
rect 149 -100 150 -99
rect 352 -100 353 -99
rect 366 -100 367 -99
rect 569 -100 570 -99
rect 758 -100 759 -99
rect 898 -100 899 -99
rect 933 -100 934 -99
rect 1101 -100 1102 -99
rect 1118 -100 1119 -99
rect 1185 -100 1186 -99
rect 152 -102 153 -101
rect 289 -102 290 -101
rect 310 -102 311 -101
rect 859 -102 860 -101
rect 870 -102 871 -101
rect 982 -102 983 -101
rect 996 -102 997 -101
rect 1094 -102 1095 -101
rect 156 -104 157 -103
rect 317 -104 318 -103
rect 380 -104 381 -103
rect 492 -104 493 -103
rect 730 -104 731 -103
rect 758 -104 759 -103
rect 779 -104 780 -103
rect 908 -104 909 -103
rect 912 -104 913 -103
rect 982 -104 983 -103
rect 1003 -104 1004 -103
rect 1164 -104 1165 -103
rect 163 -106 164 -105
rect 698 -106 699 -105
rect 789 -106 790 -105
rect 800 -106 801 -105
rect 803 -106 804 -105
rect 954 -106 955 -105
rect 968 -106 969 -105
rect 1017 -106 1018 -105
rect 1027 -106 1028 -105
rect 1234 -106 1235 -105
rect 170 -108 171 -107
rect 408 -108 409 -107
rect 411 -108 412 -107
rect 415 -108 416 -107
rect 422 -108 423 -107
rect 548 -108 549 -107
rect 807 -108 808 -107
rect 1003 -108 1004 -107
rect 1010 -108 1011 -107
rect 1143 -108 1144 -107
rect 177 -110 178 -109
rect 534 -110 535 -109
rect 548 -110 549 -109
rect 744 -110 745 -109
rect 807 -110 808 -109
rect 926 -110 927 -109
rect 933 -110 934 -109
rect 1199 -110 1200 -109
rect 184 -112 185 -111
rect 656 -112 657 -111
rect 744 -112 745 -111
rect 842 -112 843 -111
rect 947 -112 948 -111
rect 996 -112 997 -111
rect 1017 -112 1018 -111
rect 1059 -112 1060 -111
rect 1073 -112 1074 -111
rect 1220 -112 1221 -111
rect 198 -114 199 -113
rect 219 -114 220 -113
rect 229 -114 230 -113
rect 317 -114 318 -113
rect 373 -114 374 -113
rect 730 -114 731 -113
rect 814 -114 815 -113
rect 877 -114 878 -113
rect 912 -114 913 -113
rect 947 -114 948 -113
rect 1024 -114 1025 -113
rect 1059 -114 1060 -113
rect 1080 -114 1081 -113
rect 1178 -114 1179 -113
rect 198 -116 199 -115
rect 474 -116 475 -115
rect 492 -116 493 -115
rect 765 -116 766 -115
rect 891 -116 892 -115
rect 1080 -116 1081 -115
rect 1087 -116 1088 -115
rect 1206 -116 1207 -115
rect 205 -118 206 -117
rect 467 -118 468 -117
rect 534 -118 535 -117
rect 1076 -118 1077 -117
rect 1087 -118 1088 -117
rect 1248 -118 1249 -117
rect 212 -120 213 -119
rect 387 -120 388 -119
rect 390 -120 391 -119
rect 569 -120 570 -119
rect 597 -120 598 -119
rect 891 -120 892 -119
rect 1038 -120 1039 -119
rect 1111 -120 1112 -119
rect 261 -122 262 -121
rect 677 -122 678 -121
rect 681 -122 682 -121
rect 1024 -122 1025 -121
rect 1045 -122 1046 -121
rect 1129 -122 1130 -121
rect 275 -124 276 -123
rect 394 -124 395 -123
rect 401 -124 402 -123
rect 485 -124 486 -123
rect 646 -124 647 -123
rect 842 -124 843 -123
rect 1052 -124 1053 -123
rect 1066 -124 1067 -123
rect 296 -126 297 -125
rect 681 -126 682 -125
rect 688 -126 689 -125
rect 814 -126 815 -125
rect 142 -128 143 -127
rect 688 -128 689 -127
rect 723 -128 724 -127
rect 1052 -128 1053 -127
rect 394 -130 395 -129
rect 737 -130 738 -129
rect 408 -132 409 -131
rect 565 -132 566 -131
rect 723 -132 724 -131
rect 793 -132 794 -131
rect 121 -134 122 -133
rect 793 -134 794 -133
rect 415 -136 416 -135
rect 464 -136 465 -135
rect 485 -136 486 -135
rect 667 -136 668 -135
rect 446 -138 447 -137
rect 590 -138 591 -137
rect 667 -138 668 -137
rect 772 -138 773 -137
rect 457 -140 458 -139
rect 506 -140 507 -139
rect 565 -140 566 -139
rect 716 -140 717 -139
rect 772 -140 773 -139
rect 1045 -140 1046 -139
rect 460 -142 461 -141
rect 1227 -142 1228 -141
rect 16 -153 17 -152
rect 261 -153 262 -152
rect 282 -153 283 -152
rect 387 -153 388 -152
rect 408 -153 409 -152
rect 695 -153 696 -152
rect 768 -153 769 -152
rect 1346 -153 1347 -152
rect 1353 -153 1354 -152
rect 1367 -153 1368 -152
rect 1374 -153 1375 -152
rect 1500 -153 1501 -152
rect 1507 -153 1508 -152
rect 1626 -153 1627 -152
rect 1640 -153 1641 -152
rect 1668 -153 1669 -152
rect 1885 -153 1886 -152
rect 1941 -153 1942 -152
rect 23 -155 24 -154
rect 107 -155 108 -154
rect 114 -155 115 -154
rect 226 -155 227 -154
rect 240 -155 241 -154
rect 268 -155 269 -154
rect 282 -155 283 -154
rect 331 -155 332 -154
rect 345 -155 346 -154
rect 530 -155 531 -154
rect 541 -155 542 -154
rect 600 -155 601 -154
rect 611 -155 612 -154
rect 737 -155 738 -154
rect 803 -155 804 -154
rect 940 -155 941 -154
rect 950 -155 951 -154
rect 1402 -155 1403 -154
rect 1423 -155 1424 -154
rect 1493 -155 1494 -154
rect 1514 -155 1515 -154
rect 1556 -155 1557 -154
rect 1566 -155 1567 -154
rect 1584 -155 1585 -154
rect 1615 -155 1616 -154
rect 1633 -155 1634 -154
rect 37 -157 38 -156
rect 257 -157 258 -156
rect 331 -157 332 -156
rect 415 -157 416 -156
rect 422 -157 423 -156
rect 443 -157 444 -156
rect 450 -157 451 -156
rect 537 -157 538 -156
rect 541 -157 542 -156
rect 555 -157 556 -156
rect 590 -157 591 -156
rect 681 -157 682 -156
rect 684 -157 685 -156
rect 926 -157 927 -156
rect 1013 -157 1014 -156
rect 1430 -157 1431 -156
rect 1542 -157 1543 -156
rect 1815 -157 1816 -156
rect 44 -159 45 -158
rect 72 -159 73 -158
rect 86 -159 87 -158
rect 765 -159 766 -158
rect 814 -159 815 -158
rect 940 -159 941 -158
rect 1076 -159 1077 -158
rect 1248 -159 1249 -158
rect 1276 -159 1277 -158
rect 1570 -159 1571 -158
rect 51 -161 52 -160
rect 79 -161 80 -160
rect 93 -161 94 -160
rect 646 -161 647 -160
rect 649 -161 650 -160
rect 1080 -161 1081 -160
rect 1090 -161 1091 -160
rect 1465 -161 1466 -160
rect 72 -163 73 -162
rect 366 -163 367 -162
rect 380 -163 381 -162
rect 408 -163 409 -162
rect 429 -163 430 -162
rect 457 -163 458 -162
rect 467 -163 468 -162
rect 1024 -163 1025 -162
rect 1073 -163 1074 -162
rect 1248 -163 1249 -162
rect 1283 -163 1284 -162
rect 1577 -163 1578 -162
rect 79 -165 80 -164
rect 93 -165 94 -164
rect 100 -165 101 -164
rect 124 -165 125 -164
rect 128 -165 129 -164
rect 152 -165 153 -164
rect 163 -165 164 -164
rect 233 -165 234 -164
rect 240 -165 241 -164
rect 1507 -165 1508 -164
rect 100 -167 101 -166
rect 565 -167 566 -166
rect 618 -167 619 -166
rect 695 -167 696 -166
rect 737 -167 738 -166
rect 1010 -167 1011 -166
rect 1073 -167 1074 -166
rect 1108 -167 1109 -166
rect 1129 -167 1130 -166
rect 1451 -167 1452 -166
rect 107 -169 108 -168
rect 569 -169 570 -168
rect 621 -169 622 -168
rect 730 -169 731 -168
rect 814 -169 815 -168
rect 838 -169 839 -168
rect 849 -169 850 -168
rect 947 -169 948 -168
rect 975 -169 976 -168
rect 1276 -169 1277 -168
rect 1290 -169 1291 -168
rect 1374 -169 1375 -168
rect 117 -171 118 -170
rect 611 -171 612 -170
rect 849 -171 850 -170
rect 877 -171 878 -170
rect 884 -171 885 -170
rect 1108 -171 1109 -170
rect 1122 -171 1123 -170
rect 1290 -171 1291 -170
rect 1304 -171 1305 -170
rect 1444 -171 1445 -170
rect 121 -173 122 -172
rect 201 -173 202 -172
rect 226 -173 227 -172
rect 772 -173 773 -172
rect 856 -173 857 -172
rect 877 -173 878 -172
rect 887 -173 888 -172
rect 1227 -173 1228 -172
rect 1311 -173 1312 -172
rect 1472 -173 1473 -172
rect 128 -175 129 -174
rect 254 -175 255 -174
rect 275 -175 276 -174
rect 429 -175 430 -174
rect 450 -175 451 -174
rect 478 -175 479 -174
rect 492 -175 493 -174
rect 597 -175 598 -174
rect 667 -175 668 -174
rect 772 -175 773 -174
rect 870 -175 871 -174
rect 1024 -175 1025 -174
rect 1059 -175 1060 -174
rect 1129 -175 1130 -174
rect 1136 -175 1137 -174
rect 1395 -175 1396 -174
rect 65 -177 66 -176
rect 254 -177 255 -176
rect 275 -177 276 -176
rect 359 -177 360 -176
rect 366 -177 367 -176
rect 894 -177 895 -176
rect 905 -177 906 -176
rect 975 -177 976 -176
rect 989 -177 990 -176
rect 1136 -177 1137 -176
rect 1150 -177 1151 -176
rect 1283 -177 1284 -176
rect 1318 -177 1319 -176
rect 1437 -177 1438 -176
rect 135 -179 136 -178
rect 261 -179 262 -178
rect 338 -179 339 -178
rect 478 -179 479 -178
rect 513 -179 514 -178
rect 562 -179 563 -178
rect 569 -179 570 -178
rect 929 -179 930 -178
rect 961 -179 962 -178
rect 1304 -179 1305 -178
rect 1325 -179 1326 -178
rect 1591 -179 1592 -178
rect 142 -181 143 -180
rect 212 -181 213 -180
rect 243 -181 244 -180
rect 271 -181 272 -180
rect 296 -181 297 -180
rect 338 -181 339 -180
rect 345 -181 346 -180
rect 485 -181 486 -180
rect 513 -181 514 -180
rect 593 -181 594 -180
rect 705 -181 706 -180
rect 1227 -181 1228 -180
rect 1325 -181 1326 -180
rect 1332 -181 1333 -180
rect 1360 -181 1361 -180
rect 1458 -181 1459 -180
rect 145 -183 146 -182
rect 156 -183 157 -182
rect 163 -183 164 -182
rect 390 -183 391 -182
rect 401 -183 402 -182
rect 415 -183 416 -182
rect 471 -183 472 -182
rect 1010 -183 1011 -182
rect 1017 -183 1018 -182
rect 1122 -183 1123 -182
rect 1164 -183 1165 -182
rect 1423 -183 1424 -182
rect 149 -185 150 -184
rect 716 -185 717 -184
rect 786 -185 787 -184
rect 905 -185 906 -184
rect 919 -185 920 -184
rect 1059 -185 1060 -184
rect 1080 -185 1081 -184
rect 1115 -185 1116 -184
rect 1171 -185 1172 -184
rect 1388 -185 1389 -184
rect 156 -187 157 -186
rect 1514 -187 1515 -186
rect 170 -189 171 -188
rect 492 -189 493 -188
rect 520 -189 521 -188
rect 989 -189 990 -188
rect 1003 -189 1004 -188
rect 1360 -189 1361 -188
rect 177 -191 178 -190
rect 359 -191 360 -190
rect 373 -191 374 -190
rect 667 -191 668 -190
rect 709 -191 710 -190
rect 856 -191 857 -190
rect 912 -191 913 -190
rect 919 -191 920 -190
rect 954 -191 955 -190
rect 1164 -191 1165 -190
rect 1171 -191 1172 -190
rect 1265 -191 1266 -190
rect 177 -193 178 -192
rect 436 -193 437 -192
rect 520 -193 521 -192
rect 947 -193 948 -192
rect 968 -193 969 -192
rect 1115 -193 1116 -192
rect 1174 -193 1175 -192
rect 1241 -193 1242 -192
rect 58 -195 59 -194
rect 436 -195 437 -194
rect 527 -195 528 -194
rect 1052 -195 1053 -194
rect 1094 -195 1095 -194
rect 1521 -195 1522 -194
rect 58 -197 59 -196
rect 159 -197 160 -196
rect 184 -197 185 -196
rect 296 -197 297 -196
rect 310 -197 311 -196
rect 485 -197 486 -196
rect 506 -197 507 -196
rect 527 -197 528 -196
rect 534 -197 535 -196
rect 716 -197 717 -196
rect 758 -197 759 -196
rect 786 -197 787 -196
rect 793 -197 794 -196
rect 961 -197 962 -196
rect 1017 -197 1018 -196
rect 1150 -197 1151 -196
rect 1178 -197 1179 -196
rect 1353 -197 1354 -196
rect 170 -199 171 -198
rect 310 -199 311 -198
rect 317 -199 318 -198
rect 373 -199 374 -198
rect 394 -199 395 -198
rect 506 -199 507 -198
rect 555 -199 556 -198
rect 779 -199 780 -198
rect 821 -199 822 -198
rect 870 -199 871 -198
rect 1038 -199 1039 -198
rect 1052 -199 1053 -198
rect 1094 -199 1095 -198
rect 1143 -199 1144 -198
rect 1185 -199 1186 -198
rect 1409 -199 1410 -198
rect 184 -201 185 -200
rect 460 -201 461 -200
rect 674 -201 675 -200
rect 968 -201 969 -200
rect 1038 -201 1039 -200
rect 1549 -201 1550 -200
rect 194 -203 195 -202
rect 933 -203 934 -202
rect 1101 -203 1102 -202
rect 1416 -203 1417 -202
rect 198 -205 199 -204
rect 422 -205 423 -204
rect 660 -205 661 -204
rect 674 -205 675 -204
rect 688 -205 689 -204
rect 954 -205 955 -204
rect 1066 -205 1067 -204
rect 1101 -205 1102 -204
rect 1143 -205 1144 -204
rect 1269 -205 1270 -204
rect 30 -207 31 -206
rect 198 -207 199 -206
rect 212 -207 213 -206
rect 821 -207 822 -206
rect 898 -207 899 -206
rect 1185 -207 1186 -206
rect 1192 -207 1193 -206
rect 1528 -207 1529 -206
rect 219 -209 220 -208
rect 317 -209 318 -208
rect 324 -209 325 -208
rect 394 -209 395 -208
rect 401 -209 402 -208
rect 639 -209 640 -208
rect 698 -209 699 -208
rect 1192 -209 1193 -208
rect 1199 -209 1200 -208
rect 1486 -209 1487 -208
rect 219 -211 220 -210
rect 499 -211 500 -210
rect 548 -211 549 -210
rect 660 -211 661 -210
rect 709 -211 710 -210
rect 1234 -211 1235 -210
rect 1241 -211 1242 -210
rect 1297 -211 1298 -210
rect 247 -213 248 -212
rect 999 -213 1000 -212
rect 1031 -213 1032 -212
rect 1066 -213 1067 -212
rect 1157 -213 1158 -212
rect 1234 -213 1235 -212
rect 1255 -213 1256 -212
rect 1297 -213 1298 -212
rect 89 -215 90 -214
rect 247 -215 248 -214
rect 324 -215 325 -214
rect 1262 -215 1263 -214
rect 1269 -215 1270 -214
rect 1612 -215 1613 -214
rect 352 -217 353 -216
rect 380 -217 381 -216
rect 499 -217 500 -216
rect 751 -217 752 -216
rect 758 -217 759 -216
rect 1087 -217 1088 -216
rect 1199 -217 1200 -216
rect 1381 -217 1382 -216
rect 352 -219 353 -218
rect 523 -219 524 -218
rect 548 -219 549 -218
rect 915 -219 916 -218
rect 996 -219 997 -218
rect 1087 -219 1088 -218
rect 1202 -219 1203 -218
rect 1339 -219 1340 -218
rect 523 -221 524 -220
rect 842 -221 843 -220
rect 863 -221 864 -220
rect 1031 -221 1032 -220
rect 1045 -221 1046 -220
rect 1157 -221 1158 -220
rect 1206 -221 1207 -220
rect 1479 -221 1480 -220
rect 583 -223 584 -222
rect 751 -223 752 -222
rect 765 -223 766 -222
rect 1178 -223 1179 -222
rect 1213 -223 1214 -222
rect 1311 -223 1312 -222
rect 576 -225 577 -224
rect 583 -225 584 -224
rect 604 -225 605 -224
rect 688 -225 689 -224
rect 702 -225 703 -224
rect 863 -225 864 -224
rect 891 -225 892 -224
rect 1262 -225 1263 -224
rect 303 -227 304 -226
rect 604 -227 605 -226
rect 632 -227 633 -226
rect 842 -227 843 -226
rect 982 -227 983 -226
rect 1045 -227 1046 -226
rect 1216 -227 1217 -226
rect 1318 -227 1319 -226
rect 205 -229 206 -228
rect 303 -229 304 -228
rect 576 -229 577 -228
rect 733 -229 734 -228
rect 744 -229 745 -228
rect 793 -229 794 -228
rect 807 -229 808 -228
rect 898 -229 899 -228
rect 936 -229 937 -228
rect 982 -229 983 -228
rect 1003 -229 1004 -228
rect 1213 -229 1214 -228
rect 1220 -229 1221 -228
rect 1535 -229 1536 -228
rect 439 -231 440 -230
rect 1220 -231 1221 -230
rect 1255 -231 1256 -230
rect 1328 -231 1329 -230
rect 625 -233 626 -232
rect 632 -233 633 -232
rect 639 -233 640 -232
rect 712 -233 713 -232
rect 779 -233 780 -232
rect 1146 -233 1147 -232
rect 191 -235 192 -234
rect 625 -235 626 -234
rect 653 -235 654 -234
rect 744 -235 745 -234
rect 807 -235 808 -234
rect 884 -235 885 -234
rect 135 -237 136 -236
rect 653 -237 654 -236
rect 835 -237 836 -236
rect 1206 -237 1207 -236
rect 800 -239 801 -238
rect 835 -239 836 -238
rect 800 -241 801 -240
rect 828 -241 829 -240
rect 723 -243 724 -242
rect 828 -243 829 -242
rect 534 -245 535 -244
rect 723 -245 724 -244
rect 16 -256 17 -255
rect 194 -256 195 -255
rect 198 -256 199 -255
rect 338 -256 339 -255
rect 366 -256 367 -255
rect 747 -256 748 -255
rect 761 -256 762 -255
rect 915 -256 916 -255
rect 992 -256 993 -255
rect 1598 -256 1599 -255
rect 1612 -256 1613 -255
rect 1969 -256 1970 -255
rect 16 -258 17 -257
rect 149 -258 150 -257
rect 156 -258 157 -257
rect 537 -258 538 -257
rect 618 -258 619 -257
rect 800 -258 801 -257
rect 810 -258 811 -257
rect 1801 -258 1802 -257
rect 1815 -258 1816 -257
rect 1927 -258 1928 -257
rect 1941 -258 1942 -257
rect 1983 -258 1984 -257
rect 44 -260 45 -259
rect 208 -260 209 -259
rect 240 -260 241 -259
rect 313 -260 314 -259
rect 338 -260 339 -259
rect 408 -260 409 -259
rect 432 -260 433 -259
rect 796 -260 797 -259
rect 828 -260 829 -259
rect 845 -260 846 -259
rect 880 -260 881 -259
rect 1528 -260 1529 -259
rect 1542 -260 1543 -259
rect 1605 -260 1606 -259
rect 1615 -260 1616 -259
rect 1661 -260 1662 -259
rect 1668 -260 1669 -259
rect 1731 -260 1732 -259
rect 1962 -260 1963 -259
rect 2193 -260 2194 -259
rect 23 -262 24 -261
rect 240 -262 241 -261
rect 247 -262 248 -261
rect 436 -262 437 -261
rect 439 -262 440 -261
rect 590 -262 591 -261
rect 653 -262 654 -261
rect 884 -262 885 -261
rect 891 -262 892 -261
rect 1640 -262 1641 -261
rect 23 -264 24 -263
rect 37 -264 38 -263
rect 54 -264 55 -263
rect 1507 -264 1508 -263
rect 1514 -264 1515 -263
rect 1843 -264 1844 -263
rect 37 -266 38 -265
rect 415 -266 416 -265
rect 422 -266 423 -265
rect 590 -266 591 -265
rect 709 -266 710 -265
rect 1031 -266 1032 -265
rect 1083 -266 1084 -265
rect 1689 -266 1690 -265
rect 65 -268 66 -267
rect 128 -268 129 -267
rect 149 -268 150 -267
rect 170 -268 171 -267
rect 187 -268 188 -267
rect 254 -268 255 -267
rect 268 -268 269 -267
rect 303 -268 304 -267
rect 310 -268 311 -267
rect 982 -268 983 -267
rect 996 -268 997 -267
rect 1829 -268 1830 -267
rect 86 -270 87 -269
rect 93 -270 94 -269
rect 114 -270 115 -269
rect 142 -270 143 -269
rect 156 -270 157 -269
rect 632 -270 633 -269
rect 709 -270 710 -269
rect 814 -270 815 -269
rect 828 -270 829 -269
rect 849 -270 850 -269
rect 856 -270 857 -269
rect 996 -270 997 -269
rect 1010 -270 1011 -269
rect 1780 -270 1781 -269
rect 58 -272 59 -271
rect 142 -272 143 -271
rect 233 -272 234 -271
rect 408 -272 409 -271
rect 422 -272 423 -271
rect 457 -272 458 -271
rect 506 -272 507 -271
rect 520 -272 521 -271
rect 534 -272 535 -271
rect 940 -272 941 -271
rect 954 -272 955 -271
rect 1031 -272 1032 -271
rect 1094 -272 1095 -271
rect 1549 -272 1550 -271
rect 1552 -272 1553 -271
rect 1766 -272 1767 -271
rect 58 -274 59 -273
rect 744 -274 745 -273
rect 772 -274 773 -273
rect 814 -274 815 -273
rect 856 -274 857 -273
rect 989 -274 990 -273
rect 1010 -274 1011 -273
rect 1017 -274 1018 -273
rect 1020 -274 1021 -273
rect 1451 -274 1452 -273
rect 1465 -274 1466 -273
rect 1794 -274 1795 -273
rect 93 -276 94 -275
rect 100 -276 101 -275
rect 128 -276 129 -275
rect 261 -276 262 -275
rect 268 -276 269 -275
rect 471 -276 472 -275
rect 506 -276 507 -275
rect 779 -276 780 -275
rect 863 -276 864 -275
rect 940 -276 941 -275
rect 954 -276 955 -275
rect 1003 -276 1004 -275
rect 1101 -276 1102 -275
rect 1199 -276 1200 -275
rect 1227 -276 1228 -275
rect 1647 -276 1648 -275
rect 100 -278 101 -277
rect 177 -278 178 -277
rect 205 -278 206 -277
rect 779 -278 780 -277
rect 842 -278 843 -277
rect 863 -278 864 -277
rect 894 -278 895 -277
rect 1535 -278 1536 -277
rect 1556 -278 1557 -277
rect 1654 -278 1655 -277
rect 72 -280 73 -279
rect 177 -280 178 -279
rect 191 -280 192 -279
rect 205 -280 206 -279
rect 219 -280 220 -279
rect 534 -280 535 -279
rect 555 -280 556 -279
rect 618 -280 619 -279
rect 628 -280 629 -279
rect 1003 -280 1004 -279
rect 1153 -280 1154 -279
rect 1710 -280 1711 -279
rect 72 -282 73 -281
rect 835 -282 836 -281
rect 926 -282 927 -281
rect 1094 -282 1095 -281
rect 1178 -282 1179 -281
rect 1514 -282 1515 -281
rect 1591 -282 1592 -281
rect 1815 -282 1816 -281
rect 107 -284 108 -283
rect 261 -284 262 -283
rect 275 -284 276 -283
rect 464 -284 465 -283
rect 471 -284 472 -283
rect 485 -284 486 -283
rect 513 -284 514 -283
rect 653 -284 654 -283
rect 667 -284 668 -283
rect 849 -284 850 -283
rect 947 -284 948 -283
rect 1227 -284 1228 -283
rect 1262 -284 1263 -283
rect 1752 -284 1753 -283
rect 107 -286 108 -285
rect 212 -286 213 -285
rect 219 -286 220 -285
rect 226 -286 227 -285
rect 233 -286 234 -285
rect 894 -286 895 -285
rect 947 -286 948 -285
rect 1545 -286 1546 -285
rect 1626 -286 1627 -285
rect 1717 -286 1718 -285
rect 135 -288 136 -287
rect 303 -288 304 -287
rect 310 -288 311 -287
rect 450 -288 451 -287
rect 548 -288 549 -287
rect 555 -288 556 -287
rect 569 -288 570 -287
rect 926 -288 927 -287
rect 968 -288 969 -287
rect 982 -288 983 -287
rect 1213 -288 1214 -287
rect 1535 -288 1536 -287
rect 1633 -288 1634 -287
rect 1745 -288 1746 -287
rect 30 -290 31 -289
rect 450 -290 451 -289
rect 548 -290 549 -289
rect 912 -290 913 -289
rect 1122 -290 1123 -289
rect 1213 -290 1214 -289
rect 1276 -290 1277 -289
rect 1507 -290 1508 -289
rect 30 -292 31 -291
rect 51 -292 52 -291
rect 138 -292 139 -291
rect 170 -292 171 -291
rect 226 -292 227 -291
rect 352 -292 353 -291
rect 394 -292 395 -291
rect 457 -292 458 -291
rect 611 -292 612 -291
rect 968 -292 969 -291
rect 975 -292 976 -291
rect 1122 -292 1123 -291
rect 1136 -292 1137 -291
rect 1276 -292 1277 -291
rect 1297 -292 1298 -291
rect 1528 -292 1529 -291
rect 47 -294 48 -293
rect 51 -294 52 -293
rect 138 -294 139 -293
rect 366 -294 367 -293
rect 394 -294 395 -293
rect 481 -294 482 -293
rect 611 -294 612 -293
rect 681 -294 682 -293
rect 702 -294 703 -293
rect 1262 -294 1263 -293
rect 1318 -294 1319 -293
rect 1556 -294 1557 -293
rect 89 -296 90 -295
rect 681 -296 682 -295
rect 688 -296 689 -295
rect 702 -296 703 -295
rect 723 -296 724 -295
rect 912 -296 913 -295
rect 919 -296 920 -295
rect 1318 -296 1319 -295
rect 1328 -296 1329 -295
rect 2004 -296 2005 -295
rect 243 -298 244 -297
rect 415 -298 416 -297
rect 429 -298 430 -297
rect 464 -298 465 -297
rect 576 -298 577 -297
rect 919 -298 920 -297
rect 1108 -298 1109 -297
rect 1297 -298 1298 -297
rect 1353 -298 1354 -297
rect 1626 -298 1627 -297
rect 247 -300 248 -299
rect 404 -300 405 -299
rect 576 -300 577 -299
rect 838 -300 839 -299
rect 1024 -300 1025 -299
rect 1108 -300 1109 -299
rect 1360 -300 1361 -299
rect 1738 -300 1739 -299
rect 254 -302 255 -301
rect 271 -302 272 -301
rect 275 -302 276 -301
rect 324 -302 325 -301
rect 345 -302 346 -301
rect 569 -302 570 -301
rect 597 -302 598 -301
rect 688 -302 689 -301
rect 723 -302 724 -301
rect 758 -302 759 -301
rect 772 -302 773 -301
rect 1591 -302 1592 -301
rect 282 -304 283 -303
rect 436 -304 437 -303
rect 660 -304 661 -303
rect 667 -304 668 -303
rect 730 -304 731 -303
rect 842 -304 843 -303
rect 1171 -304 1172 -303
rect 1360 -304 1361 -303
rect 1374 -304 1375 -303
rect 1822 -304 1823 -303
rect 135 -306 136 -305
rect 282 -306 283 -305
rect 289 -306 290 -305
rect 485 -306 486 -305
rect 660 -306 661 -305
rect 1325 -306 1326 -305
rect 1381 -306 1382 -305
rect 1465 -306 1466 -305
rect 1472 -306 1473 -305
rect 1787 -306 1788 -305
rect 289 -308 290 -307
rect 387 -308 388 -307
rect 401 -308 402 -307
rect 513 -308 514 -307
rect 716 -308 717 -307
rect 730 -308 731 -307
rect 786 -308 787 -307
rect 1136 -308 1137 -307
rect 1185 -308 1186 -307
rect 1374 -308 1375 -307
rect 1388 -308 1389 -307
rect 1619 -308 1620 -307
rect 296 -310 297 -309
rect 499 -310 500 -309
rect 646 -310 647 -309
rect 716 -310 717 -309
rect 786 -310 787 -309
rect 1027 -310 1028 -309
rect 1073 -310 1074 -309
rect 1171 -310 1172 -309
rect 1185 -310 1186 -309
rect 1332 -310 1333 -309
rect 1395 -310 1396 -309
rect 1682 -310 1683 -309
rect 212 -312 213 -311
rect 646 -312 647 -311
rect 1073 -312 1074 -311
rect 1269 -312 1270 -311
rect 1402 -312 1403 -311
rect 1668 -312 1669 -311
rect 299 -314 300 -313
rect 807 -314 808 -313
rect 1076 -314 1077 -313
rect 1395 -314 1396 -313
rect 1409 -314 1410 -313
rect 1675 -314 1676 -313
rect 324 -316 325 -315
rect 541 -316 542 -315
rect 1157 -316 1158 -315
rect 1269 -316 1270 -315
rect 1311 -316 1312 -315
rect 1402 -316 1403 -315
rect 1416 -316 1417 -315
rect 1696 -316 1697 -315
rect 331 -318 332 -317
rect 499 -318 500 -317
rect 933 -318 934 -317
rect 1416 -318 1417 -317
rect 1423 -318 1424 -317
rect 1759 -318 1760 -317
rect 331 -320 332 -319
rect 800 -320 801 -319
rect 870 -320 871 -319
rect 933 -320 934 -319
rect 1104 -320 1105 -319
rect 1311 -320 1312 -319
rect 1430 -320 1431 -319
rect 1724 -320 1725 -319
rect 345 -322 346 -321
rect 527 -322 528 -321
rect 632 -322 633 -321
rect 870 -322 871 -321
rect 1157 -322 1158 -321
rect 1255 -322 1256 -321
rect 1437 -322 1438 -321
rect 1703 -322 1704 -321
rect 79 -324 80 -323
rect 527 -324 528 -323
rect 712 -324 713 -323
rect 1255 -324 1256 -323
rect 1444 -324 1445 -323
rect 1773 -324 1774 -323
rect 79 -326 80 -325
rect 163 -326 164 -325
rect 352 -326 353 -325
rect 621 -326 622 -325
rect 1164 -326 1165 -325
rect 1332 -326 1333 -325
rect 1451 -326 1452 -325
rect 1612 -326 1613 -325
rect 163 -328 164 -327
rect 166 -328 167 -327
rect 359 -328 360 -327
rect 597 -328 598 -327
rect 1017 -328 1018 -327
rect 1164 -328 1165 -327
rect 1192 -328 1193 -327
rect 1388 -328 1389 -327
rect 1472 -328 1473 -327
rect 1584 -328 1585 -327
rect 359 -330 360 -329
rect 523 -330 524 -329
rect 1066 -330 1067 -329
rect 1192 -330 1193 -329
rect 1206 -330 1207 -329
rect 1423 -330 1424 -329
rect 1486 -330 1487 -329
rect 1836 -330 1837 -329
rect 117 -332 118 -331
rect 1066 -332 1067 -331
rect 1087 -332 1088 -331
rect 1206 -332 1207 -331
rect 1220 -332 1221 -331
rect 1430 -332 1431 -331
rect 1493 -332 1494 -331
rect 1633 -332 1634 -331
rect 380 -334 381 -333
rect 387 -334 388 -333
rect 443 -334 444 -333
rect 541 -334 542 -333
rect 961 -334 962 -333
rect 1087 -334 1088 -333
rect 1234 -334 1235 -333
rect 1409 -334 1410 -333
rect 1500 -334 1501 -333
rect 1808 -334 1809 -333
rect 373 -336 374 -335
rect 380 -336 381 -335
rect 443 -336 444 -335
rect 478 -336 479 -335
rect 765 -336 766 -335
rect 961 -336 962 -335
rect 1038 -336 1039 -335
rect 1220 -336 1221 -335
rect 1248 -336 1249 -335
rect 1437 -336 1438 -335
rect 1479 -336 1480 -335
rect 1500 -336 1501 -335
rect 1563 -336 1564 -335
rect 1584 -336 1585 -335
rect 373 -338 374 -337
rect 705 -338 706 -337
rect 1038 -338 1039 -337
rect 1150 -338 1151 -337
rect 1248 -338 1249 -337
rect 1577 -338 1578 -337
rect 478 -340 479 -339
rect 1542 -340 1543 -339
rect 639 -342 640 -341
rect 765 -342 766 -341
rect 1129 -342 1130 -341
rect 1234 -342 1235 -341
rect 1283 -342 1284 -341
rect 1493 -342 1494 -341
rect 639 -344 640 -343
rect 695 -344 696 -343
rect 1045 -344 1046 -343
rect 1283 -344 1284 -343
rect 1290 -344 1291 -343
rect 1444 -344 1445 -343
rect 695 -346 696 -345
rect 737 -346 738 -345
rect 877 -346 878 -345
rect 1045 -346 1046 -345
rect 1052 -346 1053 -345
rect 1129 -346 1130 -345
rect 1150 -346 1151 -345
rect 1570 -346 1571 -345
rect 604 -348 605 -347
rect 737 -348 738 -347
rect 877 -348 878 -347
rect 1381 -348 1382 -347
rect 1458 -348 1459 -347
rect 1570 -348 1571 -347
rect 317 -350 318 -349
rect 604 -350 605 -349
rect 625 -350 626 -349
rect 1458 -350 1459 -349
rect 121 -352 122 -351
rect 317 -352 318 -351
rect 401 -352 402 -351
rect 625 -352 626 -351
rect 898 -352 899 -351
rect 1052 -352 1053 -351
rect 1304 -352 1305 -351
rect 1479 -352 1480 -351
rect 121 -354 122 -353
rect 583 -354 584 -353
rect 898 -354 899 -353
rect 1143 -354 1144 -353
rect 1339 -354 1340 -353
rect 1563 -354 1564 -353
rect 492 -356 493 -355
rect 583 -356 584 -355
rect 1024 -356 1025 -355
rect 1290 -356 1291 -355
rect 1346 -356 1347 -355
rect 1577 -356 1578 -355
rect 492 -358 493 -357
rect 562 -358 563 -357
rect 821 -358 822 -357
rect 1346 -358 1347 -357
rect 1367 -358 1368 -357
rect 1486 -358 1487 -357
rect 184 -360 185 -359
rect 562 -360 563 -359
rect 751 -360 752 -359
rect 821 -360 822 -359
rect 1059 -360 1060 -359
rect 1143 -360 1144 -359
rect 1181 -360 1182 -359
rect 1367 -360 1368 -359
rect 674 -362 675 -361
rect 751 -362 752 -361
rect 905 -362 906 -361
rect 1059 -362 1060 -361
rect 1115 -362 1116 -361
rect 1304 -362 1305 -361
rect 467 -364 468 -363
rect 674 -364 675 -363
rect 793 -364 794 -363
rect 905 -364 906 -363
rect 1080 -364 1081 -363
rect 1115 -364 1116 -363
rect 1241 -364 1242 -363
rect 1339 -364 1340 -363
rect 793 -366 794 -365
rect 1521 -366 1522 -365
rect 835 -368 836 -367
rect 1521 -368 1522 -367
rect 887 -370 888 -369
rect 1241 -370 1242 -369
rect 16 -381 17 -380
rect 621 -381 622 -380
rect 625 -381 626 -380
rect 702 -381 703 -380
rect 758 -381 759 -380
rect 1297 -381 1298 -380
rect 1353 -381 1354 -380
rect 1948 -381 1949 -380
rect 1958 -381 1959 -380
rect 2116 -381 2117 -380
rect 2193 -381 2194 -380
rect 2284 -381 2285 -380
rect 23 -383 24 -382
rect 747 -383 748 -382
rect 751 -383 752 -382
rect 758 -383 759 -382
rect 761 -383 762 -382
rect 800 -383 801 -382
rect 810 -383 811 -382
rect 828 -383 829 -382
rect 845 -383 846 -382
rect 1752 -383 1753 -382
rect 1766 -383 1767 -382
rect 1962 -383 1963 -382
rect 1969 -383 1970 -382
rect 2088 -383 2089 -382
rect 23 -385 24 -384
rect 44 -385 45 -384
rect 51 -385 52 -384
rect 79 -385 80 -384
rect 96 -385 97 -384
rect 1178 -385 1179 -384
rect 1185 -385 1186 -384
rect 1297 -385 1298 -384
rect 1353 -385 1354 -384
rect 1472 -385 1473 -384
rect 1591 -385 1592 -384
rect 1752 -385 1753 -384
rect 1773 -385 1774 -384
rect 1899 -385 1900 -384
rect 1927 -385 1928 -384
rect 1997 -385 1998 -384
rect 2004 -385 2005 -384
rect 2263 -385 2264 -384
rect 37 -387 38 -386
rect 481 -387 482 -386
rect 495 -387 496 -386
rect 562 -387 563 -386
rect 600 -387 601 -386
rect 1136 -387 1137 -386
rect 1167 -387 1168 -386
rect 1682 -387 1683 -386
rect 1710 -387 1711 -386
rect 1850 -387 1851 -386
rect 1976 -387 1977 -386
rect 1990 -387 1991 -386
rect 2011 -387 2012 -386
rect 2144 -387 2145 -386
rect 44 -389 45 -388
rect 446 -389 447 -388
rect 478 -389 479 -388
rect 856 -389 857 -388
rect 971 -389 972 -388
rect 1759 -389 1760 -388
rect 1794 -389 1795 -388
rect 1906 -389 1907 -388
rect 1983 -389 1984 -388
rect 2039 -389 2040 -388
rect 61 -391 62 -390
rect 247 -391 248 -390
rect 345 -391 346 -390
rect 478 -391 479 -390
rect 513 -391 514 -390
rect 562 -391 563 -390
rect 625 -391 626 -390
rect 884 -391 885 -390
rect 978 -391 979 -390
rect 1346 -391 1347 -390
rect 1356 -391 1357 -390
rect 1430 -391 1431 -390
rect 1440 -391 1441 -390
rect 1983 -391 1984 -390
rect 72 -393 73 -392
rect 135 -393 136 -392
rect 163 -393 164 -392
rect 1801 -393 1802 -392
rect 1808 -393 1809 -392
rect 1913 -393 1914 -392
rect 16 -395 17 -394
rect 163 -395 164 -394
rect 170 -395 171 -394
rect 215 -395 216 -394
rect 222 -395 223 -394
rect 590 -395 591 -394
rect 635 -395 636 -394
rect 1591 -395 1592 -394
rect 1612 -395 1613 -394
rect 1941 -395 1942 -394
rect 72 -397 73 -396
rect 86 -397 87 -396
rect 173 -397 174 -396
rect 205 -397 206 -396
rect 233 -397 234 -396
rect 751 -397 752 -396
rect 765 -397 766 -396
rect 891 -397 892 -396
rect 978 -397 979 -396
rect 1087 -397 1088 -396
rect 1125 -397 1126 -396
rect 1857 -397 1858 -396
rect 30 -399 31 -398
rect 233 -399 234 -398
rect 247 -399 248 -398
rect 373 -399 374 -398
rect 401 -399 402 -398
rect 506 -399 507 -398
rect 513 -399 514 -398
rect 688 -399 689 -398
rect 702 -399 703 -398
rect 1006 -399 1007 -398
rect 1017 -399 1018 -398
rect 1780 -399 1781 -398
rect 1815 -399 1816 -398
rect 1920 -399 1921 -398
rect 79 -401 80 -400
rect 611 -401 612 -400
rect 646 -401 647 -400
rect 912 -401 913 -400
rect 982 -401 983 -400
rect 1104 -401 1105 -400
rect 1136 -401 1137 -400
rect 1248 -401 1249 -400
rect 1262 -401 1263 -400
rect 1346 -401 1347 -400
rect 1360 -401 1361 -400
rect 1430 -401 1431 -400
rect 1493 -401 1494 -400
rect 1612 -401 1613 -400
rect 1633 -401 1634 -400
rect 1759 -401 1760 -400
rect 1787 -401 1788 -400
rect 1815 -401 1816 -400
rect 1836 -401 1837 -400
rect 1934 -401 1935 -400
rect 86 -403 87 -402
rect 415 -403 416 -402
rect 443 -403 444 -402
rect 506 -403 507 -402
rect 527 -403 528 -402
rect 982 -403 983 -402
rect 1020 -403 1021 -402
rect 1325 -403 1326 -402
rect 1360 -403 1361 -402
rect 1542 -403 1543 -402
rect 1549 -403 1550 -402
rect 1633 -403 1634 -402
rect 1654 -403 1655 -402
rect 1864 -403 1865 -402
rect 121 -405 122 -404
rect 205 -405 206 -404
rect 212 -405 213 -404
rect 443 -405 444 -404
rect 527 -405 528 -404
rect 548 -405 549 -404
rect 667 -405 668 -404
rect 772 -405 773 -404
rect 793 -405 794 -404
rect 1738 -405 1739 -404
rect 1745 -405 1746 -404
rect 1892 -405 1893 -404
rect 114 -407 115 -406
rect 121 -407 122 -406
rect 156 -407 157 -406
rect 765 -407 766 -406
rect 849 -407 850 -406
rect 891 -407 892 -406
rect 1024 -407 1025 -406
rect 1773 -407 1774 -406
rect 1843 -407 1844 -406
rect 1969 -407 1970 -406
rect 156 -409 157 -408
rect 191 -409 192 -408
rect 219 -409 220 -408
rect 667 -409 668 -408
rect 674 -409 675 -408
rect 828 -409 829 -408
rect 852 -409 853 -408
rect 1122 -409 1123 -408
rect 1129 -409 1130 -408
rect 1248 -409 1249 -408
rect 1388 -409 1389 -408
rect 1472 -409 1473 -408
rect 1500 -409 1501 -408
rect 1843 -409 1844 -408
rect 149 -411 150 -410
rect 191 -411 192 -410
rect 226 -411 227 -410
rect 611 -411 612 -410
rect 674 -411 675 -410
rect 709 -411 710 -410
rect 716 -411 717 -410
rect 772 -411 773 -410
rect 856 -411 857 -410
rect 985 -411 986 -410
rect 1027 -411 1028 -410
rect 1962 -411 1963 -410
rect 149 -413 150 -412
rect 432 -413 433 -412
rect 541 -413 542 -412
rect 590 -413 591 -412
rect 653 -413 654 -412
rect 709 -413 710 -412
rect 730 -413 731 -412
rect 793 -413 794 -412
rect 863 -413 864 -412
rect 912 -413 913 -412
rect 1031 -413 1032 -412
rect 1087 -413 1088 -412
rect 1164 -413 1165 -412
rect 1542 -413 1543 -412
rect 1563 -413 1564 -412
rect 1654 -413 1655 -412
rect 1661 -413 1662 -412
rect 1780 -413 1781 -412
rect 187 -415 188 -414
rect 1766 -415 1767 -414
rect 226 -417 227 -416
rect 240 -417 241 -416
rect 345 -417 346 -416
rect 464 -417 465 -416
rect 541 -417 542 -416
rect 649 -417 650 -416
rect 653 -417 654 -416
rect 1479 -417 1480 -416
rect 1507 -417 1508 -416
rect 1549 -417 1550 -416
rect 1570 -417 1571 -416
rect 1801 -417 1802 -416
rect 240 -419 241 -418
rect 268 -419 269 -418
rect 359 -419 360 -418
rect 429 -419 430 -418
rect 548 -419 549 -418
rect 569 -419 570 -418
rect 681 -419 682 -418
rect 1017 -419 1018 -418
rect 1059 -419 1060 -418
rect 1129 -419 1130 -418
rect 1178 -419 1179 -418
rect 1290 -419 1291 -418
rect 1311 -419 1312 -418
rect 1388 -419 1389 -418
rect 1402 -419 1403 -418
rect 1493 -419 1494 -418
rect 1584 -419 1585 -418
rect 1710 -419 1711 -418
rect 1724 -419 1725 -418
rect 1878 -419 1879 -418
rect 166 -421 167 -420
rect 359 -421 360 -420
rect 373 -421 374 -420
rect 436 -421 437 -420
rect 471 -421 472 -420
rect 681 -421 682 -420
rect 688 -421 689 -420
rect 957 -421 958 -420
rect 968 -421 969 -420
rect 1031 -421 1032 -420
rect 1073 -421 1074 -420
rect 1871 -421 1872 -420
rect 100 -423 101 -422
rect 436 -423 437 -422
rect 457 -423 458 -422
rect 471 -423 472 -422
rect 730 -423 731 -422
rect 807 -423 808 -422
rect 1076 -423 1077 -422
rect 1647 -423 1648 -422
rect 1668 -423 1669 -422
rect 1787 -423 1788 -422
rect 100 -425 101 -424
rect 520 -425 521 -424
rect 744 -425 745 -424
rect 1262 -425 1263 -424
rect 1328 -425 1329 -424
rect 1668 -425 1669 -424
rect 1675 -425 1676 -424
rect 1794 -425 1795 -424
rect 166 -427 167 -426
rect 331 -427 332 -426
rect 401 -427 402 -426
rect 485 -427 486 -426
rect 737 -427 738 -426
rect 744 -427 745 -426
rect 779 -427 780 -426
rect 1073 -427 1074 -426
rect 1080 -427 1081 -426
rect 1227 -427 1228 -426
rect 1332 -427 1333 -426
rect 1402 -427 1403 -426
rect 1409 -427 1410 -426
rect 1500 -427 1501 -426
rect 1556 -427 1557 -426
rect 1675 -427 1676 -426
rect 1682 -427 1683 -426
rect 1829 -427 1830 -426
rect 212 -429 213 -428
rect 1059 -429 1060 -428
rect 1083 -429 1084 -428
rect 1661 -429 1662 -428
rect 1689 -429 1690 -428
rect 1808 -429 1809 -428
rect 268 -431 269 -430
rect 905 -431 906 -430
rect 968 -431 969 -430
rect 1647 -431 1648 -430
rect 1703 -431 1704 -430
rect 1836 -431 1837 -430
rect 296 -433 297 -432
rect 779 -433 780 -432
rect 803 -433 804 -432
rect 1332 -433 1333 -432
rect 1367 -433 1368 -432
rect 1479 -433 1480 -432
rect 1486 -433 1487 -432
rect 1584 -433 1585 -432
rect 1619 -433 1620 -432
rect 1738 -433 1739 -432
rect 296 -435 297 -434
rect 786 -435 787 -434
rect 807 -435 808 -434
rect 1122 -435 1123 -434
rect 1192 -435 1193 -434
rect 1290 -435 1291 -434
rect 1437 -435 1438 -434
rect 1507 -435 1508 -434
rect 1514 -435 1515 -434
rect 1619 -435 1620 -434
rect 1626 -435 1627 -434
rect 1745 -435 1746 -434
rect 303 -437 304 -436
rect 485 -437 486 -436
rect 632 -437 633 -436
rect 786 -437 787 -436
rect 842 -437 843 -436
rect 1409 -437 1410 -436
rect 1423 -437 1424 -436
rect 1514 -437 1515 -436
rect 1521 -437 1522 -436
rect 1626 -437 1627 -436
rect 1640 -437 1641 -436
rect 1724 -437 1725 -436
rect 1731 -437 1732 -436
rect 1885 -437 1886 -436
rect 177 -439 178 -438
rect 303 -439 304 -438
rect 310 -439 311 -438
rect 569 -439 570 -438
rect 632 -439 633 -438
rect 877 -439 878 -438
rect 887 -439 888 -438
rect 1640 -439 1641 -438
rect 1717 -439 1718 -438
rect 1829 -439 1830 -438
rect 177 -441 178 -440
rect 338 -441 339 -440
rect 408 -441 409 -440
rect 520 -441 521 -440
rect 719 -441 720 -440
rect 1423 -441 1424 -440
rect 1444 -441 1445 -440
rect 1521 -441 1522 -440
rect 1577 -441 1578 -440
rect 1689 -441 1690 -440
rect 107 -443 108 -442
rect 408 -443 409 -442
rect 415 -443 416 -442
rect 639 -443 640 -442
rect 775 -443 776 -442
rect 1444 -443 1445 -442
rect 1451 -443 1452 -442
rect 1577 -443 1578 -442
rect 1598 -443 1599 -442
rect 1717 -443 1718 -442
rect 107 -445 108 -444
rect 275 -445 276 -444
rect 310 -445 311 -444
rect 366 -445 367 -444
rect 429 -445 430 -444
rect 618 -445 619 -444
rect 814 -445 815 -444
rect 842 -445 843 -444
rect 870 -445 871 -444
rect 1227 -445 1228 -444
rect 1241 -445 1242 -444
rect 1556 -445 1557 -444
rect 1605 -445 1606 -444
rect 1731 -445 1732 -444
rect 2 -447 3 -446
rect 618 -447 619 -446
rect 821 -447 822 -446
rect 877 -447 878 -446
rect 905 -447 906 -446
rect 940 -447 941 -446
rect 1010 -447 1011 -446
rect 1241 -447 1242 -446
rect 1255 -447 1256 -446
rect 1451 -447 1452 -446
rect 1458 -447 1459 -446
rect 1605 -447 1606 -446
rect 58 -449 59 -448
rect 814 -449 815 -448
rect 870 -449 871 -448
rect 1080 -449 1081 -448
rect 1083 -449 1084 -448
rect 1395 -449 1396 -448
rect 1465 -449 1466 -448
rect 1570 -449 1571 -448
rect 128 -451 129 -450
rect 366 -451 367 -450
rect 450 -451 451 -450
rect 1703 -451 1704 -450
rect 128 -453 129 -452
rect 142 -453 143 -452
rect 198 -453 199 -452
rect 639 -453 640 -452
rect 695 -453 696 -452
rect 821 -453 822 -452
rect 940 -453 941 -452
rect 1150 -453 1151 -452
rect 1181 -453 1182 -452
rect 1458 -453 1459 -452
rect 1486 -453 1487 -452
rect 1822 -453 1823 -452
rect 142 -455 143 -454
rect 926 -455 927 -454
rect 1010 -455 1011 -454
rect 1038 -455 1039 -454
rect 1066 -455 1067 -454
rect 1192 -455 1193 -454
rect 1220 -455 1221 -454
rect 1311 -455 1312 -454
rect 1318 -455 1319 -454
rect 1465 -455 1466 -454
rect 1696 -455 1697 -454
rect 1822 -455 1823 -454
rect 184 -457 185 -456
rect 695 -457 696 -456
rect 726 -457 727 -456
rect 1255 -457 1256 -456
rect 1269 -457 1270 -456
rect 1395 -457 1396 -456
rect 1535 -457 1536 -456
rect 1696 -457 1697 -456
rect 184 -459 185 -458
rect 576 -459 577 -458
rect 1038 -459 1039 -458
rect 1052 -459 1053 -458
rect 1066 -459 1067 -458
rect 1955 -459 1956 -458
rect 198 -461 199 -460
rect 352 -461 353 -460
rect 450 -461 451 -460
rect 723 -461 724 -460
rect 898 -461 899 -460
rect 1052 -461 1053 -460
rect 1101 -461 1102 -460
rect 1598 -461 1599 -460
rect 219 -463 220 -462
rect 926 -463 927 -462
rect 1045 -463 1046 -462
rect 1101 -463 1102 -462
rect 1108 -463 1109 -462
rect 1150 -463 1151 -462
rect 1199 -463 1200 -462
rect 1269 -463 1270 -462
rect 1283 -463 1284 -462
rect 1367 -463 1368 -462
rect 1416 -463 1417 -462
rect 1535 -463 1536 -462
rect 275 -465 276 -464
rect 387 -465 388 -464
rect 576 -465 577 -464
rect 604 -465 605 -464
rect 723 -465 724 -464
rect 1374 -465 1375 -464
rect 289 -467 290 -466
rect 387 -467 388 -466
rect 583 -467 584 -466
rect 604 -467 605 -466
rect 849 -467 850 -466
rect 1283 -467 1284 -466
rect 1339 -467 1340 -466
rect 1416 -467 1417 -466
rect 282 -469 283 -468
rect 289 -469 290 -468
rect 317 -469 318 -468
rect 457 -469 458 -468
rect 583 -469 584 -468
rect 796 -469 797 -468
rect 898 -469 899 -468
rect 954 -469 955 -468
rect 961 -469 962 -468
rect 1108 -469 1109 -468
rect 1115 -469 1116 -468
rect 1220 -469 1221 -468
rect 1276 -469 1277 -468
rect 1339 -469 1340 -468
rect 1374 -469 1375 -468
rect 1381 -469 1382 -468
rect 254 -471 255 -470
rect 282 -471 283 -470
rect 317 -471 318 -470
rect 716 -471 717 -470
rect 740 -471 741 -470
rect 1115 -471 1116 -470
rect 1171 -471 1172 -470
rect 1199 -471 1200 -470
rect 1206 -471 1207 -470
rect 1318 -471 1319 -470
rect 254 -473 255 -472
rect 597 -473 598 -472
rect 863 -473 864 -472
rect 954 -473 955 -472
rect 992 -473 993 -472
rect 1171 -473 1172 -472
rect 1213 -473 1214 -472
rect 1276 -473 1277 -472
rect 1304 -473 1305 -472
rect 1381 -473 1382 -472
rect 324 -475 325 -474
rect 737 -475 738 -474
rect 919 -475 920 -474
rect 1045 -475 1046 -474
rect 1143 -475 1144 -474
rect 1206 -475 1207 -474
rect 1234 -475 1235 -474
rect 1304 -475 1305 -474
rect 324 -477 325 -476
rect 422 -477 423 -476
rect 464 -477 465 -476
rect 597 -477 598 -476
rect 919 -477 920 -476
rect 989 -477 990 -476
rect 1094 -477 1095 -476
rect 1143 -477 1144 -476
rect 1157 -477 1158 -476
rect 1234 -477 1235 -476
rect 331 -479 332 -478
rect 380 -479 381 -478
rect 422 -479 423 -478
rect 534 -479 535 -478
rect 947 -479 948 -478
rect 961 -479 962 -478
rect 975 -479 976 -478
rect 1213 -479 1214 -478
rect 93 -481 94 -480
rect 380 -481 381 -480
rect 933 -481 934 -480
rect 947 -481 948 -480
rect 989 -481 990 -480
rect 1927 -481 1928 -480
rect 93 -483 94 -482
rect 534 -483 535 -482
rect 933 -483 934 -482
rect 1563 -483 1564 -482
rect 338 -485 339 -484
rect 394 -485 395 -484
rect 996 -485 997 -484
rect 1094 -485 1095 -484
rect 261 -487 262 -486
rect 394 -487 395 -486
rect 835 -487 836 -486
rect 996 -487 997 -486
rect 1003 -487 1004 -486
rect 1157 -487 1158 -486
rect 261 -489 262 -488
rect 660 -489 661 -488
rect 54 -491 55 -490
rect 660 -491 661 -490
rect 352 -493 353 -492
rect 1027 -493 1028 -492
rect 555 -495 556 -494
rect 835 -495 836 -494
rect 492 -497 493 -496
rect 555 -497 556 -496
rect 492 -499 493 -498
rect 1185 -499 1186 -498
rect 30 -510 31 -509
rect 72 -510 73 -509
rect 93 -510 94 -509
rect 173 -510 174 -509
rect 205 -510 206 -509
rect 733 -510 734 -509
rect 737 -510 738 -509
rect 1633 -510 1634 -509
rect 1682 -510 1683 -509
rect 2151 -510 2152 -509
rect 2214 -510 2215 -509
rect 2291 -510 2292 -509
rect 37 -512 38 -511
rect 646 -512 647 -511
rect 656 -512 657 -511
rect 695 -512 696 -511
rect 723 -512 724 -511
rect 772 -512 773 -511
rect 824 -512 825 -511
rect 1129 -512 1130 -511
rect 1146 -512 1147 -511
rect 1374 -512 1375 -511
rect 1535 -512 1536 -511
rect 2032 -512 2033 -511
rect 2039 -512 2040 -511
rect 2172 -512 2173 -511
rect 2263 -512 2264 -511
rect 2361 -512 2362 -511
rect 44 -514 45 -513
rect 212 -514 213 -513
rect 215 -514 216 -513
rect 1766 -514 1767 -513
rect 1836 -514 1837 -513
rect 2004 -514 2005 -513
rect 2014 -514 2015 -513
rect 2179 -514 2180 -513
rect 2284 -514 2285 -513
rect 2326 -514 2327 -513
rect 44 -516 45 -515
rect 166 -516 167 -515
rect 170 -516 171 -515
rect 450 -516 451 -515
rect 541 -516 542 -515
rect 632 -516 633 -515
rect 635 -516 636 -515
rect 772 -516 773 -515
rect 842 -516 843 -515
rect 884 -516 885 -515
rect 898 -516 899 -515
rect 968 -516 969 -515
rect 982 -516 983 -515
rect 1752 -516 1753 -515
rect 1864 -516 1865 -515
rect 2046 -516 2047 -515
rect 2088 -516 2089 -515
rect 2210 -516 2211 -515
rect 135 -518 136 -517
rect 737 -518 738 -517
rect 751 -518 752 -517
rect 754 -518 755 -517
rect 786 -518 787 -517
rect 842 -518 843 -517
rect 849 -518 850 -517
rect 919 -518 920 -517
rect 975 -518 976 -517
rect 1752 -518 1753 -517
rect 1864 -518 1865 -517
rect 1979 -518 1980 -517
rect 1983 -518 1984 -517
rect 2158 -518 2159 -517
rect 75 -520 76 -519
rect 919 -520 920 -519
rect 985 -520 986 -519
rect 1766 -520 1767 -519
rect 1794 -520 1795 -519
rect 1983 -520 1984 -519
rect 1990 -520 1991 -519
rect 2007 -520 2008 -519
rect 2116 -520 2117 -519
rect 2193 -520 2194 -519
rect 114 -522 115 -521
rect 975 -522 976 -521
rect 992 -522 993 -521
rect 1213 -522 1214 -521
rect 1269 -522 1270 -521
rect 1374 -522 1375 -521
rect 1472 -522 1473 -521
rect 1535 -522 1536 -521
rect 1612 -522 1613 -521
rect 1794 -522 1795 -521
rect 1808 -522 1809 -521
rect 1990 -522 1991 -521
rect 2116 -522 2117 -521
rect 2224 -522 2225 -521
rect 114 -524 115 -523
rect 331 -524 332 -523
rect 380 -524 381 -523
rect 989 -524 990 -523
rect 996 -524 997 -523
rect 1125 -524 1126 -523
rect 1164 -524 1165 -523
rect 2137 -524 2138 -523
rect 2144 -524 2145 -523
rect 2200 -524 2201 -523
rect 138 -526 139 -525
rect 898 -526 899 -525
rect 940 -526 941 -525
rect 996 -526 997 -525
rect 1003 -526 1004 -525
rect 1843 -526 1844 -525
rect 1871 -526 1872 -525
rect 2053 -526 2054 -525
rect 163 -528 164 -527
rect 716 -528 717 -527
rect 723 -528 724 -527
rect 1108 -528 1109 -527
rect 1167 -528 1168 -527
rect 1360 -528 1361 -527
rect 1395 -528 1396 -527
rect 1472 -528 1473 -527
rect 1619 -528 1620 -527
rect 1808 -528 1809 -527
rect 1878 -528 1879 -527
rect 2060 -528 2061 -527
rect 205 -530 206 -529
rect 1262 -530 1263 -529
rect 1290 -530 1291 -529
rect 1395 -530 1396 -529
rect 1479 -530 1480 -529
rect 1619 -530 1620 -529
rect 1633 -530 1634 -529
rect 2207 -530 2208 -529
rect 219 -532 220 -531
rect 2081 -532 2082 -531
rect 219 -534 220 -533
rect 653 -534 654 -533
rect 660 -534 661 -533
rect 1006 -534 1007 -533
rect 1017 -534 1018 -533
rect 1108 -534 1109 -533
rect 1192 -534 1193 -533
rect 1269 -534 1270 -533
rect 1290 -534 1291 -533
rect 1367 -534 1368 -533
rect 1479 -534 1480 -533
rect 2021 -534 2022 -533
rect 79 -536 80 -535
rect 653 -536 654 -535
rect 702 -536 703 -535
rect 1003 -536 1004 -535
rect 1024 -536 1025 -535
rect 1346 -536 1347 -535
rect 1367 -536 1368 -535
rect 1486 -536 1487 -535
rect 1640 -536 1641 -535
rect 1836 -536 1837 -535
rect 1885 -536 1886 -535
rect 2067 -536 2068 -535
rect 222 -538 223 -537
rect 282 -538 283 -537
rect 310 -538 311 -537
rect 663 -538 664 -537
rect 716 -538 717 -537
rect 726 -538 727 -537
rect 730 -538 731 -537
rect 989 -538 990 -537
rect 1031 -538 1032 -537
rect 1122 -538 1123 -537
rect 1136 -538 1137 -537
rect 1192 -538 1193 -537
rect 1227 -538 1228 -537
rect 1346 -538 1347 -537
rect 1493 -538 1494 -537
rect 1640 -538 1641 -537
rect 1661 -538 1662 -537
rect 2039 -538 2040 -537
rect 103 -540 104 -539
rect 1493 -540 1494 -539
rect 1710 -540 1711 -539
rect 1871 -540 1872 -539
rect 1899 -540 1900 -539
rect 2074 -540 2075 -539
rect 226 -542 227 -541
rect 236 -542 237 -541
rect 240 -542 241 -541
rect 310 -542 311 -541
rect 324 -542 325 -541
rect 492 -542 493 -541
rect 534 -542 535 -541
rect 1213 -542 1214 -541
rect 1255 -542 1256 -541
rect 1360 -542 1361 -541
rect 1717 -542 1718 -541
rect 1878 -542 1879 -541
rect 1906 -542 1907 -541
rect 2109 -542 2110 -541
rect 65 -544 66 -543
rect 226 -544 227 -543
rect 233 -544 234 -543
rect 1717 -544 1718 -543
rect 1731 -544 1732 -543
rect 2102 -544 2103 -543
rect 9 -546 10 -545
rect 65 -546 66 -545
rect 72 -546 73 -545
rect 240 -546 241 -545
rect 254 -546 255 -545
rect 597 -546 598 -545
rect 600 -546 601 -545
rect 1437 -546 1438 -545
rect 1570 -546 1571 -545
rect 1731 -546 1732 -545
rect 1738 -546 1739 -545
rect 1899 -546 1900 -545
rect 1913 -546 1914 -545
rect 2130 -546 2131 -545
rect 9 -548 10 -547
rect 198 -548 199 -547
rect 233 -548 234 -547
rect 429 -548 430 -547
rect 450 -548 451 -547
rect 513 -548 514 -547
rect 541 -548 542 -547
rect 740 -548 741 -547
rect 751 -548 752 -547
rect 905 -548 906 -547
rect 947 -548 948 -547
rect 1017 -548 1018 -547
rect 1034 -548 1035 -547
rect 1934 -548 1935 -547
rect 1941 -548 1942 -547
rect 2095 -548 2096 -547
rect 107 -550 108 -549
rect 198 -550 199 -549
rect 282 -550 283 -549
rect 387 -550 388 -549
rect 394 -550 395 -549
rect 1013 -550 1014 -549
rect 1062 -550 1063 -549
rect 2025 -550 2026 -549
rect 16 -552 17 -551
rect 107 -552 108 -551
rect 177 -552 178 -551
rect 254 -552 255 -551
rect 317 -552 318 -551
rect 324 -552 325 -551
rect 331 -552 332 -551
rect 537 -552 538 -551
rect 565 -552 566 -551
rect 1241 -552 1242 -551
rect 1262 -552 1263 -551
rect 1955 -552 1956 -551
rect 1962 -552 1963 -551
rect 2123 -552 2124 -551
rect 16 -554 17 -553
rect 156 -554 157 -553
rect 177 -554 178 -553
rect 887 -554 888 -553
rect 891 -554 892 -553
rect 968 -554 969 -553
rect 978 -554 979 -553
rect 1738 -554 1739 -553
rect 1759 -554 1760 -553
rect 1941 -554 1942 -553
rect 1948 -554 1949 -553
rect 2165 -554 2166 -553
rect 93 -556 94 -555
rect 537 -556 538 -555
rect 569 -556 570 -555
rect 593 -556 594 -555
rect 611 -556 612 -555
rect 702 -556 703 -555
rect 786 -556 787 -555
rect 1612 -556 1613 -555
rect 1675 -556 1676 -555
rect 1906 -556 1907 -555
rect 1920 -556 1921 -555
rect 1955 -556 1956 -555
rect 1969 -556 1970 -555
rect 2144 -556 2145 -555
rect 121 -558 122 -557
rect 156 -558 157 -557
rect 303 -558 304 -557
rect 317 -558 318 -557
rect 345 -558 346 -557
rect 429 -558 430 -557
rect 492 -558 493 -557
rect 562 -558 563 -557
rect 569 -558 570 -557
rect 744 -558 745 -557
rect 835 -558 836 -557
rect 891 -558 892 -557
rect 905 -558 906 -557
rect 961 -558 962 -557
rect 1031 -558 1032 -557
rect 1241 -558 1242 -557
rect 1283 -558 1284 -557
rect 1570 -558 1571 -557
rect 1591 -558 1592 -557
rect 1759 -558 1760 -557
rect 1773 -558 1774 -557
rect 1948 -558 1949 -557
rect 1976 -558 1977 -557
rect 1997 -558 1998 -557
rect 121 -560 122 -559
rect 548 -560 549 -559
rect 604 -560 605 -559
rect 611 -560 612 -559
rect 621 -560 622 -559
rect 870 -560 871 -559
rect 877 -560 878 -559
rect 1227 -560 1228 -559
rect 1297 -560 1298 -559
rect 1591 -560 1592 -559
rect 1696 -560 1697 -559
rect 1934 -560 1935 -559
rect 100 -562 101 -561
rect 548 -562 549 -561
rect 649 -562 650 -561
rect 1843 -562 1844 -561
rect 1927 -562 1928 -561
rect 2088 -562 2089 -561
rect 100 -564 101 -563
rect 639 -564 640 -563
rect 688 -564 689 -563
rect 730 -564 731 -563
rect 754 -564 755 -563
rect 961 -564 962 -563
rect 985 -564 986 -563
rect 1696 -564 1697 -563
rect 1703 -564 1704 -563
rect 1927 -564 1928 -563
rect 61 -566 62 -565
rect 688 -566 689 -565
rect 793 -566 794 -565
rect 870 -566 871 -565
rect 1073 -566 1074 -565
rect 1129 -566 1130 -565
rect 1150 -566 1151 -565
rect 1255 -566 1256 -565
rect 1297 -566 1298 -565
rect 1801 -566 1802 -565
rect 1829 -566 1830 -565
rect 1885 -566 1886 -565
rect 2 -568 3 -567
rect 61 -568 62 -567
rect 303 -568 304 -567
rect 527 -568 528 -567
rect 639 -568 640 -567
rect 709 -568 710 -567
rect 793 -568 794 -567
rect 828 -568 829 -567
rect 852 -568 853 -567
rect 1038 -568 1039 -567
rect 1080 -568 1081 -567
rect 1710 -568 1711 -567
rect 1724 -568 1725 -567
rect 1962 -568 1963 -567
rect 250 -570 251 -569
rect 1038 -570 1039 -569
rect 1083 -570 1084 -569
rect 1787 -570 1788 -569
rect 338 -572 339 -571
rect 345 -572 346 -571
rect 366 -572 367 -571
rect 380 -572 381 -571
rect 387 -572 388 -571
rect 432 -572 433 -571
rect 436 -572 437 -571
rect 604 -572 605 -571
rect 709 -572 710 -571
rect 758 -572 759 -571
rect 765 -572 766 -571
rect 828 -572 829 -571
rect 863 -572 864 -571
rect 947 -572 948 -571
rect 971 -572 972 -571
rect 1724 -572 1725 -571
rect 1745 -572 1746 -571
rect 1920 -572 1921 -571
rect 142 -574 143 -573
rect 765 -574 766 -573
rect 821 -574 822 -573
rect 835 -574 836 -573
rect 863 -574 864 -573
rect 1647 -574 1648 -573
rect 1703 -574 1704 -573
rect 1822 -574 1823 -573
rect 142 -576 143 -575
rect 401 -576 402 -575
rect 408 -576 409 -575
rect 513 -576 514 -575
rect 527 -576 528 -575
rect 555 -576 556 -575
rect 695 -576 696 -575
rect 821 -576 822 -575
rect 954 -576 955 -575
rect 1745 -576 1746 -575
rect 1780 -576 1781 -575
rect 1969 -576 1970 -575
rect 117 -578 118 -577
rect 401 -578 402 -577
rect 415 -578 416 -577
rect 810 -578 811 -577
rect 856 -578 857 -577
rect 954 -578 955 -577
rect 1010 -578 1011 -577
rect 1073 -578 1074 -577
rect 1094 -578 1095 -577
rect 1164 -578 1165 -577
rect 1216 -578 1217 -577
rect 1997 -578 1998 -577
rect 275 -580 276 -579
rect 408 -580 409 -579
rect 422 -580 423 -579
rect 436 -580 437 -579
rect 495 -580 496 -579
rect 744 -580 745 -579
rect 758 -580 759 -579
rect 779 -580 780 -579
rect 800 -580 801 -579
rect 856 -580 857 -579
rect 1010 -580 1011 -579
rect 1976 -580 1977 -579
rect 86 -582 87 -581
rect 800 -582 801 -581
rect 1094 -582 1095 -581
rect 1682 -582 1683 -581
rect 86 -584 87 -583
rect 352 -584 353 -583
rect 359 -584 360 -583
rect 422 -584 423 -583
rect 506 -584 507 -583
rect 562 -584 563 -583
rect 586 -584 587 -583
rect 1780 -584 1781 -583
rect 58 -586 59 -585
rect 352 -586 353 -585
rect 359 -586 360 -585
rect 478 -586 479 -585
rect 555 -586 556 -585
rect 681 -586 682 -585
rect 1101 -586 1102 -585
rect 1136 -586 1137 -585
rect 1220 -586 1221 -585
rect 1283 -586 1284 -585
rect 1325 -586 1326 -585
rect 1661 -586 1662 -585
rect 23 -588 24 -587
rect 1325 -588 1326 -587
rect 1332 -588 1333 -587
rect 2011 -588 2012 -587
rect 23 -590 24 -589
rect 51 -590 52 -589
rect 275 -590 276 -589
rect 457 -590 458 -589
rect 471 -590 472 -589
rect 506 -590 507 -589
rect 674 -590 675 -589
rect 779 -590 780 -589
rect 1080 -590 1081 -589
rect 1101 -590 1102 -589
rect 1199 -590 1200 -589
rect 1220 -590 1221 -589
rect 1234 -590 1235 -589
rect 1332 -590 1333 -589
rect 1353 -590 1354 -589
rect 1437 -590 1438 -589
rect 1465 -590 1466 -589
rect 1913 -590 1914 -589
rect 51 -592 52 -591
rect 625 -592 626 -591
rect 667 -592 668 -591
rect 674 -592 675 -591
rect 681 -592 682 -591
rect 1150 -592 1151 -591
rect 1248 -592 1249 -591
rect 1353 -592 1354 -591
rect 1416 -592 1417 -591
rect 1773 -592 1774 -591
rect 1850 -592 1851 -591
rect 2011 -592 2012 -591
rect 135 -594 136 -593
rect 457 -594 458 -593
rect 464 -594 465 -593
rect 625 -594 626 -593
rect 1157 -594 1158 -593
rect 1248 -594 1249 -593
rect 1318 -594 1319 -593
rect 1465 -594 1466 -593
rect 1500 -594 1501 -593
rect 1647 -594 1648 -593
rect 184 -596 185 -595
rect 464 -596 465 -595
rect 576 -596 577 -595
rect 667 -596 668 -595
rect 1087 -596 1088 -595
rect 1157 -596 1158 -595
rect 1311 -596 1312 -595
rect 1318 -596 1319 -595
rect 1402 -596 1403 -595
rect 1500 -596 1501 -595
rect 1521 -596 1522 -595
rect 1675 -596 1676 -595
rect 184 -598 185 -597
rect 261 -598 262 -597
rect 289 -598 290 -597
rect 471 -598 472 -597
rect 576 -598 577 -597
rect 590 -598 591 -597
rect 618 -598 619 -597
rect 1234 -598 1235 -597
rect 1304 -598 1305 -597
rect 1402 -598 1403 -597
rect 1416 -598 1417 -597
rect 2018 -598 2019 -597
rect 149 -600 150 -599
rect 261 -600 262 -599
rect 289 -600 290 -599
rect 933 -600 934 -599
rect 1206 -600 1207 -599
rect 1311 -600 1312 -599
rect 1430 -600 1431 -599
rect 1521 -600 1522 -599
rect 1528 -600 1529 -599
rect 1829 -600 1830 -599
rect 1857 -600 1858 -599
rect 2018 -600 2019 -599
rect 149 -602 150 -601
rect 247 -602 248 -601
rect 338 -602 339 -601
rect 940 -602 941 -601
rect 1115 -602 1116 -601
rect 1206 -602 1207 -601
rect 1440 -602 1441 -601
rect 1850 -602 1851 -601
rect 79 -604 80 -603
rect 247 -604 248 -603
rect 366 -604 367 -603
rect 849 -604 850 -603
rect 912 -604 913 -603
rect 1304 -604 1305 -603
rect 1528 -604 1529 -603
rect 1577 -604 1578 -603
rect 1598 -604 1599 -603
rect 1787 -604 1788 -603
rect 373 -606 374 -605
rect 478 -606 479 -605
rect 590 -606 591 -605
rect 877 -606 878 -605
rect 929 -606 930 -605
rect 1087 -606 1088 -605
rect 1178 -606 1179 -605
rect 1430 -606 1431 -605
rect 1458 -606 1459 -605
rect 1598 -606 1599 -605
rect 1605 -606 1606 -605
rect 1822 -606 1823 -605
rect 191 -608 192 -607
rect 373 -608 374 -607
rect 394 -608 395 -607
rect 499 -608 500 -607
rect 807 -608 808 -607
rect 912 -608 913 -607
rect 933 -608 934 -607
rect 936 -608 937 -607
rect 1045 -608 1046 -607
rect 1115 -608 1116 -607
rect 1143 -608 1144 -607
rect 1178 -608 1179 -607
rect 1388 -608 1389 -607
rect 1458 -608 1459 -607
rect 1507 -608 1508 -607
rect 1577 -608 1578 -607
rect 1668 -608 1669 -607
rect 1857 -608 1858 -607
rect 173 -610 174 -609
rect 191 -610 192 -609
rect 443 -610 444 -609
rect 618 -610 619 -609
rect 926 -610 927 -609
rect 1045 -610 1046 -609
rect 1143 -610 1144 -609
rect 1815 -610 1816 -609
rect 443 -612 444 -611
rect 520 -612 521 -611
rect 926 -612 927 -611
rect 1542 -612 1543 -611
rect 1549 -612 1550 -611
rect 1801 -612 1802 -611
rect 485 -614 486 -613
rect 520 -614 521 -613
rect 1202 -614 1203 -613
rect 1542 -614 1543 -613
rect 1626 -614 1627 -613
rect 1815 -614 1816 -613
rect 485 -616 486 -615
rect 583 -616 584 -615
rect 1276 -616 1277 -615
rect 1388 -616 1389 -615
rect 1423 -616 1424 -615
rect 1605 -616 1606 -615
rect 1668 -616 1669 -615
rect 1689 -616 1690 -615
rect 499 -618 500 -617
rect 660 -618 661 -617
rect 1185 -618 1186 -617
rect 1276 -618 1277 -617
rect 1339 -618 1340 -617
rect 1423 -618 1424 -617
rect 1444 -618 1445 -617
rect 1549 -618 1550 -617
rect 1556 -618 1557 -617
rect 1689 -618 1690 -617
rect 583 -620 584 -619
rect 1654 -620 1655 -619
rect 1059 -622 1060 -621
rect 1185 -622 1186 -621
rect 1381 -622 1382 -621
rect 1444 -622 1445 -621
rect 1451 -622 1452 -621
rect 1626 -622 1627 -621
rect 1059 -624 1060 -623
rect 2186 -624 2187 -623
rect 1066 -626 1067 -625
rect 1451 -626 1452 -625
rect 1507 -626 1508 -625
rect 1514 -626 1515 -625
rect 1556 -626 1557 -625
rect 1563 -626 1564 -625
rect 1584 -626 1585 -625
rect 1654 -626 1655 -625
rect 1052 -628 1053 -627
rect 1066 -628 1067 -627
rect 1171 -628 1172 -627
rect 1339 -628 1340 -627
rect 1409 -628 1410 -627
rect 1514 -628 1515 -627
rect 1563 -628 1564 -627
rect 2221 -628 2222 -627
rect 268 -630 269 -629
rect 1052 -630 1053 -629
rect 1199 -630 1200 -629
rect 1381 -630 1382 -629
rect 1409 -630 1410 -629
rect 1958 -630 1959 -629
rect 268 -632 269 -631
rect 415 -632 416 -631
rect 915 -632 916 -631
rect 1171 -632 1172 -631
rect 1489 -632 1490 -631
rect 1584 -632 1585 -631
rect 2 -643 3 -642
rect 121 -643 122 -642
rect 131 -643 132 -642
rect 2137 -643 2138 -642
rect 2144 -643 2145 -642
rect 2319 -643 2320 -642
rect 2326 -643 2327 -642
rect 2347 -643 2348 -642
rect 2361 -643 2362 -642
rect 2403 -643 2404 -642
rect 44 -645 45 -644
rect 1223 -645 1224 -644
rect 1300 -645 1301 -644
rect 2130 -645 2131 -644
rect 2137 -645 2138 -644
rect 2172 -645 2173 -644
rect 2193 -645 2194 -644
rect 2207 -645 2208 -644
rect 2214 -645 2215 -644
rect 2277 -645 2278 -644
rect 2291 -645 2292 -644
rect 2326 -645 2327 -644
rect 47 -647 48 -646
rect 65 -647 66 -646
rect 68 -647 69 -646
rect 754 -647 755 -646
rect 807 -647 808 -646
rect 1122 -647 1123 -646
rect 1143 -647 1144 -646
rect 1591 -647 1592 -646
rect 1703 -647 1704 -646
rect 2235 -647 2236 -646
rect 12 -649 13 -648
rect 65 -649 66 -648
rect 72 -649 73 -648
rect 1780 -649 1781 -648
rect 1843 -649 1844 -648
rect 2221 -649 2222 -648
rect 51 -651 52 -650
rect 926 -651 927 -650
rect 940 -651 941 -650
rect 1906 -651 1907 -650
rect 1955 -651 1956 -650
rect 2256 -651 2257 -650
rect 51 -653 52 -652
rect 681 -653 682 -652
rect 698 -653 699 -652
rect 982 -653 983 -652
rect 1010 -653 1011 -652
rect 2151 -653 2152 -652
rect 2158 -653 2159 -652
rect 2312 -653 2313 -652
rect 58 -655 59 -654
rect 1682 -655 1683 -654
rect 1885 -655 1886 -654
rect 2130 -655 2131 -654
rect 2200 -655 2201 -654
rect 2224 -655 2225 -654
rect 72 -657 73 -656
rect 1003 -657 1004 -656
rect 1059 -657 1060 -656
rect 1626 -657 1627 -656
rect 1885 -657 1886 -656
rect 1969 -657 1970 -656
rect 2004 -657 2005 -656
rect 2144 -657 2145 -656
rect 82 -659 83 -658
rect 1031 -659 1032 -658
rect 1059 -659 1060 -658
rect 1073 -659 1074 -658
rect 1083 -659 1084 -658
rect 1465 -659 1466 -658
rect 1486 -659 1487 -658
rect 2165 -659 2166 -658
rect 16 -661 17 -660
rect 1073 -661 1074 -660
rect 1094 -661 1095 -660
rect 2186 -661 2187 -660
rect 93 -663 94 -662
rect 562 -663 563 -662
rect 618 -663 619 -662
rect 940 -663 941 -662
rect 957 -663 958 -662
rect 1052 -663 1053 -662
rect 1062 -663 1063 -662
rect 2179 -663 2180 -662
rect 93 -665 94 -664
rect 142 -665 143 -664
rect 145 -665 146 -664
rect 943 -665 944 -664
rect 1052 -665 1053 -664
rect 1108 -665 1109 -664
rect 1150 -665 1151 -664
rect 2186 -665 2187 -664
rect 75 -667 76 -666
rect 1108 -667 1109 -666
rect 1136 -667 1137 -666
rect 1150 -667 1151 -666
rect 1174 -667 1175 -666
rect 2305 -667 2306 -666
rect 135 -669 136 -668
rect 1822 -669 1823 -668
rect 1857 -669 1858 -668
rect 2004 -669 2005 -668
rect 2011 -669 2012 -668
rect 2151 -669 2152 -668
rect 170 -671 171 -670
rect 310 -671 311 -670
rect 401 -671 402 -670
rect 1031 -671 1032 -670
rect 1101 -671 1102 -670
rect 1122 -671 1123 -670
rect 1178 -671 1179 -670
rect 1213 -671 1214 -670
rect 1216 -671 1217 -670
rect 2109 -671 2110 -670
rect 2116 -671 2117 -670
rect 2298 -671 2299 -670
rect 173 -673 174 -672
rect 1927 -673 1928 -672
rect 1983 -673 1984 -672
rect 2109 -673 2110 -672
rect 2123 -673 2124 -672
rect 2291 -673 2292 -672
rect 187 -675 188 -674
rect 702 -675 703 -674
rect 733 -675 734 -674
rect 2179 -675 2180 -674
rect 205 -677 206 -676
rect 1451 -677 1452 -676
rect 1493 -677 1494 -676
rect 1626 -677 1627 -676
rect 1717 -677 1718 -676
rect 1822 -677 1823 -676
rect 1864 -677 1865 -676
rect 2011 -677 2012 -676
rect 2018 -677 2019 -676
rect 2158 -677 2159 -676
rect 212 -679 213 -678
rect 747 -679 748 -678
rect 765 -679 766 -678
rect 1003 -679 1004 -678
rect 1101 -679 1102 -678
rect 1111 -679 1112 -678
rect 1199 -679 1200 -678
rect 1983 -679 1984 -678
rect 1990 -679 1991 -678
rect 2123 -679 2124 -678
rect 191 -681 192 -680
rect 212 -681 213 -680
rect 236 -681 237 -680
rect 1178 -681 1179 -680
rect 1213 -681 1214 -680
rect 1409 -681 1410 -680
rect 1430 -681 1431 -680
rect 1591 -681 1592 -680
rect 1605 -681 1606 -680
rect 1717 -681 1718 -680
rect 1738 -681 1739 -680
rect 1857 -681 1858 -680
rect 1990 -681 1991 -680
rect 2067 -681 2068 -680
rect 2074 -681 2075 -680
rect 2242 -681 2243 -680
rect 149 -683 150 -682
rect 191 -683 192 -682
rect 247 -683 248 -682
rect 317 -683 318 -682
rect 366 -683 367 -682
rect 765 -683 766 -682
rect 800 -683 801 -682
rect 807 -683 808 -682
rect 824 -683 825 -682
rect 2284 -683 2285 -682
rect 30 -685 31 -684
rect 317 -685 318 -684
rect 366 -685 367 -684
rect 772 -685 773 -684
rect 849 -685 850 -684
rect 863 -685 864 -684
rect 891 -685 892 -684
rect 926 -685 927 -684
rect 929 -685 930 -684
rect 1955 -685 1956 -684
rect 1962 -685 1963 -684
rect 2067 -685 2068 -684
rect 2081 -685 2082 -684
rect 2249 -685 2250 -684
rect 9 -687 10 -686
rect 863 -687 864 -686
rect 877 -687 878 -686
rect 891 -687 892 -686
rect 1080 -687 1081 -686
rect 1738 -687 1739 -686
rect 1752 -687 1753 -686
rect 2074 -687 2075 -686
rect 2088 -687 2089 -686
rect 2263 -687 2264 -686
rect 19 -689 20 -688
rect 2081 -689 2082 -688
rect 2095 -689 2096 -688
rect 2270 -689 2271 -688
rect 30 -691 31 -690
rect 37 -691 38 -690
rect 149 -691 150 -690
rect 985 -691 986 -690
rect 1080 -691 1081 -690
rect 1087 -691 1088 -690
rect 1129 -691 1130 -690
rect 1199 -691 1200 -690
rect 1360 -691 1361 -690
rect 1451 -691 1452 -690
rect 1549 -691 1550 -690
rect 1682 -691 1683 -690
rect 1759 -691 1760 -690
rect 2095 -691 2096 -690
rect 37 -693 38 -692
rect 723 -693 724 -692
rect 730 -693 731 -692
rect 1493 -693 1494 -692
rect 1556 -693 1557 -692
rect 1969 -693 1970 -692
rect 1976 -693 1977 -692
rect 2088 -693 2089 -692
rect 261 -695 262 -694
rect 362 -695 363 -694
rect 401 -695 402 -694
rect 555 -695 556 -694
rect 562 -695 563 -694
rect 667 -695 668 -694
rect 681 -695 682 -694
rect 1710 -695 1711 -694
rect 1794 -695 1795 -694
rect 1927 -695 1928 -694
rect 1997 -695 1998 -694
rect 2116 -695 2117 -694
rect 156 -697 157 -696
rect 261 -697 262 -696
rect 282 -697 283 -696
rect 583 -697 584 -696
rect 590 -697 591 -696
rect 667 -697 668 -696
rect 702 -697 703 -696
rect 1304 -697 1305 -696
rect 1360 -697 1361 -696
rect 1773 -697 1774 -696
rect 1829 -697 1830 -696
rect 1962 -697 1963 -696
rect 2025 -697 2026 -696
rect 2165 -697 2166 -696
rect 128 -699 129 -698
rect 156 -699 157 -698
rect 240 -699 241 -698
rect 282 -699 283 -698
rect 310 -699 311 -698
rect 506 -699 507 -698
rect 523 -699 524 -698
rect 1486 -699 1487 -698
rect 1507 -699 1508 -698
rect 1794 -699 1795 -698
rect 1829 -699 1830 -698
rect 1941 -699 1942 -698
rect 2039 -699 2040 -698
rect 2217 -699 2218 -698
rect 114 -701 115 -700
rect 240 -701 241 -700
rect 324 -701 325 -700
rect 506 -701 507 -700
rect 548 -701 549 -700
rect 565 -701 566 -700
rect 569 -701 570 -700
rect 800 -701 801 -700
rect 814 -701 815 -700
rect 849 -701 850 -700
rect 852 -701 853 -700
rect 1745 -701 1746 -700
rect 1808 -701 1809 -700
rect 1941 -701 1942 -700
rect 2046 -701 2047 -700
rect 2172 -701 2173 -700
rect 86 -703 87 -702
rect 114 -703 115 -702
rect 324 -703 325 -702
rect 464 -703 465 -702
rect 492 -703 493 -702
rect 684 -703 685 -702
rect 744 -703 745 -702
rect 2207 -703 2208 -702
rect 5 -705 6 -704
rect 86 -705 87 -704
rect 415 -705 416 -704
rect 464 -705 465 -704
rect 492 -705 493 -704
rect 695 -705 696 -704
rect 747 -705 748 -704
rect 2102 -705 2103 -704
rect 408 -707 409 -706
rect 415 -707 416 -706
rect 429 -707 430 -706
rect 555 -707 556 -706
rect 590 -707 591 -706
rect 1465 -707 1466 -706
rect 1584 -707 1585 -706
rect 1703 -707 1704 -706
rect 1836 -707 1837 -706
rect 1976 -707 1977 -706
rect 2053 -707 2054 -706
rect 2200 -707 2201 -706
rect 303 -709 304 -708
rect 408 -709 409 -708
rect 422 -709 423 -708
rect 429 -709 430 -708
rect 432 -709 433 -708
rect 625 -709 626 -708
rect 639 -709 640 -708
rect 1780 -709 1781 -708
rect 1850 -709 1851 -708
rect 1997 -709 1998 -708
rect 2060 -709 2061 -708
rect 2193 -709 2194 -708
rect 100 -711 101 -710
rect 639 -711 640 -710
rect 646 -711 647 -710
rect 1227 -711 1228 -710
rect 1248 -711 1249 -710
rect 1759 -711 1760 -710
rect 1871 -711 1872 -710
rect 2025 -711 2026 -710
rect 100 -713 101 -712
rect 198 -713 199 -712
rect 219 -713 220 -712
rect 303 -713 304 -712
rect 422 -713 423 -712
rect 1202 -713 1203 -712
rect 1248 -713 1249 -712
rect 1458 -713 1459 -712
rect 1528 -713 1529 -712
rect 1871 -713 1872 -712
rect 1878 -713 1879 -712
rect 2046 -713 2047 -712
rect 163 -715 164 -714
rect 198 -715 199 -714
rect 443 -715 444 -714
rect 548 -715 549 -714
rect 604 -715 605 -714
rect 618 -715 619 -714
rect 653 -715 654 -714
rect 789 -715 790 -714
rect 814 -715 815 -714
rect 870 -715 871 -714
rect 947 -715 948 -714
rect 1129 -715 1130 -714
rect 1136 -715 1137 -714
rect 1745 -715 1746 -714
rect 1899 -715 1900 -714
rect 2039 -715 2040 -714
rect 163 -717 164 -716
rect 485 -717 486 -716
rect 534 -717 535 -716
rect 569 -717 570 -716
rect 576 -717 577 -716
rect 604 -717 605 -716
rect 611 -717 612 -716
rect 625 -717 626 -716
rect 660 -717 661 -716
rect 2228 -717 2229 -716
rect 23 -719 24 -718
rect 485 -719 486 -718
rect 583 -719 584 -718
rect 947 -719 948 -718
rect 996 -719 997 -718
rect 1087 -719 1088 -718
rect 1097 -719 1098 -718
rect 1528 -719 1529 -718
rect 1598 -719 1599 -718
rect 1710 -719 1711 -718
rect 1724 -719 1725 -718
rect 1836 -719 1837 -718
rect 1920 -719 1921 -718
rect 2060 -719 2061 -718
rect 23 -721 24 -720
rect 744 -721 745 -720
rect 772 -721 773 -720
rect 779 -721 780 -720
rect 793 -721 794 -720
rect 870 -721 871 -720
rect 989 -721 990 -720
rect 996 -721 997 -720
rect 1045 -721 1046 -720
rect 1556 -721 1557 -720
rect 1598 -721 1599 -720
rect 1675 -721 1676 -720
rect 1689 -721 1690 -720
rect 1808 -721 1809 -720
rect 1920 -721 1921 -720
rect 1948 -721 1949 -720
rect 289 -723 290 -722
rect 653 -723 654 -722
rect 663 -723 664 -722
rect 709 -723 710 -722
rect 758 -723 759 -722
rect 793 -723 794 -722
rect 1045 -723 1046 -722
rect 1066 -723 1067 -722
rect 1143 -723 1144 -722
rect 2102 -723 2103 -722
rect 184 -725 185 -724
rect 758 -725 759 -724
rect 779 -725 780 -724
rect 1115 -725 1116 -724
rect 1192 -725 1193 -724
rect 1227 -725 1228 -724
rect 1255 -725 1256 -724
rect 1304 -725 1305 -724
rect 1367 -725 1368 -724
rect 1430 -725 1431 -724
rect 1437 -725 1438 -724
rect 1549 -725 1550 -724
rect 1570 -725 1571 -724
rect 1689 -725 1690 -724
rect 1731 -725 1732 -724
rect 1850 -725 1851 -724
rect 1934 -725 1935 -724
rect 2053 -725 2054 -724
rect 184 -727 185 -726
rect 716 -727 717 -726
rect 898 -727 899 -726
rect 1066 -727 1067 -726
rect 1171 -727 1172 -726
rect 1437 -727 1438 -726
rect 1577 -727 1578 -726
rect 1675 -727 1676 -726
rect 1766 -727 1767 -726
rect 1899 -727 1900 -726
rect 177 -729 178 -728
rect 716 -729 717 -728
rect 898 -729 899 -728
rect 1146 -729 1147 -728
rect 1171 -729 1172 -728
rect 1409 -729 1410 -728
rect 1423 -729 1424 -728
rect 1570 -729 1571 -728
rect 1605 -729 1606 -728
rect 1640 -729 1641 -728
rect 1647 -729 1648 -728
rect 1773 -729 1774 -728
rect 1801 -729 1802 -728
rect 1934 -729 1935 -728
rect 58 -731 59 -730
rect 1146 -731 1147 -730
rect 1234 -731 1235 -730
rect 1255 -731 1256 -730
rect 1290 -731 1291 -730
rect 1584 -731 1585 -730
rect 1612 -731 1613 -730
rect 1724 -731 1725 -730
rect 1815 -731 1816 -730
rect 1948 -731 1949 -730
rect 177 -733 178 -732
rect 1269 -733 1270 -732
rect 1339 -733 1340 -732
rect 1423 -733 1424 -732
rect 1444 -733 1445 -732
rect 1801 -733 1802 -732
rect 219 -735 220 -734
rect 1612 -735 1613 -734
rect 1619 -735 1620 -734
rect 1752 -735 1753 -734
rect 250 -737 251 -736
rect 1192 -737 1193 -736
rect 1206 -737 1207 -736
rect 1269 -737 1270 -736
rect 1353 -737 1354 -736
rect 1444 -737 1445 -736
rect 1472 -737 1473 -736
rect 1619 -737 1620 -736
rect 1633 -737 1634 -736
rect 1731 -737 1732 -736
rect 142 -739 143 -738
rect 1472 -739 1473 -738
rect 1500 -739 1501 -738
rect 1640 -739 1641 -738
rect 1654 -739 1655 -738
rect 1878 -739 1879 -738
rect 205 -741 206 -740
rect 1500 -741 1501 -740
rect 1514 -741 1515 -740
rect 1654 -741 1655 -740
rect 1668 -741 1669 -740
rect 2018 -741 2019 -740
rect 289 -743 290 -742
rect 499 -743 500 -742
rect 537 -743 538 -742
rect 989 -743 990 -742
rect 1024 -743 1025 -742
rect 1577 -743 1578 -742
rect 1696 -743 1697 -742
rect 1815 -743 1816 -742
rect 373 -745 374 -744
rect 1696 -745 1697 -744
rect 352 -747 353 -746
rect 373 -747 374 -746
rect 380 -747 381 -746
rect 576 -747 577 -746
rect 611 -747 612 -746
rect 688 -747 689 -746
rect 726 -747 727 -746
rect 1353 -747 1354 -746
rect 1370 -747 1371 -746
rect 1843 -747 1844 -746
rect 254 -749 255 -748
rect 380 -749 381 -748
rect 394 -749 395 -748
rect 534 -749 535 -748
rect 632 -749 633 -748
rect 660 -749 661 -748
rect 674 -749 675 -748
rect 709 -749 710 -748
rect 1017 -749 1018 -748
rect 1024 -749 1025 -748
rect 1038 -749 1039 -748
rect 1115 -749 1116 -748
rect 1185 -749 1186 -748
rect 1234 -749 1235 -748
rect 1241 -749 1242 -748
rect 1290 -749 1291 -748
rect 1374 -749 1375 -748
rect 1458 -749 1459 -748
rect 1514 -749 1515 -748
rect 1521 -749 1522 -748
rect 1535 -749 1536 -748
rect 1633 -749 1634 -748
rect 254 -751 255 -750
rect 520 -751 521 -750
rect 597 -751 598 -750
rect 674 -751 675 -750
rect 688 -751 689 -750
rect 1164 -751 1165 -750
rect 1185 -751 1186 -750
rect 1563 -751 1564 -750
rect 331 -753 332 -752
rect 352 -753 353 -752
rect 387 -753 388 -752
rect 597 -753 598 -752
rect 968 -753 969 -752
rect 1017 -753 1018 -752
rect 1094 -753 1095 -752
rect 1339 -753 1340 -752
rect 1346 -753 1347 -752
rect 1521 -753 1522 -752
rect 1535 -753 1536 -752
rect 1864 -753 1865 -752
rect 275 -755 276 -754
rect 331 -755 332 -754
rect 387 -755 388 -754
rect 478 -755 479 -754
rect 499 -755 500 -754
rect 513 -755 514 -754
rect 933 -755 934 -754
rect 968 -755 969 -754
rect 975 -755 976 -754
rect 1038 -755 1039 -754
rect 1139 -755 1140 -754
rect 1374 -755 1375 -754
rect 1381 -755 1382 -754
rect 1647 -755 1648 -754
rect 275 -757 276 -756
rect 296 -757 297 -756
rect 359 -757 360 -756
rect 478 -757 479 -756
rect 513 -757 514 -756
rect 919 -757 920 -756
rect 954 -757 955 -756
rect 975 -757 976 -756
rect 1153 -757 1154 -756
rect 1241 -757 1242 -756
rect 1283 -757 1284 -756
rect 1346 -757 1347 -756
rect 1395 -757 1396 -756
rect 1507 -757 1508 -756
rect 1538 -757 1539 -756
rect 1766 -757 1767 -756
rect 208 -759 209 -758
rect 919 -759 920 -758
rect 1157 -759 1158 -758
rect 1164 -759 1165 -758
rect 1206 -759 1207 -758
rect 1220 -759 1221 -758
rect 1311 -759 1312 -758
rect 1381 -759 1382 -758
rect 1395 -759 1396 -758
rect 1402 -759 1403 -758
rect 1542 -759 1543 -758
rect 1668 -759 1669 -758
rect 44 -761 45 -760
rect 1542 -761 1543 -760
rect 135 -763 136 -762
rect 208 -763 209 -762
rect 296 -763 297 -762
rect 541 -763 542 -762
rect 786 -763 787 -762
rect 954 -763 955 -762
rect 961 -763 962 -762
rect 1311 -763 1312 -762
rect 1318 -763 1319 -762
rect 1563 -763 1564 -762
rect 345 -765 346 -764
rect 359 -765 360 -764
rect 443 -765 444 -764
rect 527 -765 528 -764
rect 810 -765 811 -764
rect 1283 -765 1284 -764
rect 79 -767 80 -766
rect 527 -767 528 -766
rect 884 -767 885 -766
rect 933 -767 934 -766
rect 1157 -767 1158 -766
rect 2032 -767 2033 -766
rect 79 -769 80 -768
rect 632 -769 633 -768
rect 905 -769 906 -768
rect 961 -769 962 -768
rect 1209 -769 1210 -768
rect 2032 -769 2033 -768
rect 107 -771 108 -770
rect 884 -771 885 -770
rect 1220 -771 1221 -770
rect 2214 -771 2215 -770
rect 107 -773 108 -772
rect 821 -773 822 -772
rect 1262 -773 1263 -772
rect 1402 -773 1403 -772
rect 268 -775 269 -774
rect 905 -775 906 -774
rect 268 -777 269 -776
rect 338 -777 339 -776
rect 345 -777 346 -776
rect 649 -777 650 -776
rect 821 -777 822 -776
rect 835 -777 836 -776
rect 880 -777 881 -776
rect 1262 -777 1263 -776
rect 338 -779 339 -778
rect 751 -779 752 -778
rect 828 -779 829 -778
rect 835 -779 836 -778
rect 450 -781 451 -780
rect 730 -781 731 -780
rect 751 -781 752 -780
rect 1416 -781 1417 -780
rect 128 -783 129 -782
rect 1416 -783 1417 -782
rect 233 -785 234 -784
rect 450 -785 451 -784
rect 457 -785 458 -784
rect 541 -785 542 -784
rect 828 -785 829 -784
rect 1913 -785 1914 -784
rect 233 -787 234 -786
rect 394 -787 395 -786
rect 457 -787 458 -786
rect 842 -787 843 -786
rect 1787 -787 1788 -786
rect 1913 -787 1914 -786
rect 471 -789 472 -788
rect 646 -789 647 -788
rect 842 -789 843 -788
rect 912 -789 913 -788
rect 1661 -789 1662 -788
rect 1787 -789 1788 -788
rect 471 -791 472 -790
rect 1010 -791 1011 -790
rect 1276 -791 1277 -790
rect 1661 -791 1662 -790
rect 520 -793 521 -792
rect 1318 -793 1319 -792
rect 912 -795 913 -794
rect 1297 -795 1298 -794
rect 1276 -797 1277 -796
rect 1479 -797 1480 -796
rect 1297 -799 1298 -798
rect 1332 -799 1333 -798
rect 1388 -799 1389 -798
rect 1479 -799 1480 -798
rect 1325 -801 1326 -800
rect 1388 -801 1389 -800
rect 226 -803 227 -802
rect 1325 -803 1326 -802
rect 1332 -803 1333 -802
rect 1906 -803 1907 -802
rect 226 -805 227 -804
rect 586 -805 587 -804
rect 436 -807 437 -806
rect 586 -807 587 -806
rect 222 -809 223 -808
rect 436 -809 437 -808
rect 9 -820 10 -819
rect 1626 -820 1627 -819
rect 1661 -820 1662 -819
rect 2361 -820 2362 -819
rect 2403 -820 2404 -819
rect 2417 -820 2418 -819
rect 9 -822 10 -821
rect 93 -822 94 -821
rect 103 -822 104 -821
rect 352 -822 353 -821
rect 457 -822 458 -821
rect 590 -822 591 -821
rect 614 -822 615 -821
rect 653 -822 654 -821
rect 674 -822 675 -821
rect 747 -822 748 -821
rect 782 -822 783 -821
rect 849 -822 850 -821
rect 947 -822 948 -821
rect 1314 -822 1315 -821
rect 1332 -822 1333 -821
rect 1423 -822 1424 -821
rect 1538 -822 1539 -821
rect 2095 -822 2096 -821
rect 2326 -822 2327 -821
rect 2336 -822 2337 -821
rect 2343 -822 2344 -821
rect 2403 -822 2404 -821
rect 16 -824 17 -823
rect 191 -824 192 -823
rect 222 -824 223 -823
rect 2249 -824 2250 -823
rect 2277 -824 2278 -823
rect 2326 -824 2327 -823
rect 2347 -824 2348 -823
rect 2375 -824 2376 -823
rect 16 -826 17 -825
rect 1325 -826 1326 -825
rect 1335 -826 1336 -825
rect 1521 -826 1522 -825
rect 1598 -826 1599 -825
rect 1601 -826 1602 -825
rect 1626 -826 1627 -825
rect 1654 -826 1655 -825
rect 1661 -826 1662 -825
rect 1815 -826 1816 -825
rect 2095 -826 2096 -825
rect 2151 -826 2152 -825
rect 2277 -826 2278 -825
rect 2340 -826 2341 -825
rect 2347 -826 2348 -825
rect 2368 -826 2369 -825
rect 44 -828 45 -827
rect 1696 -828 1697 -827
rect 1815 -828 1816 -827
rect 1878 -828 1879 -827
rect 2151 -828 2152 -827
rect 2179 -828 2180 -827
rect 44 -830 45 -829
rect 940 -830 941 -829
rect 947 -830 948 -829
rect 968 -830 969 -829
rect 989 -830 990 -829
rect 1423 -830 1424 -829
rect 1598 -830 1599 -829
rect 1717 -830 1718 -829
rect 1878 -830 1879 -829
rect 1941 -830 1942 -829
rect 1990 -830 1991 -829
rect 2179 -830 2180 -829
rect 58 -832 59 -831
rect 754 -832 755 -831
rect 817 -832 818 -831
rect 1409 -832 1410 -831
rect 1601 -832 1602 -831
rect 1717 -832 1718 -831
rect 1899 -832 1900 -831
rect 1990 -832 1991 -831
rect 58 -834 59 -833
rect 135 -834 136 -833
rect 142 -834 143 -833
rect 222 -834 223 -833
rect 254 -834 255 -833
rect 590 -834 591 -833
rect 635 -834 636 -833
rect 926 -834 927 -833
rect 989 -834 990 -833
rect 1132 -834 1133 -833
rect 1136 -834 1137 -833
rect 1801 -834 1802 -833
rect 1941 -834 1942 -833
rect 1983 -834 1984 -833
rect 79 -836 80 -835
rect 261 -836 262 -835
rect 282 -836 283 -835
rect 362 -836 363 -835
rect 422 -836 423 -835
rect 849 -836 850 -835
rect 870 -836 871 -835
rect 940 -836 941 -835
rect 996 -836 997 -835
rect 1244 -836 1245 -835
rect 1248 -836 1249 -835
rect 1521 -836 1522 -835
rect 1605 -836 1606 -835
rect 1696 -836 1697 -835
rect 1983 -836 1984 -835
rect 2025 -836 2026 -835
rect 72 -838 73 -837
rect 996 -838 997 -837
rect 1020 -838 1021 -837
rect 1556 -838 1557 -837
rect 1573 -838 1574 -837
rect 2025 -838 2026 -837
rect 72 -840 73 -839
rect 667 -840 668 -839
rect 681 -840 682 -839
rect 716 -840 717 -839
rect 821 -840 822 -839
rect 870 -840 871 -839
rect 926 -840 927 -839
rect 1192 -840 1193 -839
rect 1195 -840 1196 -839
rect 2109 -840 2110 -839
rect 79 -842 80 -841
rect 324 -842 325 -841
rect 352 -842 353 -841
rect 499 -842 500 -841
rect 506 -842 507 -841
rect 723 -842 724 -841
rect 772 -842 773 -841
rect 821 -842 822 -841
rect 1010 -842 1011 -841
rect 2109 -842 2110 -841
rect 121 -844 122 -843
rect 268 -844 269 -843
rect 282 -844 283 -843
rect 1160 -844 1161 -843
rect 1174 -844 1175 -843
rect 1773 -844 1774 -843
rect 47 -846 48 -845
rect 1773 -846 1774 -845
rect 128 -848 129 -847
rect 562 -848 563 -847
rect 646 -848 647 -847
rect 831 -848 832 -847
rect 1010 -848 1011 -847
rect 1087 -848 1088 -847
rect 1094 -848 1095 -847
rect 1122 -848 1123 -847
rect 1129 -848 1130 -847
rect 2235 -848 2236 -847
rect 128 -850 129 -849
rect 1041 -850 1042 -849
rect 1045 -850 1046 -849
rect 1087 -850 1088 -849
rect 1094 -850 1095 -849
rect 1101 -850 1102 -849
rect 1111 -850 1112 -849
rect 2046 -850 2047 -849
rect 2235 -850 2236 -849
rect 2284 -850 2285 -849
rect 145 -852 146 -851
rect 800 -852 801 -851
rect 828 -852 829 -851
rect 1129 -852 1130 -851
rect 1136 -852 1137 -851
rect 1227 -852 1228 -851
rect 1248 -852 1249 -851
rect 1388 -852 1389 -851
rect 1402 -852 1403 -851
rect 1409 -852 1410 -851
rect 1430 -852 1431 -851
rect 2046 -852 2047 -851
rect 170 -854 171 -853
rect 191 -854 192 -853
rect 205 -854 206 -853
rect 1801 -854 1802 -853
rect 170 -856 171 -855
rect 271 -856 272 -855
rect 296 -856 297 -855
rect 583 -856 584 -855
rect 646 -856 647 -855
rect 1255 -856 1256 -855
rect 1272 -856 1273 -855
rect 1969 -856 1970 -855
rect 184 -858 185 -857
rect 289 -858 290 -857
rect 310 -858 311 -857
rect 376 -858 377 -857
rect 422 -858 423 -857
rect 1108 -858 1109 -857
rect 1139 -858 1140 -857
rect 1241 -858 1242 -857
rect 1255 -858 1256 -857
rect 1353 -858 1354 -857
rect 1360 -858 1361 -857
rect 2319 -858 2320 -857
rect 184 -860 185 -859
rect 758 -860 759 -859
rect 775 -860 776 -859
rect 1108 -860 1109 -859
rect 1143 -860 1144 -859
rect 2074 -860 2075 -859
rect 198 -862 199 -861
rect 289 -862 290 -861
rect 310 -862 311 -861
rect 450 -862 451 -861
rect 457 -862 458 -861
rect 548 -862 549 -861
rect 562 -862 563 -861
rect 569 -862 570 -861
rect 653 -862 654 -861
rect 1024 -862 1025 -861
rect 1045 -862 1046 -861
rect 1059 -862 1060 -861
rect 1101 -862 1102 -861
rect 1185 -862 1186 -861
rect 1206 -862 1207 -861
rect 1759 -862 1760 -861
rect 1969 -862 1970 -861
rect 2004 -862 2005 -861
rect 2074 -862 2075 -861
rect 2130 -862 2131 -861
rect 156 -864 157 -863
rect 198 -864 199 -863
rect 205 -864 206 -863
rect 233 -864 234 -863
rect 254 -864 255 -863
rect 520 -864 521 -863
rect 527 -864 528 -863
rect 1206 -864 1207 -863
rect 1209 -864 1210 -863
rect 2123 -864 2124 -863
rect 2130 -864 2131 -863
rect 2165 -864 2166 -863
rect 156 -866 157 -865
rect 443 -866 444 -865
rect 478 -866 479 -865
rect 520 -866 521 -865
rect 527 -866 528 -865
rect 807 -866 808 -865
rect 828 -866 829 -865
rect 1780 -866 1781 -865
rect 2004 -866 2005 -865
rect 2053 -866 2054 -865
rect 2123 -866 2124 -865
rect 2137 -866 2138 -865
rect 163 -868 164 -867
rect 450 -868 451 -867
rect 478 -868 479 -867
rect 772 -868 773 -867
rect 807 -868 808 -867
rect 1080 -868 1081 -867
rect 1143 -868 1144 -867
rect 1216 -868 1217 -867
rect 1220 -868 1221 -867
rect 2060 -868 2061 -867
rect 2102 -868 2103 -867
rect 2137 -868 2138 -867
rect 163 -870 164 -869
rect 331 -870 332 -869
rect 359 -870 360 -869
rect 569 -870 570 -869
rect 667 -870 668 -869
rect 2350 -870 2351 -869
rect 187 -872 188 -871
rect 1780 -872 1781 -871
rect 1787 -872 1788 -871
rect 2060 -872 2061 -871
rect 2102 -872 2103 -871
rect 2158 -872 2159 -871
rect 219 -874 220 -873
rect 800 -874 801 -873
rect 957 -874 958 -873
rect 1402 -874 1403 -873
rect 1556 -874 1557 -873
rect 1647 -874 1648 -873
rect 1654 -874 1655 -873
rect 1745 -874 1746 -873
rect 1787 -874 1788 -873
rect 1829 -874 1830 -873
rect 2053 -874 2054 -873
rect 2088 -874 2089 -873
rect 233 -876 234 -875
rect 303 -876 304 -875
rect 324 -876 325 -875
rect 373 -876 374 -875
rect 387 -876 388 -875
rect 443 -876 444 -875
rect 492 -876 493 -875
rect 968 -876 969 -875
rect 1024 -876 1025 -875
rect 1528 -876 1529 -875
rect 1605 -876 1606 -875
rect 1675 -876 1676 -875
rect 1682 -876 1683 -875
rect 1759 -876 1760 -875
rect 1829 -876 1830 -875
rect 1913 -876 1914 -875
rect 100 -878 101 -877
rect 387 -878 388 -877
rect 408 -878 409 -877
rect 548 -878 549 -877
rect 688 -878 689 -877
rect 726 -878 727 -877
rect 737 -878 738 -877
rect 758 -878 759 -877
rect 1055 -878 1056 -877
rect 2081 -878 2082 -877
rect 100 -880 101 -879
rect 936 -880 937 -879
rect 1080 -880 1081 -879
rect 1164 -880 1165 -879
rect 1185 -880 1186 -879
rect 1766 -880 1767 -879
rect 1871 -880 1872 -879
rect 2088 -880 2089 -879
rect 121 -882 122 -881
rect 373 -882 374 -881
rect 408 -882 409 -881
rect 415 -882 416 -881
rect 436 -882 437 -881
rect 506 -882 507 -881
rect 513 -882 514 -881
rect 719 -882 720 -881
rect 723 -882 724 -881
rect 1031 -882 1032 -881
rect 1146 -882 1147 -881
rect 1517 -882 1518 -881
rect 1647 -882 1648 -881
rect 1738 -882 1739 -881
rect 1745 -882 1746 -881
rect 1843 -882 1844 -881
rect 1913 -882 1914 -881
rect 1962 -882 1963 -881
rect 2081 -882 2082 -881
rect 2144 -882 2145 -881
rect 2 -884 3 -883
rect 415 -884 416 -883
rect 492 -884 493 -883
rect 765 -884 766 -883
rect 1031 -884 1032 -883
rect 1066 -884 1067 -883
rect 1157 -884 1158 -883
rect 2298 -884 2299 -883
rect 2 -886 3 -885
rect 177 -886 178 -885
rect 247 -886 248 -885
rect 303 -886 304 -885
rect 359 -886 360 -885
rect 380 -886 381 -885
rect 499 -886 500 -885
rect 530 -886 531 -885
rect 534 -886 535 -885
rect 583 -886 584 -885
rect 688 -886 689 -885
rect 709 -886 710 -885
rect 737 -886 738 -885
rect 884 -886 885 -885
rect 954 -886 955 -885
rect 2298 -886 2299 -885
rect 65 -888 66 -887
rect 1962 -888 1963 -887
rect 2144 -888 2145 -887
rect 2172 -888 2173 -887
rect 65 -890 66 -889
rect 394 -890 395 -889
rect 464 -890 465 -889
rect 534 -890 535 -889
rect 541 -890 542 -889
rect 674 -890 675 -889
rect 698 -890 699 -889
rect 919 -890 920 -889
rect 1052 -890 1053 -889
rect 1066 -890 1067 -889
rect 1157 -890 1158 -889
rect 1199 -890 1200 -889
rect 1213 -890 1214 -889
rect 2242 -890 2243 -889
rect 86 -892 87 -891
rect 394 -892 395 -891
rect 401 -892 402 -891
rect 464 -892 465 -891
rect 513 -892 514 -891
rect 597 -892 598 -891
rect 702 -892 703 -891
rect 1171 -892 1172 -891
rect 1199 -892 1200 -891
rect 1276 -892 1277 -891
rect 1286 -892 1287 -891
rect 1528 -892 1529 -891
rect 1682 -892 1683 -891
rect 1703 -892 1704 -891
rect 1738 -892 1739 -891
rect 1864 -892 1865 -891
rect 2172 -892 2173 -891
rect 2193 -892 2194 -891
rect 2207 -892 2208 -891
rect 2242 -892 2243 -891
rect 86 -894 87 -893
rect 366 -894 367 -893
rect 380 -894 381 -893
rect 611 -894 612 -893
rect 702 -894 703 -893
rect 835 -894 836 -893
rect 905 -894 906 -893
rect 1052 -894 1053 -893
rect 1125 -894 1126 -893
rect 1864 -894 1865 -893
rect 2193 -894 2194 -893
rect 2228 -894 2229 -893
rect 107 -896 108 -895
rect 905 -896 906 -895
rect 919 -896 920 -895
rect 1115 -896 1116 -895
rect 1164 -896 1165 -895
rect 1269 -896 1270 -895
rect 1290 -896 1291 -895
rect 1388 -896 1389 -895
rect 1395 -896 1396 -895
rect 1430 -896 1431 -895
rect 1766 -896 1767 -895
rect 2312 -896 2313 -895
rect 107 -898 108 -897
rect 240 -898 241 -897
rect 247 -898 248 -897
rect 1017 -898 1018 -897
rect 1038 -898 1039 -897
rect 1115 -898 1116 -897
rect 1171 -898 1172 -897
rect 2200 -898 2201 -897
rect 2207 -898 2208 -897
rect 2263 -898 2264 -897
rect 51 -900 52 -899
rect 240 -900 241 -899
rect 261 -900 262 -899
rect 632 -900 633 -899
rect 765 -900 766 -899
rect 814 -900 815 -899
rect 1192 -900 1193 -899
rect 1276 -900 1277 -899
rect 1290 -900 1291 -899
rect 1346 -900 1347 -899
rect 1353 -900 1354 -899
rect 1584 -900 1585 -899
rect 1794 -900 1795 -899
rect 1871 -900 1872 -899
rect 1892 -900 1893 -899
rect 2263 -900 2264 -899
rect 51 -902 52 -901
rect 628 -902 629 -901
rect 639 -902 640 -901
rect 1892 -902 1893 -901
rect 2018 -902 2019 -901
rect 2312 -902 2313 -901
rect 124 -904 125 -903
rect 1675 -904 1676 -903
rect 1794 -904 1795 -903
rect 1906 -904 1907 -903
rect 2018 -904 2019 -903
rect 2067 -904 2068 -903
rect 2186 -904 2187 -903
rect 2228 -904 2229 -903
rect 149 -906 150 -905
rect 436 -906 437 -905
rect 541 -906 542 -905
rect 611 -906 612 -905
rect 618 -906 619 -905
rect 632 -906 633 -905
rect 786 -906 787 -905
rect 835 -906 836 -905
rect 1213 -906 1214 -905
rect 1269 -906 1270 -905
rect 1304 -906 1305 -905
rect 2354 -906 2355 -905
rect 30 -908 31 -907
rect 786 -908 787 -907
rect 796 -908 797 -907
rect 884 -908 885 -907
rect 1220 -908 1221 -907
rect 1234 -908 1235 -907
rect 1241 -908 1242 -907
rect 1808 -908 1809 -907
rect 1843 -908 1844 -907
rect 2039 -908 2040 -907
rect 2067 -908 2068 -907
rect 2116 -908 2117 -907
rect 2200 -908 2201 -907
rect 2256 -908 2257 -907
rect 30 -910 31 -909
rect 177 -910 178 -909
rect 180 -910 181 -909
rect 709 -910 710 -909
rect 716 -910 717 -909
rect 1808 -910 1809 -909
rect 1906 -910 1907 -909
rect 1955 -910 1956 -909
rect 2039 -910 2040 -909
rect 2291 -910 2292 -909
rect 135 -912 136 -911
rect 2116 -912 2117 -911
rect 2214 -912 2215 -911
rect 2256 -912 2257 -911
rect 149 -914 150 -913
rect 1174 -914 1175 -913
rect 1223 -914 1224 -913
rect 1703 -914 1704 -913
rect 1955 -914 1956 -913
rect 1997 -914 1998 -913
rect 2214 -914 2215 -913
rect 2270 -914 2271 -913
rect 226 -916 227 -915
rect 639 -916 640 -915
rect 814 -916 815 -915
rect 1311 -916 1312 -915
rect 1325 -916 1326 -915
rect 1416 -916 1417 -915
rect 1535 -916 1536 -915
rect 2186 -916 2187 -915
rect 2270 -916 2271 -915
rect 2305 -916 2306 -915
rect 226 -918 227 -917
rect 877 -918 878 -917
rect 1178 -918 1179 -917
rect 1416 -918 1417 -917
rect 1493 -918 1494 -917
rect 2305 -918 2306 -917
rect 23 -920 24 -919
rect 877 -920 878 -919
rect 1122 -920 1123 -919
rect 1178 -920 1179 -919
rect 1227 -920 1228 -919
rect 1262 -920 1263 -919
rect 1304 -920 1305 -919
rect 1444 -920 1445 -919
rect 1493 -920 1494 -919
rect 1549 -920 1550 -919
rect 1584 -920 1585 -919
rect 1633 -920 1634 -919
rect 1997 -920 1998 -919
rect 2032 -920 2033 -919
rect 23 -922 24 -921
rect 114 -922 115 -921
rect 268 -922 269 -921
rect 2291 -922 2292 -921
rect 114 -924 115 -923
rect 485 -924 486 -923
rect 593 -924 594 -923
rect 954 -924 955 -923
rect 1234 -924 1235 -923
rect 1437 -924 1438 -923
rect 1535 -924 1536 -923
rect 1612 -924 1613 -923
rect 1633 -924 1634 -923
rect 1710 -924 1711 -923
rect 1857 -924 1858 -923
rect 2032 -924 2033 -923
rect 275 -926 276 -925
rect 296 -926 297 -925
rect 345 -926 346 -925
rect 618 -926 619 -925
rect 1262 -926 1263 -925
rect 1297 -926 1298 -925
rect 1311 -926 1312 -925
rect 2284 -926 2285 -925
rect 275 -928 276 -927
rect 429 -928 430 -927
rect 485 -928 486 -927
rect 555 -928 556 -927
rect 597 -928 598 -927
rect 604 -928 605 -927
rect 684 -928 685 -927
rect 1297 -928 1298 -927
rect 1339 -928 1340 -927
rect 1444 -928 1445 -927
rect 1549 -928 1550 -927
rect 1563 -928 1564 -927
rect 1612 -928 1613 -927
rect 1619 -928 1620 -927
rect 1710 -928 1711 -927
rect 1822 -928 1823 -927
rect 1857 -928 1858 -927
rect 1885 -928 1886 -927
rect 345 -930 346 -929
rect 660 -930 661 -929
rect 1283 -930 1284 -929
rect 1437 -930 1438 -929
rect 1563 -930 1564 -929
rect 1668 -930 1669 -929
rect 1822 -930 1823 -929
rect 1836 -930 1837 -929
rect 1885 -930 1886 -929
rect 1948 -930 1949 -929
rect 19 -932 20 -931
rect 1836 -932 1837 -931
rect 331 -934 332 -933
rect 1283 -934 1284 -933
rect 1339 -934 1340 -933
rect 1451 -934 1452 -933
rect 1500 -934 1501 -933
rect 1668 -934 1669 -933
rect 366 -936 367 -935
rect 1398 -936 1399 -935
rect 1500 -936 1501 -935
rect 1577 -936 1578 -935
rect 1619 -936 1620 -935
rect 1724 -936 1725 -935
rect 401 -938 402 -937
rect 695 -938 696 -937
rect 1059 -938 1060 -937
rect 1948 -938 1949 -937
rect 187 -940 188 -939
rect 695 -940 696 -939
rect 1318 -940 1319 -939
rect 1451 -940 1452 -939
rect 1577 -940 1578 -939
rect 1899 -940 1900 -939
rect 429 -942 430 -941
rect 1013 -942 1014 -941
rect 1318 -942 1319 -941
rect 1507 -942 1508 -941
rect 1724 -942 1725 -941
rect 1850 -942 1851 -941
rect 604 -944 605 -943
rect 842 -944 843 -943
rect 1346 -944 1347 -943
rect 1395 -944 1396 -943
rect 1507 -944 1508 -943
rect 1591 -944 1592 -943
rect 1850 -944 1851 -943
rect 1927 -944 1928 -943
rect 660 -946 661 -945
rect 912 -946 913 -945
rect 1360 -946 1361 -945
rect 1381 -946 1382 -945
rect 1591 -946 1592 -945
rect 1689 -946 1690 -945
rect 1927 -946 1928 -945
rect 1976 -946 1977 -945
rect 744 -948 745 -947
rect 1689 -948 1690 -947
rect 1976 -948 1977 -947
rect 2011 -948 2012 -947
rect 744 -950 745 -949
rect 793 -950 794 -949
rect 842 -950 843 -949
rect 933 -950 934 -949
rect 1363 -950 1364 -949
rect 2158 -950 2159 -949
rect 555 -952 556 -951
rect 933 -952 934 -951
rect 1367 -952 1368 -951
rect 1752 -952 1753 -951
rect 1920 -952 1921 -951
rect 2011 -952 2012 -951
rect 793 -954 794 -953
rect 961 -954 962 -953
rect 1017 -954 1018 -953
rect 1752 -954 1753 -953
rect 856 -956 857 -955
rect 912 -956 913 -955
rect 961 -956 962 -955
rect 982 -956 983 -955
rect 1367 -956 1368 -955
rect 1458 -956 1459 -955
rect 856 -958 857 -957
rect 891 -958 892 -957
rect 982 -958 983 -957
rect 1003 -958 1004 -957
rect 1370 -958 1371 -957
rect 2165 -958 2166 -957
rect 471 -960 472 -959
rect 891 -960 892 -959
rect 1374 -960 1375 -959
rect 1920 -960 1921 -959
rect 471 -962 472 -961
rect 576 -962 577 -961
rect 586 -962 587 -961
rect 1003 -962 1004 -961
rect 1374 -962 1375 -961
rect 1479 -962 1480 -961
rect 576 -964 577 -963
rect 625 -964 626 -963
rect 1381 -964 1382 -963
rect 1486 -964 1487 -963
rect 625 -966 626 -965
rect 2319 -966 2320 -965
rect 1458 -968 1459 -967
rect 1542 -968 1543 -967
rect 1479 -970 1480 -969
rect 1570 -970 1571 -969
rect 1486 -972 1487 -971
rect 1731 -972 1732 -971
rect 1465 -974 1466 -973
rect 1731 -974 1732 -973
rect 1465 -976 1466 -975
rect 1472 -976 1473 -975
rect 1542 -976 1543 -975
rect 1640 -976 1641 -975
rect 1073 -978 1074 -977
rect 1472 -978 1473 -977
rect 1514 -978 1515 -977
rect 1640 -978 1641 -977
rect 779 -980 780 -979
rect 1073 -980 1074 -979
rect 1514 -980 1515 -979
rect 2249 -980 2250 -979
rect 1570 -982 1571 -981
rect 2221 -982 2222 -981
rect 751 -984 752 -983
rect 2221 -984 2222 -983
rect 37 -986 38 -985
rect 751 -986 752 -985
rect 37 -988 38 -987
rect 975 -988 976 -987
rect 975 -990 976 -989
rect 1150 -990 1151 -989
rect 730 -992 731 -991
rect 1150 -992 1151 -991
rect 730 -994 731 -993
rect 863 -994 864 -993
rect 338 -996 339 -995
rect 863 -996 864 -995
rect 338 -998 339 -997
rect 390 -998 391 -997
rect 9 -1009 10 -1008
rect 761 -1009 762 -1008
rect 772 -1009 773 -1008
rect 2137 -1009 2138 -1008
rect 2284 -1009 2285 -1008
rect 2340 -1009 2341 -1008
rect 2375 -1009 2376 -1008
rect 2431 -1009 2432 -1008
rect 9 -1011 10 -1010
rect 58 -1011 59 -1010
rect 93 -1011 94 -1010
rect 2256 -1011 2257 -1010
rect 2298 -1011 2299 -1010
rect 2375 -1011 2376 -1010
rect 2382 -1011 2383 -1010
rect 2392 -1011 2393 -1010
rect 2403 -1011 2404 -1010
rect 2438 -1011 2439 -1010
rect 16 -1013 17 -1012
rect 58 -1013 59 -1012
rect 93 -1013 94 -1012
rect 842 -1013 843 -1012
rect 884 -1013 885 -1012
rect 933 -1013 934 -1012
rect 936 -1013 937 -1012
rect 1388 -1013 1389 -1012
rect 1507 -1013 1508 -1012
rect 1577 -1013 1578 -1012
rect 1703 -1013 1704 -1012
rect 2298 -1013 2299 -1012
rect 2368 -1013 2369 -1012
rect 2403 -1013 2404 -1012
rect 2417 -1013 2418 -1012
rect 2424 -1013 2425 -1012
rect 16 -1015 17 -1014
rect 331 -1015 332 -1014
rect 345 -1015 346 -1014
rect 1006 -1015 1007 -1014
rect 1020 -1015 1021 -1014
rect 2228 -1015 2229 -1014
rect 103 -1017 104 -1016
rect 1150 -1017 1151 -1016
rect 1174 -1017 1175 -1016
rect 1871 -1017 1872 -1016
rect 2123 -1017 2124 -1016
rect 2368 -1017 2369 -1016
rect 110 -1019 111 -1018
rect 317 -1019 318 -1018
rect 324 -1019 325 -1018
rect 331 -1019 332 -1018
rect 345 -1019 346 -1018
rect 443 -1019 444 -1018
rect 590 -1019 591 -1018
rect 628 -1019 629 -1018
rect 646 -1019 647 -1018
rect 954 -1019 955 -1018
rect 964 -1019 965 -1018
rect 2242 -1019 2243 -1018
rect 117 -1021 118 -1020
rect 1451 -1021 1452 -1020
rect 1514 -1021 1515 -1020
rect 1682 -1021 1683 -1020
rect 1689 -1021 1690 -1020
rect 1703 -1021 1704 -1020
rect 1787 -1021 1788 -1020
rect 2123 -1021 2124 -1020
rect 2165 -1021 2166 -1020
rect 2228 -1021 2229 -1020
rect 128 -1023 129 -1022
rect 782 -1023 783 -1022
rect 793 -1023 794 -1022
rect 1108 -1023 1109 -1022
rect 1122 -1023 1123 -1022
rect 1360 -1023 1361 -1022
rect 1514 -1023 1515 -1022
rect 1535 -1023 1536 -1022
rect 1710 -1023 1711 -1022
rect 1787 -1023 1788 -1022
rect 1801 -1023 1802 -1022
rect 2389 -1023 2390 -1022
rect 128 -1025 129 -1024
rect 261 -1025 262 -1024
rect 268 -1025 269 -1024
rect 478 -1025 479 -1024
rect 590 -1025 591 -1024
rect 667 -1025 668 -1024
rect 733 -1025 734 -1024
rect 2291 -1025 2292 -1024
rect 86 -1027 87 -1026
rect 667 -1027 668 -1026
rect 779 -1027 780 -1026
rect 1990 -1027 1991 -1026
rect 2102 -1027 2103 -1026
rect 2291 -1027 2292 -1026
rect 86 -1029 87 -1028
rect 135 -1029 136 -1028
rect 138 -1029 139 -1028
rect 1892 -1029 1893 -1028
rect 1962 -1029 1963 -1028
rect 1990 -1029 1991 -1028
rect 2172 -1029 2173 -1028
rect 2242 -1029 2243 -1028
rect 135 -1031 136 -1030
rect 1822 -1031 1823 -1030
rect 1836 -1031 1837 -1030
rect 1892 -1031 1893 -1030
rect 1962 -1031 1963 -1030
rect 2018 -1031 2019 -1030
rect 2130 -1031 2131 -1030
rect 2172 -1031 2173 -1030
rect 177 -1033 178 -1032
rect 2319 -1033 2320 -1032
rect 23 -1035 24 -1034
rect 177 -1035 178 -1034
rect 180 -1035 181 -1034
rect 464 -1035 465 -1034
rect 478 -1035 479 -1034
rect 485 -1035 486 -1034
rect 611 -1035 612 -1034
rect 2221 -1035 2222 -1034
rect 23 -1037 24 -1036
rect 44 -1037 45 -1036
rect 100 -1037 101 -1036
rect 2319 -1037 2320 -1036
rect 44 -1039 45 -1038
rect 240 -1039 241 -1038
rect 261 -1039 262 -1038
rect 275 -1039 276 -1038
rect 310 -1039 311 -1038
rect 880 -1039 881 -1038
rect 940 -1039 941 -1038
rect 1017 -1039 1018 -1038
rect 1024 -1039 1025 -1038
rect 1507 -1039 1508 -1038
rect 1517 -1039 1518 -1038
rect 2263 -1039 2264 -1038
rect 184 -1041 185 -1040
rect 254 -1041 255 -1040
rect 271 -1041 272 -1040
rect 779 -1041 780 -1040
rect 793 -1041 794 -1040
rect 856 -1041 857 -1040
rect 863 -1041 864 -1040
rect 884 -1041 885 -1040
rect 891 -1041 892 -1040
rect 940 -1041 941 -1040
rect 975 -1041 976 -1040
rect 1108 -1041 1109 -1040
rect 1125 -1041 1126 -1040
rect 2088 -1041 2089 -1040
rect 2158 -1041 2159 -1040
rect 2221 -1041 2222 -1040
rect 138 -1043 139 -1042
rect 2158 -1043 2159 -1042
rect 187 -1045 188 -1044
rect 2277 -1045 2278 -1044
rect 191 -1047 192 -1046
rect 310 -1047 311 -1046
rect 324 -1047 325 -1046
rect 681 -1047 682 -1046
rect 723 -1047 724 -1046
rect 975 -1047 976 -1046
rect 989 -1047 990 -1046
rect 1038 -1047 1039 -1046
rect 1041 -1047 1042 -1046
rect 2018 -1047 2019 -1046
rect 2067 -1047 2068 -1046
rect 2130 -1047 2131 -1046
rect 2200 -1047 2201 -1046
rect 2277 -1047 2278 -1046
rect 170 -1049 171 -1048
rect 191 -1049 192 -1048
rect 205 -1049 206 -1048
rect 317 -1049 318 -1048
rect 366 -1049 367 -1048
rect 611 -1049 612 -1048
rect 625 -1049 626 -1048
rect 1731 -1049 1732 -1048
rect 1738 -1049 1739 -1048
rect 1822 -1049 1823 -1048
rect 1843 -1049 1844 -1048
rect 2102 -1049 2103 -1048
rect 2200 -1049 2201 -1048
rect 2249 -1049 2250 -1048
rect 121 -1051 122 -1050
rect 205 -1051 206 -1050
rect 219 -1051 220 -1050
rect 653 -1051 654 -1050
rect 660 -1051 661 -1050
rect 716 -1051 717 -1050
rect 730 -1051 731 -1050
rect 856 -1051 857 -1050
rect 863 -1051 864 -1050
rect 1689 -1051 1690 -1050
rect 1710 -1051 1711 -1050
rect 2361 -1051 2362 -1050
rect 121 -1053 122 -1052
rect 359 -1053 360 -1052
rect 366 -1053 367 -1052
rect 1171 -1053 1172 -1052
rect 1181 -1053 1182 -1052
rect 1626 -1053 1627 -1052
rect 1745 -1053 1746 -1052
rect 1801 -1053 1802 -1052
rect 1843 -1053 1844 -1052
rect 1850 -1053 1851 -1052
rect 1864 -1053 1865 -1052
rect 2137 -1053 2138 -1052
rect 2186 -1053 2187 -1052
rect 2249 -1053 2250 -1052
rect 145 -1055 146 -1054
rect 730 -1055 731 -1054
rect 796 -1055 797 -1054
rect 912 -1055 913 -1054
rect 996 -1055 997 -1054
rect 1202 -1055 1203 -1054
rect 1234 -1055 1235 -1054
rect 1388 -1055 1389 -1054
rect 1437 -1055 1438 -1054
rect 1731 -1055 1732 -1054
rect 1815 -1055 1816 -1054
rect 1850 -1055 1851 -1054
rect 1871 -1055 1872 -1054
rect 1906 -1055 1907 -1054
rect 1983 -1055 1984 -1054
rect 2263 -1055 2264 -1054
rect 170 -1057 171 -1056
rect 376 -1057 377 -1056
rect 380 -1057 381 -1056
rect 775 -1057 776 -1056
rect 817 -1057 818 -1056
rect 1668 -1057 1669 -1056
rect 1675 -1057 1676 -1056
rect 1906 -1057 1907 -1056
rect 1955 -1057 1956 -1056
rect 1983 -1057 1984 -1056
rect 2004 -1057 2005 -1056
rect 2067 -1057 2068 -1056
rect 2186 -1057 2187 -1056
rect 2399 -1057 2400 -1056
rect 79 -1059 80 -1058
rect 380 -1059 381 -1058
rect 387 -1059 388 -1058
rect 814 -1059 815 -1058
rect 831 -1059 832 -1058
rect 2032 -1059 2033 -1058
rect 2039 -1059 2040 -1058
rect 2361 -1059 2362 -1058
rect 79 -1061 80 -1060
rect 114 -1061 115 -1060
rect 222 -1061 223 -1060
rect 618 -1061 619 -1060
rect 639 -1061 640 -1060
rect 723 -1061 724 -1060
rect 775 -1061 776 -1060
rect 968 -1061 969 -1060
rect 982 -1061 983 -1060
rect 996 -1061 997 -1060
rect 1003 -1061 1004 -1060
rect 1171 -1061 1172 -1060
rect 1192 -1061 1193 -1060
rect 2046 -1061 2047 -1060
rect 30 -1063 31 -1062
rect 618 -1063 619 -1062
rect 646 -1063 647 -1062
rect 709 -1063 710 -1062
rect 835 -1063 836 -1062
rect 1122 -1063 1123 -1062
rect 1136 -1063 1137 -1062
rect 1150 -1063 1151 -1062
rect 1157 -1063 1158 -1062
rect 1192 -1063 1193 -1062
rect 1234 -1063 1235 -1062
rect 1836 -1063 1837 -1062
rect 1878 -1063 1879 -1062
rect 2165 -1063 2166 -1062
rect 30 -1065 31 -1064
rect 719 -1065 720 -1064
rect 835 -1065 836 -1064
rect 947 -1065 948 -1064
rect 968 -1065 969 -1064
rect 1073 -1065 1074 -1064
rect 1129 -1065 1130 -1064
rect 1157 -1065 1158 -1064
rect 1237 -1065 1238 -1064
rect 1290 -1065 1291 -1064
rect 1307 -1065 1308 -1064
rect 2004 -1065 2005 -1064
rect 2011 -1065 2012 -1064
rect 2088 -1065 2089 -1064
rect 65 -1067 66 -1066
rect 639 -1067 640 -1066
rect 660 -1067 661 -1066
rect 758 -1067 759 -1066
rect 842 -1067 843 -1066
rect 870 -1067 871 -1066
rect 877 -1067 878 -1066
rect 912 -1067 913 -1066
rect 947 -1067 948 -1066
rect 2256 -1067 2257 -1066
rect 65 -1069 66 -1068
rect 471 -1069 472 -1068
rect 485 -1069 486 -1068
rect 534 -1069 535 -1068
rect 597 -1069 598 -1068
rect 625 -1069 626 -1068
rect 635 -1069 636 -1068
rect 1073 -1069 1074 -1068
rect 1087 -1069 1088 -1068
rect 1129 -1069 1130 -1068
rect 1136 -1069 1137 -1068
rect 1472 -1069 1473 -1068
rect 1479 -1069 1480 -1068
rect 1535 -1069 1536 -1068
rect 1542 -1069 1543 -1068
rect 1626 -1069 1627 -1068
rect 1633 -1069 1634 -1068
rect 1675 -1069 1676 -1068
rect 1815 -1069 1816 -1068
rect 2396 -1069 2397 -1068
rect 226 -1071 227 -1070
rect 464 -1071 465 -1070
rect 513 -1071 514 -1070
rect 814 -1071 815 -1070
rect 891 -1071 892 -1070
rect 898 -1071 899 -1070
rect 1003 -1071 1004 -1070
rect 1024 -1071 1025 -1070
rect 1045 -1071 1046 -1070
rect 1087 -1071 1088 -1070
rect 1241 -1071 1242 -1070
rect 2060 -1071 2061 -1070
rect 51 -1073 52 -1072
rect 513 -1073 514 -1072
rect 534 -1073 535 -1072
rect 1269 -1073 1270 -1072
rect 1272 -1073 1273 -1072
rect 2032 -1073 2033 -1072
rect 2039 -1073 2040 -1072
rect 2347 -1073 2348 -1072
rect 51 -1075 52 -1074
rect 142 -1075 143 -1074
rect 212 -1075 213 -1074
rect 226 -1075 227 -1074
rect 240 -1075 241 -1074
rect 527 -1075 528 -1074
rect 597 -1075 598 -1074
rect 1062 -1075 1063 -1074
rect 1223 -1075 1224 -1074
rect 1241 -1075 1242 -1074
rect 1244 -1075 1245 -1074
rect 2284 -1075 2285 -1074
rect 142 -1077 143 -1076
rect 989 -1077 990 -1076
rect 1010 -1077 1011 -1076
rect 1038 -1077 1039 -1076
rect 1055 -1077 1056 -1076
rect 1549 -1077 1550 -1076
rect 1598 -1077 1599 -1076
rect 1668 -1077 1669 -1076
rect 1829 -1077 1830 -1076
rect 1864 -1077 1865 -1076
rect 1878 -1077 1879 -1076
rect 1927 -1077 1928 -1076
rect 1941 -1077 1942 -1076
rect 1955 -1077 1956 -1076
rect 1969 -1077 1970 -1076
rect 2011 -1077 2012 -1076
rect 2207 -1077 2208 -1076
rect 2347 -1077 2348 -1076
rect 198 -1079 199 -1078
rect 212 -1079 213 -1078
rect 254 -1079 255 -1078
rect 541 -1079 542 -1078
rect 681 -1079 682 -1078
rect 950 -1079 951 -1078
rect 1017 -1079 1018 -1078
rect 1115 -1079 1116 -1078
rect 1248 -1079 1249 -1078
rect 1360 -1079 1361 -1078
rect 1374 -1079 1375 -1078
rect 1437 -1079 1438 -1078
rect 1486 -1079 1487 -1078
rect 1829 -1079 1830 -1078
rect 1927 -1079 1928 -1078
rect 2193 -1079 2194 -1078
rect 198 -1081 199 -1080
rect 807 -1081 808 -1080
rect 877 -1081 878 -1080
rect 1269 -1081 1270 -1080
rect 1283 -1081 1284 -1080
rect 2312 -1081 2313 -1080
rect 275 -1083 276 -1082
rect 415 -1083 416 -1082
rect 429 -1083 430 -1082
rect 1447 -1083 1448 -1082
rect 1500 -1083 1501 -1082
rect 1542 -1083 1543 -1082
rect 1580 -1083 1581 -1082
rect 1941 -1083 1942 -1082
rect 1997 -1083 1998 -1082
rect 2046 -1083 2047 -1082
rect 2109 -1083 2110 -1082
rect 2207 -1083 2208 -1082
rect 2235 -1083 2236 -1082
rect 2312 -1083 2313 -1082
rect 359 -1085 360 -1084
rect 432 -1085 433 -1084
rect 443 -1085 444 -1084
rect 499 -1085 500 -1084
rect 541 -1085 542 -1084
rect 604 -1085 605 -1084
rect 607 -1085 608 -1084
rect 2193 -1085 2194 -1084
rect 114 -1087 115 -1086
rect 499 -1087 500 -1086
rect 604 -1087 605 -1086
rect 1045 -1087 1046 -1086
rect 1059 -1087 1060 -1086
rect 1143 -1087 1144 -1086
rect 1227 -1087 1228 -1086
rect 1248 -1087 1249 -1086
rect 1286 -1087 1287 -1086
rect 1759 -1087 1760 -1086
rect 1808 -1087 1809 -1086
rect 1969 -1087 1970 -1086
rect 2151 -1087 2152 -1086
rect 2235 -1087 2236 -1086
rect 401 -1089 402 -1088
rect 404 -1089 405 -1088
rect 415 -1089 416 -1088
rect 506 -1089 507 -1088
rect 695 -1089 696 -1088
rect 982 -1089 983 -1088
rect 1080 -1089 1081 -1088
rect 1143 -1089 1144 -1088
rect 1213 -1089 1214 -1088
rect 1227 -1089 1228 -1088
rect 1314 -1089 1315 -1088
rect 1640 -1089 1641 -1088
rect 1654 -1089 1655 -1088
rect 1745 -1089 1746 -1088
rect 1857 -1089 1858 -1088
rect 2109 -1089 2110 -1088
rect 401 -1091 402 -1090
rect 408 -1091 409 -1090
rect 429 -1091 430 -1090
rect 1773 -1091 1774 -1090
rect 1794 -1091 1795 -1090
rect 1857 -1091 1858 -1090
rect 2095 -1091 2096 -1090
rect 2151 -1091 2152 -1090
rect 408 -1093 409 -1092
rect 576 -1093 577 -1092
rect 688 -1093 689 -1092
rect 695 -1093 696 -1092
rect 702 -1093 703 -1092
rect 807 -1093 808 -1092
rect 898 -1093 899 -1092
rect 1094 -1093 1095 -1092
rect 1101 -1093 1102 -1092
rect 1115 -1093 1116 -1092
rect 1213 -1093 1214 -1092
rect 2343 -1093 2344 -1092
rect 2 -1095 3 -1094
rect 688 -1095 689 -1094
rect 709 -1095 710 -1094
rect 926 -1095 927 -1094
rect 1031 -1095 1032 -1094
rect 1101 -1095 1102 -1094
rect 1318 -1095 1319 -1094
rect 1451 -1095 1452 -1094
rect 1556 -1095 1557 -1094
rect 1640 -1095 1641 -1094
rect 1696 -1095 1697 -1094
rect 1759 -1095 1760 -1094
rect 2025 -1095 2026 -1094
rect 2095 -1095 2096 -1094
rect 72 -1097 73 -1096
rect 702 -1097 703 -1096
rect 737 -1097 738 -1096
rect 1290 -1097 1291 -1096
rect 1325 -1097 1326 -1096
rect 1374 -1097 1375 -1096
rect 1381 -1097 1382 -1096
rect 1472 -1097 1473 -1096
rect 1598 -1097 1599 -1096
rect 1605 -1097 1606 -1096
rect 1717 -1097 1718 -1096
rect 1773 -1097 1774 -1096
rect 1899 -1097 1900 -1096
rect 2025 -1097 2026 -1096
rect 37 -1099 38 -1098
rect 72 -1099 73 -1098
rect 89 -1099 90 -1098
rect 1094 -1099 1095 -1098
rect 1185 -1099 1186 -1098
rect 1696 -1099 1697 -1098
rect 1717 -1099 1718 -1098
rect 1752 -1099 1753 -1098
rect 1899 -1099 1900 -1098
rect 2333 -1099 2334 -1098
rect 37 -1101 38 -1100
rect 593 -1101 594 -1100
rect 751 -1101 752 -1100
rect 870 -1101 871 -1100
rect 905 -1101 906 -1100
rect 1031 -1101 1032 -1100
rect 1066 -1101 1067 -1100
rect 1080 -1101 1081 -1100
rect 1185 -1101 1186 -1100
rect 1199 -1101 1200 -1100
rect 1206 -1101 1207 -1100
rect 1318 -1101 1319 -1100
rect 1335 -1101 1336 -1100
rect 2305 -1101 2306 -1100
rect 247 -1103 248 -1102
rect 926 -1103 927 -1102
rect 961 -1103 962 -1102
rect 1066 -1103 1067 -1102
rect 1178 -1103 1179 -1102
rect 1206 -1103 1207 -1102
rect 1255 -1103 1256 -1102
rect 1325 -1103 1326 -1102
rect 1367 -1103 1368 -1102
rect 1381 -1103 1382 -1102
rect 1395 -1103 1396 -1102
rect 1752 -1103 1753 -1102
rect 2214 -1103 2215 -1102
rect 2305 -1103 2306 -1102
rect 163 -1105 164 -1104
rect 247 -1105 248 -1104
rect 373 -1105 374 -1104
rect 1178 -1105 1179 -1104
rect 1195 -1105 1196 -1104
rect 1556 -1105 1557 -1104
rect 1724 -1105 1725 -1104
rect 1808 -1105 1809 -1104
rect 2116 -1105 2117 -1104
rect 2214 -1105 2215 -1104
rect 2270 -1105 2271 -1104
rect 2333 -1105 2334 -1104
rect 163 -1107 164 -1106
rect 338 -1107 339 -1106
rect 352 -1107 353 -1106
rect 373 -1107 374 -1106
rect 390 -1107 391 -1106
rect 737 -1107 738 -1106
rect 772 -1107 773 -1106
rect 1633 -1107 1634 -1106
rect 2053 -1107 2054 -1106
rect 2116 -1107 2117 -1106
rect 233 -1109 234 -1108
rect 961 -1109 962 -1108
rect 1052 -1109 1053 -1108
rect 1724 -1109 1725 -1108
rect 2053 -1109 2054 -1108
rect 2336 -1109 2337 -1108
rect 233 -1111 234 -1110
rect 394 -1111 395 -1110
rect 450 -1111 451 -1110
rect 471 -1111 472 -1110
rect 506 -1111 507 -1110
rect 1794 -1111 1795 -1110
rect 107 -1113 108 -1112
rect 394 -1113 395 -1112
rect 450 -1113 451 -1112
rect 492 -1113 493 -1112
rect 548 -1113 549 -1112
rect 576 -1113 577 -1112
rect 674 -1113 675 -1112
rect 751 -1113 752 -1112
rect 786 -1113 787 -1112
rect 1010 -1113 1011 -1112
rect 1199 -1113 1200 -1112
rect 1766 -1113 1767 -1112
rect 107 -1115 108 -1114
rect 2326 -1115 2327 -1114
rect 338 -1117 339 -1116
rect 520 -1117 521 -1116
rect 569 -1117 570 -1116
rect 1052 -1117 1053 -1116
rect 1220 -1117 1221 -1116
rect 1255 -1117 1256 -1116
rect 1262 -1117 1263 -1116
rect 1367 -1117 1368 -1116
rect 1402 -1117 1403 -1116
rect 2060 -1117 2061 -1116
rect 352 -1119 353 -1118
rect 866 -1119 867 -1118
rect 905 -1119 906 -1118
rect 1682 -1119 1683 -1118
rect 1766 -1119 1767 -1118
rect 1780 -1119 1781 -1118
rect 422 -1121 423 -1120
rect 569 -1121 570 -1120
rect 674 -1121 675 -1120
rect 1167 -1121 1168 -1120
rect 1220 -1121 1221 -1120
rect 2270 -1121 2271 -1120
rect 100 -1123 101 -1122
rect 422 -1123 423 -1122
rect 436 -1123 437 -1122
rect 492 -1123 493 -1122
rect 520 -1123 521 -1122
rect 583 -1123 584 -1122
rect 744 -1123 745 -1122
rect 786 -1123 787 -1122
rect 800 -1123 801 -1122
rect 1283 -1123 1284 -1122
rect 1297 -1123 1298 -1122
rect 1395 -1123 1396 -1122
rect 1423 -1123 1424 -1122
rect 1479 -1123 1480 -1122
rect 1549 -1123 1550 -1122
rect 1605 -1123 1606 -1122
rect 1661 -1123 1662 -1122
rect 1780 -1123 1781 -1122
rect 289 -1125 290 -1124
rect 583 -1125 584 -1124
rect 800 -1125 801 -1124
rect 821 -1125 822 -1124
rect 1164 -1125 1165 -1124
rect 1262 -1125 1263 -1124
rect 1297 -1125 1298 -1124
rect 2354 -1125 2355 -1124
rect 289 -1127 290 -1126
rect 296 -1127 297 -1126
rect 436 -1127 437 -1126
rect 656 -1127 657 -1126
rect 821 -1127 822 -1126
rect 1997 -1127 1998 -1126
rect 296 -1129 297 -1128
rect 303 -1129 304 -1128
rect 457 -1129 458 -1128
rect 548 -1129 549 -1128
rect 555 -1129 556 -1128
rect 744 -1129 745 -1128
rect 1164 -1129 1165 -1128
rect 1612 -1129 1613 -1128
rect 1619 -1129 1620 -1128
rect 1661 -1129 1662 -1128
rect 282 -1131 283 -1130
rect 303 -1131 304 -1130
rect 404 -1131 405 -1130
rect 457 -1131 458 -1130
rect 555 -1131 556 -1130
rect 562 -1131 563 -1130
rect 1304 -1131 1305 -1130
rect 1402 -1131 1403 -1130
rect 1416 -1131 1417 -1130
rect 1423 -1131 1424 -1130
rect 1430 -1131 1431 -1130
rect 1486 -1131 1487 -1130
rect 1584 -1131 1585 -1130
rect 1612 -1131 1613 -1130
rect 149 -1133 150 -1132
rect 282 -1133 283 -1132
rect 1304 -1133 1305 -1132
rect 1934 -1133 1935 -1132
rect 149 -1135 150 -1134
rect 425 -1135 426 -1134
rect 1311 -1135 1312 -1134
rect 2326 -1135 2327 -1134
rect 156 -1137 157 -1136
rect 562 -1137 563 -1136
rect 1311 -1137 1312 -1136
rect 1339 -1137 1340 -1136
rect 1398 -1137 1399 -1136
rect 2354 -1137 2355 -1136
rect 96 -1139 97 -1138
rect 156 -1139 157 -1138
rect 824 -1139 825 -1138
rect 1339 -1139 1340 -1138
rect 1430 -1139 1431 -1138
rect 1521 -1139 1522 -1138
rect 1528 -1139 1529 -1138
rect 1584 -1139 1585 -1138
rect 1591 -1139 1592 -1138
rect 1619 -1139 1620 -1138
rect 1934 -1139 1935 -1138
rect 2081 -1139 2082 -1138
rect 632 -1141 633 -1140
rect 1591 -1141 1592 -1140
rect 2081 -1141 2082 -1140
rect 2179 -1141 2180 -1140
rect 632 -1143 633 -1142
rect 1160 -1143 1161 -1142
rect 1444 -1143 1445 -1142
rect 1500 -1143 1501 -1142
rect 2144 -1143 2145 -1142
rect 2179 -1143 2180 -1142
rect 1458 -1145 1459 -1144
rect 1521 -1145 1522 -1144
rect 2074 -1145 2075 -1144
rect 2144 -1145 2145 -1144
rect 1276 -1147 1277 -1146
rect 1458 -1147 1459 -1146
rect 1493 -1147 1494 -1146
rect 1528 -1147 1529 -1146
rect 1976 -1147 1977 -1146
rect 2074 -1147 2075 -1146
rect 828 -1149 829 -1148
rect 1276 -1149 1277 -1148
rect 1465 -1149 1466 -1148
rect 1493 -1149 1494 -1148
rect 1948 -1149 1949 -1148
rect 1976 -1149 1977 -1148
rect 765 -1151 766 -1150
rect 828 -1151 829 -1150
rect 1465 -1151 1466 -1150
rect 1647 -1151 1648 -1150
rect 1920 -1151 1921 -1150
rect 1948 -1151 1949 -1150
rect 765 -1153 766 -1152
rect 849 -1153 850 -1152
rect 1563 -1153 1564 -1152
rect 1647 -1153 1648 -1152
rect 1913 -1153 1914 -1152
rect 1920 -1153 1921 -1152
rect 849 -1155 850 -1154
rect 1416 -1155 1417 -1154
rect 1885 -1155 1886 -1154
rect 1913 -1155 1914 -1154
rect 1353 -1157 1354 -1156
rect 1563 -1157 1564 -1156
rect 1741 -1157 1742 -1156
rect 1885 -1157 1886 -1156
rect 1346 -1159 1347 -1158
rect 1353 -1159 1354 -1158
rect 1332 -1161 1333 -1160
rect 1346 -1161 1347 -1160
rect 957 -1163 958 -1162
rect 1332 -1163 1333 -1162
rect 957 -1165 958 -1164
rect 1654 -1165 1655 -1164
rect 5 -1176 6 -1175
rect 432 -1176 433 -1175
rect 485 -1176 486 -1175
rect 653 -1176 654 -1175
rect 656 -1176 657 -1175
rect 1514 -1176 1515 -1175
rect 1549 -1176 1550 -1175
rect 2291 -1176 2292 -1175
rect 2298 -1176 2299 -1175
rect 2494 -1176 2495 -1175
rect 19 -1178 20 -1177
rect 30 -1178 31 -1177
rect 89 -1178 90 -1177
rect 856 -1178 857 -1177
rect 866 -1178 867 -1177
rect 1031 -1178 1032 -1177
rect 1041 -1178 1042 -1177
rect 2473 -1178 2474 -1177
rect 23 -1180 24 -1179
rect 821 -1180 822 -1179
rect 842 -1180 843 -1179
rect 856 -1180 857 -1179
rect 880 -1180 881 -1179
rect 1745 -1180 1746 -1179
rect 1906 -1180 1907 -1179
rect 2452 -1180 2453 -1179
rect 23 -1182 24 -1181
rect 611 -1182 612 -1181
rect 667 -1182 668 -1181
rect 849 -1182 850 -1181
rect 905 -1182 906 -1181
rect 926 -1182 927 -1181
rect 947 -1182 948 -1181
rect 1433 -1182 1434 -1181
rect 1447 -1182 1448 -1181
rect 2361 -1182 2362 -1181
rect 2368 -1182 2369 -1181
rect 2564 -1182 2565 -1181
rect 30 -1184 31 -1183
rect 677 -1184 678 -1183
rect 751 -1184 752 -1183
rect 842 -1184 843 -1183
rect 912 -1184 913 -1183
rect 1031 -1184 1032 -1183
rect 1048 -1184 1049 -1183
rect 1122 -1184 1123 -1183
rect 1157 -1184 1158 -1183
rect 2263 -1184 2264 -1183
rect 2277 -1184 2278 -1183
rect 2466 -1184 2467 -1183
rect 100 -1186 101 -1185
rect 908 -1186 909 -1185
rect 947 -1186 948 -1185
rect 1094 -1186 1095 -1185
rect 1104 -1186 1105 -1185
rect 2543 -1186 2544 -1185
rect 100 -1188 101 -1187
rect 247 -1188 248 -1187
rect 254 -1188 255 -1187
rect 912 -1188 913 -1187
rect 950 -1188 951 -1187
rect 1451 -1188 1452 -1187
rect 1458 -1188 1459 -1187
rect 1549 -1188 1550 -1187
rect 1552 -1188 1553 -1187
rect 1598 -1188 1599 -1187
rect 1605 -1188 1606 -1187
rect 1906 -1188 1907 -1187
rect 1927 -1188 1928 -1187
rect 2459 -1188 2460 -1187
rect 121 -1190 122 -1189
rect 509 -1190 510 -1189
rect 513 -1190 514 -1189
rect 611 -1190 612 -1189
rect 667 -1190 668 -1189
rect 1269 -1190 1270 -1189
rect 1307 -1190 1308 -1189
rect 2396 -1190 2397 -1189
rect 2431 -1190 2432 -1189
rect 2578 -1190 2579 -1189
rect 124 -1192 125 -1191
rect 1290 -1192 1291 -1191
rect 1335 -1192 1336 -1191
rect 2347 -1192 2348 -1191
rect 2354 -1192 2355 -1191
rect 2557 -1192 2558 -1191
rect 128 -1194 129 -1193
rect 1927 -1194 1928 -1193
rect 1969 -1194 1970 -1193
rect 2389 -1194 2390 -1193
rect 2438 -1194 2439 -1193
rect 2480 -1194 2481 -1193
rect 128 -1196 129 -1195
rect 268 -1196 269 -1195
rect 275 -1196 276 -1195
rect 782 -1196 783 -1195
rect 796 -1196 797 -1195
rect 968 -1196 969 -1195
rect 982 -1196 983 -1195
rect 1094 -1196 1095 -1195
rect 1115 -1196 1116 -1195
rect 1269 -1196 1270 -1195
rect 1339 -1196 1340 -1195
rect 1458 -1196 1459 -1195
rect 1500 -1196 1501 -1195
rect 1598 -1196 1599 -1195
rect 1605 -1196 1606 -1195
rect 1612 -1196 1613 -1195
rect 1745 -1196 1746 -1195
rect 1801 -1196 1802 -1195
rect 2060 -1196 2061 -1195
rect 2263 -1196 2264 -1195
rect 2284 -1196 2285 -1195
rect 2487 -1196 2488 -1195
rect 138 -1198 139 -1197
rect 583 -1198 584 -1197
rect 590 -1198 591 -1197
rect 1815 -1198 1816 -1197
rect 1857 -1198 1858 -1197
rect 2060 -1198 2061 -1197
rect 2095 -1198 2096 -1197
rect 2291 -1198 2292 -1197
rect 2305 -1198 2306 -1197
rect 2501 -1198 2502 -1197
rect 208 -1200 209 -1199
rect 730 -1200 731 -1199
rect 751 -1200 752 -1199
rect 884 -1200 885 -1199
rect 992 -1200 993 -1199
rect 2431 -1200 2432 -1199
rect 37 -1202 38 -1201
rect 884 -1202 885 -1201
rect 1003 -1202 1004 -1201
rect 1829 -1202 1830 -1201
rect 1962 -1202 1963 -1201
rect 2284 -1202 2285 -1201
rect 2312 -1202 2313 -1201
rect 2508 -1202 2509 -1201
rect 37 -1204 38 -1203
rect 702 -1204 703 -1203
rect 758 -1204 759 -1203
rect 1514 -1204 1515 -1203
rect 1521 -1204 1522 -1203
rect 1612 -1204 1613 -1203
rect 1668 -1204 1669 -1203
rect 1829 -1204 1830 -1203
rect 2109 -1204 2110 -1203
rect 2298 -1204 2299 -1203
rect 2319 -1204 2320 -1203
rect 2515 -1204 2516 -1203
rect 268 -1206 269 -1205
rect 2375 -1206 2376 -1205
rect 2424 -1206 2425 -1205
rect 2438 -1206 2439 -1205
rect 275 -1208 276 -1207
rect 2343 -1208 2344 -1207
rect 310 -1210 311 -1209
rect 968 -1210 969 -1209
rect 1003 -1210 1004 -1209
rect 2270 -1210 2271 -1209
rect 2333 -1210 2334 -1209
rect 2536 -1210 2537 -1209
rect 72 -1212 73 -1211
rect 310 -1212 311 -1211
rect 380 -1212 381 -1211
rect 429 -1212 430 -1211
rect 436 -1212 437 -1211
rect 513 -1212 514 -1211
rect 527 -1212 528 -1211
rect 583 -1212 584 -1211
rect 604 -1212 605 -1211
rect 821 -1212 822 -1211
rect 828 -1212 829 -1211
rect 926 -1212 927 -1211
rect 1010 -1212 1011 -1211
rect 1115 -1212 1116 -1211
rect 1164 -1212 1165 -1211
rect 2382 -1212 2383 -1211
rect 72 -1214 73 -1213
rect 443 -1214 444 -1213
rect 485 -1214 486 -1213
rect 548 -1214 549 -1213
rect 555 -1214 556 -1213
rect 590 -1214 591 -1213
rect 642 -1214 643 -1213
rect 1857 -1214 1858 -1213
rect 1920 -1214 1921 -1213
rect 2109 -1214 2110 -1213
rect 2116 -1214 2117 -1213
rect 2305 -1214 2306 -1213
rect 2340 -1214 2341 -1213
rect 2550 -1214 2551 -1213
rect 9 -1216 10 -1215
rect 555 -1216 556 -1215
rect 569 -1216 570 -1215
rect 653 -1216 654 -1215
rect 702 -1216 703 -1215
rect 957 -1216 958 -1215
rect 1038 -1216 1039 -1215
rect 1157 -1216 1158 -1215
rect 1167 -1216 1168 -1215
rect 2571 -1216 2572 -1215
rect 9 -1218 10 -1217
rect 135 -1218 136 -1217
rect 219 -1218 220 -1217
rect 1164 -1218 1165 -1217
rect 1178 -1218 1179 -1217
rect 1843 -1218 1844 -1217
rect 1934 -1218 1935 -1217
rect 2319 -1218 2320 -1217
rect 16 -1220 17 -1219
rect 443 -1220 444 -1219
rect 499 -1220 500 -1219
rect 730 -1220 731 -1219
rect 758 -1220 759 -1219
rect 786 -1220 787 -1219
rect 800 -1220 801 -1219
rect 894 -1220 895 -1219
rect 1045 -1220 1046 -1219
rect 1122 -1220 1123 -1219
rect 1185 -1220 1186 -1219
rect 1339 -1220 1340 -1219
rect 1370 -1220 1371 -1219
rect 2102 -1220 2103 -1219
rect 2116 -1220 2117 -1219
rect 2256 -1220 2257 -1219
rect 65 -1222 66 -1221
rect 569 -1222 570 -1221
rect 800 -1222 801 -1221
rect 1038 -1222 1039 -1221
rect 1045 -1222 1046 -1221
rect 1101 -1222 1102 -1221
rect 1192 -1222 1193 -1221
rect 1290 -1222 1291 -1221
rect 1311 -1222 1312 -1221
rect 1500 -1222 1501 -1221
rect 1563 -1222 1564 -1221
rect 2529 -1222 2530 -1221
rect 65 -1224 66 -1223
rect 79 -1224 80 -1223
rect 114 -1224 115 -1223
rect 2102 -1224 2103 -1223
rect 2144 -1224 2145 -1223
rect 2312 -1224 2313 -1223
rect 114 -1226 115 -1225
rect 646 -1226 647 -1225
rect 807 -1226 808 -1225
rect 810 -1226 811 -1225
rect 852 -1226 853 -1225
rect 1801 -1226 1802 -1225
rect 1815 -1226 1816 -1225
rect 1892 -1226 1893 -1225
rect 1948 -1226 1949 -1225
rect 2144 -1226 2145 -1225
rect 2151 -1226 2152 -1225
rect 2333 -1226 2334 -1225
rect 135 -1228 136 -1227
rect 681 -1228 682 -1227
rect 789 -1228 790 -1227
rect 1948 -1228 1949 -1227
rect 1955 -1228 1956 -1227
rect 2151 -1228 2152 -1227
rect 2158 -1228 2159 -1227
rect 2347 -1228 2348 -1227
rect 191 -1230 192 -1229
rect 219 -1230 220 -1229
rect 373 -1230 374 -1229
rect 499 -1230 500 -1229
rect 506 -1230 507 -1229
rect 2445 -1230 2446 -1229
rect 191 -1232 192 -1231
rect 387 -1232 388 -1231
rect 408 -1232 409 -1231
rect 607 -1232 608 -1231
rect 646 -1232 647 -1231
rect 1087 -1232 1088 -1231
rect 1192 -1232 1193 -1231
rect 1262 -1232 1263 -1231
rect 1283 -1232 1284 -1231
rect 1563 -1232 1564 -1231
rect 1570 -1232 1571 -1231
rect 1668 -1232 1669 -1231
rect 1731 -1232 1732 -1231
rect 1892 -1232 1893 -1231
rect 1955 -1232 1956 -1231
rect 2067 -1232 2068 -1231
rect 2088 -1232 2089 -1231
rect 2256 -1232 2257 -1231
rect 198 -1234 199 -1233
rect 1087 -1234 1088 -1233
rect 1234 -1234 1235 -1233
rect 2410 -1234 2411 -1233
rect 149 -1236 150 -1235
rect 1234 -1236 1235 -1235
rect 1255 -1236 1256 -1235
rect 1262 -1236 1263 -1235
rect 1283 -1236 1284 -1235
rect 1353 -1236 1354 -1235
rect 1381 -1236 1382 -1235
rect 1391 -1236 1392 -1235
rect 1416 -1236 1417 -1235
rect 1521 -1236 1522 -1235
rect 1591 -1236 1592 -1235
rect 1731 -1236 1732 -1235
rect 1738 -1236 1739 -1235
rect 2270 -1236 2271 -1235
rect 145 -1238 146 -1237
rect 149 -1238 150 -1237
rect 198 -1238 199 -1237
rect 1360 -1238 1361 -1237
rect 1381 -1238 1382 -1237
rect 1619 -1238 1620 -1237
rect 1633 -1238 1634 -1237
rect 1738 -1238 1739 -1237
rect 1741 -1238 1742 -1237
rect 2067 -1238 2068 -1237
rect 2172 -1238 2173 -1237
rect 2354 -1238 2355 -1237
rect 233 -1240 234 -1239
rect 408 -1240 409 -1239
rect 422 -1240 423 -1239
rect 1794 -1240 1795 -1239
rect 1885 -1240 1886 -1239
rect 2088 -1240 2089 -1239
rect 2179 -1240 2180 -1239
rect 2361 -1240 2362 -1239
rect 226 -1242 227 -1241
rect 233 -1242 234 -1241
rect 261 -1242 262 -1241
rect 422 -1242 423 -1241
rect 436 -1242 437 -1241
rect 674 -1242 675 -1241
rect 681 -1242 682 -1241
rect 744 -1242 745 -1241
rect 807 -1242 808 -1241
rect 1304 -1242 1305 -1241
rect 1332 -1242 1333 -1241
rect 1962 -1242 1963 -1241
rect 1983 -1242 1984 -1241
rect 2158 -1242 2159 -1241
rect 2186 -1242 2187 -1241
rect 2368 -1242 2369 -1241
rect 261 -1244 262 -1243
rect 1010 -1244 1011 -1243
rect 1059 -1244 1060 -1243
rect 1220 -1244 1221 -1243
rect 1241 -1244 1242 -1243
rect 1353 -1244 1354 -1243
rect 1384 -1244 1385 -1243
rect 2207 -1244 2208 -1243
rect 2221 -1244 2222 -1243
rect 2382 -1244 2383 -1243
rect 303 -1246 304 -1245
rect 373 -1246 374 -1245
rect 380 -1246 381 -1245
rect 457 -1246 458 -1245
rect 506 -1246 507 -1245
rect 723 -1246 724 -1245
rect 744 -1246 745 -1245
rect 954 -1246 955 -1245
rect 961 -1246 962 -1245
rect 1633 -1246 1634 -1245
rect 1654 -1246 1655 -1245
rect 1794 -1246 1795 -1245
rect 1990 -1246 1991 -1245
rect 2179 -1246 2180 -1245
rect 2193 -1246 2194 -1245
rect 2375 -1246 2376 -1245
rect 229 -1248 230 -1247
rect 457 -1248 458 -1247
rect 527 -1248 528 -1247
rect 831 -1248 832 -1247
rect 877 -1248 878 -1247
rect 2095 -1248 2096 -1247
rect 2200 -1248 2201 -1247
rect 2522 -1248 2523 -1247
rect 303 -1250 304 -1249
rect 534 -1250 535 -1249
rect 548 -1250 549 -1249
rect 1181 -1250 1182 -1249
rect 1206 -1250 1207 -1249
rect 1304 -1250 1305 -1249
rect 1325 -1250 1326 -1249
rect 1332 -1250 1333 -1249
rect 1416 -1250 1417 -1249
rect 2123 -1250 2124 -1249
rect 2137 -1250 2138 -1249
rect 2200 -1250 2201 -1249
rect 2228 -1250 2229 -1249
rect 2389 -1250 2390 -1249
rect 331 -1252 332 -1251
rect 387 -1252 388 -1251
rect 520 -1252 521 -1251
rect 534 -1252 535 -1251
rect 562 -1252 563 -1251
rect 786 -1252 787 -1251
rect 891 -1252 892 -1251
rect 961 -1252 962 -1251
rect 975 -1252 976 -1251
rect 1059 -1252 1060 -1251
rect 1073 -1252 1074 -1251
rect 1178 -1252 1179 -1251
rect 1241 -1252 1242 -1251
rect 1248 -1252 1249 -1251
rect 1255 -1252 1256 -1251
rect 1388 -1252 1389 -1251
rect 1423 -1252 1424 -1251
rect 1570 -1252 1571 -1251
rect 1591 -1252 1592 -1251
rect 1724 -1252 1725 -1251
rect 1759 -1252 1760 -1251
rect 1920 -1252 1921 -1251
rect 2004 -1252 2005 -1251
rect 2186 -1252 2187 -1251
rect 2242 -1252 2243 -1251
rect 2396 -1252 2397 -1251
rect 205 -1254 206 -1253
rect 520 -1254 521 -1253
rect 562 -1254 563 -1253
rect 639 -1254 640 -1253
rect 660 -1254 661 -1253
rect 1220 -1254 1221 -1253
rect 1276 -1254 1277 -1253
rect 1388 -1254 1389 -1253
rect 1447 -1254 1448 -1253
rect 2165 -1254 2166 -1253
rect 2249 -1254 2250 -1253
rect 2424 -1254 2425 -1253
rect 205 -1256 206 -1255
rect 2074 -1256 2075 -1255
rect 282 -1258 283 -1257
rect 331 -1258 332 -1257
rect 607 -1258 608 -1257
rect 814 -1258 815 -1257
rect 863 -1258 864 -1257
rect 2242 -1258 2243 -1257
rect 282 -1260 283 -1259
rect 464 -1260 465 -1259
rect 541 -1260 542 -1259
rect 814 -1260 815 -1259
rect 898 -1260 899 -1259
rect 975 -1260 976 -1259
rect 985 -1260 986 -1259
rect 1983 -1260 1984 -1259
rect 2004 -1260 2005 -1259
rect 2130 -1260 2131 -1259
rect 93 -1262 94 -1261
rect 898 -1262 899 -1261
rect 919 -1262 920 -1261
rect 1185 -1262 1186 -1261
rect 1276 -1262 1277 -1261
rect 1297 -1262 1298 -1261
rect 1367 -1262 1368 -1261
rect 1423 -1262 1424 -1261
rect 1451 -1262 1452 -1261
rect 1696 -1262 1697 -1261
rect 1703 -1262 1704 -1261
rect 1885 -1262 1886 -1261
rect 1913 -1262 1914 -1261
rect 2123 -1262 2124 -1261
rect 86 -1264 87 -1263
rect 93 -1264 94 -1263
rect 110 -1264 111 -1263
rect 1703 -1264 1704 -1263
rect 1752 -1264 1753 -1263
rect 1913 -1264 1914 -1263
rect 2018 -1264 2019 -1263
rect 2193 -1264 2194 -1263
rect 86 -1266 87 -1265
rect 597 -1266 598 -1265
rect 632 -1266 633 -1265
rect 674 -1266 675 -1265
rect 709 -1266 710 -1265
rect 919 -1266 920 -1265
rect 954 -1266 955 -1265
rect 964 -1266 965 -1265
rect 1073 -1266 1074 -1265
rect 1216 -1266 1217 -1265
rect 1325 -1266 1326 -1265
rect 1367 -1266 1368 -1265
rect 1402 -1266 1403 -1265
rect 2165 -1266 2166 -1265
rect 44 -1268 45 -1267
rect 709 -1268 710 -1267
rect 723 -1268 724 -1267
rect 1941 -1268 1942 -1267
rect 2032 -1268 2033 -1267
rect 2228 -1268 2229 -1267
rect 44 -1270 45 -1269
rect 324 -1270 325 -1269
rect 464 -1270 465 -1269
rect 835 -1270 836 -1269
rect 1080 -1270 1081 -1269
rect 1206 -1270 1207 -1269
rect 1402 -1270 1403 -1269
rect 1409 -1270 1410 -1269
rect 1507 -1270 1508 -1269
rect 1752 -1270 1753 -1269
rect 1766 -1270 1767 -1269
rect 2018 -1270 2019 -1269
rect 2039 -1270 2040 -1269
rect 2221 -1270 2222 -1269
rect 243 -1272 244 -1271
rect 324 -1272 325 -1271
rect 541 -1272 542 -1271
rect 618 -1272 619 -1271
rect 625 -1272 626 -1271
rect 632 -1272 633 -1271
rect 639 -1272 640 -1271
rect 2417 -1272 2418 -1271
rect 597 -1274 598 -1273
rect 880 -1274 881 -1273
rect 989 -1274 990 -1273
rect 1080 -1274 1081 -1273
rect 1143 -1274 1144 -1273
rect 1360 -1274 1361 -1273
rect 1528 -1274 1529 -1273
rect 1619 -1274 1620 -1273
rect 1626 -1274 1627 -1273
rect 1759 -1274 1760 -1273
rect 1773 -1274 1774 -1273
rect 1941 -1274 1942 -1273
rect 2046 -1274 2047 -1273
rect 2249 -1274 2250 -1273
rect 142 -1276 143 -1275
rect 2046 -1276 2047 -1275
rect 2053 -1276 2054 -1275
rect 2207 -1276 2208 -1275
rect 142 -1278 143 -1277
rect 824 -1278 825 -1277
rect 870 -1278 871 -1277
rect 989 -1278 990 -1277
rect 1136 -1278 1137 -1277
rect 1626 -1278 1627 -1277
rect 1640 -1278 1641 -1277
rect 1766 -1278 1767 -1277
rect 1780 -1278 1781 -1277
rect 1934 -1278 1935 -1277
rect 2011 -1278 2012 -1277
rect 2053 -1278 2054 -1277
rect 618 -1280 619 -1279
rect 1199 -1280 1200 -1279
rect 1227 -1280 1228 -1279
rect 1409 -1280 1410 -1279
rect 1535 -1280 1536 -1279
rect 1640 -1280 1641 -1279
rect 1647 -1280 1648 -1279
rect 1773 -1280 1774 -1279
rect 1780 -1280 1781 -1279
rect 1976 -1280 1977 -1279
rect 625 -1282 626 -1281
rect 779 -1282 780 -1281
rect 996 -1282 997 -1281
rect 1136 -1282 1137 -1281
rect 1143 -1282 1144 -1281
rect 1160 -1282 1161 -1281
rect 1171 -1282 1172 -1281
rect 1227 -1282 1228 -1281
rect 1237 -1282 1238 -1281
rect 1647 -1282 1648 -1281
rect 1661 -1282 1662 -1281
rect 1843 -1282 1844 -1281
rect 1850 -1282 1851 -1281
rect 2039 -1282 2040 -1281
rect 660 -1284 661 -1283
rect 891 -1284 892 -1283
rect 996 -1284 997 -1283
rect 2172 -1284 2173 -1283
rect 688 -1286 689 -1285
rect 835 -1286 836 -1285
rect 999 -1286 1000 -1285
rect 1199 -1286 1200 -1285
rect 1311 -1286 1312 -1285
rect 1507 -1286 1508 -1285
rect 1542 -1286 1543 -1285
rect 1654 -1286 1655 -1285
rect 1717 -1286 1718 -1285
rect 2011 -1286 2012 -1285
rect 688 -1288 689 -1287
rect 866 -1288 867 -1287
rect 1052 -1288 1053 -1287
rect 1171 -1288 1172 -1287
rect 1391 -1288 1392 -1287
rect 1528 -1288 1529 -1287
rect 1556 -1288 1557 -1287
rect 1661 -1288 1662 -1287
rect 1787 -1288 1788 -1287
rect 2277 -1288 2278 -1287
rect 765 -1290 766 -1289
rect 1248 -1290 1249 -1289
rect 1430 -1290 1431 -1289
rect 1717 -1290 1718 -1289
rect 1808 -1290 1809 -1289
rect 1990 -1290 1991 -1289
rect 695 -1292 696 -1291
rect 765 -1292 766 -1291
rect 1024 -1292 1025 -1291
rect 1052 -1292 1053 -1291
rect 1150 -1292 1151 -1291
rect 1297 -1292 1298 -1291
rect 1430 -1292 1431 -1291
rect 1969 -1292 1970 -1291
rect 695 -1294 696 -1293
rect 940 -1294 941 -1293
rect 1024 -1294 1025 -1293
rect 1066 -1294 1067 -1293
rect 1108 -1294 1109 -1293
rect 1150 -1294 1151 -1293
rect 1213 -1294 1214 -1293
rect 1787 -1294 1788 -1293
rect 1836 -1294 1837 -1293
rect 2032 -1294 2033 -1293
rect 51 -1296 52 -1295
rect 940 -1296 941 -1295
rect 1108 -1296 1109 -1295
rect 1129 -1296 1130 -1295
rect 1153 -1296 1154 -1295
rect 1836 -1296 1837 -1295
rect 1850 -1296 1851 -1295
rect 2392 -1296 2393 -1295
rect 51 -1298 52 -1297
rect 58 -1298 59 -1297
rect 450 -1298 451 -1297
rect 1066 -1298 1067 -1297
rect 1213 -1298 1214 -1297
rect 2214 -1298 2215 -1297
rect 58 -1300 59 -1299
rect 79 -1300 80 -1299
rect 450 -1300 451 -1299
rect 576 -1300 577 -1299
rect 1017 -1300 1018 -1299
rect 1129 -1300 1130 -1299
rect 1444 -1300 1445 -1299
rect 1535 -1300 1536 -1299
rect 1556 -1300 1557 -1299
rect 2403 -1300 2404 -1299
rect 352 -1302 353 -1301
rect 576 -1302 577 -1301
rect 933 -1302 934 -1301
rect 1017 -1302 1018 -1301
rect 1479 -1302 1480 -1301
rect 1976 -1302 1977 -1301
rect 2025 -1302 2026 -1301
rect 2214 -1302 2215 -1301
rect 352 -1304 353 -1303
rect 401 -1304 402 -1303
rect 793 -1304 794 -1303
rect 933 -1304 934 -1303
rect 1013 -1304 1014 -1303
rect 2025 -1304 2026 -1303
rect 2081 -1304 2082 -1303
rect 2403 -1304 2404 -1303
rect 394 -1306 395 -1305
rect 401 -1306 402 -1305
rect 761 -1306 762 -1305
rect 2081 -1306 2082 -1305
rect 212 -1308 213 -1307
rect 394 -1308 395 -1307
rect 793 -1308 794 -1307
rect 1997 -1308 1998 -1307
rect 212 -1310 213 -1309
rect 415 -1310 416 -1309
rect 1395 -1310 1396 -1309
rect 1479 -1310 1480 -1309
rect 1493 -1310 1494 -1309
rect 1542 -1310 1543 -1309
rect 1577 -1310 1578 -1309
rect 1696 -1310 1697 -1309
rect 1864 -1310 1865 -1309
rect 2074 -1310 2075 -1309
rect 170 -1312 171 -1311
rect 415 -1312 416 -1311
rect 1006 -1312 1007 -1311
rect 1864 -1312 1865 -1311
rect 1871 -1312 1872 -1311
rect 2130 -1312 2131 -1311
rect 107 -1314 108 -1313
rect 1006 -1314 1007 -1313
rect 1346 -1314 1347 -1313
rect 1493 -1314 1494 -1313
rect 1584 -1314 1585 -1313
rect 1724 -1314 1725 -1313
rect 1878 -1314 1879 -1313
rect 2137 -1314 2138 -1313
rect 170 -1316 171 -1315
rect 737 -1316 738 -1315
rect 1395 -1316 1396 -1315
rect 1437 -1316 1438 -1315
rect 1465 -1316 1466 -1315
rect 1878 -1316 1879 -1315
rect 247 -1318 248 -1317
rect 1346 -1318 1347 -1317
rect 1472 -1318 1473 -1317
rect 1577 -1318 1578 -1317
rect 1675 -1318 1676 -1317
rect 1808 -1318 1809 -1317
rect 716 -1320 717 -1319
rect 737 -1320 738 -1319
rect 779 -1320 780 -1319
rect 1465 -1320 1466 -1319
rect 1472 -1320 1473 -1319
rect 1710 -1320 1711 -1319
rect 359 -1322 360 -1321
rect 716 -1322 717 -1321
rect 1318 -1322 1319 -1321
rect 1437 -1322 1438 -1321
rect 1486 -1322 1487 -1321
rect 1584 -1322 1585 -1321
rect 1675 -1322 1676 -1321
rect 2235 -1322 2236 -1321
rect 163 -1324 164 -1323
rect 359 -1324 360 -1323
rect 1202 -1324 1203 -1323
rect 1318 -1324 1319 -1323
rect 1374 -1324 1375 -1323
rect 1486 -1324 1487 -1323
rect 1510 -1324 1511 -1323
rect 2235 -1324 2236 -1323
rect 156 -1326 157 -1325
rect 163 -1326 164 -1325
rect 177 -1326 178 -1325
rect 1374 -1326 1375 -1325
rect 1682 -1326 1683 -1325
rect 1871 -1326 1872 -1325
rect 156 -1328 157 -1327
rect 240 -1328 241 -1327
rect 1682 -1328 1683 -1327
rect 2326 -1328 2327 -1327
rect 177 -1330 178 -1329
rect 184 -1330 185 -1329
rect 240 -1330 241 -1329
rect 296 -1330 297 -1329
rect 1689 -1330 1690 -1329
rect 1997 -1330 1998 -1329
rect 184 -1332 185 -1331
rect 289 -1332 290 -1331
rect 296 -1332 297 -1331
rect 478 -1332 479 -1331
rect 1101 -1332 1102 -1331
rect 1689 -1332 1690 -1331
rect 1710 -1332 1711 -1331
rect 1899 -1332 1900 -1331
rect 289 -1334 290 -1333
rect 471 -1334 472 -1333
rect 1822 -1334 1823 -1333
rect 2326 -1334 2327 -1333
rect 317 -1336 318 -1335
rect 478 -1336 479 -1335
rect 828 -1336 829 -1335
rect 1822 -1336 1823 -1335
rect 1899 -1336 1900 -1335
rect 2340 -1336 2341 -1335
rect 317 -1338 318 -1337
rect 726 -1338 727 -1337
rect 366 -1340 367 -1339
rect 471 -1340 472 -1339
rect 345 -1342 346 -1341
rect 366 -1342 367 -1341
rect 345 -1344 346 -1343
rect 492 -1344 493 -1343
rect 338 -1346 339 -1345
rect 492 -1346 493 -1345
rect 121 -1348 122 -1347
rect 338 -1348 339 -1347
rect 2 -1359 3 -1358
rect 838 -1359 839 -1358
rect 880 -1359 881 -1358
rect 1136 -1359 1137 -1358
rect 1150 -1359 1151 -1358
rect 2263 -1359 2264 -1358
rect 2343 -1359 2344 -1358
rect 2578 -1359 2579 -1358
rect 26 -1361 27 -1360
rect 1577 -1361 1578 -1360
rect 1794 -1361 1795 -1360
rect 1797 -1361 1798 -1360
rect 2263 -1361 2264 -1360
rect 2361 -1361 2362 -1360
rect 37 -1363 38 -1362
rect 989 -1363 990 -1362
rect 996 -1363 997 -1362
rect 1717 -1363 1718 -1362
rect 1794 -1363 1795 -1362
rect 1850 -1363 1851 -1362
rect 2361 -1363 2362 -1362
rect 2424 -1363 2425 -1362
rect 40 -1365 41 -1364
rect 1983 -1365 1984 -1364
rect 44 -1367 45 -1366
rect 201 -1367 202 -1366
rect 208 -1367 209 -1366
rect 436 -1367 437 -1366
rect 464 -1367 465 -1366
rect 908 -1367 909 -1366
rect 943 -1367 944 -1366
rect 1976 -1367 1977 -1366
rect 1983 -1367 1984 -1366
rect 2368 -1367 2369 -1366
rect 44 -1369 45 -1368
rect 86 -1369 87 -1368
rect 89 -1369 90 -1368
rect 968 -1369 969 -1368
rect 989 -1369 990 -1368
rect 1115 -1369 1116 -1368
rect 1136 -1369 1137 -1368
rect 1192 -1369 1193 -1368
rect 1213 -1369 1214 -1368
rect 1556 -1369 1557 -1368
rect 1577 -1369 1578 -1368
rect 1605 -1369 1606 -1368
rect 1717 -1369 1718 -1368
rect 1766 -1369 1767 -1368
rect 1850 -1369 1851 -1368
rect 1913 -1369 1914 -1368
rect 1976 -1369 1977 -1368
rect 2039 -1369 2040 -1368
rect 2368 -1369 2369 -1368
rect 2431 -1369 2432 -1368
rect 54 -1371 55 -1370
rect 86 -1371 87 -1370
rect 93 -1371 94 -1370
rect 124 -1371 125 -1370
rect 170 -1371 171 -1370
rect 268 -1371 269 -1370
rect 317 -1371 318 -1370
rect 464 -1371 465 -1370
rect 499 -1371 500 -1370
rect 628 -1371 629 -1370
rect 642 -1371 643 -1370
rect 968 -1371 969 -1370
rect 996 -1371 997 -1370
rect 1500 -1371 1501 -1370
rect 1507 -1371 1508 -1370
rect 1773 -1371 1774 -1370
rect 1913 -1371 1914 -1370
rect 1962 -1371 1963 -1370
rect 2431 -1371 2432 -1370
rect 2480 -1371 2481 -1370
rect 58 -1373 59 -1372
rect 61 -1373 62 -1372
rect 72 -1373 73 -1372
rect 824 -1373 825 -1372
rect 831 -1373 832 -1372
rect 905 -1373 906 -1372
rect 957 -1373 958 -1372
rect 1423 -1373 1424 -1372
rect 1426 -1373 1427 -1372
rect 1864 -1373 1865 -1372
rect 1962 -1373 1963 -1372
rect 2032 -1373 2033 -1372
rect 58 -1375 59 -1374
rect 65 -1375 66 -1374
rect 79 -1375 80 -1374
rect 156 -1375 157 -1374
rect 170 -1375 171 -1374
rect 236 -1375 237 -1374
rect 240 -1375 241 -1374
rect 639 -1375 640 -1374
rect 646 -1375 647 -1374
rect 954 -1375 955 -1374
rect 982 -1375 983 -1374
rect 2480 -1375 2481 -1374
rect 82 -1377 83 -1376
rect 1752 -1377 1753 -1376
rect 1766 -1377 1767 -1376
rect 2109 -1377 2110 -1376
rect 93 -1379 94 -1378
rect 296 -1379 297 -1378
rect 317 -1379 318 -1378
rect 887 -1379 888 -1378
rect 891 -1379 892 -1378
rect 2529 -1379 2530 -1378
rect 107 -1381 108 -1380
rect 604 -1381 605 -1380
rect 646 -1381 647 -1380
rect 653 -1381 654 -1380
rect 681 -1381 682 -1380
rect 999 -1381 1000 -1380
rect 1006 -1381 1007 -1380
rect 1433 -1381 1434 -1380
rect 1472 -1381 1473 -1380
rect 1752 -1381 1753 -1380
rect 1773 -1381 1774 -1380
rect 1822 -1381 1823 -1380
rect 1864 -1381 1865 -1380
rect 1920 -1381 1921 -1380
rect 2109 -1381 2110 -1380
rect 2193 -1381 2194 -1380
rect 2529 -1381 2530 -1380
rect 2557 -1381 2558 -1380
rect 110 -1383 111 -1382
rect 1787 -1383 1788 -1382
rect 1797 -1383 1798 -1382
rect 2032 -1383 2033 -1382
rect 2193 -1383 2194 -1382
rect 2291 -1383 2292 -1382
rect 2340 -1383 2341 -1382
rect 2557 -1383 2558 -1382
rect 117 -1385 118 -1384
rect 208 -1385 209 -1384
rect 226 -1385 227 -1384
rect 1374 -1385 1375 -1384
rect 1430 -1385 1431 -1384
rect 1871 -1385 1872 -1384
rect 2200 -1385 2201 -1384
rect 2340 -1385 2341 -1384
rect 121 -1387 122 -1386
rect 1234 -1387 1235 -1386
rect 1251 -1387 1252 -1386
rect 2326 -1387 2327 -1386
rect 107 -1389 108 -1388
rect 121 -1389 122 -1388
rect 128 -1389 129 -1388
rect 653 -1389 654 -1388
rect 681 -1389 682 -1388
rect 737 -1389 738 -1388
rect 772 -1389 773 -1388
rect 782 -1389 783 -1388
rect 796 -1389 797 -1388
rect 912 -1389 913 -1388
rect 954 -1389 955 -1388
rect 975 -1389 976 -1388
rect 982 -1389 983 -1388
rect 1073 -1389 1074 -1388
rect 1087 -1389 1088 -1388
rect 1192 -1389 1193 -1388
rect 1213 -1389 1214 -1388
rect 1227 -1389 1228 -1388
rect 1234 -1389 1235 -1388
rect 1304 -1389 1305 -1388
rect 1332 -1389 1333 -1388
rect 1430 -1389 1431 -1388
rect 1472 -1389 1473 -1388
rect 1486 -1389 1487 -1388
rect 1500 -1389 1501 -1388
rect 2270 -1389 2271 -1388
rect 128 -1391 129 -1390
rect 992 -1391 993 -1390
rect 1013 -1391 1014 -1390
rect 1759 -1391 1760 -1390
rect 1787 -1391 1788 -1390
rect 1836 -1391 1837 -1390
rect 1871 -1391 1872 -1390
rect 1934 -1391 1935 -1390
rect 2200 -1391 2201 -1390
rect 2508 -1391 2509 -1390
rect 226 -1393 227 -1392
rect 485 -1393 486 -1392
rect 516 -1393 517 -1392
rect 569 -1393 570 -1392
rect 723 -1393 724 -1392
rect 1090 -1393 1091 -1392
rect 1104 -1393 1105 -1392
rect 1675 -1393 1676 -1392
rect 1759 -1393 1760 -1392
rect 1815 -1393 1816 -1392
rect 1822 -1393 1823 -1392
rect 1892 -1393 1893 -1392
rect 1934 -1393 1935 -1392
rect 1997 -1393 1998 -1392
rect 2270 -1393 2271 -1392
rect 2382 -1393 2383 -1392
rect 2508 -1393 2509 -1392
rect 2522 -1393 2523 -1392
rect 229 -1395 230 -1394
rect 1920 -1395 1921 -1394
rect 1997 -1395 1998 -1394
rect 2074 -1395 2075 -1394
rect 2116 -1395 2117 -1394
rect 2382 -1395 2383 -1394
rect 2522 -1395 2523 -1394
rect 2543 -1395 2544 -1394
rect 240 -1397 241 -1396
rect 751 -1397 752 -1396
rect 772 -1397 773 -1396
rect 842 -1397 843 -1396
rect 880 -1397 881 -1396
rect 919 -1397 920 -1396
rect 1038 -1397 1039 -1396
rect 1360 -1397 1361 -1396
rect 1370 -1397 1371 -1396
rect 2424 -1397 2425 -1396
rect 2543 -1397 2544 -1396
rect 2571 -1397 2572 -1396
rect 254 -1399 255 -1398
rect 688 -1399 689 -1398
rect 726 -1399 727 -1398
rect 866 -1399 867 -1398
rect 891 -1399 892 -1398
rect 961 -1399 962 -1398
rect 1031 -1399 1032 -1398
rect 1038 -1399 1039 -1398
rect 1041 -1399 1042 -1398
rect 2165 -1399 2166 -1398
rect 254 -1401 255 -1400
rect 618 -1401 619 -1400
rect 688 -1401 689 -1400
rect 758 -1401 759 -1400
rect 779 -1401 780 -1400
rect 1878 -1401 1879 -1400
rect 2165 -1401 2166 -1400
rect 2256 -1401 2257 -1400
rect 296 -1403 297 -1402
rect 894 -1403 895 -1402
rect 898 -1403 899 -1402
rect 975 -1403 976 -1402
rect 1066 -1403 1067 -1402
rect 1101 -1403 1102 -1402
rect 1115 -1403 1116 -1402
rect 1297 -1403 1298 -1402
rect 1304 -1403 1305 -1402
rect 1451 -1403 1452 -1402
rect 1482 -1403 1483 -1402
rect 2123 -1403 2124 -1402
rect 2256 -1403 2257 -1402
rect 2354 -1403 2355 -1402
rect 16 -1405 17 -1404
rect 1451 -1405 1452 -1404
rect 1510 -1405 1511 -1404
rect 2277 -1405 2278 -1404
rect 16 -1407 17 -1406
rect 2116 -1407 2117 -1406
rect 2123 -1407 2124 -1406
rect 2207 -1407 2208 -1406
rect 2277 -1407 2278 -1406
rect 2410 -1407 2411 -1406
rect 310 -1409 311 -1408
rect 604 -1409 605 -1408
rect 618 -1409 619 -1408
rect 702 -1409 703 -1408
rect 730 -1409 731 -1408
rect 740 -1409 741 -1408
rect 758 -1409 759 -1408
rect 870 -1409 871 -1408
rect 905 -1409 906 -1408
rect 2039 -1409 2040 -1408
rect 2207 -1409 2208 -1408
rect 2445 -1409 2446 -1408
rect 184 -1411 185 -1410
rect 310 -1411 311 -1410
rect 408 -1411 409 -1410
rect 863 -1411 864 -1410
rect 866 -1411 867 -1410
rect 2130 -1411 2131 -1410
rect 2410 -1411 2411 -1410
rect 2459 -1411 2460 -1410
rect 184 -1413 185 -1412
rect 275 -1413 276 -1412
rect 366 -1413 367 -1412
rect 408 -1413 409 -1412
rect 415 -1413 416 -1412
rect 607 -1413 608 -1412
rect 642 -1413 643 -1412
rect 2354 -1413 2355 -1412
rect 2445 -1413 2446 -1412
rect 2494 -1413 2495 -1412
rect 257 -1415 258 -1414
rect 415 -1415 416 -1414
rect 422 -1415 423 -1414
rect 593 -1415 594 -1414
rect 702 -1415 703 -1414
rect 1178 -1415 1179 -1414
rect 1227 -1415 1228 -1414
rect 1248 -1415 1249 -1414
rect 1258 -1415 1259 -1414
rect 2172 -1415 2173 -1414
rect 219 -1417 220 -1416
rect 422 -1417 423 -1416
rect 429 -1417 430 -1416
rect 569 -1417 570 -1416
rect 730 -1417 731 -1416
rect 1349 -1417 1350 -1416
rect 1384 -1417 1385 -1416
rect 1675 -1417 1676 -1416
rect 1682 -1417 1683 -1416
rect 2494 -1417 2495 -1416
rect 19 -1419 20 -1418
rect 429 -1419 430 -1418
rect 436 -1419 437 -1418
rect 1311 -1419 1312 -1418
rect 1332 -1419 1333 -1418
rect 1353 -1419 1354 -1418
rect 1556 -1419 1557 -1418
rect 1584 -1419 1585 -1418
rect 1591 -1419 1592 -1418
rect 1892 -1419 1893 -1418
rect 2172 -1419 2173 -1418
rect 2242 -1419 2243 -1418
rect 149 -1421 150 -1420
rect 219 -1421 220 -1420
rect 247 -1421 248 -1420
rect 1682 -1421 1683 -1420
rect 1780 -1421 1781 -1420
rect 2074 -1421 2075 -1420
rect 2242 -1421 2243 -1420
rect 2333 -1421 2334 -1420
rect 149 -1423 150 -1422
rect 765 -1423 766 -1422
rect 789 -1423 790 -1422
rect 2459 -1423 2460 -1422
rect 247 -1425 248 -1424
rect 352 -1425 353 -1424
rect 366 -1425 367 -1424
rect 492 -1425 493 -1424
rect 506 -1425 507 -1424
rect 751 -1425 752 -1424
rect 765 -1425 766 -1424
rect 1171 -1425 1172 -1424
rect 1178 -1425 1179 -1424
rect 1290 -1425 1291 -1424
rect 1297 -1425 1298 -1424
rect 1325 -1425 1326 -1424
rect 1353 -1425 1354 -1424
rect 1493 -1425 1494 -1424
rect 1584 -1425 1585 -1424
rect 1885 -1425 1886 -1424
rect 142 -1427 143 -1426
rect 1290 -1427 1291 -1426
rect 1311 -1427 1312 -1426
rect 1339 -1427 1340 -1426
rect 1591 -1427 1592 -1426
rect 1633 -1427 1634 -1426
rect 1780 -1427 1781 -1426
rect 1829 -1427 1830 -1426
rect 1836 -1427 1837 -1426
rect 1899 -1427 1900 -1426
rect 142 -1429 143 -1428
rect 985 -1429 986 -1428
rect 1003 -1429 1004 -1428
rect 1325 -1429 1326 -1428
rect 1605 -1429 1606 -1428
rect 1647 -1429 1648 -1428
rect 1815 -1429 1816 -1428
rect 1857 -1429 1858 -1428
rect 1878 -1429 1879 -1428
rect 1955 -1429 1956 -1428
rect 275 -1431 276 -1430
rect 359 -1431 360 -1430
rect 471 -1431 472 -1430
rect 506 -1431 507 -1430
rect 541 -1431 542 -1430
rect 1010 -1431 1011 -1430
rect 1024 -1431 1025 -1430
rect 1101 -1431 1102 -1430
rect 1150 -1431 1151 -1430
rect 1185 -1431 1186 -1430
rect 1241 -1431 1242 -1430
rect 1339 -1431 1340 -1430
rect 1619 -1431 1620 -1430
rect 1829 -1431 1830 -1430
rect 1857 -1431 1858 -1430
rect 1927 -1431 1928 -1430
rect 1955 -1431 1956 -1430
rect 2025 -1431 2026 -1430
rect 289 -1433 290 -1432
rect 492 -1433 493 -1432
rect 541 -1433 542 -1432
rect 1419 -1433 1420 -1432
rect 1489 -1433 1490 -1432
rect 1619 -1433 1620 -1432
rect 1633 -1433 1634 -1432
rect 1668 -1433 1669 -1432
rect 1885 -1433 1886 -1432
rect 1948 -1433 1949 -1432
rect 2025 -1433 2026 -1432
rect 2095 -1433 2096 -1432
rect 289 -1435 290 -1434
rect 548 -1435 549 -1434
rect 555 -1435 556 -1434
rect 779 -1435 780 -1434
rect 814 -1435 815 -1434
rect 1087 -1435 1088 -1434
rect 1153 -1435 1154 -1434
rect 2291 -1435 2292 -1434
rect 135 -1437 136 -1436
rect 548 -1437 549 -1436
rect 716 -1437 717 -1436
rect 1003 -1437 1004 -1436
rect 1010 -1437 1011 -1436
rect 1052 -1437 1053 -1436
rect 1059 -1437 1060 -1436
rect 1066 -1437 1067 -1436
rect 1185 -1437 1186 -1436
rect 1206 -1437 1207 -1436
rect 1241 -1437 1242 -1436
rect 1262 -1437 1263 -1436
rect 1283 -1437 1284 -1436
rect 1360 -1437 1361 -1436
rect 1647 -1437 1648 -1436
rect 1689 -1437 1690 -1436
rect 1899 -1437 1900 -1436
rect 2179 -1437 2180 -1436
rect 135 -1439 136 -1438
rect 667 -1439 668 -1438
rect 716 -1439 717 -1438
rect 828 -1439 829 -1438
rect 835 -1439 836 -1438
rect 1073 -1439 1074 -1438
rect 1206 -1439 1207 -1438
rect 1220 -1439 1221 -1438
rect 1248 -1439 1249 -1438
rect 2326 -1439 2327 -1438
rect 250 -1441 251 -1440
rect 1220 -1441 1221 -1440
rect 1255 -1441 1256 -1440
rect 1493 -1441 1494 -1440
rect 1668 -1441 1669 -1440
rect 1724 -1441 1725 -1440
rect 1927 -1441 1928 -1440
rect 2004 -1441 2005 -1440
rect 2067 -1441 2068 -1440
rect 2179 -1441 2180 -1440
rect 261 -1443 262 -1442
rect 555 -1443 556 -1442
rect 677 -1443 678 -1442
rect 1255 -1443 1256 -1442
rect 1262 -1443 1263 -1442
rect 1269 -1443 1270 -1442
rect 1283 -1443 1284 -1442
rect 1941 -1443 1942 -1442
rect 1948 -1443 1949 -1442
rect 2018 -1443 2019 -1442
rect 261 -1445 262 -1444
rect 520 -1445 521 -1444
rect 674 -1445 675 -1444
rect 1269 -1445 1270 -1444
rect 1381 -1445 1382 -1444
rect 1689 -1445 1690 -1444
rect 1941 -1445 1942 -1444
rect 2011 -1445 2012 -1444
rect 2018 -1445 2019 -1444
rect 2088 -1445 2089 -1444
rect 9 -1447 10 -1446
rect 520 -1447 521 -1446
rect 674 -1447 675 -1446
rect 691 -1447 692 -1446
rect 737 -1447 738 -1446
rect 2130 -1447 2131 -1446
rect 9 -1449 10 -1448
rect 1265 -1449 1266 -1448
rect 1381 -1449 1382 -1448
rect 1388 -1449 1389 -1448
rect 1503 -1449 1504 -1448
rect 1724 -1449 1725 -1448
rect 1969 -1449 1970 -1448
rect 2095 -1449 2096 -1448
rect 303 -1451 304 -1450
rect 359 -1451 360 -1450
rect 450 -1451 451 -1450
rect 667 -1451 668 -1450
rect 744 -1451 745 -1450
rect 1052 -1451 1053 -1450
rect 1388 -1451 1389 -1450
rect 1402 -1451 1403 -1450
rect 1514 -1451 1515 -1450
rect 2067 -1451 2068 -1450
rect 2088 -1451 2089 -1450
rect 2186 -1451 2187 -1450
rect 177 -1453 178 -1452
rect 303 -1453 304 -1452
rect 352 -1453 353 -1452
rect 373 -1453 374 -1452
rect 450 -1453 451 -1452
rect 597 -1453 598 -1452
rect 709 -1453 710 -1452
rect 744 -1453 745 -1452
rect 786 -1453 787 -1452
rect 2186 -1453 2187 -1452
rect 177 -1455 178 -1454
rect 191 -1455 192 -1454
rect 271 -1455 272 -1454
rect 709 -1455 710 -1454
rect 786 -1455 787 -1454
rect 947 -1455 948 -1454
rect 1024 -1455 1025 -1454
rect 1164 -1455 1165 -1454
rect 1276 -1455 1277 -1454
rect 1402 -1455 1403 -1454
rect 1969 -1455 1970 -1454
rect 2060 -1455 2061 -1454
rect 191 -1457 192 -1456
rect 345 -1457 346 -1456
rect 373 -1457 374 -1456
rect 401 -1457 402 -1456
rect 443 -1457 444 -1456
rect 597 -1457 598 -1456
rect 660 -1457 661 -1456
rect 947 -1457 948 -1456
rect 1031 -1457 1032 -1456
rect 1153 -1457 1154 -1456
rect 1157 -1457 1158 -1456
rect 1514 -1457 1515 -1456
rect 2004 -1457 2005 -1456
rect 2249 -1457 2250 -1456
rect 331 -1459 332 -1458
rect 345 -1459 346 -1458
rect 401 -1459 402 -1458
rect 1286 -1459 1287 -1458
rect 2011 -1459 2012 -1458
rect 2081 -1459 2082 -1458
rect 2249 -1459 2250 -1458
rect 2347 -1459 2348 -1458
rect 331 -1461 332 -1460
rect 590 -1461 591 -1460
rect 632 -1461 633 -1460
rect 660 -1461 661 -1460
rect 814 -1461 815 -1460
rect 926 -1461 927 -1460
rect 940 -1461 941 -1460
rect 1059 -1461 1060 -1460
rect 1122 -1461 1123 -1460
rect 1276 -1461 1277 -1460
rect 2060 -1461 2061 -1460
rect 2151 -1461 2152 -1460
rect 2347 -1461 2348 -1460
rect 2417 -1461 2418 -1460
rect 114 -1463 115 -1462
rect 632 -1463 633 -1462
rect 828 -1463 829 -1462
rect 1612 -1463 1613 -1462
rect 2081 -1463 2082 -1462
rect 2158 -1463 2159 -1462
rect 2417 -1463 2418 -1462
rect 2473 -1463 2474 -1462
rect 51 -1465 52 -1464
rect 114 -1465 115 -1464
rect 443 -1465 444 -1464
rect 796 -1465 797 -1464
rect 835 -1465 836 -1464
rect 849 -1465 850 -1464
rect 856 -1465 857 -1464
rect 898 -1465 899 -1464
rect 912 -1465 913 -1464
rect 1444 -1465 1445 -1464
rect 1612 -1465 1613 -1464
rect 1654 -1465 1655 -1464
rect 2151 -1465 2152 -1464
rect 2228 -1465 2229 -1464
rect 2473 -1465 2474 -1464
rect 2515 -1465 2516 -1464
rect 51 -1467 52 -1466
rect 842 -1467 843 -1466
rect 870 -1467 871 -1466
rect 884 -1467 885 -1466
rect 919 -1467 920 -1466
rect 1017 -1467 1018 -1466
rect 1122 -1467 1123 -1466
rect 1143 -1467 1144 -1466
rect 1157 -1467 1158 -1466
rect 2452 -1467 2453 -1466
rect 2515 -1467 2516 -1466
rect 2536 -1467 2537 -1466
rect 471 -1469 472 -1468
rect 800 -1469 801 -1468
rect 884 -1469 885 -1468
rect 1563 -1469 1564 -1468
rect 1654 -1469 1655 -1468
rect 1696 -1469 1697 -1468
rect 2158 -1469 2159 -1468
rect 2235 -1469 2236 -1468
rect 2452 -1469 2453 -1468
rect 2501 -1469 2502 -1468
rect 2536 -1469 2537 -1468
rect 2550 -1469 2551 -1468
rect 338 -1471 339 -1470
rect 800 -1471 801 -1470
rect 926 -1471 927 -1470
rect 933 -1471 934 -1470
rect 940 -1471 941 -1470
rect 2333 -1471 2334 -1470
rect 2375 -1471 2376 -1470
rect 2550 -1471 2551 -1470
rect 205 -1473 206 -1472
rect 933 -1473 934 -1472
rect 1017 -1473 1018 -1472
rect 2144 -1473 2145 -1472
rect 2228 -1473 2229 -1472
rect 2312 -1473 2313 -1472
rect 338 -1475 339 -1474
rect 457 -1475 458 -1474
rect 478 -1475 479 -1474
rect 499 -1475 500 -1474
rect 562 -1475 563 -1474
rect 856 -1475 857 -1474
rect 877 -1475 878 -1474
rect 2375 -1475 2376 -1474
rect 23 -1477 24 -1476
rect 562 -1477 563 -1476
rect 625 -1477 626 -1476
rect 849 -1477 850 -1476
rect 1143 -1477 1144 -1476
rect 1521 -1477 1522 -1476
rect 1563 -1477 1564 -1476
rect 1598 -1477 1599 -1476
rect 1696 -1477 1697 -1476
rect 1731 -1477 1732 -1476
rect 1990 -1477 1991 -1476
rect 2235 -1477 2236 -1476
rect 2312 -1477 2313 -1476
rect 2396 -1477 2397 -1476
rect 2 -1479 3 -1478
rect 625 -1479 626 -1478
rect 793 -1479 794 -1478
rect 1731 -1479 1732 -1478
rect 1990 -1479 1991 -1478
rect 2298 -1479 2299 -1478
rect 2396 -1479 2397 -1478
rect 2466 -1479 2467 -1478
rect 23 -1481 24 -1480
rect 2102 -1481 2103 -1480
rect 2144 -1481 2145 -1480
rect 2221 -1481 2222 -1480
rect 2284 -1481 2285 -1480
rect 2466 -1481 2467 -1480
rect 156 -1483 157 -1482
rect 877 -1483 878 -1482
rect 1160 -1483 1161 -1482
rect 1444 -1483 1445 -1482
rect 1486 -1483 1487 -1482
rect 2501 -1483 2502 -1482
rect 380 -1485 381 -1484
rect 457 -1485 458 -1484
rect 485 -1485 486 -1484
rect 513 -1485 514 -1484
rect 1164 -1485 1165 -1484
rect 1199 -1485 1200 -1484
rect 1521 -1485 1522 -1484
rect 1542 -1485 1543 -1484
rect 1598 -1485 1599 -1484
rect 1640 -1485 1641 -1484
rect 2046 -1485 2047 -1484
rect 2221 -1485 2222 -1484
rect 2284 -1485 2285 -1484
rect 2564 -1485 2565 -1484
rect 47 -1487 48 -1486
rect 513 -1487 514 -1486
rect 1080 -1487 1081 -1486
rect 1199 -1487 1200 -1486
rect 1367 -1487 1368 -1486
rect 1640 -1487 1641 -1486
rect 2046 -1487 2047 -1486
rect 2137 -1487 2138 -1486
rect 2298 -1487 2299 -1486
rect 2389 -1487 2390 -1486
rect 212 -1489 213 -1488
rect 380 -1489 381 -1488
rect 394 -1489 395 -1488
rect 478 -1489 479 -1488
rect 821 -1489 822 -1488
rect 1367 -1489 1368 -1488
rect 1542 -1489 1543 -1488
rect 1549 -1489 1550 -1488
rect 2053 -1489 2054 -1488
rect 2102 -1489 2103 -1488
rect 2137 -1489 2138 -1488
rect 2214 -1489 2215 -1488
rect 2389 -1489 2390 -1488
rect 2438 -1489 2439 -1488
rect 212 -1491 213 -1490
rect 807 -1491 808 -1490
rect 1080 -1491 1081 -1490
rect 1094 -1491 1095 -1490
rect 1549 -1491 1550 -1490
rect 1570 -1491 1571 -1490
rect 1801 -1491 1802 -1490
rect 2053 -1491 2054 -1490
rect 2214 -1491 2215 -1490
rect 2305 -1491 2306 -1490
rect 2438 -1491 2439 -1490
rect 2487 -1491 2488 -1490
rect 37 -1493 38 -1492
rect 2487 -1493 2488 -1492
rect 394 -1495 395 -1494
rect 534 -1495 535 -1494
rect 807 -1495 808 -1494
rect 1374 -1495 1375 -1494
rect 1535 -1495 1536 -1494
rect 2305 -1495 2306 -1494
rect 324 -1497 325 -1496
rect 534 -1497 535 -1496
rect 1094 -1497 1095 -1496
rect 1108 -1497 1109 -1496
rect 1395 -1497 1396 -1496
rect 1535 -1497 1536 -1496
rect 1570 -1497 1571 -1496
rect 1626 -1497 1627 -1496
rect 1801 -1497 1802 -1496
rect 1843 -1497 1844 -1496
rect 324 -1499 325 -1498
rect 611 -1499 612 -1498
rect 1045 -1499 1046 -1498
rect 1108 -1499 1109 -1498
rect 1395 -1499 1396 -1498
rect 1409 -1499 1410 -1498
rect 1626 -1499 1627 -1498
rect 1661 -1499 1662 -1498
rect 1843 -1499 1844 -1498
rect 1906 -1499 1907 -1498
rect 583 -1501 584 -1500
rect 611 -1501 612 -1500
rect 695 -1501 696 -1500
rect 1045 -1501 1046 -1500
rect 1409 -1501 1410 -1500
rect 1528 -1501 1529 -1500
rect 1661 -1501 1662 -1500
rect 1703 -1501 1704 -1500
rect 1745 -1501 1746 -1500
rect 1906 -1501 1907 -1500
rect 30 -1503 31 -1502
rect 583 -1503 584 -1502
rect 639 -1503 640 -1502
rect 1528 -1503 1529 -1502
rect 1703 -1503 1704 -1502
rect 1738 -1503 1739 -1502
rect 1745 -1503 1746 -1502
rect 1808 -1503 1809 -1502
rect 30 -1505 31 -1504
rect 527 -1505 528 -1504
rect 1416 -1505 1417 -1504
rect 1808 -1505 1809 -1504
rect 100 -1507 101 -1506
rect 527 -1507 528 -1506
rect 1416 -1507 1417 -1506
rect 1437 -1507 1438 -1506
rect 1710 -1507 1711 -1506
rect 1738 -1507 1739 -1506
rect 100 -1509 101 -1508
rect 198 -1509 199 -1508
rect 233 -1509 234 -1508
rect 695 -1509 696 -1508
rect 1437 -1509 1438 -1508
rect 1458 -1509 1459 -1508
rect 72 -1511 73 -1510
rect 233 -1511 234 -1510
rect 576 -1511 577 -1510
rect 1710 -1511 1711 -1510
rect 198 -1513 199 -1512
rect 1171 -1513 1172 -1512
rect 1458 -1513 1459 -1512
rect 1465 -1513 1466 -1512
rect 576 -1515 577 -1514
rect 961 -1515 962 -1514
rect 1465 -1515 1466 -1514
rect 1479 -1515 1480 -1514
rect 1318 -1517 1319 -1516
rect 1479 -1517 1480 -1516
rect 1318 -1519 1319 -1518
rect 1346 -1519 1347 -1518
rect 1346 -1521 1347 -1520
rect 2319 -1521 2320 -1520
rect 2319 -1523 2320 -1522
rect 2403 -1523 2404 -1522
rect 1678 -1525 1679 -1524
rect 2403 -1525 2404 -1524
rect 16 -1536 17 -1535
rect 89 -1536 90 -1535
rect 93 -1536 94 -1535
rect 208 -1536 209 -1535
rect 229 -1536 230 -1535
rect 1710 -1536 1711 -1535
rect 2389 -1536 2390 -1535
rect 2427 -1536 2428 -1535
rect 2431 -1536 2432 -1535
rect 2434 -1536 2435 -1535
rect 23 -1538 24 -1537
rect 499 -1538 500 -1537
rect 583 -1538 584 -1537
rect 793 -1538 794 -1537
rect 807 -1538 808 -1537
rect 1332 -1538 1333 -1537
rect 1360 -1538 1361 -1537
rect 1440 -1538 1441 -1537
rect 1479 -1538 1480 -1537
rect 1976 -1538 1977 -1537
rect 2284 -1538 2285 -1537
rect 2389 -1538 2390 -1537
rect 23 -1540 24 -1539
rect 628 -1540 629 -1539
rect 642 -1540 643 -1539
rect 709 -1540 710 -1539
rect 719 -1540 720 -1539
rect 2305 -1540 2306 -1539
rect 40 -1542 41 -1541
rect 828 -1542 829 -1541
rect 859 -1542 860 -1541
rect 1493 -1542 1494 -1541
rect 1496 -1542 1497 -1541
rect 2536 -1542 2537 -1541
rect 44 -1544 45 -1543
rect 54 -1544 55 -1543
rect 72 -1544 73 -1543
rect 936 -1544 937 -1543
rect 943 -1544 944 -1543
rect 1640 -1544 1641 -1543
rect 1710 -1544 1711 -1543
rect 1822 -1544 1823 -1543
rect 1976 -1544 1977 -1543
rect 2088 -1544 2089 -1543
rect 2284 -1544 2285 -1543
rect 2417 -1544 2418 -1543
rect 44 -1546 45 -1545
rect 100 -1546 101 -1545
rect 107 -1546 108 -1545
rect 810 -1546 811 -1545
rect 821 -1546 822 -1545
rect 2032 -1546 2033 -1545
rect 2305 -1546 2306 -1545
rect 2438 -1546 2439 -1545
rect 47 -1548 48 -1547
rect 422 -1548 423 -1547
rect 481 -1548 482 -1547
rect 527 -1548 528 -1547
rect 583 -1548 584 -1547
rect 660 -1548 661 -1547
rect 691 -1548 692 -1547
rect 814 -1548 815 -1547
rect 821 -1548 822 -1547
rect 1143 -1548 1144 -1547
rect 1150 -1548 1151 -1547
rect 1584 -1548 1585 -1547
rect 1822 -1548 1823 -1547
rect 1906 -1548 1907 -1547
rect 1990 -1548 1991 -1547
rect 2088 -1548 2089 -1547
rect 2340 -1548 2341 -1547
rect 2438 -1548 2439 -1547
rect 30 -1550 31 -1549
rect 422 -1550 423 -1549
rect 527 -1550 528 -1549
rect 779 -1550 780 -1549
rect 793 -1550 794 -1549
rect 989 -1550 990 -1549
rect 1076 -1550 1077 -1549
rect 2403 -1550 2404 -1549
rect 30 -1552 31 -1551
rect 282 -1552 283 -1551
rect 366 -1552 367 -1551
rect 499 -1552 500 -1551
rect 590 -1552 591 -1551
rect 604 -1552 605 -1551
rect 625 -1552 626 -1551
rect 2053 -1552 2054 -1551
rect 2403 -1552 2404 -1551
rect 2515 -1552 2516 -1551
rect 51 -1554 52 -1553
rect 303 -1554 304 -1553
rect 366 -1554 367 -1553
rect 408 -1554 409 -1553
rect 590 -1554 591 -1553
rect 618 -1554 619 -1553
rect 625 -1554 626 -1553
rect 849 -1554 850 -1553
rect 880 -1554 881 -1553
rect 1514 -1554 1515 -1553
rect 1538 -1554 1539 -1553
rect 2123 -1554 2124 -1553
rect 51 -1556 52 -1555
rect 65 -1556 66 -1555
rect 72 -1556 73 -1555
rect 261 -1556 262 -1555
rect 268 -1556 269 -1555
rect 796 -1556 797 -1555
rect 814 -1556 815 -1555
rect 1038 -1556 1039 -1555
rect 1090 -1556 1091 -1555
rect 2410 -1556 2411 -1555
rect 2 -1558 3 -1557
rect 261 -1558 262 -1557
rect 268 -1558 269 -1557
rect 723 -1558 724 -1557
rect 730 -1558 731 -1557
rect 1020 -1558 1021 -1557
rect 1038 -1558 1039 -1557
rect 1220 -1558 1221 -1557
rect 1248 -1558 1249 -1557
rect 2347 -1558 2348 -1557
rect 65 -1560 66 -1559
rect 429 -1560 430 -1559
rect 604 -1560 605 -1559
rect 1206 -1560 1207 -1559
rect 1220 -1560 1221 -1559
rect 1311 -1560 1312 -1559
rect 1332 -1560 1333 -1559
rect 1605 -1560 1606 -1559
rect 1878 -1560 1879 -1559
rect 2053 -1560 2054 -1559
rect 2123 -1560 2124 -1559
rect 2242 -1560 2243 -1559
rect 2347 -1560 2348 -1559
rect 2473 -1560 2474 -1559
rect 79 -1562 80 -1561
rect 709 -1562 710 -1561
rect 723 -1562 724 -1561
rect 1066 -1562 1067 -1561
rect 1129 -1562 1130 -1561
rect 1206 -1562 1207 -1561
rect 1248 -1562 1249 -1561
rect 1395 -1562 1396 -1561
rect 1402 -1562 1403 -1561
rect 2417 -1562 2418 -1561
rect 79 -1564 80 -1563
rect 226 -1564 227 -1563
rect 233 -1564 234 -1563
rect 520 -1564 521 -1563
rect 646 -1564 647 -1563
rect 660 -1564 661 -1563
rect 698 -1564 699 -1563
rect 2340 -1564 2341 -1563
rect 100 -1566 101 -1565
rect 471 -1566 472 -1565
rect 520 -1566 521 -1565
rect 681 -1566 682 -1565
rect 702 -1566 703 -1565
rect 884 -1566 885 -1565
rect 887 -1566 888 -1565
rect 1024 -1566 1025 -1565
rect 1066 -1566 1067 -1565
rect 1171 -1566 1172 -1565
rect 1192 -1566 1193 -1565
rect 1251 -1566 1252 -1565
rect 1255 -1566 1256 -1565
rect 1297 -1566 1298 -1565
rect 1311 -1566 1312 -1565
rect 1458 -1566 1459 -1565
rect 1479 -1566 1480 -1565
rect 1521 -1566 1522 -1565
rect 1584 -1566 1585 -1565
rect 1675 -1566 1676 -1565
rect 1878 -1566 1879 -1565
rect 1969 -1566 1970 -1565
rect 1990 -1566 1991 -1565
rect 2060 -1566 2061 -1565
rect 2095 -1566 2096 -1565
rect 2242 -1566 2243 -1565
rect 37 -1568 38 -1567
rect 1024 -1568 1025 -1567
rect 1111 -1568 1112 -1567
rect 1675 -1568 1676 -1567
rect 1906 -1568 1907 -1567
rect 2018 -1568 2019 -1567
rect 2032 -1568 2033 -1567
rect 2144 -1568 2145 -1567
rect 37 -1570 38 -1569
rect 1612 -1570 1613 -1569
rect 1955 -1570 1956 -1569
rect 2018 -1570 2019 -1569
rect 2095 -1570 2096 -1569
rect 2214 -1570 2215 -1569
rect 121 -1572 122 -1571
rect 460 -1572 461 -1571
rect 471 -1572 472 -1571
rect 506 -1572 507 -1571
rect 534 -1572 535 -1571
rect 681 -1572 682 -1571
rect 702 -1572 703 -1571
rect 751 -1572 752 -1571
rect 779 -1572 780 -1571
rect 870 -1572 871 -1571
rect 898 -1572 899 -1571
rect 940 -1572 941 -1571
rect 961 -1572 962 -1571
rect 2172 -1572 2173 -1571
rect 2214 -1572 2215 -1571
rect 2326 -1572 2327 -1571
rect 114 -1574 115 -1573
rect 751 -1574 752 -1573
rect 824 -1574 825 -1573
rect 877 -1574 878 -1573
rect 898 -1574 899 -1573
rect 1010 -1574 1011 -1573
rect 1129 -1574 1130 -1573
rect 1234 -1574 1235 -1573
rect 1283 -1574 1284 -1573
rect 1304 -1574 1305 -1573
rect 1360 -1574 1361 -1573
rect 1864 -1574 1865 -1573
rect 1955 -1574 1956 -1573
rect 2067 -1574 2068 -1573
rect 2172 -1574 2173 -1573
rect 2291 -1574 2292 -1573
rect 2326 -1574 2327 -1573
rect 2445 -1574 2446 -1573
rect 114 -1576 115 -1575
rect 201 -1576 202 -1575
rect 212 -1576 213 -1575
rect 646 -1576 647 -1575
rect 737 -1576 738 -1575
rect 1269 -1576 1270 -1575
rect 1297 -1576 1298 -1575
rect 1353 -1576 1354 -1575
rect 1395 -1576 1396 -1575
rect 1829 -1576 1830 -1575
rect 1864 -1576 1865 -1575
rect 1941 -1576 1942 -1575
rect 1969 -1576 1970 -1575
rect 2081 -1576 2082 -1575
rect 2291 -1576 2292 -1575
rect 2361 -1576 2362 -1575
rect 2445 -1576 2446 -1575
rect 2543 -1576 2544 -1575
rect 121 -1578 122 -1577
rect 912 -1578 913 -1577
rect 964 -1578 965 -1577
rect 1402 -1578 1403 -1577
rect 1423 -1578 1424 -1577
rect 1801 -1578 1802 -1577
rect 1829 -1578 1830 -1577
rect 1962 -1578 1963 -1577
rect 2067 -1578 2068 -1577
rect 2158 -1578 2159 -1577
rect 2361 -1578 2362 -1577
rect 2487 -1578 2488 -1577
rect 128 -1580 129 -1579
rect 131 -1580 132 -1579
rect 198 -1580 199 -1579
rect 2494 -1580 2495 -1579
rect 128 -1582 129 -1581
rect 674 -1582 675 -1581
rect 849 -1582 850 -1581
rect 919 -1582 920 -1581
rect 989 -1582 990 -1581
rect 1122 -1582 1123 -1581
rect 1143 -1582 1144 -1581
rect 1178 -1582 1179 -1581
rect 1192 -1582 1193 -1581
rect 1325 -1582 1326 -1581
rect 1353 -1582 1354 -1581
rect 1549 -1582 1550 -1581
rect 1605 -1582 1606 -1581
rect 1633 -1582 1634 -1581
rect 1766 -1582 1767 -1581
rect 1941 -1582 1942 -1581
rect 1962 -1582 1963 -1581
rect 2074 -1582 2075 -1581
rect 2081 -1582 2082 -1581
rect 2193 -1582 2194 -1581
rect 2494 -1582 2495 -1581
rect 2522 -1582 2523 -1581
rect 184 -1584 185 -1583
rect 198 -1584 199 -1583
rect 212 -1584 213 -1583
rect 576 -1584 577 -1583
rect 593 -1584 594 -1583
rect 2144 -1584 2145 -1583
rect 2193 -1584 2194 -1583
rect 2298 -1584 2299 -1583
rect 177 -1586 178 -1585
rect 184 -1586 185 -1585
rect 219 -1586 220 -1585
rect 961 -1586 962 -1585
rect 1122 -1586 1123 -1585
rect 1811 -1586 1812 -1585
rect 2074 -1586 2075 -1585
rect 2165 -1586 2166 -1585
rect 2298 -1586 2299 -1585
rect 2424 -1586 2425 -1585
rect 135 -1588 136 -1587
rect 219 -1588 220 -1587
rect 226 -1588 227 -1587
rect 1010 -1588 1011 -1587
rect 1153 -1588 1154 -1587
rect 1269 -1588 1270 -1587
rect 1286 -1588 1287 -1587
rect 1801 -1588 1802 -1587
rect 2165 -1588 2166 -1587
rect 2270 -1588 2271 -1587
rect 135 -1590 136 -1589
rect 1052 -1590 1053 -1589
rect 1157 -1590 1158 -1589
rect 2221 -1590 2222 -1589
rect 2270 -1590 2271 -1589
rect 2312 -1590 2313 -1589
rect 233 -1592 234 -1591
rect 695 -1592 696 -1591
rect 800 -1592 801 -1591
rect 2424 -1592 2425 -1591
rect 236 -1594 237 -1593
rect 478 -1594 479 -1593
rect 506 -1594 507 -1593
rect 541 -1594 542 -1593
rect 667 -1594 668 -1593
rect 800 -1594 801 -1593
rect 870 -1594 871 -1593
rect 1045 -1594 1046 -1593
rect 1157 -1594 1158 -1593
rect 1374 -1594 1375 -1593
rect 1423 -1594 1424 -1593
rect 1619 -1594 1620 -1593
rect 1633 -1594 1634 -1593
rect 1738 -1594 1739 -1593
rect 1766 -1594 1767 -1593
rect 1920 -1594 1921 -1593
rect 2221 -1594 2222 -1593
rect 2277 -1594 2278 -1593
rect 2312 -1594 2313 -1593
rect 2382 -1594 2383 -1593
rect 240 -1596 241 -1595
rect 1017 -1596 1018 -1595
rect 1045 -1596 1046 -1595
rect 1108 -1596 1109 -1595
rect 1160 -1596 1161 -1595
rect 1290 -1596 1291 -1595
rect 1304 -1596 1305 -1595
rect 1437 -1596 1438 -1595
rect 1458 -1596 1459 -1595
rect 1773 -1596 1774 -1595
rect 2277 -1596 2278 -1595
rect 2396 -1596 2397 -1595
rect 156 -1598 157 -1597
rect 240 -1598 241 -1597
rect 247 -1598 248 -1597
rect 408 -1598 409 -1597
rect 415 -1598 416 -1597
rect 737 -1598 738 -1597
rect 828 -1598 829 -1597
rect 1108 -1598 1109 -1597
rect 1171 -1598 1172 -1597
rect 1416 -1598 1417 -1597
rect 1486 -1598 1487 -1597
rect 1563 -1598 1564 -1597
rect 1612 -1598 1613 -1597
rect 1794 -1598 1795 -1597
rect 2382 -1598 2383 -1597
rect 2508 -1598 2509 -1597
rect 156 -1600 157 -1599
rect 170 -1600 171 -1599
rect 275 -1600 276 -1599
rect 453 -1600 454 -1599
rect 464 -1600 465 -1599
rect 534 -1600 535 -1599
rect 667 -1600 668 -1599
rect 933 -1600 934 -1599
rect 954 -1600 955 -1599
rect 1290 -1600 1291 -1599
rect 1325 -1600 1326 -1599
rect 1444 -1600 1445 -1599
rect 1489 -1600 1490 -1599
rect 2235 -1600 2236 -1599
rect 2396 -1600 2397 -1599
rect 2480 -1600 2481 -1599
rect 117 -1602 118 -1601
rect 464 -1602 465 -1601
rect 478 -1602 479 -1601
rect 492 -1602 493 -1601
rect 516 -1602 517 -1601
rect 1052 -1602 1053 -1601
rect 1178 -1602 1179 -1601
rect 1213 -1602 1214 -1601
rect 1265 -1602 1266 -1601
rect 1773 -1602 1774 -1601
rect 1794 -1602 1795 -1601
rect 1892 -1602 1893 -1601
rect 2235 -1602 2236 -1601
rect 2354 -1602 2355 -1601
rect 149 -1604 150 -1603
rect 492 -1604 493 -1603
rect 674 -1604 675 -1603
rect 891 -1604 892 -1603
rect 905 -1604 906 -1603
rect 1451 -1604 1452 -1603
rect 1493 -1604 1494 -1603
rect 1619 -1604 1620 -1603
rect 1738 -1604 1739 -1603
rect 1787 -1604 1788 -1603
rect 1892 -1604 1893 -1603
rect 1997 -1604 1998 -1603
rect 2207 -1604 2208 -1603
rect 2354 -1604 2355 -1603
rect 86 -1606 87 -1605
rect 149 -1606 150 -1605
rect 170 -1606 171 -1605
rect 254 -1606 255 -1605
rect 275 -1606 276 -1605
rect 296 -1606 297 -1605
rect 303 -1606 304 -1605
rect 401 -1606 402 -1605
rect 429 -1606 430 -1605
rect 443 -1606 444 -1605
rect 695 -1606 696 -1605
rect 772 -1606 773 -1605
rect 891 -1606 892 -1605
rect 975 -1606 976 -1605
rect 982 -1606 983 -1605
rect 1017 -1606 1018 -1605
rect 1213 -1606 1214 -1605
rect 1752 -1606 1753 -1605
rect 1759 -1606 1760 -1605
rect 1920 -1606 1921 -1605
rect 1983 -1606 1984 -1605
rect 2207 -1606 2208 -1605
rect 86 -1608 87 -1607
rect 142 -1608 143 -1607
rect 250 -1608 251 -1607
rect 1451 -1608 1452 -1607
rect 1503 -1608 1504 -1607
rect 2466 -1608 2467 -1607
rect 142 -1610 143 -1609
rect 642 -1610 643 -1609
rect 772 -1610 773 -1609
rect 842 -1610 843 -1609
rect 905 -1610 906 -1609
rect 1381 -1610 1382 -1609
rect 1416 -1610 1417 -1609
rect 1465 -1610 1466 -1609
rect 1507 -1610 1508 -1609
rect 1640 -1610 1641 -1609
rect 1752 -1610 1753 -1609
rect 1871 -1610 1872 -1609
rect 1997 -1610 1998 -1609
rect 2102 -1610 2103 -1609
rect 110 -1612 111 -1611
rect 1465 -1612 1466 -1611
rect 1514 -1612 1515 -1611
rect 1682 -1612 1683 -1611
rect 1759 -1612 1760 -1611
rect 1899 -1612 1900 -1611
rect 2102 -1612 2103 -1611
rect 2319 -1612 2320 -1611
rect 205 -1614 206 -1613
rect 1381 -1614 1382 -1613
rect 1444 -1614 1445 -1613
rect 1598 -1614 1599 -1613
rect 1787 -1614 1788 -1613
rect 2109 -1614 2110 -1613
rect 2319 -1614 2320 -1613
rect 2529 -1614 2530 -1613
rect 205 -1616 206 -1615
rect 653 -1616 654 -1615
rect 842 -1616 843 -1615
rect 926 -1616 927 -1615
rect 933 -1616 934 -1615
rect 1115 -1616 1116 -1615
rect 1234 -1616 1235 -1615
rect 1507 -1616 1508 -1615
rect 1531 -1616 1532 -1615
rect 2158 -1616 2159 -1615
rect 254 -1618 255 -1617
rect 1153 -1618 1154 -1617
rect 1276 -1618 1277 -1617
rect 1437 -1618 1438 -1617
rect 1549 -1618 1550 -1617
rect 1668 -1618 1669 -1617
rect 1815 -1618 1816 -1617
rect 1983 -1618 1984 -1617
rect 282 -1620 283 -1619
rect 373 -1620 374 -1619
rect 387 -1620 388 -1619
rect 807 -1620 808 -1619
rect 912 -1620 913 -1619
rect 1570 -1620 1571 -1619
rect 1668 -1620 1669 -1619
rect 1780 -1620 1781 -1619
rect 1871 -1620 1872 -1619
rect 1948 -1620 1949 -1619
rect 96 -1622 97 -1621
rect 1570 -1622 1571 -1621
rect 1899 -1622 1900 -1621
rect 2011 -1622 2012 -1621
rect 296 -1624 297 -1623
rect 611 -1624 612 -1623
rect 919 -1624 920 -1623
rect 1031 -1624 1032 -1623
rect 1034 -1624 1035 -1623
rect 1598 -1624 1599 -1623
rect 1927 -1624 1928 -1623
rect 2109 -1624 2110 -1623
rect 338 -1626 339 -1625
rect 401 -1626 402 -1625
rect 436 -1626 437 -1625
rect 940 -1626 941 -1625
rect 954 -1626 955 -1625
rect 1059 -1626 1060 -1625
rect 1115 -1626 1116 -1625
rect 1136 -1626 1137 -1625
rect 1258 -1626 1259 -1625
rect 1815 -1626 1816 -1625
rect 1927 -1626 1928 -1625
rect 2025 -1626 2026 -1625
rect 338 -1628 339 -1627
rect 345 -1628 346 -1627
rect 352 -1628 353 -1627
rect 415 -1628 416 -1627
rect 436 -1628 437 -1627
rect 1500 -1628 1501 -1627
rect 1563 -1628 1564 -1627
rect 1696 -1628 1697 -1627
rect 1948 -1628 1949 -1627
rect 2046 -1628 2047 -1627
rect 289 -1630 290 -1629
rect 352 -1630 353 -1629
rect 373 -1630 374 -1629
rect 457 -1630 458 -1629
rect 562 -1630 563 -1629
rect 611 -1630 612 -1629
rect 926 -1630 927 -1629
rect 1073 -1630 1074 -1629
rect 1136 -1630 1137 -1629
rect 1318 -1630 1319 -1629
rect 1349 -1630 1350 -1629
rect 1682 -1630 1683 -1629
rect 1689 -1630 1690 -1629
rect 1696 -1630 1697 -1629
rect 2004 -1630 2005 -1629
rect 2011 -1630 2012 -1629
rect 2025 -1630 2026 -1629
rect 2130 -1630 2131 -1629
rect 191 -1632 192 -1631
rect 289 -1632 290 -1631
rect 317 -1632 318 -1631
rect 345 -1632 346 -1631
rect 387 -1632 388 -1631
rect 1003 -1632 1004 -1631
rect 1059 -1632 1060 -1631
rect 1101 -1632 1102 -1631
rect 1262 -1632 1263 -1631
rect 1780 -1632 1781 -1631
rect 2004 -1632 2005 -1631
rect 2116 -1632 2117 -1631
rect 2130 -1632 2131 -1631
rect 2249 -1632 2250 -1631
rect 191 -1634 192 -1633
rect 618 -1634 619 -1633
rect 975 -1634 976 -1633
rect 1080 -1634 1081 -1633
rect 1101 -1634 1102 -1633
rect 1227 -1634 1228 -1633
rect 1276 -1634 1277 -1633
rect 1521 -1634 1522 -1633
rect 1689 -1634 1690 -1633
rect 1808 -1634 1809 -1633
rect 2046 -1634 2047 -1633
rect 2137 -1634 2138 -1633
rect 2249 -1634 2250 -1633
rect 2459 -1634 2460 -1633
rect 194 -1636 195 -1635
rect 1262 -1636 1263 -1635
rect 1318 -1636 1319 -1635
rect 1654 -1636 1655 -1635
rect 1808 -1636 1809 -1635
rect 2179 -1636 2180 -1635
rect 317 -1638 318 -1637
rect 359 -1638 360 -1637
rect 394 -1638 395 -1637
rect 639 -1638 640 -1637
rect 968 -1638 969 -1637
rect 1227 -1638 1228 -1637
rect 1293 -1638 1294 -1637
rect 1654 -1638 1655 -1637
rect 2116 -1638 2117 -1637
rect 2228 -1638 2229 -1637
rect 324 -1640 325 -1639
rect 457 -1640 458 -1639
rect 548 -1640 549 -1639
rect 562 -1640 563 -1639
rect 639 -1640 640 -1639
rect 2550 -1640 2551 -1639
rect 324 -1642 325 -1641
rect 555 -1642 556 -1641
rect 856 -1642 857 -1641
rect 968 -1642 969 -1641
rect 982 -1642 983 -1641
rect 1164 -1642 1165 -1641
rect 1374 -1642 1375 -1641
rect 1535 -1642 1536 -1641
rect 2137 -1642 2138 -1641
rect 2375 -1642 2376 -1641
rect 331 -1644 332 -1643
rect 359 -1644 360 -1643
rect 394 -1644 395 -1643
rect 632 -1644 633 -1643
rect 653 -1644 654 -1643
rect 856 -1644 857 -1643
rect 1003 -1644 1004 -1643
rect 1185 -1644 1186 -1643
rect 1500 -1644 1501 -1643
rect 1626 -1644 1627 -1643
rect 2200 -1644 2201 -1643
rect 2375 -1644 2376 -1643
rect 331 -1646 332 -1645
rect 485 -1646 486 -1645
rect 548 -1646 549 -1645
rect 758 -1646 759 -1645
rect 1073 -1646 1074 -1645
rect 2186 -1646 2187 -1645
rect 2200 -1646 2201 -1645
rect 2263 -1646 2264 -1645
rect 180 -1648 181 -1647
rect 2186 -1648 2187 -1647
rect 2228 -1648 2229 -1647
rect 2333 -1648 2334 -1647
rect 443 -1650 444 -1649
rect 1346 -1650 1347 -1649
rect 1468 -1650 1469 -1649
rect 2263 -1650 2264 -1649
rect 2333 -1650 2334 -1649
rect 2452 -1650 2453 -1649
rect 450 -1652 451 -1651
rect 632 -1652 633 -1651
rect 758 -1652 759 -1651
rect 835 -1652 836 -1651
rect 996 -1652 997 -1651
rect 1346 -1652 1347 -1651
rect 1430 -1652 1431 -1651
rect 2452 -1652 2453 -1651
rect 450 -1654 451 -1653
rect 730 -1654 731 -1653
rect 765 -1654 766 -1653
rect 835 -1654 836 -1653
rect 1080 -1654 1081 -1653
rect 1199 -1654 1200 -1653
rect 1430 -1654 1431 -1653
rect 1556 -1654 1557 -1653
rect 1626 -1654 1627 -1653
rect 1731 -1654 1732 -1653
rect 485 -1656 486 -1655
rect 716 -1656 717 -1655
rect 765 -1656 766 -1655
rect 1087 -1656 1088 -1655
rect 1164 -1656 1165 -1655
rect 1367 -1656 1368 -1655
rect 1528 -1656 1529 -1655
rect 2179 -1656 2180 -1655
rect 513 -1658 514 -1657
rect 996 -1658 997 -1657
rect 1087 -1658 1088 -1657
rect 1363 -1658 1364 -1657
rect 1367 -1658 1368 -1657
rect 1472 -1658 1473 -1657
rect 1535 -1658 1536 -1657
rect 2060 -1658 2061 -1657
rect 513 -1660 514 -1659
rect 688 -1660 689 -1659
rect 786 -1660 787 -1659
rect 1199 -1660 1200 -1659
rect 1388 -1660 1389 -1659
rect 1528 -1660 1529 -1659
rect 1556 -1660 1557 -1659
rect 1724 -1660 1725 -1659
rect 131 -1662 132 -1661
rect 786 -1662 787 -1661
rect 866 -1662 867 -1661
rect 1731 -1662 1732 -1661
rect 555 -1664 556 -1663
rect 2441 -1664 2442 -1663
rect 569 -1666 570 -1665
rect 716 -1666 717 -1665
rect 1185 -1666 1186 -1665
rect 1241 -1666 1242 -1665
rect 1388 -1666 1389 -1665
rect 1542 -1666 1543 -1665
rect 1724 -1666 1725 -1665
rect 1850 -1666 1851 -1665
rect 569 -1668 570 -1667
rect 863 -1668 864 -1667
rect 1241 -1668 1242 -1667
rect 1339 -1668 1340 -1667
rect 1472 -1668 1473 -1667
rect 1661 -1668 1662 -1667
rect 1850 -1668 1851 -1667
rect 1934 -1668 1935 -1667
rect 688 -1670 689 -1669
rect 744 -1670 745 -1669
rect 863 -1670 864 -1669
rect 947 -1670 948 -1669
rect 1339 -1670 1340 -1669
rect 1409 -1670 1410 -1669
rect 1542 -1670 1543 -1669
rect 1647 -1670 1648 -1669
rect 1661 -1670 1662 -1669
rect 1745 -1670 1746 -1669
rect 1934 -1670 1935 -1669
rect 2039 -1670 2040 -1669
rect 9 -1672 10 -1671
rect 744 -1672 745 -1671
rect 947 -1672 948 -1671
rect 2557 -1672 2558 -1671
rect 93 -1674 94 -1673
rect 2039 -1674 2040 -1673
rect 1409 -1676 1410 -1675
rect 1591 -1676 1592 -1675
rect 1745 -1676 1746 -1675
rect 1857 -1676 1858 -1675
rect 1510 -1678 1511 -1677
rect 1857 -1678 1858 -1677
rect 1577 -1680 1578 -1679
rect 1647 -1680 1648 -1679
rect 1577 -1682 1578 -1681
rect 1703 -1682 1704 -1681
rect 1591 -1684 1592 -1683
rect 1717 -1684 1718 -1683
rect 1703 -1686 1704 -1685
rect 2410 -1686 2411 -1685
rect 1717 -1688 1718 -1687
rect 1843 -1688 1844 -1687
rect 1843 -1690 1844 -1689
rect 1913 -1690 1914 -1689
rect 1913 -1692 1914 -1691
rect 2151 -1692 2152 -1691
rect 2151 -1694 2152 -1693
rect 2256 -1694 2257 -1693
rect 2256 -1696 2257 -1695
rect 2368 -1696 2369 -1695
rect 2368 -1698 2369 -1697
rect 2501 -1698 2502 -1697
rect 2 -1709 3 -1708
rect 387 -1709 388 -1708
rect 429 -1709 430 -1708
rect 1538 -1709 1539 -1708
rect 1629 -1709 1630 -1708
rect 2046 -1709 2047 -1708
rect 2389 -1709 2390 -1708
rect 2438 -1709 2439 -1708
rect 2445 -1709 2446 -1708
rect 2459 -1709 2460 -1708
rect 2469 -1709 2470 -1708
rect 2494 -1709 2495 -1708
rect 9 -1711 10 -1710
rect 107 -1711 108 -1710
rect 142 -1711 143 -1710
rect 145 -1711 146 -1710
rect 187 -1711 188 -1710
rect 1265 -1711 1266 -1710
rect 1276 -1711 1277 -1710
rect 2410 -1711 2411 -1710
rect 16 -1713 17 -1712
rect 614 -1713 615 -1712
rect 649 -1713 650 -1712
rect 943 -1713 944 -1712
rect 1017 -1713 1018 -1712
rect 1605 -1713 1606 -1712
rect 1664 -1713 1665 -1712
rect 2312 -1713 2313 -1712
rect 2347 -1713 2348 -1712
rect 2410 -1713 2411 -1712
rect 16 -1715 17 -1714
rect 1003 -1715 1004 -1714
rect 1020 -1715 1021 -1714
rect 1192 -1715 1193 -1714
rect 1206 -1715 1207 -1714
rect 1290 -1715 1291 -1714
rect 1293 -1715 1294 -1714
rect 2270 -1715 2271 -1714
rect 2389 -1715 2390 -1714
rect 2473 -1715 2474 -1714
rect 30 -1717 31 -1716
rect 894 -1717 895 -1716
rect 989 -1717 990 -1716
rect 1017 -1717 1018 -1716
rect 1031 -1717 1032 -1716
rect 1402 -1717 1403 -1716
rect 1437 -1717 1438 -1716
rect 1738 -1717 1739 -1716
rect 1801 -1717 1802 -1716
rect 2476 -1717 2477 -1716
rect 30 -1719 31 -1718
rect 331 -1719 332 -1718
rect 446 -1719 447 -1718
rect 807 -1719 808 -1718
rect 821 -1719 822 -1718
rect 1073 -1719 1074 -1718
rect 1108 -1719 1109 -1718
rect 2417 -1719 2418 -1718
rect 37 -1721 38 -1720
rect 96 -1721 97 -1720
rect 107 -1721 108 -1720
rect 373 -1721 374 -1720
rect 394 -1721 395 -1720
rect 807 -1721 808 -1720
rect 821 -1721 822 -1720
rect 1363 -1721 1364 -1720
rect 1367 -1721 1368 -1720
rect 1402 -1721 1403 -1720
rect 1440 -1721 1441 -1720
rect 2291 -1721 2292 -1720
rect 2361 -1721 2362 -1720
rect 2417 -1721 2418 -1720
rect 37 -1723 38 -1722
rect 443 -1723 444 -1722
rect 457 -1723 458 -1722
rect 828 -1723 829 -1722
rect 835 -1723 836 -1722
rect 908 -1723 909 -1722
rect 961 -1723 962 -1722
rect 1031 -1723 1032 -1722
rect 1059 -1723 1060 -1722
rect 1062 -1723 1063 -1722
rect 1111 -1723 1112 -1722
rect 1885 -1723 1886 -1722
rect 1997 -1723 1998 -1722
rect 2046 -1723 2047 -1722
rect 2228 -1723 2229 -1722
rect 2291 -1723 2292 -1722
rect 2305 -1723 2306 -1722
rect 2361 -1723 2362 -1722
rect 47 -1725 48 -1724
rect 51 -1725 52 -1724
rect 65 -1725 66 -1724
rect 180 -1725 181 -1724
rect 194 -1725 195 -1724
rect 1101 -1725 1102 -1724
rect 1153 -1725 1154 -1724
rect 1696 -1725 1697 -1724
rect 1706 -1725 1707 -1724
rect 2375 -1725 2376 -1724
rect 51 -1727 52 -1726
rect 240 -1727 241 -1726
rect 247 -1727 248 -1726
rect 534 -1727 535 -1726
rect 548 -1727 549 -1726
rect 856 -1727 857 -1726
rect 870 -1727 871 -1726
rect 961 -1727 962 -1726
rect 989 -1727 990 -1726
rect 1010 -1727 1011 -1726
rect 1059 -1727 1060 -1726
rect 1409 -1727 1410 -1726
rect 1440 -1727 1441 -1726
rect 1703 -1727 1704 -1726
rect 1836 -1727 1837 -1726
rect 2434 -1727 2435 -1726
rect 58 -1729 59 -1728
rect 65 -1729 66 -1728
rect 86 -1729 87 -1728
rect 159 -1729 160 -1728
rect 198 -1729 199 -1728
rect 1150 -1729 1151 -1728
rect 1192 -1729 1193 -1728
rect 1283 -1729 1284 -1728
rect 1293 -1729 1294 -1728
rect 1444 -1729 1445 -1728
rect 1458 -1729 1459 -1728
rect 1997 -1729 1998 -1728
rect 2039 -1729 2040 -1728
rect 2042 -1729 2043 -1728
rect 2228 -1729 2229 -1728
rect 2319 -1729 2320 -1728
rect 58 -1731 59 -1730
rect 898 -1731 899 -1730
rect 957 -1731 958 -1730
rect 1444 -1731 1445 -1730
rect 1468 -1731 1469 -1730
rect 2396 -1731 2397 -1730
rect 86 -1733 87 -1732
rect 135 -1733 136 -1732
rect 142 -1733 143 -1732
rect 450 -1733 451 -1732
rect 460 -1733 461 -1732
rect 632 -1733 633 -1732
rect 653 -1733 654 -1732
rect 828 -1733 829 -1732
rect 870 -1733 871 -1732
rect 891 -1733 892 -1732
rect 1003 -1733 1004 -1732
rect 1094 -1733 1095 -1732
rect 1143 -1733 1144 -1732
rect 1150 -1733 1151 -1732
rect 1209 -1733 1210 -1732
rect 1374 -1733 1375 -1732
rect 1388 -1733 1389 -1732
rect 1458 -1733 1459 -1732
rect 1468 -1733 1469 -1732
rect 2319 -1733 2320 -1732
rect 44 -1735 45 -1734
rect 1374 -1735 1375 -1734
rect 1493 -1735 1494 -1734
rect 1647 -1735 1648 -1734
rect 1696 -1735 1697 -1734
rect 1941 -1735 1942 -1734
rect 2039 -1735 2040 -1734
rect 2137 -1735 2138 -1734
rect 2235 -1735 2236 -1734
rect 2305 -1735 2306 -1734
rect 93 -1737 94 -1736
rect 926 -1737 927 -1736
rect 1143 -1737 1144 -1736
rect 1181 -1737 1182 -1736
rect 1213 -1737 1214 -1736
rect 1307 -1737 1308 -1736
rect 1325 -1737 1326 -1736
rect 1367 -1737 1368 -1736
rect 1493 -1737 1494 -1736
rect 1591 -1737 1592 -1736
rect 1647 -1737 1648 -1736
rect 1808 -1737 1809 -1736
rect 1815 -1737 1816 -1736
rect 1836 -1737 1837 -1736
rect 1850 -1737 1851 -1736
rect 1885 -1737 1886 -1736
rect 1941 -1737 1942 -1736
rect 2158 -1737 2159 -1736
rect 2179 -1737 2180 -1736
rect 2235 -1737 2236 -1736
rect 2242 -1737 2243 -1736
rect 2270 -1737 2271 -1736
rect 2284 -1737 2285 -1736
rect 2375 -1737 2376 -1736
rect 93 -1739 94 -1738
rect 380 -1739 381 -1738
rect 429 -1739 430 -1738
rect 926 -1739 927 -1738
rect 1171 -1739 1172 -1738
rect 1325 -1739 1326 -1738
rect 1360 -1739 1361 -1738
rect 2207 -1739 2208 -1738
rect 2221 -1739 2222 -1738
rect 2284 -1739 2285 -1738
rect 135 -1741 136 -1740
rect 205 -1741 206 -1740
rect 212 -1741 213 -1740
rect 863 -1741 864 -1740
rect 884 -1741 885 -1740
rect 1073 -1741 1074 -1740
rect 1164 -1741 1165 -1740
rect 1171 -1741 1172 -1740
rect 1213 -1741 1214 -1740
rect 1241 -1741 1242 -1740
rect 1262 -1741 1263 -1740
rect 2018 -1741 2019 -1740
rect 2081 -1741 2082 -1740
rect 2137 -1741 2138 -1740
rect 2151 -1741 2152 -1740
rect 2221 -1741 2222 -1740
rect 2263 -1741 2264 -1740
rect 2347 -1741 2348 -1740
rect 100 -1743 101 -1742
rect 205 -1743 206 -1742
rect 212 -1743 213 -1742
rect 758 -1743 759 -1742
rect 793 -1743 794 -1742
rect 1010 -1743 1011 -1742
rect 1227 -1743 1228 -1742
rect 1388 -1743 1389 -1742
rect 1510 -1743 1511 -1742
rect 2200 -1743 2201 -1742
rect 198 -1745 199 -1744
rect 366 -1745 367 -1744
rect 373 -1745 374 -1744
rect 565 -1745 566 -1744
rect 579 -1745 580 -1744
rect 1738 -1745 1739 -1744
rect 1745 -1745 1746 -1744
rect 2242 -1745 2243 -1744
rect 226 -1747 227 -1746
rect 912 -1747 913 -1746
rect 940 -1747 941 -1746
rect 1164 -1747 1165 -1746
rect 1185 -1747 1186 -1746
rect 1227 -1747 1228 -1746
rect 1241 -1747 1242 -1746
rect 1311 -1747 1312 -1746
rect 1353 -1747 1354 -1746
rect 1360 -1747 1361 -1746
rect 1528 -1747 1529 -1746
rect 2403 -1747 2404 -1746
rect 229 -1749 230 -1748
rect 1094 -1749 1095 -1748
rect 1248 -1749 1249 -1748
rect 1262 -1749 1263 -1748
rect 1283 -1749 1284 -1748
rect 1521 -1749 1522 -1748
rect 1528 -1749 1529 -1748
rect 1542 -1749 1543 -1748
rect 1556 -1749 1557 -1748
rect 1605 -1749 1606 -1748
rect 1724 -1749 1725 -1748
rect 1745 -1749 1746 -1748
rect 1759 -1749 1760 -1748
rect 2018 -1749 2019 -1748
rect 2102 -1749 2103 -1748
rect 2263 -1749 2264 -1748
rect 2333 -1749 2334 -1748
rect 2403 -1749 2404 -1748
rect 124 -1751 125 -1750
rect 1521 -1751 1522 -1750
rect 1531 -1751 1532 -1750
rect 2312 -1751 2313 -1750
rect 236 -1753 237 -1752
rect 954 -1753 955 -1752
rect 1052 -1753 1053 -1752
rect 1185 -1753 1186 -1752
rect 1297 -1753 1298 -1752
rect 1409 -1753 1410 -1752
rect 1535 -1753 1536 -1752
rect 2088 -1753 2089 -1752
rect 2130 -1753 2131 -1752
rect 2207 -1753 2208 -1752
rect 240 -1755 241 -1754
rect 1076 -1755 1077 -1754
rect 1234 -1755 1235 -1754
rect 1297 -1755 1298 -1754
rect 1304 -1755 1305 -1754
rect 1353 -1755 1354 -1754
rect 1535 -1755 1536 -1754
rect 1612 -1755 1613 -1754
rect 1619 -1755 1620 -1754
rect 1759 -1755 1760 -1754
rect 1773 -1755 1774 -1754
rect 1815 -1755 1816 -1754
rect 1850 -1755 1851 -1754
rect 2354 -1755 2355 -1754
rect 289 -1757 290 -1756
rect 698 -1757 699 -1756
rect 716 -1757 717 -1756
rect 2158 -1757 2159 -1756
rect 2165 -1757 2166 -1756
rect 2200 -1757 2201 -1756
rect 2298 -1757 2299 -1756
rect 2354 -1757 2355 -1756
rect 289 -1759 290 -1758
rect 324 -1759 325 -1758
rect 331 -1759 332 -1758
rect 513 -1759 514 -1758
rect 520 -1759 521 -1758
rect 639 -1759 640 -1758
rect 653 -1759 654 -1758
rect 737 -1759 738 -1758
rect 744 -1759 745 -1758
rect 1052 -1759 1053 -1758
rect 1157 -1759 1158 -1758
rect 1234 -1759 1235 -1758
rect 1290 -1759 1291 -1758
rect 2165 -1759 2166 -1758
rect 2179 -1759 2180 -1758
rect 2382 -1759 2383 -1758
rect 324 -1761 325 -1760
rect 590 -1761 591 -1760
rect 618 -1761 619 -1760
rect 1108 -1761 1109 -1760
rect 1115 -1761 1116 -1760
rect 1157 -1761 1158 -1760
rect 1304 -1761 1305 -1760
rect 1801 -1761 1802 -1760
rect 1808 -1761 1809 -1760
rect 1913 -1761 1914 -1760
rect 2053 -1761 2054 -1760
rect 2102 -1761 2103 -1760
rect 2151 -1761 2152 -1760
rect 2424 -1761 2425 -1760
rect 121 -1763 122 -1762
rect 618 -1763 619 -1762
rect 660 -1763 661 -1762
rect 737 -1763 738 -1762
rect 744 -1763 745 -1762
rect 905 -1763 906 -1762
rect 912 -1763 913 -1762
rect 1045 -1763 1046 -1762
rect 1496 -1763 1497 -1762
rect 2298 -1763 2299 -1762
rect 2340 -1763 2341 -1762
rect 2382 -1763 2383 -1762
rect 79 -1765 80 -1764
rect 121 -1765 122 -1764
rect 345 -1765 346 -1764
rect 366 -1765 367 -1764
rect 387 -1765 388 -1764
rect 513 -1765 514 -1764
rect 520 -1765 521 -1764
rect 611 -1765 612 -1764
rect 667 -1765 668 -1764
rect 835 -1765 836 -1764
rect 849 -1765 850 -1764
rect 884 -1765 885 -1764
rect 891 -1765 892 -1764
rect 1983 -1765 1984 -1764
rect 2004 -1765 2005 -1764
rect 2340 -1765 2341 -1764
rect 79 -1767 80 -1766
rect 268 -1767 269 -1766
rect 275 -1767 276 -1766
rect 345 -1767 346 -1766
rect 352 -1767 353 -1766
rect 380 -1767 381 -1766
rect 436 -1767 437 -1766
rect 534 -1767 535 -1766
rect 548 -1767 549 -1766
rect 947 -1767 948 -1766
rect 954 -1767 955 -1766
rect 1279 -1767 1280 -1766
rect 1556 -1767 1557 -1766
rect 1626 -1767 1627 -1766
rect 1724 -1767 1725 -1766
rect 1871 -1767 1872 -1766
rect 1934 -1767 1935 -1766
rect 1983 -1767 1984 -1766
rect 2025 -1767 2026 -1766
rect 2053 -1767 2054 -1766
rect 2249 -1767 2250 -1766
rect 2424 -1767 2425 -1766
rect 149 -1769 150 -1768
rect 436 -1769 437 -1768
rect 443 -1769 444 -1768
rect 1542 -1769 1543 -1768
rect 1563 -1769 1564 -1768
rect 1591 -1769 1592 -1768
rect 1598 -1769 1599 -1768
rect 1612 -1769 1613 -1768
rect 1619 -1769 1620 -1768
rect 1717 -1769 1718 -1768
rect 1773 -1769 1774 -1768
rect 1899 -1769 1900 -1768
rect 1955 -1769 1956 -1768
rect 2004 -1769 2005 -1768
rect 2042 -1769 2043 -1768
rect 2081 -1769 2082 -1768
rect 149 -1771 150 -1770
rect 184 -1771 185 -1770
rect 268 -1771 269 -1770
rect 338 -1771 339 -1770
rect 352 -1771 353 -1770
rect 408 -1771 409 -1770
rect 481 -1771 482 -1770
rect 1311 -1771 1312 -1770
rect 1465 -1771 1466 -1770
rect 1934 -1771 1935 -1770
rect 1969 -1771 1970 -1770
rect 2249 -1771 2250 -1770
rect 114 -1773 115 -1772
rect 338 -1773 339 -1772
rect 359 -1773 360 -1772
rect 394 -1773 395 -1772
rect 408 -1773 409 -1772
rect 415 -1773 416 -1772
rect 492 -1773 493 -1772
rect 660 -1773 661 -1772
rect 667 -1773 668 -1772
rect 681 -1773 682 -1772
rect 695 -1773 696 -1772
rect 2445 -1773 2446 -1772
rect 114 -1775 115 -1774
rect 1423 -1775 1424 -1774
rect 1465 -1775 1466 -1774
rect 1731 -1775 1732 -1774
rect 1787 -1775 1788 -1774
rect 2333 -1775 2334 -1774
rect 275 -1777 276 -1776
rect 282 -1777 283 -1776
rect 317 -1777 318 -1776
rect 359 -1777 360 -1776
rect 415 -1777 416 -1776
rect 597 -1777 598 -1776
rect 646 -1777 647 -1776
rect 947 -1777 948 -1776
rect 968 -1777 969 -1776
rect 1913 -1777 1914 -1776
rect 1927 -1777 1928 -1776
rect 1969 -1777 1970 -1776
rect 1976 -1777 1977 -1776
rect 2025 -1777 2026 -1776
rect 282 -1779 283 -1778
rect 569 -1779 570 -1778
rect 590 -1779 591 -1778
rect 688 -1779 689 -1778
rect 695 -1779 696 -1778
rect 730 -1779 731 -1778
rect 733 -1779 734 -1778
rect 996 -1779 997 -1778
rect 1045 -1779 1046 -1778
rect 1066 -1779 1067 -1778
rect 1269 -1779 1270 -1778
rect 1423 -1779 1424 -1778
rect 1479 -1779 1480 -1778
rect 1787 -1779 1788 -1778
rect 1843 -1779 1844 -1778
rect 1871 -1779 1872 -1778
rect 1878 -1779 1879 -1778
rect 1955 -1779 1956 -1778
rect 1976 -1779 1977 -1778
rect 2172 -1779 2173 -1778
rect 219 -1781 220 -1780
rect 1269 -1781 1270 -1780
rect 1276 -1781 1277 -1780
rect 1878 -1781 1879 -1780
rect 2123 -1781 2124 -1780
rect 2172 -1781 2173 -1780
rect 191 -1783 192 -1782
rect 219 -1783 220 -1782
rect 296 -1783 297 -1782
rect 597 -1783 598 -1782
rect 674 -1783 675 -1782
rect 856 -1783 857 -1782
rect 863 -1783 864 -1782
rect 1507 -1783 1508 -1782
rect 1563 -1783 1564 -1782
rect 1794 -1783 1795 -1782
rect 1857 -1783 1858 -1782
rect 1899 -1783 1900 -1782
rect 2074 -1783 2075 -1782
rect 2123 -1783 2124 -1782
rect 191 -1785 192 -1784
rect 485 -1785 486 -1784
rect 492 -1785 493 -1784
rect 506 -1785 507 -1784
rect 516 -1785 517 -1784
rect 1066 -1785 1067 -1784
rect 1472 -1785 1473 -1784
rect 1843 -1785 1844 -1784
rect 2074 -1785 2075 -1784
rect 2326 -1785 2327 -1784
rect 261 -1787 262 -1786
rect 296 -1787 297 -1786
rect 310 -1787 311 -1786
rect 317 -1787 318 -1786
rect 453 -1787 454 -1786
rect 688 -1787 689 -1786
rect 716 -1787 717 -1786
rect 751 -1787 752 -1786
rect 758 -1787 759 -1786
rect 982 -1787 983 -1786
rect 1430 -1787 1431 -1786
rect 1472 -1787 1473 -1786
rect 1479 -1787 1480 -1786
rect 1486 -1787 1487 -1786
rect 1507 -1787 1508 -1786
rect 1990 -1787 1991 -1786
rect 2116 -1787 2117 -1786
rect 2326 -1787 2327 -1786
rect 250 -1789 251 -1788
rect 261 -1789 262 -1788
rect 310 -1789 311 -1788
rect 527 -1789 528 -1788
rect 562 -1789 563 -1788
rect 576 -1789 577 -1788
rect 625 -1789 626 -1788
rect 751 -1789 752 -1788
rect 779 -1789 780 -1788
rect 793 -1789 794 -1788
rect 877 -1789 878 -1788
rect 968 -1789 969 -1788
rect 971 -1789 972 -1788
rect 2130 -1789 2131 -1788
rect 100 -1791 101 -1790
rect 562 -1791 563 -1790
rect 576 -1791 577 -1790
rect 740 -1791 741 -1790
rect 803 -1791 804 -1790
rect 877 -1791 878 -1790
rect 898 -1791 899 -1790
rect 1279 -1791 1280 -1790
rect 1332 -1791 1333 -1790
rect 1486 -1791 1487 -1790
rect 1570 -1791 1571 -1790
rect 1598 -1791 1599 -1790
rect 1675 -1791 1676 -1790
rect 1927 -1791 1928 -1790
rect 1948 -1791 1949 -1790
rect 1990 -1791 1991 -1790
rect 2060 -1791 2061 -1790
rect 2116 -1791 2117 -1790
rect 128 -1793 129 -1792
rect 527 -1793 528 -1792
rect 625 -1793 626 -1792
rect 646 -1793 647 -1792
rect 674 -1793 675 -1792
rect 709 -1793 710 -1792
rect 719 -1793 720 -1792
rect 1248 -1793 1249 -1792
rect 1346 -1793 1347 -1792
rect 1430 -1793 1431 -1792
rect 1451 -1793 1452 -1792
rect 1570 -1793 1571 -1792
rect 1661 -1793 1662 -1792
rect 1675 -1793 1676 -1792
rect 1717 -1793 1718 -1792
rect 1853 -1793 1854 -1792
rect 1920 -1793 1921 -1792
rect 1948 -1793 1949 -1792
rect 2032 -1793 2033 -1792
rect 2060 -1793 2061 -1792
rect 128 -1795 129 -1794
rect 233 -1795 234 -1794
rect 464 -1795 465 -1794
rect 681 -1795 682 -1794
rect 723 -1795 724 -1794
rect 1101 -1795 1102 -1794
rect 1199 -1795 1200 -1794
rect 1332 -1795 1333 -1794
rect 1346 -1795 1347 -1794
rect 1577 -1795 1578 -1794
rect 1752 -1795 1753 -1794
rect 1794 -1795 1795 -1794
rect 1822 -1795 1823 -1794
rect 1857 -1795 1858 -1794
rect 1892 -1795 1893 -1794
rect 1920 -1795 1921 -1794
rect 2032 -1795 2033 -1794
rect 2441 -1795 2442 -1794
rect 177 -1797 178 -1796
rect 709 -1797 710 -1796
rect 730 -1797 731 -1796
rect 1731 -1797 1732 -1796
rect 1892 -1797 1893 -1796
rect 2095 -1797 2096 -1796
rect 170 -1799 171 -1798
rect 177 -1799 178 -1798
rect 201 -1799 202 -1798
rect 779 -1799 780 -1798
rect 905 -1799 906 -1798
rect 2396 -1799 2397 -1798
rect 156 -1801 157 -1800
rect 170 -1801 171 -1800
rect 215 -1801 216 -1800
rect 1752 -1801 1753 -1800
rect 2011 -1801 2012 -1800
rect 2095 -1801 2096 -1800
rect 233 -1803 234 -1802
rect 485 -1803 486 -1802
rect 499 -1803 500 -1802
rect 569 -1803 570 -1802
rect 604 -1803 605 -1802
rect 723 -1803 724 -1802
rect 933 -1803 934 -1802
rect 2088 -1803 2089 -1802
rect 464 -1805 465 -1804
rect 471 -1805 472 -1804
rect 478 -1805 479 -1804
rect 604 -1805 605 -1804
rect 611 -1805 612 -1804
rect 1451 -1805 1452 -1804
rect 1577 -1805 1578 -1804
rect 1584 -1805 1585 -1804
rect 1962 -1805 1963 -1804
rect 2011 -1805 2012 -1804
rect 72 -1807 73 -1806
rect 471 -1807 472 -1806
rect 499 -1807 500 -1806
rect 555 -1807 556 -1806
rect 936 -1807 937 -1806
rect 996 -1807 997 -1806
rect 1024 -1807 1025 -1806
rect 1199 -1807 1200 -1806
rect 1514 -1807 1515 -1806
rect 1584 -1807 1585 -1806
rect 1710 -1807 1711 -1806
rect 1962 -1807 1963 -1806
rect 72 -1809 73 -1808
rect 401 -1809 402 -1808
rect 506 -1809 507 -1808
rect 814 -1809 815 -1808
rect 940 -1809 941 -1808
rect 2186 -1809 2187 -1808
rect 184 -1811 185 -1810
rect 478 -1811 479 -1810
rect 541 -1811 542 -1810
rect 933 -1811 934 -1810
rect 975 -1811 976 -1810
rect 982 -1811 983 -1810
rect 1024 -1811 1025 -1810
rect 1318 -1811 1319 -1810
rect 1381 -1811 1382 -1810
rect 1514 -1811 1515 -1810
rect 1689 -1811 1690 -1810
rect 1710 -1811 1711 -1810
rect 2186 -1811 2187 -1810
rect 2466 -1811 2467 -1810
rect 401 -1813 402 -1812
rect 583 -1813 584 -1812
rect 814 -1813 815 -1812
rect 842 -1813 843 -1812
rect 975 -1813 976 -1812
rect 1038 -1813 1039 -1812
rect 1136 -1813 1137 -1812
rect 1381 -1813 1382 -1812
rect 1437 -1813 1438 -1812
rect 1689 -1813 1690 -1812
rect 541 -1815 542 -1814
rect 772 -1815 773 -1814
rect 786 -1815 787 -1814
rect 842 -1815 843 -1814
rect 859 -1815 860 -1814
rect 1038 -1815 1039 -1814
rect 1136 -1815 1137 -1814
rect 1178 -1815 1179 -1814
rect 1318 -1815 1319 -1814
rect 1339 -1815 1340 -1814
rect 555 -1817 556 -1816
rect 2427 -1817 2428 -1816
rect 583 -1819 584 -1818
rect 642 -1819 643 -1818
rect 772 -1819 773 -1818
rect 800 -1819 801 -1818
rect 1178 -1819 1179 -1818
rect 1822 -1819 1823 -1818
rect 786 -1821 787 -1820
rect 1087 -1821 1088 -1820
rect 1339 -1821 1340 -1820
rect 2452 -1821 2453 -1820
rect 800 -1823 801 -1822
rect 2067 -1823 2068 -1822
rect 2193 -1823 2194 -1822
rect 2452 -1823 2453 -1822
rect 1087 -1825 1088 -1824
rect 1122 -1825 1123 -1824
rect 2067 -1825 2068 -1824
rect 2256 -1825 2257 -1824
rect 1080 -1827 1081 -1826
rect 1122 -1827 1123 -1826
rect 2144 -1827 2145 -1826
rect 2193 -1827 2194 -1826
rect 2256 -1827 2257 -1826
rect 2431 -1827 2432 -1826
rect 1080 -1829 1081 -1828
rect 1811 -1829 1812 -1828
rect 2109 -1829 2110 -1828
rect 2144 -1829 2145 -1828
rect 2368 -1829 2369 -1828
rect 2431 -1829 2432 -1828
rect 1682 -1831 1683 -1830
rect 2109 -1831 2110 -1830
rect 2277 -1831 2278 -1830
rect 2368 -1831 2369 -1830
rect 1668 -1833 1669 -1832
rect 1682 -1833 1683 -1832
rect 2214 -1833 2215 -1832
rect 2277 -1833 2278 -1832
rect 1654 -1835 1655 -1834
rect 1668 -1835 1669 -1834
rect 1906 -1835 1907 -1834
rect 2214 -1835 2215 -1834
rect 1633 -1837 1634 -1836
rect 1654 -1837 1655 -1836
rect 1864 -1837 1865 -1836
rect 1906 -1837 1907 -1836
rect 1633 -1839 1634 -1838
rect 1766 -1839 1767 -1838
rect 1766 -1841 1767 -1840
rect 1829 -1841 1830 -1840
rect 1780 -1843 1781 -1842
rect 1829 -1843 1830 -1842
rect 1395 -1845 1396 -1844
rect 1780 -1845 1781 -1844
rect 1395 -1847 1396 -1846
rect 1416 -1847 1417 -1846
rect 1416 -1849 1417 -1848
rect 1626 -1849 1627 -1848
rect 30 -1860 31 -1859
rect 611 -1860 612 -1859
rect 618 -1860 619 -1859
rect 1181 -1860 1182 -1859
rect 1206 -1860 1207 -1859
rect 1626 -1860 1627 -1859
rect 1636 -1860 1637 -1859
rect 2368 -1860 2369 -1859
rect 30 -1862 31 -1861
rect 149 -1862 150 -1861
rect 184 -1862 185 -1861
rect 1927 -1862 1928 -1861
rect 2270 -1862 2271 -1861
rect 2469 -1862 2470 -1861
rect 37 -1864 38 -1863
rect 618 -1864 619 -1863
rect 632 -1864 633 -1863
rect 1290 -1864 1291 -1863
rect 1307 -1864 1308 -1863
rect 1647 -1864 1648 -1863
rect 1664 -1864 1665 -1863
rect 2109 -1864 2110 -1863
rect 2319 -1864 2320 -1863
rect 2420 -1864 2421 -1863
rect 37 -1866 38 -1865
rect 191 -1866 192 -1865
rect 194 -1866 195 -1865
rect 614 -1866 615 -1865
rect 635 -1866 636 -1865
rect 1199 -1866 1200 -1865
rect 1206 -1866 1207 -1865
rect 1220 -1866 1221 -1865
rect 1241 -1866 1242 -1865
rect 1244 -1866 1245 -1865
rect 1276 -1866 1277 -1865
rect 1962 -1866 1963 -1865
rect 2109 -1866 2110 -1865
rect 2277 -1866 2278 -1865
rect 2319 -1866 2320 -1865
rect 2417 -1866 2418 -1865
rect 47 -1868 48 -1867
rect 2242 -1868 2243 -1867
rect 2368 -1868 2369 -1867
rect 2410 -1868 2411 -1867
rect 72 -1870 73 -1869
rect 800 -1870 801 -1869
rect 852 -1870 853 -1869
rect 1381 -1870 1382 -1869
rect 1437 -1870 1438 -1869
rect 2221 -1870 2222 -1869
rect 2410 -1870 2411 -1869
rect 2459 -1870 2460 -1869
rect 72 -1872 73 -1871
rect 128 -1872 129 -1871
rect 131 -1872 132 -1871
rect 2270 -1872 2271 -1871
rect 89 -1874 90 -1873
rect 1731 -1874 1732 -1873
rect 1734 -1874 1735 -1873
rect 2452 -1874 2453 -1873
rect 100 -1876 101 -1875
rect 187 -1876 188 -1875
rect 215 -1876 216 -1875
rect 1300 -1876 1301 -1875
rect 1332 -1876 1333 -1875
rect 1335 -1876 1336 -1875
rect 1363 -1876 1364 -1875
rect 1934 -1876 1935 -1875
rect 1962 -1876 1963 -1875
rect 1990 -1876 1991 -1875
rect 2067 -1876 2068 -1875
rect 2277 -1876 2278 -1875
rect 100 -1878 101 -1877
rect 1423 -1878 1424 -1877
rect 1468 -1878 1469 -1877
rect 2207 -1878 2208 -1877
rect 2221 -1878 2222 -1877
rect 2284 -1878 2285 -1877
rect 107 -1880 108 -1879
rect 516 -1880 517 -1879
rect 548 -1880 549 -1879
rect 1440 -1880 1441 -1879
rect 1475 -1880 1476 -1879
rect 2249 -1880 2250 -1879
rect 2256 -1880 2257 -1879
rect 2284 -1880 2285 -1879
rect 107 -1882 108 -1881
rect 135 -1882 136 -1881
rect 142 -1882 143 -1881
rect 1153 -1882 1154 -1881
rect 1164 -1882 1165 -1881
rect 1220 -1882 1221 -1881
rect 1241 -1882 1242 -1881
rect 1325 -1882 1326 -1881
rect 1332 -1882 1333 -1881
rect 1339 -1882 1340 -1881
rect 1353 -1882 1354 -1881
rect 1423 -1882 1424 -1881
rect 1489 -1882 1490 -1881
rect 1577 -1882 1578 -1881
rect 1622 -1882 1623 -1881
rect 1955 -1882 1956 -1881
rect 2067 -1882 2068 -1881
rect 2123 -1882 2124 -1881
rect 2249 -1882 2250 -1881
rect 2291 -1882 2292 -1881
rect 103 -1884 104 -1883
rect 135 -1884 136 -1883
rect 142 -1884 143 -1883
rect 380 -1884 381 -1883
rect 401 -1884 402 -1883
rect 649 -1884 650 -1883
rect 688 -1884 689 -1883
rect 730 -1884 731 -1883
rect 737 -1884 738 -1883
rect 1024 -1884 1025 -1883
rect 1059 -1884 1060 -1883
rect 1069 -1884 1070 -1883
rect 1094 -1884 1095 -1883
rect 1731 -1884 1732 -1883
rect 1773 -1884 1774 -1883
rect 1990 -1884 1991 -1883
rect 2256 -1884 2257 -1883
rect 2305 -1884 2306 -1883
rect 16 -1886 17 -1885
rect 1094 -1886 1095 -1885
rect 1136 -1886 1137 -1885
rect 2088 -1886 2089 -1885
rect 16 -1888 17 -1887
rect 352 -1888 353 -1887
rect 373 -1888 374 -1887
rect 586 -1888 587 -1887
rect 611 -1888 612 -1887
rect 681 -1888 682 -1887
rect 688 -1888 689 -1887
rect 786 -1888 787 -1887
rect 894 -1888 895 -1887
rect 1997 -1888 1998 -1887
rect 124 -1890 125 -1889
rect 1101 -1890 1102 -1889
rect 1129 -1890 1130 -1889
rect 1136 -1890 1137 -1889
rect 1150 -1890 1151 -1889
rect 1199 -1890 1200 -1889
rect 1209 -1890 1210 -1889
rect 2445 -1890 2446 -1889
rect 128 -1892 129 -1891
rect 1073 -1892 1074 -1891
rect 1080 -1892 1081 -1891
rect 1101 -1892 1102 -1891
rect 1129 -1892 1130 -1891
rect 1139 -1892 1140 -1891
rect 1164 -1892 1165 -1891
rect 1458 -1892 1459 -1891
rect 1507 -1892 1508 -1891
rect 2389 -1892 2390 -1891
rect 184 -1894 185 -1893
rect 219 -1894 220 -1893
rect 233 -1894 234 -1893
rect 2123 -1894 2124 -1893
rect 2228 -1894 2229 -1893
rect 2389 -1894 2390 -1893
rect 177 -1896 178 -1895
rect 233 -1896 234 -1895
rect 250 -1896 251 -1895
rect 1430 -1896 1431 -1895
rect 1440 -1896 1441 -1895
rect 2291 -1896 2292 -1895
rect 177 -1898 178 -1897
rect 261 -1898 262 -1897
rect 275 -1898 276 -1897
rect 429 -1898 430 -1897
rect 446 -1898 447 -1897
rect 464 -1898 465 -1897
rect 478 -1898 479 -1897
rect 782 -1898 783 -1897
rect 905 -1898 906 -1897
rect 1612 -1898 1613 -1897
rect 1633 -1898 1634 -1897
rect 1997 -1898 1998 -1897
rect 2032 -1898 2033 -1897
rect 2228 -1898 2229 -1897
rect 205 -1900 206 -1899
rect 380 -1900 381 -1899
rect 401 -1900 402 -1899
rect 632 -1900 633 -1899
rect 646 -1900 647 -1899
rect 1269 -1900 1270 -1899
rect 1290 -1900 1291 -1899
rect 1297 -1900 1298 -1899
rect 1304 -1900 1305 -1899
rect 2207 -1900 2208 -1899
rect 205 -1902 206 -1901
rect 282 -1902 283 -1901
rect 303 -1902 304 -1901
rect 352 -1902 353 -1901
rect 373 -1902 374 -1901
rect 821 -1902 822 -1901
rect 908 -1902 909 -1901
rect 947 -1902 948 -1901
rect 957 -1902 958 -1901
rect 1843 -1902 1844 -1901
rect 1853 -1902 1854 -1901
rect 2424 -1902 2425 -1901
rect 51 -1904 52 -1903
rect 282 -1904 283 -1903
rect 303 -1904 304 -1903
rect 450 -1904 451 -1903
rect 464 -1904 465 -1903
rect 527 -1904 528 -1903
rect 541 -1904 542 -1903
rect 730 -1904 731 -1903
rect 744 -1904 745 -1903
rect 1276 -1904 1277 -1903
rect 1339 -1904 1340 -1903
rect 1367 -1904 1368 -1903
rect 1381 -1904 1382 -1903
rect 1416 -1904 1417 -1903
rect 1430 -1904 1431 -1903
rect 1451 -1904 1452 -1903
rect 1458 -1904 1459 -1903
rect 1472 -1904 1473 -1903
rect 1507 -1904 1508 -1903
rect 1584 -1904 1585 -1903
rect 1605 -1904 1606 -1903
rect 1612 -1904 1613 -1903
rect 1647 -1904 1648 -1903
rect 1850 -1904 1851 -1903
rect 1864 -1904 1865 -1903
rect 2403 -1904 2404 -1903
rect 51 -1906 52 -1905
rect 1605 -1906 1606 -1905
rect 1664 -1906 1665 -1905
rect 2375 -1906 2376 -1905
rect 2403 -1906 2404 -1905
rect 2438 -1906 2439 -1905
rect 219 -1908 220 -1907
rect 1521 -1908 1522 -1907
rect 1577 -1908 1578 -1907
rect 1591 -1908 1592 -1907
rect 1773 -1908 1774 -1907
rect 1822 -1908 1823 -1907
rect 1843 -1908 1844 -1907
rect 2081 -1908 2082 -1907
rect 226 -1910 227 -1909
rect 2375 -1910 2376 -1909
rect 170 -1912 171 -1911
rect 226 -1912 227 -1911
rect 261 -1912 262 -1911
rect 268 -1912 269 -1911
rect 275 -1912 276 -1911
rect 541 -1912 542 -1911
rect 562 -1912 563 -1911
rect 1108 -1912 1109 -1911
rect 1167 -1912 1168 -1911
rect 2305 -1912 2306 -1911
rect 156 -1914 157 -1913
rect 268 -1914 269 -1913
rect 394 -1914 395 -1913
rect 527 -1914 528 -1913
rect 565 -1914 566 -1913
rect 1052 -1914 1053 -1913
rect 1059 -1914 1060 -1913
rect 1346 -1914 1347 -1913
rect 1353 -1914 1354 -1913
rect 1402 -1914 1403 -1913
rect 1416 -1914 1417 -1913
rect 1500 -1914 1501 -1913
rect 1584 -1914 1585 -1913
rect 1619 -1914 1620 -1913
rect 1822 -1914 1823 -1913
rect 1836 -1914 1837 -1913
rect 1850 -1914 1851 -1913
rect 1878 -1914 1879 -1913
rect 1934 -1914 1935 -1913
rect 1969 -1914 1970 -1913
rect 2032 -1914 2033 -1913
rect 2144 -1914 2145 -1913
rect 170 -1916 171 -1915
rect 2158 -1916 2159 -1915
rect 173 -1918 174 -1917
rect 2158 -1918 2159 -1917
rect 229 -1920 230 -1919
rect 1836 -1920 1837 -1919
rect 1864 -1920 1865 -1919
rect 1899 -1920 1900 -1919
rect 1941 -1920 1942 -1919
rect 2144 -1920 2145 -1919
rect 240 -1922 241 -1921
rect 394 -1922 395 -1921
rect 422 -1922 423 -1921
rect 548 -1922 549 -1921
rect 569 -1922 570 -1921
rect 740 -1922 741 -1921
rect 744 -1922 745 -1921
rect 807 -1922 808 -1921
rect 821 -1922 822 -1921
rect 940 -1922 941 -1921
rect 943 -1922 944 -1921
rect 1185 -1922 1186 -1921
rect 1227 -1922 1228 -1921
rect 1269 -1922 1270 -1921
rect 1346 -1922 1347 -1921
rect 1570 -1922 1571 -1921
rect 1591 -1922 1592 -1921
rect 1780 -1922 1781 -1921
rect 1878 -1922 1879 -1921
rect 1913 -1922 1914 -1921
rect 1941 -1922 1942 -1921
rect 1983 -1922 1984 -1921
rect 2081 -1922 2082 -1921
rect 2137 -1922 2138 -1921
rect 2 -1924 3 -1923
rect 240 -1924 241 -1923
rect 422 -1924 423 -1923
rect 544 -1924 545 -1923
rect 646 -1924 647 -1923
rect 863 -1924 864 -1923
rect 919 -1924 920 -1923
rect 947 -1924 948 -1923
rect 957 -1924 958 -1923
rect 2242 -1924 2243 -1923
rect 2 -1926 3 -1925
rect 737 -1926 738 -1925
rect 807 -1926 808 -1925
rect 1010 -1926 1011 -1925
rect 1024 -1926 1025 -1925
rect 1437 -1926 1438 -1925
rect 1444 -1926 1445 -1925
rect 1570 -1926 1571 -1925
rect 1780 -1926 1781 -1925
rect 1829 -1926 1830 -1925
rect 1899 -1926 1900 -1925
rect 2466 -1926 2467 -1925
rect 159 -1928 160 -1927
rect 1010 -1928 1011 -1927
rect 1038 -1928 1039 -1927
rect 1080 -1928 1081 -1927
rect 1178 -1928 1179 -1927
rect 2333 -1928 2334 -1927
rect 9 -1930 10 -1929
rect 159 -1930 160 -1929
rect 429 -1930 430 -1929
rect 499 -1930 500 -1929
rect 506 -1930 507 -1929
rect 740 -1930 741 -1929
rect 863 -1930 864 -1929
rect 975 -1930 976 -1929
rect 978 -1930 979 -1929
rect 1510 -1930 1511 -1929
rect 1913 -1930 1914 -1929
rect 1948 -1930 1949 -1929
rect 1955 -1930 1956 -1929
rect 2011 -1930 2012 -1929
rect 2074 -1930 2075 -1929
rect 2333 -1930 2334 -1929
rect 9 -1932 10 -1931
rect 198 -1932 199 -1931
rect 324 -1932 325 -1931
rect 499 -1932 500 -1931
rect 506 -1932 507 -1931
rect 877 -1932 878 -1931
rect 919 -1932 920 -1931
rect 1122 -1932 1123 -1931
rect 1178 -1932 1179 -1931
rect 1629 -1932 1630 -1931
rect 1696 -1932 1697 -1931
rect 1948 -1932 1949 -1931
rect 1969 -1932 1970 -1931
rect 2004 -1932 2005 -1931
rect 2011 -1932 2012 -1931
rect 2060 -1932 2061 -1931
rect 2074 -1932 2075 -1931
rect 2130 -1932 2131 -1931
rect 2137 -1932 2138 -1931
rect 2193 -1932 2194 -1931
rect 58 -1934 59 -1933
rect 1038 -1934 1039 -1933
rect 1062 -1934 1063 -1933
rect 2298 -1934 2299 -1933
rect 23 -1936 24 -1935
rect 58 -1936 59 -1935
rect 198 -1936 199 -1935
rect 1003 -1936 1004 -1935
rect 1066 -1936 1067 -1935
rect 1619 -1936 1620 -1935
rect 1696 -1936 1697 -1935
rect 1703 -1936 1704 -1935
rect 1983 -1936 1984 -1935
rect 2025 -1936 2026 -1935
rect 2060 -1936 2061 -1935
rect 2116 -1936 2117 -1935
rect 2130 -1936 2131 -1935
rect 2172 -1936 2173 -1935
rect 2298 -1936 2299 -1935
rect 2312 -1936 2313 -1935
rect 23 -1938 24 -1937
rect 114 -1938 115 -1937
rect 324 -1938 325 -1937
rect 1465 -1938 1466 -1937
rect 1472 -1938 1473 -1937
rect 2424 -1938 2425 -1937
rect 114 -1940 115 -1939
rect 758 -1940 759 -1939
rect 828 -1940 829 -1939
rect 877 -1940 878 -1939
rect 926 -1940 927 -1939
rect 1304 -1940 1305 -1939
rect 1367 -1940 1368 -1939
rect 1409 -1940 1410 -1939
rect 1444 -1940 1445 -1939
rect 1479 -1940 1480 -1939
rect 1486 -1940 1487 -1939
rect 1500 -1940 1501 -1939
rect 1703 -1940 1704 -1939
rect 1885 -1940 1886 -1939
rect 1892 -1940 1893 -1939
rect 2116 -1940 2117 -1939
rect 2312 -1940 2313 -1939
rect 2347 -1940 2348 -1939
rect 432 -1942 433 -1941
rect 569 -1942 570 -1941
rect 674 -1942 675 -1941
rect 681 -1942 682 -1941
rect 695 -1942 696 -1941
rect 1003 -1942 1004 -1941
rect 1066 -1942 1067 -1941
rect 1115 -1942 1116 -1941
rect 1185 -1942 1186 -1941
rect 1318 -1942 1319 -1941
rect 1335 -1942 1336 -1941
rect 1409 -1942 1410 -1941
rect 1451 -1942 1452 -1941
rect 1598 -1942 1599 -1941
rect 1724 -1942 1725 -1941
rect 2025 -1942 2026 -1941
rect 2347 -1942 2348 -1941
rect 2382 -1942 2383 -1941
rect 191 -1944 192 -1943
rect 674 -1944 675 -1943
rect 702 -1944 703 -1943
rect 954 -1944 955 -1943
rect 975 -1944 976 -1943
rect 1752 -1944 1753 -1943
rect 1766 -1944 1767 -1943
rect 1885 -1944 1886 -1943
rect 1892 -1944 1893 -1943
rect 2165 -1944 2166 -1943
rect 2179 -1944 2180 -1943
rect 2382 -1944 2383 -1943
rect 450 -1946 451 -1945
rect 590 -1946 591 -1945
rect 660 -1946 661 -1945
rect 695 -1946 696 -1945
rect 702 -1946 703 -1945
rect 996 -1946 997 -1945
rect 1073 -1946 1074 -1945
rect 1867 -1946 1868 -1945
rect 1976 -1946 1977 -1945
rect 2172 -1946 2173 -1945
rect 2179 -1946 2180 -1945
rect 2235 -1946 2236 -1945
rect 121 -1948 122 -1947
rect 660 -1948 661 -1947
rect 709 -1948 710 -1947
rect 940 -1948 941 -1947
rect 982 -1948 983 -1947
rect 996 -1948 997 -1947
rect 1087 -1948 1088 -1947
rect 1115 -1948 1116 -1947
rect 1125 -1948 1126 -1947
rect 1976 -1948 1977 -1947
rect 2004 -1948 2005 -1947
rect 2053 -1948 2054 -1947
rect 86 -1950 87 -1949
rect 982 -1950 983 -1949
rect 1111 -1950 1112 -1949
rect 2193 -1950 2194 -1949
rect 121 -1952 122 -1951
rect 296 -1952 297 -1951
rect 443 -1952 444 -1951
rect 1087 -1952 1088 -1951
rect 1227 -1952 1228 -1951
rect 2235 -1952 2236 -1951
rect 296 -1954 297 -1953
rect 359 -1954 360 -1953
rect 443 -1954 444 -1953
rect 555 -1954 556 -1953
rect 590 -1954 591 -1953
rect 726 -1954 727 -1953
rect 772 -1954 773 -1953
rect 954 -1954 955 -1953
rect 1248 -1954 1249 -1953
rect 1829 -1954 1830 -1953
rect 2053 -1954 2054 -1953
rect 2102 -1954 2103 -1953
rect 289 -1956 290 -1955
rect 555 -1956 556 -1955
rect 653 -1956 654 -1955
rect 709 -1956 710 -1955
rect 723 -1956 724 -1955
rect 758 -1956 759 -1955
rect 772 -1956 773 -1955
rect 922 -1956 923 -1955
rect 926 -1956 927 -1955
rect 1045 -1956 1046 -1955
rect 1213 -1956 1214 -1955
rect 1248 -1956 1249 -1955
rect 1395 -1956 1396 -1955
rect 1402 -1956 1403 -1955
rect 1465 -1956 1466 -1955
rect 1633 -1956 1634 -1955
rect 1654 -1956 1655 -1955
rect 1724 -1956 1725 -1955
rect 1752 -1956 1753 -1955
rect 1759 -1956 1760 -1955
rect 1766 -1956 1767 -1955
rect 1815 -1956 1816 -1955
rect 2102 -1956 2103 -1955
rect 2151 -1956 2152 -1955
rect 289 -1958 290 -1957
rect 849 -1958 850 -1957
rect 933 -1958 934 -1957
rect 1318 -1958 1319 -1957
rect 1360 -1958 1361 -1957
rect 1395 -1958 1396 -1957
rect 1486 -1958 1487 -1957
rect 1927 -1958 1928 -1957
rect 2151 -1958 2152 -1957
rect 2200 -1958 2201 -1957
rect 359 -1960 360 -1959
rect 436 -1960 437 -1959
rect 478 -1960 479 -1959
rect 604 -1960 605 -1959
rect 653 -1960 654 -1959
rect 842 -1960 843 -1959
rect 849 -1960 850 -1959
rect 898 -1960 899 -1959
rect 933 -1960 934 -1959
rect 2473 -1960 2474 -1959
rect 436 -1962 437 -1961
rect 597 -1962 598 -1961
rect 604 -1962 605 -1961
rect 751 -1962 752 -1961
rect 842 -1962 843 -1961
rect 856 -1962 857 -1961
rect 1017 -1962 1018 -1961
rect 1045 -1962 1046 -1961
rect 1213 -1962 1214 -1961
rect 1234 -1962 1235 -1961
rect 1279 -1962 1280 -1961
rect 1815 -1962 1816 -1961
rect 310 -1964 311 -1963
rect 1017 -1964 1018 -1963
rect 1234 -1964 1235 -1963
rect 1311 -1964 1312 -1963
rect 1360 -1964 1361 -1963
rect 2088 -1964 2089 -1963
rect 310 -1966 311 -1965
rect 317 -1966 318 -1965
rect 485 -1966 486 -1965
rect 562 -1966 563 -1965
rect 576 -1966 577 -1965
rect 856 -1966 857 -1965
rect 1297 -1966 1298 -1965
rect 2200 -1966 2201 -1965
rect 212 -1968 213 -1967
rect 317 -1968 318 -1967
rect 485 -1968 486 -1967
rect 492 -1968 493 -1967
rect 513 -1968 514 -1967
rect 803 -1968 804 -1967
rect 1311 -1968 1312 -1967
rect 1661 -1968 1662 -1967
rect 1675 -1968 1676 -1967
rect 1759 -1968 1760 -1967
rect 1801 -1968 1802 -1967
rect 2165 -1968 2166 -1967
rect 149 -1970 150 -1969
rect 212 -1970 213 -1969
rect 247 -1970 248 -1969
rect 492 -1970 493 -1969
rect 534 -1970 535 -1969
rect 597 -1970 598 -1969
rect 625 -1970 626 -1969
rect 898 -1970 899 -1969
rect 1549 -1970 1550 -1969
rect 1598 -1970 1599 -1969
rect 1654 -1970 1655 -1969
rect 1745 -1970 1746 -1969
rect 1801 -1970 1802 -1969
rect 1857 -1970 1858 -1969
rect 86 -1972 87 -1971
rect 247 -1972 248 -1971
rect 387 -1972 388 -1971
rect 513 -1972 514 -1971
rect 576 -1972 577 -1971
rect 793 -1972 794 -1971
rect 1524 -1972 1525 -1971
rect 1745 -1972 1746 -1971
rect 93 -1974 94 -1973
rect 534 -1974 535 -1973
rect 716 -1974 717 -1973
rect 723 -1974 724 -1973
rect 751 -1974 752 -1973
rect 891 -1974 892 -1973
rect 1535 -1974 1536 -1973
rect 1857 -1974 1858 -1973
rect 93 -1976 94 -1975
rect 338 -1976 339 -1975
rect 387 -1976 388 -1975
rect 415 -1976 416 -1975
rect 457 -1976 458 -1975
rect 625 -1976 626 -1975
rect 639 -1976 640 -1975
rect 716 -1976 717 -1975
rect 793 -1976 794 -1975
rect 1108 -1976 1109 -1975
rect 1549 -1976 1550 -1975
rect 2340 -1976 2341 -1975
rect 79 -1978 80 -1977
rect 639 -1978 640 -1977
rect 828 -1978 829 -1977
rect 2340 -1978 2341 -1977
rect 79 -1980 80 -1979
rect 831 -1980 832 -1979
rect 870 -1980 871 -1979
rect 891 -1980 892 -1979
rect 1052 -1980 1053 -1979
rect 1535 -1980 1536 -1979
rect 1661 -1980 1662 -1979
rect 2326 -1980 2327 -1979
rect 254 -1982 255 -1981
rect 457 -1982 458 -1981
rect 870 -1982 871 -1981
rect 912 -1982 913 -1981
rect 1675 -1982 1676 -1981
rect 1682 -1982 1683 -1981
rect 2326 -1982 2327 -1981
rect 2361 -1982 2362 -1981
rect 44 -1984 45 -1983
rect 254 -1984 255 -1983
rect 331 -1984 332 -1983
rect 338 -1984 339 -1983
rect 345 -1984 346 -1983
rect 415 -1984 416 -1983
rect 583 -1984 584 -1983
rect 912 -1984 913 -1983
rect 1682 -1984 1683 -1983
rect 1689 -1984 1690 -1983
rect 2361 -1984 2362 -1983
rect 2396 -1984 2397 -1983
rect 44 -1986 45 -1985
rect 65 -1986 66 -1985
rect 331 -1986 332 -1985
rect 1262 -1986 1263 -1985
rect 1689 -1986 1690 -1985
rect 1710 -1986 1711 -1985
rect 1787 -1986 1788 -1985
rect 2396 -1986 2397 -1985
rect 65 -1988 66 -1987
rect 1374 -1988 1375 -1987
rect 1563 -1988 1564 -1987
rect 1787 -1988 1788 -1987
rect 345 -1990 346 -1989
rect 366 -1990 367 -1989
rect 583 -1990 584 -1989
rect 786 -1990 787 -1989
rect 1255 -1990 1256 -1989
rect 1262 -1990 1263 -1989
rect 1283 -1990 1284 -1989
rect 1563 -1990 1564 -1989
rect 1710 -1990 1711 -1989
rect 1738 -1990 1739 -1989
rect 366 -1992 367 -1991
rect 408 -1992 409 -1991
rect 1171 -1992 1172 -1991
rect 1255 -1992 1256 -1991
rect 1374 -1992 1375 -1991
rect 1388 -1992 1389 -1991
rect 1640 -1992 1641 -1991
rect 1738 -1992 1739 -1991
rect 408 -1994 409 -1993
rect 471 -1994 472 -1993
rect 765 -1994 766 -1993
rect 1171 -1994 1172 -1993
rect 1192 -1994 1193 -1993
rect 1283 -1994 1284 -1993
rect 1388 -1994 1389 -1993
rect 1496 -1994 1497 -1993
rect 1556 -1994 1557 -1993
rect 1640 -1994 1641 -1993
rect 471 -1996 472 -1995
rect 520 -1996 521 -1995
rect 765 -1996 766 -1995
rect 1031 -1996 1032 -1995
rect 1157 -1996 1158 -1995
rect 1192 -1996 1193 -1995
rect 1514 -1996 1515 -1995
rect 1556 -1996 1557 -1995
rect 520 -1998 521 -1997
rect 667 -1998 668 -1997
rect 989 -1998 990 -1997
rect 1031 -1998 1032 -1997
rect 1143 -1998 1144 -1997
rect 1157 -1998 1158 -1997
rect 1514 -1998 1515 -1997
rect 1542 -1998 1543 -1997
rect 635 -2000 636 -1999
rect 667 -2000 668 -1999
rect 779 -2000 780 -1999
rect 1143 -2000 1144 -1999
rect 1493 -2000 1494 -1999
rect 1542 -2000 1543 -1999
rect 968 -2002 969 -2001
rect 989 -2002 990 -2001
rect 1493 -2002 1494 -2001
rect 2214 -2002 2215 -2001
rect 884 -2004 885 -2003
rect 968 -2004 969 -2003
rect 2214 -2004 2215 -2003
rect 2263 -2004 2264 -2003
rect 884 -2006 885 -2005
rect 1668 -2006 1669 -2005
rect 2039 -2006 2040 -2005
rect 2263 -2006 2264 -2005
rect 1668 -2008 1669 -2007
rect 1794 -2008 1795 -2007
rect 2039 -2008 2040 -2007
rect 2095 -2008 2096 -2007
rect 1794 -2010 1795 -2009
rect 2018 -2010 2019 -2009
rect 2095 -2010 2096 -2009
rect 2354 -2010 2355 -2009
rect 1808 -2012 1809 -2011
rect 2018 -2012 2019 -2011
rect 2354 -2012 2355 -2011
rect 2431 -2012 2432 -2011
rect 1808 -2014 1809 -2013
rect 1871 -2014 1872 -2013
rect 1871 -2016 1872 -2015
rect 1906 -2016 1907 -2015
rect 1906 -2018 1907 -2017
rect 1920 -2018 1921 -2017
rect 1920 -2020 1921 -2019
rect 2046 -2020 2047 -2019
rect 1717 -2022 1718 -2021
rect 2046 -2022 2047 -2021
rect 779 -2024 780 -2023
rect 1717 -2024 1718 -2023
rect 9 -2035 10 -2034
rect 761 -2035 762 -2034
rect 800 -2035 801 -2034
rect 849 -2035 850 -2034
rect 898 -2035 899 -2034
rect 1108 -2035 1109 -2034
rect 1111 -2035 1112 -2034
rect 1206 -2035 1207 -2034
rect 1230 -2035 1231 -2034
rect 1300 -2035 1301 -2034
rect 1335 -2035 1336 -2034
rect 1976 -2035 1977 -2034
rect 2403 -2035 2404 -2034
rect 2417 -2035 2418 -2034
rect 9 -2037 10 -2036
rect 44 -2037 45 -2036
rect 51 -2037 52 -2036
rect 65 -2037 66 -2036
rect 86 -2037 87 -2036
rect 135 -2037 136 -2036
rect 138 -2037 139 -2036
rect 1017 -2037 1018 -2036
rect 1024 -2037 1025 -2036
rect 1108 -2037 1109 -2036
rect 1122 -2037 1123 -2036
rect 1423 -2037 1424 -2036
rect 1437 -2037 1438 -2036
rect 2424 -2037 2425 -2036
rect 37 -2039 38 -2038
rect 831 -2039 832 -2038
rect 898 -2039 899 -2038
rect 1304 -2039 1305 -2038
rect 1360 -2039 1361 -2038
rect 1640 -2039 1641 -2038
rect 1713 -2039 1714 -2038
rect 1969 -2039 1970 -2038
rect 37 -2041 38 -2040
rect 240 -2041 241 -2040
rect 296 -2041 297 -2040
rect 1062 -2041 1063 -2040
rect 1073 -2041 1074 -2040
rect 1206 -2041 1207 -2040
rect 1297 -2041 1298 -2040
rect 1857 -2041 1858 -2040
rect 1934 -2041 1935 -2040
rect 2403 -2041 2404 -2040
rect 30 -2043 31 -2042
rect 240 -2043 241 -2042
rect 296 -2043 297 -2042
rect 471 -2043 472 -2042
rect 492 -2043 493 -2042
rect 1017 -2043 1018 -2042
rect 1024 -2043 1025 -2042
rect 1430 -2043 1431 -2042
rect 1437 -2043 1438 -2042
rect 1444 -2043 1445 -2042
rect 1472 -2043 1473 -2042
rect 1878 -2043 1879 -2042
rect 1969 -2043 1970 -2042
rect 2375 -2043 2376 -2042
rect 16 -2045 17 -2044
rect 471 -2045 472 -2044
rect 499 -2045 500 -2044
rect 541 -2045 542 -2044
rect 569 -2045 570 -2044
rect 1122 -2045 1123 -2044
rect 1150 -2045 1151 -2044
rect 2291 -2045 2292 -2044
rect 2340 -2045 2341 -2044
rect 2375 -2045 2376 -2044
rect 16 -2047 17 -2046
rect 807 -2047 808 -2046
rect 828 -2047 829 -2046
rect 1409 -2047 1410 -2046
rect 1430 -2047 1431 -2046
rect 1983 -2047 1984 -2046
rect 2249 -2047 2250 -2046
rect 2291 -2047 2292 -2046
rect 2298 -2047 2299 -2046
rect 2340 -2047 2341 -2046
rect 30 -2049 31 -2048
rect 72 -2049 73 -2048
rect 89 -2049 90 -2048
rect 884 -2049 885 -2048
rect 919 -2049 920 -2048
rect 926 -2049 927 -2048
rect 954 -2049 955 -2048
rect 2354 -2049 2355 -2048
rect 44 -2051 45 -2050
rect 695 -2051 696 -2050
rect 751 -2051 752 -2050
rect 849 -2051 850 -2050
rect 922 -2051 923 -2050
rect 1031 -2051 1032 -2050
rect 1153 -2051 1154 -2050
rect 1395 -2051 1396 -2050
rect 1402 -2051 1403 -2050
rect 1423 -2051 1424 -2050
rect 1440 -2051 1441 -2050
rect 2116 -2051 2117 -2050
rect 2214 -2051 2215 -2050
rect 2249 -2051 2250 -2050
rect 2 -2053 3 -2052
rect 1153 -2053 1154 -2052
rect 1171 -2053 1172 -2052
rect 1342 -2053 1343 -2052
rect 1363 -2053 1364 -2052
rect 2228 -2053 2229 -2052
rect 51 -2055 52 -2054
rect 1696 -2055 1697 -2054
rect 1766 -2055 1767 -2054
rect 2424 -2055 2425 -2054
rect 58 -2057 59 -2056
rect 1360 -2057 1361 -2056
rect 1384 -2057 1385 -2056
rect 1598 -2057 1599 -2056
rect 1605 -2057 1606 -2056
rect 1696 -2057 1697 -2056
rect 1808 -2057 1809 -2056
rect 1878 -2057 1879 -2056
rect 2095 -2057 2096 -2056
rect 2354 -2057 2355 -2056
rect 58 -2059 59 -2058
rect 96 -2059 97 -2058
rect 100 -2059 101 -2058
rect 107 -2059 108 -2058
rect 156 -2059 157 -2058
rect 2305 -2059 2306 -2058
rect 65 -2061 66 -2060
rect 702 -2061 703 -2060
rect 758 -2061 759 -2060
rect 803 -2061 804 -2060
rect 807 -2061 808 -2060
rect 1318 -2061 1319 -2060
rect 1402 -2061 1403 -2060
rect 2025 -2061 2026 -2060
rect 2095 -2061 2096 -2060
rect 2186 -2061 2187 -2060
rect 2228 -2061 2229 -2060
rect 2284 -2061 2285 -2060
rect 2305 -2061 2306 -2060
rect 2312 -2061 2313 -2060
rect 72 -2063 73 -2062
rect 961 -2063 962 -2062
rect 1031 -2063 1032 -2062
rect 1129 -2063 1130 -2062
rect 1178 -2063 1179 -2062
rect 1640 -2063 1641 -2062
rect 1654 -2063 1655 -2062
rect 1808 -2063 1809 -2062
rect 1815 -2063 1816 -2062
rect 1976 -2063 1977 -2062
rect 2046 -2063 2047 -2062
rect 2312 -2063 2313 -2062
rect 100 -2065 101 -2064
rect 1405 -2065 1406 -2064
rect 1409 -2065 1410 -2064
rect 1885 -2065 1886 -2064
rect 1920 -2065 1921 -2064
rect 2046 -2065 2047 -2064
rect 2116 -2065 2117 -2064
rect 2130 -2065 2131 -2064
rect 2172 -2065 2173 -2064
rect 2214 -2065 2215 -2064
rect 2256 -2065 2257 -2064
rect 2284 -2065 2285 -2064
rect 107 -2067 108 -2066
rect 1167 -2067 1168 -2066
rect 1178 -2067 1179 -2066
rect 1192 -2067 1193 -2066
rect 1220 -2067 1221 -2066
rect 1318 -2067 1319 -2066
rect 1486 -2067 1487 -2066
rect 1990 -2067 1991 -2066
rect 2074 -2067 2075 -2066
rect 2130 -2067 2131 -2066
rect 2137 -2067 2138 -2066
rect 2172 -2067 2173 -2066
rect 2186 -2067 2187 -2066
rect 2347 -2067 2348 -2066
rect 156 -2069 157 -2068
rect 457 -2069 458 -2068
rect 516 -2069 517 -2068
rect 1003 -2069 1004 -2068
rect 1038 -2069 1039 -2068
rect 1129 -2069 1130 -2068
rect 1192 -2069 1193 -2068
rect 1290 -2069 1291 -2068
rect 1297 -2069 1298 -2068
rect 1307 -2069 1308 -2068
rect 1486 -2069 1487 -2068
rect 1724 -2069 1725 -2068
rect 1745 -2069 1746 -2068
rect 1815 -2069 1816 -2068
rect 1871 -2069 1872 -2068
rect 1920 -2069 1921 -2068
rect 1948 -2069 1949 -2068
rect 1990 -2069 1991 -2068
rect 2018 -2069 2019 -2068
rect 2074 -2069 2075 -2068
rect 2081 -2069 2082 -2068
rect 2137 -2069 2138 -2068
rect 2207 -2069 2208 -2068
rect 2256 -2069 2257 -2068
rect 2333 -2069 2334 -2068
rect 2347 -2069 2348 -2068
rect 159 -2071 160 -2070
rect 905 -2071 906 -2070
rect 1003 -2071 1004 -2070
rect 1255 -2071 1256 -2070
rect 1269 -2071 1270 -2070
rect 1983 -2071 1984 -2070
rect 173 -2073 174 -2072
rect 1241 -2073 1242 -2072
rect 1276 -2073 1277 -2072
rect 1395 -2073 1396 -2072
rect 1489 -2073 1490 -2072
rect 2298 -2073 2299 -2072
rect 191 -2075 192 -2074
rect 506 -2075 507 -2074
rect 569 -2075 570 -2074
rect 978 -2075 979 -2074
rect 1038 -2075 1039 -2074
rect 1066 -2075 1067 -2074
rect 1080 -2075 1081 -2074
rect 1171 -2075 1172 -2074
rect 1234 -2075 1235 -2074
rect 1444 -2075 1445 -2074
rect 1521 -2075 1522 -2074
rect 1759 -2075 1760 -2074
rect 1843 -2075 1844 -2074
rect 2081 -2075 2082 -2074
rect 191 -2077 192 -2076
rect 586 -2077 587 -2076
rect 590 -2077 591 -2076
rect 656 -2077 657 -2076
rect 670 -2077 671 -2076
rect 744 -2077 745 -2076
rect 758 -2077 759 -2076
rect 884 -2077 885 -2076
rect 891 -2077 892 -2076
rect 905 -2077 906 -2076
rect 978 -2077 979 -2076
rect 1822 -2077 1823 -2076
rect 1871 -2077 1872 -2076
rect 1941 -2077 1942 -2076
rect 1955 -2077 1956 -2076
rect 2018 -2077 2019 -2076
rect 170 -2079 171 -2078
rect 590 -2079 591 -2078
rect 604 -2079 605 -2078
rect 779 -2079 780 -2078
rect 786 -2079 787 -2078
rect 800 -2079 801 -2078
rect 828 -2079 829 -2078
rect 968 -2079 969 -2078
rect 989 -2079 990 -2078
rect 1234 -2079 1235 -2078
rect 1283 -2079 1284 -2078
rect 1290 -2079 1291 -2078
rect 1304 -2079 1305 -2078
rect 1416 -2079 1417 -2078
rect 1521 -2079 1522 -2078
rect 1612 -2079 1613 -2078
rect 1622 -2079 1623 -2078
rect 2032 -2079 2033 -2078
rect 170 -2081 171 -2080
rect 730 -2081 731 -2080
rect 740 -2081 741 -2080
rect 2025 -2081 2026 -2080
rect 194 -2083 195 -2082
rect 1724 -2083 1725 -2082
rect 1752 -2083 1753 -2082
rect 1822 -2083 1823 -2082
rect 1899 -2083 1900 -2082
rect 1941 -2083 1942 -2082
rect 1955 -2083 1956 -2082
rect 2389 -2083 2390 -2082
rect 212 -2085 213 -2084
rect 317 -2085 318 -2084
rect 331 -2085 332 -2084
rect 961 -2085 962 -2084
rect 1059 -2085 1060 -2084
rect 2333 -2085 2334 -2084
rect 2361 -2085 2362 -2084
rect 2389 -2085 2390 -2084
rect 93 -2087 94 -2086
rect 331 -2087 332 -2086
rect 338 -2087 339 -2086
rect 457 -2087 458 -2086
rect 464 -2087 465 -2086
rect 604 -2087 605 -2086
rect 618 -2087 619 -2086
rect 751 -2087 752 -2086
rect 793 -2087 794 -2086
rect 926 -2087 927 -2086
rect 940 -2087 941 -2086
rect 989 -2087 990 -2086
rect 1066 -2087 1067 -2086
rect 1664 -2087 1665 -2086
rect 1689 -2087 1690 -2086
rect 1766 -2087 1767 -2086
rect 1773 -2087 1774 -2086
rect 1843 -2087 1844 -2086
rect 1850 -2087 1851 -2086
rect 1899 -2087 1900 -2086
rect 1906 -2087 1907 -2086
rect 1948 -2087 1949 -2086
rect 2326 -2087 2327 -2086
rect 2361 -2087 2362 -2086
rect 93 -2089 94 -2088
rect 1465 -2089 1466 -2088
rect 1479 -2089 1480 -2088
rect 1752 -2089 1753 -2088
rect 1780 -2089 1781 -2088
rect 1850 -2089 1851 -2088
rect 2004 -2089 2005 -2088
rect 2326 -2089 2327 -2088
rect 103 -2091 104 -2090
rect 1773 -2091 1774 -2090
rect 1780 -2091 1781 -2090
rect 1913 -2091 1914 -2090
rect 114 -2093 115 -2092
rect 793 -2093 794 -2092
rect 835 -2093 836 -2092
rect 919 -2093 920 -2092
rect 940 -2093 941 -2092
rect 982 -2093 983 -2092
rect 1080 -2093 1081 -2092
rect 1094 -2093 1095 -2092
rect 1143 -2093 1144 -2092
rect 1241 -2093 1242 -2092
rect 1311 -2093 1312 -2092
rect 1416 -2093 1417 -2092
rect 1451 -2093 1452 -2092
rect 1689 -2093 1690 -2092
rect 1703 -2093 1704 -2092
rect 1906 -2093 1907 -2092
rect 114 -2095 115 -2094
rect 352 -2095 353 -2094
rect 366 -2095 367 -2094
rect 464 -2095 465 -2094
rect 562 -2095 563 -2094
rect 618 -2095 619 -2094
rect 653 -2095 654 -2094
rect 954 -2095 955 -2094
rect 1094 -2095 1095 -2094
rect 1101 -2095 1102 -2094
rect 1136 -2095 1137 -2094
rect 1311 -2095 1312 -2094
rect 1332 -2095 1333 -2094
rect 1465 -2095 1466 -2094
rect 1500 -2095 1501 -2094
rect 1612 -2095 1613 -2094
rect 1626 -2095 1627 -2094
rect 1745 -2095 1746 -2094
rect 1794 -2095 1795 -2094
rect 2032 -2095 2033 -2094
rect 205 -2097 206 -2096
rect 352 -2097 353 -2096
rect 404 -2097 405 -2096
rect 968 -2097 969 -2096
rect 1010 -2097 1011 -2096
rect 1101 -2097 1102 -2096
rect 1136 -2097 1137 -2096
rect 1213 -2097 1214 -2096
rect 1325 -2097 1326 -2096
rect 1500 -2097 1501 -2096
rect 1528 -2097 1529 -2096
rect 1654 -2097 1655 -2096
rect 1703 -2097 1704 -2096
rect 1864 -2097 1865 -2096
rect 177 -2099 178 -2098
rect 205 -2099 206 -2098
rect 215 -2099 216 -2098
rect 1731 -2099 1732 -2098
rect 1801 -2099 1802 -2098
rect 1864 -2099 1865 -2098
rect 163 -2101 164 -2100
rect 177 -2101 178 -2100
rect 219 -2101 220 -2100
rect 1059 -2101 1060 -2100
rect 1143 -2101 1144 -2100
rect 1223 -2101 1224 -2100
rect 1262 -2101 1263 -2100
rect 1325 -2101 1326 -2100
rect 1332 -2101 1333 -2100
rect 2270 -2101 2271 -2100
rect 124 -2103 125 -2102
rect 163 -2103 164 -2102
rect 219 -2103 220 -2102
rect 1650 -2103 1651 -2102
rect 2221 -2103 2222 -2102
rect 2270 -2103 2271 -2102
rect 236 -2105 237 -2104
rect 681 -2105 682 -2104
rect 688 -2105 689 -2104
rect 1276 -2105 1277 -2104
rect 1353 -2105 1354 -2104
rect 1528 -2105 1529 -2104
rect 1535 -2105 1536 -2104
rect 1962 -2105 1963 -2104
rect 2179 -2105 2180 -2104
rect 2221 -2105 2222 -2104
rect 247 -2107 248 -2106
rect 1759 -2107 1760 -2106
rect 1927 -2107 1928 -2106
rect 1962 -2107 1963 -2106
rect 2165 -2107 2166 -2106
rect 2179 -2107 2180 -2106
rect 247 -2109 248 -2108
rect 289 -2109 290 -2108
rect 303 -2109 304 -2108
rect 506 -2109 507 -2108
rect 583 -2109 584 -2108
rect 611 -2109 612 -2108
rect 625 -2109 626 -2108
rect 681 -2109 682 -2108
rect 695 -2109 696 -2108
rect 957 -2109 958 -2108
rect 1010 -2109 1011 -2108
rect 1045 -2109 1046 -2108
rect 1164 -2109 1165 -2108
rect 2004 -2109 2005 -2108
rect 2123 -2109 2124 -2108
rect 2165 -2109 2166 -2108
rect 261 -2111 262 -2110
rect 317 -2111 318 -2110
rect 338 -2111 339 -2110
rect 1552 -2111 1553 -2110
rect 1563 -2111 1564 -2110
rect 1934 -2111 1935 -2110
rect 2067 -2111 2068 -2110
rect 2123 -2111 2124 -2110
rect 142 -2113 143 -2112
rect 261 -2113 262 -2112
rect 275 -2113 276 -2112
rect 688 -2113 689 -2112
rect 702 -2113 703 -2112
rect 1258 -2113 1259 -2112
rect 1262 -2113 1263 -2112
rect 1475 -2113 1476 -2112
rect 1538 -2113 1539 -2112
rect 1927 -2113 1928 -2112
rect 2011 -2113 2012 -2112
rect 2067 -2113 2068 -2112
rect 142 -2115 143 -2114
rect 1580 -2115 1581 -2114
rect 1584 -2115 1585 -2114
rect 1794 -2115 1795 -2114
rect 275 -2117 276 -2116
rect 548 -2117 549 -2116
rect 597 -2117 598 -2116
rect 611 -2117 612 -2116
rect 625 -2117 626 -2116
rect 856 -2117 857 -2116
rect 863 -2117 864 -2116
rect 1269 -2117 1270 -2116
rect 1367 -2117 1368 -2116
rect 1535 -2117 1536 -2116
rect 1542 -2117 1543 -2116
rect 1913 -2117 1914 -2116
rect 289 -2119 290 -2118
rect 387 -2119 388 -2118
rect 422 -2119 423 -2118
rect 1073 -2119 1074 -2118
rect 1164 -2119 1165 -2118
rect 1199 -2119 1200 -2118
rect 1213 -2119 1214 -2118
rect 1493 -2119 1494 -2118
rect 1549 -2119 1550 -2118
rect 2109 -2119 2110 -2118
rect 226 -2121 227 -2120
rect 387 -2121 388 -2120
rect 436 -2121 437 -2120
rect 597 -2121 598 -2120
rect 653 -2121 654 -2120
rect 2207 -2121 2208 -2120
rect 226 -2123 227 -2122
rect 646 -2123 647 -2122
rect 660 -2123 661 -2122
rect 1626 -2123 1627 -2122
rect 1636 -2123 1637 -2122
rect 2011 -2123 2012 -2122
rect 2060 -2123 2061 -2122
rect 2109 -2123 2110 -2122
rect 233 -2125 234 -2124
rect 422 -2125 423 -2124
rect 443 -2125 444 -2124
rect 646 -2125 647 -2124
rect 660 -2125 661 -2124
rect 975 -2125 976 -2124
rect 1188 -2125 1189 -2124
rect 1283 -2125 1284 -2124
rect 1339 -2125 1340 -2124
rect 1493 -2125 1494 -2124
rect 1549 -2125 1550 -2124
rect 1633 -2125 1634 -2124
rect 2060 -2125 2061 -2124
rect 2263 -2125 2264 -2124
rect 303 -2127 304 -2126
rect 555 -2127 556 -2126
rect 576 -2127 577 -2126
rect 863 -2127 864 -2126
rect 891 -2127 892 -2126
rect 1619 -2127 1620 -2126
rect 1633 -2127 1634 -2126
rect 1710 -2127 1711 -2126
rect 2235 -2127 2236 -2126
rect 2263 -2127 2264 -2126
rect 23 -2129 24 -2128
rect 1619 -2129 1620 -2128
rect 2193 -2129 2194 -2128
rect 2235 -2129 2236 -2128
rect 23 -2131 24 -2130
rect 131 -2131 132 -2130
rect 345 -2131 346 -2130
rect 366 -2131 367 -2130
rect 373 -2131 374 -2130
rect 548 -2131 549 -2130
rect 555 -2131 556 -2130
rect 870 -2131 871 -2130
rect 933 -2131 934 -2130
rect 1045 -2131 1046 -2130
rect 1188 -2131 1189 -2130
rect 1997 -2131 1998 -2130
rect 2151 -2131 2152 -2130
rect 2193 -2131 2194 -2130
rect 131 -2133 132 -2132
rect 212 -2133 213 -2132
rect 345 -2133 346 -2132
rect 401 -2133 402 -2132
rect 443 -2133 444 -2132
rect 996 -2133 997 -2132
rect 1199 -2133 1200 -2132
rect 2319 -2133 2320 -2132
rect 149 -2135 150 -2134
rect 870 -2135 871 -2134
rect 947 -2135 948 -2134
rect 982 -2135 983 -2134
rect 1248 -2135 1249 -2134
rect 1353 -2135 1354 -2134
rect 1381 -2135 1382 -2134
rect 1542 -2135 1543 -2134
rect 1563 -2135 1564 -2134
rect 1787 -2135 1788 -2134
rect 2151 -2135 2152 -2134
rect 2382 -2135 2383 -2134
rect 54 -2137 55 -2136
rect 149 -2137 150 -2136
rect 373 -2137 374 -2136
rect 1202 -2137 1203 -2136
rect 1381 -2137 1382 -2136
rect 1997 -2137 1998 -2136
rect 2144 -2137 2145 -2136
rect 2382 -2137 2383 -2136
rect 394 -2139 395 -2138
rect 436 -2139 437 -2138
rect 450 -2139 451 -2138
rect 632 -2139 633 -2138
rect 639 -2139 640 -2138
rect 996 -2139 997 -2138
rect 1157 -2139 1158 -2138
rect 1248 -2139 1249 -2138
rect 1570 -2139 1571 -2138
rect 1801 -2139 1802 -2138
rect 2088 -2139 2089 -2138
rect 2144 -2139 2145 -2138
rect 79 -2141 80 -2140
rect 394 -2141 395 -2140
rect 401 -2141 402 -2140
rect 408 -2141 409 -2140
rect 492 -2141 493 -2140
rect 562 -2141 563 -2140
rect 632 -2141 633 -2140
rect 1055 -2141 1056 -2140
rect 1125 -2141 1126 -2140
rect 1157 -2141 1158 -2140
rect 1458 -2141 1459 -2140
rect 1570 -2141 1571 -2140
rect 1577 -2141 1578 -2140
rect 1885 -2141 1886 -2140
rect 2039 -2141 2040 -2140
rect 2088 -2141 2089 -2140
rect 79 -2143 80 -2142
rect 534 -2143 535 -2142
rect 674 -2143 675 -2142
rect 856 -2143 857 -2142
rect 1052 -2143 1053 -2142
rect 1458 -2143 1459 -2142
rect 1584 -2143 1585 -2142
rect 1591 -2143 1592 -2142
rect 1598 -2143 1599 -2142
rect 1682 -2143 1683 -2142
rect 1787 -2143 1788 -2142
rect 2396 -2143 2397 -2142
rect 121 -2145 122 -2144
rect 450 -2145 451 -2144
rect 527 -2145 528 -2144
rect 576 -2145 577 -2144
rect 709 -2145 710 -2144
rect 779 -2145 780 -2144
rect 821 -2145 822 -2144
rect 1451 -2145 1452 -2144
rect 1556 -2145 1557 -2144
rect 1591 -2145 1592 -2144
rect 1605 -2145 1606 -2144
rect 1675 -2145 1676 -2144
rect 1682 -2145 1683 -2144
rect 1829 -2145 1830 -2144
rect 2396 -2145 2397 -2144
rect 2410 -2145 2411 -2144
rect 135 -2147 136 -2146
rect 527 -2147 528 -2146
rect 534 -2147 535 -2146
rect 1339 -2147 1340 -2146
rect 1507 -2147 1508 -2146
rect 1675 -2147 1676 -2146
rect 2102 -2147 2103 -2146
rect 2410 -2147 2411 -2146
rect 254 -2149 255 -2148
rect 674 -2149 675 -2148
rect 716 -2149 717 -2148
rect 786 -2149 787 -2148
rect 842 -2149 843 -2148
rect 947 -2149 948 -2148
rect 1052 -2149 1053 -2148
rect 1738 -2149 1739 -2148
rect 2053 -2149 2054 -2148
rect 2102 -2149 2103 -2148
rect 257 -2151 258 -2150
rect 821 -2151 822 -2150
rect 1185 -2151 1186 -2150
rect 2039 -2151 2040 -2150
rect 268 -2153 269 -2152
rect 639 -2153 640 -2152
rect 723 -2153 724 -2152
rect 835 -2153 836 -2152
rect 1185 -2153 1186 -2152
rect 2242 -2153 2243 -2152
rect 268 -2155 269 -2154
rect 1367 -2155 1368 -2154
rect 1374 -2155 1375 -2154
rect 1507 -2155 1508 -2154
rect 1556 -2155 1557 -2154
rect 1717 -2155 1718 -2154
rect 2200 -2155 2201 -2154
rect 2242 -2155 2243 -2154
rect 408 -2157 409 -2156
rect 415 -2157 416 -2156
rect 478 -2157 479 -2156
rect 709 -2157 710 -2156
rect 730 -2157 731 -2156
rect 877 -2157 878 -2156
rect 1230 -2157 1231 -2156
rect 1738 -2157 1739 -2156
rect 2158 -2157 2159 -2156
rect 2200 -2157 2201 -2156
rect 233 -2159 234 -2158
rect 478 -2159 479 -2158
rect 513 -2159 514 -2158
rect 723 -2159 724 -2158
rect 747 -2159 748 -2158
rect 933 -2159 934 -2158
rect 1255 -2159 1256 -2158
rect 1374 -2159 1375 -2158
rect 1647 -2159 1648 -2158
rect 2053 -2159 2054 -2158
rect 282 -2161 283 -2160
rect 513 -2161 514 -2160
rect 520 -2161 521 -2160
rect 716 -2161 717 -2160
rect 765 -2161 766 -2160
rect 1479 -2161 1480 -2160
rect 1647 -2161 1648 -2160
rect 2277 -2161 2278 -2160
rect 282 -2163 283 -2162
rect 324 -2163 325 -2162
rect 359 -2163 360 -2162
rect 520 -2163 521 -2162
rect 765 -2163 766 -2162
rect 772 -2163 773 -2162
rect 814 -2163 815 -2162
rect 842 -2163 843 -2162
rect 877 -2163 878 -2162
rect 1661 -2163 1662 -2162
rect 1668 -2163 1669 -2162
rect 1829 -2163 1830 -2162
rect 1892 -2163 1893 -2162
rect 2158 -2163 2159 -2162
rect 324 -2165 325 -2164
rect 429 -2165 430 -2164
rect 667 -2165 668 -2164
rect 814 -2165 815 -2164
rect 1346 -2165 1347 -2164
rect 1668 -2165 1669 -2164
rect 1717 -2165 1718 -2164
rect 1857 -2165 1858 -2164
rect 359 -2167 360 -2166
rect 485 -2167 486 -2166
rect 499 -2167 500 -2166
rect 667 -2167 668 -2166
rect 772 -2167 773 -2166
rect 912 -2167 913 -2166
rect 1346 -2167 1347 -2166
rect 1388 -2167 1389 -2166
rect 1496 -2167 1497 -2166
rect 2277 -2167 2278 -2166
rect 198 -2169 199 -2168
rect 485 -2169 486 -2168
rect 737 -2169 738 -2168
rect 1388 -2169 1389 -2168
rect 1514 -2169 1515 -2168
rect 1661 -2169 1662 -2168
rect 1836 -2169 1837 -2168
rect 1892 -2169 1893 -2168
rect 184 -2171 185 -2170
rect 198 -2171 199 -2170
rect 380 -2171 381 -2170
rect 415 -2171 416 -2170
rect 429 -2171 430 -2170
rect 744 -2171 745 -2170
rect 912 -2171 913 -2170
rect 1577 -2171 1578 -2170
rect 1836 -2171 1837 -2170
rect 2319 -2171 2320 -2170
rect 121 -2173 122 -2172
rect 380 -2173 381 -2172
rect 737 -2173 738 -2172
rect 1489 -2173 1490 -2172
rect 184 -2175 185 -2174
rect 243 -2175 244 -2174
rect 1220 -2175 1221 -2174
rect 1514 -2175 1515 -2174
rect 2 -2186 3 -2185
rect 674 -2186 675 -2185
rect 744 -2186 745 -2185
rect 1234 -2186 1235 -2185
rect 1258 -2186 1259 -2185
rect 2312 -2186 2313 -2185
rect 2343 -2186 2344 -2185
rect 2396 -2186 2397 -2185
rect 9 -2188 10 -2187
rect 51 -2188 52 -2187
rect 54 -2188 55 -2187
rect 1388 -2188 1389 -2187
rect 1398 -2188 1399 -2187
rect 1885 -2188 1886 -2187
rect 1937 -2188 1938 -2187
rect 2298 -2188 2299 -2187
rect 37 -2190 38 -2189
rect 996 -2190 997 -2189
rect 1038 -2190 1039 -2189
rect 1223 -2190 1224 -2189
rect 1227 -2190 1228 -2189
rect 2305 -2190 2306 -2189
rect 51 -2192 52 -2191
rect 1031 -2192 1032 -2191
rect 1080 -2192 1081 -2191
rect 1150 -2192 1151 -2191
rect 1157 -2192 1158 -2191
rect 1388 -2192 1389 -2191
rect 1405 -2192 1406 -2191
rect 1437 -2192 1438 -2191
rect 1489 -2192 1490 -2191
rect 2403 -2192 2404 -2191
rect 65 -2194 66 -2193
rect 1041 -2194 1042 -2193
rect 1080 -2194 1081 -2193
rect 1101 -2194 1102 -2193
rect 1115 -2194 1116 -2193
rect 1139 -2194 1140 -2193
rect 1143 -2194 1144 -2193
rect 1234 -2194 1235 -2193
rect 1293 -2194 1294 -2193
rect 1983 -2194 1984 -2193
rect 2151 -2194 2152 -2193
rect 2305 -2194 2306 -2193
rect 65 -2196 66 -2195
rect 1276 -2196 1277 -2195
rect 1304 -2196 1305 -2195
rect 1927 -2196 1928 -2195
rect 1969 -2196 1970 -2195
rect 2298 -2196 2299 -2195
rect 93 -2198 94 -2197
rect 1479 -2198 1480 -2197
rect 1496 -2198 1497 -2197
rect 1752 -2198 1753 -2197
rect 1780 -2198 1781 -2197
rect 1783 -2198 1784 -2197
rect 1836 -2198 1837 -2197
rect 1871 -2198 1872 -2197
rect 1885 -2198 1886 -2197
rect 1962 -2198 1963 -2197
rect 1969 -2198 1970 -2197
rect 2032 -2198 2033 -2197
rect 2151 -2198 2152 -2197
rect 2270 -2198 2271 -2197
rect 93 -2200 94 -2199
rect 1360 -2200 1361 -2199
rect 1367 -2200 1368 -2199
rect 2172 -2200 2173 -2199
rect 2228 -2200 2229 -2199
rect 2336 -2200 2337 -2199
rect 96 -2202 97 -2201
rect 926 -2202 927 -2201
rect 936 -2202 937 -2201
rect 1010 -2202 1011 -2201
rect 1031 -2202 1032 -2201
rect 1045 -2202 1046 -2201
rect 1094 -2202 1095 -2201
rect 1157 -2202 1158 -2201
rect 1192 -2202 1193 -2201
rect 1255 -2202 1256 -2201
rect 1304 -2202 1305 -2201
rect 1416 -2202 1417 -2201
rect 1437 -2202 1438 -2201
rect 1514 -2202 1515 -2201
rect 1521 -2202 1522 -2201
rect 1752 -2202 1753 -2201
rect 1780 -2202 1781 -2201
rect 1843 -2202 1844 -2201
rect 1860 -2202 1861 -2201
rect 2368 -2202 2369 -2201
rect 107 -2204 108 -2203
rect 128 -2204 129 -2203
rect 131 -2204 132 -2203
rect 257 -2204 258 -2203
rect 296 -2204 297 -2203
rect 656 -2204 657 -2203
rect 674 -2204 675 -2203
rect 1895 -2204 1896 -2203
rect 1927 -2204 1928 -2203
rect 1990 -2204 1991 -2203
rect 2032 -2204 2033 -2203
rect 2102 -2204 2103 -2203
rect 107 -2206 108 -2205
rect 506 -2206 507 -2205
rect 527 -2206 528 -2205
rect 1384 -2206 1385 -2205
rect 1416 -2206 1417 -2205
rect 1493 -2206 1494 -2205
rect 1521 -2206 1522 -2205
rect 1626 -2206 1627 -2205
rect 1629 -2206 1630 -2205
rect 2249 -2206 2250 -2205
rect 121 -2208 122 -2207
rect 1710 -2208 1711 -2207
rect 1843 -2208 1844 -2207
rect 1906 -2208 1907 -2207
rect 1962 -2208 1963 -2207
rect 2025 -2208 2026 -2207
rect 2060 -2208 2061 -2207
rect 2228 -2208 2229 -2207
rect 16 -2210 17 -2209
rect 121 -2210 122 -2209
rect 124 -2210 125 -2209
rect 387 -2210 388 -2209
rect 450 -2210 451 -2209
rect 495 -2210 496 -2209
rect 506 -2210 507 -2209
rect 779 -2210 780 -2209
rect 782 -2210 783 -2209
rect 992 -2210 993 -2209
rect 996 -2210 997 -2209
rect 1941 -2210 1942 -2209
rect 1983 -2210 1984 -2209
rect 2046 -2210 2047 -2209
rect 2060 -2210 2061 -2209
rect 2130 -2210 2131 -2209
rect 16 -2212 17 -2211
rect 86 -2212 87 -2211
rect 128 -2212 129 -2211
rect 1188 -2212 1189 -2211
rect 1192 -2212 1193 -2211
rect 1269 -2212 1270 -2211
rect 1332 -2212 1333 -2211
rect 1346 -2212 1347 -2211
rect 1367 -2212 1368 -2211
rect 1535 -2212 1536 -2211
rect 1545 -2212 1546 -2211
rect 2347 -2212 2348 -2211
rect 86 -2214 87 -2213
rect 625 -2214 626 -2213
rect 681 -2214 682 -2213
rect 744 -2214 745 -2213
rect 800 -2214 801 -2213
rect 1185 -2214 1186 -2213
rect 1202 -2214 1203 -2213
rect 1276 -2214 1277 -2213
rect 1283 -2214 1284 -2213
rect 1346 -2214 1347 -2213
rect 1381 -2214 1382 -2213
rect 1549 -2214 1550 -2213
rect 1580 -2214 1581 -2213
rect 2116 -2214 2117 -2213
rect 2130 -2214 2131 -2213
rect 2256 -2214 2257 -2213
rect 138 -2216 139 -2215
rect 2263 -2216 2264 -2215
rect 145 -2218 146 -2217
rect 856 -2218 857 -2217
rect 877 -2218 878 -2217
rect 1503 -2218 1504 -2217
rect 1517 -2218 1518 -2217
rect 2347 -2218 2348 -2217
rect 166 -2220 167 -2219
rect 2207 -2220 2208 -2219
rect 2256 -2220 2257 -2219
rect 2354 -2220 2355 -2219
rect 236 -2222 237 -2221
rect 940 -2222 941 -2221
rect 975 -2222 976 -2221
rect 1759 -2222 1760 -2221
rect 1783 -2222 1784 -2221
rect 1906 -2222 1907 -2221
rect 1941 -2222 1942 -2221
rect 1997 -2222 1998 -2221
rect 2025 -2222 2026 -2221
rect 2088 -2222 2089 -2221
rect 2102 -2222 2103 -2221
rect 2200 -2222 2201 -2221
rect 2207 -2222 2208 -2221
rect 2340 -2222 2341 -2221
rect 243 -2224 244 -2223
rect 884 -2224 885 -2223
rect 912 -2224 913 -2223
rect 1010 -2224 1011 -2223
rect 1094 -2224 1095 -2223
rect 1171 -2224 1172 -2223
rect 1185 -2224 1186 -2223
rect 1262 -2224 1263 -2223
rect 1269 -2224 1270 -2223
rect 1290 -2224 1291 -2223
rect 1342 -2224 1343 -2223
rect 1430 -2224 1431 -2223
rect 1479 -2224 1480 -2223
rect 1787 -2224 1788 -2223
rect 1871 -2224 1872 -2223
rect 1948 -2224 1949 -2223
rect 1990 -2224 1991 -2223
rect 2053 -2224 2054 -2223
rect 2088 -2224 2089 -2223
rect 2165 -2224 2166 -2223
rect 2200 -2224 2201 -2223
rect 2333 -2224 2334 -2223
rect 156 -2226 157 -2225
rect 1171 -2226 1172 -2225
rect 1220 -2226 1221 -2225
rect 2284 -2226 2285 -2225
rect 40 -2228 41 -2227
rect 156 -2228 157 -2227
rect 250 -2228 251 -2227
rect 1220 -2228 1221 -2227
rect 1227 -2228 1228 -2227
rect 1451 -2228 1452 -2227
rect 1535 -2228 1536 -2227
rect 1668 -2228 1669 -2227
rect 1759 -2228 1760 -2227
rect 1815 -2228 1816 -2227
rect 1934 -2228 1935 -2227
rect 2165 -2228 2166 -2227
rect 2186 -2228 2187 -2227
rect 2284 -2228 2285 -2227
rect 289 -2230 290 -2229
rect 779 -2230 780 -2229
rect 821 -2230 822 -2229
rect 926 -2230 927 -2229
rect 940 -2230 941 -2229
rect 954 -2230 955 -2229
rect 975 -2230 976 -2229
rect 1979 -2230 1980 -2229
rect 1997 -2230 1998 -2229
rect 2067 -2230 2068 -2229
rect 2116 -2230 2117 -2229
rect 2221 -2230 2222 -2229
rect 289 -2232 290 -2231
rect 352 -2232 353 -2231
rect 359 -2232 360 -2231
rect 1055 -2232 1056 -2231
rect 1101 -2232 1102 -2231
rect 1129 -2232 1130 -2231
rect 1136 -2232 1137 -2231
rect 1332 -2232 1333 -2231
rect 1381 -2232 1382 -2231
rect 1465 -2232 1466 -2231
rect 1549 -2232 1550 -2231
rect 1591 -2232 1592 -2231
rect 1647 -2232 1648 -2231
rect 2263 -2232 2264 -2231
rect 261 -2234 262 -2233
rect 359 -2234 360 -2233
rect 457 -2234 458 -2233
rect 516 -2234 517 -2233
rect 527 -2234 528 -2233
rect 583 -2234 584 -2233
rect 590 -2234 591 -2233
rect 954 -2234 955 -2233
rect 978 -2234 979 -2233
rect 2312 -2234 2313 -2233
rect 100 -2236 101 -2235
rect 261 -2236 262 -2235
rect 296 -2236 297 -2235
rect 604 -2236 605 -2235
rect 618 -2236 619 -2235
rect 667 -2236 668 -2235
rect 681 -2236 682 -2235
rect 709 -2236 710 -2235
rect 726 -2236 727 -2235
rect 2172 -2236 2173 -2235
rect 2186 -2236 2187 -2235
rect 2417 -2236 2418 -2235
rect 100 -2238 101 -2237
rect 1017 -2238 1018 -2237
rect 1115 -2238 1116 -2237
rect 1696 -2238 1697 -2237
rect 1787 -2238 1788 -2237
rect 1850 -2238 1851 -2237
rect 1934 -2238 1935 -2237
rect 2179 -2238 2180 -2237
rect 2221 -2238 2222 -2237
rect 2319 -2238 2320 -2237
rect 170 -2240 171 -2239
rect 457 -2240 458 -2239
rect 492 -2240 493 -2239
rect 1073 -2240 1074 -2239
rect 1129 -2240 1130 -2239
rect 1164 -2240 1165 -2239
rect 1248 -2240 1249 -2239
rect 1360 -2240 1361 -2239
rect 1423 -2240 1424 -2239
rect 1451 -2240 1452 -2239
rect 1465 -2240 1466 -2239
rect 1570 -2240 1571 -2239
rect 1591 -2240 1592 -2239
rect 1689 -2240 1690 -2239
rect 1703 -2240 1704 -2239
rect 1850 -2240 1851 -2239
rect 1948 -2240 1949 -2239
rect 2004 -2240 2005 -2239
rect 2046 -2240 2047 -2239
rect 2333 -2240 2334 -2239
rect 79 -2242 80 -2241
rect 492 -2242 493 -2241
rect 555 -2242 556 -2241
rect 1230 -2242 1231 -2241
rect 1248 -2242 1249 -2241
rect 2270 -2242 2271 -2241
rect 79 -2244 80 -2243
rect 639 -2244 640 -2243
rect 653 -2244 654 -2243
rect 1136 -2244 1137 -2243
rect 1143 -2244 1144 -2243
rect 1206 -2244 1207 -2243
rect 1255 -2244 1256 -2243
rect 1374 -2244 1375 -2243
rect 1423 -2244 1424 -2243
rect 1514 -2244 1515 -2243
rect 1570 -2244 1571 -2243
rect 1661 -2244 1662 -2243
rect 1682 -2244 1683 -2243
rect 1815 -2244 1816 -2243
rect 1857 -2244 1858 -2243
rect 2004 -2244 2005 -2243
rect 2053 -2244 2054 -2243
rect 2123 -2244 2124 -2243
rect 2179 -2244 2180 -2243
rect 2291 -2244 2292 -2243
rect 170 -2246 171 -2245
rect 177 -2246 178 -2245
rect 338 -2246 339 -2245
rect 450 -2246 451 -2245
rect 576 -2246 577 -2245
rect 618 -2246 619 -2245
rect 621 -2246 622 -2245
rect 1577 -2246 1578 -2245
rect 1605 -2246 1606 -2245
rect 1689 -2246 1690 -2245
rect 1703 -2246 1704 -2245
rect 1766 -2246 1767 -2245
rect 1857 -2246 1858 -2245
rect 1920 -2246 1921 -2245
rect 2067 -2246 2068 -2245
rect 2137 -2246 2138 -2245
rect 177 -2248 178 -2247
rect 1685 -2248 1686 -2247
rect 1766 -2248 1767 -2247
rect 1822 -2248 1823 -2247
rect 2123 -2248 2124 -2247
rect 2235 -2248 2236 -2247
rect 317 -2250 318 -2249
rect 338 -2250 339 -2249
rect 352 -2250 353 -2249
rect 366 -2250 367 -2249
rect 394 -2250 395 -2249
rect 555 -2250 556 -2249
rect 583 -2250 584 -2249
rect 597 -2250 598 -2249
rect 604 -2250 605 -2249
rect 695 -2250 696 -2249
rect 709 -2250 710 -2249
rect 919 -2250 920 -2249
rect 978 -2250 979 -2249
rect 2291 -2250 2292 -2249
rect 275 -2252 276 -2251
rect 597 -2252 598 -2251
rect 639 -2252 640 -2251
rect 891 -2252 892 -2251
rect 912 -2252 913 -2251
rect 989 -2252 990 -2251
rect 1073 -2252 1074 -2251
rect 1122 -2252 1123 -2251
rect 1164 -2252 1165 -2251
rect 1241 -2252 1242 -2251
rect 1262 -2252 1263 -2251
rect 1395 -2252 1396 -2251
rect 1430 -2252 1431 -2251
rect 1500 -2252 1501 -2251
rect 1605 -2252 1606 -2251
rect 1640 -2252 1641 -2251
rect 1647 -2252 1648 -2251
rect 1808 -2252 1809 -2251
rect 2074 -2252 2075 -2251
rect 2235 -2252 2236 -2251
rect 275 -2254 276 -2253
rect 625 -2254 626 -2253
rect 688 -2254 689 -2253
rect 821 -2254 822 -2253
rect 828 -2254 829 -2253
rect 884 -2254 885 -2253
rect 982 -2254 983 -2253
rect 1045 -2254 1046 -2253
rect 1087 -2254 1088 -2253
rect 1122 -2254 1123 -2253
rect 1178 -2254 1179 -2253
rect 1241 -2254 1242 -2253
rect 1283 -2254 1284 -2253
rect 1318 -2254 1319 -2253
rect 1339 -2254 1340 -2253
rect 1822 -2254 1823 -2253
rect 2018 -2254 2019 -2253
rect 2074 -2254 2075 -2253
rect 310 -2256 311 -2255
rect 317 -2256 318 -2255
rect 324 -2256 325 -2255
rect 394 -2256 395 -2255
rect 443 -2256 444 -2255
rect 891 -2256 892 -2255
rect 961 -2256 962 -2255
rect 1087 -2256 1088 -2255
rect 1178 -2256 1179 -2255
rect 1444 -2256 1445 -2255
rect 1486 -2256 1487 -2255
rect 1920 -2256 1921 -2255
rect 2018 -2256 2019 -2255
rect 2361 -2256 2362 -2255
rect 114 -2258 115 -2257
rect 324 -2258 325 -2257
rect 366 -2258 367 -2257
rect 663 -2258 664 -2257
rect 695 -2258 696 -2257
rect 1307 -2258 1308 -2257
rect 1318 -2258 1319 -2257
rect 2410 -2258 2411 -2257
rect 114 -2260 115 -2259
rect 226 -2260 227 -2259
rect 310 -2260 311 -2259
rect 541 -2260 542 -2259
rect 590 -2260 591 -2259
rect 870 -2260 871 -2259
rect 933 -2260 934 -2259
rect 961 -2260 962 -2259
rect 989 -2260 990 -2259
rect 2424 -2260 2425 -2259
rect 163 -2262 164 -2261
rect 226 -2262 227 -2261
rect 380 -2262 381 -2261
rect 688 -2262 689 -2261
rect 751 -2262 752 -2261
rect 1017 -2262 1018 -2261
rect 1206 -2262 1207 -2261
rect 1297 -2262 1298 -2261
rect 1339 -2262 1340 -2261
rect 1458 -2262 1459 -2261
rect 1472 -2262 1473 -2261
rect 1486 -2262 1487 -2261
rect 1500 -2262 1501 -2261
rect 2382 -2262 2383 -2261
rect 163 -2264 164 -2263
rect 2249 -2264 2250 -2263
rect 380 -2266 381 -2265
rect 835 -2266 836 -2265
rect 856 -2266 857 -2265
rect 1976 -2266 1977 -2265
rect 443 -2268 444 -2267
rect 471 -2268 472 -2267
rect 478 -2268 479 -2267
rect 576 -2268 577 -2267
rect 593 -2268 594 -2267
rect 2039 -2268 2040 -2267
rect 142 -2270 143 -2269
rect 471 -2270 472 -2269
rect 478 -2270 479 -2269
rect 919 -2270 920 -2269
rect 1290 -2270 1291 -2269
rect 1913 -2270 1914 -2269
rect 2039 -2270 2040 -2269
rect 2109 -2270 2110 -2269
rect 142 -2272 143 -2271
rect 254 -2272 255 -2271
rect 513 -2272 514 -2271
rect 870 -2272 871 -2271
rect 1297 -2272 1298 -2271
rect 1353 -2272 1354 -2271
rect 1370 -2272 1371 -2271
rect 1458 -2272 1459 -2271
rect 1472 -2272 1473 -2271
rect 1955 -2272 1956 -2271
rect 2109 -2272 2110 -2271
rect 2214 -2272 2215 -2271
rect 513 -2274 514 -2273
rect 534 -2274 535 -2273
rect 541 -2274 542 -2273
rect 548 -2274 549 -2273
rect 737 -2274 738 -2273
rect 751 -2274 752 -2273
rect 758 -2274 759 -2273
rect 1668 -2274 1669 -2273
rect 1808 -2274 1809 -2273
rect 2011 -2274 2012 -2273
rect 2095 -2274 2096 -2273
rect 2214 -2274 2215 -2273
rect 422 -2276 423 -2275
rect 534 -2276 535 -2275
rect 548 -2276 549 -2275
rect 716 -2276 717 -2275
rect 758 -2276 759 -2275
rect 863 -2276 864 -2275
rect 1353 -2276 1354 -2275
rect 1528 -2276 1529 -2275
rect 1563 -2276 1564 -2275
rect 1955 -2276 1956 -2275
rect 2011 -2276 2012 -2275
rect 2081 -2276 2082 -2275
rect 2095 -2276 2096 -2275
rect 2193 -2276 2194 -2275
rect 184 -2278 185 -2277
rect 716 -2278 717 -2277
rect 765 -2278 766 -2277
rect 877 -2278 878 -2277
rect 1059 -2278 1060 -2277
rect 1528 -2278 1529 -2277
rect 1563 -2278 1564 -2277
rect 1654 -2278 1655 -2277
rect 1661 -2278 1662 -2277
rect 1738 -2278 1739 -2277
rect 1892 -2278 1893 -2277
rect 1913 -2278 1914 -2277
rect 2081 -2278 2082 -2277
rect 2158 -2278 2159 -2277
rect 149 -2280 150 -2279
rect 184 -2280 185 -2279
rect 219 -2280 220 -2279
rect 422 -2280 423 -2279
rect 485 -2280 486 -2279
rect 737 -2280 738 -2279
rect 772 -2280 773 -2279
rect 800 -2280 801 -2279
rect 814 -2280 815 -2279
rect 863 -2280 864 -2279
rect 1059 -2280 1060 -2279
rect 1335 -2280 1336 -2279
rect 1374 -2280 1375 -2279
rect 1542 -2280 1543 -2279
rect 1619 -2280 1620 -2279
rect 1696 -2280 1697 -2279
rect 1738 -2280 1739 -2279
rect 1794 -2280 1795 -2279
rect 135 -2282 136 -2281
rect 149 -2282 150 -2281
rect 191 -2282 192 -2281
rect 219 -2282 220 -2281
rect 373 -2282 374 -2281
rect 765 -2282 766 -2281
rect 786 -2282 787 -2281
rect 2319 -2282 2320 -2281
rect 135 -2284 136 -2283
rect 569 -2284 570 -2283
rect 611 -2284 612 -2283
rect 814 -2284 815 -2283
rect 828 -2284 829 -2283
rect 842 -2284 843 -2283
rect 859 -2284 860 -2283
rect 2137 -2284 2138 -2283
rect 191 -2286 192 -2285
rect 1066 -2286 1067 -2285
rect 1321 -2286 1322 -2285
rect 2193 -2286 2194 -2285
rect 373 -2288 374 -2287
rect 520 -2288 521 -2287
rect 569 -2288 570 -2287
rect 723 -2288 724 -2287
rect 786 -2288 787 -2287
rect 1003 -2288 1004 -2287
rect 1066 -2288 1067 -2287
rect 1108 -2288 1109 -2287
rect 1395 -2288 1396 -2287
rect 1976 -2288 1977 -2287
rect 415 -2290 416 -2289
rect 520 -2290 521 -2289
rect 646 -2290 647 -2289
rect 772 -2290 773 -2289
rect 807 -2290 808 -2289
rect 842 -2290 843 -2289
rect 968 -2290 969 -2289
rect 1542 -2290 1543 -2289
rect 1619 -2290 1620 -2289
rect 1717 -2290 1718 -2289
rect 1794 -2290 1795 -2289
rect 1864 -2290 1865 -2289
rect 331 -2292 332 -2291
rect 415 -2292 416 -2291
rect 436 -2292 437 -2291
rect 485 -2292 486 -2291
rect 499 -2292 500 -2291
rect 611 -2292 612 -2291
rect 646 -2292 647 -2291
rect 660 -2292 661 -2291
rect 723 -2292 724 -2291
rect 982 -2292 983 -2291
rect 1052 -2292 1053 -2291
rect 1108 -2292 1109 -2291
rect 1402 -2292 1403 -2291
rect 2158 -2292 2159 -2291
rect 233 -2294 234 -2293
rect 499 -2294 500 -2293
rect 562 -2294 563 -2293
rect 1402 -2294 1403 -2293
rect 1409 -2294 1410 -2293
rect 1864 -2294 1865 -2293
rect 233 -2296 234 -2295
rect 705 -2296 706 -2295
rect 730 -2296 731 -2295
rect 1052 -2296 1053 -2295
rect 1409 -2296 1410 -2295
rect 1626 -2296 1627 -2295
rect 1633 -2296 1634 -2295
rect 1717 -2296 1718 -2295
rect 268 -2298 269 -2297
rect 436 -2298 437 -2297
rect 730 -2298 731 -2297
rect 898 -2298 899 -2297
rect 905 -2298 906 -2297
rect 968 -2298 969 -2297
rect 1444 -2298 1445 -2297
rect 1584 -2298 1585 -2297
rect 1633 -2298 1634 -2297
rect 1724 -2298 1725 -2297
rect 205 -2300 206 -2299
rect 898 -2300 899 -2299
rect 905 -2300 906 -2299
rect 1325 -2300 1326 -2299
rect 1584 -2300 1585 -2299
rect 1675 -2300 1676 -2299
rect 44 -2302 45 -2301
rect 205 -2302 206 -2301
rect 212 -2302 213 -2301
rect 268 -2302 269 -2301
rect 331 -2302 332 -2301
rect 345 -2302 346 -2301
rect 429 -2302 430 -2301
rect 562 -2302 563 -2301
rect 747 -2302 748 -2301
rect 1003 -2302 1004 -2301
rect 1024 -2302 1025 -2301
rect 1724 -2302 1725 -2301
rect 44 -2304 45 -2303
rect 58 -2304 59 -2303
rect 72 -2304 73 -2303
rect 1024 -2304 1025 -2303
rect 1325 -2304 1326 -2303
rect 1612 -2304 1613 -2303
rect 1640 -2304 1641 -2303
rect 1731 -2304 1732 -2303
rect 23 -2306 24 -2305
rect 58 -2306 59 -2305
rect 72 -2306 73 -2305
rect 401 -2306 402 -2305
rect 807 -2306 808 -2305
rect 849 -2306 850 -2305
rect 1507 -2306 1508 -2305
rect 1612 -2306 1613 -2305
rect 1650 -2306 1651 -2305
rect 2326 -2306 2327 -2305
rect 23 -2308 24 -2307
rect 198 -2308 199 -2307
rect 212 -2308 213 -2307
rect 247 -2308 248 -2307
rect 282 -2308 283 -2307
rect 345 -2308 346 -2307
rect 401 -2308 402 -2307
rect 464 -2308 465 -2307
rect 835 -2308 836 -2307
rect 1213 -2308 1214 -2307
rect 1507 -2308 1508 -2307
rect 1556 -2308 1557 -2307
rect 1675 -2308 1676 -2307
rect 1745 -2308 1746 -2307
rect 2277 -2308 2278 -2307
rect 2326 -2308 2327 -2307
rect 198 -2310 199 -2309
rect 670 -2310 671 -2309
rect 793 -2310 794 -2309
rect 1213 -2310 1214 -2309
rect 1556 -2310 1557 -2309
rect 1598 -2310 1599 -2309
rect 1731 -2310 1732 -2309
rect 2144 -2310 2145 -2309
rect 2277 -2310 2278 -2309
rect 2389 -2310 2390 -2309
rect 247 -2312 248 -2311
rect 429 -2312 430 -2311
rect 464 -2312 465 -2311
rect 632 -2312 633 -2311
rect 789 -2312 790 -2311
rect 1598 -2312 1599 -2311
rect 1745 -2312 1746 -2311
rect 1801 -2312 1802 -2311
rect 2144 -2312 2145 -2311
rect 2242 -2312 2243 -2311
rect 282 -2314 283 -2313
rect 303 -2314 304 -2313
rect 387 -2314 388 -2313
rect 670 -2314 671 -2313
rect 793 -2314 794 -2313
rect 1493 -2314 1494 -2313
rect 1801 -2314 1802 -2313
rect 1878 -2314 1879 -2313
rect 2242 -2314 2243 -2313
rect 2375 -2314 2376 -2313
rect 303 -2316 304 -2315
rect 408 -2316 409 -2315
rect 632 -2316 633 -2315
rect 702 -2316 703 -2315
rect 849 -2316 850 -2315
rect 1311 -2316 1312 -2315
rect 1773 -2316 1774 -2315
rect 1878 -2316 1879 -2315
rect 30 -2318 31 -2317
rect 408 -2318 409 -2317
rect 660 -2318 661 -2317
rect 1311 -2318 1312 -2317
rect 1773 -2318 1774 -2317
rect 1829 -2318 1830 -2317
rect 702 -2320 703 -2319
rect 1654 -2320 1655 -2319
rect 1829 -2320 1830 -2319
rect 1899 -2320 1900 -2319
rect 1199 -2322 1200 -2321
rect 1899 -2322 1900 -2321
rect 33 -2324 34 -2323
rect 1199 -2324 1200 -2323
rect 5 -2335 6 -2334
rect 65 -2335 66 -2334
rect 163 -2335 164 -2334
rect 1024 -2335 1025 -2334
rect 1038 -2335 1039 -2334
rect 1360 -2335 1361 -2334
rect 1363 -2335 1364 -2334
rect 2221 -2335 2222 -2334
rect 2326 -2335 2327 -2334
rect 2343 -2335 2344 -2334
rect 9 -2337 10 -2336
rect 873 -2337 874 -2336
rect 905 -2337 906 -2336
rect 1248 -2337 1249 -2336
rect 1272 -2337 1273 -2336
rect 2074 -2337 2075 -2336
rect 2165 -2337 2166 -2336
rect 2333 -2337 2334 -2336
rect 23 -2339 24 -2338
rect 145 -2339 146 -2338
rect 170 -2339 171 -2338
rect 173 -2339 174 -2338
rect 226 -2339 227 -2338
rect 593 -2339 594 -2338
rect 597 -2339 598 -2338
rect 726 -2339 727 -2338
rect 782 -2339 783 -2338
rect 1535 -2339 1536 -2338
rect 1542 -2339 1543 -2338
rect 1878 -2339 1879 -2338
rect 1892 -2339 1893 -2338
rect 1948 -2339 1949 -2338
rect 1976 -2339 1977 -2338
rect 2039 -2339 2040 -2338
rect 2165 -2339 2166 -2338
rect 2193 -2339 2194 -2338
rect 2221 -2339 2222 -2338
rect 2242 -2339 2243 -2338
rect 16 -2341 17 -2340
rect 226 -2341 227 -2340
rect 240 -2341 241 -2340
rect 607 -2341 608 -2340
rect 618 -2341 619 -2340
rect 1318 -2341 1319 -2340
rect 1374 -2341 1375 -2340
rect 1395 -2341 1396 -2340
rect 1398 -2341 1399 -2340
rect 1409 -2341 1410 -2340
rect 1493 -2341 1494 -2340
rect 2235 -2341 2236 -2340
rect 2242 -2341 2243 -2340
rect 2291 -2341 2292 -2340
rect 16 -2343 17 -2342
rect 37 -2343 38 -2342
rect 51 -2343 52 -2342
rect 1024 -2343 1025 -2342
rect 1041 -2343 1042 -2342
rect 1493 -2343 1494 -2342
rect 1517 -2343 1518 -2342
rect 1906 -2343 1907 -2342
rect 1934 -2343 1935 -2342
rect 2284 -2343 2285 -2342
rect 30 -2345 31 -2344
rect 1080 -2345 1081 -2344
rect 1108 -2345 1109 -2344
rect 1979 -2345 1980 -2344
rect 2039 -2345 2040 -2344
rect 2088 -2345 2089 -2344
rect 2186 -2345 2187 -2344
rect 2291 -2345 2292 -2344
rect 33 -2347 34 -2346
rect 44 -2347 45 -2346
rect 51 -2347 52 -2346
rect 1577 -2347 1578 -2346
rect 1580 -2347 1581 -2346
rect 2256 -2347 2257 -2346
rect 44 -2349 45 -2348
rect 114 -2349 115 -2348
rect 170 -2349 171 -2348
rect 177 -2349 178 -2348
rect 243 -2349 244 -2348
rect 506 -2349 507 -2348
rect 569 -2349 570 -2348
rect 618 -2349 619 -2348
rect 625 -2349 626 -2348
rect 891 -2349 892 -2348
rect 905 -2349 906 -2348
rect 940 -2349 941 -2348
rect 954 -2349 955 -2348
rect 1321 -2349 1322 -2348
rect 1377 -2349 1378 -2348
rect 1451 -2349 1452 -2348
rect 1542 -2349 1543 -2348
rect 1598 -2349 1599 -2348
rect 1682 -2349 1683 -2348
rect 2228 -2349 2229 -2348
rect 2235 -2349 2236 -2348
rect 2277 -2349 2278 -2348
rect 65 -2351 66 -2350
rect 275 -2351 276 -2350
rect 282 -2351 283 -2350
rect 1076 -2351 1077 -2350
rect 1080 -2351 1081 -2350
rect 1612 -2351 1613 -2350
rect 1682 -2351 1683 -2350
rect 1745 -2351 1746 -2350
rect 1850 -2351 1851 -2350
rect 1853 -2351 1854 -2350
rect 1878 -2351 1879 -2350
rect 2102 -2351 2103 -2350
rect 2179 -2351 2180 -2350
rect 2186 -2351 2187 -2350
rect 2193 -2351 2194 -2350
rect 2207 -2351 2208 -2350
rect 2228 -2351 2229 -2350
rect 2263 -2351 2264 -2350
rect 114 -2353 115 -2352
rect 261 -2353 262 -2352
rect 275 -2353 276 -2352
rect 387 -2353 388 -2352
rect 408 -2353 409 -2352
rect 765 -2353 766 -2352
rect 775 -2353 776 -2352
rect 940 -2353 941 -2352
rect 978 -2353 979 -2352
rect 1213 -2353 1214 -2352
rect 1248 -2353 1249 -2352
rect 1262 -2353 1263 -2352
rect 1276 -2353 1277 -2352
rect 1356 -2353 1357 -2352
rect 1451 -2353 1452 -2352
rect 1528 -2353 1529 -2352
rect 1685 -2353 1686 -2352
rect 2158 -2353 2159 -2352
rect 2207 -2353 2208 -2352
rect 2280 -2353 2281 -2352
rect 166 -2355 167 -2354
rect 2179 -2355 2180 -2354
rect 2256 -2355 2257 -2354
rect 2312 -2355 2313 -2354
rect 247 -2357 248 -2356
rect 842 -2357 843 -2356
rect 859 -2357 860 -2356
rect 1612 -2357 1613 -2356
rect 1745 -2357 1746 -2356
rect 1773 -2357 1774 -2356
rect 1850 -2357 1851 -2356
rect 1885 -2357 1886 -2356
rect 1895 -2357 1896 -2356
rect 2214 -2357 2215 -2356
rect 2263 -2357 2264 -2356
rect 2319 -2357 2320 -2356
rect 247 -2359 248 -2358
rect 478 -2359 479 -2358
rect 481 -2359 482 -2358
rect 1629 -2359 1630 -2358
rect 1773 -2359 1774 -2358
rect 1787 -2359 1788 -2358
rect 1885 -2359 1886 -2358
rect 1941 -2359 1942 -2358
rect 1948 -2359 1949 -2358
rect 2116 -2359 2117 -2358
rect 261 -2361 262 -2360
rect 401 -2361 402 -2360
rect 408 -2361 409 -2360
rect 485 -2361 486 -2360
rect 492 -2361 493 -2360
rect 506 -2361 507 -2360
rect 527 -2361 528 -2360
rect 569 -2361 570 -2360
rect 576 -2361 577 -2360
rect 779 -2361 780 -2360
rect 786 -2361 787 -2360
rect 954 -2361 955 -2360
rect 982 -2361 983 -2360
rect 1038 -2361 1039 -2360
rect 1055 -2361 1056 -2360
rect 1486 -2361 1487 -2360
rect 1528 -2361 1529 -2360
rect 1591 -2361 1592 -2360
rect 1787 -2361 1788 -2360
rect 1843 -2361 1844 -2360
rect 1853 -2361 1854 -2360
rect 1941 -2361 1942 -2360
rect 2011 -2361 2012 -2360
rect 2116 -2361 2117 -2360
rect 282 -2363 283 -2362
rect 835 -2363 836 -2362
rect 842 -2363 843 -2362
rect 912 -2363 913 -2362
rect 919 -2363 920 -2362
rect 1696 -2363 1697 -2362
rect 1843 -2363 1844 -2362
rect 1857 -2363 1858 -2362
rect 1906 -2363 1907 -2362
rect 1927 -2363 1928 -2362
rect 1934 -2363 1935 -2362
rect 1997 -2363 1998 -2362
rect 2011 -2363 2012 -2362
rect 2067 -2363 2068 -2362
rect 2088 -2363 2089 -2362
rect 2305 -2363 2306 -2362
rect 296 -2365 297 -2364
rect 723 -2365 724 -2364
rect 730 -2365 731 -2364
rect 1409 -2365 1410 -2364
rect 1486 -2365 1487 -2364
rect 1570 -2365 1571 -2364
rect 1591 -2365 1592 -2364
rect 1822 -2365 1823 -2364
rect 1836 -2365 1837 -2364
rect 1857 -2365 1858 -2364
rect 1927 -2365 1928 -2364
rect 1990 -2365 1991 -2364
rect 1997 -2365 1998 -2364
rect 2060 -2365 2061 -2364
rect 2102 -2365 2103 -2364
rect 2130 -2365 2131 -2364
rect 2305 -2365 2306 -2364
rect 2347 -2365 2348 -2364
rect 191 -2367 192 -2366
rect 723 -2367 724 -2366
rect 730 -2367 731 -2366
rect 793 -2367 794 -2366
rect 796 -2367 797 -2366
rect 1668 -2367 1669 -2366
rect 1678 -2367 1679 -2366
rect 1696 -2367 1697 -2366
rect 1836 -2367 1837 -2366
rect 1983 -2367 1984 -2366
rect 1990 -2367 1991 -2366
rect 2123 -2367 2124 -2366
rect 72 -2369 73 -2368
rect 191 -2369 192 -2368
rect 296 -2369 297 -2368
rect 1052 -2369 1053 -2368
rect 1108 -2369 1109 -2368
rect 1150 -2369 1151 -2368
rect 1262 -2369 1263 -2368
rect 1304 -2369 1305 -2368
rect 1318 -2369 1319 -2368
rect 1381 -2369 1382 -2368
rect 1668 -2369 1669 -2368
rect 1738 -2369 1739 -2368
rect 1983 -2369 1984 -2368
rect 2053 -2369 2054 -2368
rect 2060 -2369 2061 -2368
rect 2109 -2369 2110 -2368
rect 2123 -2369 2124 -2368
rect 2137 -2369 2138 -2368
rect 310 -2371 311 -2370
rect 429 -2371 430 -2370
rect 457 -2371 458 -2370
rect 856 -2371 857 -2370
rect 859 -2371 860 -2370
rect 1332 -2371 1333 -2370
rect 1381 -2371 1382 -2370
rect 1437 -2371 1438 -2370
rect 1738 -2371 1739 -2370
rect 1766 -2371 1767 -2370
rect 1969 -2371 1970 -2370
rect 2109 -2371 2110 -2370
rect 2137 -2371 2138 -2370
rect 2151 -2371 2152 -2370
rect 268 -2373 269 -2372
rect 310 -2373 311 -2372
rect 387 -2373 388 -2372
rect 856 -2373 857 -2372
rect 863 -2373 864 -2372
rect 982 -2373 983 -2372
rect 1052 -2373 1053 -2372
rect 2074 -2373 2075 -2372
rect 2151 -2373 2152 -2372
rect 2172 -2373 2173 -2372
rect 401 -2375 402 -2374
rect 681 -2375 682 -2374
rect 716 -2375 717 -2374
rect 2067 -2375 2068 -2374
rect 2172 -2375 2173 -2374
rect 2200 -2375 2201 -2374
rect 37 -2377 38 -2376
rect 2200 -2377 2201 -2376
rect 100 -2379 101 -2378
rect 716 -2379 717 -2378
rect 786 -2379 787 -2378
rect 1164 -2379 1165 -2378
rect 1227 -2379 1228 -2378
rect 1304 -2379 1305 -2378
rect 1437 -2379 1438 -2378
rect 1444 -2379 1445 -2378
rect 1766 -2379 1767 -2378
rect 1829 -2379 1830 -2378
rect 2018 -2379 2019 -2378
rect 2214 -2379 2215 -2378
rect 100 -2381 101 -2380
rect 961 -2381 962 -2380
rect 1087 -2381 1088 -2380
rect 1164 -2381 1165 -2380
rect 1227 -2381 1228 -2380
rect 1255 -2381 1256 -2380
rect 1276 -2381 1277 -2380
rect 1545 -2381 1546 -2380
rect 1647 -2381 1648 -2380
rect 1829 -2381 1830 -2380
rect 2046 -2381 2047 -2380
rect 2284 -2381 2285 -2380
rect 422 -2383 423 -2382
rect 768 -2383 769 -2382
rect 821 -2383 822 -2382
rect 978 -2383 979 -2382
rect 1087 -2383 1088 -2382
rect 1129 -2383 1130 -2382
rect 1136 -2383 1137 -2382
rect 1297 -2383 1298 -2382
rect 1444 -2383 1445 -2382
rect 1479 -2383 1480 -2382
rect 1549 -2383 1550 -2382
rect 1647 -2383 1648 -2382
rect 1801 -2383 1802 -2382
rect 1969 -2383 1970 -2382
rect 2053 -2383 2054 -2382
rect 2095 -2383 2096 -2382
rect 110 -2385 111 -2384
rect 1136 -2385 1137 -2384
rect 1150 -2385 1151 -2384
rect 1185 -2385 1186 -2384
rect 1293 -2385 1294 -2384
rect 1752 -2385 1753 -2384
rect 1899 -2385 1900 -2384
rect 2095 -2385 2096 -2384
rect 324 -2387 325 -2386
rect 422 -2387 423 -2386
rect 457 -2387 458 -2386
rect 646 -2387 647 -2386
rect 660 -2387 661 -2386
rect 758 -2387 759 -2386
rect 821 -2387 822 -2386
rect 877 -2387 878 -2386
rect 884 -2387 885 -2386
rect 891 -2387 892 -2386
rect 912 -2387 913 -2386
rect 1335 -2387 1336 -2386
rect 1479 -2387 1480 -2386
rect 1703 -2387 1704 -2386
rect 1752 -2387 1753 -2386
rect 1780 -2387 1781 -2386
rect 1801 -2387 1802 -2386
rect 1899 -2387 1900 -2386
rect 324 -2389 325 -2388
rect 394 -2389 395 -2388
rect 464 -2389 465 -2388
rect 485 -2389 486 -2388
rect 492 -2389 493 -2388
rect 1311 -2389 1312 -2388
rect 1465 -2389 1466 -2388
rect 1780 -2389 1781 -2388
rect 303 -2391 304 -2390
rect 394 -2391 395 -2390
rect 464 -2391 465 -2390
rect 1017 -2391 1018 -2390
rect 1115 -2391 1116 -2390
rect 1535 -2391 1536 -2390
rect 1703 -2391 1704 -2390
rect 1717 -2391 1718 -2390
rect 303 -2393 304 -2392
rect 331 -2393 332 -2392
rect 520 -2393 521 -2392
rect 681 -2393 682 -2392
rect 702 -2393 703 -2392
rect 1185 -2393 1186 -2392
rect 1311 -2393 1312 -2392
rect 1339 -2393 1340 -2392
rect 1710 -2393 1711 -2392
rect 1717 -2393 1718 -2392
rect 331 -2395 332 -2394
rect 352 -2395 353 -2394
rect 380 -2395 381 -2394
rect 520 -2395 521 -2394
rect 527 -2395 528 -2394
rect 1251 -2395 1252 -2394
rect 1339 -2395 1340 -2394
rect 1388 -2395 1389 -2394
rect 1598 -2395 1599 -2394
rect 1710 -2395 1711 -2394
rect 345 -2397 346 -2396
rect 352 -2397 353 -2396
rect 380 -2397 381 -2396
rect 436 -2397 437 -2396
rect 499 -2397 500 -2396
rect 702 -2397 703 -2396
rect 758 -2397 759 -2396
rect 1059 -2397 1060 -2396
rect 1115 -2397 1116 -2396
rect 1192 -2397 1193 -2396
rect 1367 -2397 1368 -2396
rect 1388 -2397 1389 -2396
rect 219 -2399 220 -2398
rect 345 -2399 346 -2398
rect 436 -2399 437 -2398
rect 471 -2399 472 -2398
rect 499 -2399 500 -2398
rect 534 -2399 535 -2398
rect 576 -2399 577 -2398
rect 740 -2399 741 -2398
rect 814 -2399 815 -2398
rect 1059 -2399 1060 -2398
rect 1129 -2399 1130 -2398
rect 1402 -2399 1403 -2398
rect 149 -2401 150 -2400
rect 219 -2401 220 -2400
rect 233 -2401 234 -2400
rect 534 -2401 535 -2400
rect 590 -2401 591 -2400
rect 611 -2401 612 -2400
rect 621 -2401 622 -2400
rect 2130 -2401 2131 -2400
rect 149 -2403 150 -2402
rect 163 -2403 164 -2402
rect 233 -2403 234 -2402
rect 450 -2403 451 -2402
rect 597 -2403 598 -2402
rect 1031 -2403 1032 -2402
rect 1171 -2403 1172 -2402
rect 1465 -2403 1466 -2402
rect 359 -2405 360 -2404
rect 450 -2405 451 -2404
rect 611 -2405 612 -2404
rect 632 -2405 633 -2404
rect 646 -2405 647 -2404
rect 737 -2405 738 -2404
rect 814 -2405 815 -2404
rect 870 -2405 871 -2404
rect 884 -2405 885 -2404
rect 1374 -2405 1375 -2404
rect 198 -2407 199 -2406
rect 359 -2407 360 -2406
rect 443 -2407 444 -2406
rect 471 -2407 472 -2406
rect 478 -2407 479 -2406
rect 870 -2407 871 -2406
rect 919 -2407 920 -2406
rect 2249 -2407 2250 -2406
rect 184 -2409 185 -2408
rect 198 -2409 199 -2408
rect 443 -2409 444 -2408
rect 604 -2409 605 -2408
rect 628 -2409 629 -2408
rect 800 -2409 801 -2408
rect 828 -2409 829 -2408
rect 877 -2409 878 -2408
rect 922 -2409 923 -2408
rect 2312 -2409 2313 -2408
rect 135 -2411 136 -2410
rect 604 -2411 605 -2410
rect 632 -2411 633 -2410
rect 709 -2411 710 -2410
rect 737 -2411 738 -2410
rect 1514 -2411 1515 -2410
rect 135 -2413 136 -2412
rect 415 -2413 416 -2412
rect 660 -2413 661 -2412
rect 989 -2413 990 -2412
rect 1013 -2413 1014 -2412
rect 1402 -2413 1403 -2412
rect 184 -2415 185 -2414
rect 639 -2415 640 -2414
rect 670 -2415 671 -2414
rect 2270 -2415 2271 -2414
rect 268 -2417 269 -2416
rect 670 -2417 671 -2416
rect 800 -2417 801 -2416
rect 807 -2417 808 -2416
rect 828 -2417 829 -2416
rect 898 -2417 899 -2416
rect 922 -2417 923 -2416
rect 1724 -2417 1725 -2416
rect 2270 -2417 2271 -2416
rect 2298 -2417 2299 -2416
rect 366 -2419 367 -2418
rect 709 -2419 710 -2418
rect 835 -2419 836 -2418
rect 1003 -2419 1004 -2418
rect 1017 -2419 1018 -2418
rect 1157 -2419 1158 -2418
rect 1171 -2419 1172 -2418
rect 1913 -2419 1914 -2418
rect 121 -2421 122 -2420
rect 1003 -2421 1004 -2420
rect 1031 -2421 1032 -2420
rect 1731 -2421 1732 -2420
rect 1808 -2421 1809 -2420
rect 1913 -2421 1914 -2420
rect 121 -2423 122 -2422
rect 667 -2423 668 -2422
rect 863 -2423 864 -2422
rect 947 -2423 948 -2422
rect 957 -2423 958 -2422
rect 1157 -2423 1158 -2422
rect 1174 -2423 1175 -2422
rect 1297 -2423 1298 -2422
rect 1332 -2423 1333 -2422
rect 2298 -2423 2299 -2422
rect 107 -2425 108 -2424
rect 667 -2425 668 -2424
rect 898 -2425 899 -2424
rect 968 -2425 969 -2424
rect 975 -2425 976 -2424
rect 1549 -2425 1550 -2424
rect 1633 -2425 1634 -2424
rect 1808 -2425 1809 -2424
rect 107 -2427 108 -2426
rect 128 -2427 129 -2426
rect 156 -2427 157 -2426
rect 366 -2427 367 -2426
rect 415 -2427 416 -2426
rect 513 -2427 514 -2426
rect 555 -2427 556 -2426
rect 807 -2427 808 -2426
rect 933 -2427 934 -2426
rect 2158 -2427 2159 -2426
rect 79 -2429 80 -2428
rect 555 -2429 556 -2428
rect 639 -2429 640 -2428
rect 744 -2429 745 -2428
rect 936 -2429 937 -2428
rect 1626 -2429 1627 -2428
rect 1724 -2429 1725 -2428
rect 1937 -2429 1938 -2428
rect 2 -2431 3 -2430
rect 79 -2431 80 -2430
rect 86 -2431 87 -2430
rect 933 -2431 934 -2430
rect 947 -2431 948 -2430
rect 1066 -2431 1067 -2430
rect 1139 -2431 1140 -2430
rect 2249 -2431 2250 -2430
rect 2 -2433 3 -2432
rect 72 -2433 73 -2432
rect 86 -2433 87 -2432
rect 1500 -2433 1501 -2432
rect 1507 -2433 1508 -2432
rect 1633 -2433 1634 -2432
rect 1731 -2433 1732 -2432
rect 1864 -2433 1865 -2432
rect 128 -2435 129 -2434
rect 548 -2435 549 -2434
rect 695 -2435 696 -2434
rect 744 -2435 745 -2434
rect 961 -2435 962 -2434
rect 1122 -2435 1123 -2434
rect 1178 -2435 1179 -2434
rect 1255 -2435 1256 -2434
rect 1346 -2435 1347 -2434
rect 1864 -2435 1865 -2434
rect 96 -2437 97 -2436
rect 1178 -2437 1179 -2436
rect 1192 -2437 1193 -2436
rect 1325 -2437 1326 -2436
rect 1346 -2437 1347 -2436
rect 1423 -2437 1424 -2436
rect 1500 -2437 1501 -2436
rect 1584 -2437 1585 -2436
rect 1605 -2437 1606 -2436
rect 1626 -2437 1627 -2436
rect 58 -2439 59 -2438
rect 96 -2439 97 -2438
rect 156 -2439 157 -2438
rect 212 -2439 213 -2438
rect 513 -2439 514 -2438
rect 562 -2439 563 -2438
rect 688 -2439 689 -2438
rect 695 -2439 696 -2438
rect 968 -2439 969 -2438
rect 1010 -2439 1011 -2438
rect 1066 -2439 1067 -2438
rect 1143 -2439 1144 -2438
rect 1213 -2439 1214 -2438
rect 1605 -2439 1606 -2438
rect 58 -2441 59 -2440
rect 996 -2441 997 -2440
rect 1010 -2441 1011 -2440
rect 1101 -2441 1102 -2440
rect 1122 -2441 1123 -2440
rect 1206 -2441 1207 -2440
rect 1325 -2441 1326 -2440
rect 1496 -2441 1497 -2440
rect 1507 -2441 1508 -2440
rect 1556 -2441 1557 -2440
rect 1584 -2441 1585 -2440
rect 1654 -2441 1655 -2440
rect 142 -2443 143 -2442
rect 562 -2443 563 -2442
rect 793 -2443 794 -2442
rect 1101 -2443 1102 -2442
rect 1143 -2443 1144 -2442
rect 1521 -2443 1522 -2442
rect 1556 -2443 1557 -2442
rect 1619 -2443 1620 -2442
rect 93 -2445 94 -2444
rect 142 -2445 143 -2444
rect 205 -2445 206 -2444
rect 688 -2445 689 -2444
rect 975 -2445 976 -2444
rect 2018 -2445 2019 -2444
rect 93 -2447 94 -2446
rect 1822 -2447 1823 -2446
rect 205 -2449 206 -2448
rect 674 -2449 675 -2448
rect 996 -2449 997 -2448
rect 1045 -2449 1046 -2448
rect 1206 -2449 1207 -2448
rect 1234 -2449 1235 -2448
rect 1353 -2449 1354 -2448
rect 1423 -2449 1424 -2448
rect 1458 -2449 1459 -2448
rect 1619 -2449 1620 -2448
rect 212 -2451 213 -2450
rect 289 -2451 290 -2450
rect 548 -2451 549 -2450
rect 1804 -2451 1805 -2450
rect 289 -2453 290 -2452
rect 338 -2453 339 -2452
rect 674 -2453 675 -2452
rect 992 -2453 993 -2452
rect 1045 -2453 1046 -2452
rect 1094 -2453 1095 -2452
rect 1234 -2453 1235 -2452
rect 2336 -2453 2337 -2452
rect 338 -2455 339 -2454
rect 541 -2455 542 -2454
rect 926 -2455 927 -2454
rect 1094 -2455 1095 -2454
rect 1353 -2455 1354 -2454
rect 2144 -2455 2145 -2454
rect 541 -2457 542 -2456
rect 849 -2457 850 -2456
rect 992 -2457 993 -2456
rect 2046 -2457 2047 -2456
rect 772 -2459 773 -2458
rect 926 -2459 927 -2458
rect 1199 -2459 1200 -2458
rect 2144 -2459 2145 -2458
rect 23 -2461 24 -2460
rect 772 -2461 773 -2460
rect 849 -2461 850 -2460
rect 1290 -2461 1291 -2460
rect 1367 -2461 1368 -2460
rect 1430 -2461 1431 -2460
rect 1458 -2461 1459 -2460
rect 1577 -2461 1578 -2460
rect 1199 -2463 1200 -2462
rect 1283 -2463 1284 -2462
rect 1430 -2463 1431 -2462
rect 1640 -2463 1641 -2462
rect 1283 -2465 1284 -2464
rect 1416 -2465 1417 -2464
rect 1521 -2465 1522 -2464
rect 1661 -2465 1662 -2464
rect 373 -2467 374 -2466
rect 1661 -2467 1662 -2466
rect 373 -2469 374 -2468
rect 583 -2469 584 -2468
rect 1416 -2469 1417 -2468
rect 1472 -2469 1473 -2468
rect 1563 -2469 1564 -2468
rect 1654 -2469 1655 -2468
rect 583 -2471 584 -2470
rect 653 -2471 654 -2470
rect 1472 -2471 1473 -2470
rect 1601 -2471 1602 -2470
rect 1640 -2471 1641 -2470
rect 1815 -2471 1816 -2470
rect 653 -2473 654 -2472
rect 751 -2473 752 -2472
rect 1563 -2473 1564 -2472
rect 1689 -2473 1690 -2472
rect 1815 -2473 1816 -2472
rect 1871 -2473 1872 -2472
rect 751 -2475 752 -2474
rect 1073 -2475 1074 -2474
rect 1689 -2475 1690 -2474
rect 1759 -2475 1760 -2474
rect 1871 -2475 1872 -2474
rect 1920 -2475 1921 -2474
rect 1073 -2477 1074 -2476
rect 1955 -2477 1956 -2476
rect 1759 -2479 1760 -2478
rect 1794 -2479 1795 -2478
rect 1920 -2479 1921 -2478
rect 1962 -2479 1963 -2478
rect 1675 -2481 1676 -2480
rect 1794 -2481 1795 -2480
rect 1955 -2481 1956 -2480
rect 2004 -2481 2005 -2480
rect 1962 -2483 1963 -2482
rect 2025 -2483 2026 -2482
rect 1083 -2485 1084 -2484
rect 2025 -2485 2026 -2484
rect 2004 -2487 2005 -2486
rect 2032 -2487 2033 -2486
rect 2032 -2489 2033 -2488
rect 2081 -2489 2082 -2488
rect 1220 -2491 1221 -2490
rect 2081 -2491 2082 -2490
rect 1220 -2493 1221 -2492
rect 1241 -2493 1242 -2492
rect 1241 -2495 1242 -2494
rect 1269 -2495 1270 -2494
rect 1269 -2497 1270 -2496
rect 1570 -2497 1571 -2496
rect 5 -2508 6 -2507
rect 415 -2508 416 -2507
rect 464 -2508 465 -2507
rect 989 -2508 990 -2507
rect 992 -2508 993 -2507
rect 1073 -2508 1074 -2507
rect 1080 -2508 1081 -2507
rect 1794 -2508 1795 -2507
rect 1801 -2508 1802 -2507
rect 1934 -2508 1935 -2507
rect 2088 -2508 2089 -2507
rect 2091 -2508 2092 -2507
rect 9 -2510 10 -2509
rect 1409 -2510 1410 -2509
rect 1510 -2510 1511 -2509
rect 2053 -2510 2054 -2509
rect 2088 -2510 2089 -2509
rect 2158 -2510 2159 -2509
rect 9 -2512 10 -2511
rect 51 -2512 52 -2511
rect 54 -2512 55 -2511
rect 765 -2512 766 -2511
rect 775 -2512 776 -2511
rect 877 -2512 878 -2511
rect 926 -2512 927 -2511
rect 1083 -2512 1084 -2511
rect 1188 -2512 1189 -2511
rect 1696 -2512 1697 -2511
rect 1794 -2512 1795 -2511
rect 1885 -2512 1886 -2511
rect 1934 -2512 1935 -2511
rect 2025 -2512 2026 -2511
rect 2053 -2512 2054 -2511
rect 2130 -2512 2131 -2511
rect 16 -2514 17 -2513
rect 37 -2514 38 -2513
rect 40 -2514 41 -2513
rect 1248 -2514 1249 -2513
rect 1290 -2514 1291 -2513
rect 1808 -2514 1809 -2513
rect 1885 -2514 1886 -2513
rect 1997 -2514 1998 -2513
rect 2025 -2514 2026 -2513
rect 2102 -2514 2103 -2513
rect 2130 -2514 2131 -2513
rect 2193 -2514 2194 -2513
rect 33 -2516 34 -2515
rect 933 -2516 934 -2515
rect 950 -2516 951 -2515
rect 1290 -2516 1291 -2515
rect 1335 -2516 1336 -2515
rect 2109 -2516 2110 -2515
rect 37 -2518 38 -2517
rect 51 -2518 52 -2517
rect 58 -2518 59 -2517
rect 1465 -2518 1466 -2517
rect 1580 -2518 1581 -2517
rect 1647 -2518 1648 -2517
rect 1678 -2518 1679 -2517
rect 1969 -2518 1970 -2517
rect 1997 -2518 1998 -2517
rect 2060 -2518 2061 -2517
rect 2102 -2518 2103 -2517
rect 2242 -2518 2243 -2517
rect 44 -2520 45 -2519
rect 75 -2520 76 -2519
rect 93 -2520 94 -2519
rect 1150 -2520 1151 -2519
rect 1195 -2520 1196 -2519
rect 1906 -2520 1907 -2519
rect 1969 -2520 1970 -2519
rect 2032 -2520 2033 -2519
rect 2109 -2520 2110 -2519
rect 2172 -2520 2173 -2519
rect 2242 -2520 2243 -2519
rect 2291 -2520 2292 -2519
rect 44 -2522 45 -2521
rect 527 -2522 528 -2521
rect 541 -2522 542 -2521
rect 978 -2522 979 -2521
rect 989 -2522 990 -2521
rect 1174 -2522 1175 -2521
rect 1199 -2522 1200 -2521
rect 1332 -2522 1333 -2521
rect 1356 -2522 1357 -2521
rect 1696 -2522 1697 -2521
rect 1804 -2522 1805 -2521
rect 2186 -2522 2187 -2521
rect 58 -2524 59 -2523
rect 61 -2524 62 -2523
rect 72 -2524 73 -2523
rect 1237 -2524 1238 -2523
rect 1332 -2524 1333 -2523
rect 1416 -2524 1417 -2523
rect 1458 -2524 1459 -2523
rect 2032 -2524 2033 -2523
rect 2172 -2524 2173 -2523
rect 2235 -2524 2236 -2523
rect 72 -2526 73 -2525
rect 366 -2526 367 -2525
rect 373 -2526 374 -2525
rect 789 -2526 790 -2525
rect 817 -2526 818 -2525
rect 2060 -2526 2061 -2525
rect 2186 -2526 2187 -2525
rect 2256 -2526 2257 -2525
rect 93 -2528 94 -2527
rect 114 -2528 115 -2527
rect 128 -2528 129 -2527
rect 810 -2528 811 -2527
rect 859 -2528 860 -2527
rect 1675 -2528 1676 -2527
rect 1808 -2528 1809 -2527
rect 1871 -2528 1872 -2527
rect 2235 -2528 2236 -2527
rect 2284 -2528 2285 -2527
rect 107 -2530 108 -2529
rect 261 -2530 262 -2529
rect 268 -2530 269 -2529
rect 870 -2530 871 -2529
rect 877 -2530 878 -2529
rect 1311 -2530 1312 -2529
rect 1360 -2530 1361 -2529
rect 2116 -2530 2117 -2529
rect 110 -2532 111 -2531
rect 1360 -2532 1361 -2531
rect 1374 -2532 1375 -2531
rect 1941 -2532 1942 -2531
rect 2116 -2532 2117 -2531
rect 2123 -2532 2124 -2531
rect 131 -2534 132 -2533
rect 968 -2534 969 -2533
rect 1006 -2534 1007 -2533
rect 1031 -2534 1032 -2533
rect 1038 -2534 1039 -2533
rect 1150 -2534 1151 -2533
rect 1216 -2534 1217 -2533
rect 2270 -2534 2271 -2533
rect 19 -2536 20 -2535
rect 1031 -2536 1032 -2535
rect 1038 -2536 1039 -2535
rect 1157 -2536 1158 -2535
rect 1311 -2536 1312 -2535
rect 1843 -2536 1844 -2535
rect 1871 -2536 1872 -2535
rect 1927 -2536 1928 -2535
rect 1941 -2536 1942 -2535
rect 2165 -2536 2166 -2535
rect 2270 -2536 2271 -2535
rect 2312 -2536 2313 -2535
rect 149 -2538 150 -2537
rect 268 -2538 269 -2537
rect 275 -2538 276 -2537
rect 793 -2538 794 -2537
rect 898 -2538 899 -2537
rect 933 -2538 934 -2537
rect 940 -2538 941 -2537
rect 1199 -2538 1200 -2537
rect 1377 -2538 1378 -2537
rect 1654 -2538 1655 -2537
rect 1843 -2538 1844 -2537
rect 1899 -2538 1900 -2537
rect 2123 -2538 2124 -2537
rect 2179 -2538 2180 -2537
rect 103 -2540 104 -2539
rect 898 -2540 899 -2539
rect 919 -2540 920 -2539
rect 968 -2540 969 -2539
rect 1010 -2540 1011 -2539
rect 1122 -2540 1123 -2539
rect 1402 -2540 1403 -2539
rect 1405 -2540 1406 -2539
rect 1416 -2540 1417 -2539
rect 1437 -2540 1438 -2539
rect 1458 -2540 1459 -2539
rect 1514 -2540 1515 -2539
rect 1580 -2540 1581 -2539
rect 2004 -2540 2005 -2539
rect 2165 -2540 2166 -2539
rect 2228 -2540 2229 -2539
rect 128 -2542 129 -2541
rect 940 -2542 941 -2541
rect 1013 -2542 1014 -2541
rect 1374 -2542 1375 -2541
rect 1402 -2542 1403 -2541
rect 1444 -2542 1445 -2541
rect 1465 -2542 1466 -2541
rect 1542 -2542 1543 -2541
rect 1601 -2542 1602 -2541
rect 2095 -2542 2096 -2541
rect 2179 -2542 2180 -2541
rect 2249 -2542 2250 -2541
rect 149 -2544 150 -2543
rect 429 -2544 430 -2543
rect 478 -2544 479 -2543
rect 1661 -2544 1662 -2543
rect 1766 -2544 1767 -2543
rect 2228 -2544 2229 -2543
rect 163 -2546 164 -2545
rect 177 -2546 178 -2545
rect 191 -2546 192 -2545
rect 261 -2546 262 -2545
rect 303 -2546 304 -2545
rect 411 -2546 412 -2545
rect 429 -2546 430 -2545
rect 1440 -2546 1441 -2545
rect 1444 -2546 1445 -2545
rect 1619 -2546 1620 -2545
rect 1647 -2546 1648 -2545
rect 1710 -2546 1711 -2545
rect 1899 -2546 1900 -2545
rect 1962 -2546 1963 -2545
rect 163 -2548 164 -2547
rect 1353 -2548 1354 -2547
rect 1437 -2548 1438 -2547
rect 1703 -2548 1704 -2547
rect 1710 -2548 1711 -2547
rect 1920 -2548 1921 -2547
rect 96 -2550 97 -2549
rect 1353 -2550 1354 -2549
rect 1500 -2550 1501 -2549
rect 1514 -2550 1515 -2549
rect 1542 -2550 1543 -2549
rect 1563 -2550 1564 -2549
rect 1612 -2550 1613 -2549
rect 1927 -2550 1928 -2549
rect 177 -2552 178 -2551
rect 583 -2552 584 -2551
rect 604 -2552 605 -2551
rect 891 -2552 892 -2551
rect 894 -2552 895 -2551
rect 1766 -2552 1767 -2551
rect 1920 -2552 1921 -2551
rect 2011 -2552 2012 -2551
rect 191 -2554 192 -2553
rect 1577 -2554 1578 -2553
rect 1619 -2554 1620 -2553
rect 1976 -2554 1977 -2553
rect 201 -2556 202 -2555
rect 607 -2556 608 -2555
rect 632 -2556 633 -2555
rect 1213 -2556 1214 -2555
rect 1272 -2556 1273 -2555
rect 1703 -2556 1704 -2555
rect 1948 -2556 1949 -2555
rect 2011 -2556 2012 -2555
rect 205 -2558 206 -2557
rect 275 -2558 276 -2557
rect 310 -2558 311 -2557
rect 1269 -2558 1270 -2557
rect 1314 -2558 1315 -2557
rect 2095 -2558 2096 -2557
rect 198 -2560 199 -2559
rect 205 -2560 206 -2559
rect 240 -2560 241 -2559
rect 541 -2560 542 -2559
rect 555 -2560 556 -2559
rect 740 -2560 741 -2559
rect 751 -2560 752 -2559
rect 772 -2560 773 -2559
rect 926 -2560 927 -2559
rect 1297 -2560 1298 -2559
rect 1451 -2560 1452 -2559
rect 1612 -2560 1613 -2559
rect 1654 -2560 1655 -2559
rect 1755 -2560 1756 -2559
rect 1948 -2560 1949 -2559
rect 2039 -2560 2040 -2559
rect 198 -2562 199 -2561
rect 611 -2562 612 -2561
rect 709 -2562 710 -2561
rect 1052 -2562 1053 -2561
rect 1066 -2562 1067 -2561
rect 1409 -2562 1410 -2561
rect 1451 -2562 1452 -2561
rect 1570 -2562 1571 -2561
rect 1661 -2562 1662 -2561
rect 1738 -2562 1739 -2561
rect 1976 -2562 1977 -2561
rect 2046 -2562 2047 -2561
rect 240 -2564 241 -2563
rect 415 -2564 416 -2563
rect 457 -2564 458 -2563
rect 611 -2564 612 -2563
rect 709 -2564 710 -2563
rect 730 -2564 731 -2563
rect 737 -2564 738 -2563
rect 2004 -2564 2005 -2563
rect 2046 -2564 2047 -2563
rect 2207 -2564 2208 -2563
rect 254 -2566 255 -2565
rect 303 -2566 304 -2565
rect 310 -2566 311 -2565
rect 422 -2566 423 -2565
rect 457 -2566 458 -2565
rect 558 -2566 559 -2565
rect 562 -2566 563 -2565
rect 765 -2566 766 -2565
rect 873 -2566 874 -2565
rect 2039 -2566 2040 -2565
rect 2091 -2566 2092 -2565
rect 2158 -2566 2159 -2565
rect 135 -2568 136 -2567
rect 254 -2568 255 -2567
rect 352 -2568 353 -2567
rect 1010 -2568 1011 -2567
rect 1017 -2568 1018 -2567
rect 2193 -2568 2194 -2567
rect 135 -2570 136 -2569
rect 247 -2570 248 -2569
rect 352 -2570 353 -2569
rect 450 -2570 451 -2569
rect 492 -2570 493 -2569
rect 1157 -2570 1158 -2569
rect 1185 -2570 1186 -2569
rect 1962 -2570 1963 -2569
rect 184 -2572 185 -2571
rect 492 -2572 493 -2571
rect 562 -2572 563 -2571
rect 863 -2572 864 -2571
rect 1017 -2572 1018 -2571
rect 1108 -2572 1109 -2571
rect 1122 -2572 1123 -2571
rect 1423 -2572 1424 -2571
rect 1479 -2572 1480 -2571
rect 1563 -2572 1564 -2571
rect 1570 -2572 1571 -2571
rect 1605 -2572 1606 -2571
rect 1738 -2572 1739 -2571
rect 1787 -2572 1788 -2571
rect 142 -2574 143 -2573
rect 863 -2574 864 -2573
rect 1052 -2574 1053 -2573
rect 1115 -2574 1116 -2573
rect 1213 -2574 1214 -2573
rect 1325 -2574 1326 -2573
rect 1423 -2574 1424 -2573
rect 1528 -2574 1529 -2573
rect 1605 -2574 1606 -2573
rect 1682 -2574 1683 -2573
rect 1787 -2574 1788 -2573
rect 1864 -2574 1865 -2573
rect 142 -2576 143 -2575
rect 891 -2576 892 -2575
rect 1066 -2576 1067 -2575
rect 1318 -2576 1319 -2575
rect 1479 -2576 1480 -2575
rect 1486 -2576 1487 -2575
rect 1500 -2576 1501 -2575
rect 1584 -2576 1585 -2575
rect 1682 -2576 1683 -2575
rect 1759 -2576 1760 -2575
rect 1850 -2576 1851 -2575
rect 1864 -2576 1865 -2575
rect 184 -2578 185 -2577
rect 975 -2578 976 -2577
rect 1073 -2578 1074 -2577
rect 1094 -2578 1095 -2577
rect 1269 -2578 1270 -2577
rect 1388 -2578 1389 -2577
rect 1486 -2578 1487 -2577
rect 1549 -2578 1550 -2577
rect 1584 -2578 1585 -2577
rect 1626 -2578 1627 -2577
rect 1731 -2578 1732 -2577
rect 1759 -2578 1760 -2577
rect 1850 -2578 1851 -2577
rect 1955 -2578 1956 -2577
rect 219 -2580 220 -2579
rect 422 -2580 423 -2579
rect 450 -2580 451 -2579
rect 828 -2580 829 -2579
rect 842 -2580 843 -2579
rect 975 -2580 976 -2579
rect 1080 -2580 1081 -2579
rect 1087 -2580 1088 -2579
rect 1094 -2580 1095 -2579
rect 1143 -2580 1144 -2579
rect 1297 -2580 1298 -2579
rect 1395 -2580 1396 -2579
rect 1528 -2580 1529 -2579
rect 1633 -2580 1634 -2579
rect 1955 -2580 1956 -2579
rect 2018 -2580 2019 -2579
rect 86 -2582 87 -2581
rect 842 -2582 843 -2581
rect 1087 -2582 1088 -2581
rect 1381 -2582 1382 -2581
rect 1388 -2582 1389 -2581
rect 1493 -2582 1494 -2581
rect 1549 -2582 1550 -2581
rect 1745 -2582 1746 -2581
rect 1990 -2582 1991 -2581
rect 2018 -2582 2019 -2581
rect 86 -2584 87 -2583
rect 922 -2584 923 -2583
rect 1143 -2584 1144 -2583
rect 1220 -2584 1221 -2583
rect 1234 -2584 1235 -2583
rect 1381 -2584 1382 -2583
rect 1395 -2584 1396 -2583
rect 1829 -2584 1830 -2583
rect 1878 -2584 1879 -2583
rect 1990 -2584 1991 -2583
rect 26 -2586 27 -2585
rect 1878 -2586 1879 -2585
rect 219 -2588 220 -2587
rect 317 -2588 318 -2587
rect 359 -2588 360 -2587
rect 1363 -2588 1364 -2587
rect 1430 -2588 1431 -2587
rect 1493 -2588 1494 -2587
rect 1591 -2588 1592 -2587
rect 1731 -2588 1732 -2587
rect 1745 -2588 1746 -2587
rect 1815 -2588 1816 -2587
rect 1829 -2588 1830 -2587
rect 1836 -2588 1837 -2587
rect 212 -2590 213 -2589
rect 317 -2590 318 -2589
rect 331 -2590 332 -2589
rect 359 -2590 360 -2589
rect 366 -2590 367 -2589
rect 506 -2590 507 -2589
rect 569 -2590 570 -2589
rect 632 -2590 633 -2589
rect 646 -2590 647 -2589
rect 1185 -2590 1186 -2589
rect 1220 -2590 1221 -2589
rect 1339 -2590 1340 -2589
rect 1430 -2590 1431 -2589
rect 1598 -2590 1599 -2589
rect 1626 -2590 1627 -2589
rect 1689 -2590 1690 -2589
rect 1815 -2590 1816 -2589
rect 1857 -2590 1858 -2589
rect 212 -2592 213 -2591
rect 597 -2592 598 -2591
rect 646 -2592 647 -2591
rect 688 -2592 689 -2591
rect 716 -2592 717 -2591
rect 793 -2592 794 -2591
rect 828 -2592 829 -2591
rect 1304 -2592 1305 -2591
rect 1318 -2592 1319 -2591
rect 1535 -2592 1536 -2591
rect 1591 -2592 1592 -2591
rect 1773 -2592 1774 -2591
rect 1836 -2592 1837 -2591
rect 1892 -2592 1893 -2591
rect 68 -2594 69 -2593
rect 688 -2594 689 -2593
rect 716 -2594 717 -2593
rect 1206 -2594 1207 -2593
rect 1234 -2594 1235 -2593
rect 1262 -2594 1263 -2593
rect 1339 -2594 1340 -2593
rect 1398 -2594 1399 -2593
rect 1472 -2594 1473 -2593
rect 1535 -2594 1536 -2593
rect 1598 -2594 1599 -2593
rect 1668 -2594 1669 -2593
rect 1773 -2594 1774 -2593
rect 1822 -2594 1823 -2593
rect 1857 -2594 1858 -2593
rect 2074 -2594 2075 -2593
rect 226 -2596 227 -2595
rect 247 -2596 248 -2595
rect 282 -2596 283 -2595
rect 1115 -2596 1116 -2595
rect 1171 -2596 1172 -2595
rect 1892 -2596 1893 -2595
rect 2074 -2596 2075 -2595
rect 2144 -2596 2145 -2595
rect 170 -2598 171 -2597
rect 226 -2598 227 -2597
rect 282 -2598 283 -2597
rect 670 -2598 671 -2597
rect 723 -2598 724 -2597
rect 737 -2598 738 -2597
rect 751 -2598 752 -2597
rect 1125 -2598 1126 -2597
rect 1171 -2598 1172 -2597
rect 1255 -2598 1256 -2597
rect 1262 -2598 1263 -2597
rect 1346 -2598 1347 -2597
rect 1412 -2598 1413 -2597
rect 1472 -2598 1473 -2597
rect 1633 -2598 1634 -2597
rect 2280 -2598 2281 -2597
rect 166 -2600 167 -2599
rect 170 -2600 171 -2599
rect 331 -2600 332 -2599
rect 345 -2600 346 -2599
rect 373 -2600 374 -2599
rect 394 -2600 395 -2599
rect 401 -2600 402 -2599
rect 856 -2600 857 -2599
rect 954 -2600 955 -2599
rect 1346 -2600 1347 -2599
rect 1640 -2600 1641 -2599
rect 1689 -2600 1690 -2599
rect 1822 -2600 1823 -2599
rect 1913 -2600 1914 -2599
rect 2144 -2600 2145 -2599
rect 2214 -2600 2215 -2599
rect 30 -2602 31 -2601
rect 345 -2602 346 -2601
rect 380 -2602 381 -2601
rect 527 -2602 528 -2601
rect 569 -2602 570 -2601
rect 814 -2602 815 -2601
rect 824 -2602 825 -2601
rect 1304 -2602 1305 -2601
rect 1640 -2602 1641 -2601
rect 1724 -2602 1725 -2601
rect 1913 -2602 1914 -2601
rect 1983 -2602 1984 -2601
rect 2214 -2602 2215 -2601
rect 2263 -2602 2264 -2601
rect 30 -2604 31 -2603
rect 485 -2604 486 -2603
rect 506 -2604 507 -2603
rect 849 -2604 850 -2603
rect 1178 -2604 1179 -2603
rect 1983 -2604 1984 -2603
rect 2263 -2604 2264 -2603
rect 2305 -2604 2306 -2603
rect 79 -2606 80 -2605
rect 856 -2606 857 -2605
rect 1003 -2606 1004 -2605
rect 1178 -2606 1179 -2605
rect 1206 -2606 1207 -2605
rect 1283 -2606 1284 -2605
rect 1447 -2606 1448 -2605
rect 1724 -2606 1725 -2605
rect 79 -2608 80 -2607
rect 548 -2608 549 -2607
rect 583 -2608 584 -2607
rect 800 -2608 801 -2607
rect 807 -2608 808 -2607
rect 1003 -2608 1004 -2607
rect 1255 -2608 1256 -2607
rect 1577 -2608 1578 -2607
rect 1668 -2608 1669 -2607
rect 1752 -2608 1753 -2607
rect 156 -2610 157 -2609
rect 401 -2610 402 -2609
rect 408 -2610 409 -2609
rect 464 -2610 465 -2609
rect 485 -2610 486 -2609
rect 639 -2610 640 -2609
rect 726 -2610 727 -2609
rect 2081 -2610 2082 -2609
rect 156 -2612 157 -2611
rect 555 -2612 556 -2611
rect 597 -2612 598 -2611
rect 957 -2612 958 -2611
rect 1752 -2612 1753 -2611
rect 2298 -2612 2299 -2611
rect 289 -2614 290 -2613
rect 408 -2614 409 -2613
rect 520 -2614 521 -2613
rect 954 -2614 955 -2613
rect 2081 -2614 2082 -2613
rect 2151 -2614 2152 -2613
rect 65 -2616 66 -2615
rect 289 -2616 290 -2615
rect 380 -2616 381 -2615
rect 660 -2616 661 -2615
rect 730 -2616 731 -2615
rect 982 -2616 983 -2615
rect 2151 -2616 2152 -2615
rect 2221 -2616 2222 -2615
rect 65 -2618 66 -2617
rect 2067 -2618 2068 -2617
rect 387 -2620 388 -2619
rect 478 -2620 479 -2619
rect 513 -2620 514 -2619
rect 660 -2620 661 -2619
rect 758 -2620 759 -2619
rect 1108 -2620 1109 -2619
rect 2067 -2620 2068 -2619
rect 2137 -2620 2138 -2619
rect 338 -2622 339 -2621
rect 387 -2622 388 -2621
rect 394 -2622 395 -2621
rect 1055 -2622 1056 -2621
rect 2137 -2622 2138 -2621
rect 2200 -2622 2201 -2621
rect 338 -2624 339 -2623
rect 499 -2624 500 -2623
rect 513 -2624 514 -2623
rect 695 -2624 696 -2623
rect 786 -2624 787 -2623
rect 1283 -2624 1284 -2623
rect 443 -2626 444 -2625
rect 499 -2626 500 -2625
rect 520 -2626 521 -2625
rect 576 -2626 577 -2625
rect 590 -2626 591 -2625
rect 758 -2626 759 -2625
rect 800 -2626 801 -2625
rect 1556 -2626 1557 -2625
rect 233 -2628 234 -2627
rect 443 -2628 444 -2627
rect 534 -2628 535 -2627
rect 590 -2628 591 -2627
rect 618 -2628 619 -2627
rect 814 -2628 815 -2627
rect 849 -2628 850 -2627
rect 1101 -2628 1102 -2627
rect 1507 -2628 1508 -2627
rect 1556 -2628 1557 -2627
rect 233 -2630 234 -2629
rect 674 -2630 675 -2629
rect 695 -2630 696 -2629
rect 996 -2630 997 -2629
rect 1101 -2630 1102 -2629
rect 1136 -2630 1137 -2629
rect 1248 -2630 1249 -2629
rect 1507 -2630 1508 -2629
rect 324 -2632 325 -2631
rect 534 -2632 535 -2631
rect 548 -2632 549 -2631
rect 835 -2632 836 -2631
rect 982 -2632 983 -2631
rect 1059 -2632 1060 -2631
rect 1136 -2632 1137 -2631
rect 2221 -2632 2222 -2631
rect 324 -2634 325 -2633
rect 471 -2634 472 -2633
rect 576 -2634 577 -2633
rect 786 -2634 787 -2633
rect 796 -2634 797 -2633
rect 1059 -2634 1060 -2633
rect 23 -2636 24 -2635
rect 471 -2636 472 -2635
rect 618 -2636 619 -2635
rect 884 -2636 885 -2635
rect 996 -2636 997 -2635
rect 1045 -2636 1046 -2635
rect 639 -2638 640 -2637
rect 681 -2638 682 -2637
rect 779 -2638 780 -2637
rect 835 -2638 836 -2637
rect 884 -2638 885 -2637
rect 905 -2638 906 -2637
rect 1045 -2638 1046 -2637
rect 1276 -2638 1277 -2637
rect 121 -2640 122 -2639
rect 779 -2640 780 -2639
rect 1241 -2640 1242 -2639
rect 1276 -2640 1277 -2639
rect 481 -2642 482 -2641
rect 905 -2642 906 -2641
rect 1241 -2642 1242 -2641
rect 1780 -2642 1781 -2641
rect 625 -2644 626 -2643
rect 681 -2644 682 -2643
rect 1013 -2644 1014 -2643
rect 1780 -2644 1781 -2643
rect 625 -2646 626 -2645
rect 912 -2646 913 -2645
rect 667 -2648 668 -2647
rect 2200 -2648 2201 -2647
rect 667 -2650 668 -2649
rect 702 -2650 703 -2649
rect 912 -2650 913 -2649
rect 1129 -2650 1130 -2649
rect 674 -2652 675 -2651
rect 821 -2652 822 -2651
rect 1129 -2652 1130 -2651
rect 1164 -2652 1165 -2651
rect 114 -2654 115 -2653
rect 821 -2654 822 -2653
rect 1164 -2654 1165 -2653
rect 1227 -2654 1228 -2653
rect 702 -2656 703 -2655
rect 744 -2656 745 -2655
rect 1227 -2656 1228 -2655
rect 1367 -2656 1368 -2655
rect 744 -2658 745 -2657
rect 961 -2658 962 -2657
rect 1192 -2658 1193 -2657
rect 1367 -2658 1368 -2657
rect 947 -2660 948 -2659
rect 961 -2660 962 -2659
rect 1192 -2660 1193 -2659
rect 1906 -2660 1907 -2659
rect 296 -2662 297 -2661
rect 947 -2662 948 -2661
rect 296 -2664 297 -2663
rect 436 -2664 437 -2663
rect 436 -2666 437 -2665
rect 653 -2666 654 -2665
rect 100 -2668 101 -2667
rect 653 -2668 654 -2667
rect 100 -2670 101 -2669
rect 121 -2670 122 -2669
rect 2 -2681 3 -2680
rect 68 -2681 69 -2680
rect 103 -2681 104 -2680
rect 338 -2681 339 -2680
rect 432 -2681 433 -2680
rect 464 -2681 465 -2680
rect 506 -2681 507 -2680
rect 733 -2681 734 -2680
rect 758 -2681 759 -2680
rect 838 -2681 839 -2680
rect 915 -2681 916 -2680
rect 2046 -2681 2047 -2680
rect 2224 -2681 2225 -2680
rect 2270 -2681 2271 -2680
rect 16 -2683 17 -2682
rect 250 -2683 251 -2682
rect 338 -2683 339 -2682
rect 345 -2683 346 -2682
rect 506 -2683 507 -2682
rect 779 -2683 780 -2682
rect 786 -2683 787 -2682
rect 1150 -2683 1151 -2682
rect 1185 -2683 1186 -2682
rect 1885 -2683 1886 -2682
rect 1927 -2683 1928 -2682
rect 2259 -2683 2260 -2682
rect 16 -2685 17 -2684
rect 695 -2685 696 -2684
rect 709 -2685 710 -2684
rect 957 -2685 958 -2684
rect 978 -2685 979 -2684
rect 1283 -2685 1284 -2684
rect 1286 -2685 1287 -2684
rect 1458 -2685 1459 -2684
rect 1489 -2685 1490 -2684
rect 1591 -2685 1592 -2684
rect 1619 -2685 1620 -2684
rect 1885 -2685 1886 -2684
rect 23 -2687 24 -2686
rect 135 -2687 136 -2686
rect 156 -2687 157 -2686
rect 1055 -2687 1056 -2686
rect 1062 -2687 1063 -2686
rect 1136 -2687 1137 -2686
rect 1139 -2687 1140 -2686
rect 1479 -2687 1480 -2686
rect 1577 -2687 1578 -2686
rect 2249 -2687 2250 -2686
rect 23 -2689 24 -2688
rect 520 -2689 521 -2688
rect 548 -2689 549 -2688
rect 817 -2689 818 -2688
rect 821 -2689 822 -2688
rect 933 -2689 934 -2688
rect 954 -2689 955 -2688
rect 1143 -2689 1144 -2688
rect 1185 -2689 1186 -2688
rect 1206 -2689 1207 -2688
rect 1234 -2689 1235 -2688
rect 2004 -2689 2005 -2688
rect 26 -2691 27 -2690
rect 842 -2691 843 -2690
rect 919 -2691 920 -2690
rect 1955 -2691 1956 -2690
rect 65 -2693 66 -2692
rect 86 -2693 87 -2692
rect 110 -2693 111 -2692
rect 282 -2693 283 -2692
rect 345 -2693 346 -2692
rect 359 -2693 360 -2692
rect 387 -2693 388 -2692
rect 520 -2693 521 -2692
rect 555 -2693 556 -2692
rect 632 -2693 633 -2692
rect 681 -2693 682 -2692
rect 723 -2693 724 -2692
rect 765 -2693 766 -2692
rect 950 -2693 951 -2692
rect 954 -2693 955 -2692
rect 975 -2693 976 -2692
rect 1013 -2693 1014 -2692
rect 2102 -2693 2103 -2692
rect 65 -2695 66 -2694
rect 996 -2695 997 -2694
rect 1041 -2695 1042 -2694
rect 1871 -2695 1872 -2694
rect 1955 -2695 1956 -2694
rect 1976 -2695 1977 -2694
rect 2102 -2695 2103 -2694
rect 2137 -2695 2138 -2694
rect 82 -2697 83 -2696
rect 632 -2697 633 -2696
rect 681 -2697 682 -2696
rect 716 -2697 717 -2696
rect 765 -2697 766 -2696
rect 1220 -2697 1221 -2696
rect 1234 -2697 1235 -2696
rect 1395 -2697 1396 -2696
rect 1423 -2697 1424 -2696
rect 1458 -2697 1459 -2696
rect 1479 -2697 1480 -2696
rect 1556 -2697 1557 -2696
rect 1584 -2697 1585 -2696
rect 1685 -2697 1686 -2696
rect 1755 -2697 1756 -2696
rect 2158 -2697 2159 -2696
rect 86 -2699 87 -2698
rect 1258 -2699 1259 -2698
rect 1318 -2699 1319 -2698
rect 2270 -2699 2271 -2698
rect 107 -2701 108 -2700
rect 555 -2701 556 -2700
rect 558 -2701 559 -2700
rect 660 -2701 661 -2700
rect 695 -2701 696 -2700
rect 737 -2701 738 -2700
rect 772 -2701 773 -2700
rect 891 -2701 892 -2700
rect 919 -2701 920 -2700
rect 961 -2701 962 -2700
rect 975 -2701 976 -2700
rect 1927 -2701 1928 -2700
rect 1976 -2701 1977 -2700
rect 2018 -2701 2019 -2700
rect 2130 -2701 2131 -2700
rect 2137 -2701 2138 -2700
rect 2158 -2701 2159 -2700
rect 2172 -2701 2173 -2700
rect 121 -2703 122 -2702
rect 128 -2703 129 -2702
rect 163 -2703 164 -2702
rect 548 -2703 549 -2702
rect 562 -2703 563 -2702
rect 1038 -2703 1039 -2702
rect 1066 -2703 1067 -2702
rect 1143 -2703 1144 -2702
rect 1195 -2703 1196 -2702
rect 1444 -2703 1445 -2702
rect 1556 -2703 1557 -2702
rect 1787 -2703 1788 -2702
rect 1871 -2703 1872 -2702
rect 1906 -2703 1907 -2702
rect 2011 -2703 2012 -2702
rect 2018 -2703 2019 -2702
rect 2130 -2703 2131 -2702
rect 2144 -2703 2145 -2702
rect 51 -2705 52 -2704
rect 1444 -2705 1445 -2704
rect 1584 -2705 1585 -2704
rect 1696 -2705 1697 -2704
rect 1759 -2705 1760 -2704
rect 2004 -2705 2005 -2704
rect 2144 -2705 2145 -2704
rect 2151 -2705 2152 -2704
rect 51 -2707 52 -2706
rect 982 -2707 983 -2706
rect 996 -2707 997 -2706
rect 1213 -2707 1214 -2706
rect 1220 -2707 1221 -2706
rect 1262 -2707 1263 -2706
rect 1360 -2707 1361 -2706
rect 1591 -2707 1592 -2706
rect 1619 -2707 1620 -2706
rect 1633 -2707 1634 -2706
rect 1647 -2707 1648 -2706
rect 1706 -2707 1707 -2706
rect 1759 -2707 1760 -2706
rect 1766 -2707 1767 -2706
rect 1899 -2707 1900 -2706
rect 1906 -2707 1907 -2706
rect 2151 -2707 2152 -2706
rect 2165 -2707 2166 -2706
rect 121 -2709 122 -2708
rect 667 -2709 668 -2708
rect 730 -2709 731 -2708
rect 1038 -2709 1039 -2708
rect 1066 -2709 1067 -2708
rect 1129 -2709 1130 -2708
rect 1206 -2709 1207 -2708
rect 1227 -2709 1228 -2708
rect 1241 -2709 1242 -2708
rect 1892 -2709 1893 -2708
rect 1899 -2709 1900 -2708
rect 1913 -2709 1914 -2708
rect 2165 -2709 2166 -2708
rect 2179 -2709 2180 -2708
rect 128 -2711 129 -2710
rect 436 -2711 437 -2710
rect 457 -2711 458 -2710
rect 562 -2711 563 -2710
rect 576 -2711 577 -2710
rect 709 -2711 710 -2710
rect 730 -2711 731 -2710
rect 2179 -2711 2180 -2710
rect 93 -2713 94 -2712
rect 436 -2713 437 -2712
rect 513 -2713 514 -2712
rect 737 -2713 738 -2712
rect 772 -2713 773 -2712
rect 1171 -2713 1172 -2712
rect 1213 -2713 1214 -2712
rect 1269 -2713 1270 -2712
rect 1276 -2713 1277 -2712
rect 1360 -2713 1361 -2712
rect 1374 -2713 1375 -2712
rect 1507 -2713 1508 -2712
rect 1598 -2713 1599 -2712
rect 1633 -2713 1634 -2712
rect 1647 -2713 1648 -2712
rect 1654 -2713 1655 -2712
rect 1668 -2713 1669 -2712
rect 1696 -2713 1697 -2712
rect 1766 -2713 1767 -2712
rect 2053 -2713 2054 -2712
rect 93 -2715 94 -2714
rect 114 -2715 115 -2714
rect 163 -2715 164 -2714
rect 352 -2715 353 -2714
rect 366 -2715 367 -2714
rect 660 -2715 661 -2714
rect 663 -2715 664 -2714
rect 1276 -2715 1277 -2714
rect 1388 -2715 1389 -2714
rect 1423 -2715 1424 -2714
rect 1430 -2715 1431 -2714
rect 1983 -2715 1984 -2714
rect 2053 -2715 2054 -2714
rect 2081 -2715 2082 -2714
rect 114 -2717 115 -2716
rect 478 -2717 479 -2716
rect 513 -2717 514 -2716
rect 1031 -2717 1032 -2716
rect 1073 -2717 1074 -2716
rect 1283 -2717 1284 -2716
rect 1395 -2717 1396 -2716
rect 2221 -2717 2222 -2716
rect 184 -2719 185 -2718
rect 1391 -2719 1392 -2718
rect 1398 -2719 1399 -2718
rect 2011 -2719 2012 -2718
rect 2060 -2719 2061 -2718
rect 2081 -2719 2082 -2718
rect 2221 -2719 2222 -2718
rect 2263 -2719 2264 -2718
rect 75 -2721 76 -2720
rect 184 -2721 185 -2720
rect 226 -2721 227 -2720
rect 387 -2721 388 -2720
rect 478 -2721 479 -2720
rect 856 -2721 857 -2720
rect 877 -2721 878 -2720
rect 1129 -2721 1130 -2720
rect 1227 -2721 1228 -2720
rect 1314 -2721 1315 -2720
rect 1433 -2721 1434 -2720
rect 2228 -2721 2229 -2720
rect 44 -2723 45 -2722
rect 856 -2723 857 -2722
rect 877 -2723 878 -2722
rect 1087 -2723 1088 -2722
rect 1097 -2723 1098 -2722
rect 2032 -2723 2033 -2722
rect 2060 -2723 2061 -2722
rect 2088 -2723 2089 -2722
rect 2214 -2723 2215 -2722
rect 2228 -2723 2229 -2722
rect 44 -2725 45 -2724
rect 471 -2725 472 -2724
rect 576 -2725 577 -2724
rect 646 -2725 647 -2724
rect 667 -2725 668 -2724
rect 702 -2725 703 -2724
rect 779 -2725 780 -2724
rect 849 -2725 850 -2724
rect 912 -2725 913 -2724
rect 1171 -2725 1172 -2724
rect 1262 -2725 1263 -2724
rect 1290 -2725 1291 -2724
rect 1437 -2725 1438 -2724
rect 1864 -2725 1865 -2724
rect 1962 -2725 1963 -2724
rect 1983 -2725 1984 -2724
rect 2088 -2725 2089 -2724
rect 2095 -2725 2096 -2724
rect 135 -2727 136 -2726
rect 912 -2727 913 -2726
rect 933 -2727 934 -2726
rect 1003 -2727 1004 -2726
rect 1010 -2727 1011 -2726
rect 1241 -2727 1242 -2726
rect 1244 -2727 1245 -2726
rect 1864 -2727 1865 -2726
rect 2095 -2727 2096 -2726
rect 2109 -2727 2110 -2726
rect 142 -2729 143 -2728
rect 646 -2729 647 -2728
rect 688 -2729 689 -2728
rect 1892 -2729 1893 -2728
rect 142 -2731 143 -2730
rect 170 -2731 171 -2730
rect 226 -2731 227 -2730
rect 331 -2731 332 -2730
rect 352 -2731 353 -2730
rect 541 -2731 542 -2730
rect 604 -2731 605 -2730
rect 1192 -2731 1193 -2730
rect 1269 -2731 1270 -2730
rect 1297 -2731 1298 -2730
rect 1437 -2731 1438 -2730
rect 1486 -2731 1487 -2730
rect 1500 -2731 1501 -2730
rect 1507 -2731 1508 -2730
rect 1528 -2731 1529 -2730
rect 1598 -2731 1599 -2730
rect 1626 -2731 1627 -2730
rect 1654 -2731 1655 -2730
rect 1668 -2731 1669 -2730
rect 1682 -2731 1683 -2730
rect 1780 -2731 1781 -2730
rect 2032 -2731 2033 -2730
rect 79 -2733 80 -2732
rect 604 -2733 605 -2732
rect 625 -2733 626 -2732
rect 758 -2733 759 -2732
rect 786 -2733 787 -2732
rect 2172 -2733 2173 -2732
rect 9 -2735 10 -2734
rect 79 -2735 80 -2734
rect 149 -2735 150 -2734
rect 331 -2735 332 -2734
rect 415 -2735 416 -2734
rect 1010 -2735 1011 -2734
rect 1073 -2735 1074 -2734
rect 1157 -2735 1158 -2734
rect 1192 -2735 1193 -2734
rect 1353 -2735 1354 -2734
rect 1440 -2735 1441 -2734
rect 2214 -2735 2215 -2734
rect 9 -2737 10 -2736
rect 863 -2737 864 -2736
rect 870 -2737 871 -2736
rect 1157 -2737 1158 -2736
rect 1290 -2737 1291 -2736
rect 1332 -2737 1333 -2736
rect 1353 -2737 1354 -2736
rect 1367 -2737 1368 -2736
rect 1472 -2737 1473 -2736
rect 2263 -2737 2264 -2736
rect 30 -2739 31 -2738
rect 415 -2739 416 -2738
rect 471 -2739 472 -2738
rect 492 -2739 493 -2738
rect 527 -2739 528 -2738
rect 863 -2739 864 -2738
rect 870 -2739 871 -2738
rect 1045 -2739 1046 -2738
rect 1087 -2739 1088 -2738
rect 1101 -2739 1102 -2738
rect 1108 -2739 1109 -2738
rect 1150 -2739 1151 -2738
rect 1332 -2739 1333 -2738
rect 2207 -2739 2208 -2738
rect 30 -2741 31 -2740
rect 254 -2741 255 -2740
rect 261 -2741 262 -2740
rect 359 -2741 360 -2740
rect 408 -2741 409 -2740
rect 1108 -2741 1109 -2740
rect 1115 -2741 1116 -2740
rect 1311 -2741 1312 -2740
rect 1314 -2741 1315 -2740
rect 2207 -2741 2208 -2740
rect 54 -2743 55 -2742
rect 1045 -2743 1046 -2742
rect 1101 -2743 1102 -2742
rect 1325 -2743 1326 -2742
rect 1367 -2743 1368 -2742
rect 1402 -2743 1403 -2742
rect 1451 -2743 1452 -2742
rect 1472 -2743 1473 -2742
rect 1521 -2743 1522 -2742
rect 1528 -2743 1529 -2742
rect 1580 -2743 1581 -2742
rect 1962 -2743 1963 -2742
rect 37 -2745 38 -2744
rect 1402 -2745 1403 -2744
rect 1521 -2745 1522 -2744
rect 1549 -2745 1550 -2744
rect 1626 -2745 1627 -2744
rect 1640 -2745 1641 -2744
rect 1850 -2745 1851 -2744
rect 2109 -2745 2110 -2744
rect 37 -2747 38 -2746
rect 450 -2747 451 -2746
rect 492 -2747 493 -2746
rect 726 -2747 727 -2746
rect 793 -2747 794 -2746
rect 842 -2747 843 -2746
rect 849 -2747 850 -2746
rect 1255 -2747 1256 -2746
rect 1549 -2747 1550 -2746
rect 1570 -2747 1571 -2746
rect 1689 -2747 1690 -2746
rect 1850 -2747 1851 -2746
rect 54 -2749 55 -2748
rect 1913 -2749 1914 -2748
rect 131 -2751 132 -2750
rect 149 -2751 150 -2750
rect 156 -2751 157 -2750
rect 1433 -2751 1434 -2750
rect 1570 -2751 1571 -2750
rect 1661 -2751 1662 -2750
rect 1689 -2751 1690 -2750
rect 1717 -2751 1718 -2750
rect 170 -2753 171 -2752
rect 317 -2753 318 -2752
rect 408 -2753 409 -2752
rect 422 -2753 423 -2752
rect 450 -2753 451 -2752
rect 597 -2753 598 -2752
rect 625 -2753 626 -2752
rect 964 -2753 965 -2752
rect 968 -2753 969 -2752
rect 1374 -2753 1375 -2752
rect 1542 -2753 1543 -2752
rect 1717 -2753 1718 -2752
rect 205 -2755 206 -2754
rect 254 -2755 255 -2754
rect 282 -2755 283 -2754
rect 310 -2755 311 -2754
rect 317 -2755 318 -2754
rect 443 -2755 444 -2754
rect 527 -2755 528 -2754
rect 751 -2755 752 -2754
rect 793 -2755 794 -2754
rect 1510 -2755 1511 -2754
rect 1542 -2755 1543 -2754
rect 1563 -2755 1564 -2754
rect 1661 -2755 1662 -2754
rect 1675 -2755 1676 -2754
rect 205 -2757 206 -2756
rect 1752 -2757 1753 -2756
rect 233 -2759 234 -2758
rect 261 -2759 262 -2758
rect 289 -2759 290 -2758
rect 366 -2759 367 -2758
rect 411 -2759 412 -2758
rect 1325 -2759 1326 -2758
rect 1675 -2759 1676 -2758
rect 1731 -2759 1732 -2758
rect 240 -2761 241 -2760
rect 1178 -2761 1179 -2760
rect 1255 -2761 1256 -2760
rect 1514 -2761 1515 -2760
rect 1731 -2761 1732 -2760
rect 1857 -2761 1858 -2760
rect 243 -2763 244 -2762
rect 401 -2763 402 -2762
rect 443 -2763 444 -2762
rect 705 -2763 706 -2762
rect 744 -2763 745 -2762
rect 968 -2763 969 -2762
rect 982 -2763 983 -2762
rect 1017 -2763 1018 -2762
rect 1059 -2763 1060 -2762
rect 1178 -2763 1179 -2762
rect 1514 -2763 1515 -2762
rect 1724 -2763 1725 -2762
rect 1857 -2763 1858 -2762
rect 1878 -2763 1879 -2762
rect 212 -2765 213 -2764
rect 401 -2765 402 -2764
rect 464 -2765 465 -2764
rect 1059 -2765 1060 -2764
rect 1115 -2765 1116 -2764
rect 1164 -2765 1165 -2764
rect 1724 -2765 1725 -2764
rect 1738 -2765 1739 -2764
rect 1878 -2765 1879 -2764
rect 2123 -2765 2124 -2764
rect 212 -2767 213 -2766
rect 303 -2767 304 -2766
rect 310 -2767 311 -2766
rect 590 -2767 591 -2766
rect 597 -2767 598 -2766
rect 1465 -2767 1466 -2766
rect 1738 -2767 1739 -2766
rect 1745 -2767 1746 -2766
rect 177 -2769 178 -2768
rect 590 -2769 591 -2768
rect 621 -2769 622 -2768
rect 751 -2769 752 -2768
rect 789 -2769 790 -2768
rect 2123 -2769 2124 -2768
rect 177 -2771 178 -2770
rect 898 -2771 899 -2770
rect 943 -2771 944 -2770
rect 1787 -2771 1788 -2770
rect 247 -2773 248 -2772
rect 303 -2773 304 -2772
rect 324 -2773 325 -2772
rect 422 -2773 423 -2772
rect 541 -2773 542 -2772
rect 1318 -2773 1319 -2772
rect 1465 -2773 1466 -2772
rect 1493 -2773 1494 -2772
rect 1496 -2773 1497 -2772
rect 1745 -2773 1746 -2772
rect 289 -2775 290 -2774
rect 569 -2775 570 -2774
rect 639 -2775 640 -2774
rect 716 -2775 717 -2774
rect 744 -2775 745 -2774
rect 1577 -2775 1578 -2774
rect 296 -2777 297 -2776
rect 324 -2777 325 -2776
rect 569 -2777 570 -2776
rect 674 -2777 675 -2776
rect 688 -2777 689 -2776
rect 940 -2777 941 -2776
rect 947 -2777 948 -2776
rect 1031 -2777 1032 -2776
rect 1122 -2777 1123 -2776
rect 1297 -2777 1298 -2776
rect 1493 -2777 1494 -2776
rect 1710 -2777 1711 -2776
rect 72 -2779 73 -2778
rect 296 -2779 297 -2778
rect 460 -2779 461 -2778
rect 1122 -2779 1123 -2778
rect 1125 -2779 1126 -2778
rect 1843 -2779 1844 -2778
rect 72 -2781 73 -2780
rect 236 -2781 237 -2780
rect 268 -2781 269 -2780
rect 674 -2781 675 -2780
rect 702 -2781 703 -2780
rect 1500 -2781 1501 -2780
rect 1710 -2781 1711 -2780
rect 1801 -2781 1802 -2780
rect 198 -2783 199 -2782
rect 947 -2783 948 -2782
rect 961 -2783 962 -2782
rect 2039 -2783 2040 -2782
rect 198 -2785 199 -2784
rect 1451 -2785 1452 -2784
rect 1794 -2785 1795 -2784
rect 1801 -2785 1802 -2784
rect 2039 -2785 2040 -2784
rect 2074 -2785 2075 -2784
rect 219 -2787 220 -2786
rect 268 -2787 269 -2786
rect 611 -2787 612 -2786
rect 639 -2787 640 -2786
rect 789 -2787 790 -2786
rect 1640 -2787 1641 -2786
rect 1794 -2787 1795 -2786
rect 1808 -2787 1809 -2786
rect 2074 -2787 2075 -2786
rect 2116 -2787 2117 -2786
rect 100 -2789 101 -2788
rect 611 -2789 612 -2788
rect 800 -2789 801 -2788
rect 1328 -2789 1329 -2788
rect 1703 -2789 1704 -2788
rect 1808 -2789 1809 -2788
rect 100 -2791 101 -2790
rect 247 -2791 248 -2790
rect 380 -2791 381 -2790
rect 800 -2791 801 -2790
rect 807 -2791 808 -2790
rect 2046 -2791 2047 -2790
rect 219 -2793 220 -2792
rect 898 -2793 899 -2792
rect 940 -2793 941 -2792
rect 1843 -2793 1844 -2792
rect 380 -2795 381 -2794
rect 618 -2795 619 -2794
rect 807 -2795 808 -2794
rect 828 -2795 829 -2794
rect 835 -2795 836 -2794
rect 922 -2795 923 -2794
rect 1003 -2795 1004 -2794
rect 1024 -2795 1025 -2794
rect 1164 -2795 1165 -2794
rect 1199 -2795 1200 -2794
rect 810 -2797 811 -2796
rect 2193 -2797 2194 -2796
rect 814 -2799 815 -2798
rect 1381 -2799 1382 -2798
rect 2186 -2799 2187 -2798
rect 2193 -2799 2194 -2798
rect 544 -2801 545 -2800
rect 2186 -2801 2187 -2800
rect 814 -2803 815 -2802
rect 884 -2803 885 -2802
rect 1017 -2803 1018 -2802
rect 1080 -2803 1081 -2802
rect 1199 -2803 1200 -2802
rect 1339 -2803 1340 -2802
rect 1381 -2803 1382 -2802
rect 1612 -2803 1613 -2802
rect 394 -2805 395 -2804
rect 884 -2805 885 -2804
rect 1024 -2805 1025 -2804
rect 1755 -2805 1756 -2804
rect 394 -2807 395 -2806
rect 457 -2807 458 -2806
rect 821 -2807 822 -2806
rect 905 -2807 906 -2806
rect 1080 -2807 1081 -2806
rect 1248 -2807 1249 -2806
rect 1339 -2807 1340 -2806
rect 1346 -2807 1347 -2806
rect 1409 -2807 1410 -2806
rect 1612 -2807 1613 -2806
rect 618 -2809 619 -2808
rect 1248 -2809 1249 -2808
rect 1346 -2809 1347 -2808
rect 1969 -2809 1970 -2808
rect 824 -2811 825 -2810
rect 1780 -2811 1781 -2810
rect 1969 -2811 1970 -2810
rect 1990 -2811 1991 -2810
rect 828 -2813 829 -2812
rect 1052 -2813 1053 -2812
rect 1409 -2813 1410 -2812
rect 1416 -2813 1417 -2812
rect 1815 -2813 1816 -2812
rect 1990 -2813 1991 -2812
rect 835 -2815 836 -2814
rect 926 -2815 927 -2814
rect 1052 -2815 1053 -2814
rect 1836 -2815 1837 -2814
rect 191 -2817 192 -2816
rect 926 -2817 927 -2816
rect 1815 -2817 1816 -2816
rect 1822 -2817 1823 -2816
rect 1836 -2817 1837 -2816
rect 1920 -2817 1921 -2816
rect 191 -2819 192 -2818
rect 534 -2819 535 -2818
rect 866 -2819 867 -2818
rect 2116 -2819 2117 -2818
rect 275 -2821 276 -2820
rect 534 -2821 535 -2820
rect 894 -2821 895 -2820
rect 1416 -2821 1417 -2820
rect 1535 -2821 1536 -2820
rect 1920 -2821 1921 -2820
rect 275 -2823 276 -2822
rect 499 -2823 500 -2822
rect 905 -2823 906 -2822
rect 1304 -2823 1305 -2822
rect 1822 -2823 1823 -2822
rect 1829 -2823 1830 -2822
rect 485 -2825 486 -2824
rect 499 -2825 500 -2824
rect 989 -2825 990 -2824
rect 1535 -2825 1536 -2824
rect 1829 -2825 1830 -2824
rect 1997 -2825 1998 -2824
rect 429 -2827 430 -2826
rect 485 -2827 486 -2826
rect 989 -2827 990 -2826
rect 1094 -2827 1095 -2826
rect 1304 -2827 1305 -2826
rect 1311 -2827 1312 -2826
rect 1997 -2827 1998 -2826
rect 2025 -2827 2026 -2826
rect 240 -2829 241 -2828
rect 1094 -2829 1095 -2828
rect 2025 -2829 2026 -2828
rect 2067 -2829 2068 -2828
rect 1941 -2831 1942 -2830
rect 2067 -2831 2068 -2830
rect 222 -2833 223 -2832
rect 1941 -2833 1942 -2832
rect 23 -2844 24 -2843
rect 467 -2844 468 -2843
rect 541 -2844 542 -2843
rect 1496 -2844 1497 -2843
rect 1500 -2844 1501 -2843
rect 2256 -2844 2257 -2843
rect 23 -2846 24 -2845
rect 184 -2846 185 -2845
rect 219 -2846 220 -2845
rect 380 -2846 381 -2845
rect 429 -2846 430 -2845
rect 492 -2846 493 -2845
rect 548 -2846 549 -2845
rect 786 -2846 787 -2845
rect 814 -2846 815 -2845
rect 940 -2846 941 -2845
rect 943 -2846 944 -2845
rect 1332 -2846 1333 -2845
rect 1346 -2846 1347 -2845
rect 1633 -2846 1634 -2845
rect 1682 -2846 1683 -2845
rect 2137 -2846 2138 -2845
rect 2221 -2846 2222 -2845
rect 2249 -2846 2250 -2845
rect 30 -2848 31 -2847
rect 544 -2848 545 -2847
rect 548 -2848 549 -2847
rect 891 -2848 892 -2847
rect 919 -2848 920 -2847
rect 1139 -2848 1140 -2847
rect 1202 -2848 1203 -2847
rect 1209 -2848 1210 -2847
rect 1255 -2848 1256 -2847
rect 1325 -2848 1326 -2847
rect 1332 -2848 1333 -2847
rect 1619 -2848 1620 -2847
rect 1682 -2848 1683 -2847
rect 2060 -2848 2061 -2847
rect 2074 -2848 2075 -2847
rect 2137 -2848 2138 -2847
rect 30 -2850 31 -2849
rect 257 -2850 258 -2849
rect 317 -2850 318 -2849
rect 789 -2850 790 -2849
rect 828 -2850 829 -2849
rect 891 -2850 892 -2849
rect 922 -2850 923 -2849
rect 1500 -2850 1501 -2849
rect 1566 -2850 1567 -2849
rect 2004 -2850 2005 -2849
rect 2060 -2850 2061 -2849
rect 2207 -2850 2208 -2849
rect 51 -2852 52 -2851
rect 478 -2852 479 -2851
rect 492 -2852 493 -2851
rect 527 -2852 528 -2851
rect 544 -2852 545 -2851
rect 912 -2852 913 -2851
rect 964 -2852 965 -2851
rect 1234 -2852 1235 -2851
rect 1258 -2852 1259 -2851
rect 1920 -2852 1921 -2851
rect 2004 -2852 2005 -2851
rect 2102 -2852 2103 -2851
rect 82 -2854 83 -2853
rect 408 -2854 409 -2853
rect 457 -2854 458 -2853
rect 499 -2854 500 -2853
rect 527 -2854 528 -2853
rect 737 -2854 738 -2853
rect 744 -2854 745 -2853
rect 842 -2854 843 -2853
rect 863 -2854 864 -2853
rect 1983 -2854 1984 -2853
rect 2074 -2854 2075 -2853
rect 2214 -2854 2215 -2853
rect 103 -2856 104 -2855
rect 352 -2856 353 -2855
rect 373 -2856 374 -2855
rect 408 -2856 409 -2855
rect 460 -2856 461 -2855
rect 555 -2856 556 -2855
rect 565 -2856 566 -2855
rect 940 -2856 941 -2855
rect 968 -2856 969 -2855
rect 971 -2856 972 -2855
rect 975 -2856 976 -2855
rect 1374 -2856 1375 -2855
rect 1391 -2856 1392 -2855
rect 1850 -2856 1851 -2855
rect 1983 -2856 1984 -2855
rect 2088 -2856 2089 -2855
rect 2098 -2856 2099 -2855
rect 2102 -2856 2103 -2855
rect 107 -2858 108 -2857
rect 387 -2858 388 -2857
rect 401 -2858 402 -2857
rect 814 -2858 815 -2857
rect 835 -2858 836 -2857
rect 926 -2858 927 -2857
rect 968 -2858 969 -2857
rect 982 -2858 983 -2857
rect 1017 -2858 1018 -2857
rect 1059 -2858 1060 -2857
rect 1062 -2858 1063 -2857
rect 1087 -2858 1088 -2857
rect 1136 -2858 1137 -2857
rect 1619 -2858 1620 -2857
rect 1703 -2858 1704 -2857
rect 2032 -2858 2033 -2857
rect 2088 -2858 2089 -2857
rect 2235 -2858 2236 -2857
rect 117 -2860 118 -2859
rect 1892 -2860 1893 -2859
rect 2032 -2860 2033 -2859
rect 2151 -2860 2152 -2859
rect 124 -2862 125 -2861
rect 856 -2862 857 -2861
rect 866 -2862 867 -2861
rect 1097 -2862 1098 -2861
rect 1234 -2862 1235 -2861
rect 1290 -2862 1291 -2861
rect 1314 -2862 1315 -2861
rect 1556 -2862 1557 -2861
rect 1703 -2862 1704 -2861
rect 1773 -2862 1774 -2861
rect 1850 -2862 1851 -2861
rect 1997 -2862 1998 -2861
rect 191 -2864 192 -2863
rect 401 -2864 402 -2863
rect 485 -2864 486 -2863
rect 555 -2864 556 -2863
rect 597 -2864 598 -2863
rect 660 -2864 661 -2863
rect 674 -2864 675 -2863
rect 926 -2864 927 -2863
rect 971 -2864 972 -2863
rect 982 -2864 983 -2863
rect 1017 -2864 1018 -2863
rect 1136 -2864 1137 -2863
rect 1283 -2864 1284 -2863
rect 1381 -2864 1382 -2863
rect 1433 -2864 1434 -2863
rect 1717 -2864 1718 -2863
rect 1731 -2864 1732 -2863
rect 1920 -2864 1921 -2863
rect 128 -2866 129 -2865
rect 597 -2866 598 -2865
rect 611 -2866 612 -2865
rect 1125 -2866 1126 -2865
rect 1286 -2866 1287 -2865
rect 1696 -2866 1697 -2865
rect 1706 -2866 1707 -2865
rect 2018 -2866 2019 -2865
rect 86 -2868 87 -2867
rect 128 -2868 129 -2867
rect 191 -2868 192 -2867
rect 212 -2868 213 -2867
rect 219 -2868 220 -2867
rect 443 -2868 444 -2867
rect 485 -2868 486 -2867
rect 520 -2868 521 -2867
rect 583 -2868 584 -2867
rect 611 -2868 612 -2867
rect 621 -2868 622 -2867
rect 800 -2868 801 -2867
rect 856 -2868 857 -2867
rect 1241 -2868 1242 -2867
rect 1290 -2868 1291 -2867
rect 1339 -2868 1340 -2867
rect 1346 -2868 1347 -2867
rect 1472 -2868 1473 -2867
rect 1486 -2868 1487 -2867
rect 2109 -2868 2110 -2867
rect 86 -2870 87 -2869
rect 247 -2870 248 -2869
rect 250 -2870 251 -2869
rect 1402 -2870 1403 -2869
rect 1419 -2870 1420 -2869
rect 1472 -2870 1473 -2869
rect 1489 -2870 1490 -2869
rect 1633 -2870 1634 -2869
rect 1696 -2870 1697 -2869
rect 1815 -2870 1816 -2869
rect 1878 -2870 1879 -2869
rect 1997 -2870 1998 -2869
rect 2018 -2870 2019 -2869
rect 2123 -2870 2124 -2869
rect 72 -2872 73 -2871
rect 247 -2872 248 -2871
rect 289 -2872 290 -2871
rect 317 -2872 318 -2871
rect 324 -2872 325 -2871
rect 429 -2872 430 -2871
rect 443 -2872 444 -2871
rect 471 -2872 472 -2871
rect 499 -2872 500 -2871
rect 604 -2872 605 -2871
rect 674 -2872 675 -2871
rect 1311 -2872 1312 -2871
rect 1314 -2872 1315 -2871
rect 2200 -2872 2201 -2871
rect 58 -2874 59 -2873
rect 72 -2874 73 -2873
rect 135 -2874 136 -2873
rect 604 -2874 605 -2873
rect 681 -2874 682 -2873
rect 912 -2874 913 -2873
rect 1038 -2874 1039 -2873
rect 1349 -2874 1350 -2873
rect 1360 -2874 1361 -2873
rect 1363 -2874 1364 -2873
rect 1374 -2874 1375 -2873
rect 1423 -2874 1424 -2873
rect 1451 -2874 1452 -2873
rect 2193 -2874 2194 -2873
rect 58 -2876 59 -2875
rect 1248 -2876 1249 -2875
rect 1339 -2876 1340 -2875
rect 1367 -2876 1368 -2875
rect 1381 -2876 1382 -2875
rect 1437 -2876 1438 -2875
rect 1493 -2876 1494 -2875
rect 1685 -2876 1686 -2875
rect 1717 -2876 1718 -2875
rect 1857 -2876 1858 -2875
rect 1892 -2876 1893 -2875
rect 1976 -2876 1977 -2875
rect 2109 -2876 2110 -2875
rect 2242 -2876 2243 -2875
rect 100 -2878 101 -2877
rect 1367 -2878 1368 -2877
rect 1402 -2878 1403 -2877
rect 1409 -2878 1410 -2877
rect 1437 -2878 1438 -2877
rect 2270 -2878 2271 -2877
rect 100 -2880 101 -2879
rect 1731 -2880 1732 -2879
rect 1752 -2880 1753 -2879
rect 1906 -2880 1907 -2879
rect 1976 -2880 1977 -2879
rect 2179 -2880 2180 -2879
rect 110 -2882 111 -2881
rect 1409 -2882 1410 -2881
rect 1493 -2882 1494 -2881
rect 1542 -2882 1543 -2881
rect 1556 -2882 1557 -2881
rect 1640 -2882 1641 -2881
rect 1752 -2882 1753 -2881
rect 1871 -2882 1872 -2881
rect 1906 -2882 1907 -2881
rect 2011 -2882 2012 -2881
rect 2123 -2882 2124 -2881
rect 2224 -2882 2225 -2881
rect 135 -2884 136 -2883
rect 576 -2884 577 -2883
rect 583 -2884 584 -2883
rect 849 -2884 850 -2883
rect 880 -2884 881 -2883
rect 1101 -2884 1102 -2883
rect 1115 -2884 1116 -2883
rect 1423 -2884 1424 -2883
rect 1444 -2884 1445 -2883
rect 1542 -2884 1543 -2883
rect 1640 -2884 1641 -2883
rect 1759 -2884 1760 -2883
rect 1773 -2884 1774 -2883
rect 1885 -2884 1886 -2883
rect 2011 -2884 2012 -2883
rect 2116 -2884 2117 -2883
rect 65 -2886 66 -2885
rect 849 -2886 850 -2885
rect 961 -2886 962 -2885
rect 2116 -2886 2117 -2885
rect 205 -2888 206 -2887
rect 478 -2888 479 -2887
rect 520 -2888 521 -2887
rect 1052 -2888 1053 -2887
rect 1059 -2888 1060 -2887
rect 1458 -2888 1459 -2887
rect 1755 -2888 1756 -2887
rect 1990 -2888 1991 -2887
rect 2 -2890 3 -2889
rect 205 -2890 206 -2889
rect 212 -2890 213 -2889
rect 632 -2890 633 -2889
rect 642 -2890 643 -2889
rect 1451 -2890 1452 -2889
rect 1759 -2890 1760 -2889
rect 1829 -2890 1830 -2889
rect 1871 -2890 1872 -2889
rect 2259 -2890 2260 -2889
rect 222 -2892 223 -2891
rect 2046 -2892 2047 -2891
rect 233 -2894 234 -2893
rect 303 -2894 304 -2893
rect 310 -2894 311 -2893
rect 352 -2894 353 -2893
rect 373 -2894 374 -2893
rect 415 -2894 416 -2893
rect 576 -2894 577 -2893
rect 1416 -2894 1417 -2893
rect 1444 -2894 1445 -2893
rect 1479 -2894 1480 -2893
rect 1801 -2894 1802 -2893
rect 1878 -2894 1879 -2893
rect 1990 -2894 1991 -2893
rect 2095 -2894 2096 -2893
rect 233 -2896 234 -2895
rect 268 -2896 269 -2895
rect 289 -2896 290 -2895
rect 534 -2896 535 -2895
rect 590 -2896 591 -2895
rect 681 -2896 682 -2895
rect 688 -2896 689 -2895
rect 828 -2896 829 -2895
rect 961 -2896 962 -2895
rect 2151 -2896 2152 -2895
rect 163 -2898 164 -2897
rect 268 -2898 269 -2897
rect 275 -2898 276 -2897
rect 534 -2898 535 -2897
rect 590 -2898 591 -2897
rect 807 -2898 808 -2897
rect 978 -2898 979 -2897
rect 1885 -2898 1886 -2897
rect 2046 -2898 2047 -2897
rect 2165 -2898 2166 -2897
rect 163 -2900 164 -2899
rect 933 -2900 934 -2899
rect 1010 -2900 1011 -2899
rect 1458 -2900 1459 -2899
rect 1479 -2900 1480 -2899
rect 1598 -2900 1599 -2899
rect 1801 -2900 1802 -2899
rect 1941 -2900 1942 -2899
rect 236 -2902 237 -2901
rect 303 -2902 304 -2901
rect 310 -2902 311 -2901
rect 422 -2902 423 -2901
rect 632 -2902 633 -2901
rect 723 -2902 724 -2901
rect 730 -2902 731 -2901
rect 1388 -2902 1389 -2901
rect 1598 -2902 1599 -2901
rect 1612 -2902 1613 -2901
rect 1815 -2902 1816 -2901
rect 1836 -2902 1837 -2901
rect 1941 -2902 1942 -2901
rect 2039 -2902 2040 -2901
rect 16 -2904 17 -2903
rect 730 -2904 731 -2903
rect 744 -2904 745 -2903
rect 1073 -2904 1074 -2903
rect 1087 -2904 1088 -2903
rect 1122 -2904 1123 -2903
rect 1199 -2904 1200 -2903
rect 1857 -2904 1858 -2903
rect 2039 -2904 2040 -2903
rect 2158 -2904 2159 -2903
rect 37 -2906 38 -2905
rect 723 -2906 724 -2905
rect 747 -2906 748 -2905
rect 947 -2906 948 -2905
rect 954 -2906 955 -2905
rect 1122 -2906 1123 -2905
rect 1241 -2906 1242 -2905
rect 1297 -2906 1298 -2905
rect 1360 -2906 1361 -2905
rect 1521 -2906 1522 -2905
rect 1612 -2906 1613 -2905
rect 1675 -2906 1676 -2905
rect 1829 -2906 1830 -2905
rect 1948 -2906 1949 -2905
rect 37 -2908 38 -2907
rect 142 -2908 143 -2907
rect 275 -2908 276 -2907
rect 366 -2908 367 -2907
rect 380 -2908 381 -2907
rect 733 -2908 734 -2907
rect 737 -2908 738 -2907
rect 1675 -2908 1676 -2907
rect 1836 -2908 1837 -2907
rect 1913 -2908 1914 -2907
rect 142 -2910 143 -2909
rect 765 -2910 766 -2909
rect 772 -2910 773 -2909
rect 863 -2910 864 -2909
rect 933 -2910 934 -2909
rect 1094 -2910 1095 -2909
rect 1101 -2910 1102 -2909
rect 1143 -2910 1144 -2909
rect 1248 -2910 1249 -2909
rect 1276 -2910 1277 -2909
rect 1297 -2910 1298 -2909
rect 1395 -2910 1396 -2909
rect 1521 -2910 1522 -2909
rect 1626 -2910 1627 -2909
rect 1913 -2910 1914 -2909
rect 2025 -2910 2026 -2909
rect 324 -2912 325 -2911
rect 394 -2912 395 -2911
rect 415 -2912 416 -2911
rect 1055 -2912 1056 -2911
rect 1066 -2912 1067 -2911
rect 1325 -2912 1326 -2911
rect 1388 -2912 1389 -2911
rect 1465 -2912 1466 -2911
rect 2025 -2912 2026 -2911
rect 2130 -2912 2131 -2911
rect 44 -2914 45 -2913
rect 1066 -2914 1067 -2913
rect 1069 -2914 1070 -2913
rect 1654 -2914 1655 -2913
rect 2130 -2914 2131 -2913
rect 2263 -2914 2264 -2913
rect 44 -2916 45 -2915
rect 618 -2916 619 -2915
rect 646 -2916 647 -2915
rect 807 -2916 808 -2915
rect 842 -2916 843 -2915
rect 1199 -2916 1200 -2915
rect 1276 -2916 1277 -2915
rect 1353 -2916 1354 -2915
rect 1395 -2916 1396 -2915
rect 1507 -2916 1508 -2915
rect 1654 -2916 1655 -2915
rect 1689 -2916 1690 -2915
rect 9 -2918 10 -2917
rect 618 -2918 619 -2917
rect 660 -2918 661 -2917
rect 1626 -2918 1627 -2917
rect 1689 -2918 1690 -2917
rect 1745 -2918 1746 -2917
rect 198 -2920 199 -2919
rect 394 -2920 395 -2919
rect 422 -2920 423 -2919
rect 464 -2920 465 -2919
rect 562 -2920 563 -2919
rect 646 -2920 647 -2919
rect 663 -2920 664 -2919
rect 947 -2920 948 -2919
rect 954 -2920 955 -2919
rect 1038 -2920 1039 -2919
rect 1045 -2920 1046 -2919
rect 1486 -2920 1487 -2919
rect 1507 -2920 1508 -2919
rect 1591 -2920 1592 -2919
rect 1745 -2920 1746 -2919
rect 1864 -2920 1865 -2919
rect 65 -2922 66 -2921
rect 464 -2922 465 -2921
rect 506 -2922 507 -2921
rect 562 -2922 563 -2921
rect 663 -2922 664 -2921
rect 1178 -2922 1179 -2921
rect 1465 -2922 1466 -2921
rect 1577 -2922 1578 -2921
rect 1710 -2922 1711 -2921
rect 1864 -2922 1865 -2921
rect 121 -2924 122 -2923
rect 506 -2924 507 -2923
rect 688 -2924 689 -2923
rect 1171 -2924 1172 -2923
rect 1178 -2924 1179 -2923
rect 1304 -2924 1305 -2923
rect 1430 -2924 1431 -2923
rect 1577 -2924 1578 -2923
rect 1710 -2924 1711 -2923
rect 1794 -2924 1795 -2923
rect 121 -2926 122 -2925
rect 184 -2926 185 -2925
rect 331 -2926 332 -2925
rect 471 -2926 472 -2925
rect 702 -2926 703 -2925
rect 1157 -2926 1158 -2925
rect 1171 -2926 1172 -2925
rect 1213 -2926 1214 -2925
rect 1304 -2926 1305 -2925
rect 1843 -2926 1844 -2925
rect 149 -2928 150 -2927
rect 198 -2928 199 -2927
rect 240 -2928 241 -2927
rect 331 -2928 332 -2927
rect 345 -2928 346 -2927
rect 366 -2928 367 -2927
rect 387 -2928 388 -2927
rect 1055 -2928 1056 -2927
rect 1073 -2928 1074 -2927
rect 1129 -2928 1130 -2927
rect 1213 -2928 1214 -2927
rect 1262 -2928 1263 -2927
rect 1430 -2928 1431 -2927
rect 1528 -2928 1529 -2927
rect 1570 -2928 1571 -2927
rect 1591 -2928 1592 -2927
rect 1794 -2928 1795 -2927
rect 1955 -2928 1956 -2927
rect 149 -2930 150 -2929
rect 1024 -2930 1025 -2929
rect 1031 -2930 1032 -2929
rect 1045 -2930 1046 -2929
rect 1080 -2930 1081 -2929
rect 1353 -2930 1354 -2929
rect 1528 -2930 1529 -2929
rect 1584 -2930 1585 -2929
rect 1843 -2930 1844 -2929
rect 1962 -2930 1963 -2929
rect 156 -2932 157 -2931
rect 240 -2932 241 -2931
rect 345 -2932 346 -2931
rect 793 -2932 794 -2931
rect 989 -2932 990 -2931
rect 1024 -2932 1025 -2931
rect 1080 -2932 1081 -2931
rect 1661 -2932 1662 -2931
rect 1955 -2932 1956 -2931
rect 2067 -2932 2068 -2931
rect 513 -2934 514 -2933
rect 1129 -2934 1130 -2933
rect 1192 -2934 1193 -2933
rect 1262 -2934 1263 -2933
rect 1514 -2934 1515 -2933
rect 1584 -2934 1585 -2933
rect 1661 -2934 1662 -2933
rect 1738 -2934 1739 -2933
rect 1962 -2934 1963 -2933
rect 2081 -2934 2082 -2933
rect 296 -2936 297 -2935
rect 513 -2936 514 -2935
rect 569 -2936 570 -2935
rect 702 -2936 703 -2935
rect 705 -2936 706 -2935
rect 884 -2936 885 -2935
rect 989 -2936 990 -2935
rect 1031 -2936 1032 -2935
rect 1094 -2936 1095 -2935
rect 1143 -2936 1144 -2935
rect 1192 -2936 1193 -2935
rect 1269 -2936 1270 -2935
rect 1514 -2936 1515 -2935
rect 1605 -2936 1606 -2935
rect 1738 -2936 1739 -2935
rect 2095 -2936 2096 -2935
rect 54 -2938 55 -2937
rect 1269 -2938 1270 -2937
rect 1605 -2938 1606 -2937
rect 1668 -2938 1669 -2937
rect 2067 -2938 2068 -2937
rect 2186 -2938 2187 -2937
rect 170 -2940 171 -2939
rect 569 -2940 570 -2939
rect 709 -2940 710 -2939
rect 884 -2940 885 -2939
rect 1010 -2940 1011 -2939
rect 1206 -2940 1207 -2939
rect 1668 -2940 1669 -2939
rect 1787 -2940 1788 -2939
rect 2081 -2940 2082 -2939
rect 2228 -2940 2229 -2939
rect 170 -2942 171 -2941
rect 261 -2942 262 -2941
rect 296 -2942 297 -2941
rect 338 -2942 339 -2941
rect 695 -2942 696 -2941
rect 709 -2942 710 -2941
rect 740 -2942 741 -2941
rect 1948 -2942 1949 -2941
rect 254 -2944 255 -2943
rect 338 -2944 339 -2943
rect 667 -2944 668 -2943
rect 695 -2944 696 -2943
rect 751 -2944 752 -2943
rect 1563 -2944 1564 -2943
rect 1787 -2944 1788 -2943
rect 1934 -2944 1935 -2943
rect 16 -2946 17 -2945
rect 254 -2946 255 -2945
rect 261 -2946 262 -2945
rect 359 -2946 360 -2945
rect 667 -2946 668 -2945
rect 1570 -2946 1571 -2945
rect 177 -2948 178 -2947
rect 751 -2948 752 -2947
rect 765 -2948 766 -2947
rect 1150 -2948 1151 -2947
rect 1157 -2948 1158 -2947
rect 1934 -2948 1935 -2947
rect 177 -2950 178 -2949
rect 215 -2950 216 -2949
rect 226 -2950 227 -2949
rect 359 -2950 360 -2949
rect 772 -2950 773 -2949
rect 1003 -2950 1004 -2949
rect 1115 -2950 1116 -2949
rect 1164 -2950 1165 -2949
rect 1206 -2950 1207 -2949
rect 1535 -2950 1536 -2949
rect 1563 -2950 1564 -2949
rect 1647 -2950 1648 -2949
rect 159 -2952 160 -2951
rect 226 -2952 227 -2951
rect 779 -2952 780 -2951
rect 800 -2952 801 -2951
rect 870 -2952 871 -2951
rect 1003 -2952 1004 -2951
rect 1150 -2952 1151 -2951
rect 1185 -2952 1186 -2951
rect 1535 -2952 1536 -2951
rect 1724 -2952 1725 -2951
rect 779 -2954 780 -2953
rect 877 -2954 878 -2953
rect 905 -2954 906 -2953
rect 1164 -2954 1165 -2953
rect 1185 -2954 1186 -2953
rect 1220 -2954 1221 -2953
rect 1647 -2954 1648 -2953
rect 1780 -2954 1781 -2953
rect 93 -2956 94 -2955
rect 905 -2956 906 -2955
rect 1097 -2956 1098 -2955
rect 1220 -2956 1221 -2955
rect 1724 -2956 1725 -2955
rect 1822 -2956 1823 -2955
rect 79 -2958 80 -2957
rect 93 -2958 94 -2957
rect 793 -2958 794 -2957
rect 821 -2958 822 -2957
rect 870 -2958 871 -2957
rect 898 -2958 899 -2957
rect 1780 -2958 1781 -2957
rect 1927 -2958 1928 -2957
rect 79 -2960 80 -2959
rect 996 -2960 997 -2959
rect 1822 -2960 1823 -2959
rect 1969 -2960 1970 -2959
rect 114 -2962 115 -2961
rect 898 -2962 899 -2961
rect 996 -2962 997 -2961
rect 1108 -2962 1109 -2961
rect 1927 -2962 1928 -2961
rect 2053 -2962 2054 -2961
rect 114 -2964 115 -2963
rect 450 -2964 451 -2963
rect 758 -2964 759 -2963
rect 821 -2964 822 -2963
rect 1108 -2964 1109 -2963
rect 1227 -2964 1228 -2963
rect 1808 -2964 1809 -2963
rect 2053 -2964 2054 -2963
rect 450 -2966 451 -2965
rect 1041 -2966 1042 -2965
rect 1227 -2966 1228 -2965
rect 1318 -2966 1319 -2965
rect 1808 -2966 1809 -2965
rect 1899 -2966 1900 -2965
rect 1969 -2966 1970 -2965
rect 2172 -2966 2173 -2965
rect 653 -2968 654 -2967
rect 758 -2968 759 -2967
rect 1318 -2968 1319 -2967
rect 1549 -2968 1550 -2967
rect 1766 -2968 1767 -2967
rect 1899 -2968 1900 -2967
rect 639 -2970 640 -2969
rect 653 -2970 654 -2969
rect 1160 -2970 1161 -2969
rect 1549 -2970 1550 -2969
rect 282 -2972 283 -2971
rect 639 -2972 640 -2971
rect 282 -2974 283 -2973
rect 625 -2974 626 -2973
rect 625 -2976 626 -2975
rect 716 -2976 717 -2975
rect 716 -2978 717 -2977
rect 985 -2978 986 -2977
rect 16 -2989 17 -2988
rect 110 -2989 111 -2988
rect 114 -2989 115 -2988
rect 387 -2989 388 -2988
rect 422 -2989 423 -2988
rect 460 -2989 461 -2988
rect 471 -2989 472 -2988
rect 562 -2989 563 -2988
rect 569 -2989 570 -2988
rect 975 -2989 976 -2988
rect 1041 -2989 1042 -2988
rect 2060 -2989 2061 -2988
rect 2095 -2989 2096 -2988
rect 2137 -2989 2138 -2988
rect 51 -2991 52 -2990
rect 72 -2991 73 -2990
rect 100 -2991 101 -2990
rect 933 -2991 934 -2990
rect 961 -2991 962 -2990
rect 968 -2991 969 -2990
rect 1052 -2991 1053 -2990
rect 1325 -2991 1326 -2990
rect 1360 -2991 1361 -2990
rect 1409 -2991 1410 -2990
rect 1416 -2991 1417 -2990
rect 1857 -2991 1858 -2990
rect 1871 -2991 1872 -2990
rect 1874 -2991 1875 -2990
rect 2098 -2991 2099 -2990
rect 2116 -2991 2117 -2990
rect 37 -2993 38 -2992
rect 72 -2993 73 -2992
rect 93 -2993 94 -2992
rect 100 -2993 101 -2992
rect 107 -2993 108 -2992
rect 779 -2993 780 -2992
rect 880 -2993 881 -2992
rect 1689 -2993 1690 -2992
rect 1769 -2993 1770 -2992
rect 1815 -2993 1816 -2992
rect 1836 -2993 1837 -2992
rect 1857 -2993 1858 -2992
rect 1871 -2993 1872 -2992
rect 1990 -2993 1991 -2992
rect 30 -2995 31 -2994
rect 93 -2995 94 -2994
rect 142 -2995 143 -2994
rect 919 -2995 920 -2994
rect 964 -2995 965 -2994
rect 1031 -2995 1032 -2994
rect 1055 -2995 1056 -2994
rect 1836 -2995 1837 -2994
rect 1892 -2995 1893 -2994
rect 1990 -2995 1991 -2994
rect 30 -2997 31 -2996
rect 58 -2997 59 -2996
rect 65 -2997 66 -2996
rect 565 -2997 566 -2996
rect 572 -2997 573 -2996
rect 961 -2997 962 -2996
rect 968 -2997 969 -2996
rect 1087 -2997 1088 -2996
rect 1125 -2997 1126 -2996
rect 1493 -2997 1494 -2996
rect 1566 -2997 1567 -2996
rect 1885 -2997 1886 -2996
rect 37 -2999 38 -2998
rect 520 -2999 521 -2998
rect 541 -2999 542 -2998
rect 814 -2999 815 -2998
rect 884 -2999 885 -2998
rect 933 -2999 934 -2998
rect 1031 -2999 1032 -2998
rect 1185 -2999 1186 -2998
rect 1199 -2999 1200 -2998
rect 1976 -2999 1977 -2998
rect 44 -3001 45 -3000
rect 65 -3001 66 -3000
rect 135 -3001 136 -3000
rect 541 -3001 542 -3000
rect 590 -3001 591 -3000
rect 915 -3001 916 -3000
rect 954 -3001 955 -3000
rect 1185 -3001 1186 -3000
rect 1199 -3001 1200 -3000
rect 1248 -3001 1249 -3000
rect 1318 -3001 1319 -3000
rect 1416 -3001 1417 -3000
rect 1419 -3001 1420 -3000
rect 1920 -3001 1921 -3000
rect 1976 -3001 1977 -3000
rect 2102 -3001 2103 -3000
rect 58 -3003 59 -3002
rect 198 -3003 199 -3002
rect 208 -3003 209 -3002
rect 443 -3003 444 -3002
rect 471 -3003 472 -3002
rect 880 -3003 881 -3002
rect 894 -3003 895 -3002
rect 1878 -3003 1879 -3002
rect 1885 -3003 1886 -3002
rect 1983 -3003 1984 -3002
rect 142 -3005 143 -3004
rect 205 -3005 206 -3004
rect 212 -3005 213 -3004
rect 338 -3005 339 -3004
rect 422 -3005 423 -3004
rect 429 -3005 430 -3004
rect 443 -3005 444 -3004
rect 1276 -3005 1277 -3004
rect 1318 -3005 1319 -3004
rect 1339 -3005 1340 -3004
rect 1398 -3005 1399 -3004
rect 1941 -3005 1942 -3004
rect 86 -3007 87 -3006
rect 212 -3007 213 -3006
rect 236 -3007 237 -3006
rect 618 -3007 619 -3006
rect 642 -3007 643 -3006
rect 758 -3007 759 -3006
rect 786 -3007 787 -3006
rect 954 -3007 955 -3006
rect 1055 -3007 1056 -3006
rect 1703 -3007 1704 -3006
rect 1808 -3007 1809 -3006
rect 1881 -3007 1882 -3006
rect 1920 -3007 1921 -3006
rect 2025 -3007 2026 -3006
rect 86 -3009 87 -3008
rect 219 -3009 220 -3008
rect 240 -3009 241 -3008
rect 429 -3009 430 -3008
rect 478 -3009 479 -3008
rect 618 -3009 619 -3008
rect 688 -3009 689 -3008
rect 1038 -3009 1039 -3008
rect 1066 -3009 1067 -3008
rect 1094 -3009 1095 -3008
rect 1139 -3009 1140 -3008
rect 1633 -3009 1634 -3008
rect 1654 -3009 1655 -3008
rect 1941 -3009 1942 -3008
rect 131 -3011 132 -3010
rect 786 -3011 787 -3010
rect 905 -3011 906 -3010
rect 919 -3011 920 -3010
rect 1038 -3011 1039 -3010
rect 1220 -3011 1221 -3010
rect 1325 -3011 1326 -3010
rect 1559 -3011 1560 -3010
rect 1570 -3011 1571 -3010
rect 1864 -3011 1865 -3010
rect 149 -3013 150 -3012
rect 464 -3013 465 -3012
rect 478 -3013 479 -3012
rect 667 -3013 668 -3012
rect 688 -3013 689 -3012
rect 1255 -3013 1256 -3012
rect 1339 -3013 1340 -3012
rect 1430 -3013 1431 -3012
rect 1486 -3013 1487 -3012
rect 1766 -3013 1767 -3012
rect 1808 -3013 1809 -3012
rect 2053 -3013 2054 -3012
rect 138 -3015 139 -3014
rect 149 -3015 150 -3014
rect 156 -3015 157 -3014
rect 663 -3015 664 -3014
rect 667 -3015 668 -3014
rect 695 -3015 696 -3014
rect 716 -3015 717 -3014
rect 719 -3015 720 -3014
rect 730 -3015 731 -3014
rect 922 -3015 923 -3014
rect 1045 -3015 1046 -3014
rect 1066 -3015 1067 -3014
rect 1069 -3015 1070 -3014
rect 1213 -3015 1214 -3014
rect 1220 -3015 1221 -3014
rect 1227 -3015 1228 -3014
rect 1255 -3015 1256 -3014
rect 1269 -3015 1270 -3014
rect 1402 -3015 1403 -3014
rect 1405 -3015 1406 -3014
rect 1430 -3015 1431 -3014
rect 1500 -3015 1501 -3014
rect 1570 -3015 1571 -3014
rect 1605 -3015 1606 -3014
rect 1633 -3015 1634 -3014
rect 1675 -3015 1676 -3014
rect 1689 -3015 1690 -3014
rect 1773 -3015 1774 -3014
rect 1815 -3015 1816 -3014
rect 1948 -3015 1949 -3014
rect 156 -3017 157 -3016
rect 191 -3017 192 -3016
rect 198 -3017 199 -3016
rect 261 -3017 262 -3016
rect 282 -3017 283 -3016
rect 569 -3017 570 -3016
rect 590 -3017 591 -3016
rect 702 -3017 703 -3016
rect 716 -3017 717 -3016
rect 800 -3017 801 -3016
rect 849 -3017 850 -3016
rect 905 -3017 906 -3016
rect 1045 -3017 1046 -3016
rect 1143 -3017 1144 -3016
rect 1160 -3017 1161 -3016
rect 1353 -3017 1354 -3016
rect 1402 -3017 1403 -3016
rect 1528 -3017 1529 -3016
rect 1549 -3017 1550 -3016
rect 1675 -3017 1676 -3016
rect 1703 -3017 1704 -3016
rect 1780 -3017 1781 -3016
rect 1864 -3017 1865 -3016
rect 2039 -3017 2040 -3016
rect 128 -3019 129 -3018
rect 1160 -3019 1161 -3018
rect 1178 -3019 1179 -3018
rect 1206 -3019 1207 -3018
rect 1213 -3019 1214 -3018
rect 1423 -3019 1424 -3018
rect 1486 -3019 1487 -3018
rect 1563 -3019 1564 -3018
rect 1573 -3019 1574 -3018
rect 2130 -3019 2131 -3018
rect 159 -3021 160 -3020
rect 1073 -3021 1074 -3020
rect 1076 -3021 1077 -3020
rect 1437 -3021 1438 -3020
rect 1493 -3021 1494 -3020
rect 1521 -3021 1522 -3020
rect 1528 -3021 1529 -3020
rect 1682 -3021 1683 -3020
rect 1759 -3021 1760 -3020
rect 1780 -3021 1781 -3020
rect 1874 -3021 1875 -3020
rect 1892 -3021 1893 -3020
rect 1948 -3021 1949 -3020
rect 2088 -3021 2089 -3020
rect 163 -3023 164 -3022
rect 520 -3023 521 -3022
rect 597 -3023 598 -3022
rect 639 -3023 640 -3022
rect 695 -3023 696 -3022
rect 709 -3023 710 -3022
rect 730 -3023 731 -3022
rect 1080 -3023 1081 -3022
rect 1083 -3023 1084 -3022
rect 1934 -3023 1935 -3022
rect 166 -3025 167 -3024
rect 926 -3025 927 -3024
rect 1087 -3025 1088 -3024
rect 1115 -3025 1116 -3024
rect 1143 -3025 1144 -3024
rect 1304 -3025 1305 -3024
rect 1353 -3025 1354 -3024
rect 1395 -3025 1396 -3024
rect 1423 -3025 1424 -3024
rect 1479 -3025 1480 -3024
rect 1500 -3025 1501 -3024
rect 1556 -3025 1557 -3024
rect 1654 -3025 1655 -3024
rect 1745 -3025 1746 -3024
rect 1759 -3025 1760 -3024
rect 1850 -3025 1851 -3024
rect 1934 -3025 1935 -3024
rect 2011 -3025 2012 -3024
rect 79 -3027 80 -3026
rect 926 -3027 927 -3026
rect 985 -3027 986 -3026
rect 1850 -3027 1851 -3026
rect 170 -3029 171 -3028
rect 261 -3029 262 -3028
rect 282 -3029 283 -3028
rect 380 -3029 381 -3028
rect 457 -3029 458 -3028
rect 597 -3029 598 -3028
rect 614 -3029 615 -3028
rect 898 -3029 899 -3028
rect 1178 -3029 1179 -3028
rect 1241 -3029 1242 -3028
rect 1269 -3029 1270 -3028
rect 1290 -3029 1291 -3028
rect 1304 -3029 1305 -3028
rect 1472 -3029 1473 -3028
rect 1549 -3029 1550 -3028
rect 1612 -3029 1613 -3028
rect 1661 -3029 1662 -3028
rect 1685 -3029 1686 -3028
rect 1745 -3029 1746 -3028
rect 1955 -3029 1956 -3028
rect 173 -3031 174 -3030
rect 604 -3031 605 -3030
rect 625 -3031 626 -3030
rect 1115 -3031 1116 -3030
rect 1192 -3031 1193 -3030
rect 1605 -3031 1606 -3030
rect 1612 -3031 1613 -3030
rect 1640 -3031 1641 -3030
rect 1661 -3031 1662 -3030
rect 1724 -3031 1725 -3030
rect 1766 -3031 1767 -3030
rect 1843 -3031 1844 -3030
rect 184 -3033 185 -3032
rect 191 -3033 192 -3032
rect 219 -3033 220 -3032
rect 373 -3033 374 -3032
rect 457 -3033 458 -3032
rect 975 -3033 976 -3032
rect 1164 -3033 1165 -3032
rect 1192 -3033 1193 -3032
rect 1202 -3033 1203 -3032
rect 1409 -3033 1410 -3032
rect 1437 -3033 1438 -3032
rect 1514 -3033 1515 -3032
rect 1598 -3033 1599 -3032
rect 1640 -3033 1641 -3032
rect 1682 -3033 1683 -3032
rect 1983 -3033 1984 -3032
rect 184 -3035 185 -3034
rect 205 -3035 206 -3034
rect 215 -3035 216 -3034
rect 373 -3035 374 -3034
rect 485 -3035 486 -3034
rect 737 -3035 738 -3034
rect 740 -3035 741 -3034
rect 870 -3035 871 -3034
rect 1136 -3035 1137 -3034
rect 1598 -3035 1599 -3034
rect 1724 -3035 1725 -3034
rect 2074 -3035 2075 -3034
rect 240 -3037 241 -3036
rect 268 -3037 269 -3036
rect 296 -3037 297 -3036
rect 660 -3037 661 -3036
rect 702 -3037 703 -3036
rect 723 -3037 724 -3036
rect 737 -3037 738 -3036
rect 912 -3037 913 -3036
rect 1136 -3037 1137 -3036
rect 1234 -3037 1235 -3036
rect 1241 -3037 1242 -3036
rect 1388 -3037 1389 -3036
rect 1451 -3037 1452 -3036
rect 1521 -3037 1522 -3036
rect 1773 -3037 1774 -3036
rect 1822 -3037 1823 -3036
rect 1843 -3037 1844 -3036
rect 2004 -3037 2005 -3036
rect 2074 -3037 2075 -3036
rect 2151 -3037 2152 -3036
rect 254 -3039 255 -3038
rect 1367 -3039 1368 -3038
rect 1388 -3039 1389 -3038
rect 1717 -3039 1718 -3038
rect 1822 -3039 1823 -3038
rect 2018 -3039 2019 -3038
rect 247 -3041 248 -3040
rect 254 -3041 255 -3040
rect 268 -3041 269 -3040
rect 1059 -3041 1060 -3040
rect 1157 -3041 1158 -3040
rect 1367 -3041 1368 -3040
rect 1451 -3041 1452 -3040
rect 1731 -3041 1732 -3040
rect 2004 -3041 2005 -3040
rect 2081 -3041 2082 -3040
rect 103 -3043 104 -3042
rect 247 -3043 248 -3042
rect 296 -3043 297 -3042
rect 401 -3043 402 -3042
rect 415 -3043 416 -3042
rect 723 -3043 724 -3042
rect 758 -3043 759 -3042
rect 817 -3043 818 -3042
rect 870 -3043 871 -3042
rect 947 -3043 948 -3042
rect 1017 -3043 1018 -3042
rect 1731 -3043 1732 -3042
rect 275 -3045 276 -3044
rect 401 -3045 402 -3044
rect 415 -3045 416 -3044
rect 506 -3045 507 -3044
rect 513 -3045 514 -3044
rect 779 -3045 780 -3044
rect 835 -3045 836 -3044
rect 947 -3045 948 -3044
rect 1003 -3045 1004 -3044
rect 1017 -3045 1018 -3044
rect 1059 -3045 1060 -3044
rect 1101 -3045 1102 -3044
rect 1164 -3045 1165 -3044
rect 1237 -3045 1238 -3044
rect 1283 -3045 1284 -3044
rect 1290 -3045 1291 -3044
rect 1332 -3045 1333 -3044
rect 1479 -3045 1480 -3044
rect 1514 -3045 1515 -3044
rect 1542 -3045 1543 -3044
rect 1717 -3045 1718 -3044
rect 1794 -3045 1795 -3044
rect 275 -3047 276 -3046
rect 324 -3047 325 -3046
rect 338 -3047 339 -3046
rect 366 -3047 367 -3046
rect 485 -3047 486 -3046
rect 555 -3047 556 -3046
rect 625 -3047 626 -3046
rect 674 -3047 675 -3046
rect 709 -3047 710 -3046
rect 1062 -3047 1063 -3046
rect 1097 -3047 1098 -3046
rect 1332 -3047 1333 -3046
rect 1465 -3047 1466 -3046
rect 1955 -3047 1956 -3046
rect 289 -3049 290 -3048
rect 555 -3049 556 -3048
rect 660 -3049 661 -3048
rect 681 -3049 682 -3048
rect 765 -3049 766 -3048
rect 849 -3049 850 -3048
rect 884 -3049 885 -3048
rect 1234 -3049 1235 -3048
rect 1283 -3049 1284 -3048
rect 1297 -3049 1298 -3048
rect 1465 -3049 1466 -3048
rect 1738 -3049 1739 -3048
rect 1794 -3049 1795 -3048
rect 1927 -3049 1928 -3048
rect 289 -3051 290 -3050
rect 632 -3051 633 -3050
rect 674 -3051 675 -3050
rect 1129 -3051 1130 -3050
rect 1227 -3051 1228 -3050
rect 1262 -3051 1263 -3050
rect 1297 -3051 1298 -3050
rect 1311 -3051 1312 -3050
rect 1472 -3051 1473 -3050
rect 1965 -3051 1966 -3050
rect 310 -3053 311 -3052
rect 387 -3053 388 -3052
rect 506 -3053 507 -3052
rect 996 -3053 997 -3052
rect 1024 -3053 1025 -3052
rect 1262 -3053 1263 -3052
rect 1311 -3053 1312 -3052
rect 1535 -3053 1536 -3052
rect 1542 -3053 1543 -3052
rect 1584 -3053 1585 -3052
rect 1738 -3053 1739 -3052
rect 1801 -3053 1802 -3052
rect 1927 -3053 1928 -3052
rect 2067 -3053 2068 -3052
rect 310 -3055 311 -3054
rect 1073 -3055 1074 -3054
rect 1101 -3055 1102 -3054
rect 1150 -3055 1151 -3054
rect 1535 -3055 1536 -3054
rect 1591 -3055 1592 -3054
rect 1801 -3055 1802 -3054
rect 1906 -3055 1907 -3054
rect 324 -3057 325 -3056
rect 499 -3057 500 -3056
rect 513 -3057 514 -3056
rect 534 -3057 535 -3056
rect 548 -3057 549 -3056
rect 1157 -3057 1158 -3056
rect 1584 -3057 1585 -3056
rect 1619 -3057 1620 -3056
rect 1906 -3057 1907 -3056
rect 2032 -3057 2033 -3056
rect 226 -3059 227 -3058
rect 534 -3059 535 -3058
rect 632 -3059 633 -3058
rect 828 -3059 829 -3058
rect 835 -3059 836 -3058
rect 1381 -3059 1382 -3058
rect 1591 -3059 1592 -3058
rect 1626 -3059 1627 -3058
rect 2032 -3059 2033 -3058
rect 2109 -3059 2110 -3058
rect 121 -3061 122 -3060
rect 226 -3061 227 -3060
rect 352 -3061 353 -3060
rect 548 -3061 549 -3060
rect 681 -3061 682 -3060
rect 842 -3061 843 -3060
rect 940 -3061 941 -3060
rect 1003 -3061 1004 -3060
rect 1024 -3061 1025 -3060
rect 1108 -3061 1109 -3060
rect 1122 -3061 1123 -3060
rect 1150 -3061 1151 -3060
rect 1381 -3061 1382 -3060
rect 1444 -3061 1445 -3060
rect 1619 -3061 1620 -3060
rect 1647 -3061 1648 -3060
rect 121 -3063 122 -3062
rect 576 -3063 577 -3062
rect 765 -3063 766 -3062
rect 856 -3063 857 -3062
rect 940 -3063 941 -3062
rect 1374 -3063 1375 -3062
rect 1626 -3063 1627 -3062
rect 1696 -3063 1697 -3062
rect 124 -3065 125 -3064
rect 352 -3065 353 -3064
rect 359 -3065 360 -3064
rect 380 -3065 381 -3064
rect 450 -3065 451 -3064
rect 828 -3065 829 -3064
rect 856 -3065 857 -3064
rect 863 -3065 864 -3064
rect 996 -3065 997 -3064
rect 1216 -3065 1217 -3064
rect 1556 -3065 1557 -3064
rect 1696 -3065 1697 -3064
rect 359 -3067 360 -3066
rect 544 -3067 545 -3066
rect 576 -3067 577 -3066
rect 653 -3067 654 -3066
rect 772 -3067 773 -3066
rect 898 -3067 899 -3066
rect 1010 -3067 1011 -3066
rect 1108 -3067 1109 -3066
rect 1129 -3067 1130 -3066
rect 1171 -3067 1172 -3066
rect 1647 -3067 1648 -3066
rect 1710 -3067 1711 -3066
rect 366 -3069 367 -3068
rect 394 -3069 395 -3068
rect 450 -3069 451 -3068
rect 492 -3069 493 -3068
rect 499 -3069 500 -3068
rect 1363 -3069 1364 -3068
rect 1710 -3069 1711 -3068
rect 1787 -3069 1788 -3068
rect 317 -3071 318 -3070
rect 394 -3071 395 -3070
rect 492 -3071 493 -3070
rect 646 -3071 647 -3070
rect 653 -3071 654 -3070
rect 891 -3071 892 -3070
rect 1034 -3071 1035 -3070
rect 1374 -3071 1375 -3070
rect 1787 -3071 1788 -3070
rect 1899 -3071 1900 -3070
rect 177 -3073 178 -3072
rect 317 -3073 318 -3072
rect 527 -3073 528 -3072
rect 604 -3073 605 -3072
rect 611 -3073 612 -3072
rect 646 -3073 647 -3072
rect 744 -3073 745 -3072
rect 1010 -3073 1011 -3072
rect 1171 -3073 1172 -3072
rect 1314 -3073 1315 -3072
rect 1899 -3073 1900 -3072
rect 1997 -3073 1998 -3072
rect 23 -3075 24 -3074
rect 611 -3075 612 -3074
rect 772 -3075 773 -3074
rect 821 -3075 822 -3074
rect 863 -3075 864 -3074
rect 1969 -3075 1970 -3074
rect 23 -3077 24 -3076
rect 982 -3077 983 -3076
rect 1507 -3077 1508 -3076
rect 1969 -3077 1970 -3076
rect 177 -3079 178 -3078
rect 303 -3079 304 -3078
rect 331 -3079 332 -3078
rect 821 -3079 822 -3078
rect 982 -3079 983 -3078
rect 989 -3079 990 -3078
rect 1507 -3079 1508 -3078
rect 1577 -3079 1578 -3078
rect 1913 -3079 1914 -3078
rect 1997 -3079 1998 -3078
rect 233 -3081 234 -3080
rect 303 -3081 304 -3080
rect 331 -3081 332 -3080
rect 345 -3081 346 -3080
rect 583 -3081 584 -3080
rect 744 -3081 745 -3080
rect 807 -3081 808 -3080
rect 842 -3081 843 -3080
rect 877 -3081 878 -3080
rect 1577 -3081 1578 -3080
rect 1913 -3081 1914 -3080
rect 2046 -3081 2047 -3080
rect 345 -3083 346 -3082
rect 408 -3083 409 -3082
rect 583 -3083 584 -3082
rect 751 -3083 752 -3082
rect 793 -3083 794 -3082
rect 807 -3083 808 -3082
rect 989 -3083 990 -3082
rect 1458 -3083 1459 -3082
rect 2046 -3083 2047 -3082
rect 2123 -3083 2124 -3082
rect 117 -3085 118 -3084
rect 408 -3085 409 -3084
rect 751 -3085 752 -3084
rect 912 -3085 913 -3084
rect 1458 -3085 1459 -3084
rect 1668 -3085 1669 -3084
rect 793 -3087 794 -3086
rect 1209 -3087 1210 -3086
rect 1668 -3087 1669 -3086
rect 1752 -3087 1753 -3086
rect 1752 -3089 1753 -3088
rect 1829 -3089 1830 -3088
rect 1829 -3091 1830 -3090
rect 1962 -3091 1963 -3090
rect 1962 -3093 1963 -3092
rect 2144 -3093 2145 -3092
rect 23 -3104 24 -3103
rect 208 -3104 209 -3103
rect 212 -3104 213 -3103
rect 233 -3104 234 -3103
rect 380 -3104 381 -3103
rect 457 -3104 458 -3103
rect 520 -3104 521 -3103
rect 817 -3104 818 -3103
rect 821 -3104 822 -3103
rect 1311 -3104 1312 -3103
rect 1381 -3104 1382 -3103
rect 1402 -3104 1403 -3103
rect 1461 -3104 1462 -3103
rect 1864 -3104 1865 -3103
rect 1962 -3104 1963 -3103
rect 2046 -3104 2047 -3103
rect 30 -3106 31 -3105
rect 205 -3106 206 -3105
rect 212 -3106 213 -3105
rect 1167 -3106 1168 -3105
rect 1199 -3106 1200 -3105
rect 1258 -3106 1259 -3105
rect 1276 -3106 1277 -3105
rect 1451 -3106 1452 -3105
rect 1465 -3106 1466 -3105
rect 1563 -3106 1564 -3105
rect 1566 -3106 1567 -3105
rect 1682 -3106 1683 -3105
rect 1853 -3106 1854 -3105
rect 1892 -3106 1893 -3105
rect 1997 -3106 1998 -3105
rect 2018 -3106 2019 -3105
rect 2046 -3106 2047 -3105
rect 2074 -3106 2075 -3105
rect 58 -3108 59 -3107
rect 131 -3108 132 -3107
rect 187 -3108 188 -3107
rect 688 -3108 689 -3107
rect 737 -3108 738 -3107
rect 1444 -3108 1445 -3107
rect 1451 -3108 1452 -3107
rect 1535 -3108 1536 -3107
rect 1640 -3108 1641 -3107
rect 1878 -3108 1879 -3107
rect 1892 -3108 1893 -3107
rect 1948 -3108 1949 -3107
rect 65 -3110 66 -3109
rect 1111 -3110 1112 -3109
rect 1199 -3110 1200 -3109
rect 1304 -3110 1305 -3109
rect 1311 -3110 1312 -3109
rect 1703 -3110 1704 -3109
rect 1864 -3110 1865 -3109
rect 1871 -3110 1872 -3109
rect 1878 -3110 1879 -3109
rect 1899 -3110 1900 -3109
rect 72 -3112 73 -3111
rect 236 -3112 237 -3111
rect 289 -3112 290 -3111
rect 821 -3112 822 -3111
rect 835 -3112 836 -3111
rect 1122 -3112 1123 -3111
rect 1216 -3112 1217 -3111
rect 1605 -3112 1606 -3111
rect 1671 -3112 1672 -3111
rect 1857 -3112 1858 -3111
rect 79 -3114 80 -3113
rect 674 -3114 675 -3113
rect 681 -3114 682 -3113
rect 1160 -3114 1161 -3113
rect 1234 -3114 1235 -3113
rect 1346 -3114 1347 -3113
rect 1381 -3114 1382 -3113
rect 1633 -3114 1634 -3113
rect 1675 -3114 1676 -3113
rect 1962 -3114 1963 -3113
rect 86 -3116 87 -3115
rect 138 -3116 139 -3115
rect 194 -3116 195 -3115
rect 282 -3116 283 -3115
rect 289 -3116 290 -3115
rect 425 -3116 426 -3115
rect 506 -3116 507 -3115
rect 737 -3116 738 -3115
rect 758 -3116 759 -3115
rect 1643 -3116 1644 -3115
rect 1857 -3116 1858 -3115
rect 1885 -3116 1886 -3115
rect 93 -3118 94 -3117
rect 142 -3118 143 -3117
rect 254 -3118 255 -3117
rect 282 -3118 283 -3117
rect 352 -3118 353 -3117
rect 1346 -3118 1347 -3117
rect 1395 -3118 1396 -3117
rect 1472 -3118 1473 -3117
rect 1486 -3118 1487 -3117
rect 1556 -3118 1557 -3117
rect 1605 -3118 1606 -3117
rect 1850 -3118 1851 -3117
rect 1885 -3118 1886 -3117
rect 1920 -3118 1921 -3117
rect 107 -3120 108 -3119
rect 880 -3120 881 -3119
rect 891 -3120 892 -3119
rect 1115 -3120 1116 -3119
rect 1122 -3120 1123 -3119
rect 1325 -3120 1326 -3119
rect 1395 -3120 1396 -3119
rect 1710 -3120 1711 -3119
rect 1920 -3120 1921 -3119
rect 1976 -3120 1977 -3119
rect 107 -3122 108 -3121
rect 177 -3122 178 -3121
rect 226 -3122 227 -3121
rect 352 -3122 353 -3121
rect 380 -3122 381 -3121
rect 579 -3122 580 -3121
rect 604 -3122 605 -3121
rect 877 -3122 878 -3121
rect 898 -3122 899 -3121
rect 1115 -3122 1116 -3121
rect 1237 -3122 1238 -3121
rect 1409 -3122 1410 -3121
rect 1437 -3122 1438 -3121
rect 1563 -3122 1564 -3121
rect 1633 -3122 1634 -3121
rect 1787 -3122 1788 -3121
rect 1976 -3122 1977 -3121
rect 2004 -3122 2005 -3121
rect 114 -3124 115 -3123
rect 166 -3124 167 -3123
rect 177 -3124 178 -3123
rect 807 -3124 808 -3123
rect 828 -3124 829 -3123
rect 891 -3124 892 -3123
rect 943 -3124 944 -3123
rect 1724 -3124 1725 -3123
rect 100 -3126 101 -3125
rect 114 -3126 115 -3125
rect 121 -3126 122 -3125
rect 208 -3126 209 -3125
rect 254 -3126 255 -3125
rect 359 -3126 360 -3125
rect 401 -3126 402 -3125
rect 530 -3126 531 -3125
rect 555 -3126 556 -3125
rect 873 -3126 874 -3125
rect 877 -3126 878 -3125
rect 1447 -3126 1448 -3125
rect 1465 -3126 1466 -3125
rect 1612 -3126 1613 -3125
rect 1647 -3126 1648 -3125
rect 1724 -3126 1725 -3125
rect 100 -3128 101 -3127
rect 310 -3128 311 -3127
rect 359 -3128 360 -3127
rect 366 -3128 367 -3127
rect 373 -3128 374 -3127
rect 555 -3128 556 -3127
rect 569 -3128 570 -3127
rect 817 -3128 818 -3127
rect 828 -3128 829 -3127
rect 1206 -3128 1207 -3127
rect 1248 -3128 1249 -3127
rect 1269 -3128 1270 -3127
rect 1276 -3128 1277 -3127
rect 1881 -3128 1882 -3127
rect 121 -3130 122 -3129
rect 156 -3130 157 -3129
rect 191 -3130 192 -3129
rect 226 -3130 227 -3129
rect 275 -3130 276 -3129
rect 401 -3130 402 -3129
rect 404 -3130 405 -3129
rect 457 -3130 458 -3129
rect 471 -3130 472 -3129
rect 604 -3130 605 -3129
rect 625 -3130 626 -3129
rect 1083 -3130 1084 -3129
rect 1094 -3130 1095 -3129
rect 1125 -3130 1126 -3129
rect 1185 -3130 1186 -3129
rect 1269 -3130 1270 -3129
rect 1297 -3130 1298 -3129
rect 1314 -3130 1315 -3129
rect 1318 -3130 1319 -3129
rect 1640 -3130 1641 -3129
rect 1647 -3130 1648 -3129
rect 1955 -3130 1956 -3129
rect 135 -3132 136 -3131
rect 275 -3132 276 -3131
rect 296 -3132 297 -3131
rect 373 -3132 374 -3131
rect 471 -3132 472 -3131
rect 534 -3132 535 -3131
rect 541 -3132 542 -3131
rect 569 -3132 570 -3131
rect 625 -3132 626 -3131
rect 709 -3132 710 -3131
rect 716 -3132 717 -3131
rect 835 -3132 836 -3131
rect 863 -3132 864 -3131
rect 919 -3132 920 -3131
rect 961 -3132 962 -3131
rect 1703 -3132 1704 -3131
rect 135 -3134 136 -3133
rect 268 -3134 269 -3133
rect 310 -3134 311 -3133
rect 317 -3134 318 -3133
rect 366 -3134 367 -3133
rect 429 -3134 430 -3133
rect 443 -3134 444 -3133
rect 709 -3134 710 -3133
rect 758 -3134 759 -3133
rect 954 -3134 955 -3133
rect 961 -3134 962 -3133
rect 1031 -3134 1032 -3133
rect 1045 -3134 1046 -3133
rect 1710 -3134 1711 -3133
rect 142 -3136 143 -3135
rect 912 -3136 913 -3135
rect 968 -3136 969 -3135
rect 1559 -3136 1560 -3135
rect 1612 -3136 1613 -3135
rect 1822 -3136 1823 -3135
rect 156 -3138 157 -3137
rect 191 -3138 192 -3137
rect 219 -3138 220 -3137
rect 296 -3138 297 -3137
rect 317 -3138 318 -3137
rect 331 -3138 332 -3137
rect 429 -3138 430 -3137
rect 597 -3138 598 -3137
rect 632 -3138 633 -3137
rect 807 -3138 808 -3137
rect 856 -3138 857 -3137
rect 919 -3138 920 -3137
rect 968 -3138 969 -3137
rect 1227 -3138 1228 -3137
rect 1248 -3138 1249 -3137
rect 1367 -3138 1368 -3137
rect 1402 -3138 1403 -3137
rect 1549 -3138 1550 -3137
rect 1556 -3138 1557 -3137
rect 1906 -3138 1907 -3137
rect 173 -3140 174 -3139
rect 1045 -3140 1046 -3139
rect 1073 -3140 1074 -3139
rect 1304 -3140 1305 -3139
rect 1318 -3140 1319 -3139
rect 1717 -3140 1718 -3139
rect 1766 -3140 1767 -3139
rect 1822 -3140 1823 -3139
rect 1906 -3140 1907 -3139
rect 1934 -3140 1935 -3139
rect 205 -3142 206 -3141
rect 632 -3142 633 -3141
rect 639 -3142 640 -3141
rect 866 -3142 867 -3141
rect 912 -3142 913 -3141
rect 1374 -3142 1375 -3141
rect 1409 -3142 1410 -3141
rect 1542 -3142 1543 -3141
rect 1549 -3142 1550 -3141
rect 1626 -3142 1627 -3141
rect 1661 -3142 1662 -3141
rect 1766 -3142 1767 -3141
rect 219 -3144 220 -3143
rect 261 -3144 262 -3143
rect 268 -3144 269 -3143
rect 345 -3144 346 -3143
rect 394 -3144 395 -3143
rect 639 -3144 640 -3143
rect 681 -3144 682 -3143
rect 702 -3144 703 -3143
rect 765 -3144 766 -3143
rect 1031 -3144 1032 -3143
rect 1073 -3144 1074 -3143
rect 1171 -3144 1172 -3143
rect 1185 -3144 1186 -3143
rect 1360 -3144 1361 -3143
rect 1367 -3144 1368 -3143
rect 1577 -3144 1578 -3143
rect 1626 -3144 1627 -3143
rect 1927 -3144 1928 -3143
rect 261 -3146 262 -3145
rect 1157 -3146 1158 -3145
rect 1171 -3146 1172 -3145
rect 1458 -3146 1459 -3145
rect 1472 -3146 1473 -3145
rect 1668 -3146 1669 -3145
rect 1675 -3146 1676 -3145
rect 1850 -3146 1851 -3145
rect 331 -3148 332 -3147
rect 583 -3148 584 -3147
rect 597 -3148 598 -3147
rect 618 -3148 619 -3147
rect 688 -3148 689 -3147
rect 793 -3148 794 -3147
rect 800 -3148 801 -3147
rect 856 -3148 857 -3147
rect 1017 -3148 1018 -3147
rect 1052 -3148 1053 -3147
rect 1076 -3148 1077 -3147
rect 1657 -3148 1658 -3147
rect 1661 -3148 1662 -3147
rect 1843 -3148 1844 -3147
rect 338 -3150 339 -3149
rect 345 -3150 346 -3149
rect 394 -3150 395 -3149
rect 660 -3150 661 -3149
rect 702 -3150 703 -3149
rect 1024 -3150 1025 -3149
rect 1094 -3150 1095 -3149
rect 1220 -3150 1221 -3149
rect 1227 -3150 1228 -3149
rect 1332 -3150 1333 -3149
rect 1360 -3150 1361 -3149
rect 1507 -3150 1508 -3149
rect 1535 -3150 1536 -3149
rect 1591 -3150 1592 -3149
rect 338 -3152 339 -3151
rect 450 -3152 451 -3151
rect 485 -3152 486 -3151
rect 541 -3152 542 -3151
rect 576 -3152 577 -3151
rect 716 -3152 717 -3151
rect 768 -3152 769 -3151
rect 1192 -3152 1193 -3151
rect 1206 -3152 1207 -3151
rect 1216 -3152 1217 -3151
rect 1220 -3152 1221 -3151
rect 1241 -3152 1242 -3151
rect 1262 -3152 1263 -3151
rect 1444 -3152 1445 -3151
rect 1486 -3152 1487 -3151
rect 1654 -3152 1655 -3151
rect 37 -3154 38 -3153
rect 576 -3154 577 -3153
rect 583 -3154 584 -3153
rect 1055 -3154 1056 -3153
rect 1101 -3154 1102 -3153
rect 1213 -3154 1214 -3153
rect 1241 -3154 1242 -3153
rect 1416 -3154 1417 -3153
rect 1437 -3154 1438 -3153
rect 1685 -3154 1686 -3153
rect 418 -3156 419 -3155
rect 450 -3156 451 -3155
rect 485 -3156 486 -3155
rect 723 -3156 724 -3155
rect 793 -3156 794 -3155
rect 842 -3156 843 -3155
rect 985 -3156 986 -3155
rect 1507 -3156 1508 -3155
rect 1542 -3156 1543 -3155
rect 1815 -3156 1816 -3155
rect 443 -3158 444 -3157
rect 1213 -3158 1214 -3157
rect 1262 -3158 1263 -3157
rect 1493 -3158 1494 -3157
rect 1570 -3158 1571 -3157
rect 1717 -3158 1718 -3157
rect 1738 -3158 1739 -3157
rect 1815 -3158 1816 -3157
rect 506 -3160 507 -3159
rect 933 -3160 934 -3159
rect 989 -3160 990 -3159
rect 1192 -3160 1193 -3159
rect 1297 -3160 1298 -3159
rect 1965 -3160 1966 -3159
rect 520 -3162 521 -3161
rect 1398 -3162 1399 -3161
rect 1416 -3162 1417 -3161
rect 1584 -3162 1585 -3161
rect 1591 -3162 1592 -3161
rect 1801 -3162 1802 -3161
rect 1965 -3162 1966 -3161
rect 2032 -3162 2033 -3161
rect 527 -3164 528 -3163
rect 884 -3164 885 -3163
rect 905 -3164 906 -3163
rect 989 -3164 990 -3163
rect 1003 -3164 1004 -3163
rect 1017 -3164 1018 -3163
rect 1024 -3164 1025 -3163
rect 1059 -3164 1060 -3163
rect 1101 -3164 1102 -3163
rect 1136 -3164 1137 -3163
rect 1157 -3164 1158 -3163
rect 1290 -3164 1291 -3163
rect 1325 -3164 1326 -3163
rect 1514 -3164 1515 -3163
rect 1521 -3164 1522 -3163
rect 1738 -3164 1739 -3163
rect 324 -3166 325 -3165
rect 1290 -3166 1291 -3165
rect 1332 -3166 1333 -3165
rect 1479 -3166 1480 -3165
rect 1493 -3166 1494 -3165
rect 1689 -3166 1690 -3165
rect 324 -3168 325 -3167
rect 387 -3168 388 -3167
rect 527 -3168 528 -3167
rect 744 -3168 745 -3167
rect 786 -3168 787 -3167
rect 884 -3168 885 -3167
rect 905 -3168 906 -3167
rect 975 -3168 976 -3167
rect 1003 -3168 1004 -3167
rect 1066 -3168 1067 -3167
rect 1143 -3168 1144 -3167
rect 1479 -3168 1480 -3167
rect 1500 -3168 1501 -3167
rect 1570 -3168 1571 -3167
rect 1577 -3168 1578 -3167
rect 1941 -3168 1942 -3167
rect 387 -3170 388 -3169
rect 513 -3170 514 -3169
rect 534 -3170 535 -3169
rect 772 -3170 773 -3169
rect 800 -3170 801 -3169
rect 1689 -3170 1690 -3169
rect 464 -3172 465 -3171
rect 744 -3172 745 -3171
rect 814 -3172 815 -3171
rect 1374 -3172 1375 -3171
rect 1500 -3172 1501 -3171
rect 1598 -3172 1599 -3171
rect 1650 -3172 1651 -3171
rect 1685 -3172 1686 -3171
rect 163 -3174 164 -3173
rect 464 -3174 465 -3173
rect 492 -3174 493 -3173
rect 975 -3174 976 -3173
rect 1059 -3174 1060 -3173
rect 1150 -3174 1151 -3173
rect 1356 -3174 1357 -3173
rect 1521 -3174 1522 -3173
rect 1584 -3174 1585 -3173
rect 1731 -3174 1732 -3173
rect 163 -3176 164 -3175
rect 765 -3176 766 -3175
rect 933 -3176 934 -3175
rect 982 -3176 983 -3175
rect 1066 -3176 1067 -3175
rect 1108 -3176 1109 -3175
rect 1143 -3176 1144 -3175
rect 1178 -3176 1179 -3175
rect 1514 -3176 1515 -3175
rect 1696 -3176 1697 -3175
rect 1731 -3176 1732 -3175
rect 1745 -3176 1746 -3175
rect 415 -3178 416 -3177
rect 492 -3178 493 -3177
rect 513 -3178 514 -3177
rect 590 -3178 591 -3177
rect 611 -3178 612 -3177
rect 786 -3178 787 -3177
rect 940 -3178 941 -3177
rect 1136 -3178 1137 -3177
rect 1150 -3178 1151 -3177
rect 1283 -3178 1284 -3177
rect 1598 -3178 1599 -3177
rect 1836 -3178 1837 -3177
rect 415 -3180 416 -3179
rect 898 -3180 899 -3179
rect 954 -3180 955 -3179
rect 1178 -3180 1179 -3179
rect 1283 -3180 1284 -3179
rect 1339 -3180 1340 -3179
rect 1654 -3180 1655 -3179
rect 1969 -3180 1970 -3179
rect 184 -3182 185 -3181
rect 1339 -3182 1340 -3181
rect 1696 -3182 1697 -3181
rect 1808 -3182 1809 -3181
rect 1969 -3182 1970 -3181
rect 1983 -3182 1984 -3181
rect 590 -3184 591 -3183
rect 695 -3184 696 -3183
rect 730 -3184 731 -3183
rect 814 -3184 815 -3183
rect 1108 -3184 1109 -3183
rect 1353 -3184 1354 -3183
rect 1745 -3184 1746 -3183
rect 1759 -3184 1760 -3183
rect 1780 -3184 1781 -3183
rect 1808 -3184 1809 -3183
rect 1983 -3184 1984 -3183
rect 1990 -3184 1991 -3183
rect 82 -3186 83 -3185
rect 730 -3186 731 -3185
rect 772 -3186 773 -3185
rect 1353 -3186 1354 -3185
rect 1752 -3186 1753 -3185
rect 1759 -3186 1760 -3185
rect 1773 -3186 1774 -3185
rect 1780 -3186 1781 -3185
rect 562 -3188 563 -3187
rect 695 -3188 696 -3187
rect 1752 -3188 1753 -3187
rect 1794 -3188 1795 -3187
rect 499 -3190 500 -3189
rect 562 -3190 563 -3189
rect 611 -3190 612 -3189
rect 667 -3190 668 -3189
rect 674 -3190 675 -3189
rect 723 -3190 724 -3189
rect 1773 -3190 1774 -3189
rect 1829 -3190 1830 -3189
rect 499 -3192 500 -3191
rect 779 -3192 780 -3191
rect 614 -3194 615 -3193
rect 940 -3194 941 -3193
rect 247 -3196 248 -3195
rect 614 -3196 615 -3195
rect 618 -3196 619 -3195
rect 646 -3196 647 -3195
rect 653 -3196 654 -3195
rect 842 -3196 843 -3195
rect 240 -3198 241 -3197
rect 247 -3198 248 -3197
rect 478 -3198 479 -3197
rect 653 -3198 654 -3197
rect 660 -3198 661 -3197
rect 1080 -3198 1081 -3197
rect 170 -3200 171 -3199
rect 240 -3200 241 -3199
rect 408 -3200 409 -3199
rect 478 -3200 479 -3199
rect 548 -3200 549 -3199
rect 646 -3200 647 -3199
rect 667 -3200 668 -3199
rect 870 -3200 871 -3199
rect 170 -3202 171 -3201
rect 751 -3202 752 -3201
rect 779 -3202 780 -3201
rect 947 -3202 948 -3201
rect 128 -3204 129 -3203
rect 751 -3204 752 -3203
rect 849 -3204 850 -3203
rect 1080 -3204 1081 -3203
rect 128 -3206 129 -3205
rect 149 -3206 150 -3205
rect 408 -3206 409 -3205
rect 422 -3206 423 -3205
rect 548 -3206 549 -3205
rect 747 -3206 748 -3205
rect 849 -3206 850 -3205
rect 1038 -3206 1039 -3205
rect 149 -3208 150 -3207
rect 460 -3208 461 -3207
rect 947 -3208 948 -3207
rect 996 -3208 997 -3207
rect 1038 -3208 1039 -3207
rect 1087 -3208 1088 -3207
rect 996 -3210 997 -3209
rect 1010 -3210 1011 -3209
rect 1087 -3210 1088 -3209
rect 1255 -3210 1256 -3209
rect 1010 -3212 1011 -3211
rect 1458 -3212 1459 -3211
rect 1255 -3214 1256 -3213
rect 1423 -3214 1424 -3213
rect 1164 -3216 1165 -3215
rect 1423 -3216 1424 -3215
rect 1164 -3218 1165 -3217
rect 1528 -3218 1529 -3217
rect 1430 -3220 1431 -3219
rect 1528 -3220 1529 -3219
rect 1430 -3222 1431 -3221
rect 1619 -3222 1620 -3221
rect 1619 -3224 1620 -3223
rect 1913 -3224 1914 -3223
rect 93 -3235 94 -3234
rect 173 -3235 174 -3234
rect 184 -3235 185 -3234
rect 537 -3235 538 -3234
rect 548 -3235 549 -3234
rect 600 -3235 601 -3234
rect 642 -3235 643 -3234
rect 772 -3235 773 -3234
rect 800 -3235 801 -3234
rect 1444 -3235 1445 -3234
rect 1563 -3235 1564 -3234
rect 1643 -3235 1644 -3234
rect 1668 -3235 1669 -3234
rect 1727 -3235 1728 -3234
rect 1738 -3235 1739 -3234
rect 1965 -3235 1966 -3234
rect 2018 -3235 2019 -3234
rect 2025 -3235 2026 -3234
rect 2032 -3235 2033 -3234
rect 2046 -3235 2047 -3234
rect 107 -3237 108 -3236
rect 677 -3237 678 -3236
rect 688 -3237 689 -3236
rect 1164 -3237 1165 -3236
rect 1213 -3237 1214 -3236
rect 1598 -3237 1599 -3236
rect 1640 -3237 1641 -3236
rect 1745 -3237 1746 -3236
rect 1766 -3237 1767 -3236
rect 1787 -3237 1788 -3236
rect 1808 -3237 1809 -3236
rect 1850 -3237 1851 -3236
rect 1871 -3237 1872 -3236
rect 1885 -3237 1886 -3236
rect 1962 -3237 1963 -3236
rect 1983 -3237 1984 -3236
rect 121 -3239 122 -3238
rect 205 -3239 206 -3238
rect 208 -3239 209 -3238
rect 226 -3239 227 -3238
rect 233 -3239 234 -3238
rect 257 -3239 258 -3238
rect 275 -3239 276 -3238
rect 782 -3239 783 -3238
rect 800 -3239 801 -3238
rect 898 -3239 899 -3238
rect 929 -3239 930 -3238
rect 1605 -3239 1606 -3238
rect 1689 -3239 1690 -3238
rect 1794 -3239 1795 -3238
rect 1815 -3239 1816 -3238
rect 1843 -3239 1844 -3238
rect 1962 -3239 1963 -3238
rect 1976 -3239 1977 -3238
rect 100 -3241 101 -3240
rect 226 -3241 227 -3240
rect 247 -3241 248 -3240
rect 275 -3241 276 -3240
rect 282 -3241 283 -3240
rect 415 -3241 416 -3240
rect 464 -3241 465 -3240
rect 870 -3241 871 -3240
rect 873 -3241 874 -3240
rect 1465 -3241 1466 -3240
rect 1528 -3241 1529 -3240
rect 1605 -3241 1606 -3240
rect 1703 -3241 1704 -3240
rect 1801 -3241 1802 -3240
rect 1815 -3241 1816 -3240
rect 1850 -3241 1851 -3240
rect 128 -3243 129 -3242
rect 187 -3243 188 -3242
rect 191 -3243 192 -3242
rect 1584 -3243 1585 -3242
rect 1598 -3243 1599 -3242
rect 1633 -3243 1634 -3242
rect 1717 -3243 1718 -3242
rect 1738 -3243 1739 -3242
rect 1745 -3243 1746 -3242
rect 1773 -3243 1774 -3242
rect 1822 -3243 1823 -3242
rect 1836 -3243 1837 -3242
rect 135 -3245 136 -3244
rect 719 -3245 720 -3244
rect 751 -3245 752 -3244
rect 943 -3245 944 -3244
rect 957 -3245 958 -3244
rect 996 -3245 997 -3244
rect 1104 -3245 1105 -3244
rect 1220 -3245 1221 -3244
rect 1237 -3245 1238 -3244
rect 1619 -3245 1620 -3244
rect 1717 -3245 1718 -3244
rect 1731 -3245 1732 -3244
rect 1759 -3245 1760 -3244
rect 1766 -3245 1767 -3244
rect 156 -3247 157 -3246
rect 170 -3247 171 -3246
rect 191 -3247 192 -3246
rect 1647 -3247 1648 -3246
rect 1731 -3247 1732 -3246
rect 1752 -3247 1753 -3246
rect 205 -3249 206 -3248
rect 212 -3249 213 -3248
rect 215 -3249 216 -3248
rect 1069 -3249 1070 -3248
rect 1108 -3249 1109 -3248
rect 1682 -3249 1683 -3248
rect 1724 -3249 1725 -3248
rect 1752 -3249 1753 -3248
rect 219 -3251 220 -3250
rect 803 -3251 804 -3250
rect 814 -3251 815 -3250
rect 1010 -3251 1011 -3250
rect 1108 -3251 1109 -3250
rect 1129 -3251 1130 -3250
rect 1216 -3251 1217 -3250
rect 1409 -3251 1410 -3250
rect 1465 -3251 1466 -3250
rect 1654 -3251 1655 -3250
rect 219 -3253 220 -3252
rect 415 -3253 416 -3252
rect 464 -3253 465 -3252
rect 506 -3253 507 -3252
rect 513 -3253 514 -3252
rect 614 -3253 615 -3252
rect 632 -3253 633 -3252
rect 1129 -3253 1130 -3252
rect 1216 -3253 1217 -3252
rect 1346 -3253 1347 -3252
rect 1353 -3253 1354 -3252
rect 1591 -3253 1592 -3252
rect 1654 -3253 1655 -3252
rect 1696 -3253 1697 -3252
rect 240 -3255 241 -3254
rect 506 -3255 507 -3254
rect 576 -3255 577 -3254
rect 1650 -3255 1651 -3254
rect 240 -3257 241 -3256
rect 639 -3257 640 -3256
rect 653 -3257 654 -3256
rect 688 -3257 689 -3256
rect 716 -3257 717 -3256
rect 1332 -3257 1333 -3256
rect 1346 -3257 1347 -3256
rect 1486 -3257 1487 -3256
rect 1549 -3257 1550 -3256
rect 1591 -3257 1592 -3256
rect 247 -3259 248 -3258
rect 261 -3259 262 -3258
rect 282 -3259 283 -3258
rect 660 -3259 661 -3258
rect 674 -3259 675 -3258
rect 702 -3259 703 -3258
rect 716 -3259 717 -3258
rect 992 -3259 993 -3258
rect 1080 -3259 1081 -3258
rect 1353 -3259 1354 -3258
rect 1374 -3259 1375 -3258
rect 1444 -3259 1445 -3258
rect 1472 -3259 1473 -3258
rect 1528 -3259 1529 -3258
rect 1563 -3259 1564 -3258
rect 1661 -3259 1662 -3258
rect 254 -3261 255 -3260
rect 261 -3261 262 -3260
rect 331 -3261 332 -3260
rect 744 -3261 745 -3260
rect 751 -3261 752 -3260
rect 807 -3261 808 -3260
rect 856 -3261 857 -3260
rect 982 -3261 983 -3260
rect 985 -3261 986 -3260
rect 1269 -3261 1270 -3260
rect 1290 -3261 1291 -3260
rect 1458 -3261 1459 -3260
rect 1486 -3261 1487 -3260
rect 1580 -3261 1581 -3260
rect 1661 -3261 1662 -3260
rect 1675 -3261 1676 -3260
rect 268 -3263 269 -3262
rect 331 -3263 332 -3262
rect 338 -3263 339 -3262
rect 726 -3263 727 -3262
rect 772 -3263 773 -3262
rect 793 -3263 794 -3262
rect 807 -3263 808 -3262
rect 947 -3263 948 -3262
rect 957 -3263 958 -3262
rect 1164 -3263 1165 -3262
rect 1167 -3263 1168 -3262
rect 1472 -3263 1473 -3262
rect 268 -3265 269 -3264
rect 289 -3265 290 -3264
rect 338 -3265 339 -3264
rect 604 -3265 605 -3264
rect 653 -3265 654 -3264
rect 695 -3265 696 -3264
rect 702 -3265 703 -3264
rect 1255 -3265 1256 -3264
rect 1269 -3265 1270 -3264
rect 1612 -3265 1613 -3264
rect 289 -3267 290 -3266
rect 345 -3267 346 -3266
rect 352 -3267 353 -3266
rect 418 -3267 419 -3266
rect 485 -3267 486 -3266
rect 513 -3267 514 -3266
rect 562 -3267 563 -3266
rect 856 -3267 857 -3266
rect 863 -3267 864 -3266
rect 870 -3267 871 -3266
rect 898 -3267 899 -3266
rect 1094 -3267 1095 -3266
rect 1115 -3267 1116 -3266
rect 1234 -3267 1235 -3266
rect 1237 -3267 1238 -3266
rect 1685 -3267 1686 -3266
rect 345 -3269 346 -3268
rect 646 -3269 647 -3268
rect 660 -3269 661 -3268
rect 667 -3269 668 -3268
rect 695 -3269 696 -3268
rect 730 -3269 731 -3268
rect 793 -3269 794 -3268
rect 1031 -3269 1032 -3268
rect 1115 -3269 1116 -3268
rect 1192 -3269 1193 -3268
rect 1220 -3269 1221 -3268
rect 1493 -3269 1494 -3268
rect 352 -3271 353 -3270
rect 443 -3271 444 -3270
rect 485 -3271 486 -3270
rect 786 -3271 787 -3270
rect 912 -3271 913 -3270
rect 1010 -3271 1011 -3270
rect 1031 -3271 1032 -3270
rect 1150 -3271 1151 -3270
rect 1171 -3271 1172 -3270
rect 1255 -3271 1256 -3270
rect 1290 -3271 1291 -3270
rect 1311 -3271 1312 -3270
rect 1332 -3271 1333 -3270
rect 1339 -3271 1340 -3270
rect 1374 -3271 1375 -3270
rect 1514 -3271 1515 -3270
rect 229 -3273 230 -3272
rect 443 -3273 444 -3272
rect 495 -3273 496 -3272
rect 579 -3273 580 -3272
rect 583 -3273 584 -3272
rect 639 -3273 640 -3272
rect 646 -3273 647 -3272
rect 681 -3273 682 -3272
rect 786 -3273 787 -3272
rect 1059 -3273 1060 -3272
rect 1066 -3273 1067 -3272
rect 1493 -3273 1494 -3272
rect 1500 -3273 1501 -3272
rect 1514 -3273 1515 -3272
rect 359 -3275 360 -3274
rect 422 -3275 423 -3274
rect 499 -3275 500 -3274
rect 733 -3275 734 -3274
rect 912 -3275 913 -3274
rect 933 -3275 934 -3274
rect 947 -3275 948 -3274
rect 1003 -3275 1004 -3274
rect 1059 -3275 1060 -3274
rect 1178 -3275 1179 -3274
rect 1192 -3275 1193 -3274
rect 1262 -3275 1263 -3274
rect 1283 -3275 1284 -3274
rect 1500 -3275 1501 -3274
rect 177 -3277 178 -3276
rect 499 -3277 500 -3276
rect 527 -3277 528 -3276
rect 681 -3277 682 -3276
rect 709 -3277 710 -3276
rect 1003 -3277 1004 -3276
rect 1066 -3277 1067 -3276
rect 1227 -3277 1228 -3276
rect 1262 -3277 1263 -3276
rect 1556 -3277 1557 -3276
rect 177 -3279 178 -3278
rect 198 -3279 199 -3278
rect 359 -3279 360 -3278
rect 436 -3279 437 -3278
rect 527 -3279 528 -3278
rect 817 -3279 818 -3278
rect 919 -3279 920 -3278
rect 933 -3279 934 -3278
rect 968 -3279 969 -3278
rect 996 -3279 997 -3278
rect 1150 -3279 1151 -3278
rect 1297 -3279 1298 -3278
rect 1311 -3279 1312 -3278
rect 1318 -3279 1319 -3278
rect 1409 -3279 1410 -3278
rect 1853 -3279 1854 -3278
rect 163 -3281 164 -3280
rect 198 -3281 199 -3280
rect 366 -3281 367 -3280
rect 422 -3281 423 -3280
rect 555 -3281 556 -3280
rect 1339 -3281 1340 -3280
rect 1458 -3281 1459 -3280
rect 1542 -3281 1543 -3280
rect 1853 -3281 1854 -3280
rect 1864 -3281 1865 -3280
rect 142 -3283 143 -3282
rect 163 -3283 164 -3282
rect 324 -3283 325 -3282
rect 366 -3283 367 -3282
rect 373 -3283 374 -3282
rect 436 -3283 437 -3282
rect 478 -3283 479 -3282
rect 555 -3283 556 -3282
rect 562 -3283 563 -3282
rect 597 -3283 598 -3282
rect 604 -3283 605 -3282
rect 737 -3283 738 -3282
rect 919 -3283 920 -3282
rect 954 -3283 955 -3282
rect 968 -3283 969 -3282
rect 1122 -3283 1123 -3282
rect 1157 -3283 1158 -3282
rect 1227 -3283 1228 -3282
rect 1283 -3283 1284 -3282
rect 1381 -3283 1382 -3282
rect 1535 -3283 1536 -3282
rect 1556 -3283 1557 -3282
rect 1864 -3283 1865 -3282
rect 1892 -3283 1893 -3282
rect 117 -3285 118 -3284
rect 142 -3285 143 -3284
rect 310 -3285 311 -3284
rect 597 -3285 598 -3284
rect 667 -3285 668 -3284
rect 779 -3285 780 -3284
rect 1122 -3285 1123 -3284
rect 1206 -3285 1207 -3284
rect 1297 -3285 1298 -3284
rect 1367 -3285 1368 -3284
rect 1892 -3285 1893 -3284
rect 1906 -3285 1907 -3284
rect 310 -3287 311 -3286
rect 317 -3287 318 -3286
rect 324 -3287 325 -3286
rect 429 -3287 430 -3286
rect 576 -3287 577 -3286
rect 940 -3287 941 -3286
rect 1143 -3287 1144 -3286
rect 1157 -3287 1158 -3286
rect 1171 -3287 1172 -3286
rect 1388 -3287 1389 -3286
rect 1906 -3287 1907 -3286
rect 1920 -3287 1921 -3286
rect 317 -3289 318 -3288
rect 625 -3289 626 -3288
rect 709 -3289 710 -3288
rect 835 -3289 836 -3288
rect 940 -3289 941 -3288
rect 1024 -3289 1025 -3288
rect 1178 -3289 1179 -3288
rect 1416 -3289 1417 -3288
rect 373 -3291 374 -3290
rect 450 -3291 451 -3290
rect 583 -3291 584 -3290
rect 611 -3291 612 -3290
rect 625 -3291 626 -3290
rect 1094 -3291 1095 -3290
rect 1206 -3291 1207 -3290
rect 1437 -3291 1438 -3290
rect 149 -3293 150 -3292
rect 611 -3293 612 -3292
rect 737 -3293 738 -3292
rect 1017 -3293 1018 -3292
rect 1024 -3293 1025 -3292
rect 1052 -3293 1053 -3292
rect 1318 -3293 1319 -3292
rect 1430 -3293 1431 -3292
rect 383 -3295 384 -3294
rect 863 -3295 864 -3294
rect 961 -3295 962 -3294
rect 1388 -3295 1389 -3294
rect 1402 -3295 1403 -3294
rect 1437 -3295 1438 -3294
rect 387 -3297 388 -3296
rect 492 -3297 493 -3296
rect 590 -3297 591 -3296
rect 632 -3297 633 -3296
rect 765 -3297 766 -3296
rect 1017 -3297 1018 -3296
rect 1038 -3297 1039 -3296
rect 1052 -3297 1053 -3296
rect 1136 -3297 1137 -3296
rect 1402 -3297 1403 -3296
rect 387 -3299 388 -3298
rect 471 -3299 472 -3298
rect 590 -3299 591 -3298
rect 1087 -3299 1088 -3298
rect 1136 -3299 1137 -3298
rect 1199 -3299 1200 -3298
rect 1325 -3299 1326 -3298
rect 1430 -3299 1431 -3298
rect 394 -3301 395 -3300
rect 548 -3301 549 -3300
rect 765 -3301 766 -3300
rect 905 -3301 906 -3300
rect 961 -3301 962 -3300
rect 989 -3301 990 -3300
rect 1038 -3301 1039 -3300
rect 1080 -3301 1081 -3300
rect 1087 -3301 1088 -3300
rect 1185 -3301 1186 -3300
rect 1199 -3301 1200 -3300
rect 1360 -3301 1361 -3300
rect 1367 -3301 1368 -3300
rect 1570 -3301 1571 -3300
rect 394 -3303 395 -3302
rect 408 -3303 409 -3302
rect 429 -3303 430 -3302
rect 534 -3303 535 -3302
rect 723 -3303 724 -3302
rect 1185 -3303 1186 -3302
rect 1325 -3303 1326 -3302
rect 1521 -3303 1522 -3302
rect 380 -3305 381 -3304
rect 408 -3305 409 -3304
rect 450 -3305 451 -3304
rect 618 -3305 619 -3304
rect 779 -3305 780 -3304
rect 1276 -3305 1277 -3304
rect 1451 -3305 1452 -3304
rect 1521 -3305 1522 -3304
rect 380 -3307 381 -3306
rect 478 -3307 479 -3306
rect 534 -3307 535 -3306
rect 1671 -3307 1672 -3306
rect 401 -3309 402 -3308
rect 618 -3309 619 -3308
rect 821 -3309 822 -3308
rect 835 -3309 836 -3308
rect 884 -3309 885 -3308
rect 1360 -3309 1361 -3308
rect 1451 -3309 1452 -3308
rect 1507 -3309 1508 -3308
rect 296 -3311 297 -3310
rect 401 -3311 402 -3310
rect 404 -3311 405 -3310
rect 457 -3311 458 -3310
rect 471 -3311 472 -3310
rect 975 -3311 976 -3310
rect 978 -3311 979 -3310
rect 1143 -3311 1144 -3310
rect 1248 -3311 1249 -3310
rect 1276 -3311 1277 -3310
rect 1423 -3311 1424 -3310
rect 1507 -3311 1508 -3310
rect 296 -3313 297 -3312
rect 768 -3313 769 -3312
rect 821 -3313 822 -3312
rect 842 -3313 843 -3312
rect 849 -3313 850 -3312
rect 884 -3313 885 -3312
rect 905 -3313 906 -3312
rect 1234 -3313 1235 -3312
rect 1248 -3313 1249 -3312
rect 1479 -3313 1480 -3312
rect 457 -3315 458 -3314
rect 520 -3315 521 -3314
rect 842 -3315 843 -3314
rect 877 -3315 878 -3314
rect 989 -3315 990 -3314
rect 1626 -3315 1627 -3314
rect 520 -3317 521 -3316
rect 758 -3317 759 -3316
rect 877 -3317 878 -3316
rect 891 -3317 892 -3316
rect 1304 -3317 1305 -3316
rect 1423 -3317 1424 -3316
rect 1479 -3317 1480 -3316
rect 1724 -3317 1725 -3316
rect 758 -3319 759 -3318
rect 849 -3319 850 -3318
rect 1304 -3319 1305 -3318
rect 1395 -3319 1396 -3318
rect 1626 -3319 1627 -3318
rect 1710 -3319 1711 -3318
rect 828 -3321 829 -3320
rect 891 -3321 892 -3320
rect 1073 -3321 1074 -3320
rect 1395 -3321 1396 -3320
rect 828 -3323 829 -3322
rect 926 -3323 927 -3322
rect 1073 -3323 1074 -3322
rect 1241 -3323 1242 -3322
rect 254 -3325 255 -3324
rect 926 -3325 927 -3324
rect 1045 -3325 1046 -3324
rect 1241 -3325 1242 -3324
rect 1045 -3327 1046 -3326
rect 1101 -3327 1102 -3326
rect 142 -3338 143 -3337
rect 173 -3338 174 -3337
rect 177 -3338 178 -3337
rect 236 -3338 237 -3337
rect 257 -3338 258 -3337
rect 373 -3338 374 -3337
rect 394 -3338 395 -3337
rect 537 -3338 538 -3337
rect 541 -3338 542 -3337
rect 544 -3338 545 -3337
rect 590 -3338 591 -3337
rect 779 -3338 780 -3337
rect 814 -3338 815 -3337
rect 1125 -3338 1126 -3337
rect 1160 -3338 1161 -3337
rect 1227 -3338 1228 -3337
rect 1234 -3338 1235 -3337
rect 1451 -3338 1452 -3337
rect 1521 -3338 1522 -3337
rect 1584 -3338 1585 -3337
rect 1591 -3338 1592 -3337
rect 1612 -3338 1613 -3337
rect 1647 -3338 1648 -3337
rect 1661 -3338 1662 -3337
rect 1717 -3338 1718 -3337
rect 1727 -3338 1728 -3337
rect 1752 -3338 1753 -3337
rect 1759 -3338 1760 -3337
rect 1766 -3338 1767 -3337
rect 1769 -3338 1770 -3337
rect 1787 -3338 1788 -3337
rect 1811 -3338 1812 -3337
rect 1829 -3338 1830 -3337
rect 1843 -3338 1844 -3337
rect 1885 -3338 1886 -3337
rect 1906 -3338 1907 -3337
rect 1955 -3338 1956 -3337
rect 1962 -3338 1963 -3337
rect 2025 -3338 2026 -3337
rect 2028 -3338 2029 -3337
rect 163 -3340 164 -3339
rect 390 -3340 391 -3339
rect 415 -3340 416 -3339
rect 485 -3340 486 -3339
rect 488 -3340 489 -3339
rect 506 -3340 507 -3339
rect 513 -3340 514 -3339
rect 992 -3340 993 -3339
rect 1034 -3340 1035 -3339
rect 1220 -3340 1221 -3339
rect 1234 -3340 1235 -3339
rect 1283 -3340 1284 -3339
rect 1339 -3340 1340 -3339
rect 1458 -3340 1459 -3339
rect 1521 -3340 1522 -3339
rect 1528 -3340 1529 -3339
rect 1549 -3340 1550 -3339
rect 1626 -3340 1627 -3339
rect 1724 -3340 1725 -3339
rect 1745 -3340 1746 -3339
rect 1787 -3340 1788 -3339
rect 1850 -3340 1851 -3339
rect 1888 -3340 1889 -3339
rect 1892 -3340 1893 -3339
rect 1962 -3340 1963 -3339
rect 1969 -3340 1970 -3339
rect 2025 -3340 2026 -3339
rect 2032 -3340 2033 -3339
rect 170 -3342 171 -3341
rect 180 -3342 181 -3341
rect 212 -3342 213 -3341
rect 408 -3342 409 -3341
rect 429 -3342 430 -3341
rect 926 -3342 927 -3341
rect 968 -3342 969 -3341
rect 1332 -3342 1333 -3341
rect 1367 -3342 1368 -3341
rect 1493 -3342 1494 -3341
rect 1528 -3342 1529 -3341
rect 1563 -3342 1564 -3341
rect 1605 -3342 1606 -3341
rect 1654 -3342 1655 -3341
rect 1794 -3342 1795 -3341
rect 1822 -3342 1823 -3341
rect 1836 -3342 1837 -3341
rect 1843 -3342 1844 -3341
rect 1850 -3342 1851 -3341
rect 1857 -3342 1858 -3341
rect 215 -3344 216 -3343
rect 803 -3344 804 -3343
rect 821 -3344 822 -3343
rect 936 -3344 937 -3343
rect 968 -3344 969 -3343
rect 1003 -3344 1004 -3343
rect 1031 -3344 1032 -3343
rect 1220 -3344 1221 -3343
rect 1237 -3344 1238 -3343
rect 1297 -3344 1298 -3343
rect 1332 -3344 1333 -3343
rect 1374 -3344 1375 -3343
rect 1381 -3344 1382 -3343
rect 1444 -3344 1445 -3343
rect 1451 -3344 1452 -3343
rect 1486 -3344 1487 -3343
rect 1552 -3344 1553 -3343
rect 1598 -3344 1599 -3343
rect 1608 -3344 1609 -3343
rect 1668 -3344 1669 -3343
rect 1801 -3344 1802 -3343
rect 1836 -3344 1837 -3343
rect 1857 -3344 1858 -3343
rect 1871 -3344 1872 -3343
rect 240 -3346 241 -3345
rect 506 -3346 507 -3345
rect 541 -3346 542 -3345
rect 576 -3346 577 -3345
rect 597 -3346 598 -3345
rect 1083 -3346 1084 -3345
rect 1097 -3346 1098 -3345
rect 1311 -3346 1312 -3345
rect 1374 -3346 1375 -3345
rect 1458 -3346 1459 -3345
rect 1556 -3346 1557 -3345
rect 1587 -3346 1588 -3345
rect 1654 -3346 1655 -3345
rect 1853 -3346 1854 -3345
rect 1864 -3346 1865 -3345
rect 1871 -3346 1872 -3345
rect 275 -3348 276 -3347
rect 373 -3348 374 -3347
rect 422 -3348 423 -3347
rect 429 -3348 430 -3347
rect 474 -3348 475 -3347
rect 1370 -3348 1371 -3347
rect 1384 -3348 1385 -3347
rect 1423 -3348 1424 -3347
rect 1801 -3348 1802 -3347
rect 1815 -3348 1816 -3347
rect 1864 -3348 1865 -3347
rect 1878 -3348 1879 -3347
rect 2028 -3348 2029 -3347
rect 2032 -3348 2033 -3347
rect 205 -3350 206 -3349
rect 422 -3350 423 -3349
rect 548 -3350 549 -3349
rect 1031 -3350 1032 -3349
rect 1066 -3350 1067 -3349
rect 1430 -3350 1431 -3349
rect 282 -3352 283 -3351
rect 859 -3352 860 -3351
rect 877 -3352 878 -3351
rect 1003 -3352 1004 -3351
rect 1080 -3352 1081 -3351
rect 1136 -3352 1137 -3351
rect 1199 -3352 1200 -3351
rect 1227 -3352 1228 -3351
rect 1269 -3352 1270 -3351
rect 1353 -3352 1354 -3351
rect 1388 -3352 1389 -3351
rect 1419 -3352 1420 -3351
rect 296 -3354 297 -3353
rect 383 -3354 384 -3353
rect 492 -3354 493 -3353
rect 548 -3354 549 -3353
rect 555 -3354 556 -3353
rect 590 -3354 591 -3353
rect 597 -3354 598 -3353
rect 646 -3354 647 -3353
rect 653 -3354 654 -3353
rect 877 -3354 878 -3353
rect 891 -3354 892 -3353
rect 954 -3354 955 -3353
rect 961 -3354 962 -3353
rect 1080 -3354 1081 -3353
rect 1101 -3354 1102 -3353
rect 1178 -3354 1179 -3353
rect 1199 -3354 1200 -3353
rect 1325 -3354 1326 -3353
rect 1416 -3354 1417 -3353
rect 1437 -3354 1438 -3353
rect 268 -3356 269 -3355
rect 296 -3356 297 -3355
rect 317 -3356 318 -3355
rect 408 -3356 409 -3355
rect 450 -3356 451 -3355
rect 492 -3356 493 -3355
rect 534 -3356 535 -3355
rect 646 -3356 647 -3355
rect 674 -3356 675 -3355
rect 1027 -3356 1028 -3355
rect 1045 -3356 1046 -3355
rect 1178 -3356 1179 -3355
rect 1213 -3356 1214 -3355
rect 1402 -3356 1403 -3355
rect 359 -3358 360 -3357
rect 513 -3358 514 -3357
rect 534 -3358 535 -3357
rect 583 -3358 584 -3357
rect 618 -3358 619 -3357
rect 639 -3358 640 -3357
rect 660 -3358 661 -3357
rect 674 -3358 675 -3357
rect 681 -3358 682 -3357
rect 1066 -3358 1067 -3357
rect 1157 -3358 1158 -3357
rect 1213 -3358 1214 -3357
rect 1269 -3358 1270 -3357
rect 1472 -3358 1473 -3357
rect 303 -3360 304 -3359
rect 359 -3360 360 -3359
rect 366 -3360 367 -3359
rect 394 -3360 395 -3359
rect 478 -3360 479 -3359
rect 555 -3360 556 -3359
rect 562 -3360 563 -3359
rect 681 -3360 682 -3359
rect 723 -3360 724 -3359
rect 1395 -3360 1396 -3359
rect 1472 -3360 1473 -3359
rect 1514 -3360 1515 -3359
rect 331 -3362 332 -3361
rect 478 -3362 479 -3361
rect 562 -3362 563 -3361
rect 726 -3362 727 -3361
rect 730 -3362 731 -3361
rect 1808 -3362 1809 -3361
rect 198 -3364 199 -3363
rect 331 -3364 332 -3363
rect 345 -3364 346 -3363
rect 660 -3364 661 -3363
rect 723 -3364 724 -3363
rect 758 -3364 759 -3363
rect 772 -3364 773 -3363
rect 814 -3364 815 -3363
rect 821 -3364 822 -3363
rect 1059 -3364 1060 -3363
rect 1272 -3364 1273 -3363
rect 1283 -3364 1284 -3363
rect 1290 -3364 1291 -3363
rect 1297 -3364 1298 -3363
rect 289 -3366 290 -3365
rect 345 -3366 346 -3365
rect 387 -3366 388 -3365
rect 450 -3366 451 -3365
rect 583 -3366 584 -3365
rect 667 -3366 668 -3365
rect 737 -3366 738 -3365
rect 961 -3366 962 -3365
rect 978 -3366 979 -3365
rect 1024 -3366 1025 -3365
rect 1045 -3366 1046 -3365
rect 1143 -3366 1144 -3365
rect 1255 -3366 1256 -3365
rect 1290 -3366 1291 -3365
rect 219 -3368 220 -3367
rect 387 -3368 388 -3367
rect 443 -3368 444 -3367
rect 730 -3368 731 -3367
rect 751 -3368 752 -3367
rect 1094 -3368 1095 -3367
rect 1192 -3368 1193 -3367
rect 1255 -3368 1256 -3367
rect 352 -3370 353 -3369
rect 667 -3370 668 -3369
rect 772 -3370 773 -3369
rect 800 -3370 801 -3369
rect 835 -3370 836 -3369
rect 849 -3370 850 -3369
rect 852 -3370 853 -3369
rect 1010 -3370 1011 -3369
rect 1024 -3370 1025 -3369
rect 1038 -3370 1039 -3369
rect 1059 -3370 1060 -3369
rect 1073 -3370 1074 -3369
rect 1094 -3370 1095 -3369
rect 1241 -3370 1242 -3369
rect 401 -3372 402 -3371
rect 443 -3372 444 -3371
rect 471 -3372 472 -3371
rect 737 -3372 738 -3371
rect 779 -3372 780 -3371
rect 975 -3372 976 -3371
rect 982 -3372 983 -3371
rect 1104 -3372 1105 -3371
rect 1192 -3372 1193 -3371
rect 1465 -3372 1466 -3371
rect 401 -3374 402 -3373
rect 751 -3374 752 -3373
rect 793 -3374 794 -3373
rect 835 -3374 836 -3373
rect 842 -3374 843 -3373
rect 957 -3374 958 -3373
rect 989 -3374 990 -3373
rect 1360 -3374 1361 -3373
rect 1465 -3374 1466 -3373
rect 1507 -3374 1508 -3373
rect 600 -3376 601 -3375
rect 1073 -3376 1074 -3375
rect 1241 -3376 1242 -3375
rect 1304 -3376 1305 -3375
rect 1346 -3376 1347 -3375
rect 1360 -3376 1361 -3375
rect 604 -3378 605 -3377
rect 758 -3378 759 -3377
rect 800 -3378 801 -3377
rect 1377 -3378 1378 -3377
rect 604 -3380 605 -3379
rect 611 -3380 612 -3379
rect 618 -3380 619 -3379
rect 709 -3380 710 -3379
rect 842 -3380 843 -3379
rect 1206 -3380 1207 -3379
rect 1318 -3380 1319 -3379
rect 1346 -3380 1347 -3379
rect 520 -3382 521 -3381
rect 709 -3382 710 -3381
rect 849 -3382 850 -3381
rect 1150 -3382 1151 -3381
rect 1185 -3382 1186 -3381
rect 1304 -3382 1305 -3381
rect 418 -3384 419 -3383
rect 520 -3384 521 -3383
rect 527 -3384 528 -3383
rect 611 -3384 612 -3383
rect 625 -3384 626 -3383
rect 653 -3384 654 -3383
rect 688 -3384 689 -3383
rect 793 -3384 794 -3383
rect 856 -3384 857 -3383
rect 982 -3384 983 -3383
rect 989 -3384 990 -3383
rect 1248 -3384 1249 -3383
rect 457 -3386 458 -3385
rect 625 -3386 626 -3385
rect 688 -3386 689 -3385
rect 786 -3386 787 -3385
rect 870 -3386 871 -3385
rect 975 -3386 976 -3385
rect 1108 -3386 1109 -3385
rect 1206 -3386 1207 -3385
rect 1209 -3386 1210 -3385
rect 1248 -3386 1249 -3385
rect 310 -3388 311 -3387
rect 457 -3388 458 -3387
rect 527 -3388 528 -3387
rect 569 -3388 570 -3387
rect 786 -3388 787 -3387
rect 884 -3388 885 -3387
rect 891 -3388 892 -3387
rect 1122 -3388 1123 -3387
rect 1185 -3388 1186 -3387
rect 1479 -3388 1480 -3387
rect 184 -3390 185 -3389
rect 569 -3390 570 -3389
rect 807 -3390 808 -3389
rect 1108 -3390 1109 -3389
rect 1122 -3390 1123 -3389
rect 1381 -3390 1382 -3389
rect 261 -3392 262 -3391
rect 310 -3392 311 -3391
rect 695 -3392 696 -3391
rect 807 -3392 808 -3391
rect 863 -3392 864 -3391
rect 884 -3392 885 -3391
rect 898 -3392 899 -3391
rect 1038 -3392 1039 -3391
rect 324 -3394 325 -3393
rect 695 -3394 696 -3393
rect 744 -3394 745 -3393
rect 863 -3394 864 -3393
rect 870 -3394 871 -3393
rect 905 -3394 906 -3393
rect 919 -3394 920 -3393
rect 1010 -3394 1011 -3393
rect 702 -3396 703 -3395
rect 744 -3396 745 -3395
rect 901 -3396 902 -3395
rect 1276 -3396 1277 -3395
rect 464 -3398 465 -3397
rect 702 -3398 703 -3397
rect 905 -3398 906 -3397
rect 1115 -3398 1116 -3397
rect 436 -3400 437 -3399
rect 464 -3400 465 -3399
rect 912 -3400 913 -3399
rect 919 -3400 920 -3399
rect 926 -3400 927 -3399
rect 1129 -3400 1130 -3399
rect 380 -3402 381 -3401
rect 436 -3402 437 -3401
rect 765 -3402 766 -3401
rect 912 -3402 913 -3401
rect 940 -3402 941 -3401
rect 1143 -3402 1144 -3401
rect 247 -3404 248 -3403
rect 380 -3404 381 -3403
rect 632 -3404 633 -3403
rect 765 -3404 766 -3403
rect 940 -3404 941 -3403
rect 1216 -3404 1217 -3403
rect 499 -3406 500 -3405
rect 632 -3406 633 -3405
rect 947 -3406 948 -3405
rect 1136 -3406 1137 -3405
rect 338 -3408 339 -3407
rect 499 -3408 500 -3407
rect 828 -3408 829 -3407
rect 947 -3408 948 -3407
rect 954 -3408 955 -3407
rect 996 -3408 997 -3407
rect 1052 -3408 1053 -3407
rect 1115 -3408 1116 -3407
rect 191 -3410 192 -3409
rect 338 -3410 339 -3409
rect 828 -3410 829 -3409
rect 933 -3410 934 -3409
rect 996 -3410 997 -3409
rect 1171 -3410 1172 -3409
rect 933 -3412 934 -3411
rect 1017 -3412 1018 -3411
rect 1052 -3412 1053 -3411
rect 1087 -3412 1088 -3411
rect 1171 -3412 1172 -3411
rect 1262 -3412 1263 -3411
rect 971 -3414 972 -3413
rect 1017 -3414 1018 -3413
rect 1087 -3414 1088 -3413
rect 1164 -3414 1165 -3413
rect 1262 -3414 1263 -3413
rect 1409 -3414 1410 -3413
rect 173 -3425 174 -3424
rect 268 -3425 269 -3424
rect 296 -3425 297 -3424
rect 317 -3425 318 -3424
rect 338 -3425 339 -3424
rect 474 -3425 475 -3424
rect 478 -3425 479 -3424
rect 593 -3425 594 -3424
rect 621 -3425 622 -3424
rect 632 -3425 633 -3424
rect 639 -3425 640 -3424
rect 723 -3425 724 -3424
rect 726 -3425 727 -3424
rect 940 -3425 941 -3424
rect 961 -3425 962 -3424
rect 1206 -3425 1207 -3424
rect 1213 -3425 1214 -3424
rect 1286 -3425 1287 -3424
rect 1297 -3425 1298 -3424
rect 1307 -3425 1308 -3424
rect 1311 -3425 1312 -3424
rect 1332 -3425 1333 -3424
rect 1346 -3425 1347 -3424
rect 1374 -3425 1375 -3424
rect 1437 -3425 1438 -3424
rect 1451 -3425 1452 -3424
rect 1458 -3425 1459 -3424
rect 1493 -3425 1494 -3424
rect 1514 -3425 1515 -3424
rect 1528 -3425 1529 -3424
rect 1584 -3425 1585 -3424
rect 1808 -3425 1809 -3424
rect 1822 -3425 1823 -3424
rect 1860 -3425 1861 -3424
rect 170 -3427 171 -3426
rect 173 -3427 174 -3426
rect 310 -3427 311 -3426
rect 324 -3427 325 -3426
rect 345 -3427 346 -3426
rect 390 -3427 391 -3426
rect 394 -3427 395 -3426
rect 401 -3427 402 -3426
rect 404 -3427 405 -3426
rect 415 -3427 416 -3426
rect 429 -3427 430 -3426
rect 467 -3427 468 -3426
rect 492 -3427 493 -3426
rect 628 -3427 629 -3426
rect 646 -3427 647 -3426
rect 723 -3427 724 -3426
rect 758 -3427 759 -3426
rect 800 -3427 801 -3426
rect 807 -3427 808 -3426
rect 842 -3427 843 -3426
rect 884 -3427 885 -3426
rect 922 -3427 923 -3426
rect 975 -3427 976 -3426
rect 1024 -3427 1025 -3426
rect 1066 -3427 1067 -3426
rect 1199 -3427 1200 -3426
rect 1206 -3427 1207 -3426
rect 1234 -3427 1235 -3426
rect 1248 -3427 1249 -3426
rect 1307 -3427 1308 -3426
rect 1321 -3427 1322 -3426
rect 1332 -3427 1333 -3426
rect 1444 -3427 1445 -3426
rect 1465 -3427 1466 -3426
rect 1612 -3427 1613 -3426
rect 1629 -3427 1630 -3426
rect 1640 -3427 1641 -3426
rect 1647 -3427 1648 -3426
rect 1724 -3427 1725 -3426
rect 1727 -3427 1728 -3426
rect 1738 -3427 1739 -3426
rect 1748 -3427 1749 -3426
rect 1759 -3427 1760 -3426
rect 1766 -3427 1767 -3426
rect 1794 -3427 1795 -3426
rect 1801 -3427 1802 -3426
rect 1822 -3427 1823 -3426
rect 1829 -3427 1830 -3426
rect 1857 -3427 1858 -3426
rect 1867 -3427 1868 -3426
rect 373 -3429 374 -3428
rect 471 -3429 472 -3428
rect 492 -3429 493 -3428
rect 562 -3429 563 -3428
rect 611 -3429 612 -3428
rect 639 -3429 640 -3428
rect 653 -3429 654 -3428
rect 656 -3429 657 -3428
rect 684 -3429 685 -3428
rect 716 -3429 717 -3428
rect 744 -3429 745 -3428
rect 758 -3429 759 -3428
rect 807 -3429 808 -3428
rect 989 -3429 990 -3428
rect 992 -3429 993 -3428
rect 1052 -3429 1053 -3428
rect 1066 -3429 1067 -3428
rect 1101 -3429 1102 -3428
rect 1108 -3429 1109 -3428
rect 1199 -3429 1200 -3428
rect 1220 -3429 1221 -3428
rect 1458 -3429 1459 -3428
rect 1461 -3429 1462 -3428
rect 1654 -3429 1655 -3428
rect 1724 -3429 1725 -3428
rect 1731 -3429 1732 -3428
rect 1766 -3429 1767 -3428
rect 1787 -3429 1788 -3428
rect 1829 -3429 1830 -3428
rect 1843 -3429 1844 -3428
rect 1857 -3429 1858 -3428
rect 1864 -3429 1865 -3428
rect 408 -3431 409 -3430
rect 488 -3431 489 -3430
rect 499 -3431 500 -3430
rect 611 -3431 612 -3430
rect 625 -3431 626 -3430
rect 667 -3431 668 -3430
rect 695 -3431 696 -3430
rect 1031 -3431 1032 -3430
rect 1052 -3431 1053 -3430
rect 1087 -3431 1088 -3430
rect 1101 -3431 1102 -3430
rect 1185 -3431 1186 -3430
rect 1255 -3431 1256 -3430
rect 1318 -3431 1319 -3430
rect 1325 -3431 1326 -3430
rect 1367 -3431 1368 -3430
rect 1381 -3431 1382 -3430
rect 1465 -3431 1466 -3430
rect 1836 -3431 1837 -3430
rect 1843 -3431 1844 -3430
rect 1864 -3431 1865 -3430
rect 1871 -3431 1872 -3430
rect 450 -3433 451 -3432
rect 485 -3433 486 -3432
rect 506 -3433 507 -3432
rect 646 -3433 647 -3432
rect 653 -3433 654 -3432
rect 688 -3433 689 -3432
rect 702 -3433 703 -3432
rect 922 -3433 923 -3432
rect 1003 -3433 1004 -3432
rect 1031 -3433 1032 -3432
rect 1069 -3433 1070 -3432
rect 1125 -3433 1126 -3432
rect 1136 -3433 1137 -3432
rect 1220 -3433 1221 -3432
rect 1276 -3433 1277 -3432
rect 1283 -3433 1284 -3432
rect 1451 -3433 1452 -3432
rect 1472 -3433 1473 -3432
rect 422 -3435 423 -3434
rect 506 -3435 507 -3434
rect 548 -3435 549 -3434
rect 579 -3435 580 -3434
rect 660 -3435 661 -3434
rect 695 -3435 696 -3434
rect 702 -3435 703 -3434
rect 786 -3435 787 -3434
rect 814 -3435 815 -3434
rect 845 -3435 846 -3434
rect 863 -3435 864 -3434
rect 884 -3435 885 -3434
rect 901 -3435 902 -3434
rect 1094 -3435 1095 -3434
rect 1108 -3435 1109 -3434
rect 1192 -3435 1193 -3434
rect 1867 -3435 1868 -3434
rect 1871 -3435 1872 -3434
rect 380 -3437 381 -3436
rect 422 -3437 423 -3436
rect 464 -3437 465 -3436
rect 499 -3437 500 -3436
rect 555 -3437 556 -3436
rect 604 -3437 605 -3436
rect 660 -3437 661 -3436
rect 705 -3437 706 -3436
rect 709 -3437 710 -3436
rect 898 -3437 899 -3436
rect 912 -3437 913 -3436
rect 975 -3437 976 -3436
rect 1010 -3437 1011 -3436
rect 1122 -3437 1123 -3436
rect 1143 -3437 1144 -3436
rect 1234 -3437 1235 -3436
rect 331 -3439 332 -3438
rect 464 -3439 465 -3438
rect 541 -3439 542 -3438
rect 555 -3439 556 -3438
rect 558 -3439 559 -3438
rect 779 -3439 780 -3438
rect 814 -3439 815 -3438
rect 828 -3439 829 -3438
rect 835 -3439 836 -3438
rect 859 -3439 860 -3438
rect 915 -3439 916 -3438
rect 968 -3439 969 -3438
rect 982 -3439 983 -3438
rect 1010 -3439 1011 -3438
rect 1034 -3439 1035 -3438
rect 1094 -3439 1095 -3438
rect 1115 -3439 1116 -3438
rect 1181 -3439 1182 -3438
rect 1185 -3439 1186 -3438
rect 1262 -3439 1263 -3438
rect 359 -3441 360 -3440
rect 380 -3441 381 -3440
rect 541 -3441 542 -3440
rect 618 -3441 619 -3440
rect 674 -3441 675 -3440
rect 709 -3441 710 -3440
rect 737 -3441 738 -3440
rect 828 -3441 829 -3440
rect 835 -3441 836 -3440
rect 870 -3441 871 -3440
rect 919 -3441 920 -3440
rect 954 -3441 955 -3440
rect 1073 -3441 1074 -3440
rect 1248 -3441 1249 -3440
rect 562 -3443 563 -3442
rect 597 -3443 598 -3442
rect 604 -3443 605 -3442
rect 625 -3443 626 -3442
rect 681 -3443 682 -3442
rect 737 -3443 738 -3442
rect 744 -3443 745 -3442
rect 821 -3443 822 -3442
rect 842 -3443 843 -3442
rect 891 -3443 892 -3442
rect 947 -3443 948 -3442
rect 1003 -3443 1004 -3442
rect 1059 -3443 1060 -3442
rect 1073 -3443 1074 -3442
rect 1080 -3443 1081 -3442
rect 1129 -3443 1130 -3442
rect 1164 -3443 1165 -3442
rect 1626 -3443 1627 -3442
rect 520 -3445 521 -3444
rect 681 -3445 682 -3444
rect 751 -3445 752 -3444
rect 1125 -3445 1126 -3444
rect 1192 -3445 1193 -3444
rect 1241 -3445 1242 -3444
rect 436 -3447 437 -3446
rect 520 -3447 521 -3446
rect 569 -3447 570 -3446
rect 716 -3447 717 -3446
rect 751 -3447 752 -3446
rect 849 -3447 850 -3446
rect 877 -3447 878 -3446
rect 1080 -3447 1081 -3446
rect 1083 -3447 1084 -3446
rect 1171 -3447 1172 -3446
rect 1227 -3447 1228 -3446
rect 1241 -3447 1242 -3446
rect 527 -3449 528 -3448
rect 569 -3449 570 -3448
rect 583 -3449 584 -3448
rect 597 -3449 598 -3448
rect 632 -3449 633 -3448
rect 1059 -3449 1060 -3448
rect 1087 -3449 1088 -3448
rect 1304 -3449 1305 -3448
rect 513 -3451 514 -3450
rect 583 -3451 584 -3450
rect 590 -3451 591 -3450
rect 674 -3451 675 -3450
rect 730 -3451 731 -3450
rect 849 -3451 850 -3450
rect 877 -3451 878 -3450
rect 905 -3451 906 -3450
rect 954 -3451 955 -3450
rect 996 -3451 997 -3450
rect 1171 -3451 1172 -3450
rect 1269 -3451 1270 -3450
rect 457 -3453 458 -3452
rect 513 -3453 514 -3452
rect 730 -3453 731 -3452
rect 926 -3453 927 -3452
rect 996 -3453 997 -3452
rect 1045 -3453 1046 -3452
rect 1178 -3453 1179 -3452
rect 1227 -3453 1228 -3452
rect 443 -3455 444 -3454
rect 457 -3455 458 -3454
rect 590 -3455 591 -3454
rect 1045 -3455 1046 -3454
rect 1178 -3455 1179 -3454
rect 1213 -3455 1214 -3454
rect 439 -3457 440 -3456
rect 443 -3457 444 -3456
rect 765 -3457 766 -3456
rect 821 -3457 822 -3456
rect 772 -3459 773 -3458
rect 779 -3459 780 -3458
rect 271 -3470 272 -3469
rect 366 -3470 367 -3469
rect 369 -3470 370 -3469
rect 394 -3470 395 -3469
rect 415 -3470 416 -3469
rect 429 -3470 430 -3469
rect 439 -3470 440 -3469
rect 443 -3470 444 -3469
rect 457 -3470 458 -3469
rect 464 -3470 465 -3469
rect 478 -3470 479 -3469
rect 492 -3470 493 -3469
rect 499 -3470 500 -3469
rect 551 -3470 552 -3469
rect 569 -3470 570 -3469
rect 639 -3470 640 -3469
rect 642 -3470 643 -3469
rect 751 -3470 752 -3469
rect 765 -3470 766 -3469
rect 807 -3470 808 -3469
rect 828 -3470 829 -3469
rect 912 -3470 913 -3469
rect 919 -3470 920 -3469
rect 954 -3470 955 -3469
rect 975 -3470 976 -3469
rect 978 -3470 979 -3469
rect 1031 -3470 1032 -3469
rect 1062 -3470 1063 -3469
rect 1080 -3470 1081 -3469
rect 1108 -3470 1109 -3469
rect 1122 -3470 1123 -3469
rect 1185 -3470 1186 -3469
rect 1199 -3470 1200 -3469
rect 1318 -3470 1319 -3469
rect 1430 -3470 1431 -3469
rect 1444 -3470 1445 -3469
rect 1458 -3470 1459 -3469
rect 1570 -3470 1571 -3469
rect 1745 -3470 1746 -3469
rect 1766 -3470 1767 -3469
rect 1790 -3470 1791 -3469
rect 1794 -3470 1795 -3469
rect 1829 -3470 1830 -3469
rect 1836 -3470 1837 -3469
rect 1839 -3470 1840 -3469
rect 1850 -3470 1851 -3469
rect 1860 -3470 1861 -3469
rect 1864 -3470 1865 -3469
rect 1958 -3470 1959 -3469
rect 1962 -3470 1963 -3469
rect 2025 -3470 2026 -3469
rect 2028 -3470 2029 -3469
rect 324 -3472 325 -3471
rect 331 -3472 332 -3471
rect 380 -3472 381 -3471
rect 387 -3472 388 -3471
rect 422 -3472 423 -3471
rect 467 -3472 468 -3471
rect 485 -3472 486 -3471
rect 523 -3472 524 -3471
rect 541 -3472 542 -3471
rect 569 -3472 570 -3471
rect 579 -3472 580 -3471
rect 604 -3472 605 -3471
rect 618 -3472 619 -3471
rect 628 -3472 629 -3471
rect 639 -3472 640 -3471
rect 653 -3472 654 -3471
rect 667 -3472 668 -3471
rect 705 -3472 706 -3471
rect 730 -3472 731 -3471
rect 737 -3472 738 -3471
rect 772 -3472 773 -3471
rect 779 -3472 780 -3471
rect 789 -3472 790 -3471
rect 814 -3472 815 -3471
rect 828 -3472 829 -3471
rect 842 -3472 843 -3471
rect 849 -3472 850 -3471
rect 922 -3472 923 -3471
rect 975 -3472 976 -3471
rect 996 -3472 997 -3471
rect 1017 -3472 1018 -3471
rect 1031 -3472 1032 -3471
rect 1059 -3472 1060 -3471
rect 1073 -3472 1074 -3471
rect 1083 -3472 1084 -3471
rect 1171 -3472 1172 -3471
rect 1178 -3472 1179 -3471
rect 1206 -3472 1207 -3471
rect 1213 -3472 1214 -3471
rect 1272 -3472 1273 -3471
rect 1276 -3472 1277 -3471
rect 1286 -3472 1287 -3471
rect 1307 -3472 1308 -3471
rect 1311 -3472 1312 -3471
rect 1433 -3472 1434 -3471
rect 1451 -3472 1452 -3471
rect 1500 -3472 1501 -3471
rect 1503 -3472 1504 -3471
rect 1507 -3472 1508 -3471
rect 1514 -3472 1515 -3471
rect 1843 -3472 1844 -3471
rect 1850 -3472 1851 -3471
rect 1864 -3472 1865 -3471
rect 1871 -3472 1872 -3471
rect 2025 -3472 2026 -3471
rect 2032 -3472 2033 -3471
rect 471 -3474 472 -3473
rect 523 -3474 524 -3473
rect 562 -3474 563 -3473
rect 604 -3474 605 -3473
rect 653 -3474 654 -3473
rect 744 -3474 745 -3473
rect 800 -3474 801 -3473
rect 887 -3474 888 -3473
rect 1010 -3474 1011 -3473
rect 1017 -3474 1018 -3473
rect 1045 -3474 1046 -3473
rect 1500 -3474 1501 -3473
rect 1822 -3474 1823 -3473
rect 1843 -3474 1844 -3473
rect 2028 -3474 2029 -3473
rect 2032 -3474 2033 -3473
rect 485 -3476 486 -3475
rect 632 -3476 633 -3475
rect 674 -3476 675 -3475
rect 702 -3476 703 -3475
rect 709 -3476 710 -3475
rect 744 -3476 745 -3475
rect 814 -3476 815 -3475
rect 835 -3476 836 -3475
rect 866 -3476 867 -3475
rect 1087 -3476 1088 -3475
rect 1094 -3476 1095 -3475
rect 1125 -3476 1126 -3475
rect 1129 -3476 1130 -3475
rect 1143 -3476 1144 -3475
rect 1178 -3476 1179 -3475
rect 1192 -3476 1193 -3475
rect 1234 -3476 1235 -3475
rect 1262 -3476 1263 -3475
rect 1269 -3476 1270 -3475
rect 1325 -3476 1326 -3475
rect 1493 -3476 1494 -3475
rect 1514 -3476 1515 -3475
rect 506 -3478 507 -3477
rect 541 -3478 542 -3477
rect 590 -3478 591 -3477
rect 597 -3478 598 -3477
rect 632 -3478 633 -3477
rect 660 -3478 661 -3477
rect 681 -3478 682 -3477
rect 751 -3478 752 -3477
rect 821 -3478 822 -3477
rect 842 -3478 843 -3477
rect 870 -3478 871 -3477
rect 877 -3478 878 -3477
rect 884 -3478 885 -3477
rect 915 -3478 916 -3477
rect 1003 -3478 1004 -3477
rect 1010 -3478 1011 -3477
rect 1038 -3478 1039 -3477
rect 1045 -3478 1046 -3477
rect 1059 -3478 1060 -3477
rect 1101 -3478 1102 -3477
rect 1157 -3478 1158 -3477
rect 1192 -3478 1193 -3477
rect 1220 -3478 1221 -3477
rect 1234 -3478 1235 -3477
rect 1255 -3478 1256 -3477
rect 1304 -3478 1305 -3477
rect 1311 -3478 1312 -3477
rect 1332 -3478 1333 -3477
rect 1465 -3478 1466 -3477
rect 1493 -3478 1494 -3477
rect 520 -3480 521 -3479
rect 898 -3480 899 -3479
rect 1024 -3480 1025 -3479
rect 1038 -3480 1039 -3479
rect 1248 -3480 1249 -3479
rect 1304 -3480 1305 -3479
rect 534 -3482 535 -3481
rect 590 -3482 591 -3481
rect 611 -3482 612 -3481
rect 681 -3482 682 -3481
rect 695 -3482 696 -3481
rect 786 -3482 787 -3481
rect 1024 -3482 1025 -3481
rect 1164 -3482 1165 -3481
rect 1241 -3482 1242 -3481
rect 1248 -3482 1249 -3481
rect 1283 -3482 1284 -3481
rect 1290 -3482 1291 -3481
rect 513 -3484 514 -3483
rect 534 -3484 535 -3483
rect 555 -3484 556 -3483
rect 611 -3484 612 -3483
rect 716 -3484 717 -3483
rect 779 -3484 780 -3483
rect 1227 -3484 1228 -3483
rect 1241 -3484 1242 -3483
rect 1290 -3484 1291 -3483
rect 1727 -3484 1728 -3483
rect 688 -3486 689 -3485
rect 716 -3486 717 -3485
rect 737 -3486 738 -3485
rect 758 -3486 759 -3485
rect 723 -3488 724 -3487
rect 758 -3488 759 -3487
rect 331 -3499 332 -3498
rect 338 -3499 339 -3498
rect 394 -3499 395 -3498
rect 429 -3499 430 -3498
rect 432 -3499 433 -3498
rect 471 -3499 472 -3498
rect 523 -3499 524 -3498
rect 653 -3499 654 -3498
rect 681 -3499 682 -3498
rect 709 -3499 710 -3498
rect 716 -3499 717 -3498
rect 730 -3499 731 -3498
rect 775 -3499 776 -3498
rect 891 -3499 892 -3498
rect 968 -3499 969 -3498
rect 975 -3499 976 -3498
rect 996 -3499 997 -3498
rect 1003 -3499 1004 -3498
rect 1038 -3499 1039 -3498
rect 1062 -3499 1063 -3498
rect 1122 -3499 1123 -3498
rect 1290 -3499 1291 -3498
rect 1304 -3499 1305 -3498
rect 1367 -3499 1368 -3498
rect 1430 -3499 1431 -3498
rect 1437 -3499 1438 -3498
rect 1500 -3499 1501 -3498
rect 1507 -3499 1508 -3498
rect 1570 -3499 1571 -3498
rect 1612 -3499 1613 -3498
rect 1724 -3499 1725 -3498
rect 1731 -3499 1732 -3498
rect 1780 -3499 1781 -3498
rect 1790 -3499 1791 -3498
rect 1850 -3499 1851 -3498
rect 1860 -3499 1861 -3498
rect 387 -3501 388 -3500
rect 394 -3501 395 -3500
rect 429 -3501 430 -3500
rect 485 -3501 486 -3500
rect 534 -3501 535 -3500
rect 548 -3501 549 -3500
rect 569 -3501 570 -3500
rect 576 -3501 577 -3500
rect 625 -3501 626 -3500
rect 632 -3501 633 -3500
rect 646 -3501 647 -3500
rect 656 -3501 657 -3500
rect 779 -3501 780 -3500
rect 800 -3501 801 -3500
rect 810 -3501 811 -3500
rect 828 -3501 829 -3500
rect 842 -3501 843 -3500
rect 866 -3501 867 -3500
rect 884 -3501 885 -3500
rect 1024 -3501 1025 -3500
rect 1038 -3501 1039 -3500
rect 1045 -3501 1046 -3500
rect 1143 -3501 1144 -3500
rect 1150 -3501 1151 -3500
rect 1160 -3501 1161 -3500
rect 1178 -3501 1179 -3500
rect 1192 -3501 1193 -3500
rect 1206 -3501 1207 -3500
rect 1234 -3501 1235 -3500
rect 1251 -3501 1252 -3500
rect 1262 -3501 1263 -3500
rect 1276 -3501 1277 -3500
rect 1283 -3501 1284 -3500
rect 1311 -3501 1312 -3500
rect 1493 -3501 1494 -3500
rect 1507 -3501 1508 -3500
rect 1843 -3501 1844 -3500
rect 1850 -3501 1851 -3500
rect 1857 -3501 1858 -3500
rect 1864 -3501 1865 -3500
rect 611 -3503 612 -3502
rect 632 -3503 633 -3502
rect 751 -3503 752 -3502
rect 779 -3503 780 -3502
rect 789 -3503 790 -3502
rect 814 -3503 815 -3502
rect 863 -3503 864 -3502
rect 870 -3503 871 -3502
rect 898 -3503 899 -3502
rect 1024 -3503 1025 -3502
rect 1031 -3503 1032 -3502
rect 1045 -3503 1046 -3502
rect 1234 -3503 1235 -3502
rect 1255 -3503 1256 -3502
rect 611 -3505 612 -3504
rect 618 -3505 619 -3504
rect 751 -3505 752 -3504
rect 758 -3505 759 -3504
rect 1031 -3505 1032 -3504
rect 1059 -3505 1060 -3504
rect 1241 -3505 1242 -3504
rect 1248 -3505 1249 -3504
rect 604 -3507 605 -3506
rect 618 -3507 619 -3506
rect 744 -3507 745 -3506
rect 758 -3507 759 -3506
rect 1059 -3507 1060 -3506
rect 1066 -3507 1067 -3506
rect 590 -3509 591 -3508
rect 604 -3509 605 -3508
rect 744 -3509 745 -3508
rect 765 -3509 766 -3508
rect 1066 -3509 1067 -3508
rect 1080 -3509 1081 -3508
rect 765 -3511 766 -3510
rect 772 -3511 773 -3510
rect 408 -3522 409 -3521
rect 429 -3522 430 -3521
rect 618 -3522 619 -3521
rect 635 -3522 636 -3521
rect 709 -3522 710 -3521
rect 716 -3522 717 -3521
rect 723 -3522 724 -3521
rect 737 -3522 738 -3521
rect 751 -3522 752 -3521
rect 786 -3522 787 -3521
rect 800 -3522 801 -3521
rect 810 -3522 811 -3521
rect 891 -3522 892 -3521
rect 926 -3522 927 -3521
rect 968 -3522 969 -3521
rect 971 -3522 972 -3521
rect 1017 -3522 1018 -3521
rect 1027 -3522 1028 -3521
rect 1038 -3522 1039 -3521
rect 1041 -3522 1042 -3521
rect 1059 -3522 1060 -3521
rect 1066 -3522 1067 -3521
rect 1150 -3522 1151 -3521
rect 1157 -3522 1158 -3521
rect 1206 -3522 1207 -3521
rect 1213 -3522 1214 -3521
rect 1223 -3522 1224 -3521
rect 1234 -3522 1235 -3521
rect 1360 -3522 1361 -3521
rect 1367 -3522 1368 -3521
rect 1507 -3522 1508 -3521
rect 1510 -3522 1511 -3521
rect 1612 -3522 1613 -3521
rect 1633 -3522 1634 -3521
rect 1850 -3522 1851 -3521
rect 1857 -3522 1858 -3521
rect 611 -3524 612 -3523
rect 618 -3524 619 -3523
rect 632 -3524 633 -3523
rect 646 -3524 647 -3523
rect 709 -3524 710 -3523
rect 740 -3524 741 -3523
rect 758 -3524 759 -3523
rect 775 -3524 776 -3523
rect 779 -3524 780 -3523
rect 786 -3524 787 -3523
rect 1024 -3524 1025 -3523
rect 1160 -3524 1161 -3523
rect 1507 -3524 1508 -3523
rect 1514 -3524 1515 -3523
rect 604 -3526 605 -3525
rect 611 -3526 612 -3525
rect 765 -3526 766 -3525
rect 789 -3526 790 -3525
rect 1010 -3526 1011 -3525
rect 1024 -3526 1025 -3525
rect 1038 -3526 1039 -3525
rect 1045 -3526 1046 -3525
rect 1052 -3526 1053 -3525
rect 1059 -3526 1060 -3525
rect 1066 -3526 1067 -3525
rect 1122 -3526 1123 -3525
rect 604 -3528 605 -3527
rect 625 -3528 626 -3527
rect 765 -3528 766 -3527
rect 772 -3528 773 -3527
rect 1003 -3528 1004 -3527
rect 1010 -3528 1011 -3527
rect 1510 -3528 1511 -3527
rect 1514 -3528 1515 -3527
rect 625 -3530 626 -3529
rect 632 -3530 633 -3529
rect 394 -3541 395 -3540
rect 401 -3541 402 -3540
rect 464 -3541 465 -3540
rect 474 -3541 475 -3540
rect 548 -3541 549 -3540
rect 555 -3541 556 -3540
rect 583 -3541 584 -3540
rect 590 -3541 591 -3540
rect 635 -3541 636 -3540
rect 639 -3541 640 -3540
rect 702 -3541 703 -3540
rect 709 -3541 710 -3540
rect 730 -3541 731 -3540
rect 740 -3541 741 -3540
rect 758 -3541 759 -3540
rect 765 -3541 766 -3540
rect 786 -3541 787 -3540
rect 789 -3541 790 -3540
rect 926 -3541 927 -3540
rect 968 -3541 969 -3540
rect 1010 -3541 1011 -3540
rect 1020 -3541 1021 -3540
rect 1027 -3541 1028 -3540
rect 1031 -3541 1032 -3540
rect 1038 -3541 1039 -3540
rect 1045 -3541 1046 -3540
rect 1213 -3541 1214 -3540
rect 1223 -3541 1224 -3540
rect 1507 -3541 1508 -3540
rect 1510 -3541 1511 -3540
rect 1640 -3541 1641 -3540
rect 1647 -3541 1648 -3540
rect 471 -3543 472 -3542
rect 478 -3543 479 -3542
rect 576 -3543 577 -3542
rect 583 -3543 584 -3542
rect 730 -3543 731 -3542
rect 744 -3543 745 -3542
rect 1038 -3543 1039 -3542
rect 1066 -3543 1067 -3542
rect 1507 -3543 1508 -3542
rect 1521 -3543 1522 -3542
rect 1633 -3543 1634 -3542
rect 1640 -3543 1641 -3542
rect 1510 -3545 1511 -3544
rect 1521 -3545 1522 -3544
rect 401 -3556 402 -3555
rect 404 -3556 405 -3555
rect 541 -3556 542 -3555
rect 548 -3556 549 -3555
rect 551 -3556 552 -3555
rect 555 -3556 556 -3555
rect 586 -3556 587 -3555
rect 590 -3556 591 -3555
rect 604 -3556 605 -3555
rect 607 -3556 608 -3555
rect 646 -3556 647 -3555
rect 649 -3556 650 -3555
rect 789 -3556 790 -3555
rect 793 -3556 794 -3555
rect 1017 -3556 1018 -3555
rect 1038 -3556 1039 -3555
rect 1059 -3556 1060 -3555
rect 1066 -3556 1067 -3555
rect 1517 -3556 1518 -3555
rect 1521 -3556 1522 -3555
rect 2028 -3556 2029 -3555
rect 2032 -3556 2033 -3555
rect 401 -3558 402 -3557
rect 408 -3558 409 -3557
rect 604 -3558 605 -3557
rect 611 -3558 612 -3557
rect 1514 -3558 1515 -3557
rect 1521 -3558 1522 -3557
rect 607 -3560 608 -3559
rect 611 -3560 612 -3559
rect 1507 -3560 1508 -3559
rect 1514 -3560 1515 -3559
rect 401 -3571 402 -3570
rect 404 -3571 405 -3570
rect 1062 -3571 1063 -3570
rect 1066 -3571 1067 -3570
rect 1514 -3571 1515 -3570
rect 1521 -3571 1522 -3570
rect 401 -3573 402 -3572
rect 408 -3573 409 -3572
rect 404 -3575 405 -3574
rect 408 -3575 409 -3574
rect 394 -3586 395 -3585
rect 401 -3586 402 -3585
rect 618 -3586 619 -3585
rect 621 -3586 622 -3585
rect 723 -3586 724 -3585
rect 726 -3586 727 -3585
rect 401 -3588 402 -3587
rect 408 -3588 409 -3587
rect 716 -3588 717 -3587
rect 723 -3588 724 -3587
rect 723 -3599 724 -3598
rect 730 -3599 731 -3598
rect 695 -3610 696 -3609
rect 705 -3610 706 -3609
rect 1640 -3610 1641 -3609
rect 1643 -3610 1644 -3609
rect 758 -3621 759 -3620
rect 765 -3621 766 -3620
rect 1640 -3621 1641 -3620
rect 1647 -3621 1648 -3620
rect 761 -3632 762 -3631
rect 765 -3632 766 -3631
rect 394 -3654 395 -3653
rect 397 -3654 398 -3653
rect 695 -3654 696 -3653
rect 698 -3654 699 -3653
rect 394 -3656 395 -3655
rect 401 -3656 402 -3655
rect 397 -3658 398 -3657
rect 401 -3658 402 -3657
rect 397 -3669 398 -3668
rect 401 -3669 402 -3668
rect 604 -3669 605 -3668
rect 611 -3669 612 -3668
<< metal2 >>
rect 254 -19 255 1
rect 432 -19 433 1
rect 485 -19 486 1
rect 632 -19 633 1
rect 635 -19 636 1
rect 772 -19 773 1
rect 796 -19 797 1
rect 814 -19 815 1
rect 824 -19 825 1
rect 961 -19 962 1
rect 968 -19 969 1
rect 1206 -19 1207 1
rect 352 -19 353 -1
rect 572 -19 573 -1
rect 576 -19 577 -1
rect 681 -19 682 -1
rect 688 -19 689 -1
rect 765 -19 766 -1
rect 800 -19 801 -1
rect 891 -19 892 -1
rect 978 -19 979 -1
rect 982 -19 983 -1
rect 1038 -19 1039 -1
rect 1437 -19 1438 -1
rect 397 -19 398 -3
rect 548 -19 549 -3
rect 555 -19 556 -3
rect 583 -19 584 -3
rect 604 -19 605 -3
rect 842 -19 843 -3
rect 863 -19 864 -3
rect 919 -19 920 -3
rect 1073 -19 1074 -3
rect 1129 -19 1130 -3
rect 415 -19 416 -5
rect 422 -19 423 -5
rect 611 -19 612 -5
rect 625 -19 626 -5
rect 639 -19 640 -5
rect 845 -19 846 -5
rect 884 -19 885 -5
rect 1087 -19 1088 -5
rect 1094 -19 1095 -5
rect 1125 -19 1126 -5
rect 618 -19 619 -7
rect 852 -19 853 -7
rect 646 -19 647 -9
rect 705 -19 706 -9
rect 709 -19 710 -9
rect 915 -19 916 -9
rect 663 -19 664 -11
rect 989 -19 990 -11
rect 716 -19 717 -13
rect 821 -19 822 -13
rect 828 -19 829 -13
rect 887 -19 888 -13
rect 730 -19 731 -15
rect 803 -19 804 -15
rect 810 -19 811 -15
rect 870 -19 871 -15
rect 835 -19 836 -17
rect 859 -19 860 -17
rect 184 -66 185 -28
rect 212 -29 213 -27
rect 240 -66 241 -28
rect 397 -29 398 -27
rect 404 -66 405 -28
rect 478 -66 479 -28
rect 492 -66 493 -28
rect 618 -29 619 -27
rect 646 -29 647 -27
rect 723 -66 724 -28
rect 737 -66 738 -28
rect 758 -66 759 -28
rect 765 -66 766 -28
rect 828 -29 829 -27
rect 842 -29 843 -27
rect 1220 -66 1221 -28
rect 1234 -66 1235 -28
rect 1360 -66 1361 -28
rect 1437 -29 1438 -27
rect 1486 -66 1487 -28
rect 1629 -29 1630 -27
rect 1633 -66 1634 -28
rect 198 -66 199 -30
rect 254 -31 255 -27
rect 275 -66 276 -30
rect 313 -66 314 -30
rect 317 -66 318 -30
rect 660 -31 661 -27
rect 667 -66 668 -30
rect 740 -66 741 -30
rect 744 -66 745 -30
rect 863 -31 864 -27
rect 870 -31 871 -27
rect 884 -66 885 -30
rect 908 -66 909 -30
rect 947 -66 948 -30
rect 961 -31 962 -27
rect 1045 -66 1046 -30
rect 1066 -66 1067 -30
rect 1101 -66 1102 -30
rect 1108 -66 1109 -30
rect 1150 -66 1151 -30
rect 1206 -31 1207 -27
rect 1290 -66 1291 -30
rect 1321 -66 1322 -30
rect 1332 -66 1333 -30
rect 1440 -31 1441 -27
rect 1759 -66 1760 -30
rect 296 -66 297 -32
rect 352 -33 353 -27
rect 355 -66 356 -32
rect 464 -66 465 -32
rect 471 -66 472 -32
rect 611 -33 612 -27
rect 618 -66 619 -32
rect 625 -33 626 -27
rect 660 -66 661 -32
rect 695 -66 696 -32
rect 702 -33 703 -27
rect 821 -66 822 -32
rect 828 -66 829 -32
rect 1038 -33 1039 -27
rect 1087 -33 1088 -27
rect 1178 -66 1179 -32
rect 394 -66 395 -34
rect 485 -35 486 -27
rect 499 -66 500 -34
rect 639 -35 640 -27
rect 677 -66 678 -34
rect 975 -66 976 -34
rect 978 -35 979 -27
rect 1003 -66 1004 -34
rect 1010 -66 1011 -34
rect 1094 -35 1095 -27
rect 1132 -35 1133 -27
rect 1213 -66 1214 -34
rect 415 -66 416 -36
rect 422 -37 423 -27
rect 432 -37 433 -27
rect 590 -66 591 -36
rect 611 -66 612 -36
rect 656 -37 657 -27
rect 702 -66 703 -36
rect 716 -37 717 -27
rect 751 -66 752 -36
rect 887 -37 888 -27
rect 912 -37 913 -27
rect 1017 -66 1018 -36
rect 1073 -37 1074 -27
rect 1087 -66 1088 -36
rect 1094 -66 1095 -36
rect 1115 -66 1116 -36
rect 422 -66 423 -38
rect 446 -39 447 -27
rect 485 -66 486 -38
rect 604 -39 605 -27
rect 639 -66 640 -38
rect 653 -39 654 -27
rect 716 -66 717 -38
rect 807 -39 808 -27
rect 842 -66 843 -38
rect 898 -39 899 -27
rect 926 -66 927 -38
rect 1125 -66 1126 -38
rect 506 -66 507 -40
rect 852 -66 853 -40
rect 856 -66 857 -40
rect 1038 -66 1039 -40
rect 520 -66 521 -42
rect 576 -43 577 -27
rect 583 -43 584 -27
rect 646 -66 647 -42
rect 653 -66 654 -42
rect 961 -66 962 -42
rect 982 -43 983 -27
rect 1031 -66 1032 -42
rect 534 -66 535 -44
rect 688 -45 689 -27
rect 768 -45 769 -27
rect 863 -66 864 -44
rect 870 -66 871 -44
rect 919 -45 920 -27
rect 982 -66 983 -44
rect 1069 -66 1070 -44
rect 548 -47 549 -27
rect 597 -66 598 -46
rect 604 -66 605 -46
rect 901 -66 902 -46
rect 989 -47 990 -27
rect 1059 -66 1060 -46
rect 548 -66 549 -48
rect 572 -49 573 -27
rect 583 -66 584 -48
rect 933 -66 934 -48
rect 1024 -66 1025 -48
rect 1073 -66 1074 -48
rect 569 -51 570 -27
rect 779 -66 780 -50
rect 793 -66 794 -50
rect 835 -51 836 -27
rect 849 -51 850 -27
rect 1080 -66 1081 -50
rect 569 -66 570 -52
rect 674 -66 675 -52
rect 688 -66 689 -52
rect 709 -53 710 -27
rect 772 -53 773 -27
rect 835 -66 836 -52
rect 849 -66 850 -52
rect 912 -66 913 -52
rect 709 -66 710 -54
rect 730 -55 731 -27
rect 772 -66 773 -54
rect 810 -55 811 -27
rect 877 -66 878 -54
rect 940 -66 941 -54
rect 730 -66 731 -56
rect 968 -57 969 -27
rect 800 -66 801 -58
rect 919 -66 920 -58
rect 807 -66 808 -60
rect 814 -61 815 -27
rect 887 -66 888 -60
rect 1052 -66 1053 -60
rect 681 -63 682 -27
rect 814 -66 815 -62
rect 891 -63 892 -27
rect 989 -66 990 -62
rect 565 -66 566 -64
rect 681 -66 682 -64
rect 803 -66 804 -64
rect 891 -66 892 -64
rect 915 -65 916 -27
rect 968 -66 969 -64
rect 58 -143 59 -75
rect 523 -143 524 -75
rect 530 -143 531 -75
rect 1241 -143 1242 -75
rect 1290 -76 1291 -74
rect 1297 -143 1298 -75
rect 1332 -76 1333 -74
rect 1374 -143 1375 -75
rect 1486 -76 1487 -74
rect 1514 -143 1515 -75
rect 1633 -76 1634 -74
rect 1640 -143 1641 -75
rect 1759 -76 1760 -74
rect 1885 -143 1886 -75
rect 65 -143 66 -77
rect 226 -143 227 -77
rect 233 -143 234 -77
rect 849 -143 850 -77
rect 852 -78 853 -74
rect 1136 -143 1137 -77
rect 1157 -143 1158 -77
rect 1167 -78 1168 -74
rect 1171 -143 1172 -77
rect 1269 -143 1270 -77
rect 1360 -78 1361 -74
rect 1423 -143 1424 -77
rect 72 -143 73 -79
rect 401 -80 402 -74
rect 404 -80 405 -74
rect 436 -143 437 -79
rect 450 -143 451 -79
rect 520 -80 521 -74
rect 555 -143 556 -79
rect 660 -80 661 -74
rect 674 -143 675 -79
rect 709 -80 710 -74
rect 740 -143 741 -79
rect 1325 -143 1326 -79
rect 79 -143 80 -81
rect 352 -82 353 -74
rect 359 -143 360 -81
rect 422 -82 423 -74
rect 429 -143 430 -81
rect 604 -82 605 -74
rect 625 -143 626 -81
rect 828 -82 829 -74
rect 835 -82 836 -74
rect 905 -143 906 -81
rect 919 -82 920 -74
rect 940 -143 941 -81
rect 943 -82 944 -74
rect 1290 -143 1291 -81
rect 1321 -82 1322 -74
rect 1360 -143 1361 -81
rect 86 -143 87 -83
rect 264 -143 265 -83
rect 282 -143 283 -83
rect 499 -84 500 -74
rect 513 -143 514 -83
rect 541 -84 542 -74
rect 562 -143 563 -83
rect 632 -143 633 -83
rect 653 -143 654 -83
rect 765 -84 766 -74
rect 786 -143 787 -83
rect 821 -84 822 -74
rect 856 -84 857 -74
rect 1122 -143 1123 -83
rect 1125 -84 1126 -74
rect 1318 -143 1319 -83
rect 93 -143 94 -85
rect 471 -86 472 -74
rect 478 -86 479 -74
rect 478 -143 479 -85
rect 478 -86 479 -74
rect 478 -143 479 -85
rect 499 -143 500 -85
rect 527 -143 528 -85
rect 541 -143 542 -85
rect 611 -86 612 -74
rect 660 -143 661 -85
rect 751 -86 752 -74
rect 779 -86 780 -74
rect 821 -143 822 -85
rect 856 -143 857 -85
rect 1010 -86 1011 -74
rect 1031 -86 1032 -74
rect 1031 -143 1032 -85
rect 1031 -86 1032 -74
rect 1031 -143 1032 -85
rect 1038 -86 1039 -74
rect 1108 -143 1109 -85
rect 1115 -143 1116 -85
rect 1150 -86 1151 -74
rect 1178 -86 1179 -74
rect 1255 -143 1256 -85
rect 100 -143 101 -87
rect 600 -143 601 -87
rect 604 -143 605 -87
rect 618 -88 619 -74
rect 702 -88 703 -74
rect 828 -143 829 -87
rect 863 -88 864 -74
rect 884 -143 885 -87
rect 919 -143 920 -87
rect 968 -88 969 -74
rect 975 -88 976 -74
rect 1283 -143 1284 -87
rect 107 -143 108 -89
rect 184 -90 185 -74
rect 191 -143 192 -89
rect 240 -90 241 -74
rect 247 -143 248 -89
rect 443 -143 444 -89
rect 471 -143 472 -89
rect 975 -143 976 -89
rect 989 -90 990 -74
rect 1192 -143 1193 -89
rect 1213 -90 1214 -74
rect 1304 -143 1305 -89
rect 114 -143 115 -91
rect 236 -143 237 -91
rect 240 -143 241 -91
rect 275 -92 276 -74
rect 296 -92 297 -74
rect 331 -143 332 -91
rect 338 -143 339 -91
rect 649 -143 650 -91
rect 702 -143 703 -91
rect 870 -92 871 -74
rect 898 -92 899 -74
rect 1213 -143 1214 -91
rect 1220 -92 1221 -74
rect 1353 -143 1354 -91
rect 124 -143 125 -93
rect 303 -143 304 -93
rect 310 -94 311 -74
rect 324 -143 325 -93
rect 345 -143 346 -93
rect 544 -94 545 -74
rect 576 -143 577 -93
rect 639 -94 640 -74
rect 709 -143 710 -93
rect 716 -94 717 -74
rect 751 -143 752 -93
rect 1234 -94 1235 -74
rect 1237 -94 1238 -74
rect 1507 -143 1508 -93
rect 128 -143 129 -95
rect 583 -96 584 -74
rect 590 -96 591 -74
rect 611 -143 612 -95
rect 618 -143 619 -95
rect 957 -96 958 -74
rect 961 -96 962 -74
rect 1150 -143 1151 -95
rect 1227 -96 1228 -74
rect 1311 -143 1312 -95
rect 135 -143 136 -97
rect 506 -98 507 -74
rect 583 -143 584 -97
rect 597 -98 598 -74
rect 639 -143 640 -97
rect 835 -143 836 -97
rect 863 -143 864 -97
rect 877 -98 878 -74
rect 954 -98 955 -74
rect 989 -143 990 -97
rect 999 -98 1000 -74
rect 1094 -98 1095 -74
rect 1101 -98 1102 -74
rect 1276 -143 1277 -97
rect 149 -143 150 -99
rect 352 -143 353 -99
rect 366 -143 367 -99
rect 569 -100 570 -74
rect 758 -100 759 -74
rect 898 -143 899 -99
rect 933 -100 934 -74
rect 1101 -143 1102 -99
rect 1118 -100 1119 -74
rect 1185 -143 1186 -99
rect 152 -143 153 -101
rect 289 -143 290 -101
rect 310 -143 311 -101
rect 859 -102 860 -74
rect 870 -143 871 -101
rect 982 -102 983 -74
rect 996 -102 997 -74
rect 1094 -143 1095 -101
rect 156 -143 157 -103
rect 317 -104 318 -74
rect 380 -143 381 -103
rect 492 -104 493 -74
rect 730 -104 731 -74
rect 758 -143 759 -103
rect 779 -143 780 -103
rect 908 -104 909 -74
rect 912 -104 913 -74
rect 982 -143 983 -103
rect 1003 -104 1004 -74
rect 1164 -143 1165 -103
rect 163 -143 164 -105
rect 698 -143 699 -105
rect 789 -106 790 -74
rect 800 -106 801 -74
rect 803 -143 804 -105
rect 954 -143 955 -105
rect 968 -143 969 -105
rect 1017 -106 1018 -74
rect 1027 -106 1028 -74
rect 1234 -143 1235 -105
rect 170 -143 171 -107
rect 408 -108 409 -74
rect 411 -108 412 -74
rect 415 -108 416 -74
rect 422 -143 423 -107
rect 548 -108 549 -74
rect 807 -108 808 -74
rect 1003 -143 1004 -107
rect 1010 -143 1011 -107
rect 1143 -143 1144 -107
rect 177 -143 178 -109
rect 534 -110 535 -74
rect 548 -143 549 -109
rect 744 -110 745 -74
rect 807 -143 808 -109
rect 926 -110 927 -74
rect 933 -143 934 -109
rect 1199 -143 1200 -109
rect 184 -143 185 -111
rect 656 -112 657 -74
rect 744 -143 745 -111
rect 842 -112 843 -74
rect 947 -112 948 -74
rect 996 -143 997 -111
rect 1017 -143 1018 -111
rect 1059 -112 1060 -74
rect 1073 -112 1074 -74
rect 1220 -143 1221 -111
rect 198 -114 199 -74
rect 219 -143 220 -113
rect 229 -143 230 -113
rect 317 -143 318 -113
rect 373 -143 374 -113
rect 730 -143 731 -113
rect 814 -114 815 -74
rect 877 -143 878 -113
rect 912 -143 913 -113
rect 947 -143 948 -113
rect 1024 -114 1025 -74
rect 1059 -143 1060 -113
rect 1080 -114 1081 -74
rect 1178 -143 1179 -113
rect 198 -143 199 -115
rect 474 -143 475 -115
rect 492 -143 493 -115
rect 765 -143 766 -115
rect 891 -116 892 -74
rect 1080 -143 1081 -115
rect 1087 -116 1088 -74
rect 1206 -143 1207 -115
rect 205 -143 206 -117
rect 467 -143 468 -117
rect 534 -143 535 -117
rect 1076 -143 1077 -117
rect 1087 -143 1088 -117
rect 1248 -143 1249 -117
rect 212 -143 213 -119
rect 387 -143 388 -119
rect 390 -143 391 -119
rect 569 -143 570 -119
rect 597 -143 598 -119
rect 891 -143 892 -119
rect 1038 -143 1039 -119
rect 1111 -120 1112 -74
rect 261 -143 262 -121
rect 677 -122 678 -74
rect 681 -122 682 -74
rect 1024 -143 1025 -121
rect 1045 -122 1046 -74
rect 1129 -143 1130 -121
rect 275 -143 276 -123
rect 394 -124 395 -74
rect 401 -143 402 -123
rect 485 -124 486 -74
rect 646 -124 647 -74
rect 842 -143 843 -123
rect 1052 -124 1053 -74
rect 1066 -143 1067 -123
rect 296 -143 297 -125
rect 681 -143 682 -125
rect 688 -126 689 -74
rect 814 -143 815 -125
rect 142 -143 143 -127
rect 688 -143 689 -127
rect 723 -128 724 -74
rect 1052 -143 1053 -127
rect 394 -143 395 -129
rect 737 -143 738 -129
rect 408 -143 409 -131
rect 565 -132 566 -74
rect 723 -143 724 -131
rect 793 -132 794 -74
rect 121 -143 122 -133
rect 793 -143 794 -133
rect 415 -143 416 -135
rect 464 -136 465 -74
rect 485 -143 486 -135
rect 667 -136 668 -74
rect 446 -143 447 -137
rect 590 -143 591 -137
rect 667 -143 668 -137
rect 772 -138 773 -74
rect 457 -143 458 -139
rect 506 -143 507 -139
rect 565 -143 566 -139
rect 716 -143 717 -139
rect 772 -143 773 -139
rect 1045 -143 1046 -139
rect 460 -143 461 -141
rect 1227 -143 1228 -141
rect 16 -246 17 -152
rect 261 -153 262 -151
rect 282 -153 283 -151
rect 387 -246 388 -152
rect 408 -153 409 -151
rect 695 -153 696 -151
rect 768 -153 769 -151
rect 1346 -246 1347 -152
rect 1353 -153 1354 -151
rect 1367 -246 1368 -152
rect 1374 -153 1375 -151
rect 1500 -246 1501 -152
rect 1507 -153 1508 -151
rect 1626 -246 1627 -152
rect 1640 -153 1641 -151
rect 1668 -246 1669 -152
rect 1885 -153 1886 -151
rect 1941 -246 1942 -152
rect 23 -246 24 -154
rect 107 -155 108 -151
rect 114 -155 115 -151
rect 226 -155 227 -151
rect 240 -155 241 -151
rect 268 -155 269 -151
rect 282 -246 283 -154
rect 331 -155 332 -151
rect 345 -155 346 -151
rect 530 -155 531 -151
rect 541 -155 542 -151
rect 600 -155 601 -151
rect 611 -155 612 -151
rect 737 -155 738 -151
rect 803 -155 804 -151
rect 940 -155 941 -151
rect 950 -155 951 -151
rect 1402 -246 1403 -154
rect 1423 -155 1424 -151
rect 1493 -246 1494 -154
rect 1514 -155 1515 -151
rect 1556 -246 1557 -154
rect 1566 -246 1567 -154
rect 1584 -246 1585 -154
rect 1615 -246 1616 -154
rect 1633 -246 1634 -154
rect 37 -246 38 -156
rect 257 -157 258 -151
rect 289 -157 290 -151
rect 289 -246 290 -156
rect 289 -157 290 -151
rect 289 -246 290 -156
rect 331 -246 332 -156
rect 415 -157 416 -151
rect 422 -157 423 -151
rect 443 -246 444 -156
rect 450 -157 451 -151
rect 537 -246 538 -156
rect 541 -246 542 -156
rect 555 -157 556 -151
rect 590 -157 591 -151
rect 681 -246 682 -156
rect 684 -157 685 -151
rect 926 -246 927 -156
rect 1013 -246 1014 -156
rect 1430 -246 1431 -156
rect 1542 -246 1543 -156
rect 1815 -246 1816 -156
rect 44 -246 45 -158
rect 72 -159 73 -151
rect 86 -159 87 -151
rect 765 -159 766 -151
rect 814 -159 815 -151
rect 940 -246 941 -158
rect 1076 -159 1077 -151
rect 1248 -159 1249 -151
rect 1276 -159 1277 -151
rect 1570 -246 1571 -158
rect 51 -246 52 -160
rect 79 -161 80 -151
rect 93 -161 94 -151
rect 646 -246 647 -160
rect 649 -161 650 -151
rect 1080 -161 1081 -151
rect 1090 -161 1091 -151
rect 1465 -246 1466 -160
rect 72 -246 73 -162
rect 366 -163 367 -151
rect 380 -163 381 -151
rect 408 -246 409 -162
rect 429 -163 430 -151
rect 457 -246 458 -162
rect 467 -163 468 -151
rect 1024 -163 1025 -151
rect 1073 -163 1074 -151
rect 1248 -246 1249 -162
rect 1283 -163 1284 -151
rect 1577 -246 1578 -162
rect 79 -246 80 -164
rect 93 -246 94 -164
rect 100 -165 101 -151
rect 124 -165 125 -151
rect 128 -165 129 -151
rect 152 -165 153 -151
rect 163 -165 164 -151
rect 233 -246 234 -164
rect 240 -246 241 -164
rect 1507 -246 1508 -164
rect 100 -246 101 -166
rect 565 -167 566 -151
rect 618 -167 619 -151
rect 695 -246 696 -166
rect 737 -246 738 -166
rect 1010 -167 1011 -151
rect 1073 -246 1074 -166
rect 1108 -167 1109 -151
rect 1129 -167 1130 -151
rect 1451 -246 1452 -166
rect 107 -246 108 -168
rect 569 -169 570 -151
rect 621 -246 622 -168
rect 730 -246 731 -168
rect 814 -246 815 -168
rect 838 -169 839 -151
rect 849 -169 850 -151
rect 947 -169 948 -151
rect 975 -169 976 -151
rect 1276 -246 1277 -168
rect 1290 -169 1291 -151
rect 1374 -246 1375 -168
rect 117 -246 118 -170
rect 611 -246 612 -170
rect 849 -246 850 -170
rect 877 -171 878 -151
rect 884 -171 885 -151
rect 1108 -246 1109 -170
rect 1122 -171 1123 -151
rect 1290 -246 1291 -170
rect 1304 -171 1305 -151
rect 1444 -246 1445 -170
rect 121 -246 122 -172
rect 201 -246 202 -172
rect 226 -246 227 -172
rect 772 -173 773 -151
rect 856 -173 857 -151
rect 877 -246 878 -172
rect 887 -246 888 -172
rect 1227 -173 1228 -151
rect 1311 -173 1312 -151
rect 1472 -246 1473 -172
rect 128 -246 129 -174
rect 254 -175 255 -151
rect 275 -175 276 -151
rect 429 -246 430 -174
rect 450 -246 451 -174
rect 478 -175 479 -151
rect 492 -175 493 -151
rect 597 -246 598 -174
rect 667 -175 668 -151
rect 772 -246 773 -174
rect 870 -175 871 -151
rect 1024 -246 1025 -174
rect 1059 -175 1060 -151
rect 1129 -246 1130 -174
rect 1136 -175 1137 -151
rect 1395 -246 1396 -174
rect 65 -177 66 -151
rect 254 -246 255 -176
rect 275 -246 276 -176
rect 359 -177 360 -151
rect 366 -246 367 -176
rect 894 -246 895 -176
rect 905 -177 906 -151
rect 975 -246 976 -176
rect 989 -177 990 -151
rect 1136 -246 1137 -176
rect 1150 -177 1151 -151
rect 1283 -246 1284 -176
rect 1318 -177 1319 -151
rect 1437 -246 1438 -176
rect 135 -179 136 -151
rect 261 -246 262 -178
rect 338 -179 339 -151
rect 478 -246 479 -178
rect 513 -179 514 -151
rect 562 -246 563 -178
rect 569 -246 570 -178
rect 929 -179 930 -151
rect 961 -179 962 -151
rect 1304 -246 1305 -178
rect 1325 -179 1326 -151
rect 1591 -246 1592 -178
rect 142 -246 143 -180
rect 212 -181 213 -151
rect 243 -246 244 -180
rect 271 -246 272 -180
rect 296 -181 297 -151
rect 338 -246 339 -180
rect 345 -246 346 -180
rect 485 -181 486 -151
rect 513 -246 514 -180
rect 593 -246 594 -180
rect 705 -246 706 -180
rect 1227 -246 1228 -180
rect 1325 -246 1326 -180
rect 1332 -246 1333 -180
rect 1360 -181 1361 -151
rect 1458 -246 1459 -180
rect 145 -183 146 -151
rect 156 -183 157 -151
rect 163 -246 164 -182
rect 390 -183 391 -151
rect 401 -183 402 -151
rect 415 -246 416 -182
rect 471 -246 472 -182
rect 1010 -246 1011 -182
rect 1017 -183 1018 -151
rect 1122 -246 1123 -182
rect 1164 -183 1165 -151
rect 1423 -246 1424 -182
rect 149 -246 150 -184
rect 716 -185 717 -151
rect 786 -185 787 -151
rect 905 -246 906 -184
rect 919 -185 920 -151
rect 1059 -246 1060 -184
rect 1080 -246 1081 -184
rect 1115 -185 1116 -151
rect 1171 -185 1172 -151
rect 1388 -246 1389 -184
rect 156 -246 157 -186
rect 1514 -246 1515 -186
rect 170 -189 171 -151
rect 492 -246 493 -188
rect 520 -189 521 -151
rect 989 -246 990 -188
rect 1003 -189 1004 -151
rect 1360 -246 1361 -188
rect 177 -191 178 -151
rect 359 -246 360 -190
rect 373 -191 374 -151
rect 667 -246 668 -190
rect 709 -191 710 -151
rect 856 -246 857 -190
rect 912 -191 913 -151
rect 919 -246 920 -190
rect 954 -191 955 -151
rect 1164 -246 1165 -190
rect 1171 -246 1172 -190
rect 1265 -191 1266 -151
rect 177 -246 178 -192
rect 436 -193 437 -151
rect 520 -246 521 -192
rect 947 -246 948 -192
rect 968 -193 969 -151
rect 1115 -246 1116 -192
rect 1174 -193 1175 -151
rect 1241 -193 1242 -151
rect 58 -195 59 -151
rect 436 -246 437 -194
rect 527 -195 528 -151
rect 1052 -195 1053 -151
rect 1094 -195 1095 -151
rect 1521 -246 1522 -194
rect 58 -246 59 -196
rect 159 -246 160 -196
rect 184 -197 185 -151
rect 296 -246 297 -196
rect 310 -197 311 -151
rect 485 -246 486 -196
rect 506 -197 507 -151
rect 527 -246 528 -196
rect 534 -197 535 -151
rect 716 -246 717 -196
rect 758 -197 759 -151
rect 786 -246 787 -196
rect 793 -197 794 -151
rect 961 -246 962 -196
rect 1017 -246 1018 -196
rect 1150 -246 1151 -196
rect 1178 -197 1179 -151
rect 1353 -246 1354 -196
rect 170 -246 171 -198
rect 310 -246 311 -198
rect 317 -199 318 -151
rect 373 -246 374 -198
rect 394 -199 395 -151
rect 506 -246 507 -198
rect 555 -246 556 -198
rect 779 -199 780 -151
rect 821 -199 822 -151
rect 870 -246 871 -198
rect 1038 -199 1039 -151
rect 1052 -246 1053 -198
rect 1094 -246 1095 -198
rect 1143 -199 1144 -151
rect 1185 -199 1186 -151
rect 1409 -246 1410 -198
rect 184 -246 185 -200
rect 460 -201 461 -151
rect 674 -201 675 -151
rect 968 -246 969 -200
rect 1038 -246 1039 -200
rect 1549 -246 1550 -200
rect 194 -246 195 -202
rect 933 -246 934 -202
rect 1101 -203 1102 -151
rect 1416 -246 1417 -202
rect 198 -205 199 -151
rect 422 -246 423 -204
rect 660 -205 661 -151
rect 674 -246 675 -204
rect 688 -205 689 -151
rect 954 -246 955 -204
rect 1066 -205 1067 -151
rect 1101 -246 1102 -204
rect 1143 -246 1144 -204
rect 1269 -205 1270 -151
rect 30 -246 31 -206
rect 198 -246 199 -206
rect 212 -246 213 -206
rect 821 -246 822 -206
rect 898 -207 899 -151
rect 1185 -246 1186 -206
rect 1192 -207 1193 -151
rect 1528 -246 1529 -206
rect 219 -209 220 -151
rect 317 -246 318 -208
rect 324 -209 325 -151
rect 394 -246 395 -208
rect 401 -246 402 -208
rect 639 -209 640 -151
rect 698 -209 699 -151
rect 1192 -246 1193 -208
rect 1199 -209 1200 -151
rect 1486 -246 1487 -208
rect 219 -246 220 -210
rect 499 -211 500 -151
rect 548 -211 549 -151
rect 660 -246 661 -210
rect 709 -246 710 -210
rect 1234 -211 1235 -151
rect 1241 -246 1242 -210
rect 1297 -211 1298 -151
rect 247 -213 248 -151
rect 999 -246 1000 -212
rect 1031 -213 1032 -151
rect 1066 -246 1067 -212
rect 1157 -213 1158 -151
rect 1234 -246 1235 -212
rect 1255 -213 1256 -151
rect 1297 -246 1298 -212
rect 89 -246 90 -214
rect 247 -246 248 -214
rect 324 -246 325 -214
rect 1262 -215 1263 -151
rect 1269 -246 1270 -214
rect 1612 -246 1613 -214
rect 352 -217 353 -151
rect 380 -246 381 -216
rect 499 -246 500 -216
rect 751 -217 752 -151
rect 758 -246 759 -216
rect 1087 -217 1088 -151
rect 1199 -246 1200 -216
rect 1381 -246 1382 -216
rect 352 -246 353 -218
rect 523 -219 524 -151
rect 548 -246 549 -218
rect 915 -246 916 -218
rect 996 -219 997 -151
rect 1087 -246 1088 -218
rect 1202 -246 1203 -218
rect 1339 -246 1340 -218
rect 523 -246 524 -220
rect 842 -221 843 -151
rect 863 -221 864 -151
rect 1031 -246 1032 -220
rect 1045 -221 1046 -151
rect 1157 -246 1158 -220
rect 1206 -221 1207 -151
rect 1479 -246 1480 -220
rect 583 -223 584 -151
rect 751 -246 752 -222
rect 765 -246 766 -222
rect 1178 -246 1179 -222
rect 1213 -223 1214 -151
rect 1311 -246 1312 -222
rect 576 -225 577 -151
rect 583 -246 584 -224
rect 604 -225 605 -151
rect 688 -246 689 -224
rect 702 -225 703 -151
rect 863 -246 864 -224
rect 891 -225 892 -151
rect 1262 -246 1263 -224
rect 303 -227 304 -151
rect 604 -246 605 -226
rect 632 -227 633 -151
rect 842 -246 843 -226
rect 982 -227 983 -151
rect 1045 -246 1046 -226
rect 1216 -246 1217 -226
rect 1318 -246 1319 -226
rect 205 -229 206 -151
rect 303 -246 304 -228
rect 576 -246 577 -228
rect 733 -229 734 -151
rect 744 -229 745 -151
rect 793 -246 794 -228
rect 807 -229 808 -151
rect 898 -246 899 -228
rect 936 -229 937 -151
rect 982 -246 983 -228
rect 1003 -246 1004 -228
rect 1213 -246 1214 -228
rect 1220 -229 1221 -151
rect 1535 -246 1536 -228
rect 439 -246 440 -230
rect 1220 -246 1221 -230
rect 1255 -246 1256 -230
rect 1328 -246 1329 -230
rect 625 -233 626 -151
rect 632 -246 633 -232
rect 639 -246 640 -232
rect 712 -246 713 -232
rect 779 -246 780 -232
rect 1146 -233 1147 -151
rect 191 -235 192 -151
rect 625 -246 626 -234
rect 653 -235 654 -151
rect 744 -246 745 -234
rect 807 -246 808 -234
rect 884 -246 885 -234
rect 135 -246 136 -236
rect 653 -246 654 -236
rect 835 -237 836 -151
rect 1206 -246 1207 -236
rect 800 -239 801 -151
rect 835 -246 836 -238
rect 800 -246 801 -240
rect 828 -241 829 -151
rect 723 -243 724 -151
rect 828 -246 829 -242
rect 534 -246 535 -244
rect 723 -246 724 -244
rect 16 -256 17 -254
rect 194 -256 195 -254
rect 198 -371 199 -255
rect 338 -256 339 -254
rect 366 -256 367 -254
rect 747 -371 748 -255
rect 761 -371 762 -255
rect 915 -256 916 -254
rect 992 -256 993 -254
rect 1598 -371 1599 -255
rect 1612 -256 1613 -254
rect 1969 -371 1970 -255
rect 16 -371 17 -257
rect 149 -258 150 -254
rect 156 -258 157 -254
rect 537 -258 538 -254
rect 618 -258 619 -254
rect 800 -258 801 -254
rect 810 -371 811 -257
rect 1801 -371 1802 -257
rect 1815 -258 1816 -254
rect 1927 -371 1928 -257
rect 1941 -258 1942 -254
rect 1983 -371 1984 -257
rect 44 -260 45 -254
rect 208 -260 209 -254
rect 240 -260 241 -254
rect 313 -260 314 -254
rect 338 -371 339 -259
rect 408 -260 409 -254
rect 432 -371 433 -259
rect 796 -371 797 -259
rect 828 -260 829 -254
rect 845 -371 846 -259
rect 880 -371 881 -259
rect 1528 -260 1529 -254
rect 1542 -260 1543 -254
rect 1605 -371 1606 -259
rect 1615 -371 1616 -259
rect 1661 -371 1662 -259
rect 1668 -260 1669 -254
rect 1731 -371 1732 -259
rect 1962 -371 1963 -259
rect 2193 -371 2194 -259
rect 23 -262 24 -254
rect 240 -371 241 -261
rect 247 -262 248 -254
rect 436 -262 437 -254
rect 439 -262 440 -254
rect 590 -262 591 -254
rect 653 -262 654 -254
rect 884 -371 885 -261
rect 891 -371 892 -261
rect 1640 -371 1641 -261
rect 23 -371 24 -263
rect 37 -264 38 -254
rect 54 -371 55 -263
rect 1507 -264 1508 -254
rect 1514 -264 1515 -254
rect 1843 -371 1844 -263
rect 37 -371 38 -265
rect 415 -266 416 -254
rect 422 -266 423 -254
rect 590 -371 591 -265
rect 709 -266 710 -254
rect 1031 -266 1032 -254
rect 1083 -371 1084 -265
rect 1689 -371 1690 -265
rect 65 -371 66 -267
rect 128 -268 129 -254
rect 149 -371 150 -267
rect 170 -268 171 -254
rect 187 -371 188 -267
rect 254 -268 255 -254
rect 268 -268 269 -254
rect 303 -268 304 -254
rect 310 -268 311 -254
rect 982 -268 983 -254
rect 996 -268 997 -254
rect 1829 -371 1830 -267
rect 86 -371 87 -269
rect 93 -270 94 -254
rect 114 -371 115 -269
rect 142 -270 143 -254
rect 156 -371 157 -269
rect 632 -270 633 -254
rect 709 -371 710 -269
rect 814 -270 815 -254
rect 828 -371 829 -269
rect 849 -270 850 -254
rect 856 -270 857 -254
rect 996 -371 997 -269
rect 1010 -270 1011 -254
rect 1780 -371 1781 -269
rect 58 -272 59 -254
rect 142 -371 143 -271
rect 233 -272 234 -254
rect 408 -371 409 -271
rect 422 -371 423 -271
rect 457 -272 458 -254
rect 506 -272 507 -254
rect 520 -371 521 -271
rect 534 -272 535 -254
rect 940 -272 941 -254
rect 954 -272 955 -254
rect 1031 -371 1032 -271
rect 1094 -272 1095 -254
rect 1549 -371 1550 -271
rect 1552 -272 1553 -254
rect 1766 -371 1767 -271
rect 58 -371 59 -273
rect 744 -274 745 -254
rect 772 -274 773 -254
rect 814 -371 815 -273
rect 856 -371 857 -273
rect 989 -371 990 -273
rect 1010 -371 1011 -273
rect 1017 -274 1018 -254
rect 1020 -371 1021 -273
rect 1451 -274 1452 -254
rect 1465 -274 1466 -254
rect 1794 -371 1795 -273
rect 93 -371 94 -275
rect 100 -276 101 -254
rect 128 -371 129 -275
rect 261 -276 262 -254
rect 268 -371 269 -275
rect 471 -276 472 -254
rect 506 -371 507 -275
rect 779 -276 780 -254
rect 863 -276 864 -254
rect 940 -371 941 -275
rect 954 -371 955 -275
rect 1003 -276 1004 -254
rect 1101 -276 1102 -254
rect 1199 -371 1200 -275
rect 1227 -276 1228 -254
rect 1647 -371 1648 -275
rect 100 -371 101 -277
rect 177 -278 178 -254
rect 205 -278 206 -254
rect 779 -371 780 -277
rect 842 -278 843 -254
rect 863 -371 864 -277
rect 894 -278 895 -254
rect 1535 -278 1536 -254
rect 1556 -278 1557 -254
rect 1654 -371 1655 -277
rect 72 -280 73 -254
rect 177 -371 178 -279
rect 191 -371 192 -279
rect 205 -371 206 -279
rect 219 -280 220 -254
rect 534 -371 535 -279
rect 555 -280 556 -254
rect 618 -371 619 -279
rect 628 -371 629 -279
rect 1003 -371 1004 -279
rect 1153 -280 1154 -254
rect 1710 -371 1711 -279
rect 72 -371 73 -281
rect 835 -282 836 -254
rect 926 -282 927 -254
rect 1094 -371 1095 -281
rect 1178 -282 1179 -254
rect 1514 -371 1515 -281
rect 1591 -282 1592 -254
rect 1815 -371 1816 -281
rect 107 -284 108 -254
rect 261 -371 262 -283
rect 275 -284 276 -254
rect 464 -284 465 -254
rect 471 -371 472 -283
rect 485 -284 486 -254
rect 513 -284 514 -254
rect 653 -371 654 -283
rect 667 -284 668 -254
rect 849 -371 850 -283
rect 947 -284 948 -254
rect 1227 -371 1228 -283
rect 1262 -284 1263 -254
rect 1752 -371 1753 -283
rect 107 -371 108 -285
rect 212 -286 213 -254
rect 219 -371 220 -285
rect 226 -286 227 -254
rect 233 -371 234 -285
rect 894 -371 895 -285
rect 947 -371 948 -285
rect 1545 -286 1546 -254
rect 1626 -286 1627 -254
rect 1717 -371 1718 -285
rect 135 -288 136 -254
rect 303 -371 304 -287
rect 310 -371 311 -287
rect 450 -288 451 -254
rect 548 -288 549 -254
rect 555 -371 556 -287
rect 569 -288 570 -254
rect 926 -371 927 -287
rect 968 -288 969 -254
rect 982 -371 983 -287
rect 1213 -288 1214 -254
rect 1535 -371 1536 -287
rect 1633 -288 1634 -254
rect 1745 -371 1746 -287
rect 30 -290 31 -254
rect 450 -371 451 -289
rect 548 -371 549 -289
rect 912 -290 913 -254
rect 1122 -290 1123 -254
rect 1213 -371 1214 -289
rect 1276 -290 1277 -254
rect 1507 -371 1508 -289
rect 30 -371 31 -291
rect 51 -292 52 -254
rect 138 -292 139 -254
rect 170 -371 171 -291
rect 226 -371 227 -291
rect 352 -292 353 -254
rect 394 -292 395 -254
rect 457 -371 458 -291
rect 611 -292 612 -254
rect 968 -371 969 -291
rect 975 -292 976 -254
rect 1122 -371 1123 -291
rect 1136 -292 1137 -254
rect 1276 -371 1277 -291
rect 1297 -292 1298 -254
rect 1528 -371 1529 -291
rect 47 -371 48 -293
rect 51 -371 52 -293
rect 138 -371 139 -293
rect 366 -371 367 -293
rect 394 -371 395 -293
rect 481 -371 482 -293
rect 611 -371 612 -293
rect 681 -294 682 -254
rect 702 -294 703 -254
rect 1262 -371 1263 -293
rect 1318 -294 1319 -254
rect 1556 -371 1557 -293
rect 89 -296 90 -254
rect 681 -371 682 -295
rect 688 -296 689 -254
rect 702 -371 703 -295
rect 723 -296 724 -254
rect 912 -371 913 -295
rect 919 -296 920 -254
rect 1318 -371 1319 -295
rect 1328 -371 1329 -295
rect 2004 -371 2005 -295
rect 243 -371 244 -297
rect 415 -371 416 -297
rect 429 -298 430 -254
rect 464 -371 465 -297
rect 576 -298 577 -254
rect 919 -371 920 -297
rect 1108 -298 1109 -254
rect 1297 -371 1298 -297
rect 1353 -298 1354 -254
rect 1626 -371 1627 -297
rect 247 -371 248 -299
rect 404 -371 405 -299
rect 576 -371 577 -299
rect 838 -371 839 -299
rect 1024 -300 1025 -254
rect 1108 -371 1109 -299
rect 1360 -300 1361 -254
rect 1738 -371 1739 -299
rect 254 -371 255 -301
rect 271 -302 272 -254
rect 275 -371 276 -301
rect 324 -302 325 -254
rect 345 -302 346 -254
rect 569 -371 570 -301
rect 597 -302 598 -254
rect 688 -371 689 -301
rect 723 -371 724 -301
rect 758 -302 759 -254
rect 772 -371 773 -301
rect 1591 -371 1592 -301
rect 282 -304 283 -254
rect 436 -371 437 -303
rect 660 -304 661 -254
rect 667 -371 668 -303
rect 730 -304 731 -254
rect 842 -371 843 -303
rect 1171 -304 1172 -254
rect 1360 -371 1361 -303
rect 1374 -304 1375 -254
rect 1822 -371 1823 -303
rect 135 -371 136 -305
rect 282 -371 283 -305
rect 289 -306 290 -254
rect 485 -371 486 -305
rect 660 -371 661 -305
rect 1325 -371 1326 -305
rect 1381 -306 1382 -254
rect 1465 -371 1466 -305
rect 1472 -306 1473 -254
rect 1787 -371 1788 -305
rect 289 -371 290 -307
rect 387 -308 388 -254
rect 401 -308 402 -254
rect 513 -371 514 -307
rect 716 -308 717 -254
rect 730 -371 731 -307
rect 786 -308 787 -254
rect 1136 -371 1137 -307
rect 1185 -308 1186 -254
rect 1374 -371 1375 -307
rect 1388 -308 1389 -254
rect 1619 -371 1620 -307
rect 296 -371 297 -309
rect 499 -310 500 -254
rect 646 -310 647 -254
rect 716 -371 717 -309
rect 786 -371 787 -309
rect 1027 -371 1028 -309
rect 1073 -310 1074 -254
rect 1171 -371 1172 -309
rect 1185 -371 1186 -309
rect 1332 -310 1333 -254
rect 1395 -310 1396 -254
rect 1682 -371 1683 -309
rect 212 -371 213 -311
rect 646 -371 647 -311
rect 1073 -371 1074 -311
rect 1269 -312 1270 -254
rect 1402 -312 1403 -254
rect 1668 -371 1669 -311
rect 299 -314 300 -254
rect 807 -314 808 -254
rect 1076 -371 1077 -313
rect 1395 -371 1396 -313
rect 1409 -314 1410 -254
rect 1675 -371 1676 -313
rect 324 -371 325 -315
rect 541 -316 542 -254
rect 1157 -316 1158 -254
rect 1269 -371 1270 -315
rect 1311 -316 1312 -254
rect 1402 -371 1403 -315
rect 1416 -316 1417 -254
rect 1696 -371 1697 -315
rect 331 -318 332 -254
rect 499 -371 500 -317
rect 933 -318 934 -254
rect 1416 -371 1417 -317
rect 1423 -318 1424 -254
rect 1759 -371 1760 -317
rect 331 -371 332 -319
rect 800 -371 801 -319
rect 870 -320 871 -254
rect 933 -371 934 -319
rect 1104 -371 1105 -319
rect 1311 -371 1312 -319
rect 1430 -320 1431 -254
rect 1724 -371 1725 -319
rect 345 -371 346 -321
rect 527 -322 528 -254
rect 632 -371 633 -321
rect 870 -371 871 -321
rect 1157 -371 1158 -321
rect 1255 -322 1256 -254
rect 1437 -322 1438 -254
rect 1703 -371 1704 -321
rect 79 -324 80 -254
rect 527 -371 528 -323
rect 712 -324 713 -254
rect 1255 -371 1256 -323
rect 1444 -324 1445 -254
rect 1773 -371 1774 -323
rect 79 -371 80 -325
rect 163 -326 164 -254
rect 352 -371 353 -325
rect 621 -326 622 -254
rect 1164 -326 1165 -254
rect 1332 -371 1333 -325
rect 1451 -371 1452 -325
rect 1612 -371 1613 -325
rect 163 -371 164 -327
rect 166 -371 167 -327
rect 359 -328 360 -254
rect 597 -371 598 -327
rect 1017 -371 1018 -327
rect 1164 -371 1165 -327
rect 1192 -328 1193 -254
rect 1388 -371 1389 -327
rect 1472 -371 1473 -327
rect 1584 -328 1585 -254
rect 359 -371 360 -329
rect 523 -330 524 -254
rect 1066 -330 1067 -254
rect 1192 -371 1193 -329
rect 1206 -330 1207 -254
rect 1423 -371 1424 -329
rect 1486 -330 1487 -254
rect 1836 -371 1837 -329
rect 117 -332 118 -254
rect 1066 -371 1067 -331
rect 1087 -332 1088 -254
rect 1206 -371 1207 -331
rect 1220 -332 1221 -254
rect 1430 -371 1431 -331
rect 1493 -332 1494 -254
rect 1633 -371 1634 -331
rect 380 -334 381 -254
rect 387 -371 388 -333
rect 443 -334 444 -254
rect 541 -371 542 -333
rect 961 -334 962 -254
rect 1087 -371 1088 -333
rect 1234 -334 1235 -254
rect 1409 -371 1410 -333
rect 1500 -334 1501 -254
rect 1808 -371 1809 -333
rect 373 -336 374 -254
rect 380 -371 381 -335
rect 443 -371 444 -335
rect 478 -336 479 -254
rect 765 -336 766 -254
rect 961 -371 962 -335
rect 1038 -336 1039 -254
rect 1220 -371 1221 -335
rect 1248 -336 1249 -254
rect 1437 -371 1438 -335
rect 1479 -336 1480 -254
rect 1500 -371 1501 -335
rect 1563 -336 1564 -254
rect 1584 -371 1585 -335
rect 373 -371 374 -337
rect 705 -338 706 -254
rect 1038 -371 1039 -337
rect 1150 -338 1151 -254
rect 1248 -371 1249 -337
rect 1577 -338 1578 -254
rect 478 -371 479 -339
rect 1542 -371 1543 -339
rect 639 -342 640 -254
rect 765 -371 766 -341
rect 1129 -342 1130 -254
rect 1234 -371 1235 -341
rect 1283 -342 1284 -254
rect 1493 -371 1494 -341
rect 639 -371 640 -343
rect 695 -344 696 -254
rect 1045 -344 1046 -254
rect 1283 -371 1284 -343
rect 1290 -344 1291 -254
rect 1444 -371 1445 -343
rect 695 -371 696 -345
rect 737 -346 738 -254
rect 877 -346 878 -254
rect 1045 -371 1046 -345
rect 1052 -346 1053 -254
rect 1129 -371 1130 -345
rect 1150 -371 1151 -345
rect 1570 -346 1571 -254
rect 604 -348 605 -254
rect 737 -371 738 -347
rect 877 -371 878 -347
rect 1381 -371 1382 -347
rect 1458 -348 1459 -254
rect 1570 -371 1571 -347
rect 317 -350 318 -254
rect 604 -371 605 -349
rect 625 -350 626 -254
rect 1458 -371 1459 -349
rect 121 -352 122 -254
rect 317 -371 318 -351
rect 401 -371 402 -351
rect 625 -371 626 -351
rect 898 -352 899 -254
rect 1052 -371 1053 -351
rect 1304 -352 1305 -254
rect 1479 -371 1480 -351
rect 121 -371 122 -353
rect 583 -354 584 -254
rect 898 -371 899 -353
rect 1143 -354 1144 -254
rect 1339 -354 1340 -254
rect 1563 -371 1564 -353
rect 492 -356 493 -254
rect 583 -371 584 -355
rect 1024 -371 1025 -355
rect 1290 -371 1291 -355
rect 1346 -356 1347 -254
rect 1577 -371 1578 -355
rect 492 -371 493 -357
rect 562 -358 563 -254
rect 821 -358 822 -254
rect 1346 -371 1347 -357
rect 1367 -358 1368 -254
rect 1486 -371 1487 -357
rect 184 -360 185 -254
rect 562 -371 563 -359
rect 751 -360 752 -254
rect 821 -371 822 -359
rect 1059 -360 1060 -254
rect 1143 -371 1144 -359
rect 1181 -371 1182 -359
rect 1367 -371 1368 -359
rect 674 -362 675 -254
rect 751 -371 752 -361
rect 905 -362 906 -254
rect 1059 -371 1060 -361
rect 1115 -362 1116 -254
rect 1304 -371 1305 -361
rect 467 -364 468 -254
rect 674 -371 675 -363
rect 793 -364 794 -254
rect 905 -371 906 -363
rect 1080 -364 1081 -254
rect 1115 -371 1116 -363
rect 1241 -364 1242 -254
rect 1339 -371 1340 -363
rect 793 -371 794 -365
rect 1521 -366 1522 -254
rect 835 -371 836 -367
rect 1521 -371 1522 -367
rect 887 -370 888 -254
rect 1241 -371 1242 -369
rect 16 -381 17 -379
rect 621 -500 622 -380
rect 625 -381 626 -379
rect 702 -381 703 -379
rect 758 -381 759 -379
rect 1297 -381 1298 -379
rect 1353 -381 1354 -379
rect 1948 -500 1949 -380
rect 1958 -500 1959 -380
rect 2116 -500 2117 -380
rect 2193 -381 2194 -379
rect 2284 -500 2285 -380
rect 23 -383 24 -379
rect 747 -383 748 -379
rect 751 -383 752 -379
rect 758 -500 759 -382
rect 761 -383 762 -379
rect 800 -500 801 -382
rect 810 -383 811 -379
rect 828 -383 829 -379
rect 845 -383 846 -379
rect 1752 -383 1753 -379
rect 1766 -383 1767 -379
rect 1962 -383 1963 -379
rect 1969 -383 1970 -379
rect 2088 -500 2089 -382
rect 23 -500 24 -384
rect 44 -385 45 -379
rect 51 -500 52 -384
rect 79 -385 80 -379
rect 96 -385 97 -379
rect 1178 -385 1179 -379
rect 1185 -385 1186 -379
rect 1297 -500 1298 -384
rect 1353 -500 1354 -384
rect 1472 -385 1473 -379
rect 1528 -385 1529 -379
rect 1528 -500 1529 -384
rect 1528 -385 1529 -379
rect 1528 -500 1529 -384
rect 1591 -385 1592 -379
rect 1752 -500 1753 -384
rect 1773 -385 1774 -379
rect 1899 -500 1900 -384
rect 1927 -385 1928 -379
rect 1997 -500 1998 -384
rect 2004 -385 2005 -379
rect 2263 -500 2264 -384
rect 37 -387 38 -379
rect 481 -387 482 -379
rect 495 -500 496 -386
rect 562 -387 563 -379
rect 600 -500 601 -386
rect 1136 -387 1137 -379
rect 1167 -500 1168 -386
rect 1682 -387 1683 -379
rect 1710 -387 1711 -379
rect 1850 -500 1851 -386
rect 1976 -500 1977 -386
rect 1990 -500 1991 -386
rect 2011 -500 2012 -386
rect 2144 -500 2145 -386
rect 44 -500 45 -388
rect 446 -389 447 -379
rect 478 -389 479 -379
rect 856 -389 857 -379
rect 971 -500 972 -388
rect 1759 -389 1760 -379
rect 1794 -389 1795 -379
rect 1906 -500 1907 -388
rect 1983 -389 1984 -379
rect 2039 -500 2040 -388
rect 61 -500 62 -390
rect 247 -391 248 -379
rect 345 -391 346 -379
rect 478 -500 479 -390
rect 499 -391 500 -379
rect 499 -500 500 -390
rect 499 -391 500 -379
rect 499 -500 500 -390
rect 513 -391 514 -379
rect 562 -500 563 -390
rect 625 -500 626 -390
rect 884 -391 885 -379
rect 978 -391 979 -379
rect 1346 -391 1347 -379
rect 1356 -391 1357 -379
rect 1430 -391 1431 -379
rect 1440 -500 1441 -390
rect 1983 -500 1984 -390
rect 65 -393 66 -379
rect 65 -500 66 -392
rect 65 -393 66 -379
rect 65 -500 66 -392
rect 72 -393 73 -379
rect 135 -500 136 -392
rect 163 -393 164 -379
rect 1801 -393 1802 -379
rect 1808 -393 1809 -379
rect 1913 -500 1914 -392
rect 16 -500 17 -394
rect 163 -500 164 -394
rect 170 -395 171 -379
rect 215 -500 216 -394
rect 222 -500 223 -394
rect 590 -395 591 -379
rect 635 -395 636 -379
rect 1591 -500 1592 -394
rect 1612 -395 1613 -379
rect 1941 -500 1942 -394
rect 72 -500 73 -396
rect 86 -397 87 -379
rect 173 -500 174 -396
rect 205 -397 206 -379
rect 233 -397 234 -379
rect 751 -500 752 -396
rect 765 -397 766 -379
rect 891 -397 892 -379
rect 978 -500 979 -396
rect 1087 -397 1088 -379
rect 1125 -500 1126 -396
rect 1857 -500 1858 -396
rect 30 -399 31 -379
rect 233 -500 234 -398
rect 247 -500 248 -398
rect 373 -399 374 -379
rect 401 -399 402 -379
rect 506 -399 507 -379
rect 513 -500 514 -398
rect 688 -399 689 -379
rect 702 -500 703 -398
rect 1006 -500 1007 -398
rect 1017 -399 1018 -379
rect 1780 -399 1781 -379
rect 1815 -399 1816 -379
rect 1920 -500 1921 -398
rect 79 -500 80 -400
rect 611 -401 612 -379
rect 646 -500 647 -400
rect 912 -401 913 -379
rect 982 -401 983 -379
rect 1104 -401 1105 -379
rect 1136 -500 1137 -400
rect 1248 -401 1249 -379
rect 1262 -401 1263 -379
rect 1346 -500 1347 -400
rect 1360 -401 1361 -379
rect 1430 -500 1431 -400
rect 1493 -401 1494 -379
rect 1612 -500 1613 -400
rect 1633 -401 1634 -379
rect 1759 -500 1760 -400
rect 1787 -401 1788 -379
rect 1815 -500 1816 -400
rect 1836 -401 1837 -379
rect 1934 -500 1935 -400
rect 86 -500 87 -402
rect 415 -403 416 -379
rect 443 -403 444 -379
rect 506 -500 507 -402
rect 527 -403 528 -379
rect 982 -500 983 -402
rect 1020 -403 1021 -379
rect 1325 -500 1326 -402
rect 1360 -500 1361 -402
rect 1542 -403 1543 -379
rect 1549 -403 1550 -379
rect 1633 -500 1634 -402
rect 1654 -403 1655 -379
rect 1864 -500 1865 -402
rect 121 -405 122 -379
rect 205 -500 206 -404
rect 212 -405 213 -379
rect 443 -500 444 -404
rect 527 -500 528 -404
rect 548 -405 549 -379
rect 667 -405 668 -379
rect 772 -405 773 -379
rect 793 -405 794 -379
rect 1738 -405 1739 -379
rect 1745 -405 1746 -379
rect 1892 -500 1893 -404
rect 114 -407 115 -379
rect 121 -500 122 -406
rect 156 -407 157 -379
rect 765 -500 766 -406
rect 849 -407 850 -379
rect 891 -500 892 -406
rect 1024 -500 1025 -406
rect 1773 -500 1774 -406
rect 1843 -407 1844 -379
rect 1969 -500 1970 -406
rect 156 -500 157 -408
rect 191 -409 192 -379
rect 219 -409 220 -379
rect 667 -500 668 -408
rect 674 -409 675 -379
rect 828 -500 829 -408
rect 852 -500 853 -408
rect 1122 -409 1123 -379
rect 1129 -409 1130 -379
rect 1248 -500 1249 -408
rect 1388 -409 1389 -379
rect 1472 -500 1473 -408
rect 1500 -409 1501 -379
rect 1843 -500 1844 -408
rect 149 -411 150 -379
rect 191 -500 192 -410
rect 226 -411 227 -379
rect 611 -500 612 -410
rect 674 -500 675 -410
rect 709 -411 710 -379
rect 716 -411 717 -379
rect 772 -500 773 -410
rect 856 -500 857 -410
rect 985 -500 986 -410
rect 1027 -411 1028 -379
rect 1962 -500 1963 -410
rect 149 -500 150 -412
rect 432 -413 433 -379
rect 541 -413 542 -379
rect 590 -500 591 -412
rect 653 -413 654 -379
rect 709 -500 710 -412
rect 730 -413 731 -379
rect 793 -500 794 -412
rect 863 -413 864 -379
rect 912 -500 913 -412
rect 1031 -413 1032 -379
rect 1087 -500 1088 -412
rect 1164 -413 1165 -379
rect 1542 -500 1543 -412
rect 1563 -413 1564 -379
rect 1654 -500 1655 -412
rect 1661 -413 1662 -379
rect 1780 -500 1781 -412
rect 187 -415 188 -379
rect 1766 -500 1767 -414
rect 226 -500 227 -416
rect 240 -417 241 -379
rect 345 -500 346 -416
rect 464 -417 465 -379
rect 541 -500 542 -416
rect 649 -417 650 -379
rect 653 -500 654 -416
rect 1479 -417 1480 -379
rect 1507 -417 1508 -379
rect 1549 -500 1550 -416
rect 1570 -417 1571 -379
rect 1801 -500 1802 -416
rect 240 -500 241 -418
rect 268 -419 269 -379
rect 359 -419 360 -379
rect 429 -419 430 -379
rect 548 -500 549 -418
rect 569 -419 570 -379
rect 681 -419 682 -379
rect 1017 -500 1018 -418
rect 1059 -419 1060 -379
rect 1129 -500 1130 -418
rect 1178 -500 1179 -418
rect 1290 -419 1291 -379
rect 1311 -419 1312 -379
rect 1388 -500 1389 -418
rect 1402 -419 1403 -379
rect 1493 -500 1494 -418
rect 1584 -419 1585 -379
rect 1710 -500 1711 -418
rect 1724 -419 1725 -379
rect 1878 -500 1879 -418
rect 166 -421 167 -379
rect 359 -500 360 -420
rect 373 -500 374 -420
rect 436 -421 437 -379
rect 471 -421 472 -379
rect 681 -500 682 -420
rect 688 -500 689 -420
rect 957 -500 958 -420
rect 968 -421 969 -379
rect 1031 -500 1032 -420
rect 1073 -421 1074 -379
rect 1871 -500 1872 -420
rect 100 -423 101 -379
rect 436 -500 437 -422
rect 457 -423 458 -379
rect 471 -500 472 -422
rect 730 -500 731 -422
rect 807 -423 808 -379
rect 1076 -423 1077 -379
rect 1647 -423 1648 -379
rect 1668 -423 1669 -379
rect 1787 -500 1788 -422
rect 100 -500 101 -424
rect 520 -425 521 -379
rect 744 -425 745 -379
rect 1262 -500 1263 -424
rect 1328 -425 1329 -379
rect 1668 -500 1669 -424
rect 1675 -425 1676 -379
rect 1794 -500 1795 -424
rect 166 -500 167 -426
rect 331 -427 332 -379
rect 401 -500 402 -426
rect 485 -427 486 -379
rect 737 -427 738 -379
rect 744 -500 745 -426
rect 779 -427 780 -379
rect 1073 -500 1074 -426
rect 1080 -427 1081 -379
rect 1227 -427 1228 -379
rect 1332 -427 1333 -379
rect 1402 -500 1403 -426
rect 1409 -427 1410 -379
rect 1500 -500 1501 -426
rect 1556 -427 1557 -379
rect 1675 -500 1676 -426
rect 1682 -500 1683 -426
rect 1829 -427 1830 -379
rect 212 -500 213 -428
rect 1059 -500 1060 -428
rect 1083 -429 1084 -379
rect 1661 -500 1662 -428
rect 1689 -429 1690 -379
rect 1808 -500 1809 -428
rect 268 -500 269 -430
rect 905 -431 906 -379
rect 968 -500 969 -430
rect 1647 -500 1648 -430
rect 1703 -431 1704 -379
rect 1836 -500 1837 -430
rect 296 -433 297 -379
rect 779 -500 780 -432
rect 803 -433 804 -379
rect 1332 -500 1333 -432
rect 1367 -433 1368 -379
rect 1479 -500 1480 -432
rect 1486 -433 1487 -379
rect 1584 -500 1585 -432
rect 1619 -433 1620 -379
rect 1738 -500 1739 -432
rect 296 -500 297 -434
rect 786 -435 787 -379
rect 807 -500 808 -434
rect 1122 -500 1123 -434
rect 1192 -435 1193 -379
rect 1290 -500 1291 -434
rect 1437 -435 1438 -379
rect 1507 -500 1508 -434
rect 1514 -435 1515 -379
rect 1619 -500 1620 -434
rect 1626 -435 1627 -379
rect 1745 -500 1746 -434
rect 303 -437 304 -379
rect 485 -500 486 -436
rect 632 -437 633 -379
rect 786 -500 787 -436
rect 842 -437 843 -379
rect 1409 -500 1410 -436
rect 1423 -437 1424 -379
rect 1514 -500 1515 -436
rect 1521 -437 1522 -379
rect 1626 -500 1627 -436
rect 1640 -437 1641 -379
rect 1724 -500 1725 -436
rect 1731 -437 1732 -379
rect 1885 -500 1886 -436
rect 177 -439 178 -379
rect 303 -500 304 -438
rect 310 -439 311 -379
rect 569 -500 570 -438
rect 632 -500 633 -438
rect 877 -439 878 -379
rect 887 -500 888 -438
rect 1640 -500 1641 -438
rect 1717 -439 1718 -379
rect 1829 -500 1830 -438
rect 177 -500 178 -440
rect 338 -441 339 -379
rect 408 -441 409 -379
rect 520 -500 521 -440
rect 719 -500 720 -440
rect 1423 -500 1424 -440
rect 1444 -441 1445 -379
rect 1521 -500 1522 -440
rect 1577 -441 1578 -379
rect 1689 -500 1690 -440
rect 107 -443 108 -379
rect 408 -500 409 -442
rect 415 -500 416 -442
rect 639 -443 640 -379
rect 775 -443 776 -379
rect 1444 -500 1445 -442
rect 1451 -443 1452 -379
rect 1577 -500 1578 -442
rect 1598 -443 1599 -379
rect 1717 -500 1718 -442
rect 107 -500 108 -444
rect 275 -445 276 -379
rect 310 -500 311 -444
rect 366 -445 367 -379
rect 429 -500 430 -444
rect 618 -445 619 -379
rect 814 -445 815 -379
rect 842 -500 843 -444
rect 870 -445 871 -379
rect 1227 -500 1228 -444
rect 1241 -445 1242 -379
rect 1556 -500 1557 -444
rect 1605 -445 1606 -379
rect 1731 -500 1732 -444
rect 2 -500 3 -446
rect 618 -500 619 -446
rect 821 -447 822 -379
rect 877 -500 878 -446
rect 905 -500 906 -446
rect 940 -447 941 -379
rect 1010 -447 1011 -379
rect 1241 -500 1242 -446
rect 1255 -447 1256 -379
rect 1451 -500 1452 -446
rect 1458 -447 1459 -379
rect 1605 -500 1606 -446
rect 58 -449 59 -379
rect 814 -500 815 -448
rect 870 -500 871 -448
rect 1080 -500 1081 -448
rect 1083 -500 1084 -448
rect 1395 -449 1396 -379
rect 1465 -449 1466 -379
rect 1570 -500 1571 -448
rect 128 -451 129 -379
rect 366 -500 367 -450
rect 450 -451 451 -379
rect 1703 -500 1704 -450
rect 128 -500 129 -452
rect 142 -453 143 -379
rect 198 -453 199 -379
rect 639 -500 640 -452
rect 695 -453 696 -379
rect 821 -500 822 -452
rect 940 -500 941 -452
rect 1150 -453 1151 -379
rect 1181 -453 1182 -379
rect 1458 -500 1459 -452
rect 1486 -500 1487 -452
rect 1822 -453 1823 -379
rect 142 -500 143 -454
rect 926 -455 927 -379
rect 1010 -500 1011 -454
rect 1038 -455 1039 -379
rect 1066 -455 1067 -379
rect 1192 -500 1193 -454
rect 1220 -455 1221 -379
rect 1311 -500 1312 -454
rect 1318 -455 1319 -379
rect 1465 -500 1466 -454
rect 1696 -455 1697 -379
rect 1822 -500 1823 -454
rect 184 -457 185 -379
rect 695 -500 696 -456
rect 726 -500 727 -456
rect 1255 -500 1256 -456
rect 1269 -457 1270 -379
rect 1395 -500 1396 -456
rect 1535 -457 1536 -379
rect 1696 -500 1697 -456
rect 184 -500 185 -458
rect 576 -459 577 -379
rect 1038 -500 1039 -458
rect 1052 -459 1053 -379
rect 1066 -500 1067 -458
rect 1955 -500 1956 -458
rect 198 -500 199 -460
rect 352 -461 353 -379
rect 450 -500 451 -460
rect 723 -461 724 -379
rect 898 -461 899 -379
rect 1052 -500 1053 -460
rect 1101 -461 1102 -379
rect 1598 -500 1599 -460
rect 219 -500 220 -462
rect 926 -500 927 -462
rect 1045 -463 1046 -379
rect 1101 -500 1102 -462
rect 1108 -463 1109 -379
rect 1150 -500 1151 -462
rect 1199 -463 1200 -379
rect 1269 -500 1270 -462
rect 1283 -463 1284 -379
rect 1367 -500 1368 -462
rect 1416 -463 1417 -379
rect 1535 -500 1536 -462
rect 275 -500 276 -464
rect 387 -465 388 -379
rect 576 -500 577 -464
rect 604 -465 605 -379
rect 723 -500 724 -464
rect 1374 -465 1375 -379
rect 289 -467 290 -379
rect 387 -500 388 -466
rect 583 -467 584 -379
rect 604 -500 605 -466
rect 849 -500 850 -466
rect 1283 -500 1284 -466
rect 1339 -467 1340 -379
rect 1416 -500 1417 -466
rect 282 -469 283 -379
rect 289 -500 290 -468
rect 317 -469 318 -379
rect 457 -500 458 -468
rect 583 -500 584 -468
rect 796 -469 797 -379
rect 898 -500 899 -468
rect 954 -469 955 -379
rect 961 -469 962 -379
rect 1108 -500 1109 -468
rect 1115 -469 1116 -379
rect 1220 -500 1221 -468
rect 1276 -469 1277 -379
rect 1339 -500 1340 -468
rect 1374 -500 1375 -468
rect 1381 -469 1382 -379
rect 254 -471 255 -379
rect 282 -500 283 -470
rect 317 -500 318 -470
rect 716 -500 717 -470
rect 740 -500 741 -470
rect 1115 -500 1116 -470
rect 1171 -471 1172 -379
rect 1199 -500 1200 -470
rect 1206 -471 1207 -379
rect 1318 -500 1319 -470
rect 254 -500 255 -472
rect 597 -473 598 -379
rect 863 -500 864 -472
rect 954 -500 955 -472
rect 992 -473 993 -379
rect 1171 -500 1172 -472
rect 1213 -473 1214 -379
rect 1276 -500 1277 -472
rect 1304 -473 1305 -379
rect 1381 -500 1382 -472
rect 324 -475 325 -379
rect 737 -500 738 -474
rect 919 -475 920 -379
rect 1045 -500 1046 -474
rect 1143 -475 1144 -379
rect 1206 -500 1207 -474
rect 1234 -475 1235 -379
rect 1304 -500 1305 -474
rect 324 -500 325 -476
rect 422 -477 423 -379
rect 464 -500 465 -476
rect 597 -500 598 -476
rect 919 -500 920 -476
rect 989 -477 990 -379
rect 1094 -477 1095 -379
rect 1143 -500 1144 -476
rect 1157 -477 1158 -379
rect 1234 -500 1235 -476
rect 331 -500 332 -478
rect 380 -479 381 -379
rect 422 -500 423 -478
rect 534 -479 535 -379
rect 947 -479 948 -379
rect 961 -500 962 -478
rect 975 -479 976 -379
rect 1213 -500 1214 -478
rect 93 -481 94 -379
rect 380 -500 381 -480
rect 933 -481 934 -379
rect 947 -500 948 -480
rect 989 -500 990 -480
rect 1927 -500 1928 -480
rect 93 -500 94 -482
rect 534 -500 535 -482
rect 933 -500 934 -482
rect 1563 -500 1564 -482
rect 338 -500 339 -484
rect 394 -485 395 -379
rect 996 -485 997 -379
rect 1094 -500 1095 -484
rect 261 -487 262 -379
rect 394 -500 395 -486
rect 835 -487 836 -379
rect 996 -500 997 -486
rect 1003 -487 1004 -379
rect 1157 -500 1158 -486
rect 261 -500 262 -488
rect 660 -489 661 -379
rect 54 -491 55 -379
rect 660 -500 661 -490
rect 352 -500 353 -492
rect 1027 -500 1028 -492
rect 555 -495 556 -379
rect 835 -500 836 -494
rect 492 -497 493 -379
rect 555 -500 556 -496
rect 492 -500 493 -498
rect 1185 -500 1186 -498
rect 30 -633 31 -509
rect 72 -510 73 -508
rect 93 -510 94 -508
rect 173 -510 174 -508
rect 205 -510 206 -508
rect 733 -633 734 -509
rect 737 -510 738 -508
rect 1633 -510 1634 -508
rect 1682 -510 1683 -508
rect 2151 -633 2152 -509
rect 2214 -633 2215 -509
rect 2291 -633 2292 -509
rect 37 -633 38 -511
rect 646 -512 647 -508
rect 656 -512 657 -508
rect 695 -512 696 -508
rect 723 -512 724 -508
rect 772 -512 773 -508
rect 814 -512 815 -508
rect 814 -633 815 -511
rect 814 -512 815 -508
rect 814 -633 815 -511
rect 824 -633 825 -511
rect 1129 -512 1130 -508
rect 1146 -633 1147 -511
rect 1374 -512 1375 -508
rect 1535 -512 1536 -508
rect 2032 -633 2033 -511
rect 2039 -512 2040 -508
rect 2172 -633 2173 -511
rect 2263 -512 2264 -508
rect 2361 -633 2362 -511
rect 44 -514 45 -508
rect 212 -633 213 -513
rect 215 -514 216 -508
rect 1766 -514 1767 -508
rect 1836 -514 1837 -508
rect 2004 -633 2005 -513
rect 2014 -514 2015 -508
rect 2179 -633 2180 -513
rect 2284 -514 2285 -508
rect 2326 -633 2327 -513
rect 44 -633 45 -515
rect 166 -516 167 -508
rect 170 -516 171 -508
rect 450 -516 451 -508
rect 541 -516 542 -508
rect 632 -633 633 -515
rect 635 -516 636 -508
rect 772 -633 773 -515
rect 842 -516 843 -508
rect 884 -633 885 -515
rect 898 -516 899 -508
rect 968 -516 969 -508
rect 982 -516 983 -508
rect 1752 -516 1753 -508
rect 1864 -516 1865 -508
rect 2046 -633 2047 -515
rect 2088 -516 2089 -508
rect 2210 -633 2211 -515
rect 128 -518 129 -508
rect 128 -633 129 -517
rect 128 -518 129 -508
rect 128 -633 129 -517
rect 135 -518 136 -508
rect 737 -633 738 -517
rect 751 -518 752 -508
rect 754 -564 755 -517
rect 786 -518 787 -508
rect 842 -633 843 -517
rect 849 -518 850 -508
rect 919 -518 920 -508
rect 975 -518 976 -508
rect 1752 -633 1753 -517
rect 1864 -633 1865 -517
rect 1979 -518 1980 -508
rect 1983 -518 1984 -508
rect 2158 -633 2159 -517
rect 75 -633 76 -519
rect 919 -633 920 -519
rect 985 -520 986 -508
rect 1766 -633 1767 -519
rect 1794 -520 1795 -508
rect 1983 -633 1984 -519
rect 1990 -520 1991 -508
rect 2007 -520 2008 -508
rect 2116 -520 2117 -508
rect 2193 -633 2194 -519
rect 114 -522 115 -508
rect 975 -633 976 -521
rect 992 -522 993 -508
rect 1213 -522 1214 -508
rect 1269 -522 1270 -508
rect 1374 -633 1375 -521
rect 1472 -522 1473 -508
rect 1535 -633 1536 -521
rect 1612 -522 1613 -508
rect 1794 -633 1795 -521
rect 1808 -522 1809 -508
rect 1990 -633 1991 -521
rect 2116 -633 2117 -521
rect 2224 -633 2225 -521
rect 114 -633 115 -523
rect 331 -524 332 -508
rect 380 -524 381 -508
rect 989 -524 990 -508
rect 996 -524 997 -508
rect 1125 -524 1126 -508
rect 1164 -524 1165 -508
rect 2137 -633 2138 -523
rect 2144 -524 2145 -508
rect 2200 -633 2201 -523
rect 138 -633 139 -525
rect 898 -633 899 -525
rect 940 -526 941 -508
rect 996 -633 997 -525
rect 1003 -526 1004 -508
rect 1843 -526 1844 -508
rect 1871 -526 1872 -508
rect 2053 -633 2054 -525
rect 163 -633 164 -527
rect 716 -528 717 -508
rect 723 -633 724 -527
rect 1108 -528 1109 -508
rect 1167 -528 1168 -508
rect 1360 -528 1361 -508
rect 1395 -528 1396 -508
rect 1472 -633 1473 -527
rect 1619 -528 1620 -508
rect 1808 -633 1809 -527
rect 1878 -528 1879 -508
rect 2060 -633 2061 -527
rect 205 -633 206 -529
rect 1262 -530 1263 -508
rect 1290 -530 1291 -508
rect 1395 -633 1396 -529
rect 1479 -530 1480 -508
rect 1619 -633 1620 -529
rect 1633 -633 1634 -529
rect 2207 -633 2208 -529
rect 219 -532 220 -508
rect 2081 -633 2082 -531
rect 219 -633 220 -533
rect 653 -534 654 -508
rect 660 -534 661 -508
rect 1006 -534 1007 -508
rect 1017 -534 1018 -508
rect 1108 -633 1109 -533
rect 1192 -534 1193 -508
rect 1269 -633 1270 -533
rect 1290 -633 1291 -533
rect 1367 -534 1368 -508
rect 1479 -633 1480 -533
rect 2021 -534 2022 -508
rect 79 -536 80 -508
rect 653 -633 654 -535
rect 702 -536 703 -508
rect 1003 -633 1004 -535
rect 1024 -633 1025 -535
rect 1346 -536 1347 -508
rect 1367 -633 1368 -535
rect 1486 -536 1487 -508
rect 1640 -536 1641 -508
rect 1836 -633 1837 -535
rect 1885 -536 1886 -508
rect 2067 -633 2068 -535
rect 222 -538 223 -508
rect 282 -538 283 -508
rect 296 -538 297 -508
rect 296 -633 297 -537
rect 296 -538 297 -508
rect 296 -633 297 -537
rect 310 -538 311 -508
rect 663 -633 664 -537
rect 716 -633 717 -537
rect 726 -538 727 -508
rect 730 -538 731 -508
rect 989 -633 990 -537
rect 1031 -538 1032 -508
rect 1122 -633 1123 -537
rect 1136 -538 1137 -508
rect 1192 -633 1193 -537
rect 1227 -538 1228 -508
rect 1346 -633 1347 -537
rect 1493 -538 1494 -508
rect 1640 -633 1641 -537
rect 1661 -538 1662 -508
rect 2039 -633 2040 -537
rect 103 -633 104 -539
rect 1493 -633 1494 -539
rect 1710 -540 1711 -508
rect 1871 -633 1872 -539
rect 1892 -540 1893 -508
rect 1892 -633 1893 -539
rect 1892 -540 1893 -508
rect 1892 -633 1893 -539
rect 1899 -540 1900 -508
rect 2074 -633 2075 -539
rect 226 -542 227 -508
rect 236 -542 237 -508
rect 240 -542 241 -508
rect 310 -633 311 -541
rect 324 -542 325 -508
rect 492 -542 493 -508
rect 534 -542 535 -508
rect 1213 -633 1214 -541
rect 1255 -542 1256 -508
rect 1360 -633 1361 -541
rect 1717 -542 1718 -508
rect 1878 -633 1879 -541
rect 1906 -542 1907 -508
rect 2109 -633 2110 -541
rect 65 -544 66 -508
rect 226 -633 227 -543
rect 233 -544 234 -508
rect 1717 -633 1718 -543
rect 1731 -544 1732 -508
rect 2102 -633 2103 -543
rect 9 -546 10 -508
rect 65 -633 66 -545
rect 72 -633 73 -545
rect 240 -633 241 -545
rect 254 -546 255 -508
rect 597 -633 598 -545
rect 600 -546 601 -508
rect 1437 -546 1438 -508
rect 1570 -546 1571 -508
rect 1731 -633 1732 -545
rect 1738 -546 1739 -508
rect 1899 -633 1900 -545
rect 1913 -546 1914 -508
rect 2130 -633 2131 -545
rect 9 -633 10 -547
rect 198 -548 199 -508
rect 233 -633 234 -547
rect 429 -548 430 -508
rect 450 -633 451 -547
rect 513 -548 514 -508
rect 541 -633 542 -547
rect 740 -548 741 -508
rect 751 -633 752 -547
rect 905 -548 906 -508
rect 947 -548 948 -508
rect 1017 -633 1018 -547
rect 1034 -633 1035 -547
rect 1934 -548 1935 -508
rect 1941 -548 1942 -508
rect 2095 -633 2096 -547
rect 107 -550 108 -508
rect 198 -633 199 -549
rect 282 -633 283 -549
rect 387 -550 388 -508
rect 394 -550 395 -508
rect 1013 -633 1014 -549
rect 1062 -633 1063 -549
rect 2025 -633 2026 -549
rect 16 -552 17 -508
rect 107 -633 108 -551
rect 177 -552 178 -508
rect 254 -633 255 -551
rect 317 -552 318 -508
rect 324 -633 325 -551
rect 331 -633 332 -551
rect 537 -552 538 -508
rect 565 -633 566 -551
rect 1241 -552 1242 -508
rect 1262 -633 1263 -551
rect 1955 -552 1956 -508
rect 1962 -552 1963 -508
rect 2123 -633 2124 -551
rect 16 -633 17 -553
rect 156 -554 157 -508
rect 177 -633 178 -553
rect 887 -554 888 -508
rect 891 -554 892 -508
rect 968 -633 969 -553
rect 978 -554 979 -508
rect 1738 -633 1739 -553
rect 1759 -554 1760 -508
rect 1941 -633 1942 -553
rect 1948 -554 1949 -508
rect 2165 -633 2166 -553
rect 93 -633 94 -555
rect 537 -633 538 -555
rect 569 -556 570 -508
rect 593 -633 594 -555
rect 611 -556 612 -508
rect 702 -633 703 -555
rect 786 -633 787 -555
rect 1612 -633 1613 -555
rect 1675 -556 1676 -508
rect 1906 -633 1907 -555
rect 1920 -556 1921 -508
rect 1955 -633 1956 -555
rect 1969 -556 1970 -508
rect 2144 -633 2145 -555
rect 121 -558 122 -508
rect 156 -633 157 -557
rect 303 -558 304 -508
rect 317 -633 318 -557
rect 345 -558 346 -508
rect 429 -633 430 -557
rect 492 -633 493 -557
rect 562 -558 563 -508
rect 569 -633 570 -557
rect 744 -558 745 -508
rect 835 -558 836 -508
rect 891 -633 892 -557
rect 905 -633 906 -557
rect 961 -558 962 -508
rect 1031 -633 1032 -557
rect 1241 -633 1242 -557
rect 1283 -558 1284 -508
rect 1570 -633 1571 -557
rect 1591 -558 1592 -508
rect 1759 -633 1760 -557
rect 1773 -558 1774 -508
rect 1948 -633 1949 -557
rect 1976 -558 1977 -508
rect 1997 -558 1998 -508
rect 121 -633 122 -559
rect 548 -560 549 -508
rect 604 -560 605 -508
rect 611 -633 612 -559
rect 621 -560 622 -508
rect 870 -560 871 -508
rect 877 -560 878 -508
rect 1227 -633 1228 -559
rect 1297 -560 1298 -508
rect 1591 -633 1592 -559
rect 1696 -560 1697 -508
rect 1934 -633 1935 -559
rect 100 -562 101 -508
rect 548 -633 549 -561
rect 649 -633 650 -561
rect 1843 -633 1844 -561
rect 1927 -562 1928 -508
rect 2088 -633 2089 -561
rect 100 -633 101 -563
rect 639 -564 640 -508
rect 688 -564 689 -508
rect 730 -633 731 -563
rect 961 -633 962 -563
rect 985 -633 986 -563
rect 1696 -633 1697 -563
rect 1703 -564 1704 -508
rect 1927 -633 1928 -563
rect 61 -566 62 -508
rect 688 -633 689 -565
rect 793 -566 794 -508
rect 870 -633 871 -565
rect 1073 -566 1074 -508
rect 1129 -633 1130 -565
rect 1150 -566 1151 -508
rect 1255 -633 1256 -565
rect 1297 -633 1298 -565
rect 1801 -566 1802 -508
rect 1829 -566 1830 -508
rect 1885 -633 1886 -565
rect 2 -568 3 -508
rect 61 -633 62 -567
rect 303 -633 304 -567
rect 527 -568 528 -508
rect 639 -633 640 -567
rect 709 -568 710 -508
rect 793 -633 794 -567
rect 828 -568 829 -508
rect 852 -633 853 -567
rect 1038 -568 1039 -508
rect 1080 -568 1081 -508
rect 1710 -633 1711 -567
rect 1724 -568 1725 -508
rect 1962 -633 1963 -567
rect 250 -633 251 -569
rect 1038 -633 1039 -569
rect 1083 -570 1084 -508
rect 1787 -570 1788 -508
rect 338 -572 339 -508
rect 345 -633 346 -571
rect 366 -572 367 -508
rect 380 -633 381 -571
rect 387 -633 388 -571
rect 432 -633 433 -571
rect 436 -572 437 -508
rect 604 -633 605 -571
rect 709 -633 710 -571
rect 758 -572 759 -508
rect 765 -572 766 -508
rect 828 -633 829 -571
rect 863 -572 864 -508
rect 947 -633 948 -571
rect 971 -572 972 -508
rect 1724 -633 1725 -571
rect 1745 -572 1746 -508
rect 1920 -633 1921 -571
rect 142 -574 143 -508
rect 765 -633 766 -573
rect 821 -574 822 -508
rect 835 -633 836 -573
rect 863 -633 864 -573
rect 1647 -574 1648 -508
rect 1703 -633 1704 -573
rect 1822 -574 1823 -508
rect 142 -633 143 -575
rect 401 -576 402 -508
rect 408 -576 409 -508
rect 513 -633 514 -575
rect 527 -633 528 -575
rect 555 -576 556 -508
rect 695 -633 696 -575
rect 821 -633 822 -575
rect 954 -576 955 -508
rect 1745 -633 1746 -575
rect 1780 -576 1781 -508
rect 1969 -633 1970 -575
rect 117 -578 118 -508
rect 401 -633 402 -577
rect 415 -578 416 -508
rect 810 -633 811 -577
rect 856 -578 857 -508
rect 954 -633 955 -577
rect 1010 -578 1011 -508
rect 1073 -633 1074 -577
rect 1094 -578 1095 -508
rect 1164 -633 1165 -577
rect 1216 -633 1217 -577
rect 1997 -633 1998 -577
rect 275 -580 276 -508
rect 408 -633 409 -579
rect 422 -580 423 -508
rect 436 -633 437 -579
rect 495 -580 496 -508
rect 744 -633 745 -579
rect 758 -633 759 -579
rect 779 -580 780 -508
rect 800 -580 801 -508
rect 856 -633 857 -579
rect 1010 -633 1011 -579
rect 1976 -633 1977 -579
rect 86 -582 87 -508
rect 800 -633 801 -581
rect 1094 -633 1095 -581
rect 1682 -633 1683 -581
rect 86 -633 87 -583
rect 352 -584 353 -508
rect 359 -584 360 -508
rect 422 -633 423 -583
rect 506 -584 507 -508
rect 562 -633 563 -583
rect 586 -633 587 -583
rect 1780 -633 1781 -583
rect 58 -633 59 -585
rect 352 -633 353 -585
rect 359 -633 360 -585
rect 478 -586 479 -508
rect 555 -633 556 -585
rect 681 -586 682 -508
rect 1101 -586 1102 -508
rect 1136 -633 1137 -585
rect 1220 -586 1221 -508
rect 1283 -633 1284 -585
rect 1325 -586 1326 -508
rect 1661 -633 1662 -585
rect 23 -588 24 -508
rect 1325 -633 1326 -587
rect 1332 -588 1333 -508
rect 2011 -588 2012 -508
rect 23 -633 24 -589
rect 51 -590 52 -508
rect 275 -633 276 -589
rect 457 -590 458 -508
rect 471 -590 472 -508
rect 506 -633 507 -589
rect 674 -590 675 -508
rect 779 -633 780 -589
rect 1080 -633 1081 -589
rect 1101 -633 1102 -589
rect 1199 -590 1200 -508
rect 1220 -633 1221 -589
rect 1234 -590 1235 -508
rect 1332 -633 1333 -589
rect 1353 -590 1354 -508
rect 1437 -633 1438 -589
rect 1465 -590 1466 -508
rect 1913 -633 1914 -589
rect 51 -633 52 -591
rect 625 -592 626 -508
rect 667 -592 668 -508
rect 674 -633 675 -591
rect 681 -633 682 -591
rect 1150 -633 1151 -591
rect 1248 -592 1249 -508
rect 1353 -633 1354 -591
rect 1416 -592 1417 -508
rect 1773 -633 1774 -591
rect 1850 -592 1851 -508
rect 2011 -633 2012 -591
rect 135 -633 136 -593
rect 457 -633 458 -593
rect 464 -594 465 -508
rect 625 -633 626 -593
rect 1157 -594 1158 -508
rect 1248 -633 1249 -593
rect 1318 -594 1319 -508
rect 1465 -633 1466 -593
rect 1500 -594 1501 -508
rect 1647 -633 1648 -593
rect 184 -596 185 -508
rect 464 -633 465 -595
rect 576 -596 577 -508
rect 667 -633 668 -595
rect 1087 -596 1088 -508
rect 1157 -633 1158 -595
rect 1311 -596 1312 -508
rect 1318 -633 1319 -595
rect 1402 -596 1403 -508
rect 1500 -633 1501 -595
rect 1521 -596 1522 -508
rect 1675 -633 1676 -595
rect 184 -633 185 -597
rect 261 -598 262 -508
rect 289 -598 290 -508
rect 471 -633 472 -597
rect 576 -633 577 -597
rect 590 -598 591 -508
rect 618 -598 619 -508
rect 1234 -633 1235 -597
rect 1304 -598 1305 -508
rect 1402 -633 1403 -597
rect 1416 -633 1417 -597
rect 2018 -598 2019 -508
rect 149 -600 150 -508
rect 261 -633 262 -599
rect 289 -633 290 -599
rect 933 -600 934 -508
rect 1206 -600 1207 -508
rect 1311 -633 1312 -599
rect 1430 -600 1431 -508
rect 1521 -633 1522 -599
rect 1528 -600 1529 -508
rect 1829 -633 1830 -599
rect 1857 -600 1858 -508
rect 2018 -633 2019 -599
rect 149 -633 150 -601
rect 247 -602 248 -508
rect 338 -633 339 -601
rect 940 -633 941 -601
rect 1115 -602 1116 -508
rect 1206 -633 1207 -601
rect 1440 -602 1441 -508
rect 1850 -633 1851 -601
rect 79 -633 80 -603
rect 247 -633 248 -603
rect 366 -633 367 -603
rect 849 -633 850 -603
rect 912 -604 913 -508
rect 1304 -633 1305 -603
rect 1528 -633 1529 -603
rect 1577 -604 1578 -508
rect 1598 -604 1599 -508
rect 1787 -633 1788 -603
rect 373 -606 374 -508
rect 478 -633 479 -605
rect 590 -633 591 -605
rect 877 -633 878 -605
rect 929 -633 930 -605
rect 1087 -633 1088 -605
rect 1178 -606 1179 -508
rect 1430 -633 1431 -605
rect 1458 -606 1459 -508
rect 1598 -633 1599 -605
rect 1605 -606 1606 -508
rect 1822 -633 1823 -605
rect 191 -608 192 -508
rect 373 -633 374 -607
rect 394 -633 395 -607
rect 499 -608 500 -508
rect 807 -608 808 -508
rect 912 -633 913 -607
rect 933 -633 934 -607
rect 936 -608 937 -508
rect 1045 -608 1046 -508
rect 1115 -633 1116 -607
rect 1143 -608 1144 -508
rect 1178 -633 1179 -607
rect 1388 -608 1389 -508
rect 1458 -633 1459 -607
rect 1507 -608 1508 -508
rect 1577 -633 1578 -607
rect 1668 -608 1669 -508
rect 1857 -633 1858 -607
rect 173 -633 174 -609
rect 191 -633 192 -609
rect 443 -610 444 -508
rect 618 -633 619 -609
rect 926 -610 927 -508
rect 1045 -633 1046 -609
rect 1143 -633 1144 -609
rect 1815 -610 1816 -508
rect 443 -633 444 -611
rect 520 -612 521 -508
rect 926 -633 927 -611
rect 1542 -612 1543 -508
rect 1549 -612 1550 -508
rect 1801 -633 1802 -611
rect 485 -614 486 -508
rect 520 -633 521 -613
rect 1202 -633 1203 -613
rect 1542 -633 1543 -613
rect 1626 -614 1627 -508
rect 1815 -633 1816 -613
rect 485 -633 486 -615
rect 583 -616 584 -508
rect 1276 -616 1277 -508
rect 1388 -633 1389 -615
rect 1423 -616 1424 -508
rect 1605 -633 1606 -615
rect 1668 -633 1669 -615
rect 1689 -616 1690 -508
rect 499 -633 500 -617
rect 660 -633 661 -617
rect 1185 -618 1186 -508
rect 1276 -633 1277 -617
rect 1339 -618 1340 -508
rect 1423 -633 1424 -617
rect 1444 -618 1445 -508
rect 1549 -633 1550 -617
rect 1556 -618 1557 -508
rect 1689 -633 1690 -617
rect 583 -633 584 -619
rect 1654 -620 1655 -508
rect 1059 -622 1060 -508
rect 1185 -633 1186 -621
rect 1381 -622 1382 -508
rect 1444 -633 1445 -621
rect 1451 -622 1452 -508
rect 1626 -633 1627 -621
rect 1059 -633 1060 -623
rect 2186 -633 2187 -623
rect 1066 -626 1067 -508
rect 1451 -633 1452 -625
rect 1507 -633 1508 -625
rect 1514 -626 1515 -508
rect 1556 -633 1557 -625
rect 1563 -626 1564 -508
rect 1584 -626 1585 -508
rect 1654 -633 1655 -625
rect 1052 -628 1053 -508
rect 1066 -633 1067 -627
rect 1171 -628 1172 -508
rect 1339 -633 1340 -627
rect 1409 -628 1410 -508
rect 1514 -633 1515 -627
rect 1563 -633 1564 -627
rect 2221 -633 2222 -627
rect 268 -630 269 -508
rect 1052 -633 1053 -629
rect 1199 -633 1200 -629
rect 1381 -633 1382 -629
rect 1409 -633 1410 -629
rect 1958 -630 1959 -508
rect 268 -633 269 -631
rect 415 -633 416 -631
rect 915 -632 916 -508
rect 1171 -633 1172 -631
rect 1489 -633 1490 -631
rect 1584 -633 1585 -631
rect 2 -810 3 -642
rect 121 -643 122 -641
rect 131 -810 132 -642
rect 2137 -643 2138 -641
rect 2144 -643 2145 -641
rect 2319 -810 2320 -642
rect 2326 -643 2327 -641
rect 2347 -810 2348 -642
rect 2361 -643 2362 -641
rect 2403 -810 2404 -642
rect 44 -645 45 -641
rect 1223 -810 1224 -644
rect 1300 -645 1301 -641
rect 2130 -645 2131 -641
rect 2137 -810 2138 -644
rect 2172 -645 2173 -641
rect 2193 -645 2194 -641
rect 2207 -645 2208 -641
rect 2214 -645 2215 -641
rect 2277 -810 2278 -644
rect 2291 -645 2292 -641
rect 2326 -810 2327 -644
rect 47 -810 48 -646
rect 65 -647 66 -641
rect 68 -810 69 -646
rect 754 -810 755 -646
rect 807 -647 808 -641
rect 1122 -647 1123 -641
rect 1143 -647 1144 -641
rect 1591 -647 1592 -641
rect 1703 -647 1704 -641
rect 2235 -810 2236 -646
rect 12 -810 13 -648
rect 65 -810 66 -648
rect 72 -649 73 -641
rect 1780 -649 1781 -641
rect 1843 -649 1844 -641
rect 2221 -810 2222 -648
rect 51 -651 52 -641
rect 926 -651 927 -641
rect 940 -651 941 -641
rect 1906 -651 1907 -641
rect 1955 -651 1956 -641
rect 2256 -810 2257 -650
rect 51 -810 52 -652
rect 681 -653 682 -641
rect 698 -810 699 -652
rect 982 -810 983 -652
rect 1010 -653 1011 -641
rect 2151 -653 2152 -641
rect 2158 -653 2159 -641
rect 2312 -810 2313 -652
rect 58 -655 59 -641
rect 1682 -655 1683 -641
rect 1885 -655 1886 -641
rect 2130 -810 2131 -654
rect 2200 -655 2201 -641
rect 2224 -655 2225 -641
rect 72 -810 73 -656
rect 1003 -657 1004 -641
rect 1059 -657 1060 -641
rect 1626 -657 1627 -641
rect 1885 -810 1886 -656
rect 1969 -657 1970 -641
rect 2004 -657 2005 -641
rect 2144 -810 2145 -656
rect 82 -810 83 -658
rect 1031 -659 1032 -641
rect 1059 -810 1060 -658
rect 1073 -659 1074 -641
rect 1083 -659 1084 -641
rect 1465 -659 1466 -641
rect 1486 -659 1487 -641
rect 2165 -659 2166 -641
rect 16 -661 17 -641
rect 1073 -810 1074 -660
rect 1094 -661 1095 -641
rect 2186 -661 2187 -641
rect 93 -663 94 -641
rect 562 -663 563 -641
rect 618 -663 619 -641
rect 940 -810 941 -662
rect 957 -810 958 -662
rect 1052 -663 1053 -641
rect 1062 -663 1063 -641
rect 2179 -663 2180 -641
rect 93 -810 94 -664
rect 142 -665 143 -641
rect 145 -810 146 -664
rect 943 -665 944 -641
rect 1052 -810 1053 -664
rect 1108 -665 1109 -641
rect 1150 -665 1151 -641
rect 2186 -810 2187 -664
rect 75 -667 76 -641
rect 1108 -810 1109 -666
rect 1136 -667 1137 -641
rect 1150 -810 1151 -666
rect 1174 -810 1175 -666
rect 2305 -810 2306 -666
rect 135 -669 136 -641
rect 1822 -669 1823 -641
rect 1857 -669 1858 -641
rect 2004 -810 2005 -668
rect 2011 -669 2012 -641
rect 2151 -810 2152 -668
rect 170 -810 171 -670
rect 310 -671 311 -641
rect 401 -671 402 -641
rect 1031 -810 1032 -670
rect 1101 -671 1102 -641
rect 1122 -810 1123 -670
rect 1178 -671 1179 -641
rect 1213 -671 1214 -641
rect 1216 -671 1217 -641
rect 2109 -671 2110 -641
rect 2116 -671 2117 -641
rect 2298 -810 2299 -670
rect 173 -673 174 -641
rect 1927 -673 1928 -641
rect 1983 -673 1984 -641
rect 2109 -810 2110 -672
rect 2123 -673 2124 -641
rect 2291 -810 2292 -672
rect 187 -810 188 -674
rect 702 -675 703 -641
rect 733 -675 734 -641
rect 2179 -810 2180 -674
rect 205 -677 206 -641
rect 1451 -677 1452 -641
rect 1493 -677 1494 -641
rect 1626 -810 1627 -676
rect 1717 -677 1718 -641
rect 1822 -810 1823 -676
rect 1864 -677 1865 -641
rect 2011 -810 2012 -676
rect 2018 -677 2019 -641
rect 2158 -810 2159 -676
rect 212 -679 213 -641
rect 747 -679 748 -641
rect 765 -679 766 -641
rect 1003 -810 1004 -678
rect 1101 -810 1102 -678
rect 1111 -810 1112 -678
rect 1199 -679 1200 -641
rect 1983 -810 1984 -678
rect 1990 -679 1991 -641
rect 2123 -810 2124 -678
rect 191 -681 192 -641
rect 212 -810 213 -680
rect 236 -810 237 -680
rect 1178 -810 1179 -680
rect 1213 -810 1214 -680
rect 1409 -681 1410 -641
rect 1430 -681 1431 -641
rect 1591 -810 1592 -680
rect 1605 -681 1606 -641
rect 1717 -810 1718 -680
rect 1738 -681 1739 -641
rect 1857 -810 1858 -680
rect 1892 -681 1893 -641
rect 1892 -810 1893 -680
rect 1892 -681 1893 -641
rect 1892 -810 1893 -680
rect 1990 -810 1991 -680
rect 2067 -681 2068 -641
rect 2074 -681 2075 -641
rect 2242 -810 2243 -680
rect 149 -683 150 -641
rect 191 -810 192 -682
rect 247 -810 248 -682
rect 317 -683 318 -641
rect 366 -683 367 -641
rect 765 -810 766 -682
rect 800 -683 801 -641
rect 807 -810 808 -682
rect 824 -683 825 -641
rect 2284 -810 2285 -682
rect 30 -685 31 -641
rect 317 -810 318 -684
rect 366 -810 367 -684
rect 772 -685 773 -641
rect 849 -685 850 -641
rect 863 -685 864 -641
rect 891 -685 892 -641
rect 926 -810 927 -684
rect 929 -685 930 -641
rect 1955 -810 1956 -684
rect 1962 -685 1963 -641
rect 2067 -810 2068 -684
rect 2081 -685 2082 -641
rect 2249 -810 2250 -684
rect 9 -687 10 -641
rect 863 -810 864 -686
rect 877 -687 878 -641
rect 891 -810 892 -686
rect 1080 -687 1081 -641
rect 1738 -810 1739 -686
rect 1752 -687 1753 -641
rect 2074 -810 2075 -686
rect 2088 -687 2089 -641
rect 2263 -810 2264 -686
rect 19 -810 20 -688
rect 2081 -810 2082 -688
rect 2095 -689 2096 -641
rect 2270 -810 2271 -688
rect 30 -810 31 -690
rect 37 -691 38 -641
rect 149 -810 150 -690
rect 985 -691 986 -641
rect 1080 -810 1081 -690
rect 1087 -691 1088 -641
rect 1129 -691 1130 -641
rect 1199 -810 1200 -690
rect 1360 -691 1361 -641
rect 1451 -810 1452 -690
rect 1549 -691 1550 -641
rect 1682 -810 1683 -690
rect 1759 -691 1760 -641
rect 2095 -810 2096 -690
rect 37 -810 38 -692
rect 723 -693 724 -641
rect 730 -693 731 -641
rect 1493 -810 1494 -692
rect 1556 -693 1557 -641
rect 1969 -810 1970 -692
rect 1976 -693 1977 -641
rect 2088 -810 2089 -692
rect 261 -695 262 -641
rect 362 -810 363 -694
rect 401 -810 402 -694
rect 555 -695 556 -641
rect 562 -810 563 -694
rect 667 -695 668 -641
rect 681 -810 682 -694
rect 1710 -695 1711 -641
rect 1794 -695 1795 -641
rect 1927 -810 1928 -694
rect 1997 -695 1998 -641
rect 2116 -810 2117 -694
rect 156 -697 157 -641
rect 261 -810 262 -696
rect 282 -697 283 -641
rect 583 -697 584 -641
rect 590 -697 591 -641
rect 667 -810 668 -696
rect 702 -810 703 -696
rect 1304 -697 1305 -641
rect 1360 -810 1361 -696
rect 1773 -697 1774 -641
rect 1829 -697 1830 -641
rect 1962 -810 1963 -696
rect 2025 -697 2026 -641
rect 2165 -810 2166 -696
rect 128 -699 129 -641
rect 156 -810 157 -698
rect 240 -699 241 -641
rect 282 -810 283 -698
rect 310 -810 311 -698
rect 506 -699 507 -641
rect 523 -810 524 -698
rect 1486 -810 1487 -698
rect 1507 -699 1508 -641
rect 1794 -810 1795 -698
rect 1829 -810 1830 -698
rect 1941 -699 1942 -641
rect 2039 -699 2040 -641
rect 2217 -699 2218 -641
rect 114 -701 115 -641
rect 240 -810 241 -700
rect 324 -701 325 -641
rect 506 -810 507 -700
rect 548 -701 549 -641
rect 565 -701 566 -641
rect 569 -701 570 -641
rect 800 -810 801 -700
rect 814 -701 815 -641
rect 849 -810 850 -700
rect 852 -701 853 -641
rect 1745 -701 1746 -641
rect 1808 -701 1809 -641
rect 1941 -810 1942 -700
rect 2046 -701 2047 -641
rect 2172 -810 2173 -700
rect 86 -703 87 -641
rect 114 -810 115 -702
rect 324 -810 325 -702
rect 464 -703 465 -641
rect 492 -703 493 -641
rect 684 -810 685 -702
rect 737 -703 738 -641
rect 737 -810 738 -702
rect 737 -703 738 -641
rect 737 -810 738 -702
rect 744 -703 745 -641
rect 2207 -810 2208 -702
rect 5 -705 6 -641
rect 86 -810 87 -704
rect 415 -705 416 -641
rect 464 -810 465 -704
rect 492 -810 493 -704
rect 695 -705 696 -641
rect 747 -810 748 -704
rect 2102 -705 2103 -641
rect 408 -707 409 -641
rect 415 -810 416 -706
rect 429 -707 430 -641
rect 555 -810 556 -706
rect 590 -810 591 -706
rect 1465 -810 1466 -706
rect 1584 -707 1585 -641
rect 1703 -810 1704 -706
rect 1836 -707 1837 -641
rect 1976 -810 1977 -706
rect 2053 -707 2054 -641
rect 2200 -810 2201 -706
rect 303 -709 304 -641
rect 408 -810 409 -708
rect 422 -709 423 -641
rect 429 -810 430 -708
rect 432 -709 433 -641
rect 625 -709 626 -641
rect 639 -709 640 -641
rect 1780 -810 1781 -708
rect 1850 -709 1851 -641
rect 1997 -810 1998 -708
rect 2060 -709 2061 -641
rect 2193 -810 2194 -708
rect 100 -711 101 -641
rect 639 -810 640 -710
rect 646 -711 647 -641
rect 1227 -711 1228 -641
rect 1248 -711 1249 -641
rect 1759 -810 1760 -710
rect 1871 -711 1872 -641
rect 2025 -810 2026 -710
rect 100 -810 101 -712
rect 198 -713 199 -641
rect 219 -713 220 -641
rect 303 -810 304 -712
rect 422 -810 423 -712
rect 1202 -713 1203 -641
rect 1248 -810 1249 -712
rect 1458 -713 1459 -641
rect 1528 -713 1529 -641
rect 1871 -810 1872 -712
rect 1878 -713 1879 -641
rect 2046 -810 2047 -712
rect 163 -715 164 -641
rect 198 -810 199 -714
rect 443 -715 444 -641
rect 548 -810 549 -714
rect 604 -715 605 -641
rect 618 -810 619 -714
rect 653 -715 654 -641
rect 789 -715 790 -641
rect 814 -810 815 -714
rect 870 -715 871 -641
rect 947 -715 948 -641
rect 1129 -810 1130 -714
rect 1136 -810 1137 -714
rect 1745 -810 1746 -714
rect 1899 -715 1900 -641
rect 2039 -810 2040 -714
rect 163 -810 164 -716
rect 485 -717 486 -641
rect 534 -717 535 -641
rect 569 -810 570 -716
rect 576 -717 577 -641
rect 604 -810 605 -716
rect 611 -717 612 -641
rect 625 -810 626 -716
rect 660 -717 661 -641
rect 2228 -810 2229 -716
rect 23 -719 24 -641
rect 485 -810 486 -718
rect 583 -810 584 -718
rect 947 -810 948 -718
rect 996 -719 997 -641
rect 1087 -810 1088 -718
rect 1097 -719 1098 -641
rect 1528 -810 1529 -718
rect 1598 -719 1599 -641
rect 1710 -810 1711 -718
rect 1724 -719 1725 -641
rect 1836 -810 1837 -718
rect 1920 -719 1921 -641
rect 2060 -810 2061 -718
rect 23 -810 24 -720
rect 744 -810 745 -720
rect 772 -810 773 -720
rect 779 -721 780 -641
rect 793 -721 794 -641
rect 870 -810 871 -720
rect 989 -721 990 -641
rect 996 -810 997 -720
rect 1045 -721 1046 -641
rect 1556 -810 1557 -720
rect 1598 -810 1599 -720
rect 1675 -721 1676 -641
rect 1689 -721 1690 -641
rect 1808 -810 1809 -720
rect 1920 -810 1921 -720
rect 1948 -721 1949 -641
rect 289 -723 290 -641
rect 653 -810 654 -722
rect 663 -723 664 -641
rect 709 -723 710 -641
rect 758 -723 759 -641
rect 793 -810 794 -722
rect 856 -723 857 -641
rect 856 -810 857 -722
rect 856 -723 857 -641
rect 856 -810 857 -722
rect 1045 -810 1046 -722
rect 1066 -723 1067 -641
rect 1143 -810 1144 -722
rect 2102 -810 2103 -722
rect 184 -725 185 -641
rect 758 -810 759 -724
rect 779 -810 780 -724
rect 1115 -725 1116 -641
rect 1192 -725 1193 -641
rect 1227 -810 1228 -724
rect 1255 -725 1256 -641
rect 1304 -810 1305 -724
rect 1367 -725 1368 -641
rect 1430 -810 1431 -724
rect 1437 -725 1438 -641
rect 1549 -810 1550 -724
rect 1570 -725 1571 -641
rect 1689 -810 1690 -724
rect 1731 -725 1732 -641
rect 1850 -810 1851 -724
rect 1934 -725 1935 -641
rect 2053 -810 2054 -724
rect 184 -810 185 -726
rect 716 -727 717 -641
rect 898 -727 899 -641
rect 1066 -810 1067 -726
rect 1171 -727 1172 -641
rect 1437 -810 1438 -726
rect 1577 -727 1578 -641
rect 1675 -810 1676 -726
rect 1766 -727 1767 -641
rect 1899 -810 1900 -726
rect 177 -729 178 -641
rect 716 -810 717 -728
rect 898 -810 899 -728
rect 1146 -729 1147 -641
rect 1171 -810 1172 -728
rect 1409 -810 1410 -728
rect 1423 -729 1424 -641
rect 1570 -810 1571 -728
rect 1605 -810 1606 -728
rect 1640 -729 1641 -641
rect 1647 -729 1648 -641
rect 1773 -810 1774 -728
rect 1801 -729 1802 -641
rect 1934 -810 1935 -728
rect 58 -810 59 -730
rect 1146 -810 1147 -730
rect 1234 -731 1235 -641
rect 1255 -810 1256 -730
rect 1290 -731 1291 -641
rect 1584 -810 1585 -730
rect 1612 -731 1613 -641
rect 1724 -810 1725 -730
rect 1815 -731 1816 -641
rect 1948 -810 1949 -730
rect 177 -810 178 -732
rect 1269 -733 1270 -641
rect 1339 -733 1340 -641
rect 1423 -810 1424 -732
rect 1444 -733 1445 -641
rect 1801 -810 1802 -732
rect 219 -810 220 -734
rect 1612 -810 1613 -734
rect 1619 -735 1620 -641
rect 1752 -810 1753 -734
rect 250 -737 251 -641
rect 1192 -810 1193 -736
rect 1206 -737 1207 -641
rect 1269 -810 1270 -736
rect 1353 -737 1354 -641
rect 1444 -810 1445 -736
rect 1472 -737 1473 -641
rect 1619 -810 1620 -736
rect 1633 -737 1634 -641
rect 1731 -810 1732 -736
rect 142 -810 143 -738
rect 1472 -810 1473 -738
rect 1500 -739 1501 -641
rect 1640 -810 1641 -738
rect 1654 -739 1655 -641
rect 1878 -810 1879 -738
rect 205 -810 206 -740
rect 1500 -810 1501 -740
rect 1514 -741 1515 -641
rect 1654 -810 1655 -740
rect 1668 -741 1669 -641
rect 2018 -810 2019 -740
rect 289 -810 290 -742
rect 499 -743 500 -641
rect 537 -743 538 -641
rect 989 -810 990 -742
rect 1024 -743 1025 -641
rect 1577 -810 1578 -742
rect 1696 -743 1697 -641
rect 1815 -810 1816 -742
rect 373 -745 374 -641
rect 1696 -810 1697 -744
rect 352 -747 353 -641
rect 373 -810 374 -746
rect 380 -747 381 -641
rect 576 -810 577 -746
rect 611 -810 612 -746
rect 688 -747 689 -641
rect 726 -810 727 -746
rect 1353 -810 1354 -746
rect 1370 -810 1371 -746
rect 1843 -810 1844 -746
rect 254 -749 255 -641
rect 380 -810 381 -748
rect 394 -749 395 -641
rect 534 -810 535 -748
rect 632 -749 633 -641
rect 660 -810 661 -748
rect 674 -749 675 -641
rect 709 -810 710 -748
rect 1017 -749 1018 -641
rect 1024 -810 1025 -748
rect 1038 -749 1039 -641
rect 1115 -810 1116 -748
rect 1185 -749 1186 -641
rect 1234 -810 1235 -748
rect 1241 -749 1242 -641
rect 1290 -810 1291 -748
rect 1374 -749 1375 -641
rect 1458 -810 1459 -748
rect 1514 -810 1515 -748
rect 1521 -749 1522 -641
rect 1535 -749 1536 -641
rect 1633 -810 1634 -748
rect 254 -810 255 -750
rect 520 -751 521 -641
rect 597 -751 598 -641
rect 674 -810 675 -750
rect 688 -810 689 -750
rect 1164 -751 1165 -641
rect 1185 -810 1186 -750
rect 1563 -751 1564 -641
rect 331 -753 332 -641
rect 352 -810 353 -752
rect 387 -753 388 -641
rect 597 -810 598 -752
rect 968 -753 969 -641
rect 1017 -810 1018 -752
rect 1094 -810 1095 -752
rect 1339 -810 1340 -752
rect 1346 -753 1347 -641
rect 1521 -810 1522 -752
rect 1535 -810 1536 -752
rect 1864 -810 1865 -752
rect 275 -755 276 -641
rect 331 -810 332 -754
rect 387 -810 388 -754
rect 478 -755 479 -641
rect 499 -810 500 -754
rect 513 -755 514 -641
rect 933 -755 934 -641
rect 968 -810 969 -754
rect 975 -755 976 -641
rect 1038 -810 1039 -754
rect 1139 -810 1140 -754
rect 1374 -810 1375 -754
rect 1381 -755 1382 -641
rect 1647 -810 1648 -754
rect 275 -810 276 -756
rect 296 -757 297 -641
rect 359 -757 360 -641
rect 478 -810 479 -756
rect 513 -810 514 -756
rect 919 -757 920 -641
rect 954 -757 955 -641
rect 975 -810 976 -756
rect 1153 -757 1154 -641
rect 1241 -810 1242 -756
rect 1283 -757 1284 -641
rect 1346 -810 1347 -756
rect 1395 -757 1396 -641
rect 1507 -810 1508 -756
rect 1538 -810 1539 -756
rect 1766 -810 1767 -756
rect 208 -759 209 -641
rect 919 -810 920 -758
rect 1157 -759 1158 -641
rect 1164 -810 1165 -758
rect 1206 -810 1207 -758
rect 1220 -759 1221 -641
rect 1311 -759 1312 -641
rect 1381 -810 1382 -758
rect 1395 -810 1396 -758
rect 1402 -759 1403 -641
rect 1542 -759 1543 -641
rect 1668 -810 1669 -758
rect 44 -810 45 -760
rect 1542 -810 1543 -760
rect 135 -810 136 -762
rect 208 -810 209 -762
rect 296 -810 297 -762
rect 541 -763 542 -641
rect 786 -810 787 -762
rect 954 -810 955 -762
rect 961 -763 962 -641
rect 1311 -810 1312 -762
rect 1318 -763 1319 -641
rect 1563 -810 1564 -762
rect 345 -765 346 -641
rect 359 -810 360 -764
rect 443 -810 444 -764
rect 527 -765 528 -641
rect 810 -765 811 -641
rect 1283 -810 1284 -764
rect 79 -767 80 -641
rect 527 -810 528 -766
rect 884 -767 885 -641
rect 933 -810 934 -766
rect 1157 -810 1158 -766
rect 2032 -767 2033 -641
rect 79 -810 80 -768
rect 632 -810 633 -768
rect 905 -769 906 -641
rect 961 -810 962 -768
rect 1209 -810 1210 -768
rect 2032 -810 2033 -768
rect 107 -771 108 -641
rect 884 -810 885 -770
rect 1220 -810 1221 -770
rect 2214 -810 2215 -770
rect 107 -810 108 -772
rect 821 -773 822 -641
rect 1262 -773 1263 -641
rect 1402 -810 1403 -772
rect 268 -775 269 -641
rect 905 -810 906 -774
rect 268 -810 269 -776
rect 338 -777 339 -641
rect 345 -810 346 -776
rect 649 -777 650 -641
rect 821 -810 822 -776
rect 835 -777 836 -641
rect 880 -810 881 -776
rect 1262 -810 1263 -776
rect 338 -810 339 -778
rect 751 -779 752 -641
rect 828 -779 829 -641
rect 835 -810 836 -778
rect 450 -781 451 -641
rect 730 -810 731 -780
rect 751 -810 752 -780
rect 1416 -781 1417 -641
rect 128 -810 129 -782
rect 1416 -810 1417 -782
rect 233 -785 234 -641
rect 450 -810 451 -784
rect 457 -785 458 -641
rect 541 -810 542 -784
rect 828 -810 829 -784
rect 1913 -785 1914 -641
rect 233 -810 234 -786
rect 394 -810 395 -786
rect 457 -810 458 -786
rect 842 -787 843 -641
rect 1787 -787 1788 -641
rect 1913 -810 1914 -786
rect 471 -789 472 -641
rect 646 -810 647 -788
rect 842 -810 843 -788
rect 912 -789 913 -641
rect 1661 -789 1662 -641
rect 1787 -810 1788 -788
rect 471 -810 472 -790
rect 1010 -810 1011 -790
rect 1276 -791 1277 -641
rect 1661 -810 1662 -790
rect 520 -810 521 -792
rect 1318 -810 1319 -792
rect 912 -810 913 -794
rect 1297 -795 1298 -641
rect 1276 -810 1277 -796
rect 1479 -797 1480 -641
rect 1297 -810 1298 -798
rect 1332 -799 1333 -641
rect 1388 -799 1389 -641
rect 1479 -810 1480 -798
rect 1325 -801 1326 -641
rect 1388 -810 1389 -800
rect 226 -803 227 -641
rect 1325 -810 1326 -802
rect 1332 -810 1333 -802
rect 1906 -810 1907 -802
rect 226 -810 227 -804
rect 586 -805 587 -641
rect 436 -807 437 -641
rect 586 -810 587 -806
rect 222 -810 223 -808
rect 436 -810 437 -808
rect 9 -820 10 -818
rect 1626 -820 1627 -818
rect 1661 -820 1662 -818
rect 2361 -999 2362 -819
rect 2403 -820 2404 -818
rect 2417 -999 2418 -819
rect 9 -999 10 -821
rect 93 -822 94 -818
rect 103 -999 104 -821
rect 352 -822 353 -818
rect 457 -822 458 -818
rect 590 -822 591 -818
rect 614 -999 615 -821
rect 653 -822 654 -818
rect 674 -822 675 -818
rect 747 -822 748 -818
rect 782 -999 783 -821
rect 849 -822 850 -818
rect 898 -822 899 -818
rect 898 -999 899 -821
rect 898 -822 899 -818
rect 898 -999 899 -821
rect 947 -822 948 -818
rect 1314 -999 1315 -821
rect 1332 -999 1333 -821
rect 1423 -822 1424 -818
rect 1538 -822 1539 -818
rect 2095 -822 2096 -818
rect 2326 -822 2327 -818
rect 2336 -999 2337 -821
rect 2343 -999 2344 -821
rect 2403 -999 2404 -821
rect 16 -824 17 -818
rect 191 -824 192 -818
rect 212 -824 213 -818
rect 212 -999 213 -823
rect 212 -824 213 -818
rect 212 -999 213 -823
rect 222 -824 223 -818
rect 2249 -824 2250 -818
rect 2277 -824 2278 -818
rect 2326 -999 2327 -823
rect 2347 -824 2348 -818
rect 2375 -999 2376 -823
rect 16 -999 17 -825
rect 1325 -826 1326 -818
rect 1335 -826 1336 -818
rect 1521 -826 1522 -818
rect 1598 -826 1599 -818
rect 1601 -832 1602 -825
rect 1626 -999 1627 -825
rect 1654 -826 1655 -818
rect 1661 -999 1662 -825
rect 1815 -826 1816 -818
rect 1934 -826 1935 -818
rect 1934 -999 1935 -825
rect 1934 -826 1935 -818
rect 1934 -999 1935 -825
rect 2095 -999 2096 -825
rect 2151 -826 2152 -818
rect 2277 -999 2278 -825
rect 2340 -999 2341 -825
rect 2347 -999 2348 -825
rect 2368 -999 2369 -825
rect 44 -828 45 -818
rect 1696 -828 1697 -818
rect 1815 -999 1816 -827
rect 1878 -828 1879 -818
rect 2151 -999 2152 -827
rect 2179 -828 2180 -818
rect 44 -999 45 -829
rect 940 -830 941 -818
rect 947 -999 948 -829
rect 968 -830 969 -818
rect 989 -830 990 -818
rect 1423 -999 1424 -829
rect 1598 -999 1599 -829
rect 1717 -830 1718 -818
rect 1878 -999 1879 -829
rect 1941 -830 1942 -818
rect 1990 -830 1991 -818
rect 2179 -999 2180 -829
rect 58 -832 59 -818
rect 754 -832 755 -818
rect 817 -999 818 -831
rect 1409 -832 1410 -818
rect 1717 -999 1718 -831
rect 1899 -832 1900 -818
rect 1990 -999 1991 -831
rect 58 -999 59 -833
rect 135 -834 136 -818
rect 142 -999 143 -833
rect 222 -999 223 -833
rect 254 -834 255 -818
rect 590 -999 591 -833
rect 635 -999 636 -833
rect 926 -834 927 -818
rect 989 -999 990 -833
rect 1132 -834 1133 -818
rect 1136 -834 1137 -818
rect 1801 -834 1802 -818
rect 1941 -999 1942 -833
rect 1983 -834 1984 -818
rect 79 -836 80 -818
rect 261 -836 262 -818
rect 282 -836 283 -818
rect 362 -836 363 -818
rect 422 -836 423 -818
rect 849 -999 850 -835
rect 870 -836 871 -818
rect 940 -999 941 -835
rect 996 -836 997 -818
rect 1244 -999 1245 -835
rect 1248 -836 1249 -818
rect 1521 -999 1522 -835
rect 1605 -836 1606 -818
rect 1696 -999 1697 -835
rect 1983 -999 1984 -835
rect 2025 -836 2026 -818
rect 72 -838 73 -818
rect 996 -999 997 -837
rect 1020 -999 1021 -837
rect 1556 -838 1557 -818
rect 1573 -999 1574 -837
rect 2025 -999 2026 -837
rect 72 -999 73 -839
rect 667 -840 668 -818
rect 681 -999 682 -839
rect 716 -840 717 -818
rect 821 -840 822 -818
rect 870 -999 871 -839
rect 926 -999 927 -839
rect 1192 -840 1193 -818
rect 1195 -999 1196 -839
rect 2109 -840 2110 -818
rect 79 -999 80 -841
rect 324 -842 325 -818
rect 352 -999 353 -841
rect 499 -842 500 -818
rect 506 -842 507 -818
rect 723 -842 724 -818
rect 772 -842 773 -818
rect 821 -999 822 -841
rect 1010 -842 1011 -818
rect 2109 -999 2110 -841
rect 121 -844 122 -818
rect 268 -844 269 -818
rect 282 -999 283 -843
rect 1160 -844 1161 -818
rect 1174 -844 1175 -818
rect 1773 -844 1774 -818
rect 47 -846 48 -818
rect 1773 -999 1774 -845
rect 128 -848 129 -818
rect 562 -848 563 -818
rect 646 -848 647 -818
rect 831 -848 832 -818
rect 1010 -999 1011 -847
rect 1087 -848 1088 -818
rect 1094 -848 1095 -818
rect 1122 -848 1123 -818
rect 1129 -848 1130 -818
rect 2235 -848 2236 -818
rect 128 -999 129 -849
rect 1041 -999 1042 -849
rect 1045 -850 1046 -818
rect 1087 -999 1088 -849
rect 1094 -999 1095 -849
rect 1101 -850 1102 -818
rect 1111 -850 1112 -818
rect 2046 -850 2047 -818
rect 2235 -999 2236 -849
rect 2284 -850 2285 -818
rect 145 -852 146 -818
rect 800 -852 801 -818
rect 828 -852 829 -818
rect 1129 -999 1130 -851
rect 1136 -999 1137 -851
rect 1227 -852 1228 -818
rect 1248 -999 1249 -851
rect 1388 -852 1389 -818
rect 1402 -852 1403 -818
rect 1409 -999 1410 -851
rect 1430 -852 1431 -818
rect 2046 -999 2047 -851
rect 170 -854 171 -818
rect 191 -999 192 -853
rect 205 -854 206 -818
rect 1801 -999 1802 -853
rect 170 -999 171 -855
rect 271 -999 272 -855
rect 296 -856 297 -818
rect 583 -856 584 -818
rect 646 -999 647 -855
rect 1255 -856 1256 -818
rect 1272 -999 1273 -855
rect 1969 -856 1970 -818
rect 184 -858 185 -818
rect 289 -858 290 -818
rect 310 -858 311 -818
rect 376 -999 377 -857
rect 422 -999 423 -857
rect 1108 -858 1109 -818
rect 1139 -858 1140 -818
rect 1241 -858 1242 -818
rect 1255 -999 1256 -857
rect 1353 -858 1354 -818
rect 1360 -858 1361 -818
rect 2319 -858 2320 -818
rect 184 -999 185 -859
rect 758 -860 759 -818
rect 775 -999 776 -859
rect 1108 -999 1109 -859
rect 1143 -860 1144 -818
rect 2074 -860 2075 -818
rect 198 -862 199 -818
rect 289 -999 290 -861
rect 310 -999 311 -861
rect 450 -862 451 -818
rect 457 -999 458 -861
rect 548 -862 549 -818
rect 562 -999 563 -861
rect 569 -862 570 -818
rect 653 -999 654 -861
rect 1024 -862 1025 -818
rect 1045 -999 1046 -861
rect 1059 -862 1060 -818
rect 1101 -999 1102 -861
rect 1185 -862 1186 -818
rect 1206 -862 1207 -818
rect 1759 -862 1760 -818
rect 1969 -999 1970 -861
rect 2004 -862 2005 -818
rect 2074 -999 2075 -861
rect 2130 -862 2131 -818
rect 156 -864 157 -818
rect 198 -999 199 -863
rect 205 -999 206 -863
rect 233 -864 234 -818
rect 254 -999 255 -863
rect 520 -864 521 -818
rect 527 -864 528 -818
rect 1206 -999 1207 -863
rect 1209 -864 1210 -818
rect 2123 -864 2124 -818
rect 2130 -999 2131 -863
rect 2165 -864 2166 -818
rect 156 -999 157 -865
rect 443 -866 444 -818
rect 478 -866 479 -818
rect 520 -999 521 -865
rect 527 -999 528 -865
rect 807 -866 808 -818
rect 828 -999 829 -865
rect 1780 -866 1781 -818
rect 2004 -999 2005 -865
rect 2053 -866 2054 -818
rect 2123 -999 2124 -865
rect 2137 -866 2138 -818
rect 163 -868 164 -818
rect 450 -999 451 -867
rect 478 -999 479 -867
rect 772 -999 773 -867
rect 807 -999 808 -867
rect 1080 -868 1081 -818
rect 1143 -999 1144 -867
rect 1216 -868 1217 -818
rect 1220 -868 1221 -818
rect 2060 -868 2061 -818
rect 2102 -868 2103 -818
rect 2137 -999 2138 -867
rect 163 -999 164 -869
rect 331 -870 332 -818
rect 359 -870 360 -818
rect 569 -999 570 -869
rect 667 -999 668 -869
rect 2350 -999 2351 -869
rect 187 -872 188 -818
rect 1780 -999 1781 -871
rect 1787 -872 1788 -818
rect 2060 -999 2061 -871
rect 2102 -999 2103 -871
rect 2158 -872 2159 -818
rect 219 -999 220 -873
rect 800 -999 801 -873
rect 957 -874 958 -818
rect 1402 -999 1403 -873
rect 1556 -999 1557 -873
rect 1647 -874 1648 -818
rect 1654 -999 1655 -873
rect 1745 -874 1746 -818
rect 1787 -999 1788 -873
rect 1829 -874 1830 -818
rect 2053 -999 2054 -873
rect 2088 -874 2089 -818
rect 233 -999 234 -875
rect 303 -876 304 -818
rect 317 -876 318 -818
rect 317 -999 318 -875
rect 317 -876 318 -818
rect 317 -999 318 -875
rect 324 -999 325 -875
rect 373 -876 374 -818
rect 387 -876 388 -818
rect 443 -999 444 -875
rect 492 -876 493 -818
rect 968 -999 969 -875
rect 1024 -999 1025 -875
rect 1528 -876 1529 -818
rect 1605 -999 1606 -875
rect 1675 -876 1676 -818
rect 1682 -876 1683 -818
rect 1759 -999 1760 -875
rect 1829 -999 1830 -875
rect 1913 -876 1914 -818
rect 100 -878 101 -818
rect 387 -999 388 -877
rect 408 -878 409 -818
rect 548 -999 549 -877
rect 688 -878 689 -818
rect 726 -878 727 -818
rect 737 -878 738 -818
rect 758 -999 759 -877
rect 1055 -999 1056 -877
rect 2081 -878 2082 -818
rect 100 -999 101 -879
rect 936 -999 937 -879
rect 1080 -999 1081 -879
rect 1164 -880 1165 -818
rect 1185 -999 1186 -879
rect 1766 -880 1767 -818
rect 1871 -880 1872 -818
rect 2088 -999 2089 -879
rect 121 -999 122 -881
rect 373 -999 374 -881
rect 408 -999 409 -881
rect 415 -882 416 -818
rect 436 -882 437 -818
rect 506 -999 507 -881
rect 513 -882 514 -818
rect 719 -999 720 -881
rect 723 -999 724 -881
rect 1031 -882 1032 -818
rect 1146 -882 1147 -818
rect 1517 -999 1518 -881
rect 1647 -999 1648 -881
rect 1738 -882 1739 -818
rect 1745 -999 1746 -881
rect 1843 -882 1844 -818
rect 1913 -999 1914 -881
rect 1962 -882 1963 -818
rect 2081 -999 2082 -881
rect 2144 -882 2145 -818
rect 2 -884 3 -818
rect 415 -999 416 -883
rect 492 -999 493 -883
rect 765 -884 766 -818
rect 1031 -999 1032 -883
rect 1066 -884 1067 -818
rect 1157 -884 1158 -818
rect 2298 -884 2299 -818
rect 2 -999 3 -885
rect 177 -886 178 -818
rect 247 -886 248 -818
rect 303 -999 304 -885
rect 359 -999 360 -885
rect 380 -886 381 -818
rect 499 -999 500 -885
rect 530 -999 531 -885
rect 534 -886 535 -818
rect 583 -999 584 -885
rect 688 -999 689 -885
rect 709 -886 710 -818
rect 737 -999 738 -885
rect 884 -886 885 -818
rect 954 -886 955 -818
rect 2298 -999 2299 -885
rect 65 -888 66 -818
rect 1962 -999 1963 -887
rect 2144 -999 2145 -887
rect 2172 -888 2173 -818
rect 65 -999 66 -889
rect 394 -890 395 -818
rect 464 -890 465 -818
rect 534 -999 535 -889
rect 541 -890 542 -818
rect 674 -999 675 -889
rect 698 -890 699 -818
rect 919 -890 920 -818
rect 1052 -890 1053 -818
rect 1066 -999 1067 -889
rect 1157 -999 1158 -889
rect 1199 -890 1200 -818
rect 1213 -890 1214 -818
rect 2242 -890 2243 -818
rect 86 -892 87 -818
rect 394 -999 395 -891
rect 401 -892 402 -818
rect 464 -999 465 -891
rect 513 -999 514 -891
rect 597 -892 598 -818
rect 702 -892 703 -818
rect 1171 -892 1172 -818
rect 1199 -999 1200 -891
rect 1276 -892 1277 -818
rect 1286 -999 1287 -891
rect 1528 -999 1529 -891
rect 1682 -999 1683 -891
rect 1703 -892 1704 -818
rect 1738 -999 1739 -891
rect 1864 -892 1865 -818
rect 2172 -999 2173 -891
rect 2193 -892 2194 -818
rect 2207 -892 2208 -818
rect 2242 -999 2243 -891
rect 86 -999 87 -893
rect 366 -894 367 -818
rect 380 -999 381 -893
rect 611 -894 612 -818
rect 702 -999 703 -893
rect 835 -894 836 -818
rect 905 -894 906 -818
rect 1052 -999 1053 -893
rect 1125 -999 1126 -893
rect 1864 -999 1865 -893
rect 2193 -999 2194 -893
rect 2228 -894 2229 -818
rect 107 -896 108 -818
rect 905 -999 906 -895
rect 919 -999 920 -895
rect 1115 -896 1116 -818
rect 1164 -999 1165 -895
rect 1269 -896 1270 -818
rect 1290 -896 1291 -818
rect 1388 -999 1389 -895
rect 1395 -896 1396 -818
rect 1430 -999 1431 -895
rect 1766 -999 1767 -895
rect 2312 -896 2313 -818
rect 107 -999 108 -897
rect 240 -898 241 -818
rect 247 -999 248 -897
rect 1017 -898 1018 -818
rect 1038 -898 1039 -818
rect 1115 -999 1116 -897
rect 1171 -999 1172 -897
rect 2200 -898 2201 -818
rect 2207 -999 2208 -897
rect 2263 -898 2264 -818
rect 51 -900 52 -818
rect 240 -999 241 -899
rect 261 -999 262 -899
rect 632 -900 633 -818
rect 765 -999 766 -899
rect 814 -900 815 -818
rect 1192 -999 1193 -899
rect 1276 -999 1277 -899
rect 1290 -999 1291 -899
rect 1346 -900 1347 -818
rect 1353 -999 1354 -899
rect 1584 -900 1585 -818
rect 1794 -900 1795 -818
rect 1871 -999 1872 -899
rect 1892 -900 1893 -818
rect 2263 -999 2264 -899
rect 51 -999 52 -901
rect 628 -999 629 -901
rect 639 -902 640 -818
rect 1892 -999 1893 -901
rect 2018 -902 2019 -818
rect 2312 -999 2313 -901
rect 124 -904 125 -818
rect 1675 -999 1676 -903
rect 1794 -999 1795 -903
rect 1906 -904 1907 -818
rect 2018 -999 2019 -903
rect 2067 -904 2068 -818
rect 2186 -904 2187 -818
rect 2228 -999 2229 -903
rect 149 -906 150 -818
rect 436 -999 437 -905
rect 541 -999 542 -905
rect 611 -999 612 -905
rect 618 -906 619 -818
rect 632 -999 633 -905
rect 786 -906 787 -818
rect 835 -999 836 -905
rect 1213 -999 1214 -905
rect 1269 -999 1270 -905
rect 1304 -906 1305 -818
rect 2354 -999 2355 -905
rect 30 -908 31 -818
rect 786 -999 787 -907
rect 796 -999 797 -907
rect 884 -999 885 -907
rect 1220 -999 1221 -907
rect 1234 -908 1235 -818
rect 1241 -999 1242 -907
rect 1808 -908 1809 -818
rect 1843 -999 1844 -907
rect 2039 -908 2040 -818
rect 2067 -999 2068 -907
rect 2116 -908 2117 -818
rect 2200 -999 2201 -907
rect 2256 -908 2257 -818
rect 30 -999 31 -909
rect 177 -999 178 -909
rect 180 -999 181 -909
rect 709 -999 710 -909
rect 716 -999 717 -909
rect 1808 -999 1809 -909
rect 1906 -999 1907 -909
rect 1955 -910 1956 -818
rect 2039 -999 2040 -909
rect 2291 -910 2292 -818
rect 135 -999 136 -911
rect 2116 -999 2117 -911
rect 2214 -912 2215 -818
rect 2256 -999 2257 -911
rect 149 -999 150 -913
rect 1174 -999 1175 -913
rect 1223 -914 1224 -818
rect 1703 -999 1704 -913
rect 1955 -999 1956 -913
rect 1997 -914 1998 -818
rect 2214 -999 2215 -913
rect 2270 -914 2271 -818
rect 226 -916 227 -818
rect 639 -999 640 -915
rect 814 -999 815 -915
rect 1311 -916 1312 -818
rect 1325 -999 1326 -915
rect 1416 -916 1417 -818
rect 1535 -916 1536 -818
rect 2186 -999 2187 -915
rect 2270 -999 2271 -915
rect 2305 -916 2306 -818
rect 226 -999 227 -917
rect 877 -918 878 -818
rect 1178 -918 1179 -818
rect 1416 -999 1417 -917
rect 1493 -918 1494 -818
rect 2305 -999 2306 -917
rect 23 -920 24 -818
rect 877 -999 878 -919
rect 1122 -999 1123 -919
rect 1178 -999 1179 -919
rect 1227 -999 1228 -919
rect 1262 -920 1263 -818
rect 1304 -999 1305 -919
rect 1444 -920 1445 -818
rect 1493 -999 1494 -919
rect 1549 -920 1550 -818
rect 1584 -999 1585 -919
rect 1633 -920 1634 -818
rect 1997 -999 1998 -919
rect 2032 -920 2033 -818
rect 23 -999 24 -921
rect 114 -922 115 -818
rect 268 -999 269 -921
rect 2291 -999 2292 -921
rect 114 -999 115 -923
rect 485 -924 486 -818
rect 593 -924 594 -818
rect 954 -999 955 -923
rect 1234 -999 1235 -923
rect 1437 -924 1438 -818
rect 1535 -999 1536 -923
rect 1612 -924 1613 -818
rect 1633 -999 1634 -923
rect 1710 -924 1711 -818
rect 1857 -924 1858 -818
rect 2032 -999 2033 -923
rect 275 -926 276 -818
rect 296 -999 297 -925
rect 345 -926 346 -818
rect 618 -999 619 -925
rect 1262 -999 1263 -925
rect 1297 -926 1298 -818
rect 1311 -999 1312 -925
rect 2284 -999 2285 -925
rect 275 -999 276 -927
rect 429 -928 430 -818
rect 485 -999 486 -927
rect 555 -928 556 -818
rect 597 -999 598 -927
rect 604 -928 605 -818
rect 684 -928 685 -818
rect 1297 -999 1298 -927
rect 1339 -928 1340 -818
rect 1444 -999 1445 -927
rect 1549 -999 1550 -927
rect 1563 -928 1564 -818
rect 1612 -999 1613 -927
rect 1619 -928 1620 -818
rect 1710 -999 1711 -927
rect 1822 -928 1823 -818
rect 1857 -999 1858 -927
rect 1885 -928 1886 -818
rect 345 -999 346 -929
rect 660 -930 661 -818
rect 1283 -930 1284 -818
rect 1437 -999 1438 -929
rect 1563 -999 1564 -929
rect 1668 -930 1669 -818
rect 1822 -999 1823 -929
rect 1836 -930 1837 -818
rect 1885 -999 1886 -929
rect 1948 -930 1949 -818
rect 19 -932 20 -818
rect 1836 -999 1837 -931
rect 331 -999 332 -933
rect 1283 -999 1284 -933
rect 1339 -999 1340 -933
rect 1451 -934 1452 -818
rect 1500 -934 1501 -818
rect 1668 -999 1669 -933
rect 366 -999 367 -935
rect 1398 -999 1399 -935
rect 1500 -999 1501 -935
rect 1577 -936 1578 -818
rect 1619 -999 1620 -935
rect 1724 -936 1725 -818
rect 401 -999 402 -937
rect 695 -938 696 -818
rect 1059 -999 1060 -937
rect 1948 -999 1949 -937
rect 187 -999 188 -939
rect 695 -999 696 -939
rect 1318 -940 1319 -818
rect 1451 -999 1452 -939
rect 1577 -999 1578 -939
rect 1899 -999 1900 -939
rect 429 -999 430 -941
rect 1013 -942 1014 -818
rect 1318 -999 1319 -941
rect 1507 -942 1508 -818
rect 1724 -999 1725 -941
rect 1850 -942 1851 -818
rect 604 -999 605 -943
rect 842 -944 843 -818
rect 1346 -999 1347 -943
rect 1395 -999 1396 -943
rect 1507 -999 1508 -943
rect 1591 -944 1592 -818
rect 1850 -999 1851 -943
rect 1927 -944 1928 -818
rect 660 -999 661 -945
rect 912 -946 913 -818
rect 1360 -999 1361 -945
rect 1381 -946 1382 -818
rect 1591 -999 1592 -945
rect 1689 -946 1690 -818
rect 1927 -999 1928 -945
rect 1976 -946 1977 -818
rect 744 -948 745 -818
rect 1689 -999 1690 -947
rect 1976 -999 1977 -947
rect 2011 -948 2012 -818
rect 744 -999 745 -949
rect 793 -950 794 -818
rect 842 -999 843 -949
rect 933 -950 934 -818
rect 1363 -950 1364 -818
rect 2158 -999 2159 -949
rect 555 -999 556 -951
rect 933 -999 934 -951
rect 1367 -952 1368 -818
rect 1752 -952 1753 -818
rect 1920 -952 1921 -818
rect 2011 -999 2012 -951
rect 793 -999 794 -953
rect 961 -954 962 -818
rect 1017 -999 1018 -953
rect 1752 -999 1753 -953
rect 856 -956 857 -818
rect 912 -999 913 -955
rect 961 -999 962 -955
rect 982 -956 983 -818
rect 1367 -999 1368 -955
rect 1458 -956 1459 -818
rect 856 -999 857 -957
rect 891 -958 892 -818
rect 982 -999 983 -957
rect 1003 -958 1004 -818
rect 1370 -958 1371 -818
rect 2165 -999 2166 -957
rect 471 -960 472 -818
rect 891 -999 892 -959
rect 1374 -960 1375 -818
rect 1920 -999 1921 -959
rect 471 -999 472 -961
rect 576 -962 577 -818
rect 586 -962 587 -818
rect 1003 -999 1004 -961
rect 1374 -999 1375 -961
rect 1479 -962 1480 -818
rect 576 -999 577 -963
rect 625 -964 626 -818
rect 1381 -999 1382 -963
rect 1486 -964 1487 -818
rect 625 -999 626 -965
rect 2319 -999 2320 -965
rect 1458 -999 1459 -967
rect 1542 -968 1543 -818
rect 1479 -999 1480 -969
rect 1570 -970 1571 -818
rect 1486 -999 1487 -971
rect 1731 -972 1732 -818
rect 1465 -974 1466 -818
rect 1731 -999 1732 -973
rect 1465 -999 1466 -975
rect 1472 -976 1473 -818
rect 1542 -999 1543 -975
rect 1640 -976 1641 -818
rect 1073 -978 1074 -818
rect 1472 -999 1473 -977
rect 1514 -978 1515 -818
rect 1640 -999 1641 -977
rect 779 -980 780 -818
rect 1073 -999 1074 -979
rect 1514 -999 1515 -979
rect 2249 -999 2250 -979
rect 1570 -999 1571 -981
rect 2221 -982 2222 -818
rect 751 -984 752 -818
rect 2221 -999 2222 -983
rect 37 -986 38 -818
rect 751 -999 752 -985
rect 37 -999 38 -987
rect 975 -988 976 -818
rect 975 -999 976 -989
rect 1150 -990 1151 -818
rect 730 -992 731 -818
rect 1150 -999 1151 -991
rect 730 -999 731 -993
rect 863 -994 864 -818
rect 338 -996 339 -818
rect 863 -999 864 -995
rect 338 -999 339 -997
rect 390 -999 391 -997
rect 9 -1009 10 -1007
rect 761 -1166 762 -1008
rect 772 -1009 773 -1007
rect 2137 -1009 2138 -1007
rect 2284 -1009 2285 -1007
rect 2340 -1166 2341 -1008
rect 2375 -1009 2376 -1007
rect 2431 -1166 2432 -1008
rect 9 -1166 10 -1010
rect 58 -1011 59 -1007
rect 93 -1011 94 -1007
rect 2256 -1011 2257 -1007
rect 2298 -1011 2299 -1007
rect 2375 -1166 2376 -1010
rect 2382 -1166 2383 -1010
rect 2392 -1166 2393 -1010
rect 2403 -1011 2404 -1007
rect 2438 -1166 2439 -1010
rect 16 -1013 17 -1007
rect 58 -1166 59 -1012
rect 93 -1166 94 -1012
rect 842 -1013 843 -1007
rect 884 -1013 885 -1007
rect 933 -1166 934 -1012
rect 936 -1013 937 -1007
rect 1388 -1013 1389 -1007
rect 1409 -1013 1410 -1007
rect 1409 -1166 1410 -1012
rect 1409 -1013 1410 -1007
rect 1409 -1166 1410 -1012
rect 1507 -1013 1508 -1007
rect 1577 -1166 1578 -1012
rect 1703 -1013 1704 -1007
rect 2298 -1166 2299 -1012
rect 2368 -1013 2369 -1007
rect 2403 -1166 2404 -1012
rect 2417 -1013 2418 -1007
rect 2424 -1166 2425 -1012
rect 16 -1166 17 -1014
rect 331 -1015 332 -1007
rect 345 -1015 346 -1007
rect 1006 -1166 1007 -1014
rect 1020 -1015 1021 -1007
rect 2228 -1015 2229 -1007
rect 103 -1017 104 -1007
rect 1150 -1017 1151 -1007
rect 1174 -1017 1175 -1007
rect 1871 -1017 1872 -1007
rect 2123 -1017 2124 -1007
rect 2368 -1166 2369 -1016
rect 110 -1166 111 -1018
rect 317 -1019 318 -1007
rect 324 -1019 325 -1007
rect 331 -1166 332 -1018
rect 345 -1166 346 -1018
rect 443 -1019 444 -1007
rect 590 -1019 591 -1007
rect 628 -1019 629 -1007
rect 646 -1019 647 -1007
rect 954 -1019 955 -1007
rect 964 -1166 965 -1018
rect 2242 -1019 2243 -1007
rect 117 -1166 118 -1020
rect 1451 -1021 1452 -1007
rect 1514 -1021 1515 -1007
rect 1682 -1021 1683 -1007
rect 1689 -1021 1690 -1007
rect 1703 -1166 1704 -1020
rect 1787 -1021 1788 -1007
rect 2123 -1166 2124 -1020
rect 2165 -1021 2166 -1007
rect 2228 -1166 2229 -1020
rect 128 -1023 129 -1007
rect 782 -1023 783 -1007
rect 793 -1023 794 -1007
rect 1108 -1023 1109 -1007
rect 1122 -1023 1123 -1007
rect 1360 -1023 1361 -1007
rect 1514 -1166 1515 -1022
rect 1535 -1023 1536 -1007
rect 1570 -1023 1571 -1007
rect 1570 -1166 1571 -1022
rect 1570 -1023 1571 -1007
rect 1570 -1166 1571 -1022
rect 1710 -1023 1711 -1007
rect 1787 -1166 1788 -1022
rect 1801 -1023 1802 -1007
rect 2389 -1166 2390 -1022
rect 128 -1166 129 -1024
rect 261 -1025 262 -1007
rect 268 -1166 269 -1024
rect 478 -1025 479 -1007
rect 590 -1166 591 -1024
rect 667 -1025 668 -1007
rect 733 -1166 734 -1024
rect 2291 -1025 2292 -1007
rect 86 -1027 87 -1007
rect 667 -1166 668 -1026
rect 779 -1027 780 -1007
rect 1990 -1027 1991 -1007
rect 2102 -1027 2103 -1007
rect 2291 -1166 2292 -1026
rect 86 -1166 87 -1028
rect 135 -1029 136 -1007
rect 138 -1029 139 -1007
rect 1892 -1029 1893 -1007
rect 1962 -1029 1963 -1007
rect 1990 -1166 1991 -1028
rect 2172 -1029 2173 -1007
rect 2242 -1166 2243 -1028
rect 135 -1166 136 -1030
rect 1822 -1031 1823 -1007
rect 1836 -1031 1837 -1007
rect 1892 -1166 1893 -1030
rect 1962 -1166 1963 -1030
rect 2018 -1031 2019 -1007
rect 2130 -1031 2131 -1007
rect 2172 -1166 2173 -1030
rect 177 -1033 178 -1007
rect 2319 -1033 2320 -1007
rect 23 -1035 24 -1007
rect 177 -1166 178 -1034
rect 180 -1035 181 -1007
rect 464 -1035 465 -1007
rect 478 -1166 479 -1034
rect 485 -1035 486 -1007
rect 611 -1035 612 -1007
rect 2221 -1035 2222 -1007
rect 23 -1166 24 -1036
rect 44 -1037 45 -1007
rect 100 -1037 101 -1007
rect 2319 -1166 2320 -1036
rect 44 -1166 45 -1038
rect 240 -1039 241 -1007
rect 261 -1166 262 -1038
rect 275 -1039 276 -1007
rect 310 -1039 311 -1007
rect 880 -1166 881 -1038
rect 919 -1039 920 -1007
rect 919 -1166 920 -1038
rect 919 -1039 920 -1007
rect 919 -1166 920 -1038
rect 940 -1039 941 -1007
rect 1017 -1039 1018 -1007
rect 1024 -1039 1025 -1007
rect 1507 -1166 1508 -1038
rect 1517 -1039 1518 -1007
rect 2263 -1039 2264 -1007
rect 184 -1166 185 -1040
rect 254 -1041 255 -1007
rect 271 -1041 272 -1007
rect 779 -1166 780 -1040
rect 793 -1166 794 -1040
rect 856 -1041 857 -1007
rect 863 -1041 864 -1007
rect 884 -1166 885 -1040
rect 891 -1041 892 -1007
rect 940 -1166 941 -1040
rect 975 -1041 976 -1007
rect 1108 -1166 1109 -1040
rect 1125 -1041 1126 -1007
rect 2088 -1041 2089 -1007
rect 2158 -1041 2159 -1007
rect 2221 -1166 2222 -1040
rect 138 -1166 139 -1042
rect 2158 -1166 2159 -1042
rect 187 -1045 188 -1007
rect 2277 -1045 2278 -1007
rect 191 -1047 192 -1007
rect 310 -1166 311 -1046
rect 324 -1166 325 -1046
rect 681 -1047 682 -1007
rect 723 -1047 724 -1007
rect 975 -1166 976 -1046
rect 989 -1047 990 -1007
rect 1038 -1047 1039 -1007
rect 1041 -1047 1042 -1007
rect 2018 -1166 2019 -1046
rect 2067 -1047 2068 -1007
rect 2130 -1166 2131 -1046
rect 2200 -1047 2201 -1007
rect 2277 -1166 2278 -1046
rect 170 -1049 171 -1007
rect 191 -1166 192 -1048
rect 205 -1049 206 -1007
rect 317 -1166 318 -1048
rect 366 -1049 367 -1007
rect 611 -1166 612 -1048
rect 625 -1049 626 -1007
rect 1731 -1049 1732 -1007
rect 1738 -1049 1739 -1007
rect 1822 -1166 1823 -1048
rect 1843 -1049 1844 -1007
rect 2102 -1166 2103 -1048
rect 2200 -1166 2201 -1048
rect 2249 -1049 2250 -1007
rect 121 -1051 122 -1007
rect 205 -1166 206 -1050
rect 219 -1166 220 -1050
rect 653 -1051 654 -1007
rect 660 -1051 661 -1007
rect 716 -1166 717 -1050
rect 730 -1051 731 -1007
rect 856 -1166 857 -1050
rect 863 -1166 864 -1050
rect 1689 -1166 1690 -1050
rect 1710 -1166 1711 -1050
rect 2361 -1051 2362 -1007
rect 121 -1166 122 -1052
rect 359 -1053 360 -1007
rect 366 -1166 367 -1052
rect 1171 -1053 1172 -1007
rect 1181 -1166 1182 -1052
rect 1626 -1053 1627 -1007
rect 1745 -1053 1746 -1007
rect 1801 -1166 1802 -1052
rect 1843 -1166 1844 -1052
rect 1850 -1053 1851 -1007
rect 1864 -1053 1865 -1007
rect 2137 -1166 2138 -1052
rect 2186 -1053 2187 -1007
rect 2249 -1166 2250 -1052
rect 145 -1166 146 -1054
rect 730 -1166 731 -1054
rect 796 -1055 797 -1007
rect 912 -1055 913 -1007
rect 996 -1055 997 -1007
rect 1202 -1166 1203 -1054
rect 1234 -1055 1235 -1007
rect 1388 -1166 1389 -1054
rect 1437 -1055 1438 -1007
rect 1731 -1166 1732 -1054
rect 1815 -1055 1816 -1007
rect 1850 -1166 1851 -1054
rect 1871 -1166 1872 -1054
rect 1906 -1055 1907 -1007
rect 1983 -1055 1984 -1007
rect 2263 -1166 2264 -1054
rect 170 -1166 171 -1056
rect 376 -1057 377 -1007
rect 380 -1057 381 -1007
rect 775 -1057 776 -1007
rect 817 -1057 818 -1007
rect 1668 -1057 1669 -1007
rect 1675 -1057 1676 -1007
rect 1906 -1166 1907 -1056
rect 1955 -1057 1956 -1007
rect 1983 -1166 1984 -1056
rect 2004 -1057 2005 -1007
rect 2067 -1166 2068 -1056
rect 2186 -1166 2187 -1056
rect 2399 -1166 2400 -1056
rect 79 -1059 80 -1007
rect 380 -1166 381 -1058
rect 387 -1166 388 -1058
rect 814 -1059 815 -1007
rect 831 -1059 832 -1007
rect 2032 -1059 2033 -1007
rect 2039 -1059 2040 -1007
rect 2361 -1166 2362 -1058
rect 79 -1166 80 -1060
rect 114 -1061 115 -1007
rect 222 -1061 223 -1007
rect 618 -1061 619 -1007
rect 639 -1061 640 -1007
rect 723 -1166 724 -1060
rect 775 -1166 776 -1060
rect 968 -1061 969 -1007
rect 982 -1061 983 -1007
rect 996 -1166 997 -1060
rect 1003 -1061 1004 -1007
rect 1171 -1166 1172 -1060
rect 1192 -1061 1193 -1007
rect 2046 -1061 2047 -1007
rect 30 -1063 31 -1007
rect 618 -1166 619 -1062
rect 646 -1166 647 -1062
rect 709 -1063 710 -1007
rect 835 -1063 836 -1007
rect 1122 -1166 1123 -1062
rect 1136 -1063 1137 -1007
rect 1150 -1166 1151 -1062
rect 1157 -1063 1158 -1007
rect 1192 -1166 1193 -1062
rect 1234 -1166 1235 -1062
rect 1836 -1166 1837 -1062
rect 1878 -1063 1879 -1007
rect 2165 -1166 2166 -1062
rect 30 -1166 31 -1064
rect 719 -1065 720 -1007
rect 835 -1166 836 -1064
rect 947 -1065 948 -1007
rect 968 -1166 969 -1064
rect 1073 -1065 1074 -1007
rect 1129 -1065 1130 -1007
rect 1157 -1166 1158 -1064
rect 1237 -1166 1238 -1064
rect 1290 -1065 1291 -1007
rect 1307 -1166 1308 -1064
rect 2004 -1166 2005 -1064
rect 2011 -1065 2012 -1007
rect 2088 -1166 2089 -1064
rect 65 -1067 66 -1007
rect 639 -1166 640 -1066
rect 660 -1166 661 -1066
rect 758 -1067 759 -1007
rect 842 -1166 843 -1066
rect 870 -1067 871 -1007
rect 877 -1067 878 -1007
rect 912 -1166 913 -1066
rect 947 -1166 948 -1066
rect 2256 -1166 2257 -1066
rect 65 -1166 66 -1068
rect 471 -1069 472 -1007
rect 485 -1166 486 -1068
rect 534 -1069 535 -1007
rect 597 -1069 598 -1007
rect 625 -1166 626 -1068
rect 635 -1069 636 -1007
rect 1073 -1166 1074 -1068
rect 1087 -1069 1088 -1007
rect 1129 -1166 1130 -1068
rect 1136 -1166 1137 -1068
rect 1472 -1069 1473 -1007
rect 1479 -1069 1480 -1007
rect 1535 -1166 1536 -1068
rect 1542 -1069 1543 -1007
rect 1626 -1166 1627 -1068
rect 1633 -1069 1634 -1007
rect 1675 -1166 1676 -1068
rect 1815 -1166 1816 -1068
rect 2396 -1166 2397 -1068
rect 226 -1071 227 -1007
rect 464 -1166 465 -1070
rect 513 -1071 514 -1007
rect 814 -1166 815 -1070
rect 891 -1166 892 -1070
rect 898 -1071 899 -1007
rect 1003 -1166 1004 -1070
rect 1024 -1166 1025 -1070
rect 1045 -1071 1046 -1007
rect 1087 -1166 1088 -1070
rect 1241 -1071 1242 -1007
rect 2060 -1071 2061 -1007
rect 51 -1073 52 -1007
rect 513 -1166 514 -1072
rect 534 -1166 535 -1072
rect 1269 -1073 1270 -1007
rect 1272 -1073 1273 -1007
rect 2032 -1166 2033 -1072
rect 2039 -1166 2040 -1072
rect 2347 -1073 2348 -1007
rect 51 -1166 52 -1074
rect 142 -1075 143 -1007
rect 212 -1075 213 -1007
rect 226 -1166 227 -1074
rect 240 -1166 241 -1074
rect 527 -1166 528 -1074
rect 597 -1166 598 -1074
rect 1062 -1075 1063 -1007
rect 1223 -1166 1224 -1074
rect 1241 -1166 1242 -1074
rect 1244 -1075 1245 -1007
rect 2284 -1166 2285 -1074
rect 142 -1166 143 -1076
rect 989 -1166 990 -1076
rect 1010 -1077 1011 -1007
rect 1038 -1166 1039 -1076
rect 1055 -1077 1056 -1007
rect 1549 -1077 1550 -1007
rect 1598 -1077 1599 -1007
rect 1668 -1166 1669 -1076
rect 1829 -1077 1830 -1007
rect 1864 -1166 1865 -1076
rect 1878 -1166 1879 -1076
rect 1927 -1077 1928 -1007
rect 1941 -1077 1942 -1007
rect 1955 -1166 1956 -1076
rect 1969 -1077 1970 -1007
rect 2011 -1166 2012 -1076
rect 2207 -1077 2208 -1007
rect 2347 -1166 2348 -1076
rect 198 -1079 199 -1007
rect 212 -1166 213 -1078
rect 254 -1166 255 -1078
rect 541 -1079 542 -1007
rect 681 -1166 682 -1078
rect 950 -1166 951 -1078
rect 1017 -1166 1018 -1078
rect 1115 -1079 1116 -1007
rect 1248 -1079 1249 -1007
rect 1360 -1166 1361 -1078
rect 1374 -1079 1375 -1007
rect 1437 -1166 1438 -1078
rect 1486 -1079 1487 -1007
rect 1829 -1166 1830 -1078
rect 1927 -1166 1928 -1078
rect 2193 -1079 2194 -1007
rect 198 -1166 199 -1080
rect 807 -1081 808 -1007
rect 877 -1166 878 -1080
rect 1269 -1166 1270 -1080
rect 1283 -1081 1284 -1007
rect 2312 -1081 2313 -1007
rect 275 -1166 276 -1082
rect 415 -1083 416 -1007
rect 429 -1083 430 -1007
rect 1447 -1166 1448 -1082
rect 1500 -1083 1501 -1007
rect 1542 -1166 1543 -1082
rect 1580 -1083 1581 -1007
rect 1941 -1166 1942 -1082
rect 1997 -1083 1998 -1007
rect 2046 -1166 2047 -1082
rect 2109 -1083 2110 -1007
rect 2207 -1166 2208 -1082
rect 2235 -1083 2236 -1007
rect 2312 -1166 2313 -1082
rect 359 -1166 360 -1084
rect 432 -1166 433 -1084
rect 443 -1166 444 -1084
rect 499 -1085 500 -1007
rect 541 -1166 542 -1084
rect 604 -1085 605 -1007
rect 607 -1166 608 -1084
rect 2193 -1166 2194 -1084
rect 114 -1166 115 -1086
rect 499 -1166 500 -1086
rect 604 -1166 605 -1086
rect 1045 -1166 1046 -1086
rect 1059 -1166 1060 -1086
rect 1143 -1087 1144 -1007
rect 1227 -1087 1228 -1007
rect 1248 -1166 1249 -1086
rect 1286 -1087 1287 -1007
rect 1759 -1087 1760 -1007
rect 1808 -1087 1809 -1007
rect 1969 -1166 1970 -1086
rect 2151 -1087 2152 -1007
rect 2235 -1166 2236 -1086
rect 401 -1089 402 -1007
rect 404 -1131 405 -1088
rect 415 -1166 416 -1088
rect 506 -1089 507 -1007
rect 695 -1089 696 -1007
rect 982 -1166 983 -1088
rect 1080 -1089 1081 -1007
rect 1143 -1166 1144 -1088
rect 1213 -1089 1214 -1007
rect 1227 -1166 1228 -1088
rect 1314 -1089 1315 -1007
rect 1640 -1089 1641 -1007
rect 1654 -1089 1655 -1007
rect 1745 -1166 1746 -1088
rect 1857 -1089 1858 -1007
rect 2109 -1166 2110 -1088
rect 401 -1166 402 -1090
rect 408 -1091 409 -1007
rect 429 -1166 430 -1090
rect 1773 -1091 1774 -1007
rect 1794 -1091 1795 -1007
rect 1857 -1166 1858 -1090
rect 2095 -1091 2096 -1007
rect 2151 -1166 2152 -1090
rect 408 -1166 409 -1092
rect 576 -1093 577 -1007
rect 688 -1093 689 -1007
rect 695 -1166 696 -1092
rect 702 -1093 703 -1007
rect 807 -1166 808 -1092
rect 898 -1166 899 -1092
rect 1094 -1093 1095 -1007
rect 1101 -1093 1102 -1007
rect 1115 -1166 1116 -1092
rect 1213 -1166 1214 -1092
rect 2343 -1093 2344 -1007
rect 2 -1095 3 -1007
rect 688 -1166 689 -1094
rect 709 -1166 710 -1094
rect 926 -1095 927 -1007
rect 1031 -1095 1032 -1007
rect 1101 -1166 1102 -1094
rect 1318 -1095 1319 -1007
rect 1451 -1166 1452 -1094
rect 1556 -1095 1557 -1007
rect 1640 -1166 1641 -1094
rect 1696 -1095 1697 -1007
rect 1759 -1166 1760 -1094
rect 2025 -1095 2026 -1007
rect 2095 -1166 2096 -1094
rect 72 -1097 73 -1007
rect 702 -1166 703 -1096
rect 737 -1097 738 -1007
rect 1290 -1166 1291 -1096
rect 1325 -1097 1326 -1007
rect 1374 -1166 1375 -1096
rect 1381 -1097 1382 -1007
rect 1472 -1166 1473 -1096
rect 1598 -1166 1599 -1096
rect 1605 -1097 1606 -1007
rect 1717 -1097 1718 -1007
rect 1773 -1166 1774 -1096
rect 1899 -1097 1900 -1007
rect 2025 -1166 2026 -1096
rect 37 -1099 38 -1007
rect 72 -1166 73 -1098
rect 89 -1166 90 -1098
rect 1094 -1166 1095 -1098
rect 1185 -1099 1186 -1007
rect 1696 -1166 1697 -1098
rect 1717 -1166 1718 -1098
rect 1752 -1099 1753 -1007
rect 1899 -1166 1900 -1098
rect 2333 -1099 2334 -1007
rect 37 -1166 38 -1100
rect 593 -1166 594 -1100
rect 751 -1101 752 -1007
rect 870 -1166 871 -1100
rect 905 -1101 906 -1007
rect 1031 -1166 1032 -1100
rect 1066 -1101 1067 -1007
rect 1080 -1166 1081 -1100
rect 1185 -1166 1186 -1100
rect 1199 -1101 1200 -1007
rect 1206 -1101 1207 -1007
rect 1318 -1166 1319 -1100
rect 1335 -1166 1336 -1100
rect 2305 -1101 2306 -1007
rect 247 -1103 248 -1007
rect 926 -1166 927 -1102
rect 961 -1103 962 -1007
rect 1066 -1166 1067 -1102
rect 1178 -1103 1179 -1007
rect 1206 -1166 1207 -1102
rect 1255 -1103 1256 -1007
rect 1325 -1166 1326 -1102
rect 1367 -1103 1368 -1007
rect 1381 -1166 1382 -1102
rect 1395 -1103 1396 -1007
rect 1752 -1166 1753 -1102
rect 2214 -1103 2215 -1007
rect 2305 -1166 2306 -1102
rect 163 -1105 164 -1007
rect 247 -1166 248 -1104
rect 373 -1105 374 -1007
rect 1178 -1166 1179 -1104
rect 1195 -1105 1196 -1007
rect 1556 -1166 1557 -1104
rect 1724 -1105 1725 -1007
rect 1808 -1166 1809 -1104
rect 2116 -1105 2117 -1007
rect 2214 -1166 2215 -1104
rect 2270 -1105 2271 -1007
rect 2333 -1166 2334 -1104
rect 163 -1166 164 -1106
rect 338 -1107 339 -1007
rect 352 -1107 353 -1007
rect 373 -1166 374 -1106
rect 390 -1107 391 -1007
rect 737 -1166 738 -1106
rect 772 -1166 773 -1106
rect 1633 -1166 1634 -1106
rect 2053 -1107 2054 -1007
rect 2116 -1166 2117 -1106
rect 233 -1109 234 -1007
rect 961 -1166 962 -1108
rect 1052 -1109 1053 -1007
rect 1724 -1166 1725 -1108
rect 2053 -1166 2054 -1108
rect 2336 -1109 2337 -1007
rect 233 -1166 234 -1110
rect 394 -1111 395 -1007
rect 450 -1111 451 -1007
rect 471 -1166 472 -1110
rect 506 -1166 507 -1110
rect 1794 -1166 1795 -1110
rect 107 -1113 108 -1007
rect 394 -1166 395 -1112
rect 450 -1166 451 -1112
rect 492 -1113 493 -1007
rect 548 -1113 549 -1007
rect 576 -1166 577 -1112
rect 674 -1113 675 -1007
rect 751 -1166 752 -1112
rect 786 -1113 787 -1007
rect 1010 -1166 1011 -1112
rect 1199 -1166 1200 -1112
rect 1766 -1113 1767 -1007
rect 107 -1166 108 -1114
rect 2326 -1115 2327 -1007
rect 338 -1166 339 -1116
rect 520 -1117 521 -1007
rect 569 -1117 570 -1007
rect 1052 -1166 1053 -1116
rect 1220 -1117 1221 -1007
rect 1255 -1166 1256 -1116
rect 1262 -1117 1263 -1007
rect 1367 -1166 1368 -1116
rect 1402 -1117 1403 -1007
rect 2060 -1166 2061 -1116
rect 352 -1166 353 -1118
rect 866 -1166 867 -1118
rect 905 -1166 906 -1118
rect 1682 -1166 1683 -1118
rect 1766 -1166 1767 -1118
rect 1780 -1119 1781 -1007
rect 422 -1121 423 -1007
rect 569 -1166 570 -1120
rect 674 -1166 675 -1120
rect 1167 -1166 1168 -1120
rect 1220 -1166 1221 -1120
rect 2270 -1166 2271 -1120
rect 100 -1166 101 -1122
rect 422 -1166 423 -1122
rect 436 -1123 437 -1007
rect 492 -1166 493 -1122
rect 520 -1166 521 -1122
rect 583 -1123 584 -1007
rect 744 -1123 745 -1007
rect 786 -1166 787 -1122
rect 800 -1123 801 -1007
rect 1283 -1166 1284 -1122
rect 1297 -1123 1298 -1007
rect 1395 -1166 1396 -1122
rect 1423 -1123 1424 -1007
rect 1479 -1166 1480 -1122
rect 1549 -1166 1550 -1122
rect 1605 -1166 1606 -1122
rect 1661 -1123 1662 -1007
rect 1780 -1166 1781 -1122
rect 289 -1125 290 -1007
rect 583 -1166 584 -1124
rect 800 -1166 801 -1124
rect 821 -1125 822 -1007
rect 1164 -1125 1165 -1007
rect 1262 -1166 1263 -1124
rect 1297 -1166 1298 -1124
rect 2354 -1125 2355 -1007
rect 289 -1166 290 -1126
rect 296 -1127 297 -1007
rect 436 -1166 437 -1126
rect 656 -1166 657 -1126
rect 821 -1166 822 -1126
rect 1997 -1166 1998 -1126
rect 296 -1166 297 -1128
rect 303 -1129 304 -1007
rect 457 -1129 458 -1007
rect 548 -1166 549 -1128
rect 555 -1129 556 -1007
rect 744 -1166 745 -1128
rect 1164 -1166 1165 -1128
rect 1612 -1129 1613 -1007
rect 1619 -1129 1620 -1007
rect 1661 -1166 1662 -1128
rect 282 -1131 283 -1007
rect 303 -1166 304 -1130
rect 457 -1166 458 -1130
rect 555 -1166 556 -1130
rect 562 -1131 563 -1007
rect 1304 -1131 1305 -1007
rect 1402 -1166 1403 -1130
rect 1416 -1131 1417 -1007
rect 1423 -1166 1424 -1130
rect 1430 -1131 1431 -1007
rect 1486 -1166 1487 -1130
rect 1584 -1131 1585 -1007
rect 1612 -1166 1613 -1130
rect 149 -1133 150 -1007
rect 282 -1166 283 -1132
rect 1304 -1166 1305 -1132
rect 1934 -1133 1935 -1007
rect 149 -1166 150 -1134
rect 425 -1166 426 -1134
rect 1311 -1135 1312 -1007
rect 2326 -1166 2327 -1134
rect 156 -1137 157 -1007
rect 562 -1166 563 -1136
rect 1311 -1166 1312 -1136
rect 1339 -1137 1340 -1007
rect 1398 -1137 1399 -1007
rect 2354 -1166 2355 -1136
rect 96 -1139 97 -1007
rect 156 -1166 157 -1138
rect 824 -1166 825 -1138
rect 1339 -1166 1340 -1138
rect 1430 -1166 1431 -1138
rect 1521 -1139 1522 -1007
rect 1528 -1139 1529 -1007
rect 1584 -1166 1585 -1138
rect 1591 -1139 1592 -1007
rect 1619 -1166 1620 -1138
rect 1934 -1166 1935 -1138
rect 2081 -1139 2082 -1007
rect 632 -1141 633 -1007
rect 1591 -1166 1592 -1140
rect 2081 -1166 2082 -1140
rect 2179 -1141 2180 -1007
rect 632 -1166 633 -1142
rect 1160 -1166 1161 -1142
rect 1444 -1143 1445 -1007
rect 1500 -1166 1501 -1142
rect 2144 -1143 2145 -1007
rect 2179 -1166 2180 -1142
rect 1458 -1145 1459 -1007
rect 1521 -1166 1522 -1144
rect 2074 -1145 2075 -1007
rect 2144 -1166 2145 -1144
rect 1276 -1147 1277 -1007
rect 1458 -1166 1459 -1146
rect 1493 -1147 1494 -1007
rect 1528 -1166 1529 -1146
rect 1976 -1147 1977 -1007
rect 2074 -1166 2075 -1146
rect 828 -1149 829 -1007
rect 1276 -1166 1277 -1148
rect 1465 -1149 1466 -1007
rect 1493 -1166 1494 -1148
rect 1948 -1149 1949 -1007
rect 1976 -1166 1977 -1148
rect 765 -1151 766 -1007
rect 828 -1166 829 -1150
rect 1465 -1166 1466 -1150
rect 1647 -1151 1648 -1007
rect 1920 -1151 1921 -1007
rect 1948 -1166 1949 -1150
rect 765 -1166 766 -1152
rect 849 -1153 850 -1007
rect 1563 -1153 1564 -1007
rect 1647 -1166 1648 -1152
rect 1913 -1153 1914 -1007
rect 1920 -1166 1921 -1152
rect 849 -1166 850 -1154
rect 1416 -1166 1417 -1154
rect 1885 -1155 1886 -1007
rect 1913 -1166 1914 -1154
rect 1353 -1157 1354 -1007
rect 1563 -1166 1564 -1156
rect 1741 -1166 1742 -1156
rect 1885 -1166 1886 -1156
rect 1346 -1159 1347 -1007
rect 1353 -1166 1354 -1158
rect 1332 -1161 1333 -1007
rect 1346 -1166 1347 -1160
rect 957 -1163 958 -1007
rect 1332 -1166 1333 -1162
rect 957 -1166 958 -1164
rect 1654 -1166 1655 -1164
rect 5 -1349 6 -1175
rect 432 -1176 433 -1174
rect 485 -1176 486 -1174
rect 653 -1176 654 -1174
rect 656 -1176 657 -1174
rect 1514 -1176 1515 -1174
rect 1549 -1176 1550 -1174
rect 2291 -1176 2292 -1174
rect 2298 -1176 2299 -1174
rect 2494 -1349 2495 -1175
rect 19 -1349 20 -1177
rect 30 -1178 31 -1174
rect 89 -1178 90 -1174
rect 856 -1178 857 -1174
rect 866 -1178 867 -1174
rect 1031 -1178 1032 -1174
rect 1041 -1349 1042 -1177
rect 2473 -1349 2474 -1177
rect 23 -1180 24 -1174
rect 821 -1180 822 -1174
rect 842 -1180 843 -1174
rect 856 -1349 857 -1179
rect 880 -1180 881 -1174
rect 1745 -1180 1746 -1174
rect 1906 -1180 1907 -1174
rect 2452 -1349 2453 -1179
rect 23 -1349 24 -1181
rect 611 -1182 612 -1174
rect 667 -1182 668 -1174
rect 849 -1349 850 -1181
rect 905 -1349 906 -1181
rect 926 -1182 927 -1174
rect 947 -1182 948 -1174
rect 1433 -1349 1434 -1181
rect 1447 -1182 1448 -1174
rect 2361 -1182 2362 -1174
rect 2368 -1182 2369 -1174
rect 2564 -1349 2565 -1181
rect 30 -1349 31 -1183
rect 677 -1349 678 -1183
rect 751 -1184 752 -1174
rect 842 -1349 843 -1183
rect 912 -1184 913 -1174
rect 1031 -1349 1032 -1183
rect 1048 -1184 1049 -1174
rect 1122 -1184 1123 -1174
rect 1157 -1184 1158 -1174
rect 2263 -1184 2264 -1174
rect 2277 -1184 2278 -1174
rect 2466 -1349 2467 -1183
rect 100 -1186 101 -1174
rect 908 -1186 909 -1174
rect 947 -1349 948 -1185
rect 1094 -1186 1095 -1174
rect 1104 -1349 1105 -1185
rect 2543 -1349 2544 -1185
rect 100 -1349 101 -1187
rect 247 -1188 248 -1174
rect 254 -1188 255 -1174
rect 912 -1349 913 -1187
rect 950 -1188 951 -1174
rect 1451 -1188 1452 -1174
rect 1458 -1188 1459 -1174
rect 1549 -1349 1550 -1187
rect 1552 -1188 1553 -1174
rect 1598 -1188 1599 -1174
rect 1605 -1188 1606 -1174
rect 1906 -1349 1907 -1187
rect 1927 -1188 1928 -1174
rect 2459 -1349 2460 -1187
rect 121 -1190 122 -1174
rect 509 -1190 510 -1174
rect 513 -1190 514 -1174
rect 611 -1349 612 -1189
rect 667 -1349 668 -1189
rect 1269 -1190 1270 -1174
rect 1307 -1190 1308 -1174
rect 2396 -1190 2397 -1174
rect 2431 -1190 2432 -1174
rect 2578 -1349 2579 -1189
rect 124 -1349 125 -1191
rect 1290 -1192 1291 -1174
rect 1335 -1192 1336 -1174
rect 2347 -1192 2348 -1174
rect 2354 -1192 2355 -1174
rect 2557 -1349 2558 -1191
rect 128 -1194 129 -1174
rect 1927 -1349 1928 -1193
rect 1969 -1194 1970 -1174
rect 2389 -1194 2390 -1174
rect 2438 -1194 2439 -1174
rect 2480 -1349 2481 -1193
rect 128 -1349 129 -1195
rect 268 -1196 269 -1174
rect 275 -1196 276 -1174
rect 782 -1349 783 -1195
rect 796 -1349 797 -1195
rect 968 -1196 969 -1174
rect 982 -1196 983 -1174
rect 1094 -1349 1095 -1195
rect 1115 -1196 1116 -1174
rect 1269 -1349 1270 -1195
rect 1339 -1196 1340 -1174
rect 1458 -1349 1459 -1195
rect 1500 -1196 1501 -1174
rect 1598 -1349 1599 -1195
rect 1605 -1349 1606 -1195
rect 1612 -1196 1613 -1174
rect 1745 -1349 1746 -1195
rect 1801 -1196 1802 -1174
rect 2060 -1196 2061 -1174
rect 2263 -1349 2264 -1195
rect 2284 -1196 2285 -1174
rect 2487 -1349 2488 -1195
rect 138 -1198 139 -1174
rect 583 -1198 584 -1174
rect 590 -1198 591 -1174
rect 1815 -1198 1816 -1174
rect 1857 -1198 1858 -1174
rect 2060 -1349 2061 -1197
rect 2095 -1198 2096 -1174
rect 2291 -1349 2292 -1197
rect 2305 -1198 2306 -1174
rect 2501 -1349 2502 -1197
rect 208 -1349 209 -1199
rect 730 -1200 731 -1174
rect 751 -1349 752 -1199
rect 884 -1200 885 -1174
rect 992 -1349 993 -1199
rect 2431 -1349 2432 -1199
rect 37 -1202 38 -1174
rect 884 -1349 885 -1201
rect 1003 -1202 1004 -1174
rect 1829 -1202 1830 -1174
rect 1962 -1202 1963 -1174
rect 2284 -1349 2285 -1201
rect 2312 -1202 2313 -1174
rect 2508 -1349 2509 -1201
rect 37 -1349 38 -1203
rect 702 -1204 703 -1174
rect 758 -1204 759 -1174
rect 1514 -1349 1515 -1203
rect 1521 -1204 1522 -1174
rect 1612 -1349 1613 -1203
rect 1668 -1204 1669 -1174
rect 1829 -1349 1830 -1203
rect 2109 -1204 2110 -1174
rect 2298 -1349 2299 -1203
rect 2319 -1204 2320 -1174
rect 2515 -1349 2516 -1203
rect 268 -1349 269 -1205
rect 2375 -1206 2376 -1174
rect 2424 -1206 2425 -1174
rect 2438 -1349 2439 -1205
rect 275 -1349 276 -1207
rect 2343 -1349 2344 -1207
rect 310 -1210 311 -1174
rect 968 -1349 969 -1209
rect 1003 -1349 1004 -1209
rect 2270 -1210 2271 -1174
rect 2333 -1210 2334 -1174
rect 2536 -1349 2537 -1209
rect 72 -1212 73 -1174
rect 310 -1349 311 -1211
rect 380 -1212 381 -1174
rect 429 -1349 430 -1211
rect 436 -1212 437 -1174
rect 513 -1349 514 -1211
rect 527 -1212 528 -1174
rect 583 -1349 584 -1211
rect 604 -1349 605 -1211
rect 821 -1349 822 -1211
rect 828 -1212 829 -1174
rect 926 -1349 927 -1211
rect 1010 -1212 1011 -1174
rect 1115 -1349 1116 -1211
rect 1164 -1212 1165 -1174
rect 2382 -1212 2383 -1174
rect 72 -1349 73 -1213
rect 443 -1214 444 -1174
rect 485 -1349 486 -1213
rect 548 -1214 549 -1174
rect 555 -1214 556 -1174
rect 590 -1349 591 -1213
rect 642 -1349 643 -1213
rect 1857 -1349 1858 -1213
rect 1920 -1214 1921 -1174
rect 2109 -1349 2110 -1213
rect 2116 -1214 2117 -1174
rect 2305 -1349 2306 -1213
rect 2340 -1214 2341 -1174
rect 2550 -1349 2551 -1213
rect 9 -1216 10 -1174
rect 555 -1349 556 -1215
rect 569 -1216 570 -1174
rect 653 -1349 654 -1215
rect 702 -1349 703 -1215
rect 957 -1349 958 -1215
rect 1038 -1216 1039 -1174
rect 1157 -1349 1158 -1215
rect 1167 -1216 1168 -1174
rect 2571 -1349 2572 -1215
rect 9 -1349 10 -1217
rect 135 -1218 136 -1174
rect 219 -1218 220 -1174
rect 1164 -1349 1165 -1217
rect 1178 -1218 1179 -1174
rect 1843 -1218 1844 -1174
rect 1934 -1218 1935 -1174
rect 2319 -1349 2320 -1217
rect 16 -1220 17 -1174
rect 443 -1349 444 -1219
rect 499 -1220 500 -1174
rect 730 -1349 731 -1219
rect 758 -1349 759 -1219
rect 786 -1220 787 -1174
rect 800 -1220 801 -1174
rect 894 -1349 895 -1219
rect 1045 -1220 1046 -1174
rect 1122 -1349 1123 -1219
rect 1185 -1220 1186 -1174
rect 1339 -1349 1340 -1219
rect 1370 -1349 1371 -1219
rect 2102 -1220 2103 -1174
rect 2116 -1349 2117 -1219
rect 2256 -1220 2257 -1174
rect 65 -1222 66 -1174
rect 569 -1349 570 -1221
rect 772 -1222 773 -1174
rect 772 -1349 773 -1221
rect 772 -1222 773 -1174
rect 772 -1349 773 -1221
rect 800 -1349 801 -1221
rect 1038 -1349 1039 -1221
rect 1045 -1349 1046 -1221
rect 1101 -1222 1102 -1174
rect 1192 -1222 1193 -1174
rect 1290 -1349 1291 -1221
rect 1311 -1222 1312 -1174
rect 1500 -1349 1501 -1221
rect 1563 -1222 1564 -1174
rect 2529 -1349 2530 -1221
rect 65 -1349 66 -1223
rect 79 -1224 80 -1174
rect 114 -1224 115 -1174
rect 2102 -1349 2103 -1223
rect 2144 -1224 2145 -1174
rect 2312 -1349 2313 -1223
rect 114 -1349 115 -1225
rect 646 -1226 647 -1174
rect 807 -1226 808 -1174
rect 810 -1288 811 -1225
rect 852 -1226 853 -1174
rect 1801 -1349 1802 -1225
rect 1815 -1349 1816 -1225
rect 1892 -1226 1893 -1174
rect 1948 -1226 1949 -1174
rect 2144 -1349 2145 -1225
rect 2151 -1226 2152 -1174
rect 2333 -1349 2334 -1225
rect 135 -1349 136 -1227
rect 681 -1228 682 -1174
rect 789 -1349 790 -1227
rect 1948 -1349 1949 -1227
rect 1955 -1228 1956 -1174
rect 2151 -1349 2152 -1227
rect 2158 -1228 2159 -1174
rect 2347 -1349 2348 -1227
rect 191 -1230 192 -1174
rect 219 -1349 220 -1229
rect 373 -1230 374 -1174
rect 499 -1349 500 -1229
rect 506 -1230 507 -1174
rect 2445 -1349 2446 -1229
rect 191 -1349 192 -1231
rect 387 -1232 388 -1174
rect 408 -1232 409 -1174
rect 607 -1232 608 -1174
rect 646 -1349 647 -1231
rect 1087 -1232 1088 -1174
rect 1192 -1349 1193 -1231
rect 1262 -1232 1263 -1174
rect 1283 -1232 1284 -1174
rect 1563 -1349 1564 -1231
rect 1570 -1232 1571 -1174
rect 1668 -1349 1669 -1231
rect 1731 -1232 1732 -1174
rect 1892 -1349 1893 -1231
rect 1955 -1349 1956 -1231
rect 2067 -1232 2068 -1174
rect 2088 -1232 2089 -1174
rect 2256 -1349 2257 -1231
rect 198 -1234 199 -1174
rect 1087 -1349 1088 -1233
rect 1234 -1234 1235 -1174
rect 2410 -1349 2411 -1233
rect 149 -1236 150 -1174
rect 1234 -1349 1235 -1235
rect 1255 -1236 1256 -1174
rect 1262 -1349 1263 -1235
rect 1283 -1349 1284 -1235
rect 1353 -1236 1354 -1174
rect 1381 -1236 1382 -1174
rect 1391 -1236 1392 -1174
rect 1416 -1236 1417 -1174
rect 1521 -1349 1522 -1235
rect 1591 -1236 1592 -1174
rect 1731 -1349 1732 -1235
rect 1738 -1236 1739 -1174
rect 2270 -1349 2271 -1235
rect 145 -1238 146 -1174
rect 149 -1349 150 -1237
rect 198 -1349 199 -1237
rect 1360 -1238 1361 -1174
rect 1381 -1349 1382 -1237
rect 1619 -1238 1620 -1174
rect 1633 -1238 1634 -1174
rect 1738 -1349 1739 -1237
rect 1741 -1238 1742 -1174
rect 2067 -1349 2068 -1237
rect 2172 -1238 2173 -1174
rect 2354 -1349 2355 -1237
rect 233 -1240 234 -1174
rect 408 -1349 409 -1239
rect 422 -1240 423 -1174
rect 1794 -1240 1795 -1174
rect 1885 -1240 1886 -1174
rect 2088 -1349 2089 -1239
rect 2179 -1240 2180 -1174
rect 2361 -1349 2362 -1239
rect 226 -1242 227 -1174
rect 233 -1349 234 -1241
rect 261 -1242 262 -1174
rect 422 -1349 423 -1241
rect 436 -1349 437 -1241
rect 674 -1242 675 -1174
rect 681 -1349 682 -1241
rect 744 -1242 745 -1174
rect 807 -1349 808 -1241
rect 1304 -1242 1305 -1174
rect 1332 -1242 1333 -1174
rect 1962 -1349 1963 -1241
rect 1983 -1242 1984 -1174
rect 2158 -1349 2159 -1241
rect 2186 -1242 2187 -1174
rect 2368 -1349 2369 -1241
rect 261 -1349 262 -1243
rect 1010 -1349 1011 -1243
rect 1059 -1244 1060 -1174
rect 1220 -1244 1221 -1174
rect 1241 -1244 1242 -1174
rect 1353 -1349 1354 -1243
rect 1384 -1349 1385 -1243
rect 2207 -1244 2208 -1174
rect 2221 -1244 2222 -1174
rect 2382 -1349 2383 -1243
rect 303 -1246 304 -1174
rect 373 -1349 374 -1245
rect 380 -1349 381 -1245
rect 457 -1246 458 -1174
rect 506 -1349 507 -1245
rect 723 -1246 724 -1174
rect 744 -1349 745 -1245
rect 954 -1246 955 -1174
rect 961 -1246 962 -1174
rect 1633 -1349 1634 -1245
rect 1654 -1246 1655 -1174
rect 1794 -1349 1795 -1245
rect 1990 -1246 1991 -1174
rect 2179 -1349 2180 -1245
rect 2193 -1246 2194 -1174
rect 2375 -1349 2376 -1245
rect 229 -1349 230 -1247
rect 457 -1349 458 -1247
rect 527 -1349 528 -1247
rect 831 -1349 832 -1247
rect 877 -1248 878 -1174
rect 2095 -1349 2096 -1247
rect 2200 -1248 2201 -1174
rect 2522 -1349 2523 -1247
rect 303 -1349 304 -1249
rect 534 -1250 535 -1174
rect 548 -1349 549 -1249
rect 1181 -1250 1182 -1174
rect 1206 -1250 1207 -1174
rect 1304 -1349 1305 -1249
rect 1325 -1250 1326 -1174
rect 1332 -1349 1333 -1249
rect 1416 -1349 1417 -1249
rect 2123 -1250 2124 -1174
rect 2137 -1250 2138 -1174
rect 2200 -1349 2201 -1249
rect 2228 -1250 2229 -1174
rect 2389 -1349 2390 -1249
rect 331 -1252 332 -1174
rect 387 -1349 388 -1251
rect 520 -1252 521 -1174
rect 534 -1349 535 -1251
rect 562 -1252 563 -1174
rect 786 -1349 787 -1251
rect 891 -1252 892 -1174
rect 961 -1349 962 -1251
rect 975 -1252 976 -1174
rect 1059 -1349 1060 -1251
rect 1073 -1252 1074 -1174
rect 1178 -1349 1179 -1251
rect 1241 -1349 1242 -1251
rect 1248 -1252 1249 -1174
rect 1255 -1349 1256 -1251
rect 1388 -1252 1389 -1174
rect 1423 -1252 1424 -1174
rect 1570 -1349 1571 -1251
rect 1591 -1349 1592 -1251
rect 1724 -1252 1725 -1174
rect 1759 -1252 1760 -1174
rect 1920 -1349 1921 -1251
rect 2004 -1252 2005 -1174
rect 2186 -1349 2187 -1251
rect 2242 -1252 2243 -1174
rect 2396 -1349 2397 -1251
rect 205 -1254 206 -1174
rect 520 -1349 521 -1253
rect 562 -1349 563 -1253
rect 639 -1254 640 -1174
rect 660 -1254 661 -1174
rect 1220 -1349 1221 -1253
rect 1276 -1254 1277 -1174
rect 1388 -1349 1389 -1253
rect 1447 -1349 1448 -1253
rect 2165 -1254 2166 -1174
rect 2249 -1254 2250 -1174
rect 2424 -1349 2425 -1253
rect 205 -1349 206 -1255
rect 2074 -1256 2075 -1174
rect 282 -1258 283 -1174
rect 331 -1349 332 -1257
rect 607 -1349 608 -1257
rect 814 -1258 815 -1174
rect 863 -1349 864 -1257
rect 2242 -1349 2243 -1257
rect 282 -1349 283 -1259
rect 464 -1260 465 -1174
rect 541 -1260 542 -1174
rect 814 -1349 815 -1259
rect 898 -1260 899 -1174
rect 975 -1349 976 -1259
rect 985 -1349 986 -1259
rect 1983 -1349 1984 -1259
rect 2004 -1349 2005 -1259
rect 2130 -1260 2131 -1174
rect 93 -1262 94 -1174
rect 898 -1349 899 -1261
rect 919 -1262 920 -1174
rect 1185 -1349 1186 -1261
rect 1276 -1349 1277 -1261
rect 1297 -1262 1298 -1174
rect 1367 -1262 1368 -1174
rect 1423 -1349 1424 -1261
rect 1451 -1349 1452 -1261
rect 1696 -1262 1697 -1174
rect 1703 -1262 1704 -1174
rect 1885 -1349 1886 -1261
rect 1913 -1262 1914 -1174
rect 2123 -1349 2124 -1261
rect 86 -1264 87 -1174
rect 93 -1349 94 -1263
rect 110 -1264 111 -1174
rect 1703 -1349 1704 -1263
rect 1752 -1264 1753 -1174
rect 1913 -1349 1914 -1263
rect 2018 -1264 2019 -1174
rect 2193 -1349 2194 -1263
rect 86 -1349 87 -1265
rect 597 -1266 598 -1174
rect 632 -1266 633 -1174
rect 674 -1349 675 -1265
rect 709 -1266 710 -1174
rect 919 -1349 920 -1265
rect 954 -1349 955 -1265
rect 964 -1266 965 -1174
rect 1073 -1349 1074 -1265
rect 1216 -1349 1217 -1265
rect 1325 -1349 1326 -1265
rect 1367 -1349 1368 -1265
rect 1402 -1266 1403 -1174
rect 2165 -1349 2166 -1265
rect 44 -1268 45 -1174
rect 709 -1349 710 -1267
rect 723 -1349 724 -1267
rect 1941 -1268 1942 -1174
rect 2032 -1268 2033 -1174
rect 2228 -1349 2229 -1267
rect 44 -1349 45 -1269
rect 324 -1270 325 -1174
rect 464 -1349 465 -1269
rect 835 -1270 836 -1174
rect 1080 -1270 1081 -1174
rect 1206 -1349 1207 -1269
rect 1402 -1349 1403 -1269
rect 1409 -1270 1410 -1174
rect 1507 -1270 1508 -1174
rect 1752 -1349 1753 -1269
rect 1766 -1270 1767 -1174
rect 2018 -1349 2019 -1269
rect 2039 -1270 2040 -1174
rect 2221 -1349 2222 -1269
rect 243 -1272 244 -1174
rect 324 -1349 325 -1271
rect 541 -1349 542 -1271
rect 618 -1272 619 -1174
rect 625 -1272 626 -1174
rect 632 -1349 633 -1271
rect 639 -1349 640 -1271
rect 2417 -1349 2418 -1271
rect 597 -1349 598 -1273
rect 880 -1349 881 -1273
rect 989 -1274 990 -1174
rect 1080 -1349 1081 -1273
rect 1143 -1274 1144 -1174
rect 1360 -1349 1361 -1273
rect 1528 -1274 1529 -1174
rect 1619 -1349 1620 -1273
rect 1626 -1274 1627 -1174
rect 1759 -1349 1760 -1273
rect 1773 -1274 1774 -1174
rect 1941 -1349 1942 -1273
rect 2046 -1274 2047 -1174
rect 2249 -1349 2250 -1273
rect 142 -1276 143 -1174
rect 2046 -1349 2047 -1275
rect 2053 -1276 2054 -1174
rect 2207 -1349 2208 -1275
rect 142 -1349 143 -1277
rect 824 -1278 825 -1174
rect 989 -1349 990 -1277
rect 1136 -1278 1137 -1174
rect 1626 -1349 1627 -1277
rect 1640 -1278 1641 -1174
rect 1766 -1349 1767 -1277
rect 1780 -1278 1781 -1174
rect 1934 -1349 1935 -1277
rect 2011 -1278 2012 -1174
rect 2053 -1349 2054 -1277
rect 618 -1349 619 -1279
rect 1199 -1280 1200 -1174
rect 1227 -1280 1228 -1174
rect 1409 -1349 1410 -1279
rect 1535 -1280 1536 -1174
rect 1640 -1349 1641 -1279
rect 1647 -1280 1648 -1174
rect 1773 -1349 1774 -1279
rect 1780 -1349 1781 -1279
rect 1976 -1280 1977 -1174
rect 625 -1349 626 -1281
rect 779 -1282 780 -1174
rect 996 -1282 997 -1174
rect 1136 -1349 1137 -1281
rect 1143 -1349 1144 -1281
rect 1160 -1282 1161 -1174
rect 1171 -1282 1172 -1174
rect 1227 -1349 1228 -1281
rect 1237 -1282 1238 -1174
rect 1647 -1349 1648 -1281
rect 1661 -1282 1662 -1174
rect 1843 -1349 1844 -1281
rect 1850 -1282 1851 -1174
rect 2039 -1349 2040 -1281
rect 660 -1349 661 -1283
rect 891 -1349 892 -1283
rect 996 -1349 997 -1283
rect 2172 -1349 2173 -1283
rect 688 -1286 689 -1174
rect 835 -1349 836 -1285
rect 999 -1349 1000 -1285
rect 1199 -1349 1200 -1285
rect 1311 -1349 1312 -1285
rect 1507 -1349 1508 -1285
rect 1542 -1286 1543 -1174
rect 1654 -1349 1655 -1285
rect 1717 -1286 1718 -1174
rect 2011 -1349 2012 -1285
rect 688 -1349 689 -1287
rect 866 -1349 867 -1287
rect 1052 -1288 1053 -1174
rect 1171 -1349 1172 -1287
rect 1391 -1349 1392 -1287
rect 1528 -1349 1529 -1287
rect 1556 -1288 1557 -1174
rect 1661 -1349 1662 -1287
rect 1787 -1288 1788 -1174
rect 2277 -1349 2278 -1287
rect 765 -1290 766 -1174
rect 1248 -1349 1249 -1289
rect 1430 -1290 1431 -1174
rect 1717 -1349 1718 -1289
rect 1808 -1290 1809 -1174
rect 1990 -1349 1991 -1289
rect 695 -1292 696 -1174
rect 765 -1349 766 -1291
rect 1024 -1292 1025 -1174
rect 1052 -1349 1053 -1291
rect 1150 -1292 1151 -1174
rect 1297 -1349 1298 -1291
rect 1430 -1349 1431 -1291
rect 1969 -1349 1970 -1291
rect 695 -1349 696 -1293
rect 940 -1294 941 -1174
rect 1024 -1349 1025 -1293
rect 1066 -1294 1067 -1174
rect 1108 -1294 1109 -1174
rect 1150 -1349 1151 -1293
rect 1213 -1294 1214 -1174
rect 1787 -1349 1788 -1293
rect 1836 -1294 1837 -1174
rect 2032 -1349 2033 -1293
rect 51 -1296 52 -1174
rect 940 -1349 941 -1295
rect 1108 -1349 1109 -1295
rect 1129 -1296 1130 -1174
rect 1153 -1349 1154 -1295
rect 1836 -1349 1837 -1295
rect 1850 -1349 1851 -1295
rect 2392 -1296 2393 -1174
rect 51 -1349 52 -1297
rect 58 -1298 59 -1174
rect 450 -1298 451 -1174
rect 1066 -1349 1067 -1297
rect 1213 -1349 1214 -1297
rect 2214 -1298 2215 -1174
rect 58 -1349 59 -1299
rect 79 -1349 80 -1299
rect 450 -1349 451 -1299
rect 576 -1300 577 -1174
rect 1017 -1300 1018 -1174
rect 1129 -1349 1130 -1299
rect 1444 -1300 1445 -1174
rect 1535 -1349 1536 -1299
rect 1556 -1349 1557 -1299
rect 2403 -1300 2404 -1174
rect 352 -1302 353 -1174
rect 576 -1349 577 -1301
rect 933 -1302 934 -1174
rect 1017 -1349 1018 -1301
rect 1479 -1302 1480 -1174
rect 1976 -1349 1977 -1301
rect 2025 -1302 2026 -1174
rect 2214 -1349 2215 -1301
rect 352 -1349 353 -1303
rect 401 -1304 402 -1174
rect 793 -1304 794 -1174
rect 933 -1349 934 -1303
rect 1013 -1349 1014 -1303
rect 2025 -1349 2026 -1303
rect 2081 -1304 2082 -1174
rect 2403 -1349 2404 -1303
rect 394 -1306 395 -1174
rect 401 -1349 402 -1305
rect 761 -1306 762 -1174
rect 2081 -1349 2082 -1305
rect 212 -1308 213 -1174
rect 394 -1349 395 -1307
rect 793 -1349 794 -1307
rect 1997 -1308 1998 -1174
rect 212 -1349 213 -1309
rect 415 -1310 416 -1174
rect 1395 -1310 1396 -1174
rect 1479 -1349 1480 -1309
rect 1493 -1310 1494 -1174
rect 1542 -1349 1543 -1309
rect 1577 -1310 1578 -1174
rect 1696 -1349 1697 -1309
rect 1864 -1310 1865 -1174
rect 2074 -1349 2075 -1309
rect 170 -1312 171 -1174
rect 415 -1349 416 -1311
rect 1006 -1312 1007 -1174
rect 1864 -1349 1865 -1311
rect 1871 -1312 1872 -1174
rect 2130 -1349 2131 -1311
rect 107 -1349 108 -1313
rect 1006 -1349 1007 -1313
rect 1346 -1314 1347 -1174
rect 1493 -1349 1494 -1313
rect 1584 -1314 1585 -1174
rect 1724 -1349 1725 -1313
rect 1878 -1314 1879 -1174
rect 2137 -1349 2138 -1313
rect 170 -1349 171 -1315
rect 737 -1316 738 -1174
rect 1395 -1349 1396 -1315
rect 1437 -1316 1438 -1174
rect 1465 -1316 1466 -1174
rect 1878 -1349 1879 -1315
rect 247 -1349 248 -1317
rect 1346 -1349 1347 -1317
rect 1472 -1318 1473 -1174
rect 1577 -1349 1578 -1317
rect 1675 -1318 1676 -1174
rect 1808 -1349 1809 -1317
rect 716 -1320 717 -1174
rect 737 -1349 738 -1319
rect 779 -1349 780 -1319
rect 1465 -1349 1466 -1319
rect 1472 -1349 1473 -1319
rect 1710 -1320 1711 -1174
rect 359 -1322 360 -1174
rect 716 -1349 717 -1321
rect 1318 -1322 1319 -1174
rect 1437 -1349 1438 -1321
rect 1486 -1322 1487 -1174
rect 1584 -1349 1585 -1321
rect 1675 -1349 1676 -1321
rect 2235 -1322 2236 -1174
rect 163 -1324 164 -1174
rect 359 -1349 360 -1323
rect 1202 -1324 1203 -1174
rect 1318 -1349 1319 -1323
rect 1374 -1324 1375 -1174
rect 1486 -1349 1487 -1323
rect 1510 -1349 1511 -1323
rect 2235 -1349 2236 -1323
rect 156 -1326 157 -1174
rect 163 -1349 164 -1325
rect 177 -1326 178 -1174
rect 1374 -1349 1375 -1325
rect 1682 -1326 1683 -1174
rect 1871 -1349 1872 -1325
rect 156 -1349 157 -1327
rect 240 -1328 241 -1174
rect 1682 -1349 1683 -1327
rect 2326 -1328 2327 -1174
rect 177 -1349 178 -1329
rect 184 -1330 185 -1174
rect 240 -1349 241 -1329
rect 296 -1330 297 -1174
rect 1689 -1330 1690 -1174
rect 1997 -1349 1998 -1329
rect 184 -1349 185 -1331
rect 289 -1332 290 -1174
rect 296 -1349 297 -1331
rect 478 -1332 479 -1174
rect 1101 -1349 1102 -1331
rect 1689 -1349 1690 -1331
rect 1710 -1349 1711 -1331
rect 1899 -1332 1900 -1174
rect 289 -1349 290 -1333
rect 471 -1334 472 -1174
rect 1822 -1334 1823 -1174
rect 2326 -1349 2327 -1333
rect 317 -1336 318 -1174
rect 478 -1349 479 -1335
rect 828 -1349 829 -1335
rect 1822 -1349 1823 -1335
rect 1899 -1349 1900 -1335
rect 2340 -1349 2341 -1335
rect 317 -1349 318 -1337
rect 726 -1349 727 -1337
rect 366 -1340 367 -1174
rect 471 -1349 472 -1339
rect 345 -1342 346 -1174
rect 366 -1349 367 -1341
rect 345 -1349 346 -1343
rect 492 -1344 493 -1174
rect 338 -1346 339 -1174
rect 492 -1349 493 -1345
rect 121 -1349 122 -1347
rect 338 -1349 339 -1347
rect 2 -1359 3 -1357
rect 838 -1359 839 -1357
rect 880 -1359 881 -1357
rect 1136 -1359 1137 -1357
rect 1150 -1359 1151 -1357
rect 2263 -1359 2264 -1357
rect 2343 -1359 2344 -1357
rect 2578 -1359 2579 -1357
rect 26 -1526 27 -1360
rect 1577 -1361 1578 -1357
rect 1794 -1361 1795 -1357
rect 1797 -1361 1798 -1357
rect 2263 -1526 2264 -1360
rect 2361 -1361 2362 -1357
rect 37 -1363 38 -1357
rect 989 -1363 990 -1357
rect 996 -1363 997 -1357
rect 1717 -1363 1718 -1357
rect 1794 -1526 1795 -1362
rect 1850 -1363 1851 -1357
rect 2361 -1526 2362 -1362
rect 2424 -1363 2425 -1357
rect 40 -1526 41 -1364
rect 1983 -1365 1984 -1357
rect 44 -1367 45 -1357
rect 201 -1526 202 -1366
rect 208 -1367 209 -1357
rect 436 -1367 437 -1357
rect 464 -1367 465 -1357
rect 908 -1526 909 -1366
rect 943 -1526 944 -1366
rect 1976 -1367 1977 -1357
rect 1983 -1526 1984 -1366
rect 2368 -1367 2369 -1357
rect 44 -1526 45 -1368
rect 86 -1369 87 -1357
rect 89 -1526 90 -1368
rect 968 -1369 969 -1357
rect 989 -1526 990 -1368
rect 1115 -1369 1116 -1357
rect 1129 -1369 1130 -1357
rect 1129 -1526 1130 -1368
rect 1129 -1369 1130 -1357
rect 1129 -1526 1130 -1368
rect 1136 -1526 1137 -1368
rect 1192 -1369 1193 -1357
rect 1213 -1369 1214 -1357
rect 1556 -1369 1557 -1357
rect 1577 -1526 1578 -1368
rect 1605 -1369 1606 -1357
rect 1717 -1526 1718 -1368
rect 1766 -1369 1767 -1357
rect 1850 -1526 1851 -1368
rect 1913 -1369 1914 -1357
rect 1976 -1526 1977 -1368
rect 2039 -1369 2040 -1357
rect 2368 -1526 2369 -1368
rect 2431 -1369 2432 -1357
rect 54 -1526 55 -1370
rect 86 -1526 87 -1370
rect 93 -1371 94 -1357
rect 124 -1371 125 -1357
rect 163 -1371 164 -1357
rect 163 -1526 164 -1370
rect 163 -1371 164 -1357
rect 163 -1526 164 -1370
rect 170 -1371 171 -1357
rect 268 -1526 269 -1370
rect 282 -1371 283 -1357
rect 282 -1526 283 -1370
rect 282 -1371 283 -1357
rect 282 -1526 283 -1370
rect 317 -1371 318 -1357
rect 464 -1526 465 -1370
rect 499 -1371 500 -1357
rect 628 -1526 629 -1370
rect 642 -1371 643 -1357
rect 968 -1526 969 -1370
rect 996 -1526 997 -1370
rect 1500 -1371 1501 -1357
rect 1507 -1526 1508 -1370
rect 1773 -1371 1774 -1357
rect 1913 -1526 1914 -1370
rect 1962 -1371 1963 -1357
rect 2431 -1526 2432 -1370
rect 2480 -1371 2481 -1357
rect 58 -1373 59 -1357
rect 61 -1383 62 -1372
rect 72 -1373 73 -1357
rect 824 -1526 825 -1372
rect 831 -1373 832 -1357
rect 905 -1373 906 -1357
rect 957 -1373 958 -1357
rect 1423 -1373 1424 -1357
rect 1426 -1526 1427 -1372
rect 1864 -1373 1865 -1357
rect 1962 -1526 1963 -1372
rect 2032 -1373 2033 -1357
rect 58 -1526 59 -1374
rect 79 -1526 80 -1374
rect 156 -1375 157 -1357
rect 170 -1526 171 -1374
rect 236 -1526 237 -1374
rect 240 -1375 241 -1357
rect 639 -1375 640 -1357
rect 646 -1375 647 -1357
rect 954 -1375 955 -1357
rect 982 -1375 983 -1357
rect 2480 -1526 2481 -1374
rect 82 -1377 83 -1357
rect 1752 -1377 1753 -1357
rect 1766 -1526 1767 -1376
rect 2109 -1377 2110 -1357
rect 93 -1526 94 -1378
rect 296 -1379 297 -1357
rect 317 -1526 318 -1378
rect 887 -1526 888 -1378
rect 891 -1379 892 -1357
rect 2529 -1379 2530 -1357
rect 107 -1381 108 -1357
rect 604 -1381 605 -1357
rect 646 -1526 647 -1380
rect 653 -1381 654 -1357
rect 681 -1381 682 -1357
rect 999 -1381 1000 -1357
rect 1006 -1381 1007 -1357
rect 1433 -1381 1434 -1357
rect 1472 -1381 1473 -1357
rect 1752 -1526 1753 -1380
rect 1773 -1526 1774 -1380
rect 1822 -1381 1823 -1357
rect 1864 -1526 1865 -1380
rect 1920 -1381 1921 -1357
rect 2109 -1526 2110 -1380
rect 2193 -1381 2194 -1357
rect 2529 -1526 2530 -1380
rect 2557 -1381 2558 -1357
rect 110 -1526 111 -1382
rect 1787 -1383 1788 -1357
rect 1797 -1526 1798 -1382
rect 2032 -1526 2033 -1382
rect 2193 -1526 2194 -1382
rect 2291 -1383 2292 -1357
rect 2340 -1383 2341 -1357
rect 2557 -1526 2558 -1382
rect 117 -1526 118 -1384
rect 208 -1526 209 -1384
rect 226 -1385 227 -1357
rect 1374 -1385 1375 -1357
rect 1430 -1385 1431 -1357
rect 1871 -1385 1872 -1357
rect 2200 -1385 2201 -1357
rect 2340 -1526 2341 -1384
rect 121 -1387 122 -1357
rect 1234 -1387 1235 -1357
rect 1251 -1526 1252 -1386
rect 2326 -1387 2327 -1357
rect 107 -1526 108 -1388
rect 121 -1526 122 -1388
rect 128 -1389 129 -1357
rect 653 -1526 654 -1388
rect 681 -1526 682 -1388
rect 737 -1389 738 -1357
rect 772 -1389 773 -1357
rect 782 -1389 783 -1357
rect 796 -1389 797 -1357
rect 912 -1389 913 -1357
rect 954 -1526 955 -1388
rect 975 -1389 976 -1357
rect 982 -1526 983 -1388
rect 1073 -1389 1074 -1357
rect 1087 -1389 1088 -1357
rect 1192 -1526 1193 -1388
rect 1213 -1526 1214 -1388
rect 1227 -1389 1228 -1357
rect 1234 -1526 1235 -1388
rect 1304 -1389 1305 -1357
rect 1332 -1389 1333 -1357
rect 1430 -1526 1431 -1388
rect 1472 -1526 1473 -1388
rect 1486 -1389 1487 -1357
rect 1500 -1526 1501 -1388
rect 2270 -1389 2271 -1357
rect 128 -1526 129 -1390
rect 992 -1391 993 -1357
rect 1013 -1391 1014 -1357
rect 1759 -1391 1760 -1357
rect 1787 -1526 1788 -1390
rect 1836 -1391 1837 -1357
rect 1871 -1526 1872 -1390
rect 1934 -1391 1935 -1357
rect 2200 -1526 2201 -1390
rect 2508 -1391 2509 -1357
rect 226 -1526 227 -1392
rect 485 -1393 486 -1357
rect 516 -1526 517 -1392
rect 569 -1393 570 -1357
rect 723 -1526 724 -1392
rect 1090 -1526 1091 -1392
rect 1104 -1393 1105 -1357
rect 1675 -1393 1676 -1357
rect 1759 -1526 1760 -1392
rect 1815 -1393 1816 -1357
rect 1822 -1526 1823 -1392
rect 1892 -1393 1893 -1357
rect 1934 -1526 1935 -1392
rect 1997 -1393 1998 -1357
rect 2270 -1526 2271 -1392
rect 2382 -1393 2383 -1357
rect 2508 -1526 2509 -1392
rect 2522 -1393 2523 -1357
rect 229 -1395 230 -1357
rect 1920 -1526 1921 -1394
rect 1997 -1526 1998 -1394
rect 2074 -1395 2075 -1357
rect 2116 -1395 2117 -1357
rect 2382 -1526 2383 -1394
rect 2522 -1526 2523 -1394
rect 2543 -1395 2544 -1357
rect 240 -1526 241 -1396
rect 751 -1397 752 -1357
rect 772 -1526 773 -1396
rect 842 -1397 843 -1357
rect 880 -1526 881 -1396
rect 919 -1397 920 -1357
rect 1038 -1397 1039 -1357
rect 1360 -1397 1361 -1357
rect 1370 -1397 1371 -1357
rect 2424 -1526 2425 -1396
rect 2543 -1526 2544 -1396
rect 2571 -1397 2572 -1357
rect 254 -1399 255 -1357
rect 688 -1399 689 -1357
rect 726 -1399 727 -1357
rect 866 -1399 867 -1357
rect 891 -1526 892 -1398
rect 961 -1399 962 -1357
rect 1031 -1399 1032 -1357
rect 1038 -1526 1039 -1398
rect 1041 -1399 1042 -1357
rect 2165 -1399 2166 -1357
rect 254 -1526 255 -1400
rect 618 -1401 619 -1357
rect 688 -1526 689 -1400
rect 758 -1401 759 -1357
rect 779 -1401 780 -1357
rect 1878 -1401 1879 -1357
rect 2165 -1526 2166 -1400
rect 2256 -1401 2257 -1357
rect 296 -1526 297 -1402
rect 894 -1403 895 -1357
rect 898 -1403 899 -1357
rect 975 -1526 976 -1402
rect 1066 -1403 1067 -1357
rect 1101 -1403 1102 -1357
rect 1115 -1526 1116 -1402
rect 1297 -1403 1298 -1357
rect 1304 -1526 1305 -1402
rect 1451 -1403 1452 -1357
rect 1482 -1526 1483 -1402
rect 2123 -1403 2124 -1357
rect 2256 -1526 2257 -1402
rect 2354 -1403 2355 -1357
rect 16 -1405 17 -1357
rect 1451 -1526 1452 -1404
rect 1510 -1405 1511 -1357
rect 2277 -1405 2278 -1357
rect 16 -1526 17 -1406
rect 2116 -1526 2117 -1406
rect 2123 -1526 2124 -1406
rect 2207 -1407 2208 -1357
rect 2277 -1526 2278 -1406
rect 2410 -1407 2411 -1357
rect 310 -1409 311 -1357
rect 604 -1526 605 -1408
rect 618 -1526 619 -1408
rect 702 -1409 703 -1357
rect 730 -1409 731 -1357
rect 740 -1526 741 -1408
rect 758 -1526 759 -1408
rect 870 -1409 871 -1357
rect 905 -1526 906 -1408
rect 2039 -1526 2040 -1408
rect 2207 -1526 2208 -1408
rect 2445 -1409 2446 -1357
rect 184 -1411 185 -1357
rect 310 -1526 311 -1410
rect 387 -1411 388 -1357
rect 387 -1526 388 -1410
rect 387 -1411 388 -1357
rect 387 -1526 388 -1410
rect 408 -1411 409 -1357
rect 863 -1526 864 -1410
rect 866 -1526 867 -1410
rect 2130 -1411 2131 -1357
rect 2410 -1526 2411 -1410
rect 2459 -1411 2460 -1357
rect 184 -1526 185 -1412
rect 275 -1413 276 -1357
rect 366 -1413 367 -1357
rect 408 -1526 409 -1412
rect 415 -1413 416 -1357
rect 607 -1413 608 -1357
rect 642 -1526 643 -1412
rect 2354 -1526 2355 -1412
rect 2445 -1526 2446 -1412
rect 2494 -1413 2495 -1357
rect 257 -1415 258 -1357
rect 415 -1526 416 -1414
rect 422 -1415 423 -1357
rect 593 -1526 594 -1414
rect 702 -1526 703 -1414
rect 1178 -1415 1179 -1357
rect 1227 -1526 1228 -1414
rect 1248 -1415 1249 -1357
rect 1258 -1526 1259 -1414
rect 2172 -1415 2173 -1357
rect 219 -1417 220 -1357
rect 422 -1526 423 -1416
rect 429 -1417 430 -1357
rect 569 -1526 570 -1416
rect 730 -1526 731 -1416
rect 1349 -1526 1350 -1416
rect 1384 -1417 1385 -1357
rect 1675 -1526 1676 -1416
rect 1682 -1417 1683 -1357
rect 2494 -1526 2495 -1416
rect 19 -1526 20 -1418
rect 429 -1526 430 -1418
rect 436 -1526 437 -1418
rect 1311 -1419 1312 -1357
rect 1332 -1526 1333 -1418
rect 1353 -1419 1354 -1357
rect 1556 -1526 1557 -1418
rect 1584 -1419 1585 -1357
rect 1591 -1419 1592 -1357
rect 1892 -1526 1893 -1418
rect 2172 -1526 2173 -1418
rect 2242 -1419 2243 -1357
rect 149 -1421 150 -1357
rect 219 -1526 220 -1420
rect 247 -1421 248 -1357
rect 1682 -1526 1683 -1420
rect 1780 -1421 1781 -1357
rect 2074 -1526 2075 -1420
rect 2242 -1526 2243 -1420
rect 2333 -1421 2334 -1357
rect 149 -1526 150 -1422
rect 765 -1423 766 -1357
rect 789 -1423 790 -1357
rect 2459 -1526 2460 -1422
rect 247 -1526 248 -1424
rect 352 -1425 353 -1357
rect 366 -1526 367 -1424
rect 492 -1425 493 -1357
rect 506 -1425 507 -1357
rect 751 -1526 752 -1424
rect 765 -1526 766 -1424
rect 1171 -1425 1172 -1357
rect 1178 -1526 1179 -1424
rect 1290 -1425 1291 -1357
rect 1297 -1526 1298 -1424
rect 1325 -1425 1326 -1357
rect 1353 -1526 1354 -1424
rect 1493 -1425 1494 -1357
rect 1584 -1526 1585 -1424
rect 1885 -1425 1886 -1357
rect 142 -1427 143 -1357
rect 1290 -1526 1291 -1426
rect 1311 -1526 1312 -1426
rect 1339 -1427 1340 -1357
rect 1591 -1526 1592 -1426
rect 1633 -1427 1634 -1357
rect 1780 -1526 1781 -1426
rect 1829 -1427 1830 -1357
rect 1836 -1526 1837 -1426
rect 1899 -1427 1900 -1357
rect 142 -1526 143 -1428
rect 985 -1429 986 -1357
rect 1003 -1429 1004 -1357
rect 1325 -1526 1326 -1428
rect 1605 -1526 1606 -1428
rect 1647 -1429 1648 -1357
rect 1815 -1526 1816 -1428
rect 1857 -1429 1858 -1357
rect 1878 -1526 1879 -1428
rect 1955 -1429 1956 -1357
rect 275 -1526 276 -1430
rect 359 -1431 360 -1357
rect 471 -1431 472 -1357
rect 506 -1526 507 -1430
rect 541 -1431 542 -1357
rect 1010 -1431 1011 -1357
rect 1024 -1431 1025 -1357
rect 1101 -1526 1102 -1430
rect 1150 -1526 1151 -1430
rect 1185 -1431 1186 -1357
rect 1241 -1431 1242 -1357
rect 1339 -1526 1340 -1430
rect 1619 -1431 1620 -1357
rect 1829 -1526 1830 -1430
rect 1857 -1526 1858 -1430
rect 1927 -1431 1928 -1357
rect 1955 -1526 1956 -1430
rect 2025 -1431 2026 -1357
rect 289 -1433 290 -1357
rect 492 -1526 493 -1432
rect 541 -1526 542 -1432
rect 1419 -1433 1420 -1357
rect 1489 -1526 1490 -1432
rect 1619 -1526 1620 -1432
rect 1633 -1526 1634 -1432
rect 1668 -1433 1669 -1357
rect 1885 -1526 1886 -1432
rect 1948 -1433 1949 -1357
rect 2025 -1526 2026 -1432
rect 2095 -1433 2096 -1357
rect 289 -1526 290 -1434
rect 548 -1435 549 -1357
rect 555 -1435 556 -1357
rect 779 -1526 780 -1434
rect 814 -1435 815 -1357
rect 1087 -1526 1088 -1434
rect 1153 -1435 1154 -1357
rect 2291 -1526 2292 -1434
rect 135 -1437 136 -1357
rect 548 -1526 549 -1436
rect 716 -1437 717 -1357
rect 1003 -1526 1004 -1436
rect 1010 -1526 1011 -1436
rect 1052 -1437 1053 -1357
rect 1059 -1437 1060 -1357
rect 1066 -1526 1067 -1436
rect 1185 -1526 1186 -1436
rect 1206 -1437 1207 -1357
rect 1241 -1526 1242 -1436
rect 1262 -1437 1263 -1357
rect 1283 -1437 1284 -1357
rect 1360 -1526 1361 -1436
rect 1647 -1526 1648 -1436
rect 1689 -1437 1690 -1357
rect 1899 -1526 1900 -1436
rect 2179 -1437 2180 -1357
rect 135 -1526 136 -1438
rect 667 -1439 668 -1357
rect 716 -1526 717 -1438
rect 828 -1439 829 -1357
rect 835 -1439 836 -1357
rect 1073 -1526 1074 -1438
rect 1206 -1526 1207 -1438
rect 1220 -1439 1221 -1357
rect 1248 -1526 1249 -1438
rect 2326 -1526 2327 -1438
rect 250 -1441 251 -1357
rect 1220 -1526 1221 -1440
rect 1255 -1441 1256 -1357
rect 1493 -1526 1494 -1440
rect 1668 -1526 1669 -1440
rect 1724 -1441 1725 -1357
rect 1927 -1526 1928 -1440
rect 2004 -1441 2005 -1357
rect 2067 -1441 2068 -1357
rect 2179 -1526 2180 -1440
rect 261 -1443 262 -1357
rect 555 -1526 556 -1442
rect 677 -1443 678 -1357
rect 1255 -1526 1256 -1442
rect 1262 -1526 1263 -1442
rect 1269 -1443 1270 -1357
rect 1283 -1526 1284 -1442
rect 1941 -1443 1942 -1357
rect 1948 -1526 1949 -1442
rect 2018 -1443 2019 -1357
rect 261 -1526 262 -1444
rect 520 -1445 521 -1357
rect 674 -1445 675 -1357
rect 1269 -1526 1270 -1444
rect 1381 -1445 1382 -1357
rect 1689 -1526 1690 -1444
rect 1941 -1526 1942 -1444
rect 2011 -1445 2012 -1357
rect 2018 -1526 2019 -1444
rect 2088 -1445 2089 -1357
rect 9 -1447 10 -1357
rect 520 -1526 521 -1446
rect 674 -1526 675 -1446
rect 691 -1526 692 -1446
rect 737 -1526 738 -1446
rect 2130 -1526 2131 -1446
rect 9 -1526 10 -1448
rect 1265 -1526 1266 -1448
rect 1381 -1526 1382 -1448
rect 1388 -1449 1389 -1357
rect 1503 -1526 1504 -1448
rect 1724 -1526 1725 -1448
rect 1969 -1449 1970 -1357
rect 2095 -1526 2096 -1448
rect 303 -1451 304 -1357
rect 359 -1526 360 -1450
rect 450 -1451 451 -1357
rect 667 -1526 668 -1450
rect 744 -1451 745 -1357
rect 1052 -1526 1053 -1450
rect 1388 -1526 1389 -1450
rect 1402 -1451 1403 -1357
rect 1514 -1451 1515 -1357
rect 2067 -1526 2068 -1450
rect 2088 -1526 2089 -1450
rect 2186 -1451 2187 -1357
rect 177 -1453 178 -1357
rect 303 -1526 304 -1452
rect 352 -1526 353 -1452
rect 373 -1453 374 -1357
rect 450 -1526 451 -1452
rect 597 -1453 598 -1357
rect 709 -1453 710 -1357
rect 744 -1526 745 -1452
rect 786 -1453 787 -1357
rect 2186 -1526 2187 -1452
rect 177 -1526 178 -1454
rect 191 -1455 192 -1357
rect 271 -1455 272 -1357
rect 709 -1526 710 -1454
rect 786 -1526 787 -1454
rect 947 -1455 948 -1357
rect 1024 -1526 1025 -1454
rect 1164 -1455 1165 -1357
rect 1276 -1455 1277 -1357
rect 1402 -1526 1403 -1454
rect 1969 -1526 1970 -1454
rect 2060 -1455 2061 -1357
rect 191 -1526 192 -1456
rect 345 -1457 346 -1357
rect 373 -1526 374 -1456
rect 401 -1457 402 -1357
rect 443 -1457 444 -1357
rect 597 -1526 598 -1456
rect 660 -1457 661 -1357
rect 947 -1526 948 -1456
rect 1031 -1526 1032 -1456
rect 1153 -1526 1154 -1456
rect 1157 -1457 1158 -1357
rect 1514 -1526 1515 -1456
rect 2004 -1526 2005 -1456
rect 2249 -1457 2250 -1357
rect 331 -1459 332 -1357
rect 345 -1526 346 -1458
rect 401 -1526 402 -1458
rect 1286 -1526 1287 -1458
rect 2011 -1526 2012 -1458
rect 2081 -1459 2082 -1357
rect 2249 -1526 2250 -1458
rect 2347 -1459 2348 -1357
rect 331 -1526 332 -1460
rect 590 -1461 591 -1357
rect 632 -1461 633 -1357
rect 660 -1526 661 -1460
rect 814 -1526 815 -1460
rect 926 -1461 927 -1357
rect 940 -1461 941 -1357
rect 1059 -1526 1060 -1460
rect 1122 -1461 1123 -1357
rect 1276 -1526 1277 -1460
rect 2060 -1526 2061 -1460
rect 2151 -1461 2152 -1357
rect 2347 -1526 2348 -1460
rect 2417 -1461 2418 -1357
rect 114 -1463 115 -1357
rect 632 -1526 633 -1462
rect 828 -1526 829 -1462
rect 1612 -1463 1613 -1357
rect 2081 -1526 2082 -1462
rect 2158 -1463 2159 -1357
rect 2417 -1526 2418 -1462
rect 2473 -1463 2474 -1357
rect 51 -1465 52 -1357
rect 114 -1526 115 -1464
rect 443 -1526 444 -1464
rect 796 -1526 797 -1464
rect 835 -1526 836 -1464
rect 849 -1465 850 -1357
rect 856 -1465 857 -1357
rect 898 -1526 899 -1464
rect 912 -1526 913 -1464
rect 1444 -1465 1445 -1357
rect 1612 -1526 1613 -1464
rect 1654 -1465 1655 -1357
rect 2151 -1526 2152 -1464
rect 2228 -1465 2229 -1357
rect 2473 -1526 2474 -1464
rect 2515 -1465 2516 -1357
rect 51 -1526 52 -1466
rect 842 -1526 843 -1466
rect 870 -1526 871 -1466
rect 884 -1467 885 -1357
rect 919 -1526 920 -1466
rect 1017 -1467 1018 -1357
rect 1122 -1526 1123 -1466
rect 1143 -1467 1144 -1357
rect 1157 -1526 1158 -1466
rect 2452 -1467 2453 -1357
rect 2515 -1526 2516 -1466
rect 2536 -1467 2537 -1357
rect 471 -1526 472 -1468
rect 800 -1469 801 -1357
rect 884 -1526 885 -1468
rect 1563 -1469 1564 -1357
rect 1654 -1526 1655 -1468
rect 1696 -1469 1697 -1357
rect 2158 -1526 2159 -1468
rect 2235 -1469 2236 -1357
rect 2452 -1526 2453 -1468
rect 2501 -1469 2502 -1357
rect 2536 -1526 2537 -1468
rect 2550 -1469 2551 -1357
rect 338 -1471 339 -1357
rect 800 -1526 801 -1470
rect 926 -1526 927 -1470
rect 933 -1471 934 -1357
rect 940 -1526 941 -1470
rect 2333 -1526 2334 -1470
rect 2375 -1471 2376 -1357
rect 2550 -1526 2551 -1470
rect 205 -1473 206 -1357
rect 933 -1526 934 -1472
rect 1017 -1526 1018 -1472
rect 2144 -1473 2145 -1357
rect 2228 -1526 2229 -1472
rect 2312 -1473 2313 -1357
rect 338 -1526 339 -1474
rect 457 -1475 458 -1357
rect 478 -1475 479 -1357
rect 499 -1526 500 -1474
rect 562 -1475 563 -1357
rect 856 -1526 857 -1474
rect 877 -1475 878 -1357
rect 2375 -1526 2376 -1474
rect 23 -1477 24 -1357
rect 562 -1526 563 -1476
rect 625 -1477 626 -1357
rect 849 -1526 850 -1476
rect 1143 -1526 1144 -1476
rect 1521 -1477 1522 -1357
rect 1563 -1526 1564 -1476
rect 1598 -1477 1599 -1357
rect 1696 -1526 1697 -1476
rect 1731 -1477 1732 -1357
rect 1990 -1477 1991 -1357
rect 2235 -1526 2236 -1476
rect 2312 -1526 2313 -1476
rect 2396 -1477 2397 -1357
rect 2 -1526 3 -1478
rect 625 -1526 626 -1478
rect 793 -1526 794 -1478
rect 1731 -1526 1732 -1478
rect 1990 -1526 1991 -1478
rect 2298 -1479 2299 -1357
rect 2396 -1526 2397 -1478
rect 2466 -1479 2467 -1357
rect 23 -1526 24 -1480
rect 2102 -1481 2103 -1357
rect 2144 -1526 2145 -1480
rect 2221 -1481 2222 -1357
rect 2284 -1481 2285 -1357
rect 2466 -1526 2467 -1480
rect 156 -1526 157 -1482
rect 877 -1526 878 -1482
rect 1160 -1526 1161 -1482
rect 1444 -1526 1445 -1482
rect 1486 -1526 1487 -1482
rect 2501 -1526 2502 -1482
rect 380 -1485 381 -1357
rect 457 -1526 458 -1484
rect 485 -1526 486 -1484
rect 513 -1485 514 -1357
rect 1164 -1526 1165 -1484
rect 1199 -1485 1200 -1357
rect 1521 -1526 1522 -1484
rect 1542 -1485 1543 -1357
rect 1598 -1526 1599 -1484
rect 1640 -1485 1641 -1357
rect 2046 -1485 2047 -1357
rect 2221 -1526 2222 -1484
rect 2284 -1526 2285 -1484
rect 2564 -1485 2565 -1357
rect 47 -1526 48 -1486
rect 513 -1526 514 -1486
rect 1080 -1487 1081 -1357
rect 1199 -1526 1200 -1486
rect 1367 -1487 1368 -1357
rect 1640 -1526 1641 -1486
rect 2046 -1526 2047 -1486
rect 2137 -1487 2138 -1357
rect 2298 -1526 2299 -1486
rect 2389 -1487 2390 -1357
rect 212 -1489 213 -1357
rect 380 -1526 381 -1488
rect 394 -1489 395 -1357
rect 478 -1526 479 -1488
rect 821 -1489 822 -1357
rect 1367 -1526 1368 -1488
rect 1542 -1526 1543 -1488
rect 1549 -1489 1550 -1357
rect 2053 -1489 2054 -1357
rect 2102 -1526 2103 -1488
rect 2137 -1526 2138 -1488
rect 2214 -1489 2215 -1357
rect 2389 -1526 2390 -1488
rect 2438 -1489 2439 -1357
rect 212 -1526 213 -1490
rect 807 -1491 808 -1357
rect 1080 -1526 1081 -1490
rect 1094 -1491 1095 -1357
rect 1549 -1526 1550 -1490
rect 1570 -1491 1571 -1357
rect 1801 -1491 1802 -1357
rect 2053 -1526 2054 -1490
rect 2214 -1526 2215 -1490
rect 2305 -1491 2306 -1357
rect 2438 -1526 2439 -1490
rect 2487 -1491 2488 -1357
rect 37 -1526 38 -1492
rect 2487 -1526 2488 -1492
rect 394 -1526 395 -1494
rect 534 -1495 535 -1357
rect 807 -1526 808 -1494
rect 1374 -1526 1375 -1494
rect 1535 -1495 1536 -1357
rect 2305 -1526 2306 -1494
rect 324 -1497 325 -1357
rect 534 -1526 535 -1496
rect 1094 -1526 1095 -1496
rect 1108 -1497 1109 -1357
rect 1395 -1497 1396 -1357
rect 1535 -1526 1536 -1496
rect 1570 -1526 1571 -1496
rect 1626 -1497 1627 -1357
rect 1801 -1526 1802 -1496
rect 1843 -1497 1844 -1357
rect 324 -1526 325 -1498
rect 611 -1499 612 -1357
rect 1045 -1499 1046 -1357
rect 1108 -1526 1109 -1498
rect 1395 -1526 1396 -1498
rect 1409 -1499 1410 -1357
rect 1626 -1526 1627 -1498
rect 1661 -1499 1662 -1357
rect 1843 -1526 1844 -1498
rect 1906 -1499 1907 -1357
rect 583 -1501 584 -1357
rect 611 -1526 612 -1500
rect 695 -1501 696 -1357
rect 1045 -1526 1046 -1500
rect 1409 -1526 1410 -1500
rect 1528 -1501 1529 -1357
rect 1661 -1526 1662 -1500
rect 1703 -1501 1704 -1357
rect 1745 -1501 1746 -1357
rect 1906 -1526 1907 -1500
rect 30 -1503 31 -1357
rect 583 -1526 584 -1502
rect 639 -1526 640 -1502
rect 1528 -1526 1529 -1502
rect 1703 -1526 1704 -1502
rect 1738 -1503 1739 -1357
rect 1745 -1526 1746 -1502
rect 1808 -1503 1809 -1357
rect 30 -1526 31 -1504
rect 527 -1505 528 -1357
rect 1416 -1505 1417 -1357
rect 1808 -1526 1809 -1504
rect 100 -1507 101 -1357
rect 527 -1526 528 -1506
rect 1416 -1526 1417 -1506
rect 1437 -1507 1438 -1357
rect 1710 -1507 1711 -1357
rect 1738 -1526 1739 -1506
rect 100 -1526 101 -1508
rect 198 -1509 199 -1357
rect 233 -1509 234 -1357
rect 695 -1526 696 -1508
rect 1437 -1526 1438 -1508
rect 1458 -1509 1459 -1357
rect 72 -1526 73 -1510
rect 233 -1526 234 -1510
rect 576 -1511 577 -1357
rect 1710 -1526 1711 -1510
rect 198 -1526 199 -1512
rect 1171 -1526 1172 -1512
rect 1458 -1526 1459 -1512
rect 1465 -1513 1466 -1357
rect 576 -1526 577 -1514
rect 961 -1526 962 -1514
rect 1465 -1526 1466 -1514
rect 1479 -1515 1480 -1357
rect 1318 -1517 1319 -1357
rect 1479 -1526 1480 -1516
rect 1318 -1526 1319 -1518
rect 1346 -1519 1347 -1357
rect 1346 -1526 1347 -1520
rect 2319 -1521 2320 -1357
rect 2319 -1526 2320 -1522
rect 2403 -1523 2404 -1357
rect 1678 -1525 1679 -1357
rect 2403 -1526 2404 -1524
rect 16 -1699 17 -1535
rect 89 -1536 90 -1534
rect 93 -1536 94 -1534
rect 208 -1536 209 -1534
rect 229 -1699 230 -1535
rect 1710 -1536 1711 -1534
rect 1836 -1536 1837 -1534
rect 1836 -1699 1837 -1535
rect 1836 -1536 1837 -1534
rect 1836 -1699 1837 -1535
rect 1885 -1536 1886 -1534
rect 1885 -1699 1886 -1535
rect 1885 -1536 1886 -1534
rect 1885 -1699 1886 -1535
rect 2389 -1536 2390 -1534
rect 2427 -1699 2428 -1535
rect 2431 -1536 2432 -1534
rect 2434 -1699 2435 -1535
rect 23 -1538 24 -1534
rect 499 -1538 500 -1534
rect 583 -1538 584 -1534
rect 793 -1538 794 -1534
rect 807 -1538 808 -1534
rect 1332 -1538 1333 -1534
rect 1360 -1538 1361 -1534
rect 1440 -1699 1441 -1537
rect 1479 -1538 1480 -1534
rect 1976 -1538 1977 -1534
rect 2284 -1538 2285 -1534
rect 2389 -1699 2390 -1537
rect 23 -1699 24 -1539
rect 628 -1540 629 -1534
rect 642 -1540 643 -1534
rect 709 -1540 710 -1534
rect 719 -1699 720 -1539
rect 2305 -1540 2306 -1534
rect 40 -1542 41 -1534
rect 828 -1542 829 -1534
rect 859 -1699 860 -1541
rect 1493 -1542 1494 -1534
rect 1496 -1699 1497 -1541
rect 2536 -1542 2537 -1534
rect 44 -1544 45 -1534
rect 54 -1662 55 -1543
rect 58 -1544 59 -1534
rect 58 -1699 59 -1543
rect 58 -1544 59 -1534
rect 58 -1699 59 -1543
rect 72 -1544 73 -1534
rect 936 -1699 937 -1543
rect 943 -1544 944 -1534
rect 1640 -1544 1641 -1534
rect 1710 -1699 1711 -1543
rect 1822 -1544 1823 -1534
rect 1976 -1699 1977 -1543
rect 2088 -1544 2089 -1534
rect 2284 -1699 2285 -1543
rect 2417 -1544 2418 -1534
rect 44 -1699 45 -1545
rect 100 -1546 101 -1534
rect 107 -1699 108 -1545
rect 810 -1546 811 -1534
rect 821 -1546 822 -1534
rect 2032 -1546 2033 -1534
rect 2305 -1699 2306 -1545
rect 2438 -1546 2439 -1534
rect 47 -1548 48 -1534
rect 422 -1548 423 -1534
rect 481 -1699 482 -1547
rect 527 -1548 528 -1534
rect 583 -1699 584 -1547
rect 660 -1548 661 -1534
rect 691 -1548 692 -1534
rect 814 -1548 815 -1534
rect 821 -1699 822 -1547
rect 1143 -1548 1144 -1534
rect 1150 -1548 1151 -1534
rect 1584 -1548 1585 -1534
rect 1822 -1699 1823 -1547
rect 1906 -1548 1907 -1534
rect 1990 -1548 1991 -1534
rect 2088 -1699 2089 -1547
rect 2340 -1548 2341 -1534
rect 2438 -1699 2439 -1547
rect 30 -1550 31 -1534
rect 422 -1699 423 -1549
rect 527 -1699 528 -1549
rect 779 -1550 780 -1534
rect 793 -1699 794 -1549
rect 989 -1550 990 -1534
rect 1076 -1699 1077 -1549
rect 2403 -1550 2404 -1534
rect 30 -1699 31 -1551
rect 282 -1552 283 -1534
rect 310 -1552 311 -1534
rect 310 -1699 311 -1551
rect 310 -1552 311 -1534
rect 310 -1699 311 -1551
rect 366 -1552 367 -1534
rect 499 -1699 500 -1551
rect 590 -1552 591 -1534
rect 604 -1552 605 -1534
rect 625 -1552 626 -1534
rect 2053 -1552 2054 -1534
rect 2403 -1699 2404 -1551
rect 2515 -1552 2516 -1534
rect 51 -1554 52 -1534
rect 303 -1554 304 -1534
rect 366 -1699 367 -1553
rect 408 -1554 409 -1534
rect 590 -1699 591 -1553
rect 618 -1554 619 -1534
rect 625 -1699 626 -1553
rect 849 -1554 850 -1534
rect 880 -1554 881 -1534
rect 1514 -1554 1515 -1534
rect 1538 -1699 1539 -1553
rect 2123 -1554 2124 -1534
rect 51 -1699 52 -1555
rect 65 -1556 66 -1534
rect 72 -1699 73 -1555
rect 261 -1556 262 -1534
rect 268 -1556 269 -1534
rect 796 -1556 797 -1534
rect 814 -1699 815 -1555
rect 1038 -1556 1039 -1534
rect 1090 -1556 1091 -1534
rect 2410 -1556 2411 -1534
rect 2 -1558 3 -1534
rect 261 -1699 262 -1557
rect 268 -1699 269 -1557
rect 723 -1558 724 -1534
rect 730 -1558 731 -1534
rect 1020 -1699 1021 -1557
rect 1038 -1699 1039 -1557
rect 1220 -1558 1221 -1534
rect 1248 -1558 1249 -1534
rect 2347 -1558 2348 -1534
rect 65 -1699 66 -1559
rect 429 -1560 430 -1534
rect 597 -1560 598 -1534
rect 597 -1699 598 -1559
rect 597 -1560 598 -1534
rect 597 -1699 598 -1559
rect 604 -1699 605 -1559
rect 1206 -1560 1207 -1534
rect 1220 -1699 1221 -1559
rect 1311 -1560 1312 -1534
rect 1332 -1699 1333 -1559
rect 1605 -1560 1606 -1534
rect 1878 -1560 1879 -1534
rect 2053 -1699 2054 -1559
rect 2123 -1699 2124 -1559
rect 2242 -1560 2243 -1534
rect 2347 -1699 2348 -1559
rect 2473 -1560 2474 -1534
rect 79 -1562 80 -1534
rect 709 -1699 710 -1561
rect 723 -1699 724 -1561
rect 1066 -1562 1067 -1534
rect 1094 -1562 1095 -1534
rect 1094 -1699 1095 -1561
rect 1094 -1562 1095 -1534
rect 1094 -1699 1095 -1561
rect 1129 -1562 1130 -1534
rect 1206 -1699 1207 -1561
rect 1248 -1699 1249 -1561
rect 1395 -1562 1396 -1534
rect 1402 -1562 1403 -1534
rect 2417 -1699 2418 -1561
rect 79 -1699 80 -1563
rect 226 -1564 227 -1534
rect 233 -1564 234 -1534
rect 520 -1564 521 -1534
rect 646 -1564 647 -1534
rect 660 -1699 661 -1563
rect 698 -1699 699 -1563
rect 2340 -1699 2341 -1563
rect 100 -1699 101 -1565
rect 471 -1566 472 -1534
rect 520 -1699 521 -1565
rect 681 -1566 682 -1534
rect 702 -1566 703 -1534
rect 884 -1699 885 -1565
rect 887 -1566 888 -1534
rect 1024 -1566 1025 -1534
rect 1066 -1699 1067 -1565
rect 1171 -1566 1172 -1534
rect 1192 -1566 1193 -1534
rect 1251 -1566 1252 -1534
rect 1255 -1699 1256 -1565
rect 1297 -1566 1298 -1534
rect 1311 -1699 1312 -1565
rect 1458 -1566 1459 -1534
rect 1479 -1699 1480 -1565
rect 1521 -1566 1522 -1534
rect 1584 -1699 1585 -1565
rect 1675 -1566 1676 -1534
rect 1878 -1699 1879 -1565
rect 1969 -1566 1970 -1534
rect 1990 -1699 1991 -1565
rect 2060 -1566 2061 -1534
rect 2095 -1566 2096 -1534
rect 2242 -1699 2243 -1565
rect 37 -1568 38 -1534
rect 1024 -1699 1025 -1567
rect 1111 -1699 1112 -1567
rect 1675 -1699 1676 -1567
rect 1906 -1699 1907 -1567
rect 2018 -1568 2019 -1534
rect 2032 -1699 2033 -1567
rect 2144 -1568 2145 -1534
rect 37 -1699 38 -1569
rect 1612 -1570 1613 -1534
rect 1955 -1570 1956 -1534
rect 2018 -1699 2019 -1569
rect 2095 -1699 2096 -1569
rect 2214 -1570 2215 -1534
rect 121 -1572 122 -1534
rect 460 -1699 461 -1571
rect 471 -1699 472 -1571
rect 506 -1572 507 -1534
rect 534 -1572 535 -1534
rect 681 -1699 682 -1571
rect 702 -1699 703 -1571
rect 751 -1572 752 -1534
rect 779 -1699 780 -1571
rect 870 -1572 871 -1534
rect 898 -1572 899 -1534
rect 940 -1572 941 -1534
rect 961 -1572 962 -1534
rect 2172 -1572 2173 -1534
rect 2214 -1699 2215 -1571
rect 2326 -1572 2327 -1534
rect 114 -1574 115 -1534
rect 751 -1699 752 -1573
rect 824 -1574 825 -1534
rect 877 -1699 878 -1573
rect 898 -1699 899 -1573
rect 1010 -1574 1011 -1534
rect 1129 -1699 1130 -1573
rect 1234 -1574 1235 -1534
rect 1283 -1699 1284 -1573
rect 1304 -1574 1305 -1534
rect 1360 -1699 1361 -1573
rect 1864 -1574 1865 -1534
rect 1955 -1699 1956 -1573
rect 2067 -1574 2068 -1534
rect 2172 -1699 2173 -1573
rect 2291 -1574 2292 -1534
rect 2326 -1699 2327 -1573
rect 2445 -1574 2446 -1534
rect 114 -1699 115 -1575
rect 201 -1576 202 -1534
rect 212 -1576 213 -1534
rect 646 -1699 647 -1575
rect 737 -1576 738 -1534
rect 1269 -1576 1270 -1534
rect 1297 -1699 1298 -1575
rect 1353 -1576 1354 -1534
rect 1395 -1699 1396 -1575
rect 1829 -1576 1830 -1534
rect 1864 -1699 1865 -1575
rect 1941 -1576 1942 -1534
rect 1969 -1699 1970 -1575
rect 2081 -1576 2082 -1534
rect 2291 -1699 2292 -1575
rect 2361 -1576 2362 -1534
rect 2445 -1699 2446 -1575
rect 2543 -1576 2544 -1534
rect 121 -1699 122 -1577
rect 912 -1578 913 -1534
rect 964 -1578 965 -1534
rect 1402 -1699 1403 -1577
rect 1423 -1578 1424 -1534
rect 1801 -1578 1802 -1534
rect 1829 -1699 1830 -1577
rect 1962 -1578 1963 -1534
rect 2067 -1699 2068 -1577
rect 2158 -1578 2159 -1534
rect 2361 -1699 2362 -1577
rect 2487 -1578 2488 -1534
rect 128 -1580 129 -1534
rect 131 -1662 132 -1579
rect 163 -1580 164 -1534
rect 163 -1699 164 -1579
rect 163 -1580 164 -1534
rect 163 -1699 164 -1579
rect 198 -1580 199 -1534
rect 2494 -1580 2495 -1534
rect 128 -1699 129 -1581
rect 674 -1582 675 -1534
rect 849 -1699 850 -1581
rect 919 -1582 920 -1534
rect 989 -1699 990 -1581
rect 1122 -1582 1123 -1534
rect 1143 -1699 1144 -1581
rect 1178 -1582 1179 -1534
rect 1192 -1699 1193 -1581
rect 1325 -1582 1326 -1534
rect 1353 -1699 1354 -1581
rect 1549 -1582 1550 -1534
rect 1605 -1699 1606 -1581
rect 1633 -1582 1634 -1534
rect 1766 -1582 1767 -1534
rect 1941 -1699 1942 -1581
rect 1962 -1699 1963 -1581
rect 2074 -1582 2075 -1534
rect 2081 -1699 2082 -1581
rect 2193 -1582 2194 -1534
rect 2494 -1699 2495 -1581
rect 2522 -1582 2523 -1534
rect 184 -1584 185 -1534
rect 198 -1699 199 -1583
rect 212 -1699 213 -1583
rect 576 -1584 577 -1534
rect 593 -1584 594 -1534
rect 2144 -1699 2145 -1583
rect 2193 -1699 2194 -1583
rect 2298 -1584 2299 -1534
rect 177 -1586 178 -1534
rect 184 -1699 185 -1585
rect 219 -1586 220 -1534
rect 961 -1699 962 -1585
rect 1122 -1699 1123 -1585
rect 1811 -1699 1812 -1585
rect 2074 -1699 2075 -1585
rect 2165 -1586 2166 -1534
rect 2298 -1699 2299 -1585
rect 2424 -1586 2425 -1534
rect 135 -1588 136 -1534
rect 219 -1699 220 -1587
rect 226 -1699 227 -1587
rect 1010 -1699 1011 -1587
rect 1153 -1588 1154 -1534
rect 1269 -1699 1270 -1587
rect 1286 -1588 1287 -1534
rect 1801 -1699 1802 -1587
rect 2165 -1699 2166 -1587
rect 2270 -1588 2271 -1534
rect 135 -1699 136 -1589
rect 1052 -1590 1053 -1534
rect 1157 -1590 1158 -1534
rect 2221 -1590 2222 -1534
rect 2270 -1699 2271 -1589
rect 2312 -1590 2313 -1534
rect 233 -1699 234 -1591
rect 695 -1592 696 -1534
rect 800 -1592 801 -1534
rect 2424 -1699 2425 -1591
rect 236 -1594 237 -1534
rect 478 -1594 479 -1534
rect 506 -1699 507 -1593
rect 541 -1594 542 -1534
rect 667 -1594 668 -1534
rect 800 -1699 801 -1593
rect 870 -1699 871 -1593
rect 1045 -1594 1046 -1534
rect 1157 -1699 1158 -1593
rect 1374 -1594 1375 -1534
rect 1423 -1699 1424 -1593
rect 1619 -1594 1620 -1534
rect 1633 -1699 1634 -1593
rect 1738 -1594 1739 -1534
rect 1766 -1699 1767 -1593
rect 1920 -1594 1921 -1534
rect 2221 -1699 2222 -1593
rect 2277 -1594 2278 -1534
rect 2312 -1699 2313 -1593
rect 2382 -1594 2383 -1534
rect 240 -1596 241 -1534
rect 1017 -1596 1018 -1534
rect 1045 -1699 1046 -1595
rect 1108 -1596 1109 -1534
rect 1160 -1596 1161 -1534
rect 1290 -1596 1291 -1534
rect 1304 -1699 1305 -1595
rect 1437 -1596 1438 -1534
rect 1458 -1699 1459 -1595
rect 1773 -1596 1774 -1534
rect 2277 -1699 2278 -1595
rect 2396 -1596 2397 -1534
rect 156 -1598 157 -1534
rect 240 -1699 241 -1597
rect 247 -1598 248 -1534
rect 408 -1699 409 -1597
rect 415 -1598 416 -1534
rect 737 -1699 738 -1597
rect 828 -1699 829 -1597
rect 1108 -1699 1109 -1597
rect 1171 -1699 1172 -1597
rect 1416 -1598 1417 -1534
rect 1486 -1699 1487 -1597
rect 1563 -1598 1564 -1534
rect 1612 -1699 1613 -1597
rect 1794 -1598 1795 -1534
rect 2382 -1699 2383 -1597
rect 2508 -1598 2509 -1534
rect 156 -1699 157 -1599
rect 170 -1600 171 -1534
rect 275 -1600 276 -1534
rect 453 -1699 454 -1599
rect 464 -1600 465 -1534
rect 534 -1699 535 -1599
rect 667 -1699 668 -1599
rect 933 -1600 934 -1534
rect 954 -1600 955 -1534
rect 1290 -1699 1291 -1599
rect 1325 -1699 1326 -1599
rect 1444 -1600 1445 -1534
rect 1489 -1600 1490 -1534
rect 2235 -1600 2236 -1534
rect 2396 -1699 2397 -1599
rect 2480 -1600 2481 -1534
rect 117 -1602 118 -1534
rect 464 -1699 465 -1601
rect 478 -1699 479 -1601
rect 492 -1602 493 -1534
rect 516 -1602 517 -1534
rect 1052 -1699 1053 -1601
rect 1178 -1699 1179 -1601
rect 1213 -1602 1214 -1534
rect 1265 -1699 1266 -1601
rect 1773 -1699 1774 -1601
rect 1794 -1699 1795 -1601
rect 1892 -1602 1893 -1534
rect 2235 -1699 2236 -1601
rect 2354 -1602 2355 -1534
rect 149 -1604 150 -1534
rect 492 -1699 493 -1603
rect 674 -1699 675 -1603
rect 891 -1604 892 -1534
rect 905 -1604 906 -1534
rect 1451 -1604 1452 -1534
rect 1493 -1699 1494 -1603
rect 1619 -1699 1620 -1603
rect 1738 -1699 1739 -1603
rect 1787 -1604 1788 -1534
rect 1892 -1699 1893 -1603
rect 1997 -1604 1998 -1534
rect 2207 -1604 2208 -1534
rect 2354 -1699 2355 -1603
rect 86 -1606 87 -1534
rect 149 -1699 150 -1605
rect 170 -1699 171 -1605
rect 254 -1606 255 -1534
rect 275 -1699 276 -1605
rect 296 -1606 297 -1534
rect 303 -1699 304 -1605
rect 401 -1606 402 -1534
rect 429 -1699 430 -1605
rect 443 -1606 444 -1534
rect 695 -1699 696 -1605
rect 772 -1606 773 -1534
rect 891 -1699 892 -1605
rect 975 -1606 976 -1534
rect 982 -1606 983 -1534
rect 1017 -1699 1018 -1605
rect 1213 -1699 1214 -1605
rect 1752 -1606 1753 -1534
rect 1759 -1606 1760 -1534
rect 1920 -1699 1921 -1605
rect 1983 -1606 1984 -1534
rect 2207 -1699 2208 -1605
rect 86 -1699 87 -1607
rect 142 -1608 143 -1534
rect 250 -1699 251 -1607
rect 1451 -1699 1452 -1607
rect 1503 -1608 1504 -1534
rect 2466 -1608 2467 -1534
rect 142 -1699 143 -1609
rect 642 -1699 643 -1609
rect 772 -1699 773 -1609
rect 842 -1610 843 -1534
rect 905 -1699 906 -1609
rect 1381 -1610 1382 -1534
rect 1416 -1699 1417 -1609
rect 1465 -1610 1466 -1534
rect 1507 -1610 1508 -1534
rect 1640 -1699 1641 -1609
rect 1752 -1699 1753 -1609
rect 1871 -1610 1872 -1534
rect 1997 -1699 1998 -1609
rect 2102 -1610 2103 -1534
rect 110 -1612 111 -1534
rect 1465 -1699 1466 -1611
rect 1514 -1699 1515 -1611
rect 1682 -1612 1683 -1534
rect 1759 -1699 1760 -1611
rect 1899 -1612 1900 -1534
rect 2102 -1699 2103 -1611
rect 2319 -1612 2320 -1534
rect 205 -1614 206 -1534
rect 1381 -1699 1382 -1613
rect 1444 -1699 1445 -1613
rect 1598 -1614 1599 -1534
rect 1787 -1699 1788 -1613
rect 2109 -1614 2110 -1534
rect 2319 -1699 2320 -1613
rect 2529 -1614 2530 -1534
rect 205 -1699 206 -1615
rect 653 -1616 654 -1534
rect 842 -1699 843 -1615
rect 926 -1616 927 -1534
rect 933 -1699 934 -1615
rect 1115 -1616 1116 -1534
rect 1234 -1699 1235 -1615
rect 1507 -1699 1508 -1615
rect 1531 -1699 1532 -1615
rect 2158 -1699 2159 -1615
rect 254 -1699 255 -1617
rect 1153 -1699 1154 -1617
rect 1276 -1618 1277 -1534
rect 1437 -1699 1438 -1617
rect 1549 -1699 1550 -1617
rect 1668 -1618 1669 -1534
rect 1815 -1618 1816 -1534
rect 1983 -1699 1984 -1617
rect 282 -1699 283 -1619
rect 373 -1620 374 -1534
rect 380 -1620 381 -1534
rect 380 -1699 381 -1619
rect 380 -1620 381 -1534
rect 380 -1699 381 -1619
rect 387 -1620 388 -1534
rect 807 -1699 808 -1619
rect 912 -1699 913 -1619
rect 1570 -1620 1571 -1534
rect 1668 -1699 1669 -1619
rect 1780 -1620 1781 -1534
rect 1871 -1699 1872 -1619
rect 1948 -1620 1949 -1534
rect 96 -1699 97 -1621
rect 1570 -1699 1571 -1621
rect 1899 -1699 1900 -1621
rect 2011 -1622 2012 -1534
rect 296 -1699 297 -1623
rect 611 -1624 612 -1534
rect 919 -1699 920 -1623
rect 1031 -1624 1032 -1534
rect 1034 -1699 1035 -1623
rect 1598 -1699 1599 -1623
rect 1927 -1624 1928 -1534
rect 2109 -1699 2110 -1623
rect 338 -1626 339 -1534
rect 401 -1699 402 -1625
rect 436 -1626 437 -1534
rect 940 -1699 941 -1625
rect 954 -1699 955 -1625
rect 1059 -1626 1060 -1534
rect 1115 -1699 1116 -1625
rect 1136 -1626 1137 -1534
rect 1258 -1626 1259 -1534
rect 1815 -1699 1816 -1625
rect 1927 -1699 1928 -1625
rect 2025 -1626 2026 -1534
rect 338 -1699 339 -1627
rect 345 -1628 346 -1534
rect 352 -1628 353 -1534
rect 415 -1699 416 -1627
rect 436 -1699 437 -1627
rect 1500 -1628 1501 -1534
rect 1563 -1699 1564 -1627
rect 1696 -1628 1697 -1534
rect 1948 -1699 1949 -1627
rect 2046 -1628 2047 -1534
rect 289 -1630 290 -1534
rect 352 -1699 353 -1629
rect 373 -1699 374 -1629
rect 457 -1630 458 -1534
rect 562 -1630 563 -1534
rect 611 -1699 612 -1629
rect 926 -1699 927 -1629
rect 1073 -1630 1074 -1534
rect 1136 -1699 1137 -1629
rect 1318 -1630 1319 -1534
rect 1349 -1630 1350 -1534
rect 1682 -1699 1683 -1629
rect 1689 -1630 1690 -1534
rect 1696 -1699 1697 -1629
rect 2004 -1630 2005 -1534
rect 2011 -1699 2012 -1629
rect 2025 -1699 2026 -1629
rect 2130 -1630 2131 -1534
rect 191 -1632 192 -1534
rect 289 -1699 290 -1631
rect 317 -1632 318 -1534
rect 345 -1699 346 -1631
rect 387 -1699 388 -1631
rect 1003 -1632 1004 -1534
rect 1059 -1699 1060 -1631
rect 1101 -1632 1102 -1534
rect 1262 -1632 1263 -1534
rect 1780 -1699 1781 -1631
rect 2004 -1699 2005 -1631
rect 2116 -1632 2117 -1534
rect 2130 -1699 2131 -1631
rect 2249 -1632 2250 -1534
rect 191 -1699 192 -1633
rect 618 -1699 619 -1633
rect 975 -1699 976 -1633
rect 1080 -1634 1081 -1534
rect 1101 -1699 1102 -1633
rect 1227 -1634 1228 -1534
rect 1276 -1699 1277 -1633
rect 1521 -1699 1522 -1633
rect 1689 -1699 1690 -1633
rect 1808 -1634 1809 -1534
rect 2046 -1699 2047 -1633
rect 2137 -1634 2138 -1534
rect 2249 -1699 2250 -1633
rect 2459 -1634 2460 -1534
rect 194 -1699 195 -1635
rect 1262 -1699 1263 -1635
rect 1318 -1699 1319 -1635
rect 1654 -1636 1655 -1534
rect 1808 -1699 1809 -1635
rect 2179 -1636 2180 -1534
rect 317 -1699 318 -1637
rect 359 -1638 360 -1534
rect 394 -1638 395 -1534
rect 639 -1638 640 -1534
rect 968 -1638 969 -1534
rect 1227 -1699 1228 -1637
rect 1293 -1699 1294 -1637
rect 1654 -1699 1655 -1637
rect 2116 -1699 2117 -1637
rect 2228 -1638 2229 -1534
rect 324 -1640 325 -1534
rect 457 -1699 458 -1639
rect 548 -1640 549 -1534
rect 562 -1699 563 -1639
rect 639 -1699 640 -1639
rect 2550 -1640 2551 -1534
rect 324 -1699 325 -1641
rect 555 -1642 556 -1534
rect 856 -1642 857 -1534
rect 968 -1699 969 -1641
rect 982 -1699 983 -1641
rect 1164 -1642 1165 -1534
rect 1374 -1699 1375 -1641
rect 1535 -1642 1536 -1534
rect 2137 -1699 2138 -1641
rect 2375 -1642 2376 -1534
rect 331 -1644 332 -1534
rect 359 -1699 360 -1643
rect 394 -1699 395 -1643
rect 632 -1644 633 -1534
rect 653 -1699 654 -1643
rect 856 -1699 857 -1643
rect 1003 -1699 1004 -1643
rect 1185 -1644 1186 -1534
rect 1500 -1699 1501 -1643
rect 1626 -1644 1627 -1534
rect 2200 -1644 2201 -1534
rect 2375 -1699 2376 -1643
rect 331 -1699 332 -1645
rect 485 -1646 486 -1534
rect 548 -1699 549 -1645
rect 758 -1646 759 -1534
rect 1073 -1699 1074 -1645
rect 2186 -1646 2187 -1534
rect 2200 -1699 2201 -1645
rect 2263 -1646 2264 -1534
rect 180 -1699 181 -1647
rect 2186 -1699 2187 -1647
rect 2228 -1699 2229 -1647
rect 2333 -1648 2334 -1534
rect 443 -1699 444 -1649
rect 1346 -1650 1347 -1534
rect 1468 -1699 1469 -1649
rect 2263 -1699 2264 -1649
rect 2333 -1699 2334 -1649
rect 2452 -1650 2453 -1534
rect 450 -1652 451 -1534
rect 632 -1699 633 -1651
rect 758 -1699 759 -1651
rect 835 -1652 836 -1534
rect 996 -1652 997 -1534
rect 1346 -1699 1347 -1651
rect 1430 -1652 1431 -1534
rect 2452 -1699 2453 -1651
rect 450 -1699 451 -1653
rect 730 -1699 731 -1653
rect 765 -1654 766 -1534
rect 835 -1699 836 -1653
rect 1080 -1699 1081 -1653
rect 1199 -1654 1200 -1534
rect 1430 -1699 1431 -1653
rect 1556 -1654 1557 -1534
rect 1626 -1699 1627 -1653
rect 1731 -1654 1732 -1534
rect 485 -1699 486 -1655
rect 716 -1656 717 -1534
rect 765 -1699 766 -1655
rect 1087 -1656 1088 -1534
rect 1164 -1699 1165 -1655
rect 1367 -1656 1368 -1534
rect 1528 -1656 1529 -1534
rect 2179 -1699 2180 -1655
rect 513 -1658 514 -1534
rect 996 -1699 997 -1657
rect 1087 -1699 1088 -1657
rect 1363 -1699 1364 -1657
rect 1367 -1699 1368 -1657
rect 1472 -1658 1473 -1534
rect 1535 -1699 1536 -1657
rect 2060 -1699 2061 -1657
rect 513 -1699 514 -1659
rect 688 -1660 689 -1534
rect 786 -1660 787 -1534
rect 1199 -1699 1200 -1659
rect 1388 -1660 1389 -1534
rect 1528 -1699 1529 -1659
rect 1556 -1699 1557 -1659
rect 1724 -1660 1725 -1534
rect 786 -1699 787 -1661
rect 866 -1662 867 -1534
rect 1731 -1699 1732 -1661
rect 555 -1699 556 -1663
rect 2441 -1699 2442 -1663
rect 569 -1666 570 -1534
rect 716 -1699 717 -1665
rect 1185 -1699 1186 -1665
rect 1241 -1666 1242 -1534
rect 1388 -1699 1389 -1665
rect 1542 -1666 1543 -1534
rect 1724 -1699 1725 -1665
rect 1850 -1666 1851 -1534
rect 569 -1699 570 -1667
rect 863 -1668 864 -1534
rect 1241 -1699 1242 -1667
rect 1339 -1668 1340 -1534
rect 1472 -1699 1473 -1667
rect 1661 -1668 1662 -1534
rect 1850 -1699 1851 -1667
rect 1934 -1668 1935 -1534
rect 688 -1699 689 -1669
rect 744 -1670 745 -1534
rect 863 -1699 864 -1669
rect 947 -1670 948 -1534
rect 1339 -1699 1340 -1669
rect 1409 -1670 1410 -1534
rect 1542 -1699 1543 -1669
rect 1647 -1670 1648 -1534
rect 1661 -1699 1662 -1669
rect 1745 -1670 1746 -1534
rect 1934 -1699 1935 -1669
rect 2039 -1670 2040 -1534
rect 9 -1672 10 -1534
rect 744 -1699 745 -1671
rect 947 -1699 948 -1671
rect 2557 -1672 2558 -1534
rect 93 -1699 94 -1673
rect 2039 -1699 2040 -1673
rect 1409 -1699 1410 -1675
rect 1591 -1676 1592 -1534
rect 1745 -1699 1746 -1675
rect 1857 -1676 1858 -1534
rect 1510 -1699 1511 -1677
rect 1857 -1699 1858 -1677
rect 1577 -1680 1578 -1534
rect 1647 -1699 1648 -1679
rect 1577 -1699 1578 -1681
rect 1703 -1682 1704 -1534
rect 1591 -1699 1592 -1683
rect 1717 -1684 1718 -1534
rect 1703 -1699 1704 -1685
rect 2410 -1699 2411 -1685
rect 1717 -1699 1718 -1687
rect 1843 -1688 1844 -1534
rect 1843 -1699 1844 -1689
rect 1913 -1690 1914 -1534
rect 1913 -1699 1914 -1691
rect 2151 -1692 2152 -1534
rect 2151 -1699 2152 -1693
rect 2256 -1694 2257 -1534
rect 2256 -1699 2257 -1695
rect 2368 -1696 2369 -1534
rect 2368 -1699 2369 -1697
rect 2501 -1698 2502 -1534
rect 2 -1850 3 -1708
rect 387 -1709 388 -1707
rect 422 -1709 423 -1707
rect 422 -1850 423 -1708
rect 422 -1709 423 -1707
rect 422 -1850 423 -1708
rect 429 -1709 430 -1707
rect 1538 -1709 1539 -1707
rect 1549 -1709 1550 -1707
rect 1549 -1850 1550 -1708
rect 1549 -1709 1550 -1707
rect 1549 -1850 1550 -1708
rect 1629 -1850 1630 -1708
rect 2046 -1709 2047 -1707
rect 2389 -1709 2390 -1707
rect 2438 -1850 2439 -1708
rect 2445 -1709 2446 -1707
rect 2459 -1850 2460 -1708
rect 2469 -1850 2470 -1708
rect 2494 -1709 2495 -1707
rect 9 -1850 10 -1710
rect 107 -1711 108 -1707
rect 142 -1711 143 -1707
rect 145 -1769 146 -1710
rect 163 -1711 164 -1707
rect 163 -1850 164 -1710
rect 163 -1711 164 -1707
rect 163 -1850 164 -1710
rect 187 -1850 188 -1710
rect 1265 -1711 1266 -1707
rect 1276 -1711 1277 -1707
rect 2410 -1711 2411 -1707
rect 16 -1713 17 -1707
rect 614 -1850 615 -1712
rect 649 -1850 650 -1712
rect 943 -1850 944 -1712
rect 1017 -1713 1018 -1707
rect 1605 -1713 1606 -1707
rect 1640 -1713 1641 -1707
rect 1640 -1850 1641 -1712
rect 1640 -1713 1641 -1707
rect 1640 -1850 1641 -1712
rect 1664 -1850 1665 -1712
rect 2312 -1713 2313 -1707
rect 2347 -1713 2348 -1707
rect 2410 -1850 2411 -1712
rect 16 -1850 17 -1714
rect 1003 -1715 1004 -1707
rect 1020 -1715 1021 -1707
rect 1192 -1715 1193 -1707
rect 1206 -1715 1207 -1707
rect 1290 -1715 1291 -1707
rect 1293 -1715 1294 -1707
rect 2270 -1715 2271 -1707
rect 2389 -1850 2390 -1714
rect 2473 -1850 2474 -1714
rect 23 -1717 24 -1707
rect 23 -1850 24 -1716
rect 23 -1717 24 -1707
rect 23 -1850 24 -1716
rect 30 -1717 31 -1707
rect 894 -1850 895 -1716
rect 919 -1717 920 -1707
rect 919 -1850 920 -1716
rect 919 -1717 920 -1707
rect 919 -1850 920 -1716
rect 989 -1717 990 -1707
rect 1017 -1850 1018 -1716
rect 1031 -1717 1032 -1707
rect 1402 -1717 1403 -1707
rect 1437 -1717 1438 -1707
rect 1738 -1717 1739 -1707
rect 1801 -1717 1802 -1707
rect 2476 -1850 2477 -1716
rect 30 -1850 31 -1718
rect 331 -1719 332 -1707
rect 446 -1850 447 -1718
rect 807 -1719 808 -1707
rect 821 -1719 822 -1707
rect 1073 -1719 1074 -1707
rect 1108 -1719 1109 -1707
rect 2417 -1719 2418 -1707
rect 37 -1721 38 -1707
rect 96 -1721 97 -1707
rect 107 -1850 108 -1720
rect 373 -1721 374 -1707
rect 394 -1721 395 -1707
rect 807 -1850 808 -1720
rect 821 -1850 822 -1720
rect 1363 -1721 1364 -1707
rect 1367 -1721 1368 -1707
rect 1402 -1850 1403 -1720
rect 1440 -1721 1441 -1707
rect 2291 -1721 2292 -1707
rect 2361 -1721 2362 -1707
rect 2417 -1850 2418 -1720
rect 37 -1850 38 -1722
rect 443 -1723 444 -1707
rect 457 -1850 458 -1722
rect 828 -1723 829 -1707
rect 835 -1723 836 -1707
rect 908 -1850 909 -1722
rect 961 -1723 962 -1707
rect 1031 -1850 1032 -1722
rect 1059 -1723 1060 -1707
rect 1062 -1769 1063 -1722
rect 1111 -1723 1112 -1707
rect 1885 -1723 1886 -1707
rect 1997 -1723 1998 -1707
rect 2046 -1850 2047 -1722
rect 2228 -1723 2229 -1707
rect 2291 -1850 2292 -1722
rect 2305 -1723 2306 -1707
rect 2361 -1850 2362 -1722
rect 47 -1850 48 -1724
rect 51 -1725 52 -1707
rect 65 -1725 66 -1707
rect 180 -1725 181 -1707
rect 194 -1725 195 -1707
rect 1101 -1725 1102 -1707
rect 1129 -1725 1130 -1707
rect 1129 -1850 1130 -1724
rect 1129 -1725 1130 -1707
rect 1129 -1850 1130 -1724
rect 1153 -1725 1154 -1707
rect 1696 -1725 1697 -1707
rect 1706 -1725 1707 -1707
rect 2375 -1725 2376 -1707
rect 51 -1850 52 -1726
rect 240 -1727 241 -1707
rect 247 -1727 248 -1707
rect 534 -1727 535 -1707
rect 548 -1727 549 -1707
rect 856 -1727 857 -1707
rect 870 -1727 871 -1707
rect 961 -1850 962 -1726
rect 989 -1850 990 -1726
rect 1010 -1727 1011 -1707
rect 1059 -1850 1060 -1726
rect 1409 -1727 1410 -1707
rect 1440 -1850 1441 -1726
rect 1703 -1850 1704 -1726
rect 1836 -1727 1837 -1707
rect 2434 -1727 2435 -1707
rect 58 -1729 59 -1707
rect 65 -1850 66 -1728
rect 86 -1729 87 -1707
rect 159 -1850 160 -1728
rect 198 -1729 199 -1707
rect 1150 -1729 1151 -1707
rect 1192 -1850 1193 -1728
rect 1283 -1729 1284 -1707
rect 1293 -1850 1294 -1728
rect 1444 -1729 1445 -1707
rect 1458 -1729 1459 -1707
rect 1997 -1850 1998 -1728
rect 2039 -1729 2040 -1707
rect 2042 -1729 2043 -1707
rect 2228 -1850 2229 -1728
rect 2319 -1729 2320 -1707
rect 58 -1850 59 -1730
rect 898 -1731 899 -1707
rect 957 -1850 958 -1730
rect 1444 -1850 1445 -1730
rect 1468 -1731 1469 -1707
rect 2396 -1731 2397 -1707
rect 86 -1850 87 -1732
rect 135 -1733 136 -1707
rect 142 -1850 143 -1732
rect 460 -1733 461 -1707
rect 632 -1733 633 -1707
rect 653 -1733 654 -1707
rect 828 -1850 829 -1732
rect 870 -1850 871 -1732
rect 891 -1733 892 -1707
rect 1003 -1850 1004 -1732
rect 1094 -1733 1095 -1707
rect 1143 -1733 1144 -1707
rect 1150 -1850 1151 -1732
rect 1209 -1850 1210 -1732
rect 1374 -1733 1375 -1707
rect 1388 -1733 1389 -1707
rect 1458 -1850 1459 -1732
rect 1468 -1850 1469 -1732
rect 2319 -1850 2320 -1732
rect 44 -1735 45 -1707
rect 1374 -1850 1375 -1734
rect 1493 -1735 1494 -1707
rect 1647 -1735 1648 -1707
rect 1696 -1850 1697 -1734
rect 1941 -1735 1942 -1707
rect 2039 -1850 2040 -1734
rect 2137 -1735 2138 -1707
rect 2235 -1735 2236 -1707
rect 2305 -1850 2306 -1734
rect 93 -1737 94 -1707
rect 926 -1737 927 -1707
rect 1143 -1850 1144 -1736
rect 1181 -1850 1182 -1736
rect 1213 -1737 1214 -1707
rect 1307 -1850 1308 -1736
rect 1325 -1737 1326 -1707
rect 1367 -1850 1368 -1736
rect 1493 -1850 1494 -1736
rect 1591 -1737 1592 -1707
rect 1647 -1850 1648 -1736
rect 1808 -1737 1809 -1707
rect 1815 -1737 1816 -1707
rect 1836 -1850 1837 -1736
rect 1850 -1737 1851 -1707
rect 1885 -1850 1886 -1736
rect 1941 -1850 1942 -1736
rect 2158 -1737 2159 -1707
rect 2179 -1737 2180 -1707
rect 2235 -1850 2236 -1736
rect 2242 -1737 2243 -1707
rect 2270 -1850 2271 -1736
rect 2284 -1737 2285 -1707
rect 2375 -1850 2376 -1736
rect 93 -1850 94 -1738
rect 380 -1739 381 -1707
rect 429 -1850 430 -1738
rect 926 -1850 927 -1738
rect 1171 -1739 1172 -1707
rect 1325 -1850 1326 -1738
rect 1360 -1739 1361 -1707
rect 2207 -1739 2208 -1707
rect 2221 -1739 2222 -1707
rect 2284 -1850 2285 -1738
rect 135 -1850 136 -1740
rect 205 -1741 206 -1707
rect 212 -1741 213 -1707
rect 863 -1741 864 -1707
rect 884 -1741 885 -1707
rect 1073 -1850 1074 -1740
rect 1164 -1741 1165 -1707
rect 1171 -1850 1172 -1740
rect 1213 -1850 1214 -1740
rect 1241 -1741 1242 -1707
rect 1255 -1741 1256 -1707
rect 1255 -1850 1256 -1740
rect 1255 -1741 1256 -1707
rect 1255 -1850 1256 -1740
rect 1262 -1741 1263 -1707
rect 2018 -1741 2019 -1707
rect 2081 -1741 2082 -1707
rect 2137 -1850 2138 -1740
rect 2151 -1741 2152 -1707
rect 2221 -1850 2222 -1740
rect 2263 -1741 2264 -1707
rect 2347 -1850 2348 -1740
rect 100 -1743 101 -1707
rect 205 -1850 206 -1742
rect 212 -1850 213 -1742
rect 758 -1743 759 -1707
rect 765 -1743 766 -1707
rect 765 -1850 766 -1742
rect 765 -1743 766 -1707
rect 765 -1850 766 -1742
rect 793 -1743 794 -1707
rect 1010 -1850 1011 -1742
rect 1220 -1743 1221 -1707
rect 1220 -1850 1221 -1742
rect 1220 -1743 1221 -1707
rect 1220 -1850 1221 -1742
rect 1227 -1743 1228 -1707
rect 1388 -1850 1389 -1742
rect 1500 -1743 1501 -1707
rect 1500 -1850 1501 -1742
rect 1500 -1743 1501 -1707
rect 1500 -1850 1501 -1742
rect 1510 -1743 1511 -1707
rect 2200 -1743 2201 -1707
rect 198 -1850 199 -1744
rect 366 -1745 367 -1707
rect 373 -1850 374 -1744
rect 565 -1850 566 -1744
rect 579 -1745 580 -1707
rect 1738 -1850 1739 -1744
rect 1745 -1745 1746 -1707
rect 2242 -1850 2243 -1744
rect 226 -1850 227 -1746
rect 912 -1747 913 -1707
rect 940 -1747 941 -1707
rect 1164 -1850 1165 -1746
rect 1185 -1747 1186 -1707
rect 1227 -1850 1228 -1746
rect 1241 -1850 1242 -1746
rect 1311 -1747 1312 -1707
rect 1353 -1747 1354 -1707
rect 1360 -1850 1361 -1746
rect 1528 -1747 1529 -1707
rect 2403 -1747 2404 -1707
rect 229 -1749 230 -1707
rect 1094 -1850 1095 -1748
rect 1248 -1749 1249 -1707
rect 1262 -1850 1263 -1748
rect 1283 -1850 1284 -1748
rect 1521 -1749 1522 -1707
rect 1528 -1850 1529 -1748
rect 1542 -1749 1543 -1707
rect 1556 -1749 1557 -1707
rect 1605 -1850 1606 -1748
rect 1724 -1749 1725 -1707
rect 1745 -1850 1746 -1748
rect 1759 -1749 1760 -1707
rect 2018 -1850 2019 -1748
rect 2102 -1749 2103 -1707
rect 2263 -1850 2264 -1748
rect 2333 -1749 2334 -1707
rect 2403 -1850 2404 -1748
rect 124 -1850 125 -1750
rect 1521 -1850 1522 -1750
rect 1531 -1751 1532 -1707
rect 2312 -1850 2313 -1750
rect 236 -1850 237 -1752
rect 954 -1753 955 -1707
rect 1052 -1753 1053 -1707
rect 1185 -1850 1186 -1752
rect 1297 -1753 1298 -1707
rect 1409 -1850 1410 -1752
rect 1535 -1753 1536 -1707
rect 2088 -1753 2089 -1707
rect 2130 -1753 2131 -1707
rect 2207 -1850 2208 -1752
rect 240 -1850 241 -1754
rect 1076 -1755 1077 -1707
rect 1234 -1755 1235 -1707
rect 1297 -1850 1298 -1754
rect 1304 -1755 1305 -1707
rect 1353 -1850 1354 -1754
rect 1535 -1850 1536 -1754
rect 1612 -1755 1613 -1707
rect 1619 -1755 1620 -1707
rect 1759 -1850 1760 -1754
rect 1773 -1755 1774 -1707
rect 1815 -1850 1816 -1754
rect 1850 -1850 1851 -1754
rect 2354 -1755 2355 -1707
rect 254 -1757 255 -1707
rect 254 -1850 255 -1756
rect 254 -1757 255 -1707
rect 254 -1850 255 -1756
rect 289 -1757 290 -1707
rect 698 -1757 699 -1707
rect 702 -1757 703 -1707
rect 702 -1850 703 -1756
rect 702 -1757 703 -1707
rect 702 -1850 703 -1756
rect 716 -1757 717 -1707
rect 2158 -1850 2159 -1756
rect 2165 -1757 2166 -1707
rect 2200 -1850 2201 -1756
rect 2298 -1757 2299 -1707
rect 2354 -1850 2355 -1756
rect 289 -1850 290 -1758
rect 324 -1759 325 -1707
rect 331 -1850 332 -1758
rect 513 -1759 514 -1707
rect 520 -1759 521 -1707
rect 639 -1850 640 -1758
rect 653 -1850 654 -1758
rect 737 -1759 738 -1707
rect 744 -1759 745 -1707
rect 1052 -1850 1053 -1758
rect 1157 -1759 1158 -1707
rect 1234 -1850 1235 -1758
rect 1290 -1850 1291 -1758
rect 2165 -1850 2166 -1758
rect 2179 -1850 2180 -1758
rect 2382 -1759 2383 -1707
rect 303 -1761 304 -1707
rect 303 -1850 304 -1760
rect 303 -1761 304 -1707
rect 303 -1850 304 -1760
rect 324 -1850 325 -1760
rect 590 -1761 591 -1707
rect 618 -1761 619 -1707
rect 1108 -1850 1109 -1760
rect 1115 -1761 1116 -1707
rect 1157 -1850 1158 -1760
rect 1304 -1850 1305 -1760
rect 1801 -1850 1802 -1760
rect 1808 -1850 1809 -1760
rect 1913 -1761 1914 -1707
rect 2053 -1761 2054 -1707
rect 2102 -1850 2103 -1760
rect 2151 -1850 2152 -1760
rect 2424 -1761 2425 -1707
rect 121 -1763 122 -1707
rect 618 -1850 619 -1762
rect 660 -1763 661 -1707
rect 737 -1850 738 -1762
rect 744 -1850 745 -1762
rect 905 -1763 906 -1707
rect 912 -1850 913 -1762
rect 1045 -1763 1046 -1707
rect 1496 -1763 1497 -1707
rect 2298 -1850 2299 -1762
rect 2340 -1763 2341 -1707
rect 2382 -1850 2383 -1762
rect 79 -1765 80 -1707
rect 121 -1850 122 -1764
rect 345 -1765 346 -1707
rect 366 -1850 367 -1764
rect 387 -1850 388 -1764
rect 513 -1850 514 -1764
rect 520 -1850 521 -1764
rect 611 -1765 612 -1707
rect 667 -1765 668 -1707
rect 835 -1850 836 -1764
rect 849 -1765 850 -1707
rect 884 -1850 885 -1764
rect 891 -1850 892 -1764
rect 1983 -1765 1984 -1707
rect 2004 -1765 2005 -1707
rect 2340 -1850 2341 -1764
rect 79 -1850 80 -1766
rect 268 -1767 269 -1707
rect 275 -1767 276 -1707
rect 345 -1850 346 -1766
rect 352 -1767 353 -1707
rect 380 -1850 381 -1766
rect 436 -1767 437 -1707
rect 534 -1850 535 -1766
rect 548 -1850 549 -1766
rect 947 -1767 948 -1707
rect 954 -1850 955 -1766
rect 1279 -1767 1280 -1707
rect 1556 -1850 1557 -1766
rect 1626 -1767 1627 -1707
rect 1724 -1850 1725 -1766
rect 1871 -1767 1872 -1707
rect 1934 -1767 1935 -1707
rect 1983 -1850 1984 -1766
rect 2025 -1767 2026 -1707
rect 2053 -1850 2054 -1766
rect 2249 -1767 2250 -1707
rect 2424 -1850 2425 -1766
rect 149 -1769 150 -1707
rect 436 -1850 437 -1768
rect 443 -1850 444 -1768
rect 1542 -1850 1543 -1768
rect 1563 -1769 1564 -1707
rect 1591 -1850 1592 -1768
rect 1598 -1769 1599 -1707
rect 1612 -1850 1613 -1768
rect 1619 -1850 1620 -1768
rect 1717 -1769 1718 -1707
rect 1773 -1850 1774 -1768
rect 1899 -1769 1900 -1707
rect 1955 -1769 1956 -1707
rect 2004 -1850 2005 -1768
rect 2042 -1850 2043 -1768
rect 2081 -1850 2082 -1768
rect 149 -1850 150 -1770
rect 184 -1771 185 -1707
rect 268 -1850 269 -1770
rect 338 -1771 339 -1707
rect 352 -1850 353 -1770
rect 408 -1771 409 -1707
rect 481 -1771 482 -1707
rect 1311 -1850 1312 -1770
rect 1465 -1771 1466 -1707
rect 1934 -1850 1935 -1770
rect 1969 -1771 1970 -1707
rect 2249 -1850 2250 -1770
rect 114 -1773 115 -1707
rect 338 -1850 339 -1772
rect 359 -1773 360 -1707
rect 394 -1850 395 -1772
rect 408 -1850 409 -1772
rect 415 -1773 416 -1707
rect 492 -1773 493 -1707
rect 660 -1850 661 -1772
rect 667 -1850 668 -1772
rect 681 -1773 682 -1707
rect 695 -1773 696 -1707
rect 2445 -1850 2446 -1772
rect 114 -1850 115 -1774
rect 1423 -1775 1424 -1707
rect 1465 -1850 1466 -1774
rect 1731 -1775 1732 -1707
rect 1787 -1775 1788 -1707
rect 2333 -1850 2334 -1774
rect 275 -1850 276 -1776
rect 282 -1777 283 -1707
rect 317 -1777 318 -1707
rect 359 -1850 360 -1776
rect 415 -1850 416 -1776
rect 597 -1777 598 -1707
rect 646 -1777 647 -1707
rect 947 -1850 948 -1776
rect 968 -1777 969 -1707
rect 1913 -1850 1914 -1776
rect 1927 -1777 1928 -1707
rect 1969 -1850 1970 -1776
rect 1976 -1777 1977 -1707
rect 2025 -1850 2026 -1776
rect 282 -1850 283 -1778
rect 569 -1779 570 -1707
rect 590 -1850 591 -1778
rect 688 -1779 689 -1707
rect 695 -1850 696 -1778
rect 730 -1779 731 -1707
rect 733 -1850 734 -1778
rect 996 -1779 997 -1707
rect 1045 -1850 1046 -1778
rect 1066 -1779 1067 -1707
rect 1269 -1779 1270 -1707
rect 1423 -1850 1424 -1778
rect 1479 -1779 1480 -1707
rect 1787 -1850 1788 -1778
rect 1843 -1779 1844 -1707
rect 1871 -1850 1872 -1778
rect 1878 -1779 1879 -1707
rect 1955 -1850 1956 -1778
rect 1976 -1850 1977 -1778
rect 2172 -1779 2173 -1707
rect 219 -1781 220 -1707
rect 1269 -1850 1270 -1780
rect 1276 -1850 1277 -1780
rect 1878 -1850 1879 -1780
rect 2123 -1781 2124 -1707
rect 2172 -1850 2173 -1780
rect 191 -1783 192 -1707
rect 219 -1850 220 -1782
rect 296 -1783 297 -1707
rect 597 -1850 598 -1782
rect 674 -1783 675 -1707
rect 856 -1850 857 -1782
rect 863 -1850 864 -1782
rect 1507 -1783 1508 -1707
rect 1563 -1850 1564 -1782
rect 1794 -1783 1795 -1707
rect 1857 -1783 1858 -1707
rect 1899 -1850 1900 -1782
rect 2074 -1783 2075 -1707
rect 2123 -1850 2124 -1782
rect 191 -1850 192 -1784
rect 485 -1785 486 -1707
rect 492 -1850 493 -1784
rect 506 -1785 507 -1707
rect 516 -1850 517 -1784
rect 1066 -1850 1067 -1784
rect 1472 -1785 1473 -1707
rect 1843 -1850 1844 -1784
rect 2074 -1850 2075 -1784
rect 2326 -1785 2327 -1707
rect 261 -1787 262 -1707
rect 296 -1850 297 -1786
rect 310 -1787 311 -1707
rect 317 -1850 318 -1786
rect 453 -1787 454 -1707
rect 688 -1850 689 -1786
rect 716 -1850 717 -1786
rect 751 -1787 752 -1707
rect 758 -1850 759 -1786
rect 982 -1787 983 -1707
rect 1430 -1787 1431 -1707
rect 1472 -1850 1473 -1786
rect 1479 -1850 1480 -1786
rect 1486 -1787 1487 -1707
rect 1507 -1850 1508 -1786
rect 1990 -1787 1991 -1707
rect 2116 -1787 2117 -1707
rect 2326 -1850 2327 -1786
rect 250 -1850 251 -1788
rect 261 -1850 262 -1788
rect 310 -1850 311 -1788
rect 527 -1789 528 -1707
rect 562 -1789 563 -1707
rect 576 -1789 577 -1707
rect 625 -1789 626 -1707
rect 751 -1850 752 -1788
rect 779 -1789 780 -1707
rect 793 -1850 794 -1788
rect 877 -1789 878 -1707
rect 968 -1850 969 -1788
rect 971 -1789 972 -1707
rect 2130 -1850 2131 -1788
rect 100 -1850 101 -1790
rect 562 -1850 563 -1790
rect 576 -1850 577 -1790
rect 740 -1850 741 -1790
rect 803 -1850 804 -1790
rect 877 -1850 878 -1790
rect 898 -1850 899 -1790
rect 1279 -1850 1280 -1790
rect 1332 -1791 1333 -1707
rect 1486 -1850 1487 -1790
rect 1570 -1791 1571 -1707
rect 1598 -1850 1599 -1790
rect 1675 -1791 1676 -1707
rect 1927 -1850 1928 -1790
rect 1948 -1791 1949 -1707
rect 1990 -1850 1991 -1790
rect 2060 -1791 2061 -1707
rect 2116 -1850 2117 -1790
rect 128 -1793 129 -1707
rect 527 -1850 528 -1792
rect 625 -1850 626 -1792
rect 646 -1850 647 -1792
rect 674 -1850 675 -1792
rect 709 -1793 710 -1707
rect 719 -1793 720 -1707
rect 1248 -1850 1249 -1792
rect 1346 -1793 1347 -1707
rect 1430 -1850 1431 -1792
rect 1451 -1793 1452 -1707
rect 1570 -1850 1571 -1792
rect 1661 -1793 1662 -1707
rect 1675 -1850 1676 -1792
rect 1717 -1850 1718 -1792
rect 1853 -1850 1854 -1792
rect 1920 -1793 1921 -1707
rect 1948 -1850 1949 -1792
rect 2032 -1793 2033 -1707
rect 2060 -1850 2061 -1792
rect 128 -1850 129 -1794
rect 233 -1795 234 -1707
rect 464 -1795 465 -1707
rect 681 -1850 682 -1794
rect 723 -1795 724 -1707
rect 1101 -1850 1102 -1794
rect 1199 -1795 1200 -1707
rect 1332 -1850 1333 -1794
rect 1346 -1850 1347 -1794
rect 1577 -1795 1578 -1707
rect 1752 -1795 1753 -1707
rect 1794 -1850 1795 -1794
rect 1822 -1795 1823 -1707
rect 1857 -1850 1858 -1794
rect 1892 -1795 1893 -1707
rect 1920 -1850 1921 -1794
rect 2032 -1850 2033 -1794
rect 2441 -1795 2442 -1707
rect 177 -1797 178 -1707
rect 709 -1850 710 -1796
rect 730 -1850 731 -1796
rect 1731 -1850 1732 -1796
rect 1892 -1850 1893 -1796
rect 2095 -1797 2096 -1707
rect 170 -1799 171 -1707
rect 177 -1850 178 -1798
rect 201 -1850 202 -1798
rect 779 -1850 780 -1798
rect 905 -1850 906 -1798
rect 2396 -1850 2397 -1798
rect 156 -1801 157 -1707
rect 170 -1850 171 -1800
rect 215 -1801 216 -1707
rect 1752 -1850 1753 -1800
rect 2011 -1801 2012 -1707
rect 2095 -1850 2096 -1800
rect 233 -1850 234 -1802
rect 485 -1850 486 -1802
rect 499 -1803 500 -1707
rect 569 -1850 570 -1802
rect 604 -1803 605 -1707
rect 723 -1850 724 -1802
rect 933 -1803 934 -1707
rect 2088 -1850 2089 -1802
rect 464 -1850 465 -1804
rect 471 -1805 472 -1707
rect 478 -1805 479 -1707
rect 604 -1850 605 -1804
rect 611 -1850 612 -1804
rect 1451 -1850 1452 -1804
rect 1577 -1850 1578 -1804
rect 1584 -1805 1585 -1707
rect 1962 -1805 1963 -1707
rect 2011 -1850 2012 -1804
rect 72 -1807 73 -1707
rect 471 -1850 472 -1806
rect 499 -1850 500 -1806
rect 555 -1807 556 -1707
rect 936 -1807 937 -1707
rect 996 -1850 997 -1806
rect 1024 -1807 1025 -1707
rect 1199 -1850 1200 -1806
rect 1514 -1807 1515 -1707
rect 1584 -1850 1585 -1806
rect 1710 -1807 1711 -1707
rect 1962 -1850 1963 -1806
rect 72 -1850 73 -1808
rect 401 -1809 402 -1707
rect 506 -1850 507 -1808
rect 814 -1809 815 -1707
rect 940 -1850 941 -1808
rect 2186 -1809 2187 -1707
rect 184 -1850 185 -1810
rect 478 -1850 479 -1810
rect 541 -1811 542 -1707
rect 933 -1850 934 -1810
rect 975 -1811 976 -1707
rect 982 -1850 983 -1810
rect 1024 -1850 1025 -1810
rect 1318 -1811 1319 -1707
rect 1381 -1811 1382 -1707
rect 1514 -1850 1515 -1810
rect 1689 -1811 1690 -1707
rect 1710 -1850 1711 -1810
rect 2186 -1850 2187 -1810
rect 2466 -1850 2467 -1810
rect 401 -1850 402 -1812
rect 583 -1813 584 -1707
rect 814 -1850 815 -1812
rect 842 -1813 843 -1707
rect 975 -1850 976 -1812
rect 1038 -1813 1039 -1707
rect 1136 -1813 1137 -1707
rect 1381 -1850 1382 -1812
rect 1437 -1850 1438 -1812
rect 1689 -1850 1690 -1812
rect 541 -1850 542 -1814
rect 772 -1815 773 -1707
rect 786 -1815 787 -1707
rect 842 -1850 843 -1814
rect 859 -1815 860 -1707
rect 1038 -1850 1039 -1814
rect 1136 -1850 1137 -1814
rect 1178 -1815 1179 -1707
rect 1318 -1850 1319 -1814
rect 1339 -1815 1340 -1707
rect 555 -1850 556 -1816
rect 2427 -1817 2428 -1707
rect 583 -1850 584 -1818
rect 642 -1819 643 -1707
rect 772 -1850 773 -1818
rect 800 -1819 801 -1707
rect 1178 -1850 1179 -1818
rect 1822 -1850 1823 -1818
rect 786 -1850 787 -1820
rect 1087 -1821 1088 -1707
rect 1339 -1850 1340 -1820
rect 2452 -1821 2453 -1707
rect 800 -1850 801 -1822
rect 2067 -1823 2068 -1707
rect 2193 -1823 2194 -1707
rect 2452 -1850 2453 -1822
rect 1087 -1850 1088 -1824
rect 1122 -1825 1123 -1707
rect 2067 -1850 2068 -1824
rect 2256 -1825 2257 -1707
rect 1080 -1827 1081 -1707
rect 1122 -1850 1123 -1826
rect 2144 -1827 2145 -1707
rect 2193 -1850 2194 -1826
rect 2256 -1850 2257 -1826
rect 2431 -1827 2432 -1707
rect 1080 -1850 1081 -1828
rect 1811 -1829 1812 -1707
rect 2109 -1829 2110 -1707
rect 2144 -1850 2145 -1828
rect 2368 -1829 2369 -1707
rect 2431 -1850 2432 -1828
rect 1682 -1831 1683 -1707
rect 2109 -1850 2110 -1830
rect 2277 -1831 2278 -1707
rect 2368 -1850 2369 -1830
rect 1668 -1833 1669 -1707
rect 1682 -1850 1683 -1832
rect 2214 -1833 2215 -1707
rect 2277 -1850 2278 -1832
rect 1654 -1835 1655 -1707
rect 1668 -1850 1669 -1834
rect 1906 -1835 1907 -1707
rect 2214 -1850 2215 -1834
rect 1633 -1837 1634 -1707
rect 1654 -1850 1655 -1836
rect 1864 -1837 1865 -1707
rect 1906 -1850 1907 -1836
rect 1633 -1850 1634 -1838
rect 1766 -1839 1767 -1707
rect 1766 -1850 1767 -1840
rect 1829 -1841 1830 -1707
rect 1780 -1843 1781 -1707
rect 1829 -1850 1830 -1842
rect 1395 -1845 1396 -1707
rect 1780 -1850 1781 -1844
rect 1395 -1850 1396 -1846
rect 1416 -1847 1417 -1707
rect 1416 -1850 1417 -1848
rect 1626 -1850 1627 -1848
rect 30 -1860 31 -1858
rect 611 -1860 612 -1858
rect 618 -1860 619 -1858
rect 1181 -1860 1182 -1858
rect 1206 -1860 1207 -1858
rect 1626 -2025 1627 -1859
rect 1636 -2025 1637 -1859
rect 2368 -1860 2369 -1858
rect 30 -2025 31 -1861
rect 149 -1862 150 -1858
rect 163 -1862 164 -1858
rect 163 -2025 164 -1861
rect 163 -1862 164 -1858
rect 163 -2025 164 -1861
rect 184 -1862 185 -1858
rect 1927 -1862 1928 -1858
rect 2186 -1862 2187 -1858
rect 2186 -2025 2187 -1861
rect 2186 -1862 2187 -1858
rect 2186 -2025 2187 -1861
rect 2270 -1862 2271 -1858
rect 2469 -1862 2470 -1858
rect 37 -1864 38 -1858
rect 618 -2025 619 -1863
rect 632 -1864 633 -1858
rect 1290 -1864 1291 -1858
rect 1307 -1864 1308 -1858
rect 1647 -1864 1648 -1858
rect 1664 -1864 1665 -1858
rect 2109 -1864 2110 -1858
rect 2319 -1864 2320 -1858
rect 2420 -2025 2421 -1863
rect 37 -2025 38 -1865
rect 191 -1866 192 -1858
rect 194 -2025 195 -1865
rect 614 -1866 615 -1858
rect 635 -1866 636 -1858
rect 1199 -1866 1200 -1858
rect 1206 -2025 1207 -1865
rect 1220 -1866 1221 -1858
rect 1241 -1866 1242 -1858
rect 1244 -1942 1245 -1865
rect 1276 -1866 1277 -1858
rect 1962 -1866 1963 -1858
rect 2109 -2025 2110 -1865
rect 2277 -1866 2278 -1858
rect 2319 -2025 2320 -1865
rect 2417 -1866 2418 -1858
rect 47 -1868 48 -1858
rect 2242 -1868 2243 -1858
rect 2368 -2025 2369 -1867
rect 2410 -1868 2411 -1858
rect 72 -1870 73 -1858
rect 800 -1870 801 -1858
rect 814 -1870 815 -1858
rect 814 -2025 815 -1869
rect 814 -1870 815 -1858
rect 814 -2025 815 -1869
rect 835 -1870 836 -1858
rect 835 -2025 836 -1869
rect 835 -1870 836 -1858
rect 835 -2025 836 -1869
rect 852 -1870 853 -1858
rect 1381 -1870 1382 -1858
rect 1437 -1870 1438 -1858
rect 2221 -1870 2222 -1858
rect 2410 -2025 2411 -1869
rect 2459 -1870 2460 -1858
rect 72 -2025 73 -1871
rect 128 -1872 129 -1858
rect 131 -2025 132 -1871
rect 2270 -2025 2271 -1871
rect 89 -2025 90 -1873
rect 1731 -1874 1732 -1858
rect 1734 -2025 1735 -1873
rect 2452 -1874 2453 -1858
rect 100 -1876 101 -1858
rect 187 -1876 188 -1858
rect 215 -2025 216 -1875
rect 1300 -2025 1301 -1875
rect 1332 -1876 1333 -1858
rect 1335 -1876 1336 -1858
rect 1363 -2025 1364 -1875
rect 1934 -1876 1935 -1858
rect 1962 -2025 1963 -1875
rect 1990 -1876 1991 -1858
rect 2067 -1876 2068 -1858
rect 2277 -2025 2278 -1875
rect 100 -2025 101 -1877
rect 1423 -1878 1424 -1858
rect 1468 -1878 1469 -1858
rect 2207 -1878 2208 -1858
rect 2221 -2025 2222 -1877
rect 2284 -1878 2285 -1858
rect 107 -1880 108 -1858
rect 516 -1880 517 -1858
rect 548 -1880 549 -1858
rect 1440 -1880 1441 -1858
rect 1475 -2025 1476 -1879
rect 2249 -1880 2250 -1858
rect 2256 -1880 2257 -1858
rect 2284 -2025 2285 -1879
rect 107 -2025 108 -1881
rect 135 -1882 136 -1858
rect 142 -1882 143 -1858
rect 1153 -2025 1154 -1881
rect 1164 -1882 1165 -1858
rect 1220 -2025 1221 -1881
rect 1241 -2025 1242 -1881
rect 1332 -2025 1333 -1881
rect 1339 -1882 1340 -1858
rect 1353 -1882 1354 -1858
rect 1423 -2025 1424 -1881
rect 1489 -2025 1490 -1881
rect 1577 -1882 1578 -1858
rect 1622 -2025 1623 -1881
rect 1955 -1882 1956 -1858
rect 2067 -2025 2068 -1881
rect 2123 -1882 2124 -1858
rect 2249 -2025 2250 -1881
rect 2291 -1882 2292 -1858
rect 103 -2025 104 -1883
rect 135 -2025 136 -1883
rect 142 -2025 143 -1883
rect 380 -1884 381 -1858
rect 401 -1884 402 -1858
rect 649 -1884 650 -1858
rect 688 -1884 689 -1858
rect 730 -1884 731 -1858
rect 737 -1884 738 -1858
rect 1024 -1884 1025 -1858
rect 1059 -1884 1060 -1858
rect 1069 -1942 1070 -1883
rect 1094 -1884 1095 -1858
rect 1731 -2025 1732 -1883
rect 1773 -1884 1774 -1858
rect 1990 -2025 1991 -1883
rect 2256 -2025 2257 -1883
rect 2305 -1884 2306 -1858
rect 16 -1886 17 -1858
rect 1094 -2025 1095 -1885
rect 1136 -1886 1137 -1858
rect 2088 -1886 2089 -1858
rect 16 -2025 17 -1887
rect 352 -1888 353 -1858
rect 373 -1888 374 -1858
rect 586 -2025 587 -1887
rect 611 -2025 612 -1887
rect 681 -1888 682 -1858
rect 688 -2025 689 -1887
rect 786 -1888 787 -1858
rect 894 -1888 895 -1858
rect 1997 -1888 1998 -1858
rect 124 -1890 125 -1858
rect 1101 -1890 1102 -1858
rect 1129 -1890 1130 -1858
rect 1136 -2025 1137 -1889
rect 1150 -1890 1151 -1858
rect 1199 -2025 1200 -1889
rect 1209 -1890 1210 -1858
rect 2445 -1890 2446 -1858
rect 128 -2025 129 -1891
rect 1073 -1892 1074 -1858
rect 1080 -1892 1081 -1858
rect 1101 -2025 1102 -1891
rect 1129 -2025 1130 -1891
rect 1139 -1892 1140 -1858
rect 1164 -2025 1165 -1891
rect 1458 -1892 1459 -1858
rect 1507 -1892 1508 -1858
rect 2389 -1892 2390 -1858
rect 184 -2025 185 -1893
rect 219 -1894 220 -1858
rect 233 -1894 234 -1858
rect 2123 -2025 2124 -1893
rect 2228 -1894 2229 -1858
rect 2389 -2025 2390 -1893
rect 177 -1896 178 -1858
rect 233 -2025 234 -1895
rect 250 -1896 251 -1858
rect 1430 -1896 1431 -1858
rect 1440 -2025 1441 -1895
rect 2291 -2025 2292 -1895
rect 177 -2025 178 -1897
rect 261 -1898 262 -1858
rect 275 -1898 276 -1858
rect 429 -1898 430 -1858
rect 446 -1898 447 -1858
rect 464 -1898 465 -1858
rect 478 -1898 479 -1858
rect 782 -2025 783 -1897
rect 905 -2025 906 -1897
rect 1612 -1898 1613 -1858
rect 1633 -1898 1634 -1858
rect 1997 -2025 1998 -1897
rect 2032 -1898 2033 -1858
rect 2228 -2025 2229 -1897
rect 205 -1900 206 -1858
rect 380 -2025 381 -1899
rect 401 -2025 402 -1899
rect 632 -2025 633 -1899
rect 646 -1900 647 -1858
rect 1269 -1900 1270 -1858
rect 1290 -2025 1291 -1899
rect 1297 -1900 1298 -1858
rect 1304 -1900 1305 -1858
rect 2207 -2025 2208 -1899
rect 205 -2025 206 -1901
rect 282 -1902 283 -1858
rect 303 -1902 304 -1858
rect 352 -2025 353 -1901
rect 373 -2025 374 -1901
rect 821 -1902 822 -1858
rect 908 -1902 909 -1858
rect 947 -1902 948 -1858
rect 957 -1902 958 -1858
rect 1843 -1902 1844 -1858
rect 1853 -1902 1854 -1858
rect 2424 -1902 2425 -1858
rect 51 -1904 52 -1858
rect 282 -2025 283 -1903
rect 303 -2025 304 -1903
rect 450 -1904 451 -1858
rect 464 -2025 465 -1903
rect 527 -1904 528 -1858
rect 541 -1904 542 -1858
rect 730 -2025 731 -1903
rect 744 -1904 745 -1858
rect 1276 -2025 1277 -1903
rect 1339 -2025 1340 -1903
rect 1367 -1904 1368 -1858
rect 1381 -2025 1382 -1903
rect 1416 -1904 1417 -1858
rect 1430 -2025 1431 -1903
rect 1451 -1904 1452 -1858
rect 1458 -2025 1459 -1903
rect 1472 -1904 1473 -1858
rect 1507 -2025 1508 -1903
rect 1584 -1904 1585 -1858
rect 1605 -1904 1606 -1858
rect 1612 -2025 1613 -1903
rect 1647 -2025 1648 -1903
rect 1850 -1904 1851 -1858
rect 1864 -1904 1865 -1858
rect 2403 -1904 2404 -1858
rect 51 -2025 52 -1905
rect 1605 -2025 1606 -1905
rect 1664 -2025 1665 -1905
rect 2375 -1906 2376 -1858
rect 2403 -2025 2404 -1905
rect 2438 -1906 2439 -1858
rect 219 -2025 220 -1907
rect 1521 -1908 1522 -1858
rect 1528 -1908 1529 -1858
rect 1528 -2025 1529 -1907
rect 1528 -1908 1529 -1858
rect 1528 -2025 1529 -1907
rect 1577 -2025 1578 -1907
rect 1591 -1908 1592 -1858
rect 1773 -2025 1774 -1907
rect 1822 -1908 1823 -1858
rect 1843 -2025 1844 -1907
rect 2081 -1908 2082 -1858
rect 226 -1910 227 -1858
rect 2375 -2025 2376 -1909
rect 170 -1912 171 -1858
rect 226 -2025 227 -1911
rect 261 -2025 262 -1911
rect 268 -1912 269 -1858
rect 275 -2025 276 -1911
rect 541 -2025 542 -1911
rect 562 -1912 563 -1858
rect 1108 -1912 1109 -1858
rect 1167 -2025 1168 -1911
rect 2305 -2025 2306 -1911
rect 156 -2025 157 -1913
rect 268 -2025 269 -1913
rect 394 -1914 395 -1858
rect 527 -2025 528 -1913
rect 565 -1914 566 -1858
rect 1052 -1914 1053 -1858
rect 1059 -2025 1060 -1913
rect 1346 -1914 1347 -1858
rect 1353 -2025 1354 -1913
rect 1402 -1914 1403 -1858
rect 1416 -2025 1417 -1913
rect 1500 -1914 1501 -1858
rect 1584 -2025 1585 -1913
rect 1619 -1914 1620 -1858
rect 1822 -2025 1823 -1913
rect 1836 -1914 1837 -1858
rect 1850 -2025 1851 -1913
rect 1878 -1914 1879 -1858
rect 1934 -2025 1935 -1913
rect 1969 -1914 1970 -1858
rect 2032 -2025 2033 -1913
rect 2144 -1914 2145 -1858
rect 170 -2025 171 -1915
rect 2158 -1916 2159 -1858
rect 173 -2025 174 -1917
rect 2158 -2025 2159 -1917
rect 229 -1920 230 -1858
rect 1836 -2025 1837 -1919
rect 1864 -2025 1865 -1919
rect 1899 -1920 1900 -1858
rect 1941 -1920 1942 -1858
rect 2144 -2025 2145 -1919
rect 240 -1922 241 -1858
rect 394 -2025 395 -1921
rect 422 -1922 423 -1858
rect 548 -2025 549 -1921
rect 569 -1922 570 -1858
rect 740 -1922 741 -1858
rect 744 -2025 745 -1921
rect 807 -1922 808 -1858
rect 821 -2025 822 -1921
rect 940 -1922 941 -1858
rect 943 -1922 944 -1858
rect 1185 -1922 1186 -1858
rect 1227 -1922 1228 -1858
rect 1269 -2025 1270 -1921
rect 1346 -2025 1347 -1921
rect 1570 -1922 1571 -1858
rect 1591 -2025 1592 -1921
rect 1780 -1922 1781 -1858
rect 1878 -2025 1879 -1921
rect 1913 -1922 1914 -1858
rect 1941 -2025 1942 -1921
rect 1983 -1922 1984 -1858
rect 2081 -2025 2082 -1921
rect 2137 -1922 2138 -1858
rect 2 -1924 3 -1858
rect 240 -2025 241 -1923
rect 422 -2025 423 -1923
rect 544 -2025 545 -1923
rect 646 -2025 647 -1923
rect 863 -1924 864 -1858
rect 919 -1924 920 -1858
rect 947 -2025 948 -1923
rect 957 -2025 958 -1923
rect 2242 -2025 2243 -1923
rect 2 -2025 3 -1925
rect 737 -2025 738 -1925
rect 807 -2025 808 -1925
rect 1010 -1926 1011 -1858
rect 1024 -2025 1025 -1925
rect 1437 -2025 1438 -1925
rect 1444 -1926 1445 -1858
rect 1570 -2025 1571 -1925
rect 1780 -2025 1781 -1925
rect 1829 -1926 1830 -1858
rect 1899 -2025 1900 -1925
rect 2466 -1926 2467 -1858
rect 159 -1928 160 -1858
rect 1010 -2025 1011 -1927
rect 1038 -1928 1039 -1858
rect 1080 -2025 1081 -1927
rect 1178 -1928 1179 -1858
rect 2333 -1928 2334 -1858
rect 9 -1930 10 -1858
rect 159 -2025 160 -1929
rect 429 -2025 430 -1929
rect 499 -1930 500 -1858
rect 506 -1930 507 -1858
rect 740 -2025 741 -1929
rect 863 -2025 864 -1929
rect 975 -1930 976 -1858
rect 978 -2025 979 -1929
rect 1510 -1930 1511 -1858
rect 1913 -2025 1914 -1929
rect 1948 -1930 1949 -1858
rect 1955 -2025 1956 -1929
rect 2011 -1930 2012 -1858
rect 2074 -1930 2075 -1858
rect 2333 -2025 2334 -1929
rect 9 -2025 10 -1931
rect 198 -1932 199 -1858
rect 324 -1932 325 -1858
rect 499 -2025 500 -1931
rect 506 -2025 507 -1931
rect 877 -1932 878 -1858
rect 919 -2025 920 -1931
rect 1122 -1932 1123 -1858
rect 1178 -2025 1179 -1931
rect 1629 -1932 1630 -1858
rect 1696 -1932 1697 -1858
rect 1948 -2025 1949 -1931
rect 1969 -2025 1970 -1931
rect 2004 -1932 2005 -1858
rect 2011 -2025 2012 -1931
rect 2060 -1932 2061 -1858
rect 2074 -2025 2075 -1931
rect 2130 -1932 2131 -1858
rect 2137 -2025 2138 -1931
rect 2193 -1932 2194 -1858
rect 58 -1934 59 -1858
rect 1038 -2025 1039 -1933
rect 1062 -2025 1063 -1933
rect 2298 -1934 2299 -1858
rect 23 -1936 24 -1858
rect 58 -2025 59 -1935
rect 198 -2025 199 -1935
rect 1003 -1936 1004 -1858
rect 1066 -1936 1067 -1858
rect 1619 -2025 1620 -1935
rect 1696 -2025 1697 -1935
rect 1703 -1936 1704 -1858
rect 1983 -2025 1984 -1935
rect 2025 -1936 2026 -1858
rect 2060 -2025 2061 -1935
rect 2116 -1936 2117 -1858
rect 2130 -2025 2131 -1935
rect 2172 -1936 2173 -1858
rect 2298 -2025 2299 -1935
rect 2312 -1936 2313 -1858
rect 23 -2025 24 -1937
rect 114 -1938 115 -1858
rect 324 -2025 325 -1937
rect 1465 -1938 1466 -1858
rect 1472 -2025 1473 -1937
rect 2424 -2025 2425 -1937
rect 114 -2025 115 -1939
rect 758 -1940 759 -1858
rect 828 -1940 829 -1858
rect 877 -2025 878 -1939
rect 926 -1940 927 -1858
rect 1304 -2025 1305 -1939
rect 1367 -2025 1368 -1939
rect 1409 -1940 1410 -1858
rect 1444 -2025 1445 -1939
rect 1479 -1940 1480 -1858
rect 1486 -1940 1487 -1858
rect 1500 -2025 1501 -1939
rect 1703 -2025 1704 -1939
rect 1885 -1940 1886 -1858
rect 1892 -1940 1893 -1858
rect 2116 -2025 2117 -1939
rect 2312 -2025 2313 -1939
rect 2347 -1940 2348 -1858
rect 432 -1942 433 -1858
rect 569 -2025 570 -1941
rect 674 -1942 675 -1858
rect 681 -2025 682 -1941
rect 695 -1942 696 -1858
rect 1003 -2025 1004 -1941
rect 1066 -2025 1067 -1941
rect 1115 -1942 1116 -1858
rect 1185 -2025 1186 -1941
rect 1318 -1942 1319 -1858
rect 1335 -2025 1336 -1941
rect 1409 -2025 1410 -1941
rect 1451 -2025 1452 -1941
rect 1598 -1942 1599 -1858
rect 1724 -1942 1725 -1858
rect 2025 -2025 2026 -1941
rect 2347 -2025 2348 -1941
rect 2382 -1942 2383 -1858
rect 191 -2025 192 -1943
rect 674 -2025 675 -1943
rect 702 -1944 703 -1858
rect 954 -1944 955 -1858
rect 961 -1944 962 -1858
rect 961 -2025 962 -1943
rect 961 -1944 962 -1858
rect 961 -2025 962 -1943
rect 975 -2025 976 -1943
rect 1752 -1944 1753 -1858
rect 1766 -1944 1767 -1858
rect 1885 -2025 1886 -1943
rect 1892 -2025 1893 -1943
rect 2165 -1944 2166 -1858
rect 2179 -1944 2180 -1858
rect 2382 -2025 2383 -1943
rect 450 -2025 451 -1945
rect 590 -1946 591 -1858
rect 660 -1946 661 -1858
rect 695 -2025 696 -1945
rect 702 -2025 703 -1945
rect 996 -1946 997 -1858
rect 1073 -2025 1074 -1945
rect 1867 -1946 1868 -1858
rect 1976 -1946 1977 -1858
rect 2172 -2025 2173 -1945
rect 2179 -2025 2180 -1945
rect 2235 -1946 2236 -1858
rect 121 -1948 122 -1858
rect 660 -2025 661 -1947
rect 709 -1948 710 -1858
rect 940 -2025 941 -1947
rect 982 -1948 983 -1858
rect 996 -2025 997 -1947
rect 1087 -1948 1088 -1858
rect 1115 -2025 1116 -1947
rect 1125 -2025 1126 -1947
rect 1976 -2025 1977 -1947
rect 2004 -2025 2005 -1947
rect 2053 -1948 2054 -1858
rect 86 -1950 87 -1858
rect 982 -2025 983 -1949
rect 1111 -2025 1112 -1949
rect 2193 -2025 2194 -1949
rect 121 -2025 122 -1951
rect 296 -1952 297 -1858
rect 443 -1952 444 -1858
rect 1087 -2025 1088 -1951
rect 1227 -2025 1228 -1951
rect 2235 -2025 2236 -1951
rect 296 -2025 297 -1953
rect 359 -1954 360 -1858
rect 443 -2025 444 -1953
rect 555 -1954 556 -1858
rect 590 -2025 591 -1953
rect 726 -1954 727 -1858
rect 772 -1954 773 -1858
rect 954 -2025 955 -1953
rect 1248 -1954 1249 -1858
rect 1829 -2025 1830 -1953
rect 2053 -2025 2054 -1953
rect 2102 -1954 2103 -1858
rect 289 -1956 290 -1858
rect 555 -2025 556 -1955
rect 653 -1956 654 -1858
rect 709 -2025 710 -1955
rect 723 -1956 724 -1858
rect 758 -2025 759 -1955
rect 772 -2025 773 -1955
rect 922 -2025 923 -1955
rect 926 -2025 927 -1955
rect 1045 -1956 1046 -1858
rect 1213 -1956 1214 -1858
rect 1248 -2025 1249 -1955
rect 1395 -1956 1396 -1858
rect 1402 -2025 1403 -1955
rect 1465 -2025 1466 -1955
rect 1633 -2025 1634 -1955
rect 1654 -1956 1655 -1858
rect 1724 -2025 1725 -1955
rect 1752 -2025 1753 -1955
rect 1759 -1956 1760 -1858
rect 1766 -2025 1767 -1955
rect 1815 -1956 1816 -1858
rect 2102 -2025 2103 -1955
rect 2151 -1956 2152 -1858
rect 289 -2025 290 -1957
rect 849 -1958 850 -1858
rect 933 -1958 934 -1858
rect 1318 -2025 1319 -1957
rect 1360 -1958 1361 -1858
rect 1395 -2025 1396 -1957
rect 1486 -2025 1487 -1957
rect 1927 -2025 1928 -1957
rect 2151 -2025 2152 -1957
rect 2200 -1958 2201 -1858
rect 359 -2025 360 -1959
rect 436 -1960 437 -1858
rect 478 -2025 479 -1959
rect 604 -1960 605 -1858
rect 653 -2025 654 -1959
rect 842 -1960 843 -1858
rect 849 -2025 850 -1959
rect 898 -1960 899 -1858
rect 933 -2025 934 -1959
rect 2473 -1960 2474 -1858
rect 436 -2025 437 -1961
rect 597 -1962 598 -1858
rect 604 -2025 605 -1961
rect 751 -1962 752 -1858
rect 842 -2025 843 -1961
rect 856 -1962 857 -1858
rect 1017 -1962 1018 -1858
rect 1045 -2025 1046 -1961
rect 1213 -2025 1214 -1961
rect 1234 -1962 1235 -1858
rect 1279 -1962 1280 -1858
rect 1815 -2025 1816 -1961
rect 310 -1964 311 -1858
rect 1017 -2025 1018 -1963
rect 1234 -2025 1235 -1963
rect 1311 -1964 1312 -1858
rect 1360 -2025 1361 -1963
rect 2088 -2025 2089 -1963
rect 310 -2025 311 -1965
rect 317 -1966 318 -1858
rect 485 -1966 486 -1858
rect 562 -2025 563 -1965
rect 576 -1966 577 -1858
rect 856 -2025 857 -1965
rect 1297 -2025 1298 -1965
rect 2200 -2025 2201 -1965
rect 212 -1968 213 -1858
rect 317 -2025 318 -1967
rect 485 -2025 486 -1967
rect 492 -1968 493 -1858
rect 513 -1968 514 -1858
rect 803 -1968 804 -1858
rect 1311 -2025 1312 -1967
rect 1661 -1968 1662 -1858
rect 1675 -1968 1676 -1858
rect 1759 -2025 1760 -1967
rect 1801 -1968 1802 -1858
rect 2165 -2025 2166 -1967
rect 149 -2025 150 -1969
rect 212 -2025 213 -1969
rect 247 -1970 248 -1858
rect 492 -2025 493 -1969
rect 534 -1970 535 -1858
rect 597 -2025 598 -1969
rect 625 -1970 626 -1858
rect 898 -2025 899 -1969
rect 1549 -1970 1550 -1858
rect 1598 -2025 1599 -1969
rect 1654 -2025 1655 -1969
rect 1745 -1970 1746 -1858
rect 1801 -2025 1802 -1969
rect 1857 -1970 1858 -1858
rect 86 -2025 87 -1971
rect 247 -2025 248 -1971
rect 387 -1972 388 -1858
rect 513 -2025 514 -1971
rect 576 -2025 577 -1971
rect 793 -1972 794 -1858
rect 1524 -2025 1525 -1971
rect 1745 -2025 1746 -1971
rect 93 -1974 94 -1858
rect 534 -2025 535 -1973
rect 716 -1974 717 -1858
rect 723 -2025 724 -1973
rect 751 -2025 752 -1973
rect 891 -1974 892 -1858
rect 1535 -1974 1536 -1858
rect 1857 -2025 1858 -1973
rect 93 -2025 94 -1975
rect 338 -1976 339 -1858
rect 387 -2025 388 -1975
rect 415 -1976 416 -1858
rect 457 -1976 458 -1858
rect 625 -2025 626 -1975
rect 639 -1976 640 -1858
rect 716 -2025 717 -1975
rect 793 -2025 794 -1975
rect 1108 -2025 1109 -1975
rect 1549 -2025 1550 -1975
rect 2340 -1976 2341 -1858
rect 79 -1978 80 -1858
rect 639 -2025 640 -1977
rect 828 -2025 829 -1977
rect 2340 -2025 2341 -1977
rect 79 -2025 80 -1979
rect 831 -2025 832 -1979
rect 870 -1980 871 -1858
rect 891 -2025 892 -1979
rect 1052 -2025 1053 -1979
rect 1535 -2025 1536 -1979
rect 1661 -2025 1662 -1979
rect 2326 -1980 2327 -1858
rect 254 -1982 255 -1858
rect 457 -2025 458 -1981
rect 870 -2025 871 -1981
rect 912 -1982 913 -1858
rect 1675 -2025 1676 -1981
rect 1682 -1982 1683 -1858
rect 2326 -2025 2327 -1981
rect 2361 -1982 2362 -1858
rect 44 -1984 45 -1858
rect 254 -2025 255 -1983
rect 331 -1984 332 -1858
rect 338 -2025 339 -1983
rect 345 -1984 346 -1858
rect 415 -2025 416 -1983
rect 583 -1984 584 -1858
rect 912 -2025 913 -1983
rect 1682 -2025 1683 -1983
rect 1689 -1984 1690 -1858
rect 2361 -2025 2362 -1983
rect 2396 -1984 2397 -1858
rect 44 -2025 45 -1985
rect 65 -1986 66 -1858
rect 331 -2025 332 -1985
rect 1262 -1986 1263 -1858
rect 1689 -2025 1690 -1985
rect 1710 -1986 1711 -1858
rect 1787 -1986 1788 -1858
rect 2396 -2025 2397 -1985
rect 65 -2025 66 -1987
rect 1374 -1988 1375 -1858
rect 1563 -1988 1564 -1858
rect 1787 -2025 1788 -1987
rect 345 -2025 346 -1989
rect 366 -1990 367 -1858
rect 583 -2025 584 -1989
rect 786 -2025 787 -1989
rect 1255 -1990 1256 -1858
rect 1262 -2025 1263 -1989
rect 1283 -1990 1284 -1858
rect 1563 -2025 1564 -1989
rect 1710 -2025 1711 -1989
rect 1738 -1990 1739 -1858
rect 366 -2025 367 -1991
rect 408 -1992 409 -1858
rect 1171 -1992 1172 -1858
rect 1255 -2025 1256 -1991
rect 1374 -2025 1375 -1991
rect 1388 -1992 1389 -1858
rect 1640 -1992 1641 -1858
rect 1738 -2025 1739 -1991
rect 408 -2025 409 -1993
rect 471 -1994 472 -1858
rect 765 -1994 766 -1858
rect 1171 -2025 1172 -1993
rect 1192 -1994 1193 -1858
rect 1283 -2025 1284 -1993
rect 1388 -2025 1389 -1993
rect 1496 -2025 1497 -1993
rect 1556 -1994 1557 -1858
rect 1640 -2025 1641 -1993
rect 471 -2025 472 -1995
rect 520 -1996 521 -1858
rect 765 -2025 766 -1995
rect 1031 -1996 1032 -1858
rect 1157 -1996 1158 -1858
rect 1192 -2025 1193 -1995
rect 1514 -1996 1515 -1858
rect 1556 -2025 1557 -1995
rect 520 -2025 521 -1997
rect 667 -1998 668 -1858
rect 989 -1998 990 -1858
rect 1031 -2025 1032 -1997
rect 1143 -1998 1144 -1858
rect 1157 -2025 1158 -1997
rect 1514 -2025 1515 -1997
rect 1542 -1998 1543 -1858
rect 635 -2025 636 -1999
rect 667 -2025 668 -1999
rect 779 -2000 780 -1858
rect 1143 -2025 1144 -1999
rect 1493 -2000 1494 -1858
rect 1542 -2025 1543 -1999
rect 968 -2002 969 -1858
rect 989 -2025 990 -2001
rect 1493 -2025 1494 -2001
rect 2214 -2002 2215 -1858
rect 884 -2004 885 -1858
rect 968 -2025 969 -2003
rect 2214 -2025 2215 -2003
rect 2263 -2004 2264 -1858
rect 884 -2025 885 -2005
rect 1668 -2006 1669 -1858
rect 2039 -2006 2040 -1858
rect 2263 -2025 2264 -2005
rect 1668 -2025 1669 -2007
rect 1794 -2008 1795 -1858
rect 2039 -2025 2040 -2007
rect 2095 -2008 2096 -1858
rect 1794 -2025 1795 -2009
rect 2018 -2010 2019 -1858
rect 2095 -2025 2096 -2009
rect 2354 -2010 2355 -1858
rect 1808 -2012 1809 -1858
rect 2018 -2025 2019 -2011
rect 2354 -2025 2355 -2011
rect 2431 -2012 2432 -1858
rect 1808 -2025 1809 -2013
rect 1871 -2014 1872 -1858
rect 1871 -2025 1872 -2015
rect 1906 -2016 1907 -1858
rect 1906 -2025 1907 -2017
rect 1920 -2018 1921 -1858
rect 1920 -2025 1921 -2019
rect 2046 -2020 2047 -1858
rect 1717 -2022 1718 -1858
rect 2046 -2025 2047 -2021
rect 779 -2025 780 -2023
rect 1717 -2025 1718 -2023
rect 9 -2035 10 -2033
rect 761 -2176 762 -2034
rect 800 -2035 801 -2033
rect 849 -2035 850 -2033
rect 898 -2035 899 -2033
rect 1108 -2035 1109 -2033
rect 1111 -2035 1112 -2033
rect 1206 -2035 1207 -2033
rect 1230 -2035 1231 -2033
rect 1300 -2035 1301 -2033
rect 1335 -2176 1336 -2034
rect 1976 -2035 1977 -2033
rect 2368 -2035 2369 -2033
rect 2368 -2176 2369 -2034
rect 2368 -2035 2369 -2033
rect 2368 -2176 2369 -2034
rect 2403 -2035 2404 -2033
rect 2417 -2176 2418 -2034
rect 9 -2176 10 -2036
rect 44 -2037 45 -2033
rect 51 -2037 52 -2033
rect 65 -2037 66 -2033
rect 86 -2176 87 -2036
rect 135 -2037 136 -2033
rect 138 -2176 139 -2036
rect 1017 -2037 1018 -2033
rect 1024 -2037 1025 -2033
rect 1108 -2176 1109 -2036
rect 1115 -2037 1116 -2033
rect 1115 -2176 1116 -2036
rect 1115 -2037 1116 -2033
rect 1115 -2176 1116 -2036
rect 1122 -2037 1123 -2033
rect 1423 -2037 1424 -2033
rect 1437 -2037 1438 -2033
rect 2424 -2037 2425 -2033
rect 37 -2039 38 -2033
rect 831 -2039 832 -2033
rect 898 -2176 899 -2038
rect 1304 -2039 1305 -2033
rect 1360 -2039 1361 -2033
rect 1640 -2039 1641 -2033
rect 1713 -2176 1714 -2038
rect 1969 -2039 1970 -2033
rect 37 -2176 38 -2040
rect 240 -2041 241 -2033
rect 296 -2041 297 -2033
rect 1062 -2041 1063 -2033
rect 1073 -2041 1074 -2033
rect 1206 -2176 1207 -2040
rect 1297 -2041 1298 -2033
rect 1857 -2041 1858 -2033
rect 1934 -2041 1935 -2033
rect 2403 -2176 2404 -2040
rect 30 -2043 31 -2033
rect 240 -2176 241 -2042
rect 296 -2176 297 -2042
rect 471 -2043 472 -2033
rect 492 -2043 493 -2033
rect 1017 -2176 1018 -2042
rect 1024 -2176 1025 -2042
rect 1430 -2043 1431 -2033
rect 1437 -2176 1438 -2042
rect 1444 -2043 1445 -2033
rect 1472 -2176 1473 -2042
rect 1878 -2043 1879 -2033
rect 1969 -2176 1970 -2042
rect 2375 -2043 2376 -2033
rect 16 -2045 17 -2033
rect 471 -2176 472 -2044
rect 499 -2045 500 -2033
rect 541 -2176 542 -2044
rect 569 -2045 570 -2033
rect 1122 -2176 1123 -2044
rect 1150 -2176 1151 -2044
rect 2291 -2045 2292 -2033
rect 2340 -2045 2341 -2033
rect 2375 -2176 2376 -2044
rect 16 -2176 17 -2046
rect 807 -2047 808 -2033
rect 828 -2047 829 -2033
rect 1409 -2047 1410 -2033
rect 1430 -2176 1431 -2046
rect 1983 -2047 1984 -2033
rect 2249 -2047 2250 -2033
rect 2291 -2176 2292 -2046
rect 2298 -2047 2299 -2033
rect 2340 -2176 2341 -2046
rect 30 -2176 31 -2048
rect 72 -2049 73 -2033
rect 89 -2049 90 -2033
rect 884 -2049 885 -2033
rect 919 -2049 920 -2033
rect 926 -2049 927 -2033
rect 954 -2049 955 -2033
rect 2354 -2049 2355 -2033
rect 44 -2176 45 -2050
rect 695 -2051 696 -2033
rect 751 -2051 752 -2033
rect 849 -2176 850 -2050
rect 922 -2051 923 -2033
rect 1031 -2051 1032 -2033
rect 1087 -2051 1088 -2033
rect 1087 -2176 1088 -2050
rect 1087 -2051 1088 -2033
rect 1087 -2176 1088 -2050
rect 1153 -2051 1154 -2033
rect 1395 -2051 1396 -2033
rect 1402 -2051 1403 -2033
rect 1423 -2176 1424 -2050
rect 1440 -2051 1441 -2033
rect 2116 -2051 2117 -2033
rect 2214 -2051 2215 -2033
rect 2249 -2176 2250 -2050
rect 2 -2053 3 -2033
rect 1153 -2176 1154 -2052
rect 1171 -2053 1172 -2033
rect 1342 -2176 1343 -2052
rect 1363 -2053 1364 -2033
rect 2228 -2053 2229 -2033
rect 51 -2176 52 -2054
rect 1696 -2055 1697 -2033
rect 1766 -2055 1767 -2033
rect 2424 -2176 2425 -2054
rect 58 -2057 59 -2033
rect 1360 -2176 1361 -2056
rect 1384 -2176 1385 -2056
rect 1598 -2057 1599 -2033
rect 1605 -2057 1606 -2033
rect 1696 -2176 1697 -2056
rect 1808 -2057 1809 -2033
rect 1878 -2176 1879 -2056
rect 2095 -2057 2096 -2033
rect 2354 -2176 2355 -2056
rect 58 -2176 59 -2058
rect 96 -2176 97 -2058
rect 100 -2059 101 -2033
rect 107 -2059 108 -2033
rect 156 -2059 157 -2033
rect 2305 -2059 2306 -2033
rect 65 -2176 66 -2060
rect 702 -2061 703 -2033
rect 758 -2061 759 -2033
rect 803 -2061 804 -2033
rect 807 -2176 808 -2060
rect 1318 -2061 1319 -2033
rect 1402 -2176 1403 -2060
rect 2025 -2061 2026 -2033
rect 2095 -2176 2096 -2060
rect 2186 -2061 2187 -2033
rect 2228 -2176 2229 -2060
rect 2284 -2061 2285 -2033
rect 2305 -2176 2306 -2060
rect 2312 -2061 2313 -2033
rect 72 -2176 73 -2062
rect 961 -2063 962 -2033
rect 1031 -2176 1032 -2062
rect 1129 -2063 1130 -2033
rect 1178 -2063 1179 -2033
rect 1640 -2176 1641 -2062
rect 1654 -2063 1655 -2033
rect 1808 -2176 1809 -2062
rect 1815 -2063 1816 -2033
rect 1976 -2176 1977 -2062
rect 2046 -2063 2047 -2033
rect 2312 -2176 2313 -2062
rect 100 -2176 101 -2064
rect 1405 -2176 1406 -2064
rect 1409 -2176 1410 -2064
rect 1885 -2065 1886 -2033
rect 1920 -2065 1921 -2033
rect 2046 -2176 2047 -2064
rect 2116 -2176 2117 -2064
rect 2130 -2065 2131 -2033
rect 2172 -2065 2173 -2033
rect 2214 -2176 2215 -2064
rect 2256 -2065 2257 -2033
rect 2284 -2176 2285 -2064
rect 107 -2176 108 -2066
rect 1167 -2067 1168 -2033
rect 1178 -2176 1179 -2066
rect 1192 -2067 1193 -2033
rect 1220 -2067 1221 -2033
rect 1318 -2176 1319 -2066
rect 1486 -2067 1487 -2033
rect 1990 -2067 1991 -2033
rect 2074 -2067 2075 -2033
rect 2130 -2176 2131 -2066
rect 2137 -2067 2138 -2033
rect 2172 -2176 2173 -2066
rect 2186 -2176 2187 -2066
rect 2347 -2067 2348 -2033
rect 156 -2176 157 -2068
rect 457 -2069 458 -2033
rect 516 -2176 517 -2068
rect 1003 -2069 1004 -2033
rect 1038 -2069 1039 -2033
rect 1129 -2176 1130 -2068
rect 1192 -2176 1193 -2068
rect 1290 -2069 1291 -2033
rect 1297 -2176 1298 -2068
rect 1307 -2176 1308 -2068
rect 1486 -2176 1487 -2068
rect 1724 -2069 1725 -2033
rect 1745 -2069 1746 -2033
rect 1815 -2176 1816 -2068
rect 1871 -2069 1872 -2033
rect 1920 -2176 1921 -2068
rect 1948 -2069 1949 -2033
rect 1990 -2176 1991 -2068
rect 2018 -2069 2019 -2033
rect 2074 -2176 2075 -2068
rect 2081 -2069 2082 -2033
rect 2137 -2176 2138 -2068
rect 2207 -2069 2208 -2033
rect 2256 -2176 2257 -2068
rect 2333 -2069 2334 -2033
rect 2347 -2176 2348 -2068
rect 159 -2071 160 -2033
rect 905 -2071 906 -2033
rect 1003 -2176 1004 -2070
rect 1255 -2071 1256 -2033
rect 1269 -2071 1270 -2033
rect 1983 -2176 1984 -2070
rect 173 -2073 174 -2033
rect 1241 -2073 1242 -2033
rect 1276 -2073 1277 -2033
rect 1395 -2176 1396 -2072
rect 1489 -2073 1490 -2033
rect 2298 -2176 2299 -2072
rect 191 -2075 192 -2033
rect 506 -2075 507 -2033
rect 569 -2176 570 -2074
rect 978 -2075 979 -2033
rect 1038 -2176 1039 -2074
rect 1066 -2075 1067 -2033
rect 1080 -2075 1081 -2033
rect 1171 -2176 1172 -2074
rect 1234 -2075 1235 -2033
rect 1444 -2176 1445 -2074
rect 1521 -2075 1522 -2033
rect 1759 -2075 1760 -2033
rect 1843 -2075 1844 -2033
rect 2081 -2176 2082 -2074
rect 191 -2176 192 -2076
rect 586 -2077 587 -2033
rect 590 -2077 591 -2033
rect 656 -2176 657 -2076
rect 670 -2176 671 -2076
rect 744 -2077 745 -2033
rect 758 -2176 759 -2076
rect 884 -2176 885 -2076
rect 891 -2077 892 -2033
rect 905 -2176 906 -2076
rect 978 -2176 979 -2076
rect 1822 -2077 1823 -2033
rect 1871 -2176 1872 -2076
rect 1941 -2077 1942 -2033
rect 1955 -2077 1956 -2033
rect 2018 -2176 2019 -2076
rect 170 -2079 171 -2033
rect 590 -2176 591 -2078
rect 604 -2079 605 -2033
rect 779 -2079 780 -2033
rect 786 -2079 787 -2033
rect 800 -2176 801 -2078
rect 828 -2176 829 -2078
rect 968 -2079 969 -2033
rect 989 -2079 990 -2033
rect 1234 -2176 1235 -2078
rect 1283 -2079 1284 -2033
rect 1290 -2176 1291 -2078
rect 1304 -2176 1305 -2078
rect 1416 -2079 1417 -2033
rect 1521 -2176 1522 -2078
rect 1612 -2079 1613 -2033
rect 1622 -2079 1623 -2033
rect 2032 -2079 2033 -2033
rect 170 -2176 171 -2080
rect 730 -2081 731 -2033
rect 740 -2081 741 -2033
rect 2025 -2176 2026 -2080
rect 194 -2083 195 -2033
rect 1724 -2176 1725 -2082
rect 1752 -2083 1753 -2033
rect 1822 -2176 1823 -2082
rect 1899 -2083 1900 -2033
rect 1941 -2176 1942 -2082
rect 1955 -2176 1956 -2082
rect 2389 -2083 2390 -2033
rect 212 -2085 213 -2033
rect 317 -2085 318 -2033
rect 331 -2085 332 -2033
rect 961 -2176 962 -2084
rect 1059 -2085 1060 -2033
rect 2333 -2176 2334 -2084
rect 2361 -2085 2362 -2033
rect 2389 -2176 2390 -2084
rect 93 -2087 94 -2033
rect 331 -2176 332 -2086
rect 338 -2087 339 -2033
rect 457 -2176 458 -2086
rect 464 -2087 465 -2033
rect 604 -2176 605 -2086
rect 618 -2087 619 -2033
rect 751 -2176 752 -2086
rect 793 -2087 794 -2033
rect 926 -2176 927 -2086
rect 940 -2087 941 -2033
rect 989 -2176 990 -2086
rect 1066 -2176 1067 -2086
rect 1664 -2087 1665 -2033
rect 1689 -2087 1690 -2033
rect 1766 -2176 1767 -2086
rect 1773 -2087 1774 -2033
rect 1843 -2176 1844 -2086
rect 1850 -2087 1851 -2033
rect 1899 -2176 1900 -2086
rect 1906 -2087 1907 -2033
rect 1948 -2176 1949 -2086
rect 2326 -2087 2327 -2033
rect 2361 -2176 2362 -2086
rect 93 -2176 94 -2088
rect 1465 -2089 1466 -2033
rect 1479 -2089 1480 -2033
rect 1752 -2176 1753 -2088
rect 1780 -2089 1781 -2033
rect 1850 -2176 1851 -2088
rect 2004 -2089 2005 -2033
rect 2326 -2176 2327 -2088
rect 103 -2091 104 -2033
rect 1773 -2176 1774 -2090
rect 1780 -2176 1781 -2090
rect 1913 -2091 1914 -2033
rect 114 -2093 115 -2033
rect 793 -2176 794 -2092
rect 835 -2093 836 -2033
rect 919 -2176 920 -2092
rect 940 -2176 941 -2092
rect 982 -2093 983 -2033
rect 1080 -2176 1081 -2092
rect 1094 -2093 1095 -2033
rect 1143 -2093 1144 -2033
rect 1241 -2176 1242 -2092
rect 1311 -2093 1312 -2033
rect 1416 -2176 1417 -2092
rect 1451 -2093 1452 -2033
rect 1689 -2176 1690 -2092
rect 1703 -2093 1704 -2033
rect 1906 -2176 1907 -2092
rect 114 -2176 115 -2094
rect 352 -2095 353 -2033
rect 366 -2095 367 -2033
rect 464 -2176 465 -2094
rect 562 -2095 563 -2033
rect 618 -2176 619 -2094
rect 653 -2095 654 -2033
rect 954 -2176 955 -2094
rect 1094 -2176 1095 -2094
rect 1101 -2095 1102 -2033
rect 1136 -2095 1137 -2033
rect 1311 -2176 1312 -2094
rect 1332 -2095 1333 -2033
rect 1465 -2176 1466 -2094
rect 1500 -2095 1501 -2033
rect 1612 -2176 1613 -2094
rect 1626 -2095 1627 -2033
rect 1745 -2176 1746 -2094
rect 1794 -2095 1795 -2033
rect 2032 -2176 2033 -2094
rect 205 -2097 206 -2033
rect 352 -2176 353 -2096
rect 404 -2176 405 -2096
rect 968 -2176 969 -2096
rect 1010 -2097 1011 -2033
rect 1101 -2176 1102 -2096
rect 1136 -2176 1137 -2096
rect 1213 -2097 1214 -2033
rect 1325 -2097 1326 -2033
rect 1500 -2176 1501 -2096
rect 1528 -2097 1529 -2033
rect 1654 -2176 1655 -2096
rect 1703 -2176 1704 -2096
rect 1864 -2097 1865 -2033
rect 177 -2099 178 -2033
rect 205 -2176 206 -2098
rect 215 -2099 216 -2033
rect 1731 -2176 1732 -2098
rect 1801 -2099 1802 -2033
rect 1864 -2176 1865 -2098
rect 163 -2101 164 -2033
rect 177 -2176 178 -2100
rect 219 -2101 220 -2033
rect 1059 -2176 1060 -2100
rect 1143 -2176 1144 -2100
rect 1223 -2176 1224 -2100
rect 1262 -2101 1263 -2033
rect 1325 -2176 1326 -2100
rect 1332 -2176 1333 -2100
rect 2270 -2101 2271 -2033
rect 124 -2176 125 -2102
rect 163 -2176 164 -2102
rect 219 -2176 220 -2102
rect 1650 -2176 1651 -2102
rect 2221 -2103 2222 -2033
rect 2270 -2176 2271 -2102
rect 236 -2176 237 -2104
rect 681 -2105 682 -2033
rect 688 -2105 689 -2033
rect 1276 -2176 1277 -2104
rect 1353 -2105 1354 -2033
rect 1528 -2176 1529 -2104
rect 1535 -2105 1536 -2033
rect 1962 -2105 1963 -2033
rect 2179 -2105 2180 -2033
rect 2221 -2176 2222 -2104
rect 247 -2107 248 -2033
rect 1759 -2176 1760 -2106
rect 1927 -2107 1928 -2033
rect 1962 -2176 1963 -2106
rect 2165 -2107 2166 -2033
rect 2179 -2176 2180 -2106
rect 247 -2176 248 -2108
rect 289 -2109 290 -2033
rect 303 -2109 304 -2033
rect 506 -2176 507 -2108
rect 583 -2176 584 -2108
rect 611 -2109 612 -2033
rect 625 -2109 626 -2033
rect 681 -2176 682 -2108
rect 695 -2176 696 -2108
rect 957 -2109 958 -2033
rect 1010 -2176 1011 -2108
rect 1045 -2109 1046 -2033
rect 1164 -2109 1165 -2033
rect 2004 -2176 2005 -2108
rect 2123 -2109 2124 -2033
rect 2165 -2176 2166 -2108
rect 261 -2111 262 -2033
rect 317 -2176 318 -2110
rect 338 -2176 339 -2110
rect 1552 -2111 1553 -2033
rect 1563 -2111 1564 -2033
rect 1934 -2176 1935 -2110
rect 2067 -2111 2068 -2033
rect 2123 -2176 2124 -2110
rect 142 -2113 143 -2033
rect 261 -2176 262 -2112
rect 275 -2113 276 -2033
rect 688 -2176 689 -2112
rect 702 -2176 703 -2112
rect 1258 -2176 1259 -2112
rect 1262 -2176 1263 -2112
rect 1475 -2113 1476 -2033
rect 1538 -2113 1539 -2033
rect 1927 -2176 1928 -2112
rect 2011 -2113 2012 -2033
rect 2067 -2176 2068 -2112
rect 142 -2176 143 -2114
rect 1580 -2176 1581 -2114
rect 1584 -2115 1585 -2033
rect 1794 -2176 1795 -2114
rect 275 -2176 276 -2116
rect 548 -2117 549 -2033
rect 597 -2117 598 -2033
rect 611 -2176 612 -2116
rect 625 -2176 626 -2116
rect 856 -2117 857 -2033
rect 863 -2117 864 -2033
rect 1269 -2176 1270 -2116
rect 1367 -2117 1368 -2033
rect 1535 -2176 1536 -2116
rect 1542 -2117 1543 -2033
rect 1913 -2176 1914 -2116
rect 289 -2176 290 -2118
rect 387 -2119 388 -2033
rect 422 -2119 423 -2033
rect 1073 -2176 1074 -2118
rect 1164 -2176 1165 -2118
rect 1199 -2119 1200 -2033
rect 1213 -2176 1214 -2118
rect 1493 -2119 1494 -2033
rect 1549 -2119 1550 -2033
rect 2109 -2119 2110 -2033
rect 226 -2121 227 -2033
rect 387 -2176 388 -2120
rect 436 -2121 437 -2033
rect 597 -2176 598 -2120
rect 653 -2176 654 -2120
rect 2207 -2176 2208 -2120
rect 226 -2176 227 -2122
rect 646 -2123 647 -2033
rect 660 -2123 661 -2033
rect 1626 -2176 1627 -2122
rect 1636 -2123 1637 -2033
rect 2011 -2176 2012 -2122
rect 2060 -2123 2061 -2033
rect 2109 -2176 2110 -2122
rect 233 -2125 234 -2033
rect 422 -2176 423 -2124
rect 443 -2125 444 -2033
rect 646 -2176 647 -2124
rect 660 -2176 661 -2124
rect 975 -2176 976 -2124
rect 1188 -2125 1189 -2033
rect 1283 -2176 1284 -2124
rect 1339 -2125 1340 -2033
rect 1493 -2176 1494 -2124
rect 1549 -2176 1550 -2124
rect 1633 -2125 1634 -2033
rect 2060 -2176 2061 -2124
rect 2263 -2125 2264 -2033
rect 303 -2176 304 -2126
rect 555 -2127 556 -2033
rect 576 -2127 577 -2033
rect 863 -2176 864 -2126
rect 891 -2176 892 -2126
rect 1619 -2127 1620 -2033
rect 1633 -2176 1634 -2126
rect 1710 -2127 1711 -2033
rect 2235 -2127 2236 -2033
rect 2263 -2176 2264 -2126
rect 23 -2129 24 -2033
rect 1619 -2176 1620 -2128
rect 2193 -2129 2194 -2033
rect 2235 -2176 2236 -2128
rect 23 -2176 24 -2130
rect 131 -2131 132 -2033
rect 310 -2131 311 -2033
rect 310 -2176 311 -2130
rect 310 -2131 311 -2033
rect 310 -2176 311 -2130
rect 345 -2131 346 -2033
rect 366 -2176 367 -2130
rect 373 -2131 374 -2033
rect 548 -2176 549 -2130
rect 555 -2176 556 -2130
rect 870 -2131 871 -2033
rect 933 -2131 934 -2033
rect 1045 -2176 1046 -2130
rect 1188 -2176 1189 -2130
rect 1997 -2131 1998 -2033
rect 2151 -2131 2152 -2033
rect 2193 -2176 2194 -2130
rect 131 -2176 132 -2132
rect 212 -2176 213 -2132
rect 345 -2176 346 -2132
rect 401 -2133 402 -2033
rect 443 -2176 444 -2132
rect 996 -2133 997 -2033
rect 1199 -2176 1200 -2132
rect 2319 -2133 2320 -2033
rect 149 -2135 150 -2033
rect 870 -2176 871 -2134
rect 947 -2135 948 -2033
rect 982 -2176 983 -2134
rect 1248 -2135 1249 -2033
rect 1353 -2176 1354 -2134
rect 1381 -2135 1382 -2033
rect 1542 -2176 1543 -2134
rect 1563 -2176 1564 -2134
rect 1787 -2135 1788 -2033
rect 2151 -2176 2152 -2134
rect 2382 -2135 2383 -2033
rect 54 -2137 55 -2033
rect 149 -2176 150 -2136
rect 373 -2176 374 -2136
rect 1202 -2176 1203 -2136
rect 1381 -2176 1382 -2136
rect 1997 -2176 1998 -2136
rect 2144 -2137 2145 -2033
rect 2382 -2176 2383 -2136
rect 394 -2139 395 -2033
rect 436 -2176 437 -2138
rect 450 -2139 451 -2033
rect 632 -2139 633 -2033
rect 639 -2139 640 -2033
rect 996 -2176 997 -2138
rect 1157 -2139 1158 -2033
rect 1248 -2176 1249 -2138
rect 1570 -2139 1571 -2033
rect 1801 -2176 1802 -2138
rect 2088 -2139 2089 -2033
rect 2144 -2176 2145 -2138
rect 79 -2141 80 -2033
rect 394 -2176 395 -2140
rect 401 -2176 402 -2140
rect 408 -2141 409 -2033
rect 492 -2176 493 -2140
rect 562 -2176 563 -2140
rect 632 -2176 633 -2140
rect 1055 -2176 1056 -2140
rect 1125 -2141 1126 -2033
rect 1157 -2176 1158 -2140
rect 1458 -2141 1459 -2033
rect 1570 -2176 1571 -2140
rect 1577 -2141 1578 -2033
rect 1885 -2176 1886 -2140
rect 2039 -2141 2040 -2033
rect 2088 -2176 2089 -2140
rect 79 -2176 80 -2142
rect 534 -2143 535 -2033
rect 674 -2143 675 -2033
rect 856 -2176 857 -2142
rect 1052 -2143 1053 -2033
rect 1458 -2176 1459 -2142
rect 1584 -2176 1585 -2142
rect 1591 -2143 1592 -2033
rect 1598 -2176 1599 -2142
rect 1682 -2143 1683 -2033
rect 1787 -2176 1788 -2142
rect 2396 -2143 2397 -2033
rect 121 -2145 122 -2033
rect 450 -2176 451 -2144
rect 527 -2145 528 -2033
rect 576 -2176 577 -2144
rect 709 -2145 710 -2033
rect 779 -2176 780 -2144
rect 821 -2145 822 -2033
rect 1451 -2176 1452 -2144
rect 1556 -2145 1557 -2033
rect 1591 -2176 1592 -2144
rect 1605 -2176 1606 -2144
rect 1675 -2145 1676 -2033
rect 1682 -2176 1683 -2144
rect 1829 -2145 1830 -2033
rect 2396 -2176 2397 -2144
rect 2410 -2145 2411 -2033
rect 135 -2176 136 -2146
rect 527 -2176 528 -2146
rect 534 -2176 535 -2146
rect 1339 -2176 1340 -2146
rect 1507 -2147 1508 -2033
rect 1675 -2176 1676 -2146
rect 2102 -2147 2103 -2033
rect 2410 -2176 2411 -2146
rect 254 -2149 255 -2033
rect 674 -2176 675 -2148
rect 716 -2149 717 -2033
rect 786 -2176 787 -2148
rect 842 -2149 843 -2033
rect 947 -2176 948 -2148
rect 1052 -2176 1053 -2148
rect 1738 -2149 1739 -2033
rect 2053 -2149 2054 -2033
rect 2102 -2176 2103 -2148
rect 257 -2176 258 -2150
rect 821 -2176 822 -2150
rect 1185 -2151 1186 -2033
rect 2039 -2176 2040 -2150
rect 268 -2153 269 -2033
rect 639 -2176 640 -2152
rect 723 -2153 724 -2033
rect 835 -2176 836 -2152
rect 1185 -2176 1186 -2152
rect 2242 -2153 2243 -2033
rect 268 -2176 269 -2154
rect 1367 -2176 1368 -2154
rect 1374 -2155 1375 -2033
rect 1507 -2176 1508 -2154
rect 1556 -2176 1557 -2154
rect 1717 -2155 1718 -2033
rect 2200 -2155 2201 -2033
rect 2242 -2176 2243 -2154
rect 408 -2176 409 -2156
rect 415 -2157 416 -2033
rect 478 -2157 479 -2033
rect 709 -2176 710 -2156
rect 730 -2176 731 -2156
rect 877 -2157 878 -2033
rect 1230 -2176 1231 -2156
rect 1738 -2176 1739 -2156
rect 2158 -2157 2159 -2033
rect 2200 -2176 2201 -2156
rect 233 -2176 234 -2158
rect 478 -2176 479 -2158
rect 513 -2159 514 -2033
rect 723 -2176 724 -2158
rect 747 -2176 748 -2158
rect 933 -2176 934 -2158
rect 1255 -2176 1256 -2158
rect 1374 -2176 1375 -2158
rect 1647 -2159 1648 -2033
rect 2053 -2176 2054 -2158
rect 282 -2161 283 -2033
rect 513 -2176 514 -2160
rect 520 -2161 521 -2033
rect 716 -2176 717 -2160
rect 765 -2161 766 -2033
rect 1479 -2176 1480 -2160
rect 1647 -2176 1648 -2160
rect 2277 -2161 2278 -2033
rect 282 -2176 283 -2162
rect 324 -2163 325 -2033
rect 359 -2163 360 -2033
rect 520 -2176 521 -2162
rect 765 -2176 766 -2162
rect 772 -2163 773 -2033
rect 814 -2163 815 -2033
rect 842 -2176 843 -2162
rect 877 -2176 878 -2162
rect 1661 -2163 1662 -2033
rect 1668 -2163 1669 -2033
rect 1829 -2176 1830 -2162
rect 1892 -2163 1893 -2033
rect 2158 -2176 2159 -2162
rect 324 -2176 325 -2164
rect 429 -2165 430 -2033
rect 667 -2165 668 -2033
rect 814 -2176 815 -2164
rect 1346 -2165 1347 -2033
rect 1668 -2176 1669 -2164
rect 1717 -2176 1718 -2164
rect 1857 -2176 1858 -2164
rect 359 -2176 360 -2166
rect 485 -2167 486 -2033
rect 499 -2176 500 -2166
rect 667 -2176 668 -2166
rect 772 -2176 773 -2166
rect 912 -2167 913 -2033
rect 1346 -2176 1347 -2166
rect 1388 -2167 1389 -2033
rect 1496 -2167 1497 -2033
rect 2277 -2176 2278 -2166
rect 198 -2169 199 -2033
rect 485 -2176 486 -2168
rect 737 -2169 738 -2033
rect 1388 -2176 1389 -2168
rect 1514 -2169 1515 -2033
rect 1661 -2176 1662 -2168
rect 1836 -2169 1837 -2033
rect 1892 -2176 1893 -2168
rect 184 -2171 185 -2033
rect 198 -2176 199 -2170
rect 380 -2171 381 -2033
rect 415 -2176 416 -2170
rect 429 -2176 430 -2170
rect 744 -2176 745 -2170
rect 912 -2176 913 -2170
rect 1577 -2176 1578 -2170
rect 1836 -2176 1837 -2170
rect 2319 -2176 2320 -2170
rect 121 -2176 122 -2172
rect 380 -2176 381 -2172
rect 737 -2176 738 -2172
rect 1489 -2176 1490 -2172
rect 184 -2176 185 -2174
rect 243 -2176 244 -2174
rect 1220 -2176 1221 -2174
rect 1514 -2176 1515 -2174
rect 2 -2325 3 -2185
rect 674 -2186 675 -2184
rect 744 -2186 745 -2184
rect 1234 -2186 1235 -2184
rect 1258 -2186 1259 -2184
rect 2312 -2186 2313 -2184
rect 2343 -2325 2344 -2185
rect 2396 -2186 2397 -2184
rect 9 -2188 10 -2184
rect 51 -2188 52 -2184
rect 54 -2188 55 -2184
rect 1388 -2188 1389 -2184
rect 1398 -2325 1399 -2187
rect 1885 -2188 1886 -2184
rect 1937 -2325 1938 -2187
rect 2298 -2188 2299 -2184
rect 37 -2325 38 -2189
rect 996 -2190 997 -2184
rect 1038 -2190 1039 -2184
rect 1223 -2190 1224 -2184
rect 1227 -2190 1228 -2184
rect 2305 -2190 2306 -2184
rect 51 -2325 52 -2191
rect 1031 -2192 1032 -2184
rect 1080 -2192 1081 -2184
rect 1150 -2325 1151 -2191
rect 1157 -2192 1158 -2184
rect 1388 -2325 1389 -2191
rect 1405 -2192 1406 -2184
rect 1437 -2192 1438 -2184
rect 1489 -2192 1490 -2184
rect 2403 -2192 2404 -2184
rect 65 -2194 66 -2184
rect 1041 -2325 1042 -2193
rect 1080 -2325 1081 -2193
rect 1101 -2194 1102 -2184
rect 1115 -2194 1116 -2184
rect 1139 -2325 1140 -2193
rect 1143 -2194 1144 -2184
rect 1234 -2325 1235 -2193
rect 1293 -2325 1294 -2193
rect 1983 -2194 1984 -2184
rect 2151 -2194 2152 -2184
rect 2305 -2325 2306 -2193
rect 65 -2325 66 -2195
rect 1276 -2196 1277 -2184
rect 1304 -2196 1305 -2184
rect 1927 -2196 1928 -2184
rect 1969 -2196 1970 -2184
rect 2298 -2325 2299 -2195
rect 93 -2198 94 -2184
rect 1479 -2198 1480 -2184
rect 1496 -2325 1497 -2197
rect 1752 -2198 1753 -2184
rect 1780 -2198 1781 -2184
rect 1783 -2222 1784 -2197
rect 1836 -2325 1837 -2197
rect 1871 -2198 1872 -2184
rect 1885 -2325 1886 -2197
rect 1962 -2198 1963 -2184
rect 1969 -2325 1970 -2197
rect 2032 -2198 2033 -2184
rect 2151 -2325 2152 -2197
rect 2270 -2198 2271 -2184
rect 93 -2325 94 -2199
rect 1360 -2200 1361 -2184
rect 1367 -2200 1368 -2184
rect 2172 -2200 2173 -2184
rect 2228 -2200 2229 -2184
rect 2336 -2325 2337 -2199
rect 96 -2202 97 -2184
rect 926 -2202 927 -2184
rect 936 -2325 937 -2201
rect 1010 -2202 1011 -2184
rect 1031 -2325 1032 -2201
rect 1045 -2202 1046 -2184
rect 1094 -2202 1095 -2184
rect 1157 -2325 1158 -2201
rect 1192 -2202 1193 -2184
rect 1255 -2202 1256 -2184
rect 1304 -2325 1305 -2201
rect 1416 -2202 1417 -2184
rect 1437 -2325 1438 -2201
rect 1514 -2202 1515 -2184
rect 1521 -2202 1522 -2184
rect 1752 -2325 1753 -2201
rect 1780 -2325 1781 -2201
rect 1843 -2202 1844 -2184
rect 1860 -2202 1861 -2184
rect 2368 -2202 2369 -2184
rect 107 -2204 108 -2184
rect 128 -2204 129 -2184
rect 131 -2204 132 -2184
rect 257 -2204 258 -2184
rect 296 -2204 297 -2184
rect 656 -2204 657 -2184
rect 674 -2325 675 -2203
rect 1895 -2325 1896 -2203
rect 1927 -2325 1928 -2203
rect 1990 -2204 1991 -2184
rect 2032 -2325 2033 -2203
rect 2102 -2204 2103 -2184
rect 107 -2325 108 -2205
rect 506 -2206 507 -2184
rect 527 -2206 528 -2184
rect 1384 -2206 1385 -2184
rect 1416 -2325 1417 -2205
rect 1493 -2206 1494 -2184
rect 1521 -2325 1522 -2205
rect 1626 -2206 1627 -2184
rect 1629 -2325 1630 -2205
rect 2249 -2206 2250 -2184
rect 121 -2208 122 -2184
rect 1710 -2325 1711 -2207
rect 1843 -2325 1844 -2207
rect 1906 -2208 1907 -2184
rect 1962 -2325 1963 -2207
rect 2025 -2208 2026 -2184
rect 2060 -2208 2061 -2184
rect 2228 -2325 2229 -2207
rect 16 -2210 17 -2184
rect 121 -2325 122 -2209
rect 124 -2210 125 -2184
rect 387 -2210 388 -2184
rect 450 -2210 451 -2184
rect 495 -2210 496 -2184
rect 506 -2325 507 -2209
rect 779 -2210 780 -2184
rect 782 -2325 783 -2209
rect 992 -2325 993 -2209
rect 996 -2325 997 -2209
rect 1941 -2210 1942 -2184
rect 1983 -2325 1984 -2209
rect 2046 -2210 2047 -2184
rect 2060 -2325 2061 -2209
rect 2130 -2210 2131 -2184
rect 16 -2325 17 -2211
rect 86 -2212 87 -2184
rect 128 -2325 129 -2211
rect 1188 -2212 1189 -2184
rect 1192 -2325 1193 -2211
rect 1269 -2212 1270 -2184
rect 1332 -2212 1333 -2184
rect 1346 -2212 1347 -2184
rect 1367 -2325 1368 -2211
rect 1535 -2212 1536 -2184
rect 1545 -2325 1546 -2211
rect 2347 -2212 2348 -2184
rect 86 -2325 87 -2213
rect 625 -2214 626 -2184
rect 681 -2214 682 -2184
rect 744 -2325 745 -2213
rect 800 -2214 801 -2184
rect 1185 -2214 1186 -2184
rect 1202 -2214 1203 -2184
rect 1276 -2325 1277 -2213
rect 1283 -2214 1284 -2184
rect 1346 -2325 1347 -2213
rect 1381 -2214 1382 -2184
rect 1549 -2214 1550 -2184
rect 1580 -2214 1581 -2184
rect 2116 -2214 2117 -2184
rect 2130 -2325 2131 -2213
rect 2256 -2214 2257 -2184
rect 138 -2216 139 -2184
rect 2263 -2216 2264 -2184
rect 145 -2325 146 -2217
rect 856 -2218 857 -2184
rect 877 -2218 878 -2184
rect 1503 -2325 1504 -2217
rect 1517 -2325 1518 -2217
rect 2347 -2325 2348 -2217
rect 166 -2325 167 -2219
rect 2207 -2220 2208 -2184
rect 2256 -2325 2257 -2219
rect 2354 -2220 2355 -2184
rect 236 -2222 237 -2184
rect 940 -2222 941 -2184
rect 947 -2222 948 -2184
rect 947 -2325 948 -2221
rect 947 -2222 948 -2184
rect 947 -2325 948 -2221
rect 975 -2222 976 -2184
rect 1759 -2222 1760 -2184
rect 1906 -2325 1907 -2221
rect 1941 -2325 1942 -2221
rect 1997 -2222 1998 -2184
rect 2025 -2325 2026 -2221
rect 2088 -2222 2089 -2184
rect 2102 -2325 2103 -2221
rect 2200 -2222 2201 -2184
rect 2207 -2325 2208 -2221
rect 2340 -2222 2341 -2184
rect 243 -2325 244 -2223
rect 884 -2224 885 -2184
rect 912 -2224 913 -2184
rect 1010 -2325 1011 -2223
rect 1094 -2325 1095 -2223
rect 1171 -2224 1172 -2184
rect 1185 -2325 1186 -2223
rect 1262 -2224 1263 -2184
rect 1269 -2325 1270 -2223
rect 1290 -2224 1291 -2184
rect 1342 -2224 1343 -2184
rect 1430 -2224 1431 -2184
rect 1479 -2325 1480 -2223
rect 1787 -2224 1788 -2184
rect 1871 -2325 1872 -2223
rect 1948 -2224 1949 -2184
rect 1990 -2325 1991 -2223
rect 2053 -2224 2054 -2184
rect 2088 -2325 2089 -2223
rect 2165 -2224 2166 -2184
rect 2200 -2325 2201 -2223
rect 2333 -2224 2334 -2184
rect 156 -2226 157 -2184
rect 1171 -2325 1172 -2225
rect 1220 -2226 1221 -2184
rect 2284 -2226 2285 -2184
rect 40 -2228 41 -2184
rect 156 -2325 157 -2227
rect 250 -2325 251 -2227
rect 1220 -2325 1221 -2227
rect 1227 -2325 1228 -2227
rect 1451 -2228 1452 -2184
rect 1535 -2325 1536 -2227
rect 1668 -2228 1669 -2184
rect 1759 -2325 1760 -2227
rect 1815 -2228 1816 -2184
rect 1934 -2228 1935 -2184
rect 2165 -2325 2166 -2227
rect 2186 -2228 2187 -2184
rect 2284 -2325 2285 -2227
rect 289 -2230 290 -2184
rect 779 -2325 780 -2229
rect 821 -2230 822 -2184
rect 926 -2325 927 -2229
rect 940 -2325 941 -2229
rect 954 -2230 955 -2184
rect 975 -2325 976 -2229
rect 1979 -2325 1980 -2229
rect 1997 -2325 1998 -2229
rect 2067 -2230 2068 -2184
rect 2116 -2325 2117 -2229
rect 2221 -2230 2222 -2184
rect 289 -2325 290 -2231
rect 352 -2232 353 -2184
rect 359 -2232 360 -2184
rect 1055 -2232 1056 -2184
rect 1101 -2325 1102 -2231
rect 1129 -2232 1130 -2184
rect 1136 -2232 1137 -2184
rect 1332 -2325 1333 -2231
rect 1381 -2325 1382 -2231
rect 1465 -2232 1466 -2184
rect 1549 -2325 1550 -2231
rect 1591 -2232 1592 -2184
rect 1647 -2232 1648 -2184
rect 2263 -2325 2264 -2231
rect 261 -2234 262 -2184
rect 359 -2325 360 -2233
rect 457 -2234 458 -2184
rect 516 -2234 517 -2184
rect 527 -2325 528 -2233
rect 583 -2234 584 -2184
rect 590 -2234 591 -2184
rect 954 -2325 955 -2233
rect 978 -2234 979 -2184
rect 2312 -2325 2313 -2233
rect 100 -2236 101 -2184
rect 261 -2325 262 -2235
rect 296 -2325 297 -2235
rect 604 -2236 605 -2184
rect 618 -2236 619 -2184
rect 667 -2325 668 -2235
rect 681 -2325 682 -2235
rect 709 -2236 710 -2184
rect 726 -2325 727 -2235
rect 2172 -2325 2173 -2235
rect 2186 -2325 2187 -2235
rect 2417 -2236 2418 -2184
rect 100 -2325 101 -2237
rect 1017 -2238 1018 -2184
rect 1115 -2325 1116 -2237
rect 1696 -2238 1697 -2184
rect 1787 -2325 1788 -2237
rect 1850 -2238 1851 -2184
rect 1934 -2325 1935 -2237
rect 2179 -2238 2180 -2184
rect 2221 -2325 2222 -2237
rect 2319 -2238 2320 -2184
rect 170 -2240 171 -2184
rect 457 -2325 458 -2239
rect 492 -2240 493 -2184
rect 1073 -2240 1074 -2184
rect 1129 -2325 1130 -2239
rect 1164 -2240 1165 -2184
rect 1248 -2240 1249 -2184
rect 1360 -2325 1361 -2239
rect 1423 -2240 1424 -2184
rect 1451 -2325 1452 -2239
rect 1465 -2325 1466 -2239
rect 1570 -2240 1571 -2184
rect 1591 -2325 1592 -2239
rect 1689 -2240 1690 -2184
rect 1703 -2240 1704 -2184
rect 1850 -2325 1851 -2239
rect 1948 -2325 1949 -2239
rect 2004 -2240 2005 -2184
rect 2046 -2325 2047 -2239
rect 2333 -2325 2334 -2239
rect 79 -2242 80 -2184
rect 492 -2325 493 -2241
rect 555 -2242 556 -2184
rect 1230 -2242 1231 -2184
rect 1248 -2325 1249 -2241
rect 2270 -2325 2271 -2241
rect 79 -2325 80 -2243
rect 639 -2244 640 -2184
rect 653 -2325 654 -2243
rect 1136 -2325 1137 -2243
rect 1143 -2325 1144 -2243
rect 1206 -2244 1207 -2184
rect 1255 -2325 1256 -2243
rect 1374 -2244 1375 -2184
rect 1423 -2325 1424 -2243
rect 1514 -2325 1515 -2243
rect 1570 -2325 1571 -2243
rect 1661 -2244 1662 -2184
rect 1682 -2244 1683 -2184
rect 1815 -2325 1816 -2243
rect 1857 -2244 1858 -2184
rect 2004 -2325 2005 -2243
rect 2053 -2325 2054 -2243
rect 2123 -2244 2124 -2184
rect 2179 -2325 2180 -2243
rect 2291 -2244 2292 -2184
rect 170 -2325 171 -2245
rect 177 -2246 178 -2184
rect 338 -2246 339 -2184
rect 450 -2325 451 -2245
rect 576 -2246 577 -2184
rect 618 -2325 619 -2245
rect 621 -2325 622 -2245
rect 1577 -2325 1578 -2245
rect 1605 -2246 1606 -2184
rect 1689 -2325 1690 -2245
rect 1703 -2325 1704 -2245
rect 1766 -2246 1767 -2184
rect 1857 -2325 1858 -2245
rect 1920 -2246 1921 -2184
rect 2067 -2325 2068 -2245
rect 2137 -2246 2138 -2184
rect 177 -2325 178 -2247
rect 1685 -2325 1686 -2247
rect 1766 -2325 1767 -2247
rect 1822 -2248 1823 -2184
rect 2123 -2325 2124 -2247
rect 2235 -2248 2236 -2184
rect 317 -2250 318 -2184
rect 338 -2325 339 -2249
rect 352 -2325 353 -2249
rect 366 -2250 367 -2184
rect 394 -2250 395 -2184
rect 555 -2325 556 -2249
rect 583 -2325 584 -2249
rect 597 -2250 598 -2184
rect 604 -2325 605 -2249
rect 695 -2250 696 -2184
rect 709 -2325 710 -2249
rect 919 -2250 920 -2184
rect 978 -2325 979 -2249
rect 2291 -2325 2292 -2249
rect 275 -2252 276 -2184
rect 597 -2325 598 -2251
rect 639 -2325 640 -2251
rect 891 -2252 892 -2184
rect 912 -2325 913 -2251
rect 989 -2252 990 -2184
rect 1073 -2325 1074 -2251
rect 1122 -2252 1123 -2184
rect 1164 -2325 1165 -2251
rect 1241 -2252 1242 -2184
rect 1262 -2325 1263 -2251
rect 1395 -2252 1396 -2184
rect 1430 -2325 1431 -2251
rect 1500 -2252 1501 -2184
rect 1605 -2325 1606 -2251
rect 1640 -2252 1641 -2184
rect 1647 -2325 1648 -2251
rect 1808 -2252 1809 -2184
rect 2074 -2252 2075 -2184
rect 2235 -2325 2236 -2251
rect 275 -2325 276 -2253
rect 625 -2325 626 -2253
rect 688 -2254 689 -2184
rect 821 -2325 822 -2253
rect 828 -2254 829 -2184
rect 884 -2325 885 -2253
rect 982 -2254 983 -2184
rect 1045 -2325 1046 -2253
rect 1087 -2254 1088 -2184
rect 1122 -2325 1123 -2253
rect 1178 -2254 1179 -2184
rect 1241 -2325 1242 -2253
rect 1283 -2325 1284 -2253
rect 1318 -2254 1319 -2184
rect 1339 -2254 1340 -2184
rect 1822 -2325 1823 -2253
rect 2018 -2254 2019 -2184
rect 2074 -2325 2075 -2253
rect 310 -2256 311 -2184
rect 317 -2325 318 -2255
rect 324 -2256 325 -2184
rect 394 -2325 395 -2255
rect 443 -2256 444 -2184
rect 891 -2325 892 -2255
rect 961 -2256 962 -2184
rect 1087 -2325 1088 -2255
rect 1178 -2325 1179 -2255
rect 1444 -2256 1445 -2184
rect 1486 -2256 1487 -2184
rect 1920 -2325 1921 -2255
rect 2018 -2325 2019 -2255
rect 2361 -2256 2362 -2184
rect 114 -2258 115 -2184
rect 324 -2325 325 -2257
rect 366 -2325 367 -2257
rect 663 -2325 664 -2257
rect 695 -2325 696 -2257
rect 1307 -2258 1308 -2184
rect 1318 -2325 1319 -2257
rect 2410 -2258 2411 -2184
rect 114 -2325 115 -2259
rect 226 -2260 227 -2184
rect 310 -2325 311 -2259
rect 541 -2260 542 -2184
rect 590 -2325 591 -2259
rect 870 -2260 871 -2184
rect 933 -2260 934 -2184
rect 961 -2325 962 -2259
rect 989 -2325 990 -2259
rect 2424 -2260 2425 -2184
rect 163 -2262 164 -2184
rect 226 -2325 227 -2261
rect 380 -2262 381 -2184
rect 688 -2325 689 -2261
rect 751 -2262 752 -2184
rect 1017 -2325 1018 -2261
rect 1206 -2325 1207 -2261
rect 1297 -2262 1298 -2184
rect 1339 -2325 1340 -2261
rect 1458 -2262 1459 -2184
rect 1472 -2262 1473 -2184
rect 1486 -2325 1487 -2261
rect 1500 -2325 1501 -2261
rect 2382 -2262 2383 -2184
rect 163 -2325 164 -2263
rect 2249 -2325 2250 -2263
rect 380 -2325 381 -2265
rect 835 -2266 836 -2184
rect 856 -2325 857 -2265
rect 1976 -2266 1977 -2184
rect 443 -2325 444 -2267
rect 471 -2268 472 -2184
rect 478 -2268 479 -2184
rect 576 -2325 577 -2267
rect 593 -2325 594 -2267
rect 2039 -2268 2040 -2184
rect 142 -2270 143 -2184
rect 471 -2325 472 -2269
rect 478 -2325 479 -2269
rect 919 -2325 920 -2269
rect 1290 -2325 1291 -2269
rect 1913 -2270 1914 -2184
rect 2039 -2325 2040 -2269
rect 2109 -2270 2110 -2184
rect 142 -2325 143 -2271
rect 254 -2325 255 -2271
rect 513 -2272 514 -2184
rect 870 -2325 871 -2271
rect 1297 -2325 1298 -2271
rect 1353 -2272 1354 -2184
rect 1370 -2272 1371 -2184
rect 1458 -2325 1459 -2271
rect 1472 -2325 1473 -2271
rect 1955 -2272 1956 -2184
rect 2109 -2325 2110 -2271
rect 2214 -2272 2215 -2184
rect 513 -2325 514 -2273
rect 534 -2274 535 -2184
rect 541 -2325 542 -2273
rect 548 -2274 549 -2184
rect 737 -2274 738 -2184
rect 751 -2325 752 -2273
rect 758 -2274 759 -2184
rect 1668 -2325 1669 -2273
rect 1808 -2325 1809 -2273
rect 2011 -2274 2012 -2184
rect 2095 -2274 2096 -2184
rect 2214 -2325 2215 -2273
rect 422 -2276 423 -2184
rect 534 -2325 535 -2275
rect 548 -2325 549 -2275
rect 716 -2276 717 -2184
rect 758 -2325 759 -2275
rect 863 -2276 864 -2184
rect 1353 -2325 1354 -2275
rect 1528 -2276 1529 -2184
rect 1563 -2276 1564 -2184
rect 1955 -2325 1956 -2275
rect 2011 -2325 2012 -2275
rect 2081 -2276 2082 -2184
rect 2095 -2325 2096 -2275
rect 2193 -2276 2194 -2184
rect 184 -2278 185 -2184
rect 716 -2325 717 -2277
rect 765 -2278 766 -2184
rect 877 -2325 878 -2277
rect 1059 -2278 1060 -2184
rect 1528 -2325 1529 -2277
rect 1563 -2325 1564 -2277
rect 1654 -2278 1655 -2184
rect 1661 -2325 1662 -2277
rect 1738 -2278 1739 -2184
rect 1892 -2278 1893 -2184
rect 1913 -2325 1914 -2277
rect 2081 -2325 2082 -2277
rect 2158 -2278 2159 -2184
rect 149 -2280 150 -2184
rect 184 -2325 185 -2279
rect 219 -2280 220 -2184
rect 422 -2325 423 -2279
rect 485 -2280 486 -2184
rect 737 -2325 738 -2279
rect 772 -2280 773 -2184
rect 800 -2325 801 -2279
rect 814 -2280 815 -2184
rect 863 -2325 864 -2279
rect 1059 -2325 1060 -2279
rect 1335 -2280 1336 -2184
rect 1374 -2325 1375 -2279
rect 1542 -2280 1543 -2184
rect 1619 -2280 1620 -2184
rect 1696 -2325 1697 -2279
rect 1738 -2325 1739 -2279
rect 1794 -2280 1795 -2184
rect 135 -2282 136 -2184
rect 149 -2325 150 -2281
rect 191 -2282 192 -2184
rect 219 -2325 220 -2281
rect 373 -2282 374 -2184
rect 765 -2325 766 -2281
rect 786 -2282 787 -2184
rect 2319 -2325 2320 -2281
rect 135 -2325 136 -2283
rect 569 -2284 570 -2184
rect 611 -2284 612 -2184
rect 814 -2325 815 -2283
rect 828 -2325 829 -2283
rect 842 -2284 843 -2184
rect 859 -2325 860 -2283
rect 2137 -2325 2138 -2283
rect 191 -2325 192 -2285
rect 1066 -2286 1067 -2184
rect 1321 -2325 1322 -2285
rect 2193 -2325 2194 -2285
rect 373 -2325 374 -2287
rect 520 -2288 521 -2184
rect 569 -2325 570 -2287
rect 723 -2288 724 -2184
rect 786 -2325 787 -2287
rect 1003 -2288 1004 -2184
rect 1066 -2325 1067 -2287
rect 1108 -2288 1109 -2184
rect 1395 -2325 1396 -2287
rect 1976 -2325 1977 -2287
rect 415 -2290 416 -2184
rect 520 -2325 521 -2289
rect 646 -2290 647 -2184
rect 772 -2325 773 -2289
rect 807 -2290 808 -2184
rect 842 -2325 843 -2289
rect 968 -2290 969 -2184
rect 1542 -2325 1543 -2289
rect 1619 -2325 1620 -2289
rect 1717 -2290 1718 -2184
rect 1794 -2325 1795 -2289
rect 1864 -2290 1865 -2184
rect 331 -2292 332 -2184
rect 415 -2325 416 -2291
rect 436 -2292 437 -2184
rect 485 -2325 486 -2291
rect 499 -2292 500 -2184
rect 611 -2325 612 -2291
rect 646 -2325 647 -2291
rect 660 -2292 661 -2184
rect 723 -2325 724 -2291
rect 982 -2325 983 -2291
rect 1052 -2292 1053 -2184
rect 1108 -2325 1109 -2291
rect 1402 -2292 1403 -2184
rect 2158 -2325 2159 -2291
rect 233 -2294 234 -2184
rect 499 -2325 500 -2293
rect 562 -2294 563 -2184
rect 1402 -2325 1403 -2293
rect 1409 -2294 1410 -2184
rect 1864 -2325 1865 -2293
rect 233 -2325 234 -2295
rect 705 -2325 706 -2295
rect 730 -2296 731 -2184
rect 1052 -2325 1053 -2295
rect 1409 -2325 1410 -2295
rect 1626 -2325 1627 -2295
rect 1633 -2296 1634 -2184
rect 1717 -2325 1718 -2295
rect 268 -2298 269 -2184
rect 436 -2325 437 -2297
rect 730 -2325 731 -2297
rect 898 -2298 899 -2184
rect 905 -2298 906 -2184
rect 968 -2325 969 -2297
rect 1444 -2325 1445 -2297
rect 1584 -2298 1585 -2184
rect 1633 -2325 1634 -2297
rect 1724 -2298 1725 -2184
rect 205 -2300 206 -2184
rect 898 -2325 899 -2299
rect 905 -2325 906 -2299
rect 1325 -2300 1326 -2184
rect 1584 -2325 1585 -2299
rect 1675 -2300 1676 -2184
rect 44 -2302 45 -2184
rect 205 -2325 206 -2301
rect 212 -2302 213 -2184
rect 268 -2325 269 -2301
rect 331 -2325 332 -2301
rect 345 -2302 346 -2184
rect 429 -2302 430 -2184
rect 562 -2325 563 -2301
rect 747 -2302 748 -2184
rect 1003 -2325 1004 -2301
rect 1024 -2302 1025 -2184
rect 1724 -2325 1725 -2301
rect 44 -2325 45 -2303
rect 58 -2304 59 -2184
rect 72 -2304 73 -2184
rect 1024 -2325 1025 -2303
rect 1325 -2325 1326 -2303
rect 1612 -2304 1613 -2184
rect 1640 -2325 1641 -2303
rect 1731 -2304 1732 -2184
rect 23 -2306 24 -2184
rect 58 -2325 59 -2305
rect 72 -2325 73 -2305
rect 401 -2306 402 -2184
rect 807 -2325 808 -2305
rect 849 -2306 850 -2184
rect 1507 -2306 1508 -2184
rect 1612 -2325 1613 -2305
rect 1650 -2306 1651 -2184
rect 2326 -2306 2327 -2184
rect 23 -2325 24 -2307
rect 198 -2308 199 -2184
rect 212 -2325 213 -2307
rect 247 -2308 248 -2184
rect 282 -2308 283 -2184
rect 345 -2325 346 -2307
rect 401 -2325 402 -2307
rect 464 -2308 465 -2184
rect 835 -2325 836 -2307
rect 1213 -2308 1214 -2184
rect 1507 -2325 1508 -2307
rect 1556 -2308 1557 -2184
rect 1675 -2325 1676 -2307
rect 1745 -2308 1746 -2184
rect 2277 -2308 2278 -2184
rect 2326 -2325 2327 -2307
rect 198 -2325 199 -2309
rect 670 -2310 671 -2184
rect 793 -2310 794 -2184
rect 1213 -2325 1214 -2309
rect 1556 -2325 1557 -2309
rect 1598 -2310 1599 -2184
rect 1731 -2325 1732 -2309
rect 2144 -2310 2145 -2184
rect 2277 -2325 2278 -2309
rect 2389 -2310 2390 -2184
rect 247 -2325 248 -2311
rect 429 -2325 430 -2311
rect 464 -2325 465 -2311
rect 632 -2312 633 -2184
rect 789 -2312 790 -2184
rect 1598 -2325 1599 -2311
rect 1745 -2325 1746 -2311
rect 1801 -2312 1802 -2184
rect 2144 -2325 2145 -2311
rect 2242 -2312 2243 -2184
rect 282 -2325 283 -2313
rect 303 -2314 304 -2184
rect 387 -2325 388 -2313
rect 670 -2325 671 -2313
rect 793 -2325 794 -2313
rect 1493 -2325 1494 -2313
rect 1801 -2325 1802 -2313
rect 1878 -2314 1879 -2184
rect 2242 -2325 2243 -2313
rect 2375 -2314 2376 -2184
rect 303 -2325 304 -2315
rect 408 -2316 409 -2184
rect 632 -2325 633 -2315
rect 702 -2316 703 -2184
rect 849 -2325 850 -2315
rect 1311 -2316 1312 -2184
rect 1773 -2316 1774 -2184
rect 1878 -2325 1879 -2315
rect 30 -2318 31 -2184
rect 408 -2325 409 -2317
rect 660 -2325 661 -2317
rect 1311 -2325 1312 -2317
rect 1773 -2325 1774 -2317
rect 1829 -2318 1830 -2184
rect 702 -2325 703 -2319
rect 1654 -2325 1655 -2319
rect 1829 -2325 1830 -2319
rect 1899 -2320 1900 -2184
rect 1199 -2322 1200 -2184
rect 1899 -2325 1900 -2321
rect 33 -2325 34 -2323
rect 1199 -2325 1200 -2323
rect 5 -2498 6 -2334
rect 65 -2335 66 -2333
rect 163 -2335 164 -2333
rect 1024 -2335 1025 -2333
rect 1038 -2335 1039 -2333
rect 1360 -2335 1361 -2333
rect 1363 -2498 1364 -2334
rect 2221 -2335 2222 -2333
rect 2326 -2335 2327 -2333
rect 2343 -2335 2344 -2333
rect 9 -2498 10 -2336
rect 873 -2498 874 -2336
rect 905 -2337 906 -2333
rect 1248 -2337 1249 -2333
rect 1272 -2498 1273 -2336
rect 2074 -2337 2075 -2333
rect 2165 -2337 2166 -2333
rect 2333 -2337 2334 -2333
rect 23 -2339 24 -2333
rect 145 -2339 146 -2333
rect 170 -2339 171 -2333
rect 173 -2361 174 -2338
rect 226 -2339 227 -2333
rect 593 -2339 594 -2333
rect 597 -2339 598 -2333
rect 726 -2339 727 -2333
rect 782 -2339 783 -2333
rect 1535 -2339 1536 -2333
rect 1542 -2339 1543 -2333
rect 1878 -2339 1879 -2333
rect 1892 -2498 1893 -2338
rect 1948 -2339 1949 -2333
rect 1976 -2498 1977 -2338
rect 2039 -2339 2040 -2333
rect 2165 -2498 2166 -2338
rect 2193 -2339 2194 -2333
rect 2221 -2498 2222 -2338
rect 2242 -2339 2243 -2333
rect 16 -2341 17 -2333
rect 226 -2498 227 -2340
rect 240 -2498 241 -2340
rect 607 -2498 608 -2340
rect 618 -2341 619 -2333
rect 1318 -2341 1319 -2333
rect 1374 -2341 1375 -2333
rect 1395 -2498 1396 -2340
rect 1398 -2341 1399 -2333
rect 1409 -2341 1410 -2333
rect 1493 -2341 1494 -2333
rect 2235 -2341 2236 -2333
rect 2242 -2498 2243 -2340
rect 2291 -2341 2292 -2333
rect 16 -2498 17 -2342
rect 37 -2343 38 -2333
rect 51 -2343 52 -2333
rect 1024 -2498 1025 -2342
rect 1041 -2343 1042 -2333
rect 1493 -2498 1494 -2342
rect 1517 -2343 1518 -2333
rect 1906 -2343 1907 -2333
rect 1934 -2343 1935 -2333
rect 2284 -2343 2285 -2333
rect 30 -2345 31 -2333
rect 1080 -2345 1081 -2333
rect 1108 -2345 1109 -2333
rect 1979 -2345 1980 -2333
rect 2039 -2498 2040 -2344
rect 2088 -2345 2089 -2333
rect 2186 -2345 2187 -2333
rect 2291 -2498 2292 -2344
rect 33 -2347 34 -2333
rect 44 -2347 45 -2333
rect 51 -2498 52 -2346
rect 1577 -2347 1578 -2333
rect 1580 -2498 1581 -2346
rect 2256 -2347 2257 -2333
rect 44 -2498 45 -2348
rect 114 -2349 115 -2333
rect 170 -2498 171 -2348
rect 243 -2349 244 -2333
rect 506 -2349 507 -2333
rect 569 -2349 570 -2333
rect 618 -2498 619 -2348
rect 625 -2498 626 -2348
rect 891 -2349 892 -2333
rect 905 -2498 906 -2348
rect 940 -2349 941 -2333
rect 954 -2349 955 -2333
rect 1321 -2349 1322 -2333
rect 1377 -2498 1378 -2348
rect 1451 -2349 1452 -2333
rect 1542 -2498 1543 -2348
rect 1598 -2349 1599 -2333
rect 1682 -2349 1683 -2333
rect 2228 -2349 2229 -2333
rect 2235 -2498 2236 -2348
rect 2277 -2349 2278 -2333
rect 65 -2498 66 -2350
rect 275 -2351 276 -2333
rect 282 -2351 283 -2333
rect 1076 -2498 1077 -2350
rect 1080 -2498 1081 -2350
rect 1612 -2351 1613 -2333
rect 1682 -2498 1683 -2350
rect 1745 -2351 1746 -2333
rect 1850 -2351 1851 -2333
rect 1853 -2351 1854 -2333
rect 1878 -2498 1879 -2350
rect 2102 -2351 2103 -2333
rect 2179 -2351 2180 -2333
rect 2186 -2498 2187 -2350
rect 2193 -2498 2194 -2350
rect 2207 -2351 2208 -2333
rect 2228 -2498 2229 -2350
rect 2263 -2351 2264 -2333
rect 114 -2498 115 -2352
rect 261 -2353 262 -2333
rect 275 -2498 276 -2352
rect 387 -2353 388 -2333
rect 408 -2353 409 -2333
rect 765 -2498 766 -2352
rect 775 -2498 776 -2352
rect 940 -2498 941 -2352
rect 978 -2353 979 -2333
rect 1213 -2353 1214 -2333
rect 1248 -2498 1249 -2352
rect 1262 -2353 1263 -2333
rect 1276 -2353 1277 -2333
rect 1356 -2498 1357 -2352
rect 1451 -2498 1452 -2352
rect 1528 -2353 1529 -2333
rect 1685 -2353 1686 -2333
rect 2158 -2353 2159 -2333
rect 2207 -2498 2208 -2352
rect 2280 -2498 2281 -2352
rect 166 -2355 167 -2333
rect 2179 -2498 2180 -2354
rect 2256 -2498 2257 -2354
rect 2312 -2355 2313 -2333
rect 247 -2357 248 -2333
rect 842 -2357 843 -2333
rect 859 -2357 860 -2333
rect 1612 -2498 1613 -2356
rect 1745 -2498 1746 -2356
rect 1773 -2357 1774 -2333
rect 1850 -2498 1851 -2356
rect 1885 -2357 1886 -2333
rect 1895 -2357 1896 -2333
rect 2214 -2357 2215 -2333
rect 2263 -2498 2264 -2356
rect 2319 -2357 2320 -2333
rect 247 -2498 248 -2358
rect 478 -2359 479 -2333
rect 481 -2498 482 -2358
rect 1629 -2359 1630 -2333
rect 1773 -2498 1774 -2358
rect 1787 -2359 1788 -2333
rect 1885 -2498 1886 -2358
rect 1941 -2359 1942 -2333
rect 1948 -2498 1949 -2358
rect 2116 -2359 2117 -2333
rect 254 -2361 255 -2333
rect 254 -2498 255 -2360
rect 254 -2361 255 -2333
rect 254 -2498 255 -2360
rect 261 -2498 262 -2360
rect 401 -2361 402 -2333
rect 408 -2498 409 -2360
rect 485 -2361 486 -2333
rect 492 -2361 493 -2333
rect 506 -2498 507 -2360
rect 527 -2361 528 -2333
rect 569 -2498 570 -2360
rect 576 -2361 577 -2333
rect 779 -2498 780 -2360
rect 786 -2361 787 -2333
rect 954 -2498 955 -2360
rect 982 -2361 983 -2333
rect 1038 -2498 1039 -2360
rect 1055 -2498 1056 -2360
rect 1486 -2361 1487 -2333
rect 1528 -2498 1529 -2360
rect 1591 -2361 1592 -2333
rect 1787 -2498 1788 -2360
rect 1843 -2361 1844 -2333
rect 1853 -2498 1854 -2360
rect 1941 -2498 1942 -2360
rect 2011 -2361 2012 -2333
rect 2116 -2498 2117 -2360
rect 282 -2498 283 -2362
rect 835 -2363 836 -2333
rect 842 -2498 843 -2362
rect 912 -2363 913 -2333
rect 919 -2363 920 -2333
rect 1696 -2363 1697 -2333
rect 1843 -2498 1844 -2362
rect 1857 -2363 1858 -2333
rect 1906 -2498 1907 -2362
rect 1927 -2363 1928 -2333
rect 1934 -2498 1935 -2362
rect 1997 -2363 1998 -2333
rect 2011 -2498 2012 -2362
rect 2067 -2363 2068 -2333
rect 2088 -2498 2089 -2362
rect 2305 -2363 2306 -2333
rect 296 -2365 297 -2333
rect 723 -2365 724 -2333
rect 730 -2365 731 -2333
rect 1409 -2498 1410 -2364
rect 1486 -2498 1487 -2364
rect 1570 -2365 1571 -2333
rect 1591 -2498 1592 -2364
rect 1822 -2365 1823 -2333
rect 1836 -2365 1837 -2333
rect 1857 -2498 1858 -2364
rect 1927 -2498 1928 -2364
rect 1990 -2365 1991 -2333
rect 1997 -2498 1998 -2364
rect 2060 -2365 2061 -2333
rect 2102 -2498 2103 -2364
rect 2130 -2365 2131 -2333
rect 2305 -2498 2306 -2364
rect 2347 -2365 2348 -2333
rect 191 -2367 192 -2333
rect 723 -2498 724 -2366
rect 730 -2498 731 -2366
rect 793 -2367 794 -2333
rect 796 -2498 797 -2366
rect 1668 -2367 1669 -2333
rect 1678 -2498 1679 -2366
rect 1696 -2498 1697 -2366
rect 1836 -2498 1837 -2366
rect 1983 -2367 1984 -2333
rect 1990 -2498 1991 -2366
rect 2123 -2367 2124 -2333
rect 72 -2369 73 -2333
rect 191 -2498 192 -2368
rect 296 -2498 297 -2368
rect 1052 -2369 1053 -2333
rect 1108 -2498 1109 -2368
rect 1150 -2369 1151 -2333
rect 1262 -2498 1263 -2368
rect 1304 -2369 1305 -2333
rect 1318 -2498 1319 -2368
rect 1381 -2369 1382 -2333
rect 1668 -2498 1669 -2368
rect 1738 -2369 1739 -2333
rect 1983 -2498 1984 -2368
rect 2053 -2369 2054 -2333
rect 2060 -2498 2061 -2368
rect 2109 -2369 2110 -2333
rect 2123 -2498 2124 -2368
rect 2137 -2369 2138 -2333
rect 310 -2371 311 -2333
rect 429 -2498 430 -2370
rect 457 -2371 458 -2333
rect 856 -2371 857 -2333
rect 859 -2498 860 -2370
rect 1332 -2371 1333 -2333
rect 1381 -2498 1382 -2370
rect 1437 -2371 1438 -2333
rect 1738 -2498 1739 -2370
rect 1766 -2371 1767 -2333
rect 1969 -2371 1970 -2333
rect 2109 -2498 2110 -2370
rect 2137 -2498 2138 -2370
rect 2151 -2371 2152 -2333
rect 268 -2373 269 -2333
rect 310 -2498 311 -2372
rect 317 -2373 318 -2333
rect 317 -2498 318 -2372
rect 317 -2373 318 -2333
rect 317 -2498 318 -2372
rect 387 -2498 388 -2372
rect 856 -2498 857 -2372
rect 863 -2373 864 -2333
rect 982 -2498 983 -2372
rect 1052 -2498 1053 -2372
rect 2074 -2498 2075 -2372
rect 2151 -2498 2152 -2372
rect 2172 -2373 2173 -2333
rect 401 -2498 402 -2374
rect 681 -2375 682 -2333
rect 716 -2375 717 -2333
rect 2067 -2498 2068 -2374
rect 2172 -2498 2173 -2374
rect 2200 -2375 2201 -2333
rect 37 -2498 38 -2376
rect 2200 -2498 2201 -2376
rect 100 -2379 101 -2333
rect 716 -2498 717 -2378
rect 786 -2498 787 -2378
rect 1164 -2379 1165 -2333
rect 1227 -2379 1228 -2333
rect 1304 -2498 1305 -2378
rect 1437 -2498 1438 -2378
rect 1444 -2379 1445 -2333
rect 1766 -2498 1767 -2378
rect 1829 -2379 1830 -2333
rect 2018 -2379 2019 -2333
rect 2214 -2498 2215 -2378
rect 100 -2498 101 -2380
rect 961 -2381 962 -2333
rect 1087 -2381 1088 -2333
rect 1164 -2498 1165 -2380
rect 1227 -2498 1228 -2380
rect 1255 -2381 1256 -2333
rect 1276 -2498 1277 -2380
rect 1545 -2381 1546 -2333
rect 1647 -2381 1648 -2333
rect 1829 -2498 1830 -2380
rect 2046 -2381 2047 -2333
rect 2284 -2498 2285 -2380
rect 422 -2383 423 -2333
rect 768 -2383 769 -2333
rect 821 -2383 822 -2333
rect 978 -2498 979 -2382
rect 1087 -2498 1088 -2382
rect 1129 -2383 1130 -2333
rect 1136 -2383 1137 -2333
rect 1297 -2383 1298 -2333
rect 1444 -2498 1445 -2382
rect 1479 -2383 1480 -2333
rect 1549 -2383 1550 -2333
rect 1647 -2498 1648 -2382
rect 1801 -2383 1802 -2333
rect 1969 -2498 1970 -2382
rect 2053 -2498 2054 -2382
rect 2095 -2383 2096 -2333
rect 110 -2498 111 -2384
rect 1136 -2498 1137 -2384
rect 1150 -2498 1151 -2384
rect 1185 -2385 1186 -2333
rect 1293 -2385 1294 -2333
rect 1752 -2385 1753 -2333
rect 1899 -2385 1900 -2333
rect 2095 -2498 2096 -2384
rect 324 -2387 325 -2333
rect 422 -2498 423 -2386
rect 457 -2498 458 -2386
rect 646 -2387 647 -2333
rect 660 -2387 661 -2333
rect 758 -2387 759 -2333
rect 821 -2498 822 -2386
rect 877 -2387 878 -2333
rect 884 -2387 885 -2333
rect 891 -2498 892 -2386
rect 912 -2498 913 -2386
rect 1335 -2498 1336 -2386
rect 1479 -2498 1480 -2386
rect 1703 -2387 1704 -2333
rect 1752 -2498 1753 -2386
rect 1780 -2387 1781 -2333
rect 1801 -2498 1802 -2386
rect 1899 -2498 1900 -2386
rect 324 -2498 325 -2388
rect 394 -2389 395 -2333
rect 464 -2389 465 -2333
rect 485 -2498 486 -2388
rect 492 -2498 493 -2388
rect 1311 -2389 1312 -2333
rect 1465 -2389 1466 -2333
rect 1780 -2498 1781 -2388
rect 303 -2391 304 -2333
rect 394 -2498 395 -2390
rect 464 -2498 465 -2390
rect 1017 -2391 1018 -2333
rect 1115 -2391 1116 -2333
rect 1535 -2498 1536 -2390
rect 1703 -2498 1704 -2390
rect 1717 -2391 1718 -2333
rect 303 -2498 304 -2392
rect 331 -2393 332 -2333
rect 520 -2393 521 -2333
rect 681 -2498 682 -2392
rect 702 -2393 703 -2333
rect 1185 -2498 1186 -2392
rect 1311 -2498 1312 -2392
rect 1339 -2393 1340 -2333
rect 1710 -2393 1711 -2333
rect 1717 -2498 1718 -2392
rect 331 -2498 332 -2394
rect 352 -2395 353 -2333
rect 380 -2395 381 -2333
rect 520 -2498 521 -2394
rect 527 -2498 528 -2394
rect 1251 -2395 1252 -2333
rect 1339 -2498 1340 -2394
rect 1388 -2395 1389 -2333
rect 1598 -2498 1599 -2394
rect 1710 -2498 1711 -2394
rect 345 -2397 346 -2333
rect 352 -2498 353 -2396
rect 380 -2498 381 -2396
rect 436 -2397 437 -2333
rect 499 -2397 500 -2333
rect 702 -2498 703 -2396
rect 758 -2498 759 -2396
rect 1059 -2397 1060 -2333
rect 1115 -2498 1116 -2396
rect 1192 -2397 1193 -2333
rect 1367 -2397 1368 -2333
rect 1388 -2498 1389 -2396
rect 219 -2399 220 -2333
rect 345 -2498 346 -2398
rect 436 -2498 437 -2398
rect 471 -2399 472 -2333
rect 499 -2498 500 -2398
rect 534 -2399 535 -2333
rect 576 -2498 577 -2398
rect 740 -2498 741 -2398
rect 814 -2399 815 -2333
rect 1059 -2498 1060 -2398
rect 1129 -2498 1130 -2398
rect 1402 -2399 1403 -2333
rect 149 -2401 150 -2333
rect 219 -2498 220 -2400
rect 233 -2401 234 -2333
rect 534 -2498 535 -2400
rect 590 -2498 591 -2400
rect 611 -2401 612 -2333
rect 621 -2401 622 -2333
rect 2130 -2498 2131 -2400
rect 149 -2498 150 -2402
rect 163 -2498 164 -2402
rect 233 -2498 234 -2402
rect 450 -2403 451 -2333
rect 597 -2498 598 -2402
rect 1031 -2403 1032 -2333
rect 1171 -2403 1172 -2333
rect 1465 -2498 1466 -2402
rect 359 -2405 360 -2333
rect 450 -2498 451 -2404
rect 611 -2498 612 -2404
rect 632 -2405 633 -2333
rect 646 -2498 647 -2404
rect 737 -2405 738 -2333
rect 814 -2498 815 -2404
rect 870 -2405 871 -2333
rect 884 -2498 885 -2404
rect 1374 -2498 1375 -2404
rect 198 -2407 199 -2333
rect 359 -2498 360 -2406
rect 443 -2407 444 -2333
rect 471 -2498 472 -2406
rect 478 -2498 479 -2406
rect 870 -2498 871 -2406
rect 919 -2498 920 -2406
rect 2249 -2407 2250 -2333
rect 184 -2409 185 -2333
rect 198 -2498 199 -2408
rect 443 -2498 444 -2408
rect 604 -2409 605 -2333
rect 628 -2409 629 -2333
rect 800 -2409 801 -2333
rect 828 -2409 829 -2333
rect 877 -2498 878 -2408
rect 922 -2409 923 -2333
rect 2312 -2498 2313 -2408
rect 135 -2411 136 -2333
rect 604 -2498 605 -2410
rect 632 -2498 633 -2410
rect 709 -2411 710 -2333
rect 737 -2498 738 -2410
rect 1514 -2498 1515 -2410
rect 135 -2498 136 -2412
rect 415 -2413 416 -2333
rect 660 -2498 661 -2412
rect 989 -2413 990 -2333
rect 1013 -2498 1014 -2412
rect 1402 -2498 1403 -2412
rect 184 -2498 185 -2414
rect 639 -2415 640 -2333
rect 670 -2415 671 -2333
rect 2270 -2415 2271 -2333
rect 268 -2498 269 -2416
rect 670 -2498 671 -2416
rect 800 -2498 801 -2416
rect 807 -2417 808 -2333
rect 828 -2498 829 -2416
rect 898 -2417 899 -2333
rect 922 -2498 923 -2416
rect 1724 -2417 1725 -2333
rect 2270 -2498 2271 -2416
rect 2298 -2417 2299 -2333
rect 366 -2419 367 -2333
rect 709 -2498 710 -2418
rect 835 -2498 836 -2418
rect 1003 -2419 1004 -2333
rect 1017 -2498 1018 -2418
rect 1157 -2419 1158 -2333
rect 1171 -2498 1172 -2418
rect 1913 -2419 1914 -2333
rect 121 -2421 122 -2333
rect 1003 -2498 1004 -2420
rect 1031 -2498 1032 -2420
rect 1731 -2421 1732 -2333
rect 1808 -2421 1809 -2333
rect 1913 -2498 1914 -2420
rect 121 -2498 122 -2422
rect 667 -2423 668 -2333
rect 863 -2498 864 -2422
rect 947 -2423 948 -2333
rect 957 -2498 958 -2422
rect 1157 -2498 1158 -2422
rect 1174 -2498 1175 -2422
rect 1297 -2498 1298 -2422
rect 1332 -2498 1333 -2422
rect 2298 -2498 2299 -2422
rect 107 -2425 108 -2333
rect 667 -2498 668 -2424
rect 898 -2498 899 -2424
rect 968 -2425 969 -2333
rect 975 -2425 976 -2333
rect 1549 -2498 1550 -2424
rect 1633 -2425 1634 -2333
rect 1808 -2498 1809 -2424
rect 107 -2498 108 -2426
rect 128 -2427 129 -2333
rect 156 -2427 157 -2333
rect 366 -2498 367 -2426
rect 415 -2498 416 -2426
rect 513 -2427 514 -2333
rect 555 -2427 556 -2333
rect 807 -2498 808 -2426
rect 933 -2427 934 -2333
rect 2158 -2498 2159 -2426
rect 79 -2429 80 -2333
rect 555 -2498 556 -2428
rect 639 -2498 640 -2428
rect 744 -2429 745 -2333
rect 936 -2429 937 -2333
rect 1626 -2429 1627 -2333
rect 1724 -2498 1725 -2428
rect 1937 -2429 1938 -2333
rect 2 -2431 3 -2333
rect 79 -2498 80 -2430
rect 86 -2431 87 -2333
rect 933 -2498 934 -2430
rect 947 -2498 948 -2430
rect 1066 -2431 1067 -2333
rect 1139 -2431 1140 -2333
rect 2249 -2498 2250 -2430
rect 2 -2498 3 -2432
rect 72 -2498 73 -2432
rect 86 -2498 87 -2432
rect 1500 -2433 1501 -2333
rect 1507 -2433 1508 -2333
rect 1633 -2498 1634 -2432
rect 1731 -2498 1732 -2432
rect 1864 -2433 1865 -2333
rect 128 -2498 129 -2434
rect 548 -2435 549 -2333
rect 695 -2435 696 -2333
rect 744 -2498 745 -2434
rect 961 -2498 962 -2434
rect 1122 -2435 1123 -2333
rect 1178 -2435 1179 -2333
rect 1255 -2498 1256 -2434
rect 1346 -2435 1347 -2333
rect 1864 -2498 1865 -2434
rect 96 -2437 97 -2333
rect 1178 -2498 1179 -2436
rect 1192 -2498 1193 -2436
rect 1325 -2437 1326 -2333
rect 1346 -2498 1347 -2436
rect 1423 -2437 1424 -2333
rect 1500 -2498 1501 -2436
rect 1584 -2437 1585 -2333
rect 1605 -2437 1606 -2333
rect 1626 -2498 1627 -2436
rect 58 -2439 59 -2333
rect 96 -2498 97 -2438
rect 156 -2498 157 -2438
rect 212 -2439 213 -2333
rect 513 -2498 514 -2438
rect 562 -2439 563 -2333
rect 688 -2439 689 -2333
rect 695 -2498 696 -2438
rect 968 -2498 969 -2438
rect 1010 -2439 1011 -2333
rect 1066 -2498 1067 -2438
rect 1143 -2439 1144 -2333
rect 1213 -2498 1214 -2438
rect 1605 -2498 1606 -2438
rect 58 -2498 59 -2440
rect 996 -2441 997 -2333
rect 1010 -2498 1011 -2440
rect 1101 -2441 1102 -2333
rect 1122 -2498 1123 -2440
rect 1206 -2441 1207 -2333
rect 1325 -2498 1326 -2440
rect 1496 -2441 1497 -2333
rect 1507 -2498 1508 -2440
rect 1556 -2441 1557 -2333
rect 1584 -2498 1585 -2440
rect 1654 -2441 1655 -2333
rect 142 -2443 143 -2333
rect 562 -2498 563 -2442
rect 793 -2498 794 -2442
rect 1101 -2498 1102 -2442
rect 1143 -2498 1144 -2442
rect 1521 -2443 1522 -2333
rect 1556 -2498 1557 -2442
rect 1619 -2443 1620 -2333
rect 93 -2445 94 -2333
rect 142 -2498 143 -2444
rect 205 -2445 206 -2333
rect 688 -2498 689 -2444
rect 975 -2498 976 -2444
rect 2018 -2498 2019 -2444
rect 93 -2498 94 -2446
rect 1822 -2498 1823 -2446
rect 205 -2498 206 -2448
rect 674 -2449 675 -2333
rect 996 -2498 997 -2448
rect 1045 -2449 1046 -2333
rect 1206 -2498 1207 -2448
rect 1234 -2449 1235 -2333
rect 1353 -2449 1354 -2333
rect 1423 -2498 1424 -2448
rect 1458 -2449 1459 -2333
rect 1619 -2498 1620 -2448
rect 212 -2498 213 -2450
rect 289 -2451 290 -2333
rect 548 -2498 549 -2450
rect 1804 -2498 1805 -2450
rect 289 -2498 290 -2452
rect 338 -2453 339 -2333
rect 674 -2498 675 -2452
rect 992 -2453 993 -2333
rect 1045 -2498 1046 -2452
rect 1094 -2453 1095 -2333
rect 1234 -2498 1235 -2452
rect 2336 -2453 2337 -2333
rect 338 -2498 339 -2454
rect 541 -2455 542 -2333
rect 926 -2455 927 -2333
rect 1094 -2498 1095 -2454
rect 1353 -2498 1354 -2454
rect 2144 -2455 2145 -2333
rect 541 -2498 542 -2456
rect 849 -2457 850 -2333
rect 992 -2498 993 -2456
rect 2046 -2498 2047 -2456
rect 772 -2459 773 -2333
rect 926 -2498 927 -2458
rect 1199 -2459 1200 -2333
rect 2144 -2498 2145 -2458
rect 23 -2498 24 -2460
rect 772 -2498 773 -2460
rect 849 -2498 850 -2460
rect 1290 -2461 1291 -2333
rect 1367 -2498 1368 -2460
rect 1430 -2461 1431 -2333
rect 1458 -2498 1459 -2460
rect 1577 -2498 1578 -2460
rect 1199 -2498 1200 -2462
rect 1283 -2463 1284 -2333
rect 1430 -2498 1431 -2462
rect 1640 -2463 1641 -2333
rect 1283 -2498 1284 -2464
rect 1416 -2465 1417 -2333
rect 1521 -2498 1522 -2464
rect 1661 -2465 1662 -2333
rect 373 -2467 374 -2333
rect 1661 -2498 1662 -2466
rect 373 -2498 374 -2468
rect 583 -2469 584 -2333
rect 1416 -2498 1417 -2468
rect 1472 -2469 1473 -2333
rect 1563 -2469 1564 -2333
rect 1654 -2498 1655 -2468
rect 583 -2498 584 -2470
rect 653 -2471 654 -2333
rect 1472 -2498 1473 -2470
rect 1601 -2498 1602 -2470
rect 1640 -2498 1641 -2470
rect 1815 -2471 1816 -2333
rect 653 -2498 654 -2472
rect 751 -2473 752 -2333
rect 1563 -2498 1564 -2472
rect 1689 -2473 1690 -2333
rect 1815 -2498 1816 -2472
rect 1871 -2473 1872 -2333
rect 751 -2498 752 -2474
rect 1073 -2475 1074 -2333
rect 1689 -2498 1690 -2474
rect 1759 -2475 1760 -2333
rect 1871 -2498 1872 -2474
rect 1920 -2475 1921 -2333
rect 1073 -2498 1074 -2476
rect 1955 -2477 1956 -2333
rect 1759 -2498 1760 -2478
rect 1794 -2479 1795 -2333
rect 1920 -2498 1921 -2478
rect 1962 -2479 1963 -2333
rect 1675 -2481 1676 -2333
rect 1794 -2498 1795 -2480
rect 1955 -2498 1956 -2480
rect 2004 -2481 2005 -2333
rect 1962 -2498 1963 -2482
rect 2025 -2483 2026 -2333
rect 1083 -2498 1084 -2484
rect 2025 -2498 2026 -2484
rect 2004 -2498 2005 -2486
rect 2032 -2487 2033 -2333
rect 2032 -2498 2033 -2488
rect 2081 -2489 2082 -2333
rect 1220 -2491 1221 -2333
rect 2081 -2498 2082 -2490
rect 1220 -2498 1221 -2492
rect 1241 -2493 1242 -2333
rect 1241 -2498 1242 -2494
rect 1269 -2495 1270 -2333
rect 1269 -2498 1270 -2496
rect 1570 -2498 1571 -2496
rect 5 -2508 6 -2506
rect 415 -2508 416 -2506
rect 464 -2508 465 -2506
rect 989 -2508 990 -2506
rect 992 -2508 993 -2506
rect 1073 -2508 1074 -2506
rect 1080 -2508 1081 -2506
rect 1794 -2508 1795 -2506
rect 1801 -2671 1802 -2507
rect 1934 -2508 1935 -2506
rect 2088 -2508 2089 -2506
rect 2091 -2566 2092 -2507
rect 9 -2510 10 -2506
rect 1409 -2510 1410 -2506
rect 1510 -2671 1511 -2509
rect 2053 -2510 2054 -2506
rect 2088 -2671 2089 -2509
rect 2158 -2510 2159 -2506
rect 9 -2671 10 -2511
rect 51 -2512 52 -2506
rect 54 -2671 55 -2511
rect 765 -2512 766 -2506
rect 775 -2512 776 -2506
rect 877 -2512 878 -2506
rect 926 -2512 927 -2506
rect 1083 -2512 1084 -2506
rect 1188 -2671 1189 -2511
rect 1696 -2512 1697 -2506
rect 1717 -2512 1718 -2506
rect 1717 -2671 1718 -2511
rect 1717 -2512 1718 -2506
rect 1717 -2671 1718 -2511
rect 1794 -2671 1795 -2511
rect 1885 -2512 1886 -2506
rect 1934 -2671 1935 -2511
rect 2025 -2512 2026 -2506
rect 2053 -2671 2054 -2511
rect 2130 -2512 2131 -2506
rect 16 -2671 17 -2513
rect 37 -2514 38 -2506
rect 40 -2514 41 -2506
rect 1248 -2514 1249 -2506
rect 1290 -2514 1291 -2506
rect 1808 -2514 1809 -2506
rect 1885 -2671 1886 -2513
rect 1997 -2514 1998 -2506
rect 2025 -2671 2026 -2513
rect 2102 -2514 2103 -2506
rect 2130 -2671 2131 -2513
rect 2193 -2514 2194 -2506
rect 33 -2516 34 -2506
rect 933 -2516 934 -2506
rect 950 -2671 951 -2515
rect 1290 -2671 1291 -2515
rect 1335 -2516 1336 -2506
rect 2109 -2516 2110 -2506
rect 37 -2671 38 -2517
rect 51 -2671 52 -2517
rect 58 -2518 59 -2506
rect 1465 -2518 1466 -2506
rect 1521 -2518 1522 -2506
rect 1521 -2671 1522 -2517
rect 1521 -2518 1522 -2506
rect 1521 -2671 1522 -2517
rect 1580 -2518 1581 -2506
rect 1647 -2518 1648 -2506
rect 1678 -2518 1679 -2506
rect 1969 -2518 1970 -2506
rect 1997 -2671 1998 -2517
rect 2060 -2518 2061 -2506
rect 2102 -2671 2103 -2517
rect 2242 -2518 2243 -2506
rect 44 -2520 45 -2506
rect 75 -2671 76 -2519
rect 93 -2520 94 -2506
rect 1150 -2520 1151 -2506
rect 1195 -2671 1196 -2519
rect 1906 -2520 1907 -2506
rect 1969 -2671 1970 -2519
rect 2032 -2520 2033 -2506
rect 2109 -2671 2110 -2519
rect 2172 -2520 2173 -2506
rect 2242 -2671 2243 -2519
rect 2291 -2520 2292 -2506
rect 44 -2671 45 -2521
rect 527 -2522 528 -2506
rect 541 -2522 542 -2506
rect 978 -2522 979 -2506
rect 989 -2671 990 -2521
rect 1174 -2522 1175 -2506
rect 1199 -2522 1200 -2506
rect 1332 -2522 1333 -2506
rect 1356 -2522 1357 -2506
rect 1696 -2671 1697 -2521
rect 1804 -2522 1805 -2506
rect 2186 -2522 2187 -2506
rect 58 -2671 59 -2523
rect 61 -2524 62 -2506
rect 72 -2524 73 -2506
rect 1237 -2671 1238 -2523
rect 1332 -2671 1333 -2523
rect 1416 -2524 1417 -2506
rect 1458 -2524 1459 -2506
rect 2032 -2671 2033 -2523
rect 2172 -2671 2173 -2523
rect 2235 -2524 2236 -2506
rect 72 -2671 73 -2525
rect 366 -2526 367 -2506
rect 373 -2526 374 -2506
rect 789 -2671 790 -2525
rect 817 -2671 818 -2525
rect 2060 -2671 2061 -2525
rect 2186 -2671 2187 -2525
rect 2256 -2526 2257 -2506
rect 93 -2671 94 -2527
rect 114 -2528 115 -2506
rect 128 -2528 129 -2506
rect 810 -2671 811 -2527
rect 859 -2528 860 -2506
rect 1675 -2671 1676 -2527
rect 1808 -2671 1809 -2527
rect 1871 -2528 1872 -2506
rect 2235 -2671 2236 -2527
rect 2284 -2528 2285 -2506
rect 107 -2671 108 -2529
rect 261 -2530 262 -2506
rect 268 -2530 269 -2506
rect 870 -2671 871 -2529
rect 877 -2671 878 -2529
rect 1311 -2530 1312 -2506
rect 1360 -2530 1361 -2506
rect 2116 -2530 2117 -2506
rect 110 -2532 111 -2506
rect 1360 -2671 1361 -2531
rect 1374 -2532 1375 -2506
rect 1941 -2532 1942 -2506
rect 2116 -2671 2117 -2531
rect 2123 -2532 2124 -2506
rect 131 -2671 132 -2533
rect 968 -2534 969 -2506
rect 1006 -2671 1007 -2533
rect 1031 -2534 1032 -2506
rect 1038 -2534 1039 -2506
rect 1150 -2671 1151 -2533
rect 1216 -2534 1217 -2506
rect 2270 -2534 2271 -2506
rect 19 -2536 20 -2506
rect 1031 -2671 1032 -2535
rect 1038 -2671 1039 -2535
rect 1157 -2536 1158 -2506
rect 1311 -2671 1312 -2535
rect 1843 -2536 1844 -2506
rect 1871 -2671 1872 -2535
rect 1927 -2536 1928 -2506
rect 1941 -2671 1942 -2535
rect 2165 -2536 2166 -2506
rect 2270 -2671 2271 -2535
rect 2312 -2536 2313 -2506
rect 149 -2538 150 -2506
rect 268 -2671 269 -2537
rect 275 -2538 276 -2506
rect 793 -2538 794 -2506
rect 898 -2538 899 -2506
rect 933 -2671 934 -2537
rect 940 -2538 941 -2506
rect 1199 -2671 1200 -2537
rect 1377 -2538 1378 -2506
rect 1654 -2538 1655 -2506
rect 1843 -2671 1844 -2537
rect 1899 -2538 1900 -2506
rect 2123 -2671 2124 -2537
rect 2179 -2538 2180 -2506
rect 103 -2671 104 -2539
rect 898 -2671 899 -2539
rect 919 -2540 920 -2506
rect 968 -2671 969 -2539
rect 1010 -2540 1011 -2506
rect 1122 -2540 1123 -2506
rect 1402 -2540 1403 -2506
rect 1405 -2566 1406 -2539
rect 1416 -2671 1417 -2539
rect 1437 -2540 1438 -2506
rect 1458 -2671 1459 -2539
rect 1514 -2540 1515 -2506
rect 1580 -2671 1581 -2539
rect 2004 -2540 2005 -2506
rect 2165 -2671 2166 -2539
rect 2228 -2540 2229 -2506
rect 128 -2671 129 -2541
rect 940 -2671 941 -2541
rect 1013 -2542 1014 -2506
rect 1374 -2671 1375 -2541
rect 1402 -2671 1403 -2541
rect 1444 -2542 1445 -2506
rect 1465 -2671 1466 -2541
rect 1542 -2542 1543 -2506
rect 1601 -2542 1602 -2506
rect 2095 -2542 2096 -2506
rect 2179 -2671 2180 -2541
rect 2249 -2542 2250 -2506
rect 149 -2671 150 -2543
rect 429 -2544 430 -2506
rect 478 -2544 479 -2506
rect 1661 -2544 1662 -2506
rect 1766 -2544 1767 -2506
rect 2228 -2671 2229 -2543
rect 163 -2546 164 -2506
rect 177 -2546 178 -2506
rect 191 -2546 192 -2506
rect 261 -2671 262 -2545
rect 303 -2546 304 -2506
rect 411 -2671 412 -2545
rect 429 -2671 430 -2545
rect 1440 -2671 1441 -2545
rect 1444 -2671 1445 -2545
rect 1619 -2546 1620 -2506
rect 1647 -2671 1648 -2545
rect 1710 -2546 1711 -2506
rect 1899 -2671 1900 -2545
rect 1962 -2546 1963 -2506
rect 163 -2671 164 -2547
rect 1353 -2548 1354 -2506
rect 1437 -2671 1438 -2547
rect 1703 -2548 1704 -2506
rect 1710 -2671 1711 -2547
rect 1920 -2548 1921 -2506
rect 96 -2550 97 -2506
rect 1353 -2671 1354 -2549
rect 1500 -2550 1501 -2506
rect 1514 -2671 1515 -2549
rect 1542 -2671 1543 -2549
rect 1563 -2550 1564 -2506
rect 1612 -2550 1613 -2506
rect 1927 -2671 1928 -2549
rect 177 -2671 178 -2551
rect 583 -2552 584 -2506
rect 604 -2671 605 -2551
rect 891 -2552 892 -2506
rect 894 -2671 895 -2551
rect 1766 -2671 1767 -2551
rect 1920 -2671 1921 -2551
rect 2011 -2552 2012 -2506
rect 191 -2671 192 -2553
rect 1577 -2554 1578 -2506
rect 1619 -2671 1620 -2553
rect 1976 -2554 1977 -2506
rect 201 -2671 202 -2555
rect 607 -2556 608 -2506
rect 632 -2556 633 -2506
rect 1213 -2556 1214 -2506
rect 1272 -2556 1273 -2506
rect 1703 -2671 1704 -2555
rect 1948 -2556 1949 -2506
rect 2011 -2671 2012 -2555
rect 205 -2558 206 -2506
rect 275 -2671 276 -2557
rect 310 -2558 311 -2506
rect 1269 -2558 1270 -2506
rect 1314 -2671 1315 -2557
rect 2095 -2671 2096 -2557
rect 198 -2560 199 -2506
rect 205 -2671 206 -2559
rect 240 -2560 241 -2506
rect 541 -2671 542 -2559
rect 555 -2560 556 -2506
rect 740 -2560 741 -2506
rect 751 -2560 752 -2506
rect 772 -2671 773 -2559
rect 926 -2671 927 -2559
rect 1297 -2560 1298 -2506
rect 1451 -2560 1452 -2506
rect 1612 -2671 1613 -2559
rect 1654 -2671 1655 -2559
rect 1755 -2671 1756 -2559
rect 1948 -2671 1949 -2559
rect 2039 -2560 2040 -2506
rect 198 -2671 199 -2561
rect 611 -2562 612 -2506
rect 709 -2562 710 -2506
rect 1052 -2562 1053 -2506
rect 1066 -2562 1067 -2506
rect 1409 -2671 1410 -2561
rect 1451 -2671 1452 -2561
rect 1570 -2562 1571 -2506
rect 1661 -2671 1662 -2561
rect 1738 -2562 1739 -2506
rect 1976 -2671 1977 -2561
rect 2046 -2562 2047 -2506
rect 240 -2671 241 -2563
rect 415 -2671 416 -2563
rect 457 -2564 458 -2506
rect 611 -2671 612 -2563
rect 709 -2671 710 -2563
rect 730 -2564 731 -2506
rect 737 -2564 738 -2506
rect 2004 -2671 2005 -2563
rect 2046 -2671 2047 -2563
rect 2207 -2564 2208 -2506
rect 254 -2566 255 -2506
rect 303 -2671 304 -2565
rect 310 -2671 311 -2565
rect 422 -2566 423 -2506
rect 457 -2671 458 -2565
rect 558 -2671 559 -2565
rect 562 -2566 563 -2506
rect 765 -2671 766 -2565
rect 873 -2566 874 -2506
rect 2039 -2671 2040 -2565
rect 2158 -2671 2159 -2565
rect 135 -2568 136 -2506
rect 254 -2671 255 -2567
rect 352 -2568 353 -2506
rect 1010 -2671 1011 -2567
rect 1017 -2568 1018 -2506
rect 2193 -2671 2194 -2567
rect 135 -2671 136 -2569
rect 247 -2570 248 -2506
rect 352 -2671 353 -2569
rect 450 -2570 451 -2506
rect 492 -2570 493 -2506
rect 1157 -2671 1158 -2569
rect 1185 -2570 1186 -2506
rect 1962 -2671 1963 -2569
rect 184 -2572 185 -2506
rect 492 -2671 493 -2571
rect 562 -2671 563 -2571
rect 863 -2572 864 -2506
rect 1017 -2671 1018 -2571
rect 1108 -2572 1109 -2506
rect 1122 -2671 1123 -2571
rect 1423 -2572 1424 -2506
rect 1479 -2572 1480 -2506
rect 1563 -2671 1564 -2571
rect 1570 -2671 1571 -2571
rect 1605 -2572 1606 -2506
rect 1738 -2671 1739 -2571
rect 1787 -2572 1788 -2506
rect 142 -2574 143 -2506
rect 863 -2671 864 -2573
rect 1024 -2574 1025 -2506
rect 1024 -2671 1025 -2573
rect 1024 -2574 1025 -2506
rect 1024 -2671 1025 -2573
rect 1052 -2671 1053 -2573
rect 1115 -2574 1116 -2506
rect 1213 -2671 1214 -2573
rect 1325 -2574 1326 -2506
rect 1423 -2671 1424 -2573
rect 1528 -2574 1529 -2506
rect 1605 -2671 1606 -2573
rect 1682 -2574 1683 -2506
rect 1787 -2671 1788 -2573
rect 1864 -2574 1865 -2506
rect 142 -2671 143 -2575
rect 891 -2671 892 -2575
rect 1066 -2671 1067 -2575
rect 1318 -2576 1319 -2506
rect 1479 -2671 1480 -2575
rect 1486 -2576 1487 -2506
rect 1500 -2671 1501 -2575
rect 1584 -2576 1585 -2506
rect 1682 -2671 1683 -2575
rect 1759 -2576 1760 -2506
rect 1850 -2576 1851 -2506
rect 1864 -2671 1865 -2575
rect 184 -2671 185 -2577
rect 975 -2578 976 -2506
rect 1073 -2671 1074 -2577
rect 1094 -2578 1095 -2506
rect 1269 -2671 1270 -2577
rect 1388 -2578 1389 -2506
rect 1486 -2671 1487 -2577
rect 1549 -2578 1550 -2506
rect 1584 -2671 1585 -2577
rect 1626 -2578 1627 -2506
rect 1731 -2578 1732 -2506
rect 1759 -2671 1760 -2577
rect 1850 -2671 1851 -2577
rect 1955 -2578 1956 -2506
rect 219 -2580 220 -2506
rect 422 -2671 423 -2579
rect 450 -2671 451 -2579
rect 828 -2580 829 -2506
rect 842 -2580 843 -2506
rect 975 -2671 976 -2579
rect 1080 -2671 1081 -2579
rect 1087 -2580 1088 -2506
rect 1094 -2671 1095 -2579
rect 1143 -2580 1144 -2506
rect 1297 -2671 1298 -2579
rect 1395 -2580 1396 -2506
rect 1528 -2671 1529 -2579
rect 1633 -2580 1634 -2506
rect 1955 -2671 1956 -2579
rect 2018 -2580 2019 -2506
rect 86 -2582 87 -2506
rect 842 -2671 843 -2581
rect 1087 -2671 1088 -2581
rect 1381 -2582 1382 -2506
rect 1388 -2671 1389 -2581
rect 1493 -2582 1494 -2506
rect 1549 -2671 1550 -2581
rect 1745 -2582 1746 -2506
rect 1990 -2582 1991 -2506
rect 2018 -2671 2019 -2581
rect 86 -2671 87 -2583
rect 922 -2584 923 -2506
rect 1143 -2671 1144 -2583
rect 1220 -2584 1221 -2506
rect 1234 -2584 1235 -2506
rect 1381 -2671 1382 -2583
rect 1395 -2671 1396 -2583
rect 1829 -2584 1830 -2506
rect 1878 -2584 1879 -2506
rect 1990 -2671 1991 -2583
rect 26 -2671 27 -2585
rect 1878 -2671 1879 -2585
rect 219 -2671 220 -2587
rect 317 -2588 318 -2506
rect 359 -2588 360 -2506
rect 1363 -2588 1364 -2506
rect 1430 -2588 1431 -2506
rect 1493 -2671 1494 -2587
rect 1591 -2588 1592 -2506
rect 1731 -2671 1732 -2587
rect 1745 -2671 1746 -2587
rect 1815 -2588 1816 -2506
rect 1829 -2671 1830 -2587
rect 1836 -2588 1837 -2506
rect 212 -2590 213 -2506
rect 317 -2671 318 -2589
rect 331 -2590 332 -2506
rect 359 -2671 360 -2589
rect 366 -2671 367 -2589
rect 506 -2590 507 -2506
rect 569 -2590 570 -2506
rect 632 -2671 633 -2589
rect 646 -2590 647 -2506
rect 1185 -2671 1186 -2589
rect 1220 -2671 1221 -2589
rect 1339 -2590 1340 -2506
rect 1430 -2671 1431 -2589
rect 1598 -2590 1599 -2506
rect 1626 -2671 1627 -2589
rect 1689 -2590 1690 -2506
rect 1815 -2671 1816 -2589
rect 1857 -2590 1858 -2506
rect 212 -2671 213 -2591
rect 597 -2592 598 -2506
rect 646 -2671 647 -2591
rect 688 -2592 689 -2506
rect 716 -2592 717 -2506
rect 793 -2671 794 -2591
rect 828 -2671 829 -2591
rect 1304 -2592 1305 -2506
rect 1318 -2671 1319 -2591
rect 1535 -2592 1536 -2506
rect 1591 -2671 1592 -2591
rect 1773 -2592 1774 -2506
rect 1836 -2671 1837 -2591
rect 1892 -2592 1893 -2506
rect 68 -2671 69 -2593
rect 688 -2671 689 -2593
rect 716 -2671 717 -2593
rect 1206 -2594 1207 -2506
rect 1234 -2671 1235 -2593
rect 1262 -2594 1263 -2506
rect 1339 -2671 1340 -2593
rect 1398 -2671 1399 -2593
rect 1472 -2594 1473 -2506
rect 1535 -2671 1536 -2593
rect 1598 -2671 1599 -2593
rect 1668 -2594 1669 -2506
rect 1773 -2671 1774 -2593
rect 1822 -2594 1823 -2506
rect 1857 -2671 1858 -2593
rect 2074 -2594 2075 -2506
rect 226 -2596 227 -2506
rect 247 -2671 248 -2595
rect 282 -2596 283 -2506
rect 1115 -2671 1116 -2595
rect 1171 -2596 1172 -2506
rect 1892 -2671 1893 -2595
rect 2074 -2671 2075 -2595
rect 2144 -2596 2145 -2506
rect 170 -2598 171 -2506
rect 226 -2671 227 -2597
rect 282 -2671 283 -2597
rect 670 -2598 671 -2506
rect 723 -2598 724 -2506
rect 737 -2671 738 -2597
rect 751 -2671 752 -2597
rect 1125 -2671 1126 -2597
rect 1171 -2671 1172 -2597
rect 1255 -2598 1256 -2506
rect 1262 -2671 1263 -2597
rect 1346 -2598 1347 -2506
rect 1412 -2671 1413 -2597
rect 1472 -2671 1473 -2597
rect 1633 -2671 1634 -2597
rect 2280 -2598 2281 -2506
rect 166 -2600 167 -2506
rect 170 -2671 171 -2599
rect 331 -2671 332 -2599
rect 345 -2600 346 -2506
rect 373 -2671 374 -2599
rect 394 -2600 395 -2506
rect 401 -2600 402 -2506
rect 856 -2600 857 -2506
rect 954 -2600 955 -2506
rect 1346 -2671 1347 -2599
rect 1640 -2600 1641 -2506
rect 1689 -2671 1690 -2599
rect 1822 -2671 1823 -2599
rect 1913 -2600 1914 -2506
rect 2144 -2671 2145 -2599
rect 2214 -2600 2215 -2506
rect 30 -2602 31 -2506
rect 345 -2671 346 -2601
rect 380 -2602 381 -2506
rect 527 -2671 528 -2601
rect 569 -2671 570 -2601
rect 814 -2602 815 -2506
rect 824 -2671 825 -2601
rect 1304 -2671 1305 -2601
rect 1640 -2671 1641 -2601
rect 1724 -2602 1725 -2506
rect 1913 -2671 1914 -2601
rect 1983 -2602 1984 -2506
rect 2214 -2671 2215 -2601
rect 2263 -2602 2264 -2506
rect 30 -2671 31 -2603
rect 485 -2604 486 -2506
rect 506 -2671 507 -2603
rect 849 -2604 850 -2506
rect 1178 -2604 1179 -2506
rect 1983 -2671 1984 -2603
rect 2263 -2671 2264 -2603
rect 2305 -2604 2306 -2506
rect 79 -2606 80 -2506
rect 856 -2671 857 -2605
rect 1003 -2606 1004 -2506
rect 1178 -2671 1179 -2605
rect 1206 -2671 1207 -2605
rect 1283 -2606 1284 -2506
rect 1447 -2671 1448 -2605
rect 1724 -2671 1725 -2605
rect 79 -2671 80 -2607
rect 548 -2608 549 -2506
rect 583 -2671 584 -2607
rect 800 -2608 801 -2506
rect 807 -2608 808 -2506
rect 1003 -2671 1004 -2607
rect 1255 -2671 1256 -2607
rect 1577 -2671 1578 -2607
rect 1668 -2671 1669 -2607
rect 1752 -2608 1753 -2506
rect 156 -2610 157 -2506
rect 401 -2671 402 -2609
rect 408 -2610 409 -2506
rect 464 -2671 465 -2609
rect 485 -2671 486 -2609
rect 639 -2610 640 -2506
rect 726 -2671 727 -2609
rect 2081 -2610 2082 -2506
rect 156 -2671 157 -2611
rect 555 -2671 556 -2611
rect 597 -2671 598 -2611
rect 957 -2612 958 -2506
rect 1752 -2671 1753 -2611
rect 2298 -2612 2299 -2506
rect 289 -2614 290 -2506
rect 408 -2671 409 -2613
rect 520 -2614 521 -2506
rect 954 -2671 955 -2613
rect 2081 -2671 2082 -2613
rect 2151 -2614 2152 -2506
rect 65 -2616 66 -2506
rect 289 -2671 290 -2615
rect 380 -2671 381 -2615
rect 660 -2616 661 -2506
rect 730 -2671 731 -2615
rect 982 -2616 983 -2506
rect 2151 -2671 2152 -2615
rect 2221 -2616 2222 -2506
rect 65 -2671 66 -2617
rect 2067 -2618 2068 -2506
rect 387 -2620 388 -2506
rect 478 -2671 479 -2619
rect 513 -2620 514 -2506
rect 660 -2671 661 -2619
rect 758 -2620 759 -2506
rect 1108 -2671 1109 -2619
rect 2067 -2671 2068 -2619
rect 2137 -2620 2138 -2506
rect 338 -2622 339 -2506
rect 387 -2671 388 -2621
rect 394 -2671 395 -2621
rect 1055 -2622 1056 -2506
rect 2137 -2671 2138 -2621
rect 2200 -2622 2201 -2506
rect 338 -2671 339 -2623
rect 499 -2624 500 -2506
rect 513 -2671 514 -2623
rect 695 -2624 696 -2506
rect 786 -2624 787 -2506
rect 1283 -2671 1284 -2623
rect 443 -2626 444 -2506
rect 499 -2671 500 -2625
rect 520 -2671 521 -2625
rect 576 -2626 577 -2506
rect 590 -2626 591 -2506
rect 758 -2671 759 -2625
rect 800 -2671 801 -2625
rect 1556 -2626 1557 -2506
rect 233 -2628 234 -2506
rect 443 -2671 444 -2627
rect 534 -2628 535 -2506
rect 590 -2671 591 -2627
rect 618 -2628 619 -2506
rect 814 -2671 815 -2627
rect 849 -2671 850 -2627
rect 1101 -2628 1102 -2506
rect 1507 -2628 1508 -2506
rect 1556 -2671 1557 -2627
rect 233 -2671 234 -2629
rect 674 -2630 675 -2506
rect 695 -2671 696 -2629
rect 996 -2630 997 -2506
rect 1101 -2671 1102 -2629
rect 1136 -2630 1137 -2506
rect 1248 -2671 1249 -2629
rect 1507 -2671 1508 -2629
rect 324 -2632 325 -2506
rect 534 -2671 535 -2631
rect 548 -2671 549 -2631
rect 835 -2632 836 -2506
rect 982 -2671 983 -2631
rect 1059 -2632 1060 -2506
rect 1136 -2671 1137 -2631
rect 2221 -2671 2222 -2631
rect 324 -2671 325 -2633
rect 471 -2634 472 -2506
rect 576 -2671 577 -2633
rect 786 -2671 787 -2633
rect 796 -2634 797 -2506
rect 1059 -2671 1060 -2633
rect 23 -2636 24 -2506
rect 471 -2671 472 -2635
rect 618 -2671 619 -2635
rect 884 -2636 885 -2506
rect 996 -2671 997 -2635
rect 1045 -2636 1046 -2506
rect 639 -2671 640 -2637
rect 681 -2638 682 -2506
rect 779 -2638 780 -2506
rect 835 -2671 836 -2637
rect 884 -2671 885 -2637
rect 905 -2638 906 -2506
rect 1045 -2671 1046 -2637
rect 1276 -2638 1277 -2506
rect 121 -2640 122 -2506
rect 779 -2671 780 -2639
rect 1241 -2640 1242 -2506
rect 1276 -2671 1277 -2639
rect 481 -2642 482 -2506
rect 905 -2671 906 -2641
rect 1241 -2671 1242 -2641
rect 1780 -2642 1781 -2506
rect 625 -2644 626 -2506
rect 681 -2671 682 -2643
rect 1013 -2671 1014 -2643
rect 1780 -2671 1781 -2643
rect 625 -2671 626 -2645
rect 912 -2646 913 -2506
rect 667 -2648 668 -2506
rect 2200 -2671 2201 -2647
rect 667 -2671 668 -2649
rect 702 -2650 703 -2506
rect 912 -2671 913 -2649
rect 1129 -2650 1130 -2506
rect 674 -2671 675 -2651
rect 821 -2652 822 -2506
rect 1129 -2671 1130 -2651
rect 1164 -2652 1165 -2506
rect 114 -2671 115 -2653
rect 821 -2671 822 -2653
rect 1164 -2671 1165 -2653
rect 1227 -2654 1228 -2506
rect 702 -2671 703 -2655
rect 744 -2656 745 -2506
rect 1227 -2671 1228 -2655
rect 1367 -2656 1368 -2506
rect 744 -2671 745 -2657
rect 961 -2658 962 -2506
rect 1192 -2658 1193 -2506
rect 1367 -2671 1368 -2657
rect 947 -2660 948 -2506
rect 961 -2671 962 -2659
rect 1192 -2671 1193 -2659
rect 1906 -2671 1907 -2659
rect 296 -2662 297 -2506
rect 947 -2671 948 -2661
rect 296 -2671 297 -2663
rect 436 -2664 437 -2506
rect 436 -2671 437 -2665
rect 653 -2666 654 -2506
rect 100 -2668 101 -2506
rect 653 -2671 654 -2667
rect 100 -2671 101 -2669
rect 121 -2671 122 -2669
rect 2 -2834 3 -2680
rect 68 -2681 69 -2679
rect 103 -2681 104 -2679
rect 338 -2681 339 -2679
rect 373 -2681 374 -2679
rect 373 -2834 374 -2680
rect 373 -2681 374 -2679
rect 373 -2834 374 -2680
rect 432 -2834 433 -2680
rect 464 -2681 465 -2679
rect 506 -2681 507 -2679
rect 733 -2834 734 -2680
rect 758 -2681 759 -2679
rect 838 -2834 839 -2680
rect 915 -2834 916 -2680
rect 2046 -2681 2047 -2679
rect 2200 -2681 2201 -2679
rect 2200 -2834 2201 -2680
rect 2200 -2681 2201 -2679
rect 2200 -2834 2201 -2680
rect 2224 -2834 2225 -2680
rect 2270 -2681 2271 -2679
rect 16 -2683 17 -2679
rect 250 -2834 251 -2682
rect 338 -2834 339 -2682
rect 345 -2683 346 -2679
rect 506 -2834 507 -2682
rect 779 -2683 780 -2679
rect 786 -2683 787 -2679
rect 1150 -2683 1151 -2679
rect 1185 -2683 1186 -2679
rect 1885 -2683 1886 -2679
rect 1927 -2683 1928 -2679
rect 2259 -2834 2260 -2682
rect 16 -2834 17 -2684
rect 695 -2685 696 -2679
rect 709 -2685 710 -2679
rect 957 -2685 958 -2679
rect 978 -2834 979 -2684
rect 1283 -2685 1284 -2679
rect 1286 -2834 1287 -2684
rect 1458 -2685 1459 -2679
rect 1489 -2834 1490 -2684
rect 1591 -2685 1592 -2679
rect 1605 -2685 1606 -2679
rect 1605 -2834 1606 -2684
rect 1605 -2685 1606 -2679
rect 1605 -2834 1606 -2684
rect 1619 -2685 1620 -2679
rect 1885 -2834 1886 -2684
rect 1934 -2685 1935 -2679
rect 1934 -2834 1935 -2684
rect 1934 -2685 1935 -2679
rect 1934 -2834 1935 -2684
rect 1948 -2685 1949 -2679
rect 1948 -2834 1949 -2684
rect 1948 -2685 1949 -2679
rect 1948 -2834 1949 -2684
rect 2235 -2685 2236 -2679
rect 2235 -2834 2236 -2684
rect 2235 -2685 2236 -2679
rect 2235 -2834 2236 -2684
rect 2242 -2685 2243 -2679
rect 2242 -2834 2243 -2684
rect 2242 -2685 2243 -2679
rect 2242 -2834 2243 -2684
rect 23 -2687 24 -2679
rect 135 -2687 136 -2679
rect 156 -2687 157 -2679
rect 1055 -2834 1056 -2686
rect 1062 -2834 1063 -2686
rect 1136 -2834 1137 -2686
rect 1139 -2687 1140 -2679
rect 1479 -2687 1480 -2679
rect 1577 -2687 1578 -2679
rect 2249 -2834 2250 -2686
rect 23 -2834 24 -2688
rect 520 -2689 521 -2679
rect 548 -2689 549 -2679
rect 817 -2689 818 -2679
rect 821 -2689 822 -2679
rect 933 -2689 934 -2679
rect 954 -2689 955 -2679
rect 1143 -2689 1144 -2679
rect 1185 -2834 1186 -2688
rect 1206 -2689 1207 -2679
rect 1234 -2689 1235 -2679
rect 2004 -2689 2005 -2679
rect 26 -2691 27 -2679
rect 842 -2691 843 -2679
rect 919 -2691 920 -2679
rect 1955 -2691 1956 -2679
rect 58 -2693 59 -2679
rect 58 -2834 59 -2692
rect 58 -2693 59 -2679
rect 58 -2834 59 -2692
rect 65 -2693 66 -2679
rect 86 -2693 87 -2679
rect 110 -2834 111 -2692
rect 282 -2693 283 -2679
rect 345 -2834 346 -2692
rect 359 -2693 360 -2679
rect 387 -2693 388 -2679
rect 520 -2834 521 -2692
rect 555 -2693 556 -2679
rect 632 -2693 633 -2679
rect 653 -2693 654 -2679
rect 653 -2834 654 -2692
rect 653 -2693 654 -2679
rect 653 -2834 654 -2692
rect 681 -2693 682 -2679
rect 723 -2834 724 -2692
rect 765 -2693 766 -2679
rect 950 -2693 951 -2679
rect 954 -2834 955 -2692
rect 975 -2693 976 -2679
rect 1013 -2693 1014 -2679
rect 2102 -2693 2103 -2679
rect 65 -2834 66 -2694
rect 996 -2695 997 -2679
rect 1041 -2695 1042 -2679
rect 1871 -2695 1872 -2679
rect 1955 -2834 1956 -2694
rect 1976 -2695 1977 -2679
rect 2102 -2834 2103 -2694
rect 2137 -2695 2138 -2679
rect 82 -2834 83 -2696
rect 632 -2834 633 -2696
rect 681 -2834 682 -2696
rect 716 -2697 717 -2679
rect 765 -2834 766 -2696
rect 1220 -2697 1221 -2679
rect 1234 -2834 1235 -2696
rect 1395 -2697 1396 -2679
rect 1423 -2697 1424 -2679
rect 1458 -2834 1459 -2696
rect 1479 -2834 1480 -2696
rect 1556 -2697 1557 -2679
rect 1584 -2697 1585 -2679
rect 1685 -2834 1686 -2696
rect 1755 -2697 1756 -2679
rect 2158 -2697 2159 -2679
rect 86 -2834 87 -2698
rect 1258 -2834 1259 -2698
rect 1318 -2699 1319 -2679
rect 2270 -2834 2271 -2698
rect 107 -2701 108 -2679
rect 555 -2834 556 -2700
rect 558 -2701 559 -2679
rect 660 -2701 661 -2679
rect 695 -2834 696 -2700
rect 737 -2701 738 -2679
rect 772 -2701 773 -2679
rect 891 -2834 892 -2700
rect 919 -2834 920 -2700
rect 961 -2701 962 -2679
rect 975 -2834 976 -2700
rect 1927 -2834 1928 -2700
rect 1976 -2834 1977 -2700
rect 2018 -2701 2019 -2679
rect 2130 -2701 2131 -2679
rect 2137 -2834 2138 -2700
rect 2158 -2834 2159 -2700
rect 2172 -2701 2173 -2679
rect 121 -2703 122 -2679
rect 128 -2703 129 -2679
rect 163 -2703 164 -2679
rect 548 -2834 549 -2702
rect 562 -2703 563 -2679
rect 1038 -2703 1039 -2679
rect 1066 -2703 1067 -2679
rect 1143 -2834 1144 -2702
rect 1195 -2703 1196 -2679
rect 1444 -2703 1445 -2679
rect 1556 -2834 1557 -2702
rect 1787 -2703 1788 -2679
rect 1871 -2834 1872 -2702
rect 1906 -2703 1907 -2679
rect 2011 -2703 2012 -2679
rect 2018 -2834 2019 -2702
rect 2130 -2834 2131 -2702
rect 2144 -2703 2145 -2679
rect 51 -2705 52 -2679
rect 1444 -2834 1445 -2704
rect 1584 -2834 1585 -2704
rect 1696 -2705 1697 -2679
rect 1759 -2705 1760 -2679
rect 2004 -2834 2005 -2704
rect 2144 -2834 2145 -2704
rect 2151 -2705 2152 -2679
rect 51 -2834 52 -2706
rect 982 -2707 983 -2679
rect 996 -2834 997 -2706
rect 1213 -2707 1214 -2679
rect 1220 -2834 1221 -2706
rect 1262 -2707 1263 -2679
rect 1360 -2707 1361 -2679
rect 1591 -2834 1592 -2706
rect 1619 -2834 1620 -2706
rect 1633 -2707 1634 -2679
rect 1647 -2707 1648 -2679
rect 1706 -2834 1707 -2706
rect 1759 -2834 1760 -2706
rect 1766 -2707 1767 -2679
rect 1773 -2707 1774 -2679
rect 1773 -2834 1774 -2706
rect 1773 -2707 1774 -2679
rect 1773 -2834 1774 -2706
rect 1899 -2707 1900 -2679
rect 1906 -2834 1907 -2706
rect 2151 -2834 2152 -2706
rect 2165 -2707 2166 -2679
rect 121 -2834 122 -2708
rect 667 -2709 668 -2679
rect 730 -2709 731 -2679
rect 1038 -2834 1039 -2708
rect 1066 -2834 1067 -2708
rect 1129 -2709 1130 -2679
rect 1206 -2834 1207 -2708
rect 1227 -2709 1228 -2679
rect 1241 -2709 1242 -2679
rect 1892 -2709 1893 -2679
rect 1899 -2834 1900 -2708
rect 1913 -2709 1914 -2679
rect 2165 -2834 2166 -2708
rect 2179 -2709 2180 -2679
rect 128 -2834 129 -2710
rect 436 -2711 437 -2679
rect 457 -2711 458 -2679
rect 562 -2834 563 -2710
rect 576 -2711 577 -2679
rect 709 -2834 710 -2710
rect 730 -2834 731 -2710
rect 2179 -2834 2180 -2710
rect 93 -2713 94 -2679
rect 436 -2834 437 -2712
rect 513 -2713 514 -2679
rect 737 -2834 738 -2712
rect 772 -2834 773 -2712
rect 1171 -2713 1172 -2679
rect 1213 -2834 1214 -2712
rect 1269 -2713 1270 -2679
rect 1276 -2713 1277 -2679
rect 1360 -2834 1361 -2712
rect 1374 -2713 1375 -2679
rect 1507 -2713 1508 -2679
rect 1598 -2713 1599 -2679
rect 1633 -2834 1634 -2712
rect 1647 -2834 1648 -2712
rect 1654 -2713 1655 -2679
rect 1668 -2713 1669 -2679
rect 1696 -2834 1697 -2712
rect 1766 -2834 1767 -2712
rect 2053 -2713 2054 -2679
rect 93 -2834 94 -2714
rect 114 -2715 115 -2679
rect 163 -2834 164 -2714
rect 352 -2715 353 -2679
rect 366 -2715 367 -2679
rect 660 -2834 661 -2714
rect 663 -2834 664 -2714
rect 1276 -2834 1277 -2714
rect 1388 -2715 1389 -2679
rect 1423 -2834 1424 -2714
rect 1430 -2715 1431 -2679
rect 1983 -2715 1984 -2679
rect 2053 -2834 2054 -2714
rect 2081 -2715 2082 -2679
rect 114 -2834 115 -2716
rect 478 -2717 479 -2679
rect 513 -2834 514 -2716
rect 1031 -2717 1032 -2679
rect 1073 -2717 1074 -2679
rect 1283 -2834 1284 -2716
rect 1395 -2834 1396 -2716
rect 2221 -2717 2222 -2679
rect 184 -2719 185 -2679
rect 1391 -2834 1392 -2718
rect 1398 -2719 1399 -2679
rect 2011 -2834 2012 -2718
rect 2060 -2719 2061 -2679
rect 2081 -2834 2082 -2718
rect 2221 -2834 2222 -2718
rect 2263 -2719 2264 -2679
rect 75 -2721 76 -2679
rect 184 -2834 185 -2720
rect 226 -2721 227 -2679
rect 387 -2834 388 -2720
rect 478 -2834 479 -2720
rect 856 -2721 857 -2679
rect 877 -2721 878 -2679
rect 1129 -2834 1130 -2720
rect 1227 -2834 1228 -2720
rect 1314 -2721 1315 -2679
rect 1433 -2721 1434 -2679
rect 2228 -2721 2229 -2679
rect 44 -2723 45 -2679
rect 856 -2834 857 -2722
rect 877 -2834 878 -2722
rect 1087 -2723 1088 -2679
rect 1097 -2834 1098 -2722
rect 2032 -2723 2033 -2679
rect 2060 -2834 2061 -2722
rect 2088 -2723 2089 -2679
rect 2214 -2723 2215 -2679
rect 2228 -2834 2229 -2722
rect 44 -2834 45 -2724
rect 471 -2725 472 -2679
rect 576 -2834 577 -2724
rect 646 -2725 647 -2679
rect 667 -2834 668 -2724
rect 702 -2725 703 -2679
rect 779 -2834 780 -2724
rect 849 -2725 850 -2679
rect 912 -2725 913 -2679
rect 1171 -2834 1172 -2724
rect 1262 -2834 1263 -2724
rect 1290 -2725 1291 -2679
rect 1437 -2725 1438 -2679
rect 1864 -2725 1865 -2679
rect 1962 -2725 1963 -2679
rect 1983 -2834 1984 -2724
rect 2088 -2834 2089 -2724
rect 2095 -2725 2096 -2679
rect 135 -2834 136 -2726
rect 912 -2834 913 -2726
rect 933 -2834 934 -2726
rect 1003 -2727 1004 -2679
rect 1010 -2727 1011 -2679
rect 1241 -2834 1242 -2726
rect 1244 -2727 1245 -2679
rect 1864 -2834 1865 -2726
rect 2095 -2834 2096 -2726
rect 2109 -2727 2110 -2679
rect 142 -2729 143 -2679
rect 646 -2834 647 -2728
rect 688 -2729 689 -2679
rect 1892 -2834 1893 -2728
rect 142 -2834 143 -2730
rect 170 -2731 171 -2679
rect 226 -2834 227 -2730
rect 331 -2731 332 -2679
rect 352 -2834 353 -2730
rect 541 -2731 542 -2679
rect 583 -2731 584 -2679
rect 583 -2834 584 -2730
rect 583 -2731 584 -2679
rect 583 -2834 584 -2730
rect 604 -2731 605 -2679
rect 1192 -2731 1193 -2679
rect 1269 -2834 1270 -2730
rect 1297 -2731 1298 -2679
rect 1437 -2834 1438 -2730
rect 1486 -2731 1487 -2679
rect 1500 -2731 1501 -2679
rect 1507 -2834 1508 -2730
rect 1528 -2731 1529 -2679
rect 1598 -2834 1599 -2730
rect 1626 -2731 1627 -2679
rect 1654 -2834 1655 -2730
rect 1668 -2834 1669 -2730
rect 1682 -2731 1683 -2679
rect 1780 -2731 1781 -2679
rect 2032 -2834 2033 -2730
rect 79 -2733 80 -2679
rect 604 -2834 605 -2732
rect 625 -2733 626 -2679
rect 758 -2834 759 -2732
rect 786 -2834 787 -2732
rect 2172 -2834 2173 -2732
rect 9 -2735 10 -2679
rect 79 -2834 80 -2734
rect 149 -2735 150 -2679
rect 331 -2834 332 -2734
rect 415 -2735 416 -2679
rect 1010 -2834 1011 -2734
rect 1073 -2834 1074 -2734
rect 1157 -2735 1158 -2679
rect 1192 -2834 1193 -2734
rect 1353 -2735 1354 -2679
rect 1440 -2735 1441 -2679
rect 2214 -2834 2215 -2734
rect 9 -2834 10 -2736
rect 863 -2737 864 -2679
rect 870 -2737 871 -2679
rect 1157 -2834 1158 -2736
rect 1290 -2834 1291 -2736
rect 1332 -2737 1333 -2679
rect 1353 -2834 1354 -2736
rect 1367 -2737 1368 -2679
rect 1472 -2737 1473 -2679
rect 2263 -2834 2264 -2736
rect 30 -2739 31 -2679
rect 415 -2834 416 -2738
rect 471 -2834 472 -2738
rect 492 -2739 493 -2679
rect 527 -2739 528 -2679
rect 863 -2834 864 -2738
rect 870 -2834 871 -2738
rect 1045 -2739 1046 -2679
rect 1087 -2834 1088 -2738
rect 1101 -2739 1102 -2679
rect 1108 -2739 1109 -2679
rect 1150 -2834 1151 -2738
rect 1332 -2834 1333 -2738
rect 2207 -2739 2208 -2679
rect 30 -2834 31 -2740
rect 254 -2741 255 -2679
rect 261 -2741 262 -2679
rect 359 -2834 360 -2740
rect 408 -2741 409 -2679
rect 1108 -2834 1109 -2740
rect 1115 -2741 1116 -2679
rect 1311 -2741 1312 -2679
rect 1314 -2834 1315 -2740
rect 2207 -2834 2208 -2740
rect 54 -2743 55 -2679
rect 1045 -2834 1046 -2742
rect 1101 -2834 1102 -2742
rect 1325 -2743 1326 -2679
rect 1367 -2834 1368 -2742
rect 1402 -2743 1403 -2679
rect 1451 -2743 1452 -2679
rect 1472 -2834 1473 -2742
rect 1521 -2743 1522 -2679
rect 1528 -2834 1529 -2742
rect 1580 -2743 1581 -2679
rect 1962 -2834 1963 -2742
rect 37 -2745 38 -2679
rect 1402 -2834 1403 -2744
rect 1521 -2834 1522 -2744
rect 1549 -2745 1550 -2679
rect 1626 -2834 1627 -2744
rect 1640 -2745 1641 -2679
rect 1850 -2745 1851 -2679
rect 2109 -2834 2110 -2744
rect 37 -2834 38 -2746
rect 450 -2747 451 -2679
rect 492 -2834 493 -2746
rect 726 -2747 727 -2679
rect 793 -2747 794 -2679
rect 842 -2834 843 -2746
rect 849 -2834 850 -2746
rect 1255 -2747 1256 -2679
rect 1549 -2834 1550 -2746
rect 1570 -2747 1571 -2679
rect 1689 -2747 1690 -2679
rect 1850 -2834 1851 -2746
rect 54 -2834 55 -2748
rect 1913 -2834 1914 -2748
rect 131 -2751 132 -2679
rect 149 -2834 150 -2750
rect 156 -2834 157 -2750
rect 1433 -2834 1434 -2750
rect 1570 -2834 1571 -2750
rect 1661 -2751 1662 -2679
rect 1689 -2834 1690 -2750
rect 1717 -2751 1718 -2679
rect 170 -2834 171 -2752
rect 317 -2753 318 -2679
rect 408 -2834 409 -2752
rect 422 -2753 423 -2679
rect 450 -2834 451 -2752
rect 597 -2753 598 -2679
rect 625 -2834 626 -2752
rect 964 -2834 965 -2752
rect 968 -2753 969 -2679
rect 1374 -2834 1375 -2752
rect 1542 -2753 1543 -2679
rect 1717 -2834 1718 -2752
rect 205 -2755 206 -2679
rect 254 -2834 255 -2754
rect 282 -2834 283 -2754
rect 310 -2755 311 -2679
rect 317 -2834 318 -2754
rect 443 -2755 444 -2679
rect 527 -2834 528 -2754
rect 751 -2755 752 -2679
rect 793 -2834 794 -2754
rect 1510 -2755 1511 -2679
rect 1542 -2834 1543 -2754
rect 1563 -2755 1564 -2679
rect 1661 -2834 1662 -2754
rect 1675 -2755 1676 -2679
rect 205 -2834 206 -2756
rect 1752 -2757 1753 -2679
rect 233 -2759 234 -2679
rect 261 -2834 262 -2758
rect 289 -2759 290 -2679
rect 366 -2834 367 -2758
rect 411 -2759 412 -2679
rect 1325 -2834 1326 -2758
rect 1675 -2834 1676 -2758
rect 1731 -2759 1732 -2679
rect 240 -2761 241 -2679
rect 1178 -2761 1179 -2679
rect 1255 -2834 1256 -2760
rect 1514 -2761 1515 -2679
rect 1731 -2834 1732 -2760
rect 1857 -2761 1858 -2679
rect 243 -2763 244 -2679
rect 401 -2763 402 -2679
rect 443 -2834 444 -2762
rect 705 -2834 706 -2762
rect 744 -2763 745 -2679
rect 968 -2834 969 -2762
rect 982 -2834 983 -2762
rect 1017 -2763 1018 -2679
rect 1059 -2763 1060 -2679
rect 1178 -2834 1179 -2762
rect 1514 -2834 1515 -2762
rect 1724 -2763 1725 -2679
rect 1857 -2834 1858 -2762
rect 1878 -2763 1879 -2679
rect 212 -2765 213 -2679
rect 401 -2834 402 -2764
rect 464 -2834 465 -2764
rect 1059 -2834 1060 -2764
rect 1115 -2834 1116 -2764
rect 1164 -2765 1165 -2679
rect 1724 -2834 1725 -2764
rect 1738 -2765 1739 -2679
rect 1878 -2834 1879 -2764
rect 2123 -2765 2124 -2679
rect 212 -2834 213 -2766
rect 303 -2767 304 -2679
rect 310 -2834 311 -2766
rect 590 -2767 591 -2679
rect 597 -2834 598 -2766
rect 1465 -2767 1466 -2679
rect 1738 -2834 1739 -2766
rect 1745 -2767 1746 -2679
rect 177 -2769 178 -2679
rect 590 -2834 591 -2768
rect 621 -2834 622 -2768
rect 751 -2834 752 -2768
rect 789 -2769 790 -2679
rect 2123 -2834 2124 -2768
rect 177 -2834 178 -2770
rect 898 -2771 899 -2679
rect 943 -2834 944 -2770
rect 1787 -2834 1788 -2770
rect 247 -2773 248 -2679
rect 303 -2834 304 -2772
rect 324 -2773 325 -2679
rect 422 -2834 423 -2772
rect 541 -2834 542 -2772
rect 1318 -2834 1319 -2772
rect 1465 -2834 1466 -2772
rect 1493 -2773 1494 -2679
rect 1496 -2834 1497 -2772
rect 1745 -2834 1746 -2772
rect 289 -2834 290 -2774
rect 569 -2775 570 -2679
rect 639 -2775 640 -2679
rect 716 -2834 717 -2774
rect 744 -2834 745 -2774
rect 1577 -2834 1578 -2774
rect 296 -2777 297 -2679
rect 324 -2834 325 -2776
rect 569 -2834 570 -2776
rect 674 -2777 675 -2679
rect 688 -2834 689 -2776
rect 940 -2777 941 -2679
rect 947 -2777 948 -2679
rect 1031 -2834 1032 -2776
rect 1122 -2777 1123 -2679
rect 1297 -2834 1298 -2776
rect 1493 -2834 1494 -2776
rect 1710 -2777 1711 -2679
rect 72 -2779 73 -2679
rect 296 -2834 297 -2778
rect 460 -2834 461 -2778
rect 1122 -2834 1123 -2778
rect 1125 -2779 1126 -2679
rect 1843 -2779 1844 -2679
rect 72 -2834 73 -2780
rect 236 -2834 237 -2780
rect 268 -2781 269 -2679
rect 674 -2834 675 -2780
rect 702 -2834 703 -2780
rect 1500 -2834 1501 -2780
rect 1710 -2834 1711 -2780
rect 1801 -2781 1802 -2679
rect 198 -2783 199 -2679
rect 947 -2834 948 -2782
rect 961 -2834 962 -2782
rect 2039 -2783 2040 -2679
rect 198 -2834 199 -2784
rect 1451 -2834 1452 -2784
rect 1794 -2785 1795 -2679
rect 1801 -2834 1802 -2784
rect 2039 -2834 2040 -2784
rect 2074 -2785 2075 -2679
rect 219 -2787 220 -2679
rect 268 -2834 269 -2786
rect 611 -2787 612 -2679
rect 639 -2834 640 -2786
rect 789 -2834 790 -2786
rect 1640 -2834 1641 -2786
rect 1794 -2834 1795 -2786
rect 1808 -2787 1809 -2679
rect 2074 -2834 2075 -2786
rect 2116 -2787 2117 -2679
rect 100 -2789 101 -2679
rect 611 -2834 612 -2788
rect 800 -2789 801 -2679
rect 1328 -2789 1329 -2679
rect 1703 -2789 1704 -2679
rect 1808 -2834 1809 -2788
rect 100 -2834 101 -2790
rect 247 -2834 248 -2790
rect 380 -2791 381 -2679
rect 800 -2834 801 -2790
rect 807 -2791 808 -2679
rect 2046 -2834 2047 -2790
rect 219 -2834 220 -2792
rect 898 -2834 899 -2792
rect 940 -2834 941 -2792
rect 1843 -2834 1844 -2792
rect 380 -2834 381 -2794
rect 618 -2795 619 -2679
rect 807 -2834 808 -2794
rect 828 -2795 829 -2679
rect 835 -2795 836 -2679
rect 922 -2795 923 -2679
rect 1003 -2834 1004 -2794
rect 1024 -2795 1025 -2679
rect 1164 -2834 1165 -2794
rect 1199 -2795 1200 -2679
rect 810 -2797 811 -2679
rect 2193 -2797 2194 -2679
rect 814 -2799 815 -2679
rect 1381 -2799 1382 -2679
rect 2186 -2799 2187 -2679
rect 2193 -2834 2194 -2798
rect 544 -2834 545 -2800
rect 2186 -2834 2187 -2800
rect 814 -2834 815 -2802
rect 884 -2803 885 -2679
rect 1017 -2834 1018 -2802
rect 1080 -2803 1081 -2679
rect 1199 -2834 1200 -2802
rect 1339 -2803 1340 -2679
rect 1381 -2834 1382 -2802
rect 1612 -2803 1613 -2679
rect 394 -2805 395 -2679
rect 884 -2834 885 -2804
rect 1024 -2834 1025 -2804
rect 1755 -2834 1756 -2804
rect 394 -2834 395 -2806
rect 457 -2834 458 -2806
rect 821 -2834 822 -2806
rect 905 -2807 906 -2679
rect 1080 -2834 1081 -2806
rect 1248 -2807 1249 -2679
rect 1339 -2834 1340 -2806
rect 1346 -2807 1347 -2679
rect 1409 -2807 1410 -2679
rect 1612 -2834 1613 -2806
rect 618 -2834 619 -2808
rect 1248 -2834 1249 -2808
rect 1346 -2834 1347 -2808
rect 1969 -2809 1970 -2679
rect 824 -2811 825 -2679
rect 1780 -2834 1781 -2810
rect 1969 -2834 1970 -2810
rect 1990 -2811 1991 -2679
rect 828 -2834 829 -2812
rect 1052 -2813 1053 -2679
rect 1409 -2834 1410 -2812
rect 1416 -2813 1417 -2679
rect 1815 -2813 1816 -2679
rect 1990 -2834 1991 -2812
rect 835 -2834 836 -2814
rect 926 -2815 927 -2679
rect 1052 -2834 1053 -2814
rect 1836 -2815 1837 -2679
rect 191 -2817 192 -2679
rect 926 -2834 927 -2816
rect 1815 -2834 1816 -2816
rect 1822 -2817 1823 -2679
rect 1836 -2834 1837 -2816
rect 1920 -2817 1921 -2679
rect 191 -2834 192 -2818
rect 534 -2819 535 -2679
rect 866 -2834 867 -2818
rect 2116 -2834 2117 -2818
rect 275 -2821 276 -2679
rect 534 -2834 535 -2820
rect 894 -2821 895 -2679
rect 1416 -2834 1417 -2820
rect 1535 -2821 1536 -2679
rect 1920 -2834 1921 -2820
rect 275 -2834 276 -2822
rect 499 -2823 500 -2679
rect 905 -2834 906 -2822
rect 1304 -2823 1305 -2679
rect 1822 -2834 1823 -2822
rect 1829 -2823 1830 -2679
rect 485 -2825 486 -2679
rect 499 -2834 500 -2824
rect 989 -2825 990 -2679
rect 1535 -2834 1536 -2824
rect 1829 -2834 1830 -2824
rect 1997 -2825 1998 -2679
rect 429 -2827 430 -2679
rect 485 -2834 486 -2826
rect 989 -2834 990 -2826
rect 1094 -2827 1095 -2679
rect 1304 -2834 1305 -2826
rect 1311 -2834 1312 -2826
rect 1997 -2834 1998 -2826
rect 2025 -2827 2026 -2679
rect 240 -2834 241 -2828
rect 1094 -2834 1095 -2828
rect 2025 -2834 2026 -2828
rect 2067 -2829 2068 -2679
rect 1941 -2831 1942 -2679
rect 2067 -2834 2068 -2830
rect 222 -2834 223 -2832
rect 1941 -2834 1942 -2832
rect 23 -2844 24 -2842
rect 467 -2979 468 -2843
rect 541 -2979 542 -2843
rect 1496 -2844 1497 -2842
rect 1500 -2844 1501 -2842
rect 2256 -2844 2257 -2842
rect 23 -2979 24 -2845
rect 184 -2846 185 -2842
rect 219 -2846 220 -2842
rect 380 -2846 381 -2842
rect 429 -2846 430 -2842
rect 492 -2846 493 -2842
rect 548 -2846 549 -2842
rect 786 -2979 787 -2845
rect 814 -2846 815 -2842
rect 940 -2846 941 -2842
rect 943 -2846 944 -2842
rect 1332 -2846 1333 -2842
rect 1346 -2846 1347 -2842
rect 1633 -2846 1634 -2842
rect 1682 -2846 1683 -2842
rect 2137 -2846 2138 -2842
rect 2144 -2846 2145 -2842
rect 2144 -2979 2145 -2845
rect 2144 -2846 2145 -2842
rect 2144 -2979 2145 -2845
rect 2221 -2846 2222 -2842
rect 2249 -2846 2250 -2842
rect 30 -2848 31 -2842
rect 544 -2848 545 -2842
rect 548 -2979 549 -2847
rect 891 -2848 892 -2842
rect 919 -2848 920 -2842
rect 1139 -2979 1140 -2847
rect 1202 -2979 1203 -2847
rect 1209 -2979 1210 -2847
rect 1255 -2979 1256 -2847
rect 1325 -2848 1326 -2842
rect 1332 -2979 1333 -2847
rect 1619 -2848 1620 -2842
rect 1682 -2979 1683 -2847
rect 2060 -2848 2061 -2842
rect 2074 -2848 2075 -2842
rect 2137 -2979 2138 -2847
rect 30 -2979 31 -2849
rect 257 -2979 258 -2849
rect 317 -2850 318 -2842
rect 789 -2850 790 -2842
rect 828 -2850 829 -2842
rect 891 -2979 892 -2849
rect 922 -2979 923 -2849
rect 1500 -2979 1501 -2849
rect 1566 -2850 1567 -2842
rect 2004 -2850 2005 -2842
rect 2060 -2979 2061 -2849
rect 2207 -2850 2208 -2842
rect 51 -2852 52 -2842
rect 478 -2852 479 -2842
rect 492 -2979 493 -2851
rect 527 -2852 528 -2842
rect 544 -2979 545 -2851
rect 912 -2852 913 -2842
rect 964 -2979 965 -2851
rect 1234 -2852 1235 -2842
rect 1258 -2852 1259 -2842
rect 1920 -2852 1921 -2842
rect 2004 -2979 2005 -2851
rect 2102 -2852 2103 -2842
rect 82 -2854 83 -2842
rect 408 -2854 409 -2842
rect 436 -2854 437 -2842
rect 436 -2979 437 -2853
rect 436 -2854 437 -2842
rect 436 -2979 437 -2853
rect 457 -2979 458 -2853
rect 499 -2854 500 -2842
rect 527 -2979 528 -2853
rect 737 -2854 738 -2842
rect 744 -2854 745 -2842
rect 842 -2854 843 -2842
rect 863 -2854 864 -2842
rect 1983 -2854 1984 -2842
rect 2074 -2979 2075 -2853
rect 2214 -2854 2215 -2842
rect 103 -2979 104 -2855
rect 352 -2856 353 -2842
rect 373 -2856 374 -2842
rect 408 -2979 409 -2855
rect 460 -2856 461 -2842
rect 555 -2856 556 -2842
rect 565 -2979 566 -2855
rect 940 -2979 941 -2855
rect 968 -2856 969 -2842
rect 971 -2864 972 -2855
rect 975 -2979 976 -2855
rect 1374 -2856 1375 -2842
rect 1391 -2856 1392 -2842
rect 1850 -2856 1851 -2842
rect 1983 -2979 1984 -2855
rect 2088 -2856 2089 -2842
rect 2098 -2979 2099 -2855
rect 2102 -2979 2103 -2855
rect 107 -2858 108 -2842
rect 387 -2858 388 -2842
rect 401 -2858 402 -2842
rect 814 -2979 815 -2857
rect 835 -2979 836 -2857
rect 926 -2858 927 -2842
rect 968 -2979 969 -2857
rect 982 -2858 983 -2842
rect 1017 -2858 1018 -2842
rect 1059 -2858 1060 -2842
rect 1062 -2979 1063 -2857
rect 1087 -2858 1088 -2842
rect 1136 -2858 1137 -2842
rect 1619 -2979 1620 -2857
rect 1703 -2858 1704 -2842
rect 2032 -2858 2033 -2842
rect 2088 -2979 2089 -2857
rect 2235 -2858 2236 -2842
rect 117 -2979 118 -2859
rect 1892 -2860 1893 -2842
rect 2032 -2979 2033 -2859
rect 2151 -2860 2152 -2842
rect 124 -2979 125 -2861
rect 856 -2862 857 -2842
rect 866 -2862 867 -2842
rect 1097 -2862 1098 -2842
rect 1234 -2979 1235 -2861
rect 1290 -2862 1291 -2842
rect 1314 -2862 1315 -2842
rect 1556 -2862 1557 -2842
rect 1703 -2979 1704 -2861
rect 1773 -2862 1774 -2842
rect 1850 -2979 1851 -2861
rect 1997 -2862 1998 -2842
rect 191 -2864 192 -2842
rect 401 -2979 402 -2863
rect 485 -2864 486 -2842
rect 555 -2979 556 -2863
rect 597 -2864 598 -2842
rect 660 -2864 661 -2842
rect 674 -2864 675 -2842
rect 926 -2979 927 -2863
rect 982 -2979 983 -2863
rect 1017 -2979 1018 -2863
rect 1136 -2979 1137 -2863
rect 1283 -2979 1284 -2863
rect 1381 -2864 1382 -2842
rect 1433 -2864 1434 -2842
rect 1717 -2864 1718 -2842
rect 1731 -2864 1732 -2842
rect 1920 -2979 1921 -2863
rect 128 -2866 129 -2842
rect 597 -2979 598 -2865
rect 611 -2866 612 -2842
rect 1125 -2979 1126 -2865
rect 1286 -2866 1287 -2842
rect 1696 -2866 1697 -2842
rect 1706 -2866 1707 -2842
rect 2018 -2866 2019 -2842
rect 86 -2868 87 -2842
rect 128 -2979 129 -2867
rect 191 -2979 192 -2867
rect 212 -2868 213 -2842
rect 219 -2979 220 -2867
rect 443 -2868 444 -2842
rect 485 -2979 486 -2867
rect 520 -2868 521 -2842
rect 583 -2868 584 -2842
rect 611 -2979 612 -2867
rect 621 -2868 622 -2842
rect 800 -2868 801 -2842
rect 856 -2979 857 -2867
rect 1241 -2868 1242 -2842
rect 1290 -2979 1291 -2867
rect 1339 -2868 1340 -2842
rect 1346 -2979 1347 -2867
rect 1472 -2868 1473 -2842
rect 1486 -2868 1487 -2842
rect 2109 -2868 2110 -2842
rect 86 -2979 87 -2869
rect 247 -2870 248 -2842
rect 250 -2870 251 -2842
rect 1402 -2870 1403 -2842
rect 1419 -2979 1420 -2869
rect 1472 -2979 1473 -2869
rect 1489 -2870 1490 -2842
rect 1633 -2979 1634 -2869
rect 1696 -2979 1697 -2869
rect 1815 -2870 1816 -2842
rect 1878 -2870 1879 -2842
rect 1997 -2979 1998 -2869
rect 2018 -2979 2019 -2869
rect 2123 -2870 2124 -2842
rect 72 -2872 73 -2842
rect 247 -2979 248 -2871
rect 289 -2872 290 -2842
rect 317 -2979 318 -2871
rect 324 -2872 325 -2842
rect 429 -2979 430 -2871
rect 443 -2979 444 -2871
rect 471 -2872 472 -2842
rect 499 -2979 500 -2871
rect 604 -2872 605 -2842
rect 674 -2979 675 -2871
rect 1311 -2872 1312 -2842
rect 1314 -2979 1315 -2871
rect 2200 -2872 2201 -2842
rect 58 -2874 59 -2842
rect 72 -2979 73 -2873
rect 135 -2874 136 -2842
rect 604 -2979 605 -2873
rect 681 -2874 682 -2842
rect 912 -2979 913 -2873
rect 1038 -2874 1039 -2842
rect 1349 -2874 1350 -2842
rect 1360 -2874 1361 -2842
rect 1363 -2979 1364 -2873
rect 1374 -2979 1375 -2873
rect 1423 -2874 1424 -2842
rect 1451 -2874 1452 -2842
rect 2193 -2874 2194 -2842
rect 58 -2979 59 -2875
rect 1248 -2876 1249 -2842
rect 1339 -2979 1340 -2875
rect 1367 -2876 1368 -2842
rect 1381 -2979 1382 -2875
rect 1437 -2876 1438 -2842
rect 1493 -2876 1494 -2842
rect 1685 -2876 1686 -2842
rect 1717 -2979 1718 -2875
rect 1857 -2876 1858 -2842
rect 1892 -2979 1893 -2875
rect 1976 -2876 1977 -2842
rect 2109 -2979 2110 -2875
rect 2242 -2876 2243 -2842
rect 100 -2878 101 -2842
rect 1367 -2979 1368 -2877
rect 1402 -2979 1403 -2877
rect 1409 -2878 1410 -2842
rect 1437 -2979 1438 -2877
rect 2270 -2878 2271 -2842
rect 100 -2979 101 -2879
rect 1731 -2979 1732 -2879
rect 1752 -2880 1753 -2842
rect 1906 -2880 1907 -2842
rect 1976 -2979 1977 -2879
rect 2179 -2880 2180 -2842
rect 110 -2979 111 -2881
rect 1409 -2979 1410 -2881
rect 1493 -2979 1494 -2881
rect 1542 -2882 1543 -2842
rect 1556 -2979 1557 -2881
rect 1640 -2882 1641 -2842
rect 1752 -2979 1753 -2881
rect 1871 -2882 1872 -2842
rect 1906 -2979 1907 -2881
rect 2011 -2882 2012 -2842
rect 2123 -2979 2124 -2881
rect 2224 -2882 2225 -2842
rect 135 -2979 136 -2883
rect 576 -2884 577 -2842
rect 583 -2979 584 -2883
rect 849 -2884 850 -2842
rect 880 -2979 881 -2883
rect 1101 -2884 1102 -2842
rect 1115 -2884 1116 -2842
rect 1423 -2979 1424 -2883
rect 1444 -2884 1445 -2842
rect 1542 -2979 1543 -2883
rect 1640 -2979 1641 -2883
rect 1759 -2884 1760 -2842
rect 1773 -2979 1774 -2883
rect 1885 -2884 1886 -2842
rect 2011 -2979 2012 -2883
rect 2116 -2884 2117 -2842
rect 65 -2886 66 -2842
rect 849 -2979 850 -2885
rect 961 -2886 962 -2842
rect 2116 -2979 2117 -2885
rect 205 -2888 206 -2842
rect 478 -2979 479 -2887
rect 520 -2979 521 -2887
rect 1052 -2888 1053 -2842
rect 1059 -2979 1060 -2887
rect 1458 -2888 1459 -2842
rect 1755 -2888 1756 -2842
rect 1990 -2888 1991 -2842
rect 2 -2890 3 -2842
rect 205 -2979 206 -2889
rect 212 -2979 213 -2889
rect 632 -2890 633 -2842
rect 642 -2979 643 -2889
rect 1451 -2979 1452 -2889
rect 1759 -2979 1760 -2889
rect 1829 -2890 1830 -2842
rect 1871 -2979 1872 -2889
rect 2259 -2890 2260 -2842
rect 222 -2892 223 -2842
rect 2046 -2892 2047 -2842
rect 233 -2894 234 -2842
rect 303 -2894 304 -2842
rect 310 -2894 311 -2842
rect 352 -2979 353 -2893
rect 373 -2979 374 -2893
rect 415 -2894 416 -2842
rect 576 -2979 577 -2893
rect 1416 -2894 1417 -2842
rect 1444 -2979 1445 -2893
rect 1479 -2894 1480 -2842
rect 1801 -2894 1802 -2842
rect 1878 -2979 1879 -2893
rect 1990 -2979 1991 -2893
rect 2095 -2894 2096 -2842
rect 233 -2979 234 -2895
rect 268 -2896 269 -2842
rect 289 -2979 290 -2895
rect 534 -2896 535 -2842
rect 590 -2896 591 -2842
rect 681 -2979 682 -2895
rect 688 -2896 689 -2842
rect 828 -2979 829 -2895
rect 961 -2979 962 -2895
rect 2151 -2979 2152 -2895
rect 163 -2898 164 -2842
rect 268 -2979 269 -2897
rect 275 -2898 276 -2842
rect 534 -2979 535 -2897
rect 590 -2979 591 -2897
rect 807 -2898 808 -2842
rect 978 -2898 979 -2842
rect 1885 -2979 1886 -2897
rect 2046 -2979 2047 -2897
rect 2165 -2898 2166 -2842
rect 163 -2979 164 -2899
rect 933 -2900 934 -2842
rect 1010 -2900 1011 -2842
rect 1458 -2979 1459 -2899
rect 1479 -2979 1480 -2899
rect 1598 -2900 1599 -2842
rect 1801 -2979 1802 -2899
rect 1941 -2900 1942 -2842
rect 236 -2902 237 -2842
rect 303 -2979 304 -2901
rect 310 -2979 311 -2901
rect 422 -2902 423 -2842
rect 632 -2979 633 -2901
rect 723 -2902 724 -2842
rect 730 -2902 731 -2842
rect 1388 -2902 1389 -2842
rect 1598 -2979 1599 -2901
rect 1612 -2902 1613 -2842
rect 1815 -2979 1816 -2901
rect 1836 -2902 1837 -2842
rect 1941 -2979 1942 -2901
rect 2039 -2902 2040 -2842
rect 16 -2904 17 -2842
rect 730 -2979 731 -2903
rect 744 -2979 745 -2903
rect 1073 -2904 1074 -2842
rect 1087 -2979 1088 -2903
rect 1122 -2904 1123 -2842
rect 1199 -2904 1200 -2842
rect 1857 -2979 1858 -2903
rect 2039 -2979 2040 -2903
rect 2158 -2904 2159 -2842
rect 37 -2906 38 -2842
rect 723 -2979 724 -2905
rect 747 -2906 748 -2842
rect 947 -2906 948 -2842
rect 954 -2906 955 -2842
rect 1122 -2979 1123 -2905
rect 1241 -2979 1242 -2905
rect 1297 -2906 1298 -2842
rect 1360 -2979 1361 -2905
rect 1521 -2906 1522 -2842
rect 1612 -2979 1613 -2905
rect 1675 -2906 1676 -2842
rect 1829 -2979 1830 -2905
rect 1948 -2906 1949 -2842
rect 37 -2979 38 -2907
rect 142 -2908 143 -2842
rect 275 -2979 276 -2907
rect 366 -2908 367 -2842
rect 380 -2979 381 -2907
rect 733 -2908 734 -2842
rect 737 -2979 738 -2907
rect 1675 -2979 1676 -2907
rect 1836 -2979 1837 -2907
rect 1913 -2908 1914 -2842
rect 142 -2979 143 -2909
rect 765 -2910 766 -2842
rect 772 -2910 773 -2842
rect 863 -2979 864 -2909
rect 933 -2979 934 -2909
rect 1094 -2910 1095 -2842
rect 1101 -2979 1102 -2909
rect 1143 -2910 1144 -2842
rect 1248 -2979 1249 -2909
rect 1276 -2910 1277 -2842
rect 1297 -2979 1298 -2909
rect 1395 -2910 1396 -2842
rect 1521 -2979 1522 -2909
rect 1626 -2910 1627 -2842
rect 1913 -2979 1914 -2909
rect 2025 -2910 2026 -2842
rect 324 -2979 325 -2911
rect 394 -2912 395 -2842
rect 415 -2979 416 -2911
rect 1055 -2912 1056 -2842
rect 1066 -2912 1067 -2842
rect 1325 -2979 1326 -2911
rect 1388 -2979 1389 -2911
rect 1465 -2912 1466 -2842
rect 2025 -2979 2026 -2911
rect 2130 -2912 2131 -2842
rect 44 -2914 45 -2842
rect 1066 -2979 1067 -2913
rect 1069 -2979 1070 -2913
rect 1654 -2914 1655 -2842
rect 2130 -2979 2131 -2913
rect 2263 -2914 2264 -2842
rect 44 -2979 45 -2915
rect 618 -2916 619 -2842
rect 646 -2916 647 -2842
rect 807 -2979 808 -2915
rect 842 -2979 843 -2915
rect 1199 -2979 1200 -2915
rect 1276 -2979 1277 -2915
rect 1353 -2916 1354 -2842
rect 1395 -2979 1396 -2915
rect 1507 -2916 1508 -2842
rect 1654 -2979 1655 -2915
rect 1689 -2916 1690 -2842
rect 9 -2918 10 -2842
rect 618 -2979 619 -2917
rect 660 -2979 661 -2917
rect 1626 -2979 1627 -2917
rect 1689 -2979 1690 -2917
rect 1745 -2918 1746 -2842
rect 198 -2920 199 -2842
rect 394 -2979 395 -2919
rect 422 -2979 423 -2919
rect 464 -2920 465 -2842
rect 562 -2920 563 -2842
rect 646 -2979 647 -2919
rect 663 -2920 664 -2842
rect 947 -2979 948 -2919
rect 954 -2979 955 -2919
rect 1038 -2979 1039 -2919
rect 1045 -2920 1046 -2842
rect 1486 -2979 1487 -2919
rect 1507 -2979 1508 -2919
rect 1591 -2920 1592 -2842
rect 1745 -2979 1746 -2919
rect 1864 -2920 1865 -2842
rect 65 -2979 66 -2921
rect 464 -2979 465 -2921
rect 506 -2922 507 -2842
rect 562 -2979 563 -2921
rect 663 -2979 664 -2921
rect 1178 -2922 1179 -2842
rect 1465 -2979 1466 -2921
rect 1577 -2922 1578 -2842
rect 1710 -2922 1711 -2842
rect 1864 -2979 1865 -2921
rect 121 -2924 122 -2842
rect 506 -2979 507 -2923
rect 688 -2979 689 -2923
rect 1171 -2924 1172 -2842
rect 1178 -2979 1179 -2923
rect 1304 -2924 1305 -2842
rect 1430 -2924 1431 -2842
rect 1577 -2979 1578 -2923
rect 1710 -2979 1711 -2923
rect 1794 -2924 1795 -2842
rect 121 -2979 122 -2925
rect 184 -2979 185 -2925
rect 331 -2926 332 -2842
rect 471 -2979 472 -2925
rect 702 -2926 703 -2842
rect 1157 -2926 1158 -2842
rect 1171 -2979 1172 -2925
rect 1213 -2926 1214 -2842
rect 1304 -2979 1305 -2925
rect 1843 -2926 1844 -2842
rect 149 -2928 150 -2842
rect 198 -2979 199 -2927
rect 240 -2928 241 -2842
rect 331 -2979 332 -2927
rect 345 -2928 346 -2842
rect 366 -2979 367 -2927
rect 387 -2979 388 -2927
rect 1055 -2979 1056 -2927
rect 1073 -2979 1074 -2927
rect 1129 -2928 1130 -2842
rect 1213 -2979 1214 -2927
rect 1262 -2928 1263 -2842
rect 1430 -2979 1431 -2927
rect 1528 -2928 1529 -2842
rect 1570 -2928 1571 -2842
rect 1591 -2979 1592 -2927
rect 1794 -2979 1795 -2927
rect 1955 -2928 1956 -2842
rect 149 -2979 150 -2929
rect 1024 -2930 1025 -2842
rect 1031 -2930 1032 -2842
rect 1045 -2979 1046 -2929
rect 1080 -2930 1081 -2842
rect 1353 -2979 1354 -2929
rect 1528 -2979 1529 -2929
rect 1584 -2930 1585 -2842
rect 1843 -2979 1844 -2929
rect 1962 -2930 1963 -2842
rect 156 -2932 157 -2842
rect 240 -2979 241 -2931
rect 345 -2979 346 -2931
rect 793 -2932 794 -2842
rect 989 -2932 990 -2842
rect 1024 -2979 1025 -2931
rect 1080 -2979 1081 -2931
rect 1661 -2932 1662 -2842
rect 1955 -2979 1956 -2931
rect 2067 -2932 2068 -2842
rect 513 -2934 514 -2842
rect 1129 -2979 1130 -2933
rect 1192 -2934 1193 -2842
rect 1262 -2979 1263 -2933
rect 1514 -2934 1515 -2842
rect 1584 -2979 1585 -2933
rect 1661 -2979 1662 -2933
rect 1738 -2934 1739 -2842
rect 1962 -2979 1963 -2933
rect 2081 -2934 2082 -2842
rect 296 -2936 297 -2842
rect 513 -2979 514 -2935
rect 569 -2936 570 -2842
rect 702 -2979 703 -2935
rect 705 -2936 706 -2842
rect 884 -2936 885 -2842
rect 989 -2979 990 -2935
rect 1031 -2979 1032 -2935
rect 1094 -2979 1095 -2935
rect 1143 -2979 1144 -2935
rect 1192 -2979 1193 -2935
rect 1269 -2936 1270 -2842
rect 1514 -2979 1515 -2935
rect 1605 -2936 1606 -2842
rect 1738 -2979 1739 -2935
rect 2095 -2979 2096 -2935
rect 54 -2979 55 -2937
rect 1269 -2979 1270 -2937
rect 1605 -2979 1606 -2937
rect 1668 -2938 1669 -2842
rect 2067 -2979 2068 -2937
rect 2186 -2938 2187 -2842
rect 170 -2940 171 -2842
rect 569 -2979 570 -2939
rect 709 -2940 710 -2842
rect 884 -2979 885 -2939
rect 1010 -2979 1011 -2939
rect 1206 -2940 1207 -2842
rect 1668 -2979 1669 -2939
rect 1787 -2940 1788 -2842
rect 2081 -2979 2082 -2939
rect 2228 -2940 2229 -2842
rect 170 -2979 171 -2941
rect 261 -2942 262 -2842
rect 296 -2979 297 -2941
rect 338 -2942 339 -2842
rect 695 -2942 696 -2842
rect 709 -2979 710 -2941
rect 740 -2979 741 -2941
rect 1948 -2979 1949 -2941
rect 254 -2944 255 -2842
rect 338 -2979 339 -2943
rect 667 -2944 668 -2842
rect 695 -2979 696 -2943
rect 751 -2944 752 -2842
rect 1563 -2944 1564 -2842
rect 1787 -2979 1788 -2943
rect 1934 -2944 1935 -2842
rect 16 -2979 17 -2945
rect 254 -2979 255 -2945
rect 261 -2979 262 -2945
rect 359 -2946 360 -2842
rect 667 -2979 668 -2945
rect 1570 -2979 1571 -2945
rect 177 -2948 178 -2842
rect 751 -2979 752 -2947
rect 765 -2979 766 -2947
rect 1150 -2948 1151 -2842
rect 1157 -2979 1158 -2947
rect 1934 -2979 1935 -2947
rect 177 -2979 178 -2949
rect 215 -2979 216 -2949
rect 226 -2950 227 -2842
rect 359 -2979 360 -2949
rect 772 -2979 773 -2949
rect 1003 -2950 1004 -2842
rect 1115 -2979 1116 -2949
rect 1164 -2950 1165 -2842
rect 1206 -2979 1207 -2949
rect 1535 -2950 1536 -2842
rect 1563 -2979 1564 -2949
rect 1647 -2950 1648 -2842
rect 159 -2979 160 -2951
rect 226 -2979 227 -2951
rect 779 -2952 780 -2842
rect 800 -2979 801 -2951
rect 870 -2952 871 -2842
rect 1003 -2979 1004 -2951
rect 1150 -2979 1151 -2951
rect 1185 -2952 1186 -2842
rect 1535 -2979 1536 -2951
rect 1724 -2952 1725 -2842
rect 779 -2979 780 -2953
rect 877 -2954 878 -2842
rect 905 -2954 906 -2842
rect 1164 -2979 1165 -2953
rect 1185 -2979 1186 -2953
rect 1220 -2954 1221 -2842
rect 1647 -2979 1648 -2953
rect 1780 -2954 1781 -2842
rect 93 -2956 94 -2842
rect 905 -2979 906 -2955
rect 1097 -2979 1098 -2955
rect 1220 -2979 1221 -2955
rect 1724 -2979 1725 -2955
rect 1822 -2956 1823 -2842
rect 79 -2958 80 -2842
rect 93 -2979 94 -2957
rect 793 -2979 794 -2957
rect 821 -2958 822 -2842
rect 870 -2979 871 -2957
rect 898 -2958 899 -2842
rect 1780 -2979 1781 -2957
rect 1927 -2958 1928 -2842
rect 79 -2979 80 -2959
rect 996 -2960 997 -2842
rect 1822 -2979 1823 -2959
rect 1969 -2960 1970 -2842
rect 114 -2962 115 -2842
rect 898 -2979 899 -2961
rect 996 -2979 997 -2961
rect 1108 -2962 1109 -2842
rect 1927 -2979 1928 -2961
rect 2053 -2962 2054 -2842
rect 114 -2979 115 -2963
rect 450 -2964 451 -2842
rect 758 -2964 759 -2842
rect 821 -2979 822 -2963
rect 1108 -2979 1109 -2963
rect 1227 -2964 1228 -2842
rect 1808 -2964 1809 -2842
rect 2053 -2979 2054 -2963
rect 450 -2979 451 -2965
rect 1041 -2979 1042 -2965
rect 1227 -2979 1228 -2965
rect 1318 -2966 1319 -2842
rect 1808 -2979 1809 -2965
rect 1899 -2966 1900 -2842
rect 1969 -2979 1970 -2965
rect 2172 -2966 2173 -2842
rect 653 -2968 654 -2842
rect 758 -2979 759 -2967
rect 1318 -2979 1319 -2967
rect 1549 -2968 1550 -2842
rect 1766 -2968 1767 -2842
rect 1899 -2979 1900 -2967
rect 639 -2970 640 -2842
rect 653 -2979 654 -2969
rect 1160 -2979 1161 -2969
rect 1549 -2979 1550 -2969
rect 282 -2972 283 -2842
rect 639 -2979 640 -2971
rect 282 -2979 283 -2973
rect 625 -2974 626 -2842
rect 625 -2979 626 -2975
rect 716 -2976 717 -2842
rect 716 -2979 717 -2977
rect 985 -2979 986 -2977
rect 16 -2989 17 -2987
rect 110 -2989 111 -2987
rect 114 -3094 115 -2988
rect 387 -2989 388 -2987
rect 422 -2989 423 -2987
rect 460 -3094 461 -2988
rect 471 -2989 472 -2987
rect 562 -3094 563 -2988
rect 569 -2989 570 -2987
rect 975 -2989 976 -2987
rect 1041 -2989 1042 -2987
rect 2060 -2989 2061 -2987
rect 2095 -2989 2096 -2987
rect 2137 -2989 2138 -2987
rect 51 -2991 52 -2987
rect 72 -2991 73 -2987
rect 100 -2991 101 -2987
rect 933 -2991 934 -2987
rect 961 -2991 962 -2987
rect 968 -2991 969 -2987
rect 1052 -2991 1053 -2987
rect 1325 -2991 1326 -2987
rect 1346 -2991 1347 -2987
rect 1346 -3094 1347 -2990
rect 1346 -2991 1347 -2987
rect 1346 -3094 1347 -2990
rect 1360 -3094 1361 -2990
rect 1409 -2991 1410 -2987
rect 1416 -2991 1417 -2987
rect 1857 -2991 1858 -2987
rect 1871 -2991 1872 -2987
rect 1874 -2991 1875 -2987
rect 2098 -2991 2099 -2987
rect 2116 -2991 2117 -2987
rect 37 -2993 38 -2987
rect 72 -3094 73 -2992
rect 93 -2993 94 -2987
rect 100 -3094 101 -2992
rect 107 -3094 108 -2992
rect 779 -2993 780 -2987
rect 880 -2993 881 -2987
rect 1689 -2993 1690 -2987
rect 1769 -2993 1770 -2987
rect 1815 -2993 1816 -2987
rect 1836 -2993 1837 -2987
rect 1857 -3094 1858 -2992
rect 1871 -3094 1872 -2992
rect 1990 -2993 1991 -2987
rect 30 -2995 31 -2987
rect 93 -3094 94 -2994
rect 142 -2995 143 -2987
rect 919 -2995 920 -2987
rect 964 -2995 965 -2987
rect 1031 -2995 1032 -2987
rect 1055 -2995 1056 -2987
rect 1836 -3094 1837 -2994
rect 1892 -2995 1893 -2987
rect 1990 -3094 1991 -2994
rect 30 -3094 31 -2996
rect 58 -2997 59 -2987
rect 65 -2997 66 -2987
rect 565 -2997 566 -2987
rect 572 -2997 573 -2987
rect 961 -3094 962 -2996
rect 968 -3094 969 -2996
rect 1087 -2997 1088 -2987
rect 1125 -2997 1126 -2987
rect 1493 -2997 1494 -2987
rect 1566 -3094 1567 -2996
rect 1885 -2997 1886 -2987
rect 37 -3094 38 -2998
rect 520 -2999 521 -2987
rect 541 -2999 542 -2987
rect 814 -2999 815 -2987
rect 884 -2999 885 -2987
rect 933 -3094 934 -2998
rect 1031 -3094 1032 -2998
rect 1185 -2999 1186 -2987
rect 1199 -2999 1200 -2987
rect 1976 -2999 1977 -2987
rect 44 -3001 45 -2987
rect 65 -3094 66 -3000
rect 135 -3001 136 -2987
rect 541 -3094 542 -3000
rect 590 -3001 591 -2987
rect 915 -3094 916 -3000
rect 954 -3001 955 -2987
rect 1185 -3094 1186 -3000
rect 1199 -3094 1200 -3000
rect 1248 -3001 1249 -2987
rect 1318 -3001 1319 -2987
rect 1416 -3094 1417 -3000
rect 1419 -3001 1420 -2987
rect 1920 -3001 1921 -2987
rect 1976 -3094 1977 -3000
rect 2102 -3001 2103 -2987
rect 58 -3094 59 -3002
rect 198 -3003 199 -2987
rect 208 -3094 209 -3002
rect 443 -3003 444 -2987
rect 471 -3094 472 -3002
rect 880 -3094 881 -3002
rect 894 -3094 895 -3002
rect 1878 -3003 1879 -2987
rect 1885 -3094 1886 -3002
rect 1983 -3003 1984 -2987
rect 142 -3094 143 -3004
rect 205 -3005 206 -2987
rect 212 -3005 213 -2987
rect 338 -3005 339 -2987
rect 422 -3094 423 -3004
rect 429 -3005 430 -2987
rect 436 -3005 437 -2987
rect 436 -3094 437 -3004
rect 436 -3005 437 -2987
rect 436 -3094 437 -3004
rect 443 -3094 444 -3004
rect 1276 -3005 1277 -2987
rect 1318 -3094 1319 -3004
rect 1339 -3005 1340 -2987
rect 1398 -3094 1399 -3004
rect 1941 -3005 1942 -2987
rect 86 -3007 87 -2987
rect 212 -3094 213 -3006
rect 236 -3094 237 -3006
rect 618 -3007 619 -2987
rect 642 -3007 643 -2987
rect 758 -3007 759 -2987
rect 786 -3007 787 -2987
rect 954 -3094 955 -3006
rect 1055 -3094 1056 -3006
rect 1703 -3007 1704 -2987
rect 1808 -3007 1809 -2987
rect 1881 -3094 1882 -3006
rect 1920 -3094 1921 -3006
rect 2025 -3007 2026 -2987
rect 86 -3094 87 -3008
rect 219 -3009 220 -2987
rect 240 -3009 241 -2987
rect 429 -3094 430 -3008
rect 478 -3009 479 -2987
rect 618 -3094 619 -3008
rect 688 -3009 689 -2987
rect 1038 -3009 1039 -2987
rect 1066 -3009 1067 -2987
rect 1094 -3094 1095 -3008
rect 1139 -3009 1140 -2987
rect 1633 -3009 1634 -2987
rect 1654 -3009 1655 -2987
rect 1941 -3094 1942 -3008
rect 131 -3094 132 -3010
rect 786 -3094 787 -3010
rect 905 -3011 906 -2987
rect 919 -3094 920 -3010
rect 1038 -3094 1039 -3010
rect 1220 -3011 1221 -2987
rect 1325 -3094 1326 -3010
rect 1559 -3094 1560 -3010
rect 1570 -3011 1571 -2987
rect 1864 -3011 1865 -2987
rect 149 -3013 150 -2987
rect 464 -3094 465 -3012
rect 478 -3094 479 -3012
rect 667 -3013 668 -2987
rect 688 -3094 689 -3012
rect 1255 -3013 1256 -2987
rect 1339 -3094 1340 -3012
rect 1430 -3013 1431 -2987
rect 1486 -3013 1487 -2987
rect 1766 -3013 1767 -2987
rect 1808 -3094 1809 -3012
rect 2053 -3013 2054 -2987
rect 138 -3094 139 -3014
rect 149 -3094 150 -3014
rect 156 -3015 157 -2987
rect 663 -3015 664 -2987
rect 667 -3094 668 -3014
rect 695 -3015 696 -2987
rect 716 -3015 717 -2987
rect 719 -3021 720 -3014
rect 730 -3015 731 -2987
rect 922 -3015 923 -2987
rect 1045 -3015 1046 -2987
rect 1066 -3094 1067 -3014
rect 1069 -3015 1070 -2987
rect 1213 -3015 1214 -2987
rect 1220 -3094 1221 -3014
rect 1227 -3015 1228 -2987
rect 1255 -3094 1256 -3014
rect 1269 -3015 1270 -2987
rect 1402 -3015 1403 -2987
rect 1405 -3094 1406 -3014
rect 1430 -3094 1431 -3014
rect 1500 -3015 1501 -2987
rect 1570 -3094 1571 -3014
rect 1605 -3015 1606 -2987
rect 1633 -3094 1634 -3014
rect 1675 -3015 1676 -2987
rect 1689 -3094 1690 -3014
rect 1773 -3015 1774 -2987
rect 1815 -3094 1816 -3014
rect 1948 -3015 1949 -2987
rect 156 -3094 157 -3016
rect 191 -3017 192 -2987
rect 198 -3094 199 -3016
rect 261 -3017 262 -2987
rect 282 -3017 283 -2987
rect 569 -3094 570 -3016
rect 590 -3094 591 -3016
rect 702 -3017 703 -2987
rect 716 -3094 717 -3016
rect 849 -3017 850 -2987
rect 905 -3094 906 -3016
rect 1045 -3094 1046 -3016
rect 1143 -3017 1144 -2987
rect 1160 -3017 1161 -2987
rect 1353 -3017 1354 -2987
rect 1402 -3094 1403 -3016
rect 1528 -3017 1529 -2987
rect 1549 -3017 1550 -2987
rect 1675 -3094 1676 -3016
rect 1703 -3094 1704 -3016
rect 1780 -3017 1781 -2987
rect 1864 -3094 1865 -3016
rect 2039 -3017 2040 -2987
rect 128 -3019 129 -2987
rect 1160 -3094 1161 -3018
rect 1178 -3019 1179 -2987
rect 1206 -3094 1207 -3018
rect 1213 -3094 1214 -3018
rect 1423 -3019 1424 -2987
rect 1486 -3094 1487 -3018
rect 1563 -3019 1564 -2987
rect 1573 -3019 1574 -2987
rect 2130 -3019 2131 -2987
rect 159 -3021 160 -2987
rect 1073 -3021 1074 -2987
rect 1076 -3094 1077 -3020
rect 1437 -3021 1438 -2987
rect 1493 -3094 1494 -3020
rect 1521 -3021 1522 -2987
rect 1528 -3094 1529 -3020
rect 1682 -3021 1683 -2987
rect 1759 -3021 1760 -2987
rect 1780 -3094 1781 -3020
rect 1874 -3094 1875 -3020
rect 1892 -3094 1893 -3020
rect 1948 -3094 1949 -3020
rect 2088 -3021 2089 -2987
rect 163 -3023 164 -2987
rect 520 -3094 521 -3022
rect 597 -3023 598 -2987
rect 639 -3094 640 -3022
rect 695 -3094 696 -3022
rect 709 -3023 710 -2987
rect 730 -3094 731 -3022
rect 1080 -3023 1081 -2987
rect 1083 -3094 1084 -3022
rect 1934 -3023 1935 -2987
rect 166 -3094 167 -3024
rect 926 -3025 927 -2987
rect 1087 -3094 1088 -3024
rect 1115 -3025 1116 -2987
rect 1143 -3094 1144 -3024
rect 1304 -3025 1305 -2987
rect 1353 -3094 1354 -3024
rect 1395 -3025 1396 -2987
rect 1423 -3094 1424 -3024
rect 1479 -3025 1480 -2987
rect 1500 -3094 1501 -3024
rect 1556 -3025 1557 -2987
rect 1654 -3094 1655 -3024
rect 1745 -3025 1746 -2987
rect 1759 -3094 1760 -3024
rect 1850 -3025 1851 -2987
rect 1934 -3094 1935 -3024
rect 2011 -3025 2012 -2987
rect 79 -3027 80 -2987
rect 926 -3094 927 -3026
rect 985 -3027 986 -2987
rect 1850 -3094 1851 -3026
rect 170 -3029 171 -2987
rect 261 -3094 262 -3028
rect 282 -3094 283 -3028
rect 380 -3029 381 -2987
rect 457 -3029 458 -2987
rect 597 -3094 598 -3028
rect 614 -3094 615 -3028
rect 898 -3029 899 -2987
rect 1178 -3094 1179 -3028
rect 1241 -3029 1242 -2987
rect 1269 -3094 1270 -3028
rect 1290 -3029 1291 -2987
rect 1304 -3094 1305 -3028
rect 1472 -3029 1473 -2987
rect 1549 -3094 1550 -3028
rect 1612 -3029 1613 -2987
rect 1661 -3029 1662 -2987
rect 1685 -3094 1686 -3028
rect 1745 -3094 1746 -3028
rect 1955 -3029 1956 -2987
rect 173 -3094 174 -3030
rect 604 -3031 605 -2987
rect 625 -3031 626 -2987
rect 1115 -3094 1116 -3030
rect 1192 -3031 1193 -2987
rect 1605 -3094 1606 -3030
rect 1612 -3094 1613 -3030
rect 1640 -3031 1641 -2987
rect 1661 -3094 1662 -3030
rect 1724 -3031 1725 -2987
rect 1766 -3094 1767 -3030
rect 1843 -3031 1844 -2987
rect 184 -3033 185 -2987
rect 191 -3094 192 -3032
rect 219 -3094 220 -3032
rect 373 -3033 374 -2987
rect 457 -3094 458 -3032
rect 975 -3094 976 -3032
rect 1164 -3033 1165 -2987
rect 1192 -3094 1193 -3032
rect 1202 -3033 1203 -2987
rect 1409 -3094 1410 -3032
rect 1437 -3094 1438 -3032
rect 1514 -3033 1515 -2987
rect 1598 -3033 1599 -2987
rect 1640 -3094 1641 -3032
rect 1682 -3094 1683 -3032
rect 1983 -3094 1984 -3032
rect 184 -3094 185 -3034
rect 205 -3094 206 -3034
rect 215 -3035 216 -2987
rect 373 -3094 374 -3034
rect 485 -3035 486 -2987
rect 737 -3035 738 -2987
rect 740 -3035 741 -2987
rect 870 -3035 871 -2987
rect 1136 -3035 1137 -2987
rect 1598 -3094 1599 -3034
rect 1724 -3094 1725 -3034
rect 2074 -3035 2075 -2987
rect 240 -3094 241 -3036
rect 268 -3037 269 -2987
rect 296 -3037 297 -2987
rect 660 -3037 661 -2987
rect 702 -3094 703 -3036
rect 723 -3037 724 -2987
rect 737 -3094 738 -3036
rect 912 -3037 913 -2987
rect 1136 -3094 1137 -3036
rect 1234 -3037 1235 -2987
rect 1241 -3094 1242 -3036
rect 1388 -3037 1389 -2987
rect 1451 -3037 1452 -2987
rect 1521 -3094 1522 -3036
rect 1773 -3094 1774 -3036
rect 1822 -3037 1823 -2987
rect 1843 -3094 1844 -3036
rect 2004 -3037 2005 -2987
rect 2074 -3094 2075 -3036
rect 2151 -3037 2152 -2987
rect 254 -3039 255 -2987
rect 1367 -3039 1368 -2987
rect 1388 -3094 1389 -3038
rect 1717 -3039 1718 -2987
rect 1822 -3094 1823 -3038
rect 2018 -3039 2019 -2987
rect 247 -3041 248 -2987
rect 254 -3094 255 -3040
rect 268 -3094 269 -3040
rect 1059 -3041 1060 -2987
rect 1157 -3041 1158 -2987
rect 1367 -3094 1368 -3040
rect 1451 -3094 1452 -3040
rect 1731 -3041 1732 -2987
rect 2004 -3094 2005 -3040
rect 2081 -3041 2082 -2987
rect 103 -3043 104 -2987
rect 247 -3094 248 -3042
rect 296 -3094 297 -3042
rect 401 -3043 402 -2987
rect 415 -3043 416 -2987
rect 723 -3094 724 -3042
rect 758 -3094 759 -3042
rect 817 -3094 818 -3042
rect 870 -3094 871 -3042
rect 947 -3043 948 -2987
rect 1017 -3043 1018 -2987
rect 1731 -3094 1732 -3042
rect 275 -3045 276 -2987
rect 401 -3094 402 -3044
rect 415 -3094 416 -3044
rect 506 -3045 507 -2987
rect 513 -3045 514 -2987
rect 779 -3094 780 -3044
rect 835 -3045 836 -2987
rect 947 -3094 948 -3044
rect 1003 -3045 1004 -2987
rect 1017 -3094 1018 -3044
rect 1059 -3094 1060 -3044
rect 1101 -3045 1102 -2987
rect 1164 -3094 1165 -3044
rect 1237 -3094 1238 -3044
rect 1283 -3045 1284 -2987
rect 1290 -3094 1291 -3044
rect 1332 -3045 1333 -2987
rect 1479 -3094 1480 -3044
rect 1514 -3094 1515 -3044
rect 1542 -3045 1543 -2987
rect 1717 -3094 1718 -3044
rect 1794 -3045 1795 -2987
rect 275 -3094 276 -3046
rect 324 -3047 325 -2987
rect 338 -3094 339 -3046
rect 366 -3047 367 -2987
rect 485 -3094 486 -3046
rect 555 -3047 556 -2987
rect 625 -3094 626 -3046
rect 674 -3047 675 -2987
rect 709 -3094 710 -3046
rect 1062 -3047 1063 -2987
rect 1097 -3047 1098 -2987
rect 1332 -3094 1333 -3046
rect 1465 -3047 1466 -2987
rect 1955 -3094 1956 -3046
rect 289 -3049 290 -2987
rect 555 -3094 556 -3048
rect 660 -3094 661 -3048
rect 681 -3049 682 -2987
rect 765 -3049 766 -2987
rect 849 -3094 850 -3048
rect 884 -3094 885 -3048
rect 1234 -3094 1235 -3048
rect 1283 -3094 1284 -3048
rect 1297 -3049 1298 -2987
rect 1465 -3094 1466 -3048
rect 1738 -3049 1739 -2987
rect 1794 -3094 1795 -3048
rect 1927 -3049 1928 -2987
rect 289 -3094 290 -3050
rect 632 -3051 633 -2987
rect 674 -3094 675 -3050
rect 1129 -3051 1130 -2987
rect 1227 -3094 1228 -3050
rect 1262 -3051 1263 -2987
rect 1297 -3094 1298 -3050
rect 1311 -3051 1312 -2987
rect 1472 -3094 1473 -3050
rect 1965 -3094 1966 -3050
rect 310 -3053 311 -2987
rect 387 -3094 388 -3052
rect 506 -3094 507 -3052
rect 996 -3053 997 -2987
rect 1024 -3053 1025 -2987
rect 1262 -3094 1263 -3052
rect 1311 -3094 1312 -3052
rect 1535 -3053 1536 -2987
rect 1542 -3094 1543 -3052
rect 1584 -3053 1585 -2987
rect 1738 -3094 1739 -3052
rect 1801 -3053 1802 -2987
rect 1927 -3094 1928 -3052
rect 2067 -3053 2068 -2987
rect 310 -3094 311 -3054
rect 1073 -3094 1074 -3054
rect 1101 -3094 1102 -3054
rect 1150 -3055 1151 -2987
rect 1535 -3094 1536 -3054
rect 1591 -3055 1592 -2987
rect 1801 -3094 1802 -3054
rect 1906 -3055 1907 -2987
rect 324 -3094 325 -3056
rect 499 -3057 500 -2987
rect 513 -3094 514 -3056
rect 534 -3057 535 -2987
rect 548 -3057 549 -2987
rect 1157 -3094 1158 -3056
rect 1584 -3094 1585 -3056
rect 1619 -3057 1620 -2987
rect 1906 -3094 1907 -3056
rect 2032 -3057 2033 -2987
rect 226 -3059 227 -2987
rect 534 -3094 535 -3058
rect 632 -3094 633 -3058
rect 828 -3059 829 -2987
rect 835 -3094 836 -3058
rect 1381 -3059 1382 -2987
rect 1591 -3094 1592 -3058
rect 1626 -3059 1627 -2987
rect 2032 -3094 2033 -3058
rect 2109 -3059 2110 -2987
rect 121 -3061 122 -2987
rect 226 -3094 227 -3060
rect 352 -3061 353 -2987
rect 548 -3094 549 -3060
rect 681 -3094 682 -3060
rect 842 -3061 843 -2987
rect 940 -3061 941 -2987
rect 1003 -3094 1004 -3060
rect 1024 -3094 1025 -3060
rect 1108 -3061 1109 -2987
rect 1122 -3094 1123 -3060
rect 1150 -3094 1151 -3060
rect 1381 -3094 1382 -3060
rect 1444 -3061 1445 -2987
rect 1619 -3094 1620 -3060
rect 1647 -3061 1648 -2987
rect 121 -3094 122 -3062
rect 576 -3063 577 -2987
rect 765 -3094 766 -3062
rect 856 -3063 857 -2987
rect 940 -3094 941 -3062
rect 1374 -3063 1375 -2987
rect 1626 -3094 1627 -3062
rect 1696 -3063 1697 -2987
rect 124 -3065 125 -2987
rect 352 -3094 353 -3064
rect 359 -3065 360 -2987
rect 380 -3094 381 -3064
rect 450 -3065 451 -2987
rect 828 -3094 829 -3064
rect 856 -3094 857 -3064
rect 863 -3065 864 -2987
rect 996 -3094 997 -3064
rect 1216 -3094 1217 -3064
rect 1556 -3094 1557 -3064
rect 1696 -3094 1697 -3064
rect 359 -3094 360 -3066
rect 544 -3067 545 -2987
rect 576 -3094 577 -3066
rect 653 -3067 654 -2987
rect 772 -3067 773 -2987
rect 898 -3094 899 -3066
rect 1010 -3067 1011 -2987
rect 1108 -3094 1109 -3066
rect 1129 -3094 1130 -3066
rect 1171 -3067 1172 -2987
rect 1647 -3094 1648 -3066
rect 1710 -3067 1711 -2987
rect 366 -3094 367 -3068
rect 394 -3069 395 -2987
rect 450 -3094 451 -3068
rect 492 -3069 493 -2987
rect 499 -3094 500 -3068
rect 1363 -3069 1364 -2987
rect 1710 -3094 1711 -3068
rect 1787 -3069 1788 -2987
rect 317 -3071 318 -2987
rect 394 -3094 395 -3070
rect 492 -3094 493 -3070
rect 646 -3071 647 -2987
rect 653 -3094 654 -3070
rect 891 -3071 892 -2987
rect 1034 -3071 1035 -2987
rect 1374 -3094 1375 -3070
rect 1787 -3094 1788 -3070
rect 1899 -3071 1900 -2987
rect 177 -3073 178 -2987
rect 317 -3094 318 -3072
rect 527 -3073 528 -2987
rect 604 -3094 605 -3072
rect 611 -3073 612 -2987
rect 646 -3094 647 -3072
rect 744 -3073 745 -2987
rect 1010 -3094 1011 -3072
rect 1171 -3094 1172 -3072
rect 1314 -3073 1315 -2987
rect 1899 -3094 1900 -3072
rect 1997 -3073 1998 -2987
rect 23 -3075 24 -2987
rect 611 -3094 612 -3074
rect 772 -3094 773 -3074
rect 821 -3075 822 -2987
rect 863 -3094 864 -3074
rect 1969 -3075 1970 -2987
rect 23 -3094 24 -3076
rect 982 -3077 983 -2987
rect 1507 -3077 1508 -2987
rect 1969 -3094 1970 -3076
rect 177 -3094 178 -3078
rect 303 -3079 304 -2987
rect 331 -3079 332 -2987
rect 821 -3094 822 -3078
rect 982 -3094 983 -3078
rect 989 -3079 990 -2987
rect 1507 -3094 1508 -3078
rect 1577 -3079 1578 -2987
rect 1913 -3079 1914 -2987
rect 1997 -3094 1998 -3078
rect 233 -3081 234 -2987
rect 303 -3094 304 -3080
rect 331 -3094 332 -3080
rect 345 -3081 346 -2987
rect 583 -3081 584 -2987
rect 744 -3094 745 -3080
rect 807 -3081 808 -2987
rect 842 -3094 843 -3080
rect 877 -3094 878 -3080
rect 1577 -3094 1578 -3080
rect 1913 -3094 1914 -3080
rect 2046 -3081 2047 -2987
rect 345 -3094 346 -3082
rect 408 -3083 409 -2987
rect 583 -3094 584 -3082
rect 751 -3083 752 -2987
rect 793 -3083 794 -2987
rect 807 -3094 808 -3082
rect 989 -3094 990 -3082
rect 1458 -3083 1459 -2987
rect 2046 -3094 2047 -3082
rect 2123 -3083 2124 -2987
rect 117 -3085 118 -2987
rect 408 -3094 409 -3084
rect 751 -3094 752 -3084
rect 912 -3094 913 -3084
rect 1458 -3094 1459 -3084
rect 1668 -3085 1669 -2987
rect 793 -3094 794 -3086
rect 1209 -3087 1210 -2987
rect 1668 -3094 1669 -3086
rect 1752 -3087 1753 -2987
rect 1752 -3094 1753 -3088
rect 1829 -3089 1830 -2987
rect 1829 -3094 1830 -3090
rect 1962 -3091 1963 -2987
rect 1962 -3094 1963 -3092
rect 2144 -3093 2145 -2987
rect 23 -3104 24 -3102
rect 208 -3104 209 -3102
rect 212 -3104 213 -3102
rect 233 -3225 234 -3103
rect 303 -3104 304 -3102
rect 303 -3225 304 -3103
rect 303 -3104 304 -3102
rect 303 -3225 304 -3103
rect 380 -3104 381 -3102
rect 457 -3104 458 -3102
rect 520 -3104 521 -3102
rect 817 -3104 818 -3102
rect 821 -3104 822 -3102
rect 1311 -3104 1312 -3102
rect 1381 -3104 1382 -3102
rect 1402 -3104 1403 -3102
rect 1461 -3225 1462 -3103
rect 1864 -3104 1865 -3102
rect 1962 -3104 1963 -3102
rect 2046 -3104 2047 -3102
rect 30 -3106 31 -3102
rect 205 -3106 206 -3102
rect 212 -3225 213 -3105
rect 1167 -3225 1168 -3105
rect 1199 -3106 1200 -3102
rect 1258 -3225 1259 -3105
rect 1276 -3106 1277 -3102
rect 1451 -3106 1452 -3102
rect 1465 -3106 1466 -3102
rect 1563 -3106 1564 -3102
rect 1566 -3106 1567 -3102
rect 1682 -3225 1683 -3105
rect 1853 -3225 1854 -3105
rect 1892 -3106 1893 -3102
rect 1997 -3106 1998 -3102
rect 2018 -3225 2019 -3105
rect 2046 -3225 2047 -3105
rect 2074 -3106 2075 -3102
rect 58 -3108 59 -3102
rect 131 -3108 132 -3102
rect 187 -3225 188 -3107
rect 688 -3108 689 -3102
rect 737 -3108 738 -3102
rect 1444 -3108 1445 -3102
rect 1451 -3225 1452 -3107
rect 1535 -3108 1536 -3102
rect 1640 -3108 1641 -3102
rect 1878 -3108 1879 -3102
rect 1892 -3225 1893 -3107
rect 1948 -3108 1949 -3102
rect 65 -3110 66 -3102
rect 1111 -3225 1112 -3109
rect 1129 -3110 1130 -3102
rect 1129 -3225 1130 -3109
rect 1129 -3110 1130 -3102
rect 1129 -3225 1130 -3109
rect 1199 -3225 1200 -3109
rect 1304 -3110 1305 -3102
rect 1311 -3225 1312 -3109
rect 1703 -3110 1704 -3102
rect 1864 -3225 1865 -3109
rect 1871 -3110 1872 -3102
rect 1878 -3225 1879 -3109
rect 1899 -3110 1900 -3102
rect 72 -3112 73 -3102
rect 236 -3112 237 -3102
rect 289 -3112 290 -3102
rect 821 -3225 822 -3111
rect 835 -3112 836 -3102
rect 1122 -3112 1123 -3102
rect 1216 -3112 1217 -3102
rect 1605 -3112 1606 -3102
rect 1671 -3225 1672 -3111
rect 1857 -3112 1858 -3102
rect 79 -3114 80 -3102
rect 674 -3114 675 -3102
rect 681 -3114 682 -3102
rect 1160 -3114 1161 -3102
rect 1234 -3114 1235 -3102
rect 1346 -3114 1347 -3102
rect 1381 -3225 1382 -3113
rect 1633 -3114 1634 -3102
rect 1675 -3114 1676 -3102
rect 1962 -3225 1963 -3113
rect 86 -3116 87 -3102
rect 138 -3116 139 -3102
rect 194 -3225 195 -3115
rect 282 -3116 283 -3102
rect 289 -3225 290 -3115
rect 425 -3225 426 -3115
rect 436 -3116 437 -3102
rect 436 -3225 437 -3115
rect 436 -3116 437 -3102
rect 436 -3225 437 -3115
rect 506 -3116 507 -3102
rect 737 -3225 738 -3115
rect 758 -3116 759 -3102
rect 1643 -3225 1644 -3115
rect 1857 -3225 1858 -3115
rect 1885 -3116 1886 -3102
rect 93 -3225 94 -3117
rect 142 -3118 143 -3102
rect 198 -3118 199 -3102
rect 198 -3225 199 -3117
rect 198 -3118 199 -3102
rect 198 -3225 199 -3117
rect 254 -3118 255 -3102
rect 282 -3225 283 -3117
rect 352 -3118 353 -3102
rect 1346 -3225 1347 -3117
rect 1388 -3118 1389 -3102
rect 1388 -3225 1389 -3117
rect 1388 -3118 1389 -3102
rect 1388 -3225 1389 -3117
rect 1395 -3118 1396 -3102
rect 1472 -3118 1473 -3102
rect 1486 -3118 1487 -3102
rect 1556 -3118 1557 -3102
rect 1605 -3225 1606 -3117
rect 1850 -3118 1851 -3102
rect 1885 -3225 1886 -3117
rect 1920 -3118 1921 -3102
rect 107 -3120 108 -3102
rect 880 -3120 881 -3102
rect 891 -3120 892 -3102
rect 1115 -3120 1116 -3102
rect 1122 -3225 1123 -3119
rect 1325 -3120 1326 -3102
rect 1395 -3225 1396 -3119
rect 1710 -3120 1711 -3102
rect 1920 -3225 1921 -3119
rect 1976 -3120 1977 -3102
rect 107 -3225 108 -3121
rect 177 -3122 178 -3102
rect 226 -3122 227 -3102
rect 352 -3225 353 -3121
rect 380 -3225 381 -3121
rect 579 -3225 580 -3121
rect 604 -3122 605 -3102
rect 877 -3122 878 -3102
rect 898 -3122 899 -3102
rect 1115 -3225 1116 -3121
rect 1237 -3122 1238 -3102
rect 1409 -3122 1410 -3102
rect 1437 -3122 1438 -3102
rect 1563 -3225 1564 -3121
rect 1633 -3225 1634 -3121
rect 1787 -3122 1788 -3102
rect 1976 -3225 1977 -3121
rect 2004 -3122 2005 -3102
rect 114 -3124 115 -3102
rect 166 -3124 167 -3102
rect 177 -3225 178 -3123
rect 807 -3124 808 -3102
rect 828 -3124 829 -3102
rect 891 -3225 892 -3123
rect 926 -3124 927 -3102
rect 926 -3225 927 -3123
rect 926 -3124 927 -3102
rect 926 -3225 927 -3123
rect 943 -3225 944 -3123
rect 1724 -3124 1725 -3102
rect 100 -3126 101 -3102
rect 114 -3225 115 -3125
rect 121 -3126 122 -3102
rect 208 -3225 209 -3125
rect 254 -3225 255 -3125
rect 359 -3126 360 -3102
rect 401 -3126 402 -3102
rect 530 -3126 531 -3102
rect 555 -3126 556 -3102
rect 873 -3225 874 -3125
rect 877 -3225 878 -3125
rect 1447 -3126 1448 -3102
rect 1465 -3225 1466 -3125
rect 1612 -3126 1613 -3102
rect 1647 -3126 1648 -3102
rect 1724 -3225 1725 -3125
rect 100 -3225 101 -3127
rect 310 -3128 311 -3102
rect 359 -3225 360 -3127
rect 366 -3128 367 -3102
rect 373 -3128 374 -3102
rect 555 -3225 556 -3127
rect 569 -3128 570 -3102
rect 817 -3225 818 -3127
rect 828 -3225 829 -3127
rect 1206 -3128 1207 -3102
rect 1248 -3128 1249 -3102
rect 1269 -3128 1270 -3102
rect 1276 -3225 1277 -3127
rect 1881 -3128 1882 -3102
rect 121 -3225 122 -3129
rect 156 -3130 157 -3102
rect 191 -3130 192 -3102
rect 226 -3225 227 -3129
rect 275 -3130 276 -3102
rect 401 -3225 402 -3129
rect 404 -3225 405 -3129
rect 457 -3225 458 -3129
rect 471 -3130 472 -3102
rect 604 -3225 605 -3129
rect 625 -3130 626 -3102
rect 1083 -3130 1084 -3102
rect 1094 -3130 1095 -3102
rect 1125 -3130 1126 -3102
rect 1185 -3130 1186 -3102
rect 1269 -3225 1270 -3129
rect 1297 -3130 1298 -3102
rect 1314 -3130 1315 -3102
rect 1318 -3130 1319 -3102
rect 1640 -3225 1641 -3129
rect 1647 -3225 1648 -3129
rect 1955 -3130 1956 -3102
rect 135 -3132 136 -3102
rect 275 -3225 276 -3131
rect 296 -3132 297 -3102
rect 373 -3225 374 -3131
rect 471 -3225 472 -3131
rect 534 -3132 535 -3102
rect 541 -3132 542 -3102
rect 569 -3225 570 -3131
rect 625 -3225 626 -3131
rect 709 -3132 710 -3102
rect 716 -3132 717 -3102
rect 835 -3225 836 -3131
rect 863 -3225 864 -3131
rect 919 -3132 920 -3102
rect 961 -3132 962 -3102
rect 1703 -3225 1704 -3131
rect 135 -3225 136 -3133
rect 268 -3134 269 -3102
rect 310 -3225 311 -3133
rect 317 -3134 318 -3102
rect 366 -3225 367 -3133
rect 429 -3134 430 -3102
rect 443 -3134 444 -3102
rect 709 -3225 710 -3133
rect 758 -3225 759 -3133
rect 954 -3134 955 -3102
rect 961 -3225 962 -3133
rect 1031 -3134 1032 -3102
rect 1045 -3134 1046 -3102
rect 1710 -3225 1711 -3133
rect 142 -3225 143 -3135
rect 912 -3136 913 -3102
rect 968 -3136 969 -3102
rect 1559 -3136 1560 -3102
rect 1612 -3225 1613 -3135
rect 1822 -3136 1823 -3102
rect 156 -3225 157 -3137
rect 191 -3225 192 -3137
rect 219 -3138 220 -3102
rect 296 -3225 297 -3137
rect 317 -3225 318 -3137
rect 331 -3138 332 -3102
rect 429 -3225 430 -3137
rect 597 -3138 598 -3102
rect 632 -3138 633 -3102
rect 807 -3225 808 -3137
rect 856 -3138 857 -3102
rect 919 -3225 920 -3137
rect 968 -3225 969 -3137
rect 1227 -3138 1228 -3102
rect 1248 -3225 1249 -3137
rect 1367 -3138 1368 -3102
rect 1402 -3225 1403 -3137
rect 1549 -3138 1550 -3102
rect 1556 -3225 1557 -3137
rect 1906 -3138 1907 -3102
rect 173 -3140 174 -3102
rect 1045 -3225 1046 -3139
rect 1073 -3140 1074 -3102
rect 1304 -3225 1305 -3139
rect 1318 -3225 1319 -3139
rect 1717 -3140 1718 -3102
rect 1766 -3140 1767 -3102
rect 1822 -3225 1823 -3139
rect 1906 -3225 1907 -3139
rect 1934 -3140 1935 -3102
rect 205 -3225 206 -3141
rect 632 -3225 633 -3141
rect 639 -3142 640 -3102
rect 866 -3142 867 -3102
rect 912 -3225 913 -3141
rect 1374 -3142 1375 -3102
rect 1409 -3225 1410 -3141
rect 1542 -3142 1543 -3102
rect 1549 -3225 1550 -3141
rect 1626 -3142 1627 -3102
rect 1661 -3142 1662 -3102
rect 1766 -3225 1767 -3141
rect 219 -3225 220 -3143
rect 261 -3144 262 -3102
rect 268 -3225 269 -3143
rect 345 -3144 346 -3102
rect 394 -3144 395 -3102
rect 639 -3225 640 -3143
rect 681 -3225 682 -3143
rect 702 -3144 703 -3102
rect 765 -3144 766 -3102
rect 1031 -3225 1032 -3143
rect 1073 -3225 1074 -3143
rect 1171 -3144 1172 -3102
rect 1185 -3225 1186 -3143
rect 1360 -3144 1361 -3102
rect 1367 -3225 1368 -3143
rect 1577 -3144 1578 -3102
rect 1626 -3225 1627 -3143
rect 1927 -3144 1928 -3102
rect 261 -3225 262 -3145
rect 1157 -3146 1158 -3102
rect 1171 -3225 1172 -3145
rect 1458 -3146 1459 -3102
rect 1472 -3225 1473 -3145
rect 1668 -3146 1669 -3102
rect 1675 -3225 1676 -3145
rect 1850 -3225 1851 -3145
rect 331 -3225 332 -3147
rect 583 -3148 584 -3102
rect 597 -3225 598 -3147
rect 618 -3148 619 -3102
rect 688 -3225 689 -3147
rect 793 -3148 794 -3102
rect 800 -3148 801 -3102
rect 856 -3225 857 -3147
rect 1017 -3148 1018 -3102
rect 1052 -3225 1053 -3147
rect 1076 -3148 1077 -3102
rect 1657 -3225 1658 -3147
rect 1661 -3225 1662 -3147
rect 1843 -3148 1844 -3102
rect 338 -3150 339 -3102
rect 345 -3225 346 -3149
rect 394 -3225 395 -3149
rect 660 -3150 661 -3102
rect 702 -3225 703 -3149
rect 1024 -3150 1025 -3102
rect 1094 -3225 1095 -3149
rect 1220 -3150 1221 -3102
rect 1227 -3225 1228 -3149
rect 1332 -3150 1333 -3102
rect 1360 -3225 1361 -3149
rect 1507 -3150 1508 -3102
rect 1535 -3225 1536 -3149
rect 1591 -3150 1592 -3102
rect 338 -3225 339 -3151
rect 450 -3152 451 -3102
rect 485 -3152 486 -3102
rect 541 -3225 542 -3151
rect 576 -3152 577 -3102
rect 716 -3225 717 -3151
rect 768 -3225 769 -3151
rect 1192 -3152 1193 -3102
rect 1206 -3225 1207 -3151
rect 1216 -3225 1217 -3151
rect 1220 -3225 1221 -3151
rect 1241 -3152 1242 -3102
rect 1262 -3152 1263 -3102
rect 1444 -3225 1445 -3151
rect 1486 -3225 1487 -3151
rect 1654 -3152 1655 -3102
rect 37 -3154 38 -3102
rect 576 -3225 577 -3153
rect 583 -3225 584 -3153
rect 1055 -3154 1056 -3102
rect 1101 -3154 1102 -3102
rect 1213 -3154 1214 -3102
rect 1241 -3225 1242 -3153
rect 1416 -3154 1417 -3102
rect 1437 -3225 1438 -3153
rect 1685 -3154 1686 -3102
rect 418 -3225 419 -3155
rect 450 -3225 451 -3155
rect 485 -3225 486 -3155
rect 723 -3156 724 -3102
rect 793 -3225 794 -3155
rect 842 -3156 843 -3102
rect 985 -3225 986 -3155
rect 1507 -3225 1508 -3155
rect 1542 -3225 1543 -3155
rect 1815 -3156 1816 -3102
rect 443 -3225 444 -3157
rect 1213 -3225 1214 -3157
rect 1262 -3225 1263 -3157
rect 1493 -3158 1494 -3102
rect 1570 -3158 1571 -3102
rect 1717 -3225 1718 -3157
rect 1738 -3158 1739 -3102
rect 1815 -3225 1816 -3157
rect 506 -3225 507 -3159
rect 933 -3160 934 -3102
rect 989 -3160 990 -3102
rect 1192 -3225 1193 -3159
rect 1297 -3225 1298 -3159
rect 1965 -3160 1966 -3102
rect 520 -3225 521 -3161
rect 1398 -3162 1399 -3102
rect 1416 -3225 1417 -3161
rect 1584 -3162 1585 -3102
rect 1591 -3225 1592 -3161
rect 1801 -3162 1802 -3102
rect 1965 -3225 1966 -3161
rect 2032 -3162 2033 -3102
rect 527 -3164 528 -3102
rect 884 -3164 885 -3102
rect 905 -3164 906 -3102
rect 989 -3225 990 -3163
rect 1003 -3164 1004 -3102
rect 1017 -3225 1018 -3163
rect 1024 -3225 1025 -3163
rect 1059 -3164 1060 -3102
rect 1101 -3225 1102 -3163
rect 1136 -3164 1137 -3102
rect 1157 -3225 1158 -3163
rect 1290 -3164 1291 -3102
rect 1325 -3225 1326 -3163
rect 1514 -3164 1515 -3102
rect 1521 -3164 1522 -3102
rect 1738 -3225 1739 -3163
rect 324 -3166 325 -3102
rect 1290 -3225 1291 -3165
rect 1332 -3225 1333 -3165
rect 1479 -3166 1480 -3102
rect 1493 -3225 1494 -3165
rect 1689 -3166 1690 -3102
rect 324 -3225 325 -3167
rect 387 -3168 388 -3102
rect 527 -3225 528 -3167
rect 744 -3168 745 -3102
rect 786 -3168 787 -3102
rect 884 -3225 885 -3167
rect 905 -3225 906 -3167
rect 975 -3168 976 -3102
rect 1003 -3225 1004 -3167
rect 1066 -3168 1067 -3102
rect 1143 -3168 1144 -3102
rect 1479 -3225 1480 -3167
rect 1500 -3168 1501 -3102
rect 1570 -3225 1571 -3167
rect 1577 -3225 1578 -3167
rect 1941 -3168 1942 -3102
rect 387 -3225 388 -3169
rect 513 -3170 514 -3102
rect 534 -3225 535 -3169
rect 772 -3170 773 -3102
rect 800 -3225 801 -3169
rect 1689 -3225 1690 -3169
rect 464 -3172 465 -3102
rect 744 -3225 745 -3171
rect 814 -3172 815 -3102
rect 1374 -3225 1375 -3171
rect 1500 -3225 1501 -3171
rect 1598 -3172 1599 -3102
rect 1650 -3225 1651 -3171
rect 1685 -3225 1686 -3171
rect 163 -3174 164 -3102
rect 464 -3225 465 -3173
rect 492 -3174 493 -3102
rect 975 -3225 976 -3173
rect 1059 -3225 1060 -3173
rect 1150 -3174 1151 -3102
rect 1356 -3225 1357 -3173
rect 1521 -3225 1522 -3173
rect 1584 -3225 1585 -3173
rect 1731 -3174 1732 -3102
rect 163 -3225 164 -3175
rect 765 -3225 766 -3175
rect 933 -3225 934 -3175
rect 982 -3176 983 -3102
rect 1066 -3225 1067 -3175
rect 1108 -3176 1109 -3102
rect 1143 -3225 1144 -3175
rect 1178 -3176 1179 -3102
rect 1514 -3225 1515 -3175
rect 1696 -3176 1697 -3102
rect 1731 -3225 1732 -3175
rect 1745 -3176 1746 -3102
rect 415 -3178 416 -3102
rect 492 -3225 493 -3177
rect 513 -3225 514 -3177
rect 590 -3178 591 -3102
rect 611 -3178 612 -3102
rect 786 -3225 787 -3177
rect 940 -3178 941 -3102
rect 1136 -3225 1137 -3177
rect 1150 -3225 1151 -3177
rect 1283 -3178 1284 -3102
rect 1598 -3225 1599 -3177
rect 1836 -3178 1837 -3102
rect 415 -3225 416 -3179
rect 898 -3225 899 -3179
rect 954 -3225 955 -3179
rect 1178 -3225 1179 -3179
rect 1283 -3225 1284 -3179
rect 1339 -3180 1340 -3102
rect 1654 -3225 1655 -3179
rect 1969 -3180 1970 -3102
rect 184 -3182 185 -3102
rect 1339 -3225 1340 -3181
rect 1696 -3225 1697 -3181
rect 1808 -3182 1809 -3102
rect 1969 -3225 1970 -3181
rect 1983 -3182 1984 -3102
rect 590 -3225 591 -3183
rect 695 -3184 696 -3102
rect 730 -3184 731 -3102
rect 814 -3225 815 -3183
rect 1108 -3225 1109 -3183
rect 1353 -3184 1354 -3102
rect 1745 -3225 1746 -3183
rect 1759 -3184 1760 -3102
rect 1780 -3184 1781 -3102
rect 1808 -3225 1809 -3183
rect 1983 -3225 1984 -3183
rect 1990 -3184 1991 -3102
rect 82 -3186 83 -3102
rect 730 -3225 731 -3185
rect 772 -3225 773 -3185
rect 1353 -3225 1354 -3185
rect 1752 -3186 1753 -3102
rect 1759 -3225 1760 -3185
rect 1773 -3186 1774 -3102
rect 1780 -3225 1781 -3185
rect 562 -3188 563 -3102
rect 695 -3225 696 -3187
rect 1752 -3225 1753 -3187
rect 1794 -3188 1795 -3102
rect 499 -3190 500 -3102
rect 562 -3225 563 -3189
rect 611 -3225 612 -3189
rect 667 -3190 668 -3102
rect 674 -3225 675 -3189
rect 723 -3225 724 -3189
rect 1773 -3225 1774 -3189
rect 1829 -3190 1830 -3102
rect 499 -3225 500 -3191
rect 779 -3192 780 -3102
rect 614 -3194 615 -3102
rect 940 -3225 941 -3193
rect 247 -3196 248 -3102
rect 614 -3225 615 -3195
rect 618 -3225 619 -3195
rect 646 -3196 647 -3102
rect 653 -3196 654 -3102
rect 842 -3225 843 -3195
rect 240 -3198 241 -3102
rect 247 -3225 248 -3197
rect 478 -3198 479 -3102
rect 653 -3225 654 -3197
rect 660 -3225 661 -3197
rect 1080 -3198 1081 -3102
rect 170 -3200 171 -3102
rect 240 -3225 241 -3199
rect 408 -3200 409 -3102
rect 478 -3225 479 -3199
rect 548 -3200 549 -3102
rect 646 -3225 647 -3199
rect 667 -3225 668 -3199
rect 870 -3200 871 -3102
rect 170 -3225 171 -3201
rect 751 -3202 752 -3102
rect 779 -3225 780 -3201
rect 947 -3202 948 -3102
rect 128 -3204 129 -3102
rect 751 -3225 752 -3203
rect 849 -3204 850 -3102
rect 1080 -3225 1081 -3203
rect 128 -3225 129 -3205
rect 149 -3206 150 -3102
rect 408 -3225 409 -3205
rect 422 -3206 423 -3102
rect 548 -3225 549 -3205
rect 747 -3225 748 -3205
rect 849 -3225 850 -3205
rect 1038 -3206 1039 -3102
rect 149 -3225 150 -3207
rect 460 -3208 461 -3102
rect 947 -3225 948 -3207
rect 996 -3208 997 -3102
rect 1038 -3225 1039 -3207
rect 1087 -3208 1088 -3102
rect 996 -3225 997 -3209
rect 1010 -3210 1011 -3102
rect 1087 -3225 1088 -3209
rect 1255 -3210 1256 -3102
rect 1010 -3225 1011 -3211
rect 1458 -3225 1459 -3211
rect 1255 -3225 1256 -3213
rect 1423 -3214 1424 -3102
rect 1164 -3216 1165 -3102
rect 1423 -3225 1424 -3215
rect 1164 -3225 1165 -3217
rect 1528 -3218 1529 -3102
rect 1430 -3220 1431 -3102
rect 1528 -3225 1529 -3219
rect 1430 -3225 1431 -3221
rect 1619 -3222 1620 -3102
rect 1619 -3225 1620 -3223
rect 1913 -3224 1914 -3102
rect 93 -3235 94 -3233
rect 173 -3235 174 -3233
rect 184 -3328 185 -3234
rect 537 -3328 538 -3234
rect 541 -3235 542 -3233
rect 541 -3328 542 -3234
rect 541 -3235 542 -3233
rect 541 -3328 542 -3234
rect 548 -3235 549 -3233
rect 600 -3328 601 -3234
rect 642 -3328 643 -3234
rect 772 -3235 773 -3233
rect 800 -3235 801 -3233
rect 1444 -3235 1445 -3233
rect 1563 -3235 1564 -3233
rect 1643 -3235 1644 -3233
rect 1668 -3328 1669 -3234
rect 1727 -3328 1728 -3234
rect 1738 -3235 1739 -3233
rect 1965 -3235 1966 -3233
rect 1969 -3235 1970 -3233
rect 1969 -3328 1970 -3234
rect 1969 -3235 1970 -3233
rect 1969 -3328 1970 -3234
rect 2018 -3235 2019 -3233
rect 2025 -3328 2026 -3234
rect 2032 -3328 2033 -3234
rect 2046 -3235 2047 -3233
rect 107 -3237 108 -3233
rect 677 -3237 678 -3233
rect 688 -3237 689 -3233
rect 1164 -3237 1165 -3233
rect 1213 -3237 1214 -3233
rect 1598 -3237 1599 -3233
rect 1640 -3237 1641 -3233
rect 1745 -3237 1746 -3233
rect 1766 -3237 1767 -3233
rect 1787 -3328 1788 -3236
rect 1808 -3237 1809 -3233
rect 1850 -3237 1851 -3233
rect 1857 -3237 1858 -3233
rect 1857 -3328 1858 -3236
rect 1857 -3237 1858 -3233
rect 1857 -3328 1858 -3236
rect 1871 -3328 1872 -3236
rect 1885 -3237 1886 -3233
rect 1962 -3237 1963 -3233
rect 1983 -3237 1984 -3233
rect 121 -3239 122 -3233
rect 205 -3239 206 -3233
rect 208 -3239 209 -3233
rect 226 -3239 227 -3233
rect 233 -3239 234 -3233
rect 257 -3328 258 -3238
rect 275 -3239 276 -3233
rect 782 -3328 783 -3238
rect 800 -3328 801 -3238
rect 898 -3239 899 -3233
rect 929 -3328 930 -3238
rect 1605 -3239 1606 -3233
rect 1689 -3239 1690 -3233
rect 1794 -3328 1795 -3238
rect 1815 -3239 1816 -3233
rect 1843 -3328 1844 -3238
rect 1878 -3239 1879 -3233
rect 1878 -3328 1879 -3238
rect 1878 -3239 1879 -3233
rect 1878 -3328 1879 -3238
rect 1962 -3328 1963 -3238
rect 1976 -3239 1977 -3233
rect 100 -3241 101 -3233
rect 226 -3328 227 -3240
rect 247 -3241 248 -3233
rect 275 -3328 276 -3240
rect 282 -3241 283 -3233
rect 415 -3241 416 -3233
rect 464 -3241 465 -3233
rect 870 -3241 871 -3233
rect 873 -3241 874 -3233
rect 1465 -3241 1466 -3233
rect 1528 -3241 1529 -3233
rect 1605 -3328 1606 -3240
rect 1703 -3241 1704 -3233
rect 1801 -3328 1802 -3240
rect 1815 -3328 1816 -3240
rect 1850 -3328 1851 -3240
rect 128 -3243 129 -3233
rect 187 -3243 188 -3233
rect 191 -3243 192 -3233
rect 1584 -3243 1585 -3233
rect 1598 -3328 1599 -3242
rect 1633 -3243 1634 -3233
rect 1717 -3243 1718 -3233
rect 1738 -3328 1739 -3242
rect 1745 -3328 1746 -3242
rect 1773 -3243 1774 -3233
rect 1780 -3243 1781 -3233
rect 1780 -3328 1781 -3242
rect 1780 -3243 1781 -3233
rect 1780 -3328 1781 -3242
rect 1822 -3243 1823 -3233
rect 1836 -3328 1837 -3242
rect 135 -3245 136 -3233
rect 719 -3245 720 -3233
rect 751 -3245 752 -3233
rect 943 -3245 944 -3233
rect 957 -3245 958 -3233
rect 996 -3245 997 -3233
rect 1104 -3328 1105 -3244
rect 1220 -3245 1221 -3233
rect 1237 -3245 1238 -3233
rect 1619 -3245 1620 -3233
rect 1717 -3328 1718 -3244
rect 1731 -3245 1732 -3233
rect 1759 -3245 1760 -3233
rect 1766 -3328 1767 -3244
rect 156 -3247 157 -3233
rect 170 -3328 171 -3246
rect 191 -3328 192 -3246
rect 1647 -3247 1648 -3233
rect 1731 -3328 1732 -3246
rect 1752 -3247 1753 -3233
rect 205 -3328 206 -3248
rect 212 -3249 213 -3233
rect 215 -3328 216 -3248
rect 1069 -3328 1070 -3248
rect 1108 -3249 1109 -3233
rect 1682 -3249 1683 -3233
rect 1724 -3249 1725 -3233
rect 1752 -3328 1753 -3248
rect 219 -3251 220 -3233
rect 803 -3251 804 -3233
rect 814 -3328 815 -3250
rect 1010 -3251 1011 -3233
rect 1108 -3328 1109 -3250
rect 1129 -3251 1130 -3233
rect 1216 -3251 1217 -3233
rect 1409 -3251 1410 -3233
rect 1465 -3328 1466 -3250
rect 1654 -3251 1655 -3233
rect 219 -3328 220 -3252
rect 415 -3328 416 -3252
rect 464 -3328 465 -3252
rect 506 -3253 507 -3233
rect 513 -3253 514 -3233
rect 614 -3253 615 -3233
rect 632 -3253 633 -3233
rect 1129 -3328 1130 -3252
rect 1216 -3328 1217 -3252
rect 1346 -3253 1347 -3233
rect 1353 -3253 1354 -3233
rect 1591 -3253 1592 -3233
rect 1654 -3328 1655 -3252
rect 1696 -3253 1697 -3233
rect 240 -3255 241 -3233
rect 506 -3328 507 -3254
rect 569 -3255 570 -3233
rect 569 -3328 570 -3254
rect 569 -3255 570 -3233
rect 569 -3328 570 -3254
rect 576 -3255 577 -3233
rect 1650 -3255 1651 -3233
rect 240 -3328 241 -3256
rect 639 -3257 640 -3233
rect 653 -3257 654 -3233
rect 688 -3328 689 -3256
rect 716 -3257 717 -3233
rect 1332 -3257 1333 -3233
rect 1346 -3328 1347 -3256
rect 1486 -3257 1487 -3233
rect 1549 -3257 1550 -3233
rect 1591 -3328 1592 -3256
rect 247 -3328 248 -3258
rect 261 -3259 262 -3233
rect 282 -3328 283 -3258
rect 660 -3259 661 -3233
rect 674 -3328 675 -3258
rect 702 -3259 703 -3233
rect 716 -3328 717 -3258
rect 992 -3328 993 -3258
rect 1080 -3259 1081 -3233
rect 1353 -3328 1354 -3258
rect 1374 -3259 1375 -3233
rect 1444 -3328 1445 -3258
rect 1472 -3259 1473 -3233
rect 1528 -3328 1529 -3258
rect 1563 -3328 1564 -3258
rect 1661 -3259 1662 -3233
rect 254 -3261 255 -3233
rect 261 -3328 262 -3260
rect 303 -3261 304 -3233
rect 303 -3328 304 -3260
rect 303 -3261 304 -3233
rect 303 -3328 304 -3260
rect 331 -3261 332 -3233
rect 744 -3328 745 -3260
rect 751 -3328 752 -3260
rect 807 -3261 808 -3233
rect 856 -3261 857 -3233
rect 982 -3328 983 -3260
rect 985 -3261 986 -3233
rect 1269 -3261 1270 -3233
rect 1290 -3261 1291 -3233
rect 1458 -3261 1459 -3233
rect 1486 -3328 1487 -3260
rect 1580 -3261 1581 -3233
rect 1661 -3328 1662 -3260
rect 1675 -3261 1676 -3233
rect 268 -3263 269 -3233
rect 331 -3328 332 -3262
rect 338 -3263 339 -3233
rect 726 -3328 727 -3262
rect 772 -3328 773 -3262
rect 793 -3263 794 -3233
rect 807 -3328 808 -3262
rect 947 -3263 948 -3233
rect 957 -3328 958 -3262
rect 1164 -3328 1165 -3262
rect 1167 -3263 1168 -3233
rect 1472 -3328 1473 -3262
rect 268 -3328 269 -3264
rect 289 -3265 290 -3233
rect 338 -3328 339 -3264
rect 604 -3265 605 -3233
rect 653 -3328 654 -3264
rect 695 -3265 696 -3233
rect 702 -3328 703 -3264
rect 1255 -3265 1256 -3233
rect 1269 -3328 1270 -3264
rect 1612 -3265 1613 -3233
rect 289 -3328 290 -3266
rect 345 -3267 346 -3233
rect 352 -3267 353 -3233
rect 418 -3267 419 -3233
rect 485 -3267 486 -3233
rect 513 -3328 514 -3266
rect 562 -3267 563 -3233
rect 856 -3328 857 -3266
rect 863 -3267 864 -3233
rect 870 -3328 871 -3266
rect 898 -3328 899 -3266
rect 1094 -3267 1095 -3233
rect 1115 -3267 1116 -3233
rect 1234 -3267 1235 -3233
rect 1237 -3328 1238 -3266
rect 1685 -3267 1686 -3233
rect 345 -3328 346 -3268
rect 646 -3269 647 -3233
rect 660 -3328 661 -3268
rect 667 -3269 668 -3233
rect 695 -3328 696 -3268
rect 730 -3269 731 -3233
rect 793 -3328 794 -3268
rect 1031 -3269 1032 -3233
rect 1115 -3328 1116 -3268
rect 1192 -3269 1193 -3233
rect 1220 -3328 1221 -3268
rect 1493 -3269 1494 -3233
rect 352 -3328 353 -3270
rect 443 -3271 444 -3233
rect 485 -3328 486 -3270
rect 786 -3271 787 -3233
rect 912 -3271 913 -3233
rect 1010 -3328 1011 -3270
rect 1031 -3328 1032 -3270
rect 1150 -3271 1151 -3233
rect 1171 -3271 1172 -3233
rect 1255 -3328 1256 -3270
rect 1290 -3328 1291 -3270
rect 1311 -3271 1312 -3233
rect 1332 -3328 1333 -3270
rect 1339 -3271 1340 -3233
rect 1374 -3328 1375 -3270
rect 1514 -3271 1515 -3233
rect 229 -3328 230 -3272
rect 443 -3328 444 -3272
rect 495 -3273 496 -3233
rect 579 -3273 580 -3233
rect 583 -3273 584 -3233
rect 639 -3328 640 -3272
rect 646 -3328 647 -3272
rect 681 -3273 682 -3233
rect 786 -3328 787 -3272
rect 1059 -3273 1060 -3233
rect 1066 -3273 1067 -3233
rect 1493 -3328 1494 -3272
rect 1500 -3273 1501 -3233
rect 1514 -3328 1515 -3272
rect 359 -3275 360 -3233
rect 422 -3275 423 -3233
rect 499 -3275 500 -3233
rect 733 -3328 734 -3274
rect 912 -3328 913 -3274
rect 933 -3275 934 -3233
rect 947 -3328 948 -3274
rect 1003 -3275 1004 -3233
rect 1059 -3328 1060 -3274
rect 1178 -3275 1179 -3233
rect 1192 -3328 1193 -3274
rect 1262 -3275 1263 -3233
rect 1283 -3275 1284 -3233
rect 1500 -3328 1501 -3274
rect 177 -3277 178 -3233
rect 499 -3328 500 -3276
rect 527 -3277 528 -3233
rect 681 -3328 682 -3276
rect 709 -3277 710 -3233
rect 1003 -3328 1004 -3276
rect 1066 -3328 1067 -3276
rect 1227 -3277 1228 -3233
rect 1262 -3328 1263 -3276
rect 1556 -3277 1557 -3233
rect 177 -3328 178 -3278
rect 198 -3279 199 -3233
rect 359 -3328 360 -3278
rect 436 -3279 437 -3233
rect 527 -3328 528 -3278
rect 817 -3279 818 -3233
rect 919 -3279 920 -3233
rect 933 -3328 934 -3278
rect 968 -3279 969 -3233
rect 996 -3328 997 -3278
rect 1150 -3328 1151 -3278
rect 1297 -3279 1298 -3233
rect 1311 -3328 1312 -3278
rect 1318 -3279 1319 -3233
rect 1409 -3328 1410 -3278
rect 1853 -3279 1854 -3233
rect 163 -3281 164 -3233
rect 198 -3328 199 -3280
rect 366 -3281 367 -3233
rect 422 -3328 423 -3280
rect 555 -3281 556 -3233
rect 1339 -3328 1340 -3280
rect 1458 -3328 1459 -3280
rect 1542 -3281 1543 -3233
rect 1853 -3328 1854 -3280
rect 1864 -3281 1865 -3233
rect 142 -3283 143 -3233
rect 163 -3328 164 -3282
rect 324 -3283 325 -3233
rect 366 -3328 367 -3282
rect 373 -3283 374 -3233
rect 436 -3328 437 -3282
rect 478 -3283 479 -3233
rect 555 -3328 556 -3282
rect 562 -3328 563 -3282
rect 597 -3283 598 -3233
rect 604 -3328 605 -3282
rect 737 -3283 738 -3233
rect 919 -3328 920 -3282
rect 954 -3283 955 -3233
rect 968 -3328 969 -3282
rect 1122 -3283 1123 -3233
rect 1157 -3283 1158 -3233
rect 1227 -3328 1228 -3282
rect 1283 -3328 1284 -3282
rect 1381 -3283 1382 -3233
rect 1535 -3283 1536 -3233
rect 1556 -3328 1557 -3282
rect 1864 -3328 1865 -3282
rect 1892 -3283 1893 -3233
rect 117 -3285 118 -3233
rect 142 -3328 143 -3284
rect 310 -3285 311 -3233
rect 597 -3328 598 -3284
rect 667 -3328 668 -3284
rect 779 -3285 780 -3233
rect 1122 -3328 1123 -3284
rect 1206 -3285 1207 -3233
rect 1297 -3328 1298 -3284
rect 1367 -3285 1368 -3233
rect 1892 -3328 1893 -3284
rect 1906 -3285 1907 -3233
rect 310 -3328 311 -3286
rect 317 -3287 318 -3233
rect 324 -3328 325 -3286
rect 429 -3287 430 -3233
rect 576 -3328 577 -3286
rect 940 -3287 941 -3233
rect 1143 -3287 1144 -3233
rect 1157 -3328 1158 -3286
rect 1171 -3328 1172 -3286
rect 1388 -3287 1389 -3233
rect 1906 -3328 1907 -3286
rect 1920 -3287 1921 -3233
rect 317 -3328 318 -3288
rect 625 -3289 626 -3233
rect 709 -3328 710 -3288
rect 835 -3289 836 -3233
rect 940 -3328 941 -3288
rect 1024 -3289 1025 -3233
rect 1178 -3328 1179 -3288
rect 1416 -3289 1417 -3233
rect 373 -3328 374 -3290
rect 450 -3291 451 -3233
rect 583 -3328 584 -3290
rect 611 -3291 612 -3233
rect 625 -3328 626 -3290
rect 1094 -3328 1095 -3290
rect 1206 -3328 1207 -3290
rect 1437 -3291 1438 -3233
rect 149 -3293 150 -3233
rect 611 -3328 612 -3292
rect 737 -3328 738 -3292
rect 1017 -3293 1018 -3233
rect 1024 -3328 1025 -3292
rect 1052 -3293 1053 -3233
rect 1318 -3328 1319 -3292
rect 1430 -3293 1431 -3233
rect 383 -3328 384 -3294
rect 863 -3328 864 -3294
rect 961 -3295 962 -3233
rect 1388 -3328 1389 -3294
rect 1402 -3295 1403 -3233
rect 1437 -3328 1438 -3294
rect 387 -3297 388 -3233
rect 492 -3328 493 -3296
rect 590 -3297 591 -3233
rect 632 -3328 633 -3296
rect 765 -3297 766 -3233
rect 1017 -3328 1018 -3296
rect 1038 -3297 1039 -3233
rect 1052 -3328 1053 -3296
rect 1136 -3297 1137 -3233
rect 1402 -3328 1403 -3296
rect 387 -3328 388 -3298
rect 471 -3299 472 -3233
rect 590 -3328 591 -3298
rect 1087 -3299 1088 -3233
rect 1136 -3328 1137 -3298
rect 1199 -3299 1200 -3233
rect 1325 -3299 1326 -3233
rect 1430 -3328 1431 -3298
rect 394 -3301 395 -3233
rect 548 -3328 549 -3300
rect 765 -3328 766 -3300
rect 905 -3301 906 -3233
rect 961 -3328 962 -3300
rect 989 -3301 990 -3233
rect 1038 -3328 1039 -3300
rect 1080 -3328 1081 -3300
rect 1087 -3328 1088 -3300
rect 1185 -3301 1186 -3233
rect 1199 -3328 1200 -3300
rect 1360 -3301 1361 -3233
rect 1367 -3328 1368 -3300
rect 1570 -3301 1571 -3233
rect 394 -3328 395 -3302
rect 408 -3303 409 -3233
rect 429 -3328 430 -3302
rect 534 -3303 535 -3233
rect 723 -3303 724 -3233
rect 1185 -3328 1186 -3302
rect 1325 -3328 1326 -3302
rect 1521 -3303 1522 -3233
rect 380 -3305 381 -3233
rect 408 -3328 409 -3304
rect 450 -3328 451 -3304
rect 618 -3305 619 -3233
rect 779 -3328 780 -3304
rect 1276 -3305 1277 -3233
rect 1451 -3305 1452 -3233
rect 1521 -3328 1522 -3304
rect 380 -3328 381 -3306
rect 478 -3328 479 -3306
rect 534 -3328 535 -3306
rect 1671 -3307 1672 -3233
rect 401 -3309 402 -3233
rect 618 -3328 619 -3308
rect 821 -3309 822 -3233
rect 835 -3328 836 -3308
rect 884 -3309 885 -3233
rect 1360 -3328 1361 -3308
rect 1451 -3328 1452 -3308
rect 1507 -3309 1508 -3233
rect 296 -3311 297 -3233
rect 401 -3328 402 -3310
rect 404 -3311 405 -3233
rect 457 -3311 458 -3233
rect 471 -3328 472 -3310
rect 975 -3311 976 -3233
rect 978 -3328 979 -3310
rect 1143 -3328 1144 -3310
rect 1248 -3311 1249 -3233
rect 1276 -3328 1277 -3310
rect 1423 -3311 1424 -3233
rect 1507 -3328 1508 -3310
rect 296 -3328 297 -3312
rect 768 -3313 769 -3233
rect 821 -3328 822 -3312
rect 842 -3313 843 -3233
rect 849 -3313 850 -3233
rect 884 -3328 885 -3312
rect 905 -3328 906 -3312
rect 1234 -3328 1235 -3312
rect 1248 -3328 1249 -3312
rect 1479 -3313 1480 -3233
rect 457 -3328 458 -3314
rect 520 -3315 521 -3233
rect 842 -3328 843 -3314
rect 877 -3315 878 -3233
rect 989 -3328 990 -3314
rect 1626 -3315 1627 -3233
rect 520 -3328 521 -3316
rect 758 -3317 759 -3233
rect 877 -3328 878 -3316
rect 891 -3317 892 -3233
rect 1304 -3317 1305 -3233
rect 1423 -3328 1424 -3316
rect 1479 -3328 1480 -3316
rect 1724 -3328 1725 -3316
rect 758 -3328 759 -3318
rect 849 -3328 850 -3318
rect 1304 -3328 1305 -3318
rect 1395 -3319 1396 -3233
rect 1626 -3328 1627 -3318
rect 1710 -3319 1711 -3233
rect 828 -3321 829 -3233
rect 891 -3328 892 -3320
rect 1073 -3321 1074 -3233
rect 1395 -3328 1396 -3320
rect 828 -3328 829 -3322
rect 926 -3323 927 -3233
rect 1073 -3328 1074 -3322
rect 1241 -3323 1242 -3233
rect 254 -3328 255 -3324
rect 926 -3328 927 -3324
rect 1045 -3325 1046 -3233
rect 1241 -3328 1242 -3324
rect 1045 -3328 1046 -3326
rect 1101 -3327 1102 -3233
rect 142 -3338 143 -3336
rect 173 -3415 174 -3337
rect 177 -3338 178 -3336
rect 236 -3338 237 -3336
rect 257 -3338 258 -3336
rect 373 -3338 374 -3336
rect 394 -3338 395 -3336
rect 537 -3338 538 -3336
rect 541 -3338 542 -3336
rect 544 -3348 545 -3337
rect 590 -3338 591 -3336
rect 779 -3338 780 -3336
rect 814 -3338 815 -3336
rect 1125 -3415 1126 -3337
rect 1160 -3415 1161 -3337
rect 1227 -3338 1228 -3336
rect 1234 -3338 1235 -3336
rect 1451 -3338 1452 -3336
rect 1500 -3338 1501 -3336
rect 1500 -3415 1501 -3337
rect 1500 -3338 1501 -3336
rect 1500 -3415 1501 -3337
rect 1521 -3338 1522 -3336
rect 1584 -3415 1585 -3337
rect 1591 -3338 1592 -3336
rect 1612 -3415 1613 -3337
rect 1647 -3415 1648 -3337
rect 1661 -3338 1662 -3336
rect 1717 -3338 1718 -3336
rect 1727 -3338 1728 -3336
rect 1731 -3338 1732 -3336
rect 1731 -3415 1732 -3337
rect 1731 -3338 1732 -3336
rect 1731 -3415 1732 -3337
rect 1738 -3338 1739 -3336
rect 1738 -3415 1739 -3337
rect 1738 -3338 1739 -3336
rect 1738 -3415 1739 -3337
rect 1752 -3338 1753 -3336
rect 1759 -3415 1760 -3337
rect 1766 -3338 1767 -3336
rect 1769 -3415 1770 -3337
rect 1780 -3338 1781 -3336
rect 1780 -3415 1781 -3337
rect 1780 -3338 1781 -3336
rect 1780 -3415 1781 -3337
rect 1787 -3338 1788 -3336
rect 1811 -3415 1812 -3337
rect 1829 -3415 1830 -3337
rect 1843 -3338 1844 -3336
rect 1885 -3338 1886 -3336
rect 1906 -3338 1907 -3336
rect 1955 -3415 1956 -3337
rect 1962 -3338 1963 -3336
rect 2025 -3338 2026 -3336
rect 2028 -3338 2029 -3336
rect 163 -3340 164 -3336
rect 390 -3415 391 -3339
rect 415 -3340 416 -3336
rect 485 -3340 486 -3336
rect 488 -3415 489 -3339
rect 506 -3340 507 -3336
rect 513 -3340 514 -3336
rect 992 -3415 993 -3339
rect 1034 -3415 1035 -3339
rect 1220 -3340 1221 -3336
rect 1234 -3415 1235 -3339
rect 1283 -3340 1284 -3336
rect 1339 -3340 1340 -3336
rect 1458 -3340 1459 -3336
rect 1521 -3415 1522 -3339
rect 1528 -3340 1529 -3336
rect 1549 -3415 1550 -3339
rect 1626 -3340 1627 -3336
rect 1724 -3415 1725 -3339
rect 1745 -3340 1746 -3336
rect 1787 -3415 1788 -3339
rect 1850 -3340 1851 -3336
rect 1888 -3340 1889 -3336
rect 1892 -3340 1893 -3336
rect 1962 -3415 1963 -3339
rect 1969 -3340 1970 -3336
rect 2025 -3415 2026 -3339
rect 2032 -3340 2033 -3336
rect 170 -3342 171 -3336
rect 180 -3415 181 -3341
rect 212 -3342 213 -3336
rect 408 -3342 409 -3336
rect 429 -3342 430 -3336
rect 926 -3342 927 -3336
rect 968 -3342 969 -3336
rect 1332 -3342 1333 -3336
rect 1367 -3415 1368 -3341
rect 1493 -3342 1494 -3336
rect 1528 -3415 1529 -3341
rect 1563 -3342 1564 -3336
rect 1605 -3342 1606 -3336
rect 1654 -3342 1655 -3336
rect 1794 -3342 1795 -3336
rect 1822 -3415 1823 -3341
rect 1836 -3342 1837 -3336
rect 1843 -3415 1844 -3341
rect 1850 -3415 1851 -3341
rect 1857 -3342 1858 -3336
rect 215 -3344 216 -3336
rect 803 -3415 804 -3343
rect 821 -3344 822 -3336
rect 936 -3415 937 -3343
rect 968 -3415 969 -3343
rect 1003 -3344 1004 -3336
rect 1031 -3344 1032 -3336
rect 1220 -3415 1221 -3343
rect 1237 -3344 1238 -3336
rect 1297 -3344 1298 -3336
rect 1332 -3415 1333 -3343
rect 1374 -3344 1375 -3336
rect 1381 -3344 1382 -3336
rect 1444 -3344 1445 -3336
rect 1451 -3415 1452 -3343
rect 1486 -3344 1487 -3336
rect 1552 -3415 1553 -3343
rect 1598 -3344 1599 -3336
rect 1608 -3344 1609 -3336
rect 1668 -3344 1669 -3336
rect 1801 -3344 1802 -3336
rect 1836 -3415 1837 -3343
rect 1857 -3415 1858 -3343
rect 1871 -3344 1872 -3336
rect 240 -3346 241 -3336
rect 506 -3415 507 -3345
rect 541 -3415 542 -3345
rect 597 -3346 598 -3336
rect 1083 -3346 1084 -3336
rect 1097 -3346 1098 -3336
rect 1311 -3346 1312 -3336
rect 1374 -3415 1375 -3345
rect 1458 -3415 1459 -3345
rect 1556 -3346 1557 -3336
rect 1587 -3415 1588 -3345
rect 1654 -3415 1655 -3345
rect 1853 -3346 1854 -3336
rect 1864 -3346 1865 -3336
rect 1871 -3415 1872 -3345
rect 275 -3348 276 -3336
rect 373 -3415 374 -3347
rect 422 -3348 423 -3336
rect 429 -3415 430 -3347
rect 474 -3415 475 -3347
rect 1370 -3348 1371 -3336
rect 1384 -3348 1385 -3336
rect 1423 -3348 1424 -3336
rect 1801 -3415 1802 -3347
rect 1815 -3348 1816 -3336
rect 1864 -3415 1865 -3347
rect 1878 -3348 1879 -3336
rect 2028 -3415 2029 -3347
rect 2032 -3415 2033 -3347
rect 205 -3350 206 -3336
rect 422 -3415 423 -3349
rect 548 -3350 549 -3336
rect 1031 -3415 1032 -3349
rect 1066 -3350 1067 -3336
rect 1430 -3350 1431 -3336
rect 282 -3352 283 -3336
rect 859 -3415 860 -3351
rect 877 -3352 878 -3336
rect 1003 -3415 1004 -3351
rect 1080 -3352 1081 -3336
rect 1136 -3352 1137 -3336
rect 1199 -3352 1200 -3336
rect 1227 -3415 1228 -3351
rect 1269 -3352 1270 -3336
rect 1353 -3352 1354 -3336
rect 1388 -3352 1389 -3336
rect 1419 -3352 1420 -3336
rect 296 -3354 297 -3336
rect 383 -3354 384 -3336
rect 492 -3354 493 -3336
rect 548 -3415 549 -3353
rect 555 -3354 556 -3336
rect 590 -3415 591 -3353
rect 597 -3415 598 -3353
rect 646 -3354 647 -3336
rect 653 -3354 654 -3336
rect 877 -3415 878 -3353
rect 891 -3354 892 -3336
rect 954 -3354 955 -3336
rect 961 -3354 962 -3336
rect 1080 -3415 1081 -3353
rect 1101 -3415 1102 -3353
rect 1178 -3354 1179 -3336
rect 1199 -3415 1200 -3353
rect 1325 -3354 1326 -3336
rect 1416 -3354 1417 -3336
rect 1437 -3354 1438 -3336
rect 268 -3356 269 -3336
rect 296 -3415 297 -3355
rect 317 -3356 318 -3336
rect 408 -3415 409 -3355
rect 450 -3356 451 -3336
rect 492 -3415 493 -3355
rect 534 -3356 535 -3336
rect 646 -3415 647 -3355
rect 674 -3356 675 -3336
rect 1027 -3415 1028 -3355
rect 1045 -3356 1046 -3336
rect 1178 -3415 1179 -3355
rect 1213 -3356 1214 -3336
rect 1402 -3356 1403 -3336
rect 359 -3358 360 -3336
rect 513 -3415 514 -3357
rect 534 -3415 535 -3357
rect 583 -3358 584 -3336
rect 618 -3358 619 -3336
rect 639 -3415 640 -3357
rect 660 -3358 661 -3336
rect 674 -3415 675 -3357
rect 681 -3358 682 -3336
rect 1066 -3415 1067 -3357
rect 1157 -3358 1158 -3336
rect 1213 -3415 1214 -3357
rect 1269 -3415 1270 -3357
rect 1472 -3358 1473 -3336
rect 303 -3360 304 -3336
rect 359 -3415 360 -3359
rect 366 -3360 367 -3336
rect 394 -3415 395 -3359
rect 478 -3360 479 -3336
rect 555 -3415 556 -3359
rect 562 -3360 563 -3336
rect 681 -3415 682 -3359
rect 716 -3360 717 -3336
rect 716 -3415 717 -3359
rect 716 -3360 717 -3336
rect 716 -3415 717 -3359
rect 723 -3360 724 -3336
rect 1395 -3360 1396 -3336
rect 1472 -3415 1473 -3359
rect 1514 -3360 1515 -3336
rect 331 -3362 332 -3336
rect 478 -3415 479 -3361
rect 562 -3415 563 -3361
rect 726 -3415 727 -3361
rect 730 -3362 731 -3336
rect 1808 -3415 1809 -3361
rect 198 -3364 199 -3336
rect 331 -3415 332 -3363
rect 345 -3364 346 -3336
rect 660 -3415 661 -3363
rect 723 -3415 724 -3363
rect 758 -3364 759 -3336
rect 772 -3364 773 -3336
rect 814 -3415 815 -3363
rect 821 -3415 822 -3363
rect 1059 -3364 1060 -3336
rect 1272 -3364 1273 -3336
rect 1283 -3415 1284 -3363
rect 1290 -3364 1291 -3336
rect 1297 -3415 1298 -3363
rect 289 -3366 290 -3336
rect 345 -3415 346 -3365
rect 387 -3366 388 -3336
rect 450 -3415 451 -3365
rect 583 -3415 584 -3365
rect 667 -3366 668 -3336
rect 737 -3366 738 -3336
rect 961 -3415 962 -3365
rect 978 -3366 979 -3336
rect 1024 -3366 1025 -3336
rect 1045 -3415 1046 -3365
rect 1143 -3366 1144 -3336
rect 1255 -3366 1256 -3336
rect 1290 -3415 1291 -3365
rect 219 -3368 220 -3336
rect 387 -3415 388 -3367
rect 443 -3368 444 -3336
rect 730 -3415 731 -3367
rect 751 -3368 752 -3336
rect 1094 -3368 1095 -3336
rect 1192 -3368 1193 -3336
rect 1255 -3415 1256 -3367
rect 352 -3370 353 -3336
rect 667 -3415 668 -3369
rect 772 -3415 773 -3369
rect 800 -3370 801 -3336
rect 835 -3370 836 -3336
rect 849 -3370 850 -3336
rect 852 -3370 853 -3336
rect 1010 -3370 1011 -3336
rect 1024 -3415 1025 -3369
rect 1038 -3370 1039 -3336
rect 1059 -3415 1060 -3369
rect 1073 -3370 1074 -3336
rect 1094 -3415 1095 -3369
rect 1241 -3370 1242 -3336
rect 401 -3372 402 -3336
rect 443 -3415 444 -3371
rect 471 -3372 472 -3336
rect 737 -3415 738 -3371
rect 779 -3415 780 -3371
rect 975 -3372 976 -3336
rect 982 -3372 983 -3336
rect 1104 -3372 1105 -3336
rect 1192 -3415 1193 -3371
rect 1465 -3372 1466 -3336
rect 401 -3415 402 -3373
rect 751 -3415 752 -3373
rect 793 -3374 794 -3336
rect 835 -3415 836 -3373
rect 842 -3374 843 -3336
rect 957 -3374 958 -3336
rect 989 -3374 990 -3336
rect 1360 -3374 1361 -3336
rect 1465 -3415 1466 -3373
rect 1507 -3374 1508 -3336
rect 600 -3376 601 -3336
rect 1073 -3415 1074 -3375
rect 1241 -3415 1242 -3375
rect 1304 -3376 1305 -3336
rect 1346 -3376 1347 -3336
rect 1360 -3415 1361 -3375
rect 604 -3378 605 -3336
rect 758 -3415 759 -3377
rect 800 -3415 801 -3377
rect 1377 -3415 1378 -3377
rect 604 -3415 605 -3379
rect 611 -3380 612 -3336
rect 618 -3415 619 -3379
rect 709 -3380 710 -3336
rect 842 -3415 843 -3379
rect 1206 -3380 1207 -3336
rect 1318 -3380 1319 -3336
rect 1346 -3415 1347 -3379
rect 520 -3382 521 -3336
rect 709 -3415 710 -3381
rect 849 -3415 850 -3381
rect 1150 -3382 1151 -3336
rect 1185 -3382 1186 -3336
rect 1304 -3415 1305 -3381
rect 418 -3384 419 -3336
rect 520 -3415 521 -3383
rect 527 -3384 528 -3336
rect 611 -3415 612 -3383
rect 625 -3384 626 -3336
rect 653 -3415 654 -3383
rect 688 -3384 689 -3336
rect 793 -3415 794 -3383
rect 856 -3384 857 -3336
rect 982 -3415 983 -3383
rect 989 -3415 990 -3383
rect 1248 -3384 1249 -3336
rect 457 -3386 458 -3336
rect 625 -3415 626 -3385
rect 688 -3415 689 -3385
rect 786 -3386 787 -3336
rect 870 -3386 871 -3336
rect 975 -3415 976 -3385
rect 1108 -3386 1109 -3336
rect 1206 -3415 1207 -3385
rect 1209 -3415 1210 -3385
rect 1248 -3415 1249 -3385
rect 310 -3388 311 -3336
rect 457 -3415 458 -3387
rect 527 -3415 528 -3387
rect 569 -3388 570 -3336
rect 786 -3415 787 -3387
rect 884 -3388 885 -3336
rect 891 -3415 892 -3387
rect 1122 -3388 1123 -3336
rect 1185 -3415 1186 -3387
rect 1479 -3388 1480 -3336
rect 184 -3390 185 -3336
rect 569 -3415 570 -3389
rect 807 -3390 808 -3336
rect 1108 -3415 1109 -3389
rect 1122 -3415 1123 -3389
rect 1381 -3415 1382 -3389
rect 261 -3392 262 -3336
rect 310 -3415 311 -3391
rect 695 -3392 696 -3336
rect 807 -3415 808 -3391
rect 863 -3392 864 -3336
rect 884 -3415 885 -3391
rect 898 -3392 899 -3336
rect 1038 -3415 1039 -3391
rect 324 -3394 325 -3336
rect 695 -3415 696 -3393
rect 744 -3394 745 -3336
rect 863 -3415 864 -3393
rect 870 -3415 871 -3393
rect 905 -3394 906 -3336
rect 919 -3394 920 -3336
rect 1010 -3415 1011 -3393
rect 702 -3396 703 -3336
rect 744 -3415 745 -3395
rect 901 -3415 902 -3395
rect 1276 -3396 1277 -3336
rect 464 -3398 465 -3336
rect 702 -3415 703 -3397
rect 905 -3415 906 -3397
rect 1115 -3398 1116 -3336
rect 436 -3400 437 -3336
rect 464 -3415 465 -3399
rect 912 -3400 913 -3336
rect 919 -3415 920 -3399
rect 926 -3415 927 -3399
rect 1129 -3400 1130 -3336
rect 380 -3402 381 -3336
rect 436 -3415 437 -3401
rect 765 -3402 766 -3336
rect 912 -3415 913 -3401
rect 940 -3402 941 -3336
rect 1143 -3415 1144 -3401
rect 247 -3404 248 -3336
rect 380 -3415 381 -3403
rect 632 -3404 633 -3336
rect 765 -3415 766 -3403
rect 940 -3415 941 -3403
rect 1216 -3404 1217 -3336
rect 499 -3406 500 -3336
rect 632 -3415 633 -3405
rect 947 -3406 948 -3336
rect 1136 -3415 1137 -3405
rect 338 -3408 339 -3336
rect 499 -3415 500 -3407
rect 828 -3408 829 -3336
rect 947 -3415 948 -3407
rect 954 -3415 955 -3407
rect 996 -3408 997 -3336
rect 1052 -3408 1053 -3336
rect 1115 -3415 1116 -3407
rect 191 -3410 192 -3336
rect 338 -3415 339 -3409
rect 828 -3415 829 -3409
rect 933 -3410 934 -3336
rect 996 -3415 997 -3409
rect 1171 -3410 1172 -3336
rect 933 -3415 934 -3411
rect 1017 -3412 1018 -3336
rect 1052 -3415 1053 -3411
rect 1087 -3412 1088 -3336
rect 1171 -3415 1172 -3411
rect 1262 -3412 1263 -3336
rect 971 -3414 972 -3336
rect 1017 -3415 1018 -3413
rect 1087 -3415 1088 -3413
rect 1164 -3414 1165 -3336
rect 1262 -3415 1263 -3413
rect 1409 -3414 1410 -3336
rect 173 -3425 174 -3423
rect 268 -3460 269 -3424
rect 296 -3425 297 -3423
rect 317 -3425 318 -3423
rect 338 -3425 339 -3423
rect 474 -3425 475 -3423
rect 478 -3425 479 -3423
rect 593 -3460 594 -3424
rect 621 -3460 622 -3424
rect 632 -3425 633 -3423
rect 639 -3425 640 -3423
rect 723 -3425 724 -3423
rect 726 -3425 727 -3423
rect 940 -3425 941 -3423
rect 961 -3425 962 -3423
rect 1206 -3425 1207 -3423
rect 1213 -3425 1214 -3423
rect 1286 -3460 1287 -3424
rect 1290 -3425 1291 -3423
rect 1290 -3460 1291 -3424
rect 1290 -3425 1291 -3423
rect 1290 -3460 1291 -3424
rect 1297 -3425 1298 -3423
rect 1307 -3425 1308 -3423
rect 1311 -3460 1312 -3424
rect 1332 -3425 1333 -3423
rect 1346 -3425 1347 -3423
rect 1374 -3425 1375 -3423
rect 1437 -3460 1438 -3424
rect 1451 -3425 1452 -3423
rect 1458 -3425 1459 -3423
rect 1493 -3460 1494 -3424
rect 1500 -3425 1501 -3423
rect 1500 -3460 1501 -3424
rect 1500 -3425 1501 -3423
rect 1500 -3460 1501 -3424
rect 1514 -3460 1515 -3424
rect 1528 -3425 1529 -3423
rect 1584 -3425 1585 -3423
rect 1808 -3425 1809 -3423
rect 1822 -3425 1823 -3423
rect 1860 -3460 1861 -3424
rect 1955 -3425 1956 -3423
rect 1955 -3460 1956 -3424
rect 1955 -3425 1956 -3423
rect 1955 -3460 1956 -3424
rect 1962 -3425 1963 -3423
rect 1962 -3460 1963 -3424
rect 1962 -3425 1963 -3423
rect 1962 -3460 1963 -3424
rect 2025 -3425 2026 -3423
rect 2025 -3460 2026 -3424
rect 2025 -3425 2026 -3423
rect 2025 -3460 2026 -3424
rect 2032 -3425 2033 -3423
rect 2032 -3460 2033 -3424
rect 2032 -3425 2033 -3423
rect 2032 -3460 2033 -3424
rect 170 -3427 171 -3423
rect 173 -3460 174 -3426
rect 310 -3427 311 -3423
rect 324 -3460 325 -3426
rect 345 -3427 346 -3423
rect 390 -3427 391 -3423
rect 394 -3427 395 -3423
rect 401 -3427 402 -3423
rect 404 -3427 405 -3423
rect 415 -3460 416 -3426
rect 429 -3427 430 -3423
rect 467 -3460 468 -3426
rect 492 -3427 493 -3423
rect 628 -3460 629 -3426
rect 646 -3427 647 -3423
rect 723 -3460 724 -3426
rect 758 -3427 759 -3423
rect 800 -3460 801 -3426
rect 807 -3427 808 -3423
rect 842 -3427 843 -3423
rect 884 -3427 885 -3423
rect 922 -3427 923 -3423
rect 975 -3427 976 -3423
rect 1024 -3460 1025 -3426
rect 1038 -3427 1039 -3423
rect 1038 -3460 1039 -3426
rect 1038 -3427 1039 -3423
rect 1038 -3460 1039 -3426
rect 1066 -3427 1067 -3423
rect 1199 -3427 1200 -3423
rect 1206 -3460 1207 -3426
rect 1234 -3427 1235 -3423
rect 1248 -3427 1249 -3423
rect 1307 -3460 1308 -3426
rect 1321 -3460 1322 -3426
rect 1332 -3460 1333 -3426
rect 1360 -3427 1361 -3423
rect 1360 -3460 1361 -3426
rect 1360 -3427 1361 -3423
rect 1360 -3460 1361 -3426
rect 1444 -3460 1445 -3426
rect 1465 -3427 1466 -3423
rect 1521 -3427 1522 -3423
rect 1521 -3460 1522 -3426
rect 1521 -3427 1522 -3423
rect 1521 -3460 1522 -3426
rect 1612 -3427 1613 -3423
rect 1629 -3460 1630 -3426
rect 1640 -3460 1641 -3426
rect 1647 -3427 1648 -3423
rect 1724 -3427 1725 -3423
rect 1727 -3435 1728 -3426
rect 1738 -3427 1739 -3423
rect 1748 -3460 1749 -3426
rect 1759 -3427 1760 -3423
rect 1766 -3427 1767 -3423
rect 1780 -3427 1781 -3423
rect 1780 -3460 1781 -3426
rect 1780 -3427 1781 -3423
rect 1780 -3460 1781 -3426
rect 1794 -3460 1795 -3426
rect 1801 -3427 1802 -3423
rect 1822 -3460 1823 -3426
rect 1829 -3427 1830 -3423
rect 1850 -3427 1851 -3423
rect 1850 -3460 1851 -3426
rect 1850 -3427 1851 -3423
rect 1850 -3460 1851 -3426
rect 1857 -3427 1858 -3423
rect 1867 -3427 1868 -3423
rect 373 -3429 374 -3423
rect 471 -3429 472 -3423
rect 492 -3460 493 -3428
rect 562 -3429 563 -3423
rect 576 -3429 577 -3423
rect 576 -3460 577 -3428
rect 576 -3429 577 -3423
rect 576 -3460 577 -3428
rect 611 -3429 612 -3423
rect 639 -3460 640 -3428
rect 653 -3429 654 -3423
rect 656 -3435 657 -3428
rect 684 -3460 685 -3428
rect 716 -3429 717 -3423
rect 744 -3429 745 -3423
rect 758 -3460 759 -3428
rect 793 -3429 794 -3423
rect 793 -3460 794 -3428
rect 793 -3429 794 -3423
rect 793 -3460 794 -3428
rect 807 -3460 808 -3428
rect 989 -3429 990 -3423
rect 992 -3429 993 -3423
rect 1052 -3429 1053 -3423
rect 1066 -3460 1067 -3428
rect 1101 -3429 1102 -3423
rect 1108 -3429 1109 -3423
rect 1199 -3460 1200 -3428
rect 1220 -3429 1221 -3423
rect 1458 -3460 1459 -3428
rect 1461 -3460 1462 -3428
rect 1654 -3429 1655 -3423
rect 1724 -3460 1725 -3428
rect 1731 -3429 1732 -3423
rect 1766 -3460 1767 -3428
rect 1787 -3429 1788 -3423
rect 1829 -3460 1830 -3428
rect 1843 -3429 1844 -3423
rect 1857 -3460 1858 -3428
rect 1864 -3429 1865 -3423
rect 408 -3431 409 -3423
rect 488 -3431 489 -3423
rect 499 -3431 500 -3423
rect 611 -3460 612 -3430
rect 625 -3431 626 -3423
rect 667 -3460 668 -3430
rect 695 -3431 696 -3423
rect 1031 -3431 1032 -3423
rect 1052 -3460 1053 -3430
rect 1087 -3431 1088 -3423
rect 1101 -3460 1102 -3430
rect 1185 -3431 1186 -3423
rect 1255 -3431 1256 -3423
rect 1318 -3460 1319 -3430
rect 1325 -3460 1326 -3430
rect 1367 -3431 1368 -3423
rect 1381 -3431 1382 -3423
rect 1465 -3460 1466 -3430
rect 1836 -3431 1837 -3423
rect 1843 -3460 1844 -3430
rect 1864 -3460 1865 -3430
rect 1871 -3431 1872 -3423
rect 450 -3433 451 -3423
rect 485 -3460 486 -3432
rect 506 -3433 507 -3423
rect 646 -3460 647 -3432
rect 653 -3460 654 -3432
rect 702 -3433 703 -3423
rect 922 -3460 923 -3432
rect 1003 -3433 1004 -3423
rect 1031 -3460 1032 -3432
rect 1069 -3433 1070 -3423
rect 1125 -3433 1126 -3423
rect 1136 -3433 1137 -3423
rect 1220 -3460 1221 -3432
rect 1276 -3433 1277 -3423
rect 1283 -3433 1284 -3423
rect 1451 -3460 1452 -3432
rect 1472 -3433 1473 -3423
rect 422 -3435 423 -3423
rect 506 -3460 507 -3434
rect 534 -3435 535 -3423
rect 534 -3460 535 -3434
rect 534 -3435 535 -3423
rect 534 -3460 535 -3434
rect 548 -3435 549 -3423
rect 579 -3460 580 -3434
rect 660 -3435 661 -3423
rect 695 -3460 696 -3434
rect 702 -3460 703 -3434
rect 786 -3435 787 -3423
rect 814 -3435 815 -3423
rect 845 -3435 846 -3423
rect 863 -3435 864 -3423
rect 884 -3460 885 -3434
rect 901 -3435 902 -3423
rect 1094 -3435 1095 -3423
rect 1108 -3460 1109 -3434
rect 1192 -3435 1193 -3423
rect 1867 -3460 1868 -3434
rect 1871 -3460 1872 -3434
rect 380 -3437 381 -3423
rect 422 -3460 423 -3436
rect 464 -3437 465 -3423
rect 499 -3460 500 -3436
rect 555 -3437 556 -3423
rect 604 -3437 605 -3423
rect 660 -3460 661 -3436
rect 705 -3460 706 -3436
rect 709 -3437 710 -3423
rect 898 -3437 899 -3423
rect 912 -3437 913 -3423
rect 975 -3460 976 -3436
rect 1010 -3437 1011 -3423
rect 1122 -3437 1123 -3423
rect 1143 -3437 1144 -3423
rect 1234 -3460 1235 -3436
rect 331 -3439 332 -3423
rect 464 -3460 465 -3438
rect 541 -3439 542 -3423
rect 555 -3460 556 -3438
rect 558 -3439 559 -3423
rect 779 -3439 780 -3423
rect 814 -3460 815 -3438
rect 828 -3439 829 -3423
rect 835 -3439 836 -3423
rect 859 -3439 860 -3423
rect 915 -3460 916 -3438
rect 968 -3439 969 -3423
rect 982 -3439 983 -3423
rect 1010 -3460 1011 -3438
rect 1017 -3439 1018 -3423
rect 1017 -3460 1018 -3438
rect 1017 -3439 1018 -3423
rect 1017 -3460 1018 -3438
rect 1034 -3439 1035 -3423
rect 1094 -3460 1095 -3438
rect 1115 -3439 1116 -3423
rect 1181 -3460 1182 -3438
rect 1185 -3460 1186 -3438
rect 1262 -3439 1263 -3423
rect 359 -3441 360 -3423
rect 380 -3460 381 -3440
rect 541 -3460 542 -3440
rect 618 -3441 619 -3423
rect 674 -3441 675 -3423
rect 709 -3460 710 -3440
rect 737 -3441 738 -3423
rect 828 -3460 829 -3440
rect 835 -3460 836 -3440
rect 870 -3441 871 -3423
rect 919 -3441 920 -3423
rect 954 -3441 955 -3423
rect 1073 -3441 1074 -3423
rect 1248 -3460 1249 -3440
rect 562 -3460 563 -3442
rect 597 -3443 598 -3423
rect 604 -3460 605 -3442
rect 625 -3460 626 -3442
rect 681 -3443 682 -3423
rect 737 -3460 738 -3442
rect 744 -3460 745 -3442
rect 821 -3443 822 -3423
rect 842 -3460 843 -3442
rect 891 -3443 892 -3423
rect 947 -3443 948 -3423
rect 1003 -3460 1004 -3442
rect 1059 -3443 1060 -3423
rect 1073 -3460 1074 -3442
rect 1080 -3443 1081 -3423
rect 1129 -3460 1130 -3442
rect 1157 -3443 1158 -3423
rect 1157 -3460 1158 -3442
rect 1157 -3443 1158 -3423
rect 1157 -3460 1158 -3442
rect 1164 -3460 1165 -3442
rect 1626 -3460 1627 -3442
rect 520 -3445 521 -3423
rect 681 -3460 682 -3444
rect 751 -3445 752 -3423
rect 1125 -3460 1126 -3444
rect 1192 -3460 1193 -3444
rect 1241 -3445 1242 -3423
rect 436 -3447 437 -3423
rect 520 -3460 521 -3446
rect 569 -3447 570 -3423
rect 716 -3460 717 -3446
rect 751 -3460 752 -3446
rect 849 -3447 850 -3423
rect 877 -3447 878 -3423
rect 1080 -3460 1081 -3446
rect 1083 -3460 1084 -3446
rect 1171 -3447 1172 -3423
rect 1227 -3447 1228 -3423
rect 1241 -3460 1242 -3446
rect 527 -3449 528 -3423
rect 569 -3460 570 -3448
rect 583 -3449 584 -3423
rect 597 -3460 598 -3448
rect 632 -3460 633 -3448
rect 1059 -3460 1060 -3448
rect 1087 -3460 1088 -3448
rect 1304 -3460 1305 -3448
rect 513 -3451 514 -3423
rect 583 -3460 584 -3450
rect 590 -3451 591 -3423
rect 674 -3460 675 -3450
rect 730 -3451 731 -3423
rect 849 -3460 850 -3450
rect 877 -3460 878 -3450
rect 905 -3451 906 -3423
rect 954 -3460 955 -3450
rect 996 -3451 997 -3423
rect 1171 -3460 1172 -3450
rect 1269 -3451 1270 -3423
rect 457 -3453 458 -3423
rect 513 -3460 514 -3452
rect 730 -3460 731 -3452
rect 926 -3453 927 -3423
rect 996 -3460 997 -3452
rect 1045 -3453 1046 -3423
rect 1178 -3453 1179 -3423
rect 1227 -3460 1228 -3452
rect 443 -3455 444 -3423
rect 457 -3460 458 -3454
rect 590 -3460 591 -3454
rect 1045 -3460 1046 -3454
rect 1178 -3460 1179 -3454
rect 1213 -3460 1214 -3454
rect 439 -3457 440 -3423
rect 443 -3460 444 -3456
rect 765 -3457 766 -3423
rect 821 -3460 822 -3456
rect 772 -3459 773 -3423
rect 779 -3460 780 -3458
rect 271 -3470 272 -3468
rect 366 -3489 367 -3469
rect 369 -3489 370 -3469
rect 394 -3489 395 -3469
rect 415 -3470 416 -3468
rect 429 -3489 430 -3469
rect 439 -3470 440 -3468
rect 443 -3470 444 -3468
rect 457 -3470 458 -3468
rect 464 -3489 465 -3469
rect 478 -3489 479 -3469
rect 492 -3470 493 -3468
rect 499 -3470 500 -3468
rect 551 -3470 552 -3468
rect 569 -3470 570 -3468
rect 639 -3470 640 -3468
rect 642 -3470 643 -3468
rect 751 -3470 752 -3468
rect 765 -3489 766 -3469
rect 807 -3470 808 -3468
rect 828 -3470 829 -3468
rect 912 -3470 913 -3468
rect 919 -3470 920 -3468
rect 954 -3470 955 -3468
rect 975 -3470 976 -3468
rect 978 -3474 979 -3469
rect 1031 -3470 1032 -3468
rect 1062 -3470 1063 -3468
rect 1066 -3470 1067 -3468
rect 1066 -3489 1067 -3469
rect 1066 -3470 1067 -3468
rect 1066 -3489 1067 -3469
rect 1080 -3489 1081 -3469
rect 1108 -3470 1109 -3468
rect 1122 -3470 1123 -3468
rect 1185 -3470 1186 -3468
rect 1199 -3470 1200 -3468
rect 1318 -3470 1319 -3468
rect 1360 -3470 1361 -3468
rect 1360 -3489 1361 -3469
rect 1360 -3470 1361 -3468
rect 1360 -3489 1361 -3469
rect 1430 -3489 1431 -3469
rect 1444 -3470 1445 -3468
rect 1458 -3470 1459 -3468
rect 1570 -3489 1571 -3469
rect 1640 -3470 1641 -3468
rect 1640 -3489 1641 -3469
rect 1640 -3470 1641 -3468
rect 1640 -3489 1641 -3469
rect 1724 -3470 1725 -3468
rect 1724 -3489 1725 -3469
rect 1724 -3470 1725 -3468
rect 1724 -3489 1725 -3469
rect 1731 -3470 1732 -3468
rect 1731 -3489 1732 -3469
rect 1731 -3470 1732 -3468
rect 1731 -3489 1732 -3469
rect 1745 -3470 1746 -3468
rect 1766 -3470 1767 -3468
rect 1780 -3470 1781 -3468
rect 1780 -3489 1781 -3469
rect 1780 -3470 1781 -3468
rect 1780 -3489 1781 -3469
rect 1790 -3489 1791 -3469
rect 1794 -3470 1795 -3468
rect 1829 -3470 1830 -3468
rect 1836 -3470 1837 -3468
rect 1839 -3470 1840 -3468
rect 1850 -3470 1851 -3468
rect 1860 -3470 1861 -3468
rect 1864 -3470 1865 -3468
rect 1955 -3470 1956 -3468
rect 1955 -3489 1956 -3469
rect 1955 -3470 1956 -3468
rect 1955 -3489 1956 -3469
rect 1958 -3489 1959 -3469
rect 1962 -3470 1963 -3468
rect 2025 -3470 2026 -3468
rect 2028 -3470 2029 -3468
rect 324 -3472 325 -3468
rect 331 -3489 332 -3471
rect 380 -3472 381 -3468
rect 387 -3489 388 -3471
rect 422 -3472 423 -3468
rect 467 -3472 468 -3468
rect 485 -3472 486 -3468
rect 523 -3472 524 -3468
rect 541 -3472 542 -3468
rect 569 -3489 570 -3471
rect 579 -3472 580 -3468
rect 604 -3472 605 -3468
rect 618 -3489 619 -3471
rect 628 -3472 629 -3468
rect 639 -3489 640 -3471
rect 653 -3472 654 -3468
rect 667 -3472 668 -3468
rect 705 -3472 706 -3468
rect 730 -3472 731 -3468
rect 737 -3472 738 -3468
rect 772 -3489 773 -3471
rect 779 -3472 780 -3468
rect 789 -3489 790 -3471
rect 814 -3472 815 -3468
rect 828 -3489 829 -3471
rect 842 -3472 843 -3468
rect 849 -3472 850 -3468
rect 922 -3472 923 -3468
rect 975 -3489 976 -3471
rect 1017 -3472 1018 -3468
rect 1031 -3489 1032 -3471
rect 1052 -3472 1053 -3468
rect 1052 -3489 1053 -3471
rect 1052 -3472 1053 -3468
rect 1052 -3489 1053 -3471
rect 1059 -3472 1060 -3468
rect 1073 -3472 1074 -3468
rect 1083 -3472 1084 -3468
rect 1171 -3472 1172 -3468
rect 1178 -3472 1179 -3468
rect 1206 -3472 1207 -3468
rect 1213 -3472 1214 -3468
rect 1272 -3489 1273 -3471
rect 1276 -3489 1277 -3471
rect 1286 -3489 1287 -3471
rect 1307 -3472 1308 -3468
rect 1311 -3472 1312 -3468
rect 1433 -3489 1434 -3471
rect 1451 -3472 1452 -3468
rect 1500 -3472 1501 -3468
rect 1503 -3489 1504 -3471
rect 1507 -3489 1508 -3471
rect 1514 -3472 1515 -3468
rect 1521 -3472 1522 -3468
rect 1521 -3489 1522 -3471
rect 1521 -3472 1522 -3468
rect 1521 -3489 1522 -3471
rect 1843 -3472 1844 -3468
rect 1850 -3489 1851 -3471
rect 1864 -3489 1865 -3471
rect 1871 -3472 1872 -3468
rect 2025 -3489 2026 -3471
rect 2032 -3472 2033 -3468
rect 471 -3489 472 -3473
rect 523 -3489 524 -3473
rect 562 -3474 563 -3468
rect 604 -3489 605 -3473
rect 646 -3474 647 -3468
rect 646 -3489 647 -3473
rect 646 -3474 647 -3468
rect 646 -3489 647 -3473
rect 653 -3489 654 -3473
rect 744 -3474 745 -3468
rect 793 -3474 794 -3468
rect 793 -3489 794 -3473
rect 793 -3474 794 -3468
rect 793 -3489 794 -3473
rect 800 -3474 801 -3468
rect 887 -3489 888 -3473
rect 1010 -3474 1011 -3468
rect 1017 -3489 1018 -3473
rect 1045 -3474 1046 -3468
rect 1500 -3489 1501 -3473
rect 1822 -3474 1823 -3468
rect 1843 -3489 1844 -3473
rect 2028 -3489 2029 -3473
rect 2032 -3489 2033 -3473
rect 485 -3489 486 -3475
rect 632 -3476 633 -3468
rect 674 -3476 675 -3468
rect 702 -3476 703 -3468
rect 709 -3476 710 -3468
rect 744 -3489 745 -3475
rect 814 -3489 815 -3475
rect 835 -3476 836 -3468
rect 866 -3489 867 -3475
rect 1087 -3476 1088 -3468
rect 1094 -3476 1095 -3468
rect 1125 -3476 1126 -3468
rect 1129 -3476 1130 -3468
rect 1143 -3489 1144 -3475
rect 1178 -3489 1179 -3475
rect 1192 -3476 1193 -3468
rect 1234 -3476 1235 -3468
rect 1262 -3489 1263 -3475
rect 1269 -3489 1270 -3475
rect 1325 -3476 1326 -3468
rect 1437 -3476 1438 -3468
rect 1437 -3489 1438 -3475
rect 1437 -3476 1438 -3468
rect 1437 -3489 1438 -3475
rect 1493 -3476 1494 -3468
rect 1514 -3489 1515 -3475
rect 506 -3478 507 -3468
rect 541 -3489 542 -3477
rect 583 -3478 584 -3468
rect 583 -3489 584 -3477
rect 583 -3478 584 -3468
rect 583 -3489 584 -3477
rect 590 -3478 591 -3468
rect 597 -3478 598 -3468
rect 632 -3489 633 -3477
rect 660 -3478 661 -3468
rect 681 -3478 682 -3468
rect 751 -3489 752 -3477
rect 821 -3478 822 -3468
rect 842 -3489 843 -3477
rect 870 -3489 871 -3477
rect 877 -3478 878 -3468
rect 884 -3478 885 -3468
rect 915 -3478 916 -3468
rect 1003 -3478 1004 -3468
rect 1010 -3489 1011 -3477
rect 1038 -3478 1039 -3468
rect 1045 -3489 1046 -3477
rect 1059 -3489 1060 -3477
rect 1101 -3478 1102 -3468
rect 1157 -3478 1158 -3468
rect 1192 -3489 1193 -3477
rect 1220 -3478 1221 -3468
rect 1234 -3489 1235 -3477
rect 1255 -3489 1256 -3477
rect 1304 -3478 1305 -3468
rect 1311 -3489 1312 -3477
rect 1332 -3478 1333 -3468
rect 1465 -3478 1466 -3468
rect 1493 -3489 1494 -3477
rect 520 -3480 521 -3468
rect 898 -3489 899 -3479
rect 1024 -3480 1025 -3468
rect 1038 -3489 1039 -3479
rect 1248 -3480 1249 -3468
rect 1304 -3489 1305 -3479
rect 534 -3482 535 -3468
rect 590 -3489 591 -3481
rect 611 -3482 612 -3468
rect 681 -3489 682 -3481
rect 695 -3482 696 -3468
rect 786 -3489 787 -3481
rect 1024 -3489 1025 -3481
rect 1164 -3482 1165 -3468
rect 1241 -3482 1242 -3468
rect 1248 -3489 1249 -3481
rect 1283 -3482 1284 -3468
rect 1290 -3482 1291 -3468
rect 513 -3484 514 -3468
rect 534 -3489 535 -3483
rect 555 -3484 556 -3468
rect 611 -3489 612 -3483
rect 716 -3484 717 -3468
rect 779 -3489 780 -3483
rect 1227 -3484 1228 -3468
rect 1241 -3489 1242 -3483
rect 1290 -3489 1291 -3483
rect 1727 -3489 1728 -3483
rect 688 -3486 689 -3468
rect 716 -3489 717 -3485
rect 737 -3489 738 -3485
rect 758 -3486 759 -3468
rect 723 -3488 724 -3468
rect 758 -3489 759 -3487
rect 331 -3499 332 -3497
rect 338 -3512 339 -3498
rect 394 -3499 395 -3497
rect 429 -3499 430 -3497
rect 432 -3499 433 -3497
rect 471 -3499 472 -3497
rect 478 -3499 479 -3497
rect 478 -3512 479 -3498
rect 478 -3499 479 -3497
rect 478 -3512 479 -3498
rect 523 -3499 524 -3497
rect 653 -3499 654 -3497
rect 681 -3499 682 -3497
rect 709 -3512 710 -3498
rect 716 -3499 717 -3497
rect 730 -3512 731 -3498
rect 737 -3499 738 -3497
rect 737 -3512 738 -3498
rect 737 -3499 738 -3497
rect 737 -3512 738 -3498
rect 775 -3512 776 -3498
rect 891 -3512 892 -3498
rect 968 -3512 969 -3498
rect 975 -3499 976 -3497
rect 996 -3499 997 -3497
rect 1003 -3512 1004 -3498
rect 1010 -3499 1011 -3497
rect 1010 -3512 1011 -3498
rect 1010 -3499 1011 -3497
rect 1010 -3512 1011 -3498
rect 1017 -3499 1018 -3497
rect 1017 -3512 1018 -3498
rect 1017 -3499 1018 -3497
rect 1017 -3512 1018 -3498
rect 1038 -3499 1039 -3497
rect 1062 -3512 1063 -3498
rect 1122 -3512 1123 -3498
rect 1290 -3499 1291 -3497
rect 1304 -3499 1305 -3497
rect 1367 -3512 1368 -3498
rect 1430 -3499 1431 -3497
rect 1437 -3499 1438 -3497
rect 1500 -3499 1501 -3497
rect 1507 -3499 1508 -3497
rect 1514 -3499 1515 -3497
rect 1514 -3512 1515 -3498
rect 1514 -3499 1515 -3497
rect 1514 -3512 1515 -3498
rect 1521 -3499 1522 -3497
rect 1521 -3512 1522 -3498
rect 1521 -3499 1522 -3497
rect 1521 -3512 1522 -3498
rect 1570 -3499 1571 -3497
rect 1612 -3512 1613 -3498
rect 1640 -3499 1641 -3497
rect 1640 -3512 1641 -3498
rect 1640 -3499 1641 -3497
rect 1640 -3512 1641 -3498
rect 1724 -3499 1725 -3497
rect 1731 -3499 1732 -3497
rect 1780 -3499 1781 -3497
rect 1790 -3499 1791 -3497
rect 1850 -3499 1851 -3497
rect 1860 -3512 1861 -3498
rect 2025 -3499 2026 -3497
rect 2025 -3512 2026 -3498
rect 2025 -3499 2026 -3497
rect 2025 -3512 2026 -3498
rect 2032 -3499 2033 -3497
rect 2032 -3512 2033 -3498
rect 2032 -3499 2033 -3497
rect 2032 -3512 2033 -3498
rect 387 -3501 388 -3497
rect 394 -3512 395 -3500
rect 429 -3512 430 -3500
rect 485 -3501 486 -3497
rect 534 -3501 535 -3497
rect 548 -3512 549 -3500
rect 569 -3501 570 -3497
rect 576 -3512 577 -3500
rect 583 -3501 584 -3497
rect 583 -3512 584 -3500
rect 583 -3501 584 -3497
rect 583 -3512 584 -3500
rect 625 -3512 626 -3500
rect 632 -3501 633 -3497
rect 639 -3501 640 -3497
rect 639 -3512 640 -3500
rect 639 -3501 640 -3497
rect 639 -3512 640 -3500
rect 646 -3501 647 -3497
rect 656 -3501 657 -3497
rect 779 -3501 780 -3497
rect 800 -3512 801 -3500
rect 810 -3512 811 -3500
rect 828 -3501 829 -3497
rect 842 -3501 843 -3497
rect 866 -3501 867 -3497
rect 884 -3501 885 -3497
rect 1024 -3501 1025 -3497
rect 1038 -3512 1039 -3500
rect 1045 -3501 1046 -3497
rect 1052 -3501 1053 -3497
rect 1052 -3512 1053 -3500
rect 1052 -3501 1053 -3497
rect 1052 -3512 1053 -3500
rect 1143 -3501 1144 -3497
rect 1150 -3512 1151 -3500
rect 1160 -3512 1161 -3500
rect 1178 -3501 1179 -3497
rect 1192 -3501 1193 -3497
rect 1206 -3512 1207 -3500
rect 1234 -3501 1235 -3497
rect 1251 -3501 1252 -3497
rect 1262 -3501 1263 -3497
rect 1276 -3501 1277 -3497
rect 1283 -3501 1284 -3497
rect 1311 -3501 1312 -3497
rect 1360 -3501 1361 -3497
rect 1360 -3512 1361 -3500
rect 1360 -3501 1361 -3497
rect 1360 -3512 1361 -3500
rect 1493 -3501 1494 -3497
rect 1507 -3512 1508 -3500
rect 1843 -3501 1844 -3497
rect 1850 -3512 1851 -3500
rect 1857 -3512 1858 -3500
rect 1864 -3501 1865 -3497
rect 464 -3503 465 -3497
rect 464 -3512 465 -3502
rect 464 -3503 465 -3497
rect 464 -3512 465 -3502
rect 541 -3503 542 -3497
rect 541 -3512 542 -3502
rect 541 -3503 542 -3497
rect 541 -3512 542 -3502
rect 611 -3503 612 -3497
rect 632 -3512 633 -3502
rect 751 -3503 752 -3497
rect 779 -3512 780 -3502
rect 789 -3512 790 -3502
rect 814 -3503 815 -3497
rect 863 -3503 864 -3497
rect 870 -3503 871 -3497
rect 898 -3503 899 -3497
rect 1024 -3512 1025 -3502
rect 1031 -3503 1032 -3497
rect 1045 -3512 1046 -3502
rect 1234 -3512 1235 -3502
rect 1255 -3503 1256 -3497
rect 611 -3512 612 -3504
rect 618 -3505 619 -3497
rect 751 -3512 752 -3504
rect 758 -3505 759 -3497
rect 793 -3505 794 -3497
rect 793 -3512 794 -3504
rect 793 -3505 794 -3497
rect 793 -3512 794 -3504
rect 1031 -3512 1032 -3504
rect 1059 -3505 1060 -3497
rect 1241 -3505 1242 -3497
rect 1248 -3505 1249 -3497
rect 604 -3507 605 -3497
rect 618 -3512 619 -3506
rect 744 -3507 745 -3497
rect 758 -3512 759 -3506
rect 1059 -3512 1060 -3506
rect 1066 -3507 1067 -3497
rect 590 -3509 591 -3497
rect 604 -3512 605 -3508
rect 744 -3512 745 -3508
rect 765 -3509 766 -3497
rect 1066 -3512 1067 -3508
rect 1080 -3509 1081 -3497
rect 765 -3512 766 -3510
rect 772 -3511 773 -3497
rect 394 -3522 395 -3520
rect 394 -3531 395 -3521
rect 394 -3522 395 -3520
rect 394 -3531 395 -3521
rect 408 -3531 409 -3521
rect 429 -3522 430 -3520
rect 464 -3522 465 -3520
rect 464 -3531 465 -3521
rect 464 -3522 465 -3520
rect 464 -3531 465 -3521
rect 478 -3522 479 -3520
rect 478 -3531 479 -3521
rect 478 -3522 479 -3520
rect 478 -3531 479 -3521
rect 541 -3522 542 -3520
rect 541 -3531 542 -3521
rect 541 -3522 542 -3520
rect 541 -3531 542 -3521
rect 548 -3522 549 -3520
rect 548 -3531 549 -3521
rect 548 -3522 549 -3520
rect 548 -3531 549 -3521
rect 576 -3522 577 -3520
rect 576 -3531 577 -3521
rect 576 -3522 577 -3520
rect 576 -3531 577 -3521
rect 583 -3522 584 -3520
rect 583 -3531 584 -3521
rect 583 -3522 584 -3520
rect 583 -3531 584 -3521
rect 618 -3522 619 -3520
rect 635 -3531 636 -3521
rect 639 -3522 640 -3520
rect 639 -3531 640 -3521
rect 639 -3522 640 -3520
rect 639 -3531 640 -3521
rect 709 -3522 710 -3520
rect 716 -3531 717 -3521
rect 723 -3531 724 -3521
rect 737 -3522 738 -3520
rect 744 -3522 745 -3520
rect 744 -3531 745 -3521
rect 744 -3522 745 -3520
rect 744 -3531 745 -3521
rect 751 -3522 752 -3520
rect 786 -3522 787 -3520
rect 793 -3522 794 -3520
rect 793 -3531 794 -3521
rect 793 -3522 794 -3520
rect 793 -3531 794 -3521
rect 800 -3522 801 -3520
rect 810 -3522 811 -3520
rect 891 -3522 892 -3520
rect 926 -3531 927 -3521
rect 968 -3522 969 -3520
rect 971 -3531 972 -3521
rect 1017 -3522 1018 -3520
rect 1027 -3531 1028 -3521
rect 1031 -3522 1032 -3520
rect 1031 -3531 1032 -3521
rect 1031 -3522 1032 -3520
rect 1031 -3531 1032 -3521
rect 1038 -3522 1039 -3520
rect 1041 -3528 1042 -3521
rect 1059 -3522 1060 -3520
rect 1066 -3522 1067 -3520
rect 1150 -3522 1151 -3520
rect 1157 -3522 1158 -3520
rect 1206 -3522 1207 -3520
rect 1213 -3531 1214 -3521
rect 1223 -3531 1224 -3521
rect 1234 -3522 1235 -3520
rect 1360 -3522 1361 -3520
rect 1367 -3522 1368 -3520
rect 1507 -3522 1508 -3520
rect 1510 -3522 1511 -3520
rect 1521 -3522 1522 -3520
rect 1521 -3531 1522 -3521
rect 1521 -3522 1522 -3520
rect 1521 -3531 1522 -3521
rect 1612 -3522 1613 -3520
rect 1633 -3531 1634 -3521
rect 1640 -3522 1641 -3520
rect 1640 -3531 1641 -3521
rect 1640 -3522 1641 -3520
rect 1640 -3531 1641 -3521
rect 1850 -3522 1851 -3520
rect 1857 -3522 1858 -3520
rect 2025 -3522 2026 -3520
rect 2025 -3531 2026 -3521
rect 2025 -3522 2026 -3520
rect 2025 -3531 2026 -3521
rect 2032 -3522 2033 -3520
rect 2032 -3531 2033 -3521
rect 2032 -3522 2033 -3520
rect 2032 -3531 2033 -3521
rect 611 -3524 612 -3520
rect 618 -3531 619 -3523
rect 632 -3524 633 -3520
rect 646 -3531 647 -3523
rect 709 -3531 710 -3523
rect 740 -3531 741 -3523
rect 758 -3524 759 -3520
rect 775 -3524 776 -3520
rect 779 -3524 780 -3520
rect 786 -3531 787 -3523
rect 1024 -3524 1025 -3520
rect 1160 -3524 1161 -3520
rect 1507 -3531 1508 -3523
rect 1514 -3524 1515 -3520
rect 604 -3526 605 -3520
rect 611 -3531 612 -3525
rect 730 -3526 731 -3520
rect 730 -3531 731 -3525
rect 730 -3526 731 -3520
rect 730 -3531 731 -3525
rect 765 -3526 766 -3520
rect 789 -3526 790 -3520
rect 1010 -3526 1011 -3520
rect 1024 -3531 1025 -3525
rect 1038 -3531 1039 -3525
rect 1052 -3526 1053 -3520
rect 1059 -3531 1060 -3525
rect 1066 -3531 1067 -3525
rect 1122 -3526 1123 -3520
rect 604 -3531 605 -3527
rect 625 -3528 626 -3520
rect 765 -3531 766 -3527
rect 772 -3528 773 -3520
rect 1003 -3528 1004 -3520
rect 1010 -3531 1011 -3527
rect 1510 -3531 1511 -3527
rect 1514 -3531 1515 -3527
rect 625 -3531 626 -3529
rect 632 -3531 633 -3529
rect 394 -3541 395 -3539
rect 401 -3546 402 -3540
rect 408 -3541 409 -3539
rect 408 -3546 409 -3540
rect 408 -3541 409 -3539
rect 408 -3546 409 -3540
rect 464 -3541 465 -3539
rect 474 -3541 475 -3539
rect 541 -3541 542 -3539
rect 541 -3546 542 -3540
rect 541 -3541 542 -3539
rect 541 -3546 542 -3540
rect 548 -3541 549 -3539
rect 555 -3546 556 -3540
rect 583 -3541 584 -3539
rect 590 -3546 591 -3540
rect 604 -3541 605 -3539
rect 604 -3546 605 -3540
rect 604 -3541 605 -3539
rect 604 -3546 605 -3540
rect 611 -3541 612 -3539
rect 611 -3546 612 -3540
rect 611 -3541 612 -3539
rect 611 -3546 612 -3540
rect 618 -3541 619 -3539
rect 618 -3546 619 -3540
rect 618 -3541 619 -3539
rect 618 -3546 619 -3540
rect 635 -3541 636 -3539
rect 639 -3541 640 -3539
rect 646 -3541 647 -3539
rect 646 -3546 647 -3540
rect 646 -3541 647 -3539
rect 646 -3546 647 -3540
rect 702 -3546 703 -3540
rect 709 -3541 710 -3539
rect 716 -3541 717 -3539
rect 716 -3546 717 -3540
rect 716 -3541 717 -3539
rect 716 -3546 717 -3540
rect 723 -3541 724 -3539
rect 723 -3546 724 -3540
rect 723 -3541 724 -3539
rect 723 -3546 724 -3540
rect 730 -3541 731 -3539
rect 740 -3541 741 -3539
rect 758 -3546 759 -3540
rect 765 -3541 766 -3539
rect 786 -3541 787 -3539
rect 789 -3546 790 -3540
rect 793 -3541 794 -3539
rect 793 -3546 794 -3540
rect 793 -3541 794 -3539
rect 793 -3546 794 -3540
rect 926 -3541 927 -3539
rect 968 -3541 969 -3539
rect 1010 -3541 1011 -3539
rect 1020 -3546 1021 -3540
rect 1027 -3541 1028 -3539
rect 1031 -3541 1032 -3539
rect 1038 -3541 1039 -3539
rect 1045 -3541 1046 -3539
rect 1059 -3541 1060 -3539
rect 1059 -3546 1060 -3540
rect 1059 -3541 1060 -3539
rect 1059 -3546 1060 -3540
rect 1213 -3541 1214 -3539
rect 1223 -3541 1224 -3539
rect 1507 -3541 1508 -3539
rect 1510 -3545 1511 -3540
rect 1514 -3541 1515 -3539
rect 1514 -3546 1515 -3540
rect 1514 -3541 1515 -3539
rect 1514 -3546 1515 -3540
rect 1640 -3541 1641 -3539
rect 1647 -3546 1648 -3540
rect 2025 -3541 2026 -3539
rect 2025 -3546 2026 -3540
rect 2025 -3541 2026 -3539
rect 2025 -3546 2026 -3540
rect 2032 -3541 2033 -3539
rect 2032 -3546 2033 -3540
rect 2032 -3541 2033 -3539
rect 2032 -3546 2033 -3540
rect 471 -3543 472 -3539
rect 478 -3543 479 -3539
rect 576 -3543 577 -3539
rect 583 -3546 584 -3542
rect 730 -3546 731 -3542
rect 744 -3543 745 -3539
rect 1038 -3546 1039 -3542
rect 1066 -3543 1067 -3539
rect 1507 -3546 1508 -3542
rect 1521 -3543 1522 -3539
rect 1633 -3543 1634 -3539
rect 1640 -3546 1641 -3542
rect 1521 -3546 1522 -3544
rect 401 -3556 402 -3554
rect 404 -3560 405 -3555
rect 541 -3556 542 -3554
rect 548 -3556 549 -3554
rect 551 -3556 552 -3554
rect 555 -3556 556 -3554
rect 586 -3556 587 -3554
rect 590 -3556 591 -3554
rect 604 -3556 605 -3554
rect 607 -3556 608 -3554
rect 618 -3556 619 -3554
rect 618 -3561 619 -3555
rect 618 -3556 619 -3554
rect 618 -3561 619 -3555
rect 646 -3556 647 -3554
rect 649 -3561 650 -3555
rect 702 -3556 703 -3554
rect 702 -3561 703 -3555
rect 702 -3556 703 -3554
rect 702 -3561 703 -3555
rect 716 -3556 717 -3554
rect 716 -3561 717 -3555
rect 716 -3556 717 -3554
rect 716 -3561 717 -3555
rect 723 -3556 724 -3554
rect 723 -3561 724 -3555
rect 723 -3556 724 -3554
rect 723 -3561 724 -3555
rect 730 -3556 731 -3554
rect 730 -3561 731 -3555
rect 730 -3556 731 -3554
rect 730 -3561 731 -3555
rect 758 -3556 759 -3554
rect 758 -3561 759 -3555
rect 758 -3556 759 -3554
rect 758 -3561 759 -3555
rect 789 -3556 790 -3554
rect 793 -3556 794 -3554
rect 1017 -3556 1018 -3554
rect 1038 -3556 1039 -3554
rect 1059 -3556 1060 -3554
rect 1066 -3561 1067 -3555
rect 1517 -3561 1518 -3555
rect 1521 -3556 1522 -3554
rect 1640 -3556 1641 -3554
rect 1640 -3561 1641 -3555
rect 1640 -3556 1641 -3554
rect 1640 -3561 1641 -3555
rect 1647 -3556 1648 -3554
rect 1647 -3561 1648 -3555
rect 1647 -3556 1648 -3554
rect 1647 -3561 1648 -3555
rect 2025 -3556 2026 -3554
rect 2025 -3561 2026 -3555
rect 2025 -3556 2026 -3554
rect 2025 -3561 2026 -3555
rect 2028 -3561 2029 -3555
rect 2032 -3556 2033 -3554
rect 401 -3561 402 -3557
rect 604 -3561 605 -3557
rect 611 -3558 612 -3554
rect 1514 -3558 1515 -3554
rect 1521 -3561 1522 -3557
rect 607 -3561 608 -3559
rect 611 -3561 612 -3559
rect 1507 -3560 1508 -3554
rect 1514 -3561 1515 -3559
rect 401 -3571 402 -3569
rect 404 -3575 405 -3570
rect 604 -3571 605 -3569
rect 604 -3576 605 -3570
rect 604 -3571 605 -3569
rect 604 -3576 605 -3570
rect 611 -3571 612 -3569
rect 611 -3576 612 -3570
rect 611 -3571 612 -3569
rect 611 -3576 612 -3570
rect 618 -3571 619 -3569
rect 618 -3576 619 -3570
rect 618 -3571 619 -3569
rect 618 -3576 619 -3570
rect 702 -3571 703 -3569
rect 702 -3576 703 -3570
rect 702 -3571 703 -3569
rect 702 -3576 703 -3570
rect 716 -3571 717 -3569
rect 716 -3576 717 -3570
rect 716 -3571 717 -3569
rect 716 -3576 717 -3570
rect 723 -3571 724 -3569
rect 723 -3576 724 -3570
rect 723 -3571 724 -3569
rect 723 -3576 724 -3570
rect 730 -3571 731 -3569
rect 730 -3576 731 -3570
rect 730 -3571 731 -3569
rect 730 -3576 731 -3570
rect 758 -3571 759 -3569
rect 758 -3576 759 -3570
rect 758 -3571 759 -3569
rect 758 -3576 759 -3570
rect 1062 -3571 1063 -3569
rect 1066 -3571 1067 -3569
rect 1514 -3571 1515 -3569
rect 1521 -3571 1522 -3569
rect 1640 -3571 1641 -3569
rect 1640 -3576 1641 -3570
rect 1640 -3571 1641 -3569
rect 1640 -3576 1641 -3570
rect 1647 -3571 1648 -3569
rect 1647 -3576 1648 -3570
rect 1647 -3571 1648 -3569
rect 1647 -3576 1648 -3570
rect 401 -3576 402 -3572
rect 408 -3573 409 -3569
rect 408 -3576 409 -3574
rect 394 -3589 395 -3585
rect 401 -3586 402 -3584
rect 604 -3586 605 -3584
rect 604 -3589 605 -3585
rect 604 -3586 605 -3584
rect 604 -3589 605 -3585
rect 611 -3586 612 -3584
rect 611 -3589 612 -3585
rect 611 -3586 612 -3584
rect 611 -3589 612 -3585
rect 618 -3586 619 -3584
rect 621 -3589 622 -3585
rect 702 -3586 703 -3584
rect 702 -3589 703 -3585
rect 702 -3586 703 -3584
rect 702 -3589 703 -3585
rect 723 -3586 724 -3584
rect 726 -3589 727 -3585
rect 730 -3586 731 -3584
rect 730 -3589 731 -3585
rect 730 -3586 731 -3584
rect 730 -3589 731 -3585
rect 758 -3586 759 -3584
rect 758 -3589 759 -3585
rect 758 -3586 759 -3584
rect 758 -3589 759 -3585
rect 1640 -3586 1641 -3584
rect 1640 -3589 1641 -3585
rect 1640 -3586 1641 -3584
rect 1640 -3589 1641 -3585
rect 1647 -3586 1648 -3584
rect 1647 -3589 1648 -3585
rect 1647 -3586 1648 -3584
rect 1647 -3589 1648 -3585
rect 401 -3589 402 -3587
rect 408 -3588 409 -3584
rect 716 -3588 717 -3584
rect 723 -3589 724 -3587
rect 394 -3599 395 -3597
rect 394 -3600 395 -3598
rect 394 -3599 395 -3597
rect 394 -3600 395 -3598
rect 401 -3599 402 -3597
rect 401 -3600 402 -3598
rect 401 -3599 402 -3597
rect 401 -3600 402 -3598
rect 604 -3599 605 -3597
rect 604 -3600 605 -3598
rect 604 -3599 605 -3597
rect 604 -3600 605 -3598
rect 611 -3599 612 -3597
rect 611 -3600 612 -3598
rect 611 -3599 612 -3597
rect 611 -3600 612 -3598
rect 702 -3599 703 -3597
rect 702 -3600 703 -3598
rect 702 -3599 703 -3597
rect 702 -3600 703 -3598
rect 723 -3599 724 -3597
rect 730 -3599 731 -3597
rect 758 -3599 759 -3597
rect 758 -3600 759 -3598
rect 758 -3599 759 -3597
rect 758 -3600 759 -3598
rect 1640 -3599 1641 -3597
rect 1640 -3600 1641 -3598
rect 1640 -3599 1641 -3597
rect 1640 -3600 1641 -3598
rect 1647 -3599 1648 -3597
rect 1647 -3600 1648 -3598
rect 1647 -3599 1648 -3597
rect 1647 -3600 1648 -3598
rect 394 -3610 395 -3608
rect 394 -3611 395 -3609
rect 394 -3610 395 -3608
rect 394 -3611 395 -3609
rect 401 -3610 402 -3608
rect 401 -3611 402 -3609
rect 401 -3610 402 -3608
rect 401 -3611 402 -3609
rect 604 -3610 605 -3608
rect 604 -3611 605 -3609
rect 604 -3610 605 -3608
rect 604 -3611 605 -3609
rect 611 -3610 612 -3608
rect 611 -3611 612 -3609
rect 611 -3610 612 -3608
rect 611 -3611 612 -3609
rect 695 -3611 696 -3609
rect 705 -3610 706 -3608
rect 758 -3610 759 -3608
rect 758 -3611 759 -3609
rect 758 -3610 759 -3608
rect 758 -3611 759 -3609
rect 1640 -3610 1641 -3608
rect 1643 -3611 1644 -3609
rect 1647 -3610 1648 -3608
rect 1647 -3611 1648 -3609
rect 1647 -3610 1648 -3608
rect 1647 -3611 1648 -3609
rect 394 -3621 395 -3619
rect 394 -3622 395 -3620
rect 394 -3621 395 -3619
rect 394 -3622 395 -3620
rect 401 -3621 402 -3619
rect 401 -3622 402 -3620
rect 401 -3621 402 -3619
rect 401 -3622 402 -3620
rect 604 -3621 605 -3619
rect 604 -3622 605 -3620
rect 604 -3621 605 -3619
rect 604 -3622 605 -3620
rect 611 -3621 612 -3619
rect 611 -3622 612 -3620
rect 611 -3621 612 -3619
rect 611 -3622 612 -3620
rect 695 -3621 696 -3619
rect 695 -3622 696 -3620
rect 695 -3621 696 -3619
rect 695 -3622 696 -3620
rect 758 -3621 759 -3619
rect 765 -3622 766 -3620
rect 1640 -3621 1641 -3619
rect 1647 -3621 1648 -3619
rect 394 -3632 395 -3630
rect 394 -3633 395 -3631
rect 394 -3632 395 -3630
rect 394 -3633 395 -3631
rect 401 -3632 402 -3630
rect 401 -3633 402 -3631
rect 401 -3632 402 -3630
rect 401 -3633 402 -3631
rect 604 -3632 605 -3630
rect 604 -3633 605 -3631
rect 604 -3632 605 -3630
rect 604 -3633 605 -3631
rect 611 -3632 612 -3630
rect 611 -3633 612 -3631
rect 611 -3632 612 -3630
rect 611 -3633 612 -3631
rect 695 -3632 696 -3630
rect 695 -3633 696 -3631
rect 695 -3632 696 -3630
rect 695 -3633 696 -3631
rect 761 -3632 762 -3630
rect 765 -3632 766 -3630
rect 394 -3643 395 -3641
rect 394 -3644 395 -3642
rect 394 -3643 395 -3641
rect 394 -3644 395 -3642
rect 401 -3643 402 -3641
rect 401 -3644 402 -3642
rect 401 -3643 402 -3641
rect 401 -3644 402 -3642
rect 604 -3643 605 -3641
rect 604 -3644 605 -3642
rect 604 -3643 605 -3641
rect 604 -3644 605 -3642
rect 611 -3643 612 -3641
rect 611 -3644 612 -3642
rect 611 -3643 612 -3641
rect 611 -3644 612 -3642
rect 695 -3643 696 -3641
rect 695 -3644 696 -3642
rect 695 -3643 696 -3641
rect 695 -3644 696 -3642
rect 394 -3654 395 -3652
rect 397 -3658 398 -3653
rect 604 -3654 605 -3652
rect 604 -3659 605 -3653
rect 604 -3654 605 -3652
rect 604 -3659 605 -3653
rect 611 -3654 612 -3652
rect 611 -3659 612 -3653
rect 611 -3654 612 -3652
rect 611 -3659 612 -3653
rect 695 -3654 696 -3652
rect 698 -3659 699 -3653
rect 394 -3659 395 -3655
rect 401 -3656 402 -3652
rect 401 -3659 402 -3657
rect 397 -3669 398 -3667
rect 401 -3669 402 -3667
rect 604 -3669 605 -3667
rect 611 -3669 612 -3667
<< labels >>
rlabel pdiffusion 3 -24 3 -24 0 cellNo=80
rlabel pdiffusion 10 -24 10 -24 0 cellNo=143
rlabel pdiffusion 17 -24 17 -24 0 cellNo=1080
rlabel pdiffusion 24 -24 24 -24 0 cellNo=1007
rlabel pdiffusion 31 -24 31 -24 0 cellNo=1002
rlabel pdiffusion 38 -24 38 -24 0 cellNo=1006
rlabel pdiffusion 45 -24 45 -24 0 cellNo=1009
rlabel pdiffusion 52 -24 52 -24 0 cellNo=1041
rlabel pdiffusion 213 -24 213 -24 0 cellNo=3
rlabel pdiffusion 255 -24 255 -24 0 feedthrough
rlabel pdiffusion 353 -24 353 -24 0 feedthrough
rlabel pdiffusion 395 -24 395 -24 0 cellNo=581
rlabel pdiffusion 416 -24 416 -24 0 cellNo=568
rlabel pdiffusion 423 -24 423 -24 0 feedthrough
rlabel pdiffusion 430 -24 430 -24 0 cellNo=352
rlabel pdiffusion 444 -24 444 -24 0 cellNo=15
rlabel pdiffusion 486 -24 486 -24 0 feedthrough
rlabel pdiffusion 549 -24 549 -24 0 feedthrough
rlabel pdiffusion 556 -24 556 -24 0 cellNo=128
rlabel pdiffusion 570 -24 570 -24 0 cellNo=671
rlabel pdiffusion 577 -24 577 -24 0 feedthrough
rlabel pdiffusion 584 -24 584 -24 0 feedthrough
rlabel pdiffusion 605 -24 605 -24 0 feedthrough
rlabel pdiffusion 612 -24 612 -24 0 cellNo=9
rlabel pdiffusion 619 -24 619 -24 0 feedthrough
rlabel pdiffusion 626 -24 626 -24 0 feedthrough
rlabel pdiffusion 633 -24 633 -24 0 cellNo=67
rlabel pdiffusion 640 -24 640 -24 0 feedthrough
rlabel pdiffusion 647 -24 647 -24 0 feedthrough
rlabel pdiffusion 654 -24 654 -24 0 cellNo=612
rlabel pdiffusion 661 -24 661 -24 0 cellNo=441
rlabel pdiffusion 682 -24 682 -24 0 cellNo=758
rlabel pdiffusion 689 -24 689 -24 0 feedthrough
rlabel pdiffusion 703 -24 703 -24 0 cellNo=170
rlabel pdiffusion 710 -24 710 -24 0 feedthrough
rlabel pdiffusion 717 -24 717 -24 0 feedthrough
rlabel pdiffusion 731 -24 731 -24 0 feedthrough
rlabel pdiffusion 766 -24 766 -24 0 cellNo=405
rlabel pdiffusion 773 -24 773 -24 0 feedthrough
rlabel pdiffusion 794 -24 794 -24 0 cellNo=965
rlabel pdiffusion 801 -24 801 -24 0 cellNo=497
rlabel pdiffusion 808 -24 808 -24 0 cellNo=575
rlabel pdiffusion 815 -24 815 -24 0 feedthrough
rlabel pdiffusion 822 -24 822 -24 0 cellNo=690
rlabel pdiffusion 829 -24 829 -24 0 feedthrough
rlabel pdiffusion 836 -24 836 -24 0 feedthrough
rlabel pdiffusion 843 -24 843 -24 0 cellNo=950
rlabel pdiffusion 850 -24 850 -24 0 cellNo=646
rlabel pdiffusion 857 -24 857 -24 0 cellNo=216
rlabel pdiffusion 864 -24 864 -24 0 cellNo=371
rlabel pdiffusion 871 -24 871 -24 0 feedthrough
rlabel pdiffusion 885 -24 885 -24 0 cellNo=635
rlabel pdiffusion 892 -24 892 -24 0 feedthrough
rlabel pdiffusion 899 -24 899 -24 0 cellNo=125
rlabel pdiffusion 913 -24 913 -24 0 cellNo=347
rlabel pdiffusion 920 -24 920 -24 0 feedthrough
rlabel pdiffusion 962 -24 962 -24 0 feedthrough
rlabel pdiffusion 969 -24 969 -24 0 cellNo=604
rlabel pdiffusion 976 -24 976 -24 0 cellNo=169
rlabel pdiffusion 983 -24 983 -24 0 feedthrough
rlabel pdiffusion 990 -24 990 -24 0 feedthrough
rlabel pdiffusion 1039 -24 1039 -24 0 feedthrough
rlabel pdiffusion 1074 -24 1074 -24 0 feedthrough
rlabel pdiffusion 1088 -24 1088 -24 0 feedthrough
rlabel pdiffusion 1095 -24 1095 -24 0 feedthrough
rlabel pdiffusion 1123 -24 1123 -24 0 cellNo=28
rlabel pdiffusion 1130 -24 1130 -24 0 cellNo=175
rlabel pdiffusion 1207 -24 1207 -24 0 feedthrough
rlabel pdiffusion 1438 -24 1438 -24 0 cellNo=661
rlabel pdiffusion 1627 -24 1627 -24 0 cellNo=5
rlabel pdiffusion 3 -71 3 -71 0 cellNo=485
rlabel pdiffusion 10 -71 10 -71 0 cellNo=1184
rlabel pdiffusion 17 -71 17 -71 0 cellNo=1012
rlabel pdiffusion 24 -71 24 -71 0 cellNo=688
rlabel pdiffusion 31 -71 31 -71 0 cellNo=1026
rlabel pdiffusion 38 -71 38 -71 0 cellNo=1010
rlabel pdiffusion 45 -71 45 -71 0 cellNo=1045
rlabel pdiffusion 52 -71 52 -71 0 cellNo=1077
rlabel pdiffusion 59 -71 59 -71 0 cellNo=1209
rlabel pdiffusion 185 -71 185 -71 0 feedthrough
rlabel pdiffusion 199 -71 199 -71 0 feedthrough
rlabel pdiffusion 241 -71 241 -71 0 feedthrough
rlabel pdiffusion 276 -71 276 -71 0 feedthrough
rlabel pdiffusion 297 -71 297 -71 0 feedthrough
rlabel pdiffusion 311 -71 311 -71 0 cellNo=404
rlabel pdiffusion 318 -71 318 -71 0 feedthrough
rlabel pdiffusion 353 -71 353 -71 0 cellNo=36
rlabel pdiffusion 395 -71 395 -71 0 feedthrough
rlabel pdiffusion 402 -71 402 -71 0 cellNo=735
rlabel pdiffusion 409 -71 409 -71 0 cellNo=732
rlabel pdiffusion 416 -71 416 -71 0 feedthrough
rlabel pdiffusion 423 -71 423 -71 0 feedthrough
rlabel pdiffusion 465 -71 465 -71 0 feedthrough
rlabel pdiffusion 472 -71 472 -71 0 feedthrough
rlabel pdiffusion 479 -71 479 -71 0 feedthrough
rlabel pdiffusion 486 -71 486 -71 0 feedthrough
rlabel pdiffusion 493 -71 493 -71 0 feedthrough
rlabel pdiffusion 500 -71 500 -71 0 feedthrough
rlabel pdiffusion 507 -71 507 -71 0 feedthrough
rlabel pdiffusion 521 -71 521 -71 0 feedthrough
rlabel pdiffusion 535 -71 535 -71 0 feedthrough
rlabel pdiffusion 542 -71 542 -71 0 cellNo=823
rlabel pdiffusion 549 -71 549 -71 0 feedthrough
rlabel pdiffusion 563 -71 563 -71 0 cellNo=387
rlabel pdiffusion 570 -71 570 -71 0 feedthrough
rlabel pdiffusion 584 -71 584 -71 0 cellNo=291
rlabel pdiffusion 591 -71 591 -71 0 feedthrough
rlabel pdiffusion 598 -71 598 -71 0 feedthrough
rlabel pdiffusion 605 -71 605 -71 0 feedthrough
rlabel pdiffusion 612 -71 612 -71 0 feedthrough
rlabel pdiffusion 619 -71 619 -71 0 feedthrough
rlabel pdiffusion 640 -71 640 -71 0 feedthrough
rlabel pdiffusion 647 -71 647 -71 0 feedthrough
rlabel pdiffusion 654 -71 654 -71 0 cellNo=911
rlabel pdiffusion 661 -71 661 -71 0 feedthrough
rlabel pdiffusion 668 -71 668 -71 0 feedthrough
rlabel pdiffusion 675 -71 675 -71 0 cellNo=864
rlabel pdiffusion 682 -71 682 -71 0 feedthrough
rlabel pdiffusion 689 -71 689 -71 0 feedthrough
rlabel pdiffusion 696 -71 696 -71 0 cellNo=854
rlabel pdiffusion 703 -71 703 -71 0 feedthrough
rlabel pdiffusion 710 -71 710 -71 0 feedthrough
rlabel pdiffusion 717 -71 717 -71 0 feedthrough
rlabel pdiffusion 724 -71 724 -71 0 feedthrough
rlabel pdiffusion 731 -71 731 -71 0 feedthrough
rlabel pdiffusion 738 -71 738 -71 0 cellNo=148
rlabel pdiffusion 745 -71 745 -71 0 feedthrough
rlabel pdiffusion 752 -71 752 -71 0 feedthrough
rlabel pdiffusion 759 -71 759 -71 0 feedthrough
rlabel pdiffusion 766 -71 766 -71 0 feedthrough
rlabel pdiffusion 773 -71 773 -71 0 feedthrough
rlabel pdiffusion 780 -71 780 -71 0 feedthrough
rlabel pdiffusion 787 -71 787 -71 0 cellNo=237
rlabel pdiffusion 794 -71 794 -71 0 feedthrough
rlabel pdiffusion 801 -71 801 -71 0 cellNo=608
rlabel pdiffusion 808 -71 808 -71 0 feedthrough
rlabel pdiffusion 815 -71 815 -71 0 feedthrough
rlabel pdiffusion 822 -71 822 -71 0 feedthrough
rlabel pdiffusion 829 -71 829 -71 0 feedthrough
rlabel pdiffusion 836 -71 836 -71 0 feedthrough
rlabel pdiffusion 843 -71 843 -71 0 feedthrough
rlabel pdiffusion 850 -71 850 -71 0 cellNo=514
rlabel pdiffusion 857 -71 857 -71 0 cellNo=991
rlabel pdiffusion 864 -71 864 -71 0 feedthrough
rlabel pdiffusion 871 -71 871 -71 0 feedthrough
rlabel pdiffusion 878 -71 878 -71 0 feedthrough
rlabel pdiffusion 885 -71 885 -71 0 cellNo=793
rlabel pdiffusion 892 -71 892 -71 0 feedthrough
rlabel pdiffusion 899 -71 899 -71 0 cellNo=317
rlabel pdiffusion 906 -71 906 -71 0 cellNo=102
rlabel pdiffusion 913 -71 913 -71 0 feedthrough
rlabel pdiffusion 920 -71 920 -71 0 feedthrough
rlabel pdiffusion 927 -71 927 -71 0 feedthrough
rlabel pdiffusion 934 -71 934 -71 0 feedthrough
rlabel pdiffusion 941 -71 941 -71 0 cellNo=233
rlabel pdiffusion 948 -71 948 -71 0 feedthrough
rlabel pdiffusion 955 -71 955 -71 0 cellNo=902
rlabel pdiffusion 962 -71 962 -71 0 feedthrough
rlabel pdiffusion 969 -71 969 -71 0 feedthrough
rlabel pdiffusion 976 -71 976 -71 0 feedthrough
rlabel pdiffusion 983 -71 983 -71 0 feedthrough
rlabel pdiffusion 990 -71 990 -71 0 feedthrough
rlabel pdiffusion 997 -71 997 -71 0 cellNo=746
rlabel pdiffusion 1004 -71 1004 -71 0 feedthrough
rlabel pdiffusion 1011 -71 1011 -71 0 feedthrough
rlabel pdiffusion 1018 -71 1018 -71 0 feedthrough
rlabel pdiffusion 1025 -71 1025 -71 0 cellNo=770
rlabel pdiffusion 1032 -71 1032 -71 0 feedthrough
rlabel pdiffusion 1039 -71 1039 -71 0 feedthrough
rlabel pdiffusion 1046 -71 1046 -71 0 feedthrough
rlabel pdiffusion 1053 -71 1053 -71 0 feedthrough
rlabel pdiffusion 1060 -71 1060 -71 0 feedthrough
rlabel pdiffusion 1067 -71 1067 -71 0 cellNo=76
rlabel pdiffusion 1074 -71 1074 -71 0 feedthrough
rlabel pdiffusion 1081 -71 1081 -71 0 feedthrough
rlabel pdiffusion 1088 -71 1088 -71 0 feedthrough
rlabel pdiffusion 1095 -71 1095 -71 0 feedthrough
rlabel pdiffusion 1102 -71 1102 -71 0 feedthrough
rlabel pdiffusion 1109 -71 1109 -71 0 cellNo=663
rlabel pdiffusion 1116 -71 1116 -71 0 cellNo=51
rlabel pdiffusion 1123 -71 1123 -71 0 cellNo=195
rlabel pdiffusion 1151 -71 1151 -71 0 feedthrough
rlabel pdiffusion 1165 -71 1165 -71 0 cellNo=449
rlabel pdiffusion 1179 -71 1179 -71 0 feedthrough
rlabel pdiffusion 1214 -71 1214 -71 0 feedthrough
rlabel pdiffusion 1221 -71 1221 -71 0 feedthrough
rlabel pdiffusion 1228 -71 1228 -71 0 cellNo=926
rlabel pdiffusion 1235 -71 1235 -71 0 cellNo=453
rlabel pdiffusion 1291 -71 1291 -71 0 feedthrough
rlabel pdiffusion 1319 -71 1319 -71 0 cellNo=309
rlabel pdiffusion 1333 -71 1333 -71 0 feedthrough
rlabel pdiffusion 1361 -71 1361 -71 0 feedthrough
rlabel pdiffusion 1487 -71 1487 -71 0 feedthrough
rlabel pdiffusion 1634 -71 1634 -71 0 feedthrough
rlabel pdiffusion 1760 -71 1760 -71 0 feedthrough
rlabel pdiffusion 3 -148 3 -148 0 cellNo=1001
rlabel pdiffusion 10 -148 10 -148 0 cellNo=1037
rlabel pdiffusion 59 -148 59 -148 0 feedthrough
rlabel pdiffusion 66 -148 66 -148 0 feedthrough
rlabel pdiffusion 73 -148 73 -148 0 feedthrough
rlabel pdiffusion 80 -148 80 -148 0 feedthrough
rlabel pdiffusion 87 -148 87 -148 0 feedthrough
rlabel pdiffusion 94 -148 94 -148 0 feedthrough
rlabel pdiffusion 101 -148 101 -148 0 feedthrough
rlabel pdiffusion 108 -148 108 -148 0 feedthrough
rlabel pdiffusion 115 -148 115 -148 0 feedthrough
rlabel pdiffusion 122 -148 122 -148 0 cellNo=64
rlabel pdiffusion 129 -148 129 -148 0 feedthrough
rlabel pdiffusion 136 -148 136 -148 0 feedthrough
rlabel pdiffusion 143 -148 143 -148 0 cellNo=323
rlabel pdiffusion 150 -148 150 -148 0 cellNo=632
rlabel pdiffusion 157 -148 157 -148 0 feedthrough
rlabel pdiffusion 164 -148 164 -148 0 feedthrough
rlabel pdiffusion 171 -148 171 -148 0 feedthrough
rlabel pdiffusion 178 -148 178 -148 0 feedthrough
rlabel pdiffusion 185 -148 185 -148 0 feedthrough
rlabel pdiffusion 192 -148 192 -148 0 feedthrough
rlabel pdiffusion 199 -148 199 -148 0 feedthrough
rlabel pdiffusion 206 -148 206 -148 0 feedthrough
rlabel pdiffusion 213 -148 213 -148 0 feedthrough
rlabel pdiffusion 220 -148 220 -148 0 feedthrough
rlabel pdiffusion 227 -148 227 -148 0 cellNo=666
rlabel pdiffusion 234 -148 234 -148 0 cellNo=200
rlabel pdiffusion 241 -148 241 -148 0 feedthrough
rlabel pdiffusion 248 -148 248 -148 0 feedthrough
rlabel pdiffusion 255 -148 255 -148 0 cellNo=205
rlabel pdiffusion 262 -148 262 -148 0 cellNo=81
rlabel pdiffusion 269 -148 269 -148 0 cellNo=775
rlabel pdiffusion 276 -148 276 -148 0 feedthrough
rlabel pdiffusion 283 -148 283 -148 0 feedthrough
rlabel pdiffusion 290 -148 290 -148 0 feedthrough
rlabel pdiffusion 297 -148 297 -148 0 feedthrough
rlabel pdiffusion 304 -148 304 -148 0 feedthrough
rlabel pdiffusion 311 -148 311 -148 0 feedthrough
rlabel pdiffusion 318 -148 318 -148 0 feedthrough
rlabel pdiffusion 325 -148 325 -148 0 feedthrough
rlabel pdiffusion 332 -148 332 -148 0 feedthrough
rlabel pdiffusion 339 -148 339 -148 0 feedthrough
rlabel pdiffusion 346 -148 346 -148 0 feedthrough
rlabel pdiffusion 353 -148 353 -148 0 feedthrough
rlabel pdiffusion 360 -148 360 -148 0 feedthrough
rlabel pdiffusion 367 -148 367 -148 0 feedthrough
rlabel pdiffusion 374 -148 374 -148 0 feedthrough
rlabel pdiffusion 381 -148 381 -148 0 feedthrough
rlabel pdiffusion 388 -148 388 -148 0 cellNo=724
rlabel pdiffusion 395 -148 395 -148 0 feedthrough
rlabel pdiffusion 402 -148 402 -148 0 feedthrough
rlabel pdiffusion 409 -148 409 -148 0 feedthrough
rlabel pdiffusion 416 -148 416 -148 0 feedthrough
rlabel pdiffusion 423 -148 423 -148 0 feedthrough
rlabel pdiffusion 430 -148 430 -148 0 feedthrough
rlabel pdiffusion 437 -148 437 -148 0 feedthrough
rlabel pdiffusion 444 -148 444 -148 0 cellNo=694
rlabel pdiffusion 451 -148 451 -148 0 feedthrough
rlabel pdiffusion 458 -148 458 -148 0 cellNo=711
rlabel pdiffusion 465 -148 465 -148 0 cellNo=253
rlabel pdiffusion 472 -148 472 -148 0 cellNo=801
rlabel pdiffusion 479 -148 479 -148 0 feedthrough
rlabel pdiffusion 486 -148 486 -148 0 feedthrough
rlabel pdiffusion 493 -148 493 -148 0 feedthrough
rlabel pdiffusion 500 -148 500 -148 0 feedthrough
rlabel pdiffusion 507 -148 507 -148 0 feedthrough
rlabel pdiffusion 514 -148 514 -148 0 feedthrough
rlabel pdiffusion 521 -148 521 -148 0 cellNo=966
rlabel pdiffusion 528 -148 528 -148 0 cellNo=86
rlabel pdiffusion 535 -148 535 -148 0 feedthrough
rlabel pdiffusion 542 -148 542 -148 0 feedthrough
rlabel pdiffusion 549 -148 549 -148 0 feedthrough
rlabel pdiffusion 556 -148 556 -148 0 feedthrough
rlabel pdiffusion 563 -148 563 -148 0 cellNo=783
rlabel pdiffusion 570 -148 570 -148 0 feedthrough
rlabel pdiffusion 577 -148 577 -148 0 feedthrough
rlabel pdiffusion 584 -148 584 -148 0 feedthrough
rlabel pdiffusion 591 -148 591 -148 0 feedthrough
rlabel pdiffusion 598 -148 598 -148 0 cellNo=208
rlabel pdiffusion 605 -148 605 -148 0 feedthrough
rlabel pdiffusion 612 -148 612 -148 0 feedthrough
rlabel pdiffusion 619 -148 619 -148 0 feedthrough
rlabel pdiffusion 626 -148 626 -148 0 feedthrough
rlabel pdiffusion 633 -148 633 -148 0 feedthrough
rlabel pdiffusion 640 -148 640 -148 0 feedthrough
rlabel pdiffusion 647 -148 647 -148 0 cellNo=993
rlabel pdiffusion 654 -148 654 -148 0 feedthrough
rlabel pdiffusion 661 -148 661 -148 0 feedthrough
rlabel pdiffusion 668 -148 668 -148 0 feedthrough
rlabel pdiffusion 675 -148 675 -148 0 cellNo=160
rlabel pdiffusion 682 -148 682 -148 0 cellNo=284
rlabel pdiffusion 689 -148 689 -148 0 feedthrough
rlabel pdiffusion 696 -148 696 -148 0 cellNo=312
rlabel pdiffusion 703 -148 703 -148 0 feedthrough
rlabel pdiffusion 710 -148 710 -148 0 feedthrough
rlabel pdiffusion 717 -148 717 -148 0 feedthrough
rlabel pdiffusion 724 -148 724 -148 0 feedthrough
rlabel pdiffusion 731 -148 731 -148 0 cellNo=795
rlabel pdiffusion 738 -148 738 -148 0 cellNo=268
rlabel pdiffusion 745 -148 745 -148 0 feedthrough
rlabel pdiffusion 752 -148 752 -148 0 feedthrough
rlabel pdiffusion 759 -148 759 -148 0 feedthrough
rlabel pdiffusion 766 -148 766 -148 0 cellNo=365
rlabel pdiffusion 773 -148 773 -148 0 cellNo=706
rlabel pdiffusion 780 -148 780 -148 0 feedthrough
rlabel pdiffusion 787 -148 787 -148 0 feedthrough
rlabel pdiffusion 794 -148 794 -148 0 feedthrough
rlabel pdiffusion 801 -148 801 -148 0 cellNo=640
rlabel pdiffusion 808 -148 808 -148 0 feedthrough
rlabel pdiffusion 815 -148 815 -148 0 feedthrough
rlabel pdiffusion 822 -148 822 -148 0 feedthrough
rlabel pdiffusion 829 -148 829 -148 0 feedthrough
rlabel pdiffusion 836 -148 836 -148 0 cellNo=553
rlabel pdiffusion 843 -148 843 -148 0 feedthrough
rlabel pdiffusion 850 -148 850 -148 0 feedthrough
rlabel pdiffusion 857 -148 857 -148 0 feedthrough
rlabel pdiffusion 864 -148 864 -148 0 feedthrough
rlabel pdiffusion 871 -148 871 -148 0 feedthrough
rlabel pdiffusion 878 -148 878 -148 0 feedthrough
rlabel pdiffusion 885 -148 885 -148 0 feedthrough
rlabel pdiffusion 892 -148 892 -148 0 feedthrough
rlabel pdiffusion 899 -148 899 -148 0 feedthrough
rlabel pdiffusion 906 -148 906 -148 0 feedthrough
rlabel pdiffusion 913 -148 913 -148 0 feedthrough
rlabel pdiffusion 920 -148 920 -148 0 feedthrough
rlabel pdiffusion 927 -148 927 -148 0 cellNo=948
rlabel pdiffusion 934 -148 934 -148 0 cellNo=474
rlabel pdiffusion 941 -148 941 -148 0 feedthrough
rlabel pdiffusion 948 -148 948 -148 0 cellNo=620
rlabel pdiffusion 955 -148 955 -148 0 feedthrough
rlabel pdiffusion 962 -148 962 -148 0 cellNo=678
rlabel pdiffusion 969 -148 969 -148 0 feedthrough
rlabel pdiffusion 976 -148 976 -148 0 cellNo=369
rlabel pdiffusion 983 -148 983 -148 0 feedthrough
rlabel pdiffusion 990 -148 990 -148 0 feedthrough
rlabel pdiffusion 997 -148 997 -148 0 feedthrough
rlabel pdiffusion 1004 -148 1004 -148 0 feedthrough
rlabel pdiffusion 1011 -148 1011 -148 0 feedthrough
rlabel pdiffusion 1018 -148 1018 -148 0 feedthrough
rlabel pdiffusion 1025 -148 1025 -148 0 feedthrough
rlabel pdiffusion 1032 -148 1032 -148 0 feedthrough
rlabel pdiffusion 1039 -148 1039 -148 0 feedthrough
rlabel pdiffusion 1046 -148 1046 -148 0 feedthrough
rlabel pdiffusion 1053 -148 1053 -148 0 feedthrough
rlabel pdiffusion 1060 -148 1060 -148 0 feedthrough
rlabel pdiffusion 1067 -148 1067 -148 0 feedthrough
rlabel pdiffusion 1074 -148 1074 -148 0 cellNo=885
rlabel pdiffusion 1081 -148 1081 -148 0 feedthrough
rlabel pdiffusion 1088 -148 1088 -148 0 cellNo=591
rlabel pdiffusion 1095 -148 1095 -148 0 feedthrough
rlabel pdiffusion 1102 -148 1102 -148 0 feedthrough
rlabel pdiffusion 1109 -148 1109 -148 0 feedthrough
rlabel pdiffusion 1116 -148 1116 -148 0 feedthrough
rlabel pdiffusion 1123 -148 1123 -148 0 feedthrough
rlabel pdiffusion 1130 -148 1130 -148 0 feedthrough
rlabel pdiffusion 1137 -148 1137 -148 0 feedthrough
rlabel pdiffusion 1144 -148 1144 -148 0 cellNo=631
rlabel pdiffusion 1151 -148 1151 -148 0 feedthrough
rlabel pdiffusion 1158 -148 1158 -148 0 feedthrough
rlabel pdiffusion 1165 -148 1165 -148 0 feedthrough
rlabel pdiffusion 1172 -148 1172 -148 0 cellNo=493
rlabel pdiffusion 1179 -148 1179 -148 0 feedthrough
rlabel pdiffusion 1186 -148 1186 -148 0 feedthrough
rlabel pdiffusion 1193 -148 1193 -148 0 feedthrough
rlabel pdiffusion 1200 -148 1200 -148 0 feedthrough
rlabel pdiffusion 1207 -148 1207 -148 0 feedthrough
rlabel pdiffusion 1214 -148 1214 -148 0 feedthrough
rlabel pdiffusion 1221 -148 1221 -148 0 feedthrough
rlabel pdiffusion 1228 -148 1228 -148 0 feedthrough
rlabel pdiffusion 1235 -148 1235 -148 0 feedthrough
rlabel pdiffusion 1242 -148 1242 -148 0 feedthrough
rlabel pdiffusion 1249 -148 1249 -148 0 feedthrough
rlabel pdiffusion 1256 -148 1256 -148 0 feedthrough
rlabel pdiffusion 1263 -148 1263 -148 0 cellNo=97
rlabel pdiffusion 1270 -148 1270 -148 0 feedthrough
rlabel pdiffusion 1277 -148 1277 -148 0 feedthrough
rlabel pdiffusion 1284 -148 1284 -148 0 feedthrough
rlabel pdiffusion 1291 -148 1291 -148 0 feedthrough
rlabel pdiffusion 1298 -148 1298 -148 0 feedthrough
rlabel pdiffusion 1305 -148 1305 -148 0 feedthrough
rlabel pdiffusion 1312 -148 1312 -148 0 feedthrough
rlabel pdiffusion 1319 -148 1319 -148 0 feedthrough
rlabel pdiffusion 1326 -148 1326 -148 0 feedthrough
rlabel pdiffusion 1354 -148 1354 -148 0 feedthrough
rlabel pdiffusion 1361 -148 1361 -148 0 feedthrough
rlabel pdiffusion 1375 -148 1375 -148 0 feedthrough
rlabel pdiffusion 1424 -148 1424 -148 0 feedthrough
rlabel pdiffusion 1508 -148 1508 -148 0 feedthrough
rlabel pdiffusion 1515 -148 1515 -148 0 feedthrough
rlabel pdiffusion 1641 -148 1641 -148 0 feedthrough
rlabel pdiffusion 1886 -148 1886 -148 0 feedthrough
rlabel pdiffusion 3 -251 3 -251 0 cellNo=1011
rlabel pdiffusion 10 -251 10 -251 0 cellNo=1150
rlabel pdiffusion 17 -251 17 -251 0 feedthrough
rlabel pdiffusion 24 -251 24 -251 0 feedthrough
rlabel pdiffusion 31 -251 31 -251 0 feedthrough
rlabel pdiffusion 38 -251 38 -251 0 feedthrough
rlabel pdiffusion 45 -251 45 -251 0 feedthrough
rlabel pdiffusion 52 -251 52 -251 0 feedthrough
rlabel pdiffusion 59 -251 59 -251 0 feedthrough
rlabel pdiffusion 66 -251 66 -251 0 cellNo=1052
rlabel pdiffusion 73 -251 73 -251 0 feedthrough
rlabel pdiffusion 80 -251 80 -251 0 cellNo=856
rlabel pdiffusion 87 -251 87 -251 0 cellNo=183
rlabel pdiffusion 94 -251 94 -251 0 feedthrough
rlabel pdiffusion 101 -251 101 -251 0 feedthrough
rlabel pdiffusion 108 -251 108 -251 0 feedthrough
rlabel pdiffusion 115 -251 115 -251 0 cellNo=84
rlabel pdiffusion 122 -251 122 -251 0 feedthrough
rlabel pdiffusion 129 -251 129 -251 0 feedthrough
rlabel pdiffusion 136 -251 136 -251 0 cellNo=482
rlabel pdiffusion 143 -251 143 -251 0 feedthrough
rlabel pdiffusion 150 -251 150 -251 0 feedthrough
rlabel pdiffusion 157 -251 157 -251 0 cellNo=636
rlabel pdiffusion 164 -251 164 -251 0 feedthrough
rlabel pdiffusion 171 -251 171 -251 0 feedthrough
rlabel pdiffusion 178 -251 178 -251 0 feedthrough
rlabel pdiffusion 185 -251 185 -251 0 feedthrough
rlabel pdiffusion 192 -251 192 -251 0 cellNo=386
rlabel pdiffusion 199 -251 199 -251 0 cellNo=820
rlabel pdiffusion 206 -251 206 -251 0 cellNo=144
rlabel pdiffusion 213 -251 213 -251 0 cellNo=651
rlabel pdiffusion 220 -251 220 -251 0 feedthrough
rlabel pdiffusion 227 -251 227 -251 0 feedthrough
rlabel pdiffusion 234 -251 234 -251 0 feedthrough
rlabel pdiffusion 241 -251 241 -251 0 cellNo=590
rlabel pdiffusion 248 -251 248 -251 0 feedthrough
rlabel pdiffusion 255 -251 255 -251 0 feedthrough
rlabel pdiffusion 262 -251 262 -251 0 feedthrough
rlabel pdiffusion 269 -251 269 -251 0 cellNo=714
rlabel pdiffusion 276 -251 276 -251 0 feedthrough
rlabel pdiffusion 283 -251 283 -251 0 feedthrough
rlabel pdiffusion 290 -251 290 -251 0 feedthrough
rlabel pdiffusion 297 -251 297 -251 0 cellNo=357
rlabel pdiffusion 304 -251 304 -251 0 feedthrough
rlabel pdiffusion 311 -251 311 -251 0 cellNo=251
rlabel pdiffusion 318 -251 318 -251 0 feedthrough
rlabel pdiffusion 325 -251 325 -251 0 feedthrough
rlabel pdiffusion 332 -251 332 -251 0 feedthrough
rlabel pdiffusion 339 -251 339 -251 0 feedthrough
rlabel pdiffusion 346 -251 346 -251 0 feedthrough
rlabel pdiffusion 353 -251 353 -251 0 feedthrough
rlabel pdiffusion 360 -251 360 -251 0 feedthrough
rlabel pdiffusion 367 -251 367 -251 0 feedthrough
rlabel pdiffusion 374 -251 374 -251 0 feedthrough
rlabel pdiffusion 381 -251 381 -251 0 feedthrough
rlabel pdiffusion 388 -251 388 -251 0 feedthrough
rlabel pdiffusion 395 -251 395 -251 0 feedthrough
rlabel pdiffusion 402 -251 402 -251 0 feedthrough
rlabel pdiffusion 409 -251 409 -251 0 feedthrough
rlabel pdiffusion 416 -251 416 -251 0 feedthrough
rlabel pdiffusion 423 -251 423 -251 0 feedthrough
rlabel pdiffusion 430 -251 430 -251 0 feedthrough
rlabel pdiffusion 437 -251 437 -251 0 cellNo=425
rlabel pdiffusion 444 -251 444 -251 0 feedthrough
rlabel pdiffusion 451 -251 451 -251 0 feedthrough
rlabel pdiffusion 458 -251 458 -251 0 feedthrough
rlabel pdiffusion 465 -251 465 -251 0 cellNo=615
rlabel pdiffusion 472 -251 472 -251 0 feedthrough
rlabel pdiffusion 479 -251 479 -251 0 feedthrough
rlabel pdiffusion 486 -251 486 -251 0 feedthrough
rlabel pdiffusion 493 -251 493 -251 0 feedthrough
rlabel pdiffusion 500 -251 500 -251 0 feedthrough
rlabel pdiffusion 507 -251 507 -251 0 feedthrough
rlabel pdiffusion 514 -251 514 -251 0 feedthrough
rlabel pdiffusion 521 -251 521 -251 0 cellNo=643
rlabel pdiffusion 528 -251 528 -251 0 feedthrough
rlabel pdiffusion 535 -251 535 -251 0 cellNo=884
rlabel pdiffusion 542 -251 542 -251 0 feedthrough
rlabel pdiffusion 549 -251 549 -251 0 feedthrough
rlabel pdiffusion 556 -251 556 -251 0 feedthrough
rlabel pdiffusion 563 -251 563 -251 0 feedthrough
rlabel pdiffusion 570 -251 570 -251 0 feedthrough
rlabel pdiffusion 577 -251 577 -251 0 feedthrough
rlabel pdiffusion 584 -251 584 -251 0 feedthrough
rlabel pdiffusion 591 -251 591 -251 0 cellNo=478
rlabel pdiffusion 598 -251 598 -251 0 feedthrough
rlabel pdiffusion 605 -251 605 -251 0 feedthrough
rlabel pdiffusion 612 -251 612 -251 0 feedthrough
rlabel pdiffusion 619 -251 619 -251 0 cellNo=778
rlabel pdiffusion 626 -251 626 -251 0 feedthrough
rlabel pdiffusion 633 -251 633 -251 0 feedthrough
rlabel pdiffusion 640 -251 640 -251 0 feedthrough
rlabel pdiffusion 647 -251 647 -251 0 feedthrough
rlabel pdiffusion 654 -251 654 -251 0 feedthrough
rlabel pdiffusion 661 -251 661 -251 0 feedthrough
rlabel pdiffusion 668 -251 668 -251 0 feedthrough
rlabel pdiffusion 675 -251 675 -251 0 feedthrough
rlabel pdiffusion 682 -251 682 -251 0 feedthrough
rlabel pdiffusion 689 -251 689 -251 0 feedthrough
rlabel pdiffusion 696 -251 696 -251 0 feedthrough
rlabel pdiffusion 703 -251 703 -251 0 cellNo=120
rlabel pdiffusion 710 -251 710 -251 0 cellNo=342
rlabel pdiffusion 717 -251 717 -251 0 feedthrough
rlabel pdiffusion 724 -251 724 -251 0 feedthrough
rlabel pdiffusion 731 -251 731 -251 0 feedthrough
rlabel pdiffusion 738 -251 738 -251 0 feedthrough
rlabel pdiffusion 745 -251 745 -251 0 feedthrough
rlabel pdiffusion 752 -251 752 -251 0 feedthrough
rlabel pdiffusion 759 -251 759 -251 0 feedthrough
rlabel pdiffusion 766 -251 766 -251 0 feedthrough
rlabel pdiffusion 773 -251 773 -251 0 feedthrough
rlabel pdiffusion 780 -251 780 -251 0 feedthrough
rlabel pdiffusion 787 -251 787 -251 0 feedthrough
rlabel pdiffusion 794 -251 794 -251 0 feedthrough
rlabel pdiffusion 801 -251 801 -251 0 feedthrough
rlabel pdiffusion 808 -251 808 -251 0 feedthrough
rlabel pdiffusion 815 -251 815 -251 0 feedthrough
rlabel pdiffusion 822 -251 822 -251 0 feedthrough
rlabel pdiffusion 829 -251 829 -251 0 feedthrough
rlabel pdiffusion 836 -251 836 -251 0 feedthrough
rlabel pdiffusion 843 -251 843 -251 0 feedthrough
rlabel pdiffusion 850 -251 850 -251 0 feedthrough
rlabel pdiffusion 857 -251 857 -251 0 feedthrough
rlabel pdiffusion 864 -251 864 -251 0 feedthrough
rlabel pdiffusion 871 -251 871 -251 0 feedthrough
rlabel pdiffusion 878 -251 878 -251 0 feedthrough
rlabel pdiffusion 885 -251 885 -251 0 cellNo=766
rlabel pdiffusion 892 -251 892 -251 0 cellNo=281
rlabel pdiffusion 899 -251 899 -251 0 feedthrough
rlabel pdiffusion 906 -251 906 -251 0 feedthrough
rlabel pdiffusion 913 -251 913 -251 0 cellNo=218
rlabel pdiffusion 920 -251 920 -251 0 feedthrough
rlabel pdiffusion 927 -251 927 -251 0 feedthrough
rlabel pdiffusion 934 -251 934 -251 0 feedthrough
rlabel pdiffusion 941 -251 941 -251 0 feedthrough
rlabel pdiffusion 948 -251 948 -251 0 feedthrough
rlabel pdiffusion 955 -251 955 -251 0 feedthrough
rlabel pdiffusion 962 -251 962 -251 0 feedthrough
rlabel pdiffusion 969 -251 969 -251 0 feedthrough
rlabel pdiffusion 976 -251 976 -251 0 feedthrough
rlabel pdiffusion 983 -251 983 -251 0 feedthrough
rlabel pdiffusion 990 -251 990 -251 0 cellNo=112
rlabel pdiffusion 997 -251 997 -251 0 cellNo=492
rlabel pdiffusion 1004 -251 1004 -251 0 feedthrough
rlabel pdiffusion 1011 -251 1011 -251 0 cellNo=521
rlabel pdiffusion 1018 -251 1018 -251 0 feedthrough
rlabel pdiffusion 1025 -251 1025 -251 0 feedthrough
rlabel pdiffusion 1032 -251 1032 -251 0 feedthrough
rlabel pdiffusion 1039 -251 1039 -251 0 feedthrough
rlabel pdiffusion 1046 -251 1046 -251 0 feedthrough
rlabel pdiffusion 1053 -251 1053 -251 0 feedthrough
rlabel pdiffusion 1060 -251 1060 -251 0 feedthrough
rlabel pdiffusion 1067 -251 1067 -251 0 feedthrough
rlabel pdiffusion 1074 -251 1074 -251 0 feedthrough
rlabel pdiffusion 1081 -251 1081 -251 0 feedthrough
rlabel pdiffusion 1088 -251 1088 -251 0 feedthrough
rlabel pdiffusion 1095 -251 1095 -251 0 feedthrough
rlabel pdiffusion 1102 -251 1102 -251 0 feedthrough
rlabel pdiffusion 1109 -251 1109 -251 0 feedthrough
rlabel pdiffusion 1116 -251 1116 -251 0 feedthrough
rlabel pdiffusion 1123 -251 1123 -251 0 feedthrough
rlabel pdiffusion 1130 -251 1130 -251 0 feedthrough
rlabel pdiffusion 1137 -251 1137 -251 0 feedthrough
rlabel pdiffusion 1144 -251 1144 -251 0 feedthrough
rlabel pdiffusion 1151 -251 1151 -251 0 cellNo=602
rlabel pdiffusion 1158 -251 1158 -251 0 feedthrough
rlabel pdiffusion 1165 -251 1165 -251 0 feedthrough
rlabel pdiffusion 1172 -251 1172 -251 0 feedthrough
rlabel pdiffusion 1179 -251 1179 -251 0 cellNo=38
rlabel pdiffusion 1186 -251 1186 -251 0 feedthrough
rlabel pdiffusion 1193 -251 1193 -251 0 feedthrough
rlabel pdiffusion 1200 -251 1200 -251 0 cellNo=587
rlabel pdiffusion 1207 -251 1207 -251 0 feedthrough
rlabel pdiffusion 1214 -251 1214 -251 0 cellNo=303
rlabel pdiffusion 1221 -251 1221 -251 0 feedthrough
rlabel pdiffusion 1228 -251 1228 -251 0 feedthrough
rlabel pdiffusion 1235 -251 1235 -251 0 feedthrough
rlabel pdiffusion 1242 -251 1242 -251 0 feedthrough
rlabel pdiffusion 1249 -251 1249 -251 0 feedthrough
rlabel pdiffusion 1256 -251 1256 -251 0 feedthrough
rlabel pdiffusion 1263 -251 1263 -251 0 feedthrough
rlabel pdiffusion 1270 -251 1270 -251 0 feedthrough
rlabel pdiffusion 1277 -251 1277 -251 0 feedthrough
rlabel pdiffusion 1284 -251 1284 -251 0 feedthrough
rlabel pdiffusion 1291 -251 1291 -251 0 feedthrough
rlabel pdiffusion 1298 -251 1298 -251 0 feedthrough
rlabel pdiffusion 1305 -251 1305 -251 0 feedthrough
rlabel pdiffusion 1312 -251 1312 -251 0 feedthrough
rlabel pdiffusion 1319 -251 1319 -251 0 feedthrough
rlabel pdiffusion 1326 -251 1326 -251 0 cellNo=446
rlabel pdiffusion 1333 -251 1333 -251 0 feedthrough
rlabel pdiffusion 1340 -251 1340 -251 0 feedthrough
rlabel pdiffusion 1347 -251 1347 -251 0 feedthrough
rlabel pdiffusion 1354 -251 1354 -251 0 feedthrough
rlabel pdiffusion 1361 -251 1361 -251 0 feedthrough
rlabel pdiffusion 1368 -251 1368 -251 0 feedthrough
rlabel pdiffusion 1375 -251 1375 -251 0 feedthrough
rlabel pdiffusion 1382 -251 1382 -251 0 feedthrough
rlabel pdiffusion 1389 -251 1389 -251 0 feedthrough
rlabel pdiffusion 1396 -251 1396 -251 0 feedthrough
rlabel pdiffusion 1403 -251 1403 -251 0 feedthrough
rlabel pdiffusion 1410 -251 1410 -251 0 feedthrough
rlabel pdiffusion 1417 -251 1417 -251 0 feedthrough
rlabel pdiffusion 1424 -251 1424 -251 0 feedthrough
rlabel pdiffusion 1431 -251 1431 -251 0 feedthrough
rlabel pdiffusion 1438 -251 1438 -251 0 feedthrough
rlabel pdiffusion 1445 -251 1445 -251 0 feedthrough
rlabel pdiffusion 1452 -251 1452 -251 0 feedthrough
rlabel pdiffusion 1459 -251 1459 -251 0 feedthrough
rlabel pdiffusion 1466 -251 1466 -251 0 feedthrough
rlabel pdiffusion 1473 -251 1473 -251 0 feedthrough
rlabel pdiffusion 1480 -251 1480 -251 0 feedthrough
rlabel pdiffusion 1487 -251 1487 -251 0 feedthrough
rlabel pdiffusion 1494 -251 1494 -251 0 feedthrough
rlabel pdiffusion 1501 -251 1501 -251 0 feedthrough
rlabel pdiffusion 1508 -251 1508 -251 0 feedthrough
rlabel pdiffusion 1515 -251 1515 -251 0 feedthrough
rlabel pdiffusion 1522 -251 1522 -251 0 feedthrough
rlabel pdiffusion 1529 -251 1529 -251 0 feedthrough
rlabel pdiffusion 1536 -251 1536 -251 0 feedthrough
rlabel pdiffusion 1543 -251 1543 -251 0 cellNo=675
rlabel pdiffusion 1550 -251 1550 -251 0 cellNo=278
rlabel pdiffusion 1557 -251 1557 -251 0 feedthrough
rlabel pdiffusion 1564 -251 1564 -251 0 cellNo=420
rlabel pdiffusion 1571 -251 1571 -251 0 feedthrough
rlabel pdiffusion 1578 -251 1578 -251 0 feedthrough
rlabel pdiffusion 1585 -251 1585 -251 0 feedthrough
rlabel pdiffusion 1592 -251 1592 -251 0 feedthrough
rlabel pdiffusion 1613 -251 1613 -251 0 cellNo=468
rlabel pdiffusion 1627 -251 1627 -251 0 feedthrough
rlabel pdiffusion 1634 -251 1634 -251 0 feedthrough
rlabel pdiffusion 1669 -251 1669 -251 0 feedthrough
rlabel pdiffusion 1816 -251 1816 -251 0 feedthrough
rlabel pdiffusion 1942 -251 1942 -251 0 feedthrough
rlabel pdiffusion 3 -376 3 -376 0 cellNo=1035
rlabel pdiffusion 10 -376 10 -376 0 cellNo=1193
rlabel pdiffusion 17 -376 17 -376 0 feedthrough
rlabel pdiffusion 24 -376 24 -376 0 feedthrough
rlabel pdiffusion 31 -376 31 -376 0 feedthrough
rlabel pdiffusion 38 -376 38 -376 0 feedthrough
rlabel pdiffusion 45 -376 45 -376 0 cellNo=709
rlabel pdiffusion 52 -376 52 -376 0 cellNo=667
rlabel pdiffusion 59 -376 59 -376 0 feedthrough
rlabel pdiffusion 66 -376 66 -376 0 feedthrough
rlabel pdiffusion 73 -376 73 -376 0 feedthrough
rlabel pdiffusion 80 -376 80 -376 0 feedthrough
rlabel pdiffusion 87 -376 87 -376 0 feedthrough
rlabel pdiffusion 94 -376 94 -376 0 cellNo=157
rlabel pdiffusion 101 -376 101 -376 0 feedthrough
rlabel pdiffusion 108 -376 108 -376 0 feedthrough
rlabel pdiffusion 115 -376 115 -376 0 feedthrough
rlabel pdiffusion 122 -376 122 -376 0 feedthrough
rlabel pdiffusion 129 -376 129 -376 0 feedthrough
rlabel pdiffusion 136 -376 136 -376 0 cellNo=137
rlabel pdiffusion 143 -376 143 -376 0 feedthrough
rlabel pdiffusion 150 -376 150 -376 0 feedthrough
rlabel pdiffusion 157 -376 157 -376 0 feedthrough
rlabel pdiffusion 164 -376 164 -376 0 cellNo=782
rlabel pdiffusion 171 -376 171 -376 0 feedthrough
rlabel pdiffusion 178 -376 178 -376 0 feedthrough
rlabel pdiffusion 185 -376 185 -376 0 cellNo=264
rlabel pdiffusion 192 -376 192 -376 0 cellNo=57
rlabel pdiffusion 199 -376 199 -376 0 feedthrough
rlabel pdiffusion 206 -376 206 -376 0 feedthrough
rlabel pdiffusion 213 -376 213 -376 0 feedthrough
rlabel pdiffusion 220 -376 220 -376 0 feedthrough
rlabel pdiffusion 227 -376 227 -376 0 feedthrough
rlabel pdiffusion 234 -376 234 -376 0 feedthrough
rlabel pdiffusion 241 -376 241 -376 0 cellNo=272
rlabel pdiffusion 248 -376 248 -376 0 feedthrough
rlabel pdiffusion 255 -376 255 -376 0 feedthrough
rlabel pdiffusion 262 -376 262 -376 0 feedthrough
rlabel pdiffusion 269 -376 269 -376 0 feedthrough
rlabel pdiffusion 276 -376 276 -376 0 feedthrough
rlabel pdiffusion 283 -376 283 -376 0 feedthrough
rlabel pdiffusion 290 -376 290 -376 0 feedthrough
rlabel pdiffusion 297 -376 297 -376 0 feedthrough
rlabel pdiffusion 304 -376 304 -376 0 feedthrough
rlabel pdiffusion 311 -376 311 -376 0 feedthrough
rlabel pdiffusion 318 -376 318 -376 0 feedthrough
rlabel pdiffusion 325 -376 325 -376 0 feedthrough
rlabel pdiffusion 332 -376 332 -376 0 feedthrough
rlabel pdiffusion 339 -376 339 -376 0 feedthrough
rlabel pdiffusion 346 -376 346 -376 0 feedthrough
rlabel pdiffusion 353 -376 353 -376 0 feedthrough
rlabel pdiffusion 360 -376 360 -376 0 feedthrough
rlabel pdiffusion 367 -376 367 -376 0 feedthrough
rlabel pdiffusion 374 -376 374 -376 0 feedthrough
rlabel pdiffusion 381 -376 381 -376 0 feedthrough
rlabel pdiffusion 388 -376 388 -376 0 feedthrough
rlabel pdiffusion 395 -376 395 -376 0 feedthrough
rlabel pdiffusion 402 -376 402 -376 0 cellNo=132
rlabel pdiffusion 409 -376 409 -376 0 feedthrough
rlabel pdiffusion 416 -376 416 -376 0 feedthrough
rlabel pdiffusion 423 -376 423 -376 0 feedthrough
rlabel pdiffusion 430 -376 430 -376 0 cellNo=394
rlabel pdiffusion 437 -376 437 -376 0 feedthrough
rlabel pdiffusion 444 -376 444 -376 0 cellNo=345
rlabel pdiffusion 451 -376 451 -376 0 feedthrough
rlabel pdiffusion 458 -376 458 -376 0 feedthrough
rlabel pdiffusion 465 -376 465 -376 0 feedthrough
rlabel pdiffusion 472 -376 472 -376 0 feedthrough
rlabel pdiffusion 479 -376 479 -376 0 cellNo=563
rlabel pdiffusion 486 -376 486 -376 0 feedthrough
rlabel pdiffusion 493 -376 493 -376 0 feedthrough
rlabel pdiffusion 500 -376 500 -376 0 feedthrough
rlabel pdiffusion 507 -376 507 -376 0 feedthrough
rlabel pdiffusion 514 -376 514 -376 0 feedthrough
rlabel pdiffusion 521 -376 521 -376 0 feedthrough
rlabel pdiffusion 528 -376 528 -376 0 feedthrough
rlabel pdiffusion 535 -376 535 -376 0 feedthrough
rlabel pdiffusion 542 -376 542 -376 0 feedthrough
rlabel pdiffusion 549 -376 549 -376 0 feedthrough
rlabel pdiffusion 556 -376 556 -376 0 feedthrough
rlabel pdiffusion 563 -376 563 -376 0 feedthrough
rlabel pdiffusion 570 -376 570 -376 0 feedthrough
rlabel pdiffusion 577 -376 577 -376 0 feedthrough
rlabel pdiffusion 584 -376 584 -376 0 feedthrough
rlabel pdiffusion 591 -376 591 -376 0 feedthrough
rlabel pdiffusion 598 -376 598 -376 0 feedthrough
rlabel pdiffusion 605 -376 605 -376 0 feedthrough
rlabel pdiffusion 612 -376 612 -376 0 feedthrough
rlabel pdiffusion 619 -376 619 -376 0 feedthrough
rlabel pdiffusion 626 -376 626 -376 0 cellNo=115
rlabel pdiffusion 633 -376 633 -376 0 cellNo=811
rlabel pdiffusion 640 -376 640 -376 0 feedthrough
rlabel pdiffusion 647 -376 647 -376 0 cellNo=509
rlabel pdiffusion 654 -376 654 -376 0 feedthrough
rlabel pdiffusion 661 -376 661 -376 0 feedthrough
rlabel pdiffusion 668 -376 668 -376 0 feedthrough
rlabel pdiffusion 675 -376 675 -376 0 feedthrough
rlabel pdiffusion 682 -376 682 -376 0 feedthrough
rlabel pdiffusion 689 -376 689 -376 0 feedthrough
rlabel pdiffusion 696 -376 696 -376 0 feedthrough
rlabel pdiffusion 703 -376 703 -376 0 feedthrough
rlabel pdiffusion 710 -376 710 -376 0 feedthrough
rlabel pdiffusion 717 -376 717 -376 0 feedthrough
rlabel pdiffusion 724 -376 724 -376 0 feedthrough
rlabel pdiffusion 731 -376 731 -376 0 feedthrough
rlabel pdiffusion 738 -376 738 -376 0 feedthrough
rlabel pdiffusion 745 -376 745 -376 0 cellNo=159
rlabel pdiffusion 752 -376 752 -376 0 feedthrough
rlabel pdiffusion 759 -376 759 -376 0 cellNo=85
rlabel pdiffusion 766 -376 766 -376 0 feedthrough
rlabel pdiffusion 773 -376 773 -376 0 cellNo=109
rlabel pdiffusion 780 -376 780 -376 0 feedthrough
rlabel pdiffusion 787 -376 787 -376 0 feedthrough
rlabel pdiffusion 794 -376 794 -376 0 cellNo=414
rlabel pdiffusion 801 -376 801 -376 0 cellNo=275
rlabel pdiffusion 808 -376 808 -376 0 cellNo=181
rlabel pdiffusion 815 -376 815 -376 0 feedthrough
rlabel pdiffusion 822 -376 822 -376 0 feedthrough
rlabel pdiffusion 829 -376 829 -376 0 feedthrough
rlabel pdiffusion 836 -376 836 -376 0 cellNo=458
rlabel pdiffusion 843 -376 843 -376 0 cellNo=263
rlabel pdiffusion 850 -376 850 -376 0 feedthrough
rlabel pdiffusion 857 -376 857 -376 0 feedthrough
rlabel pdiffusion 864 -376 864 -376 0 feedthrough
rlabel pdiffusion 871 -376 871 -376 0 feedthrough
rlabel pdiffusion 878 -376 878 -376 0 cellNo=308
rlabel pdiffusion 885 -376 885 -376 0 feedthrough
rlabel pdiffusion 892 -376 892 -376 0 cellNo=91
rlabel pdiffusion 899 -376 899 -376 0 feedthrough
rlabel pdiffusion 906 -376 906 -376 0 feedthrough
rlabel pdiffusion 913 -376 913 -376 0 feedthrough
rlabel pdiffusion 920 -376 920 -376 0 feedthrough
rlabel pdiffusion 927 -376 927 -376 0 feedthrough
rlabel pdiffusion 934 -376 934 -376 0 feedthrough
rlabel pdiffusion 941 -376 941 -376 0 feedthrough
rlabel pdiffusion 948 -376 948 -376 0 feedthrough
rlabel pdiffusion 955 -376 955 -376 0 feedthrough
rlabel pdiffusion 962 -376 962 -376 0 feedthrough
rlabel pdiffusion 969 -376 969 -376 0 feedthrough
rlabel pdiffusion 976 -376 976 -376 0 cellNo=215
rlabel pdiffusion 983 -376 983 -376 0 feedthrough
rlabel pdiffusion 990 -376 990 -376 0 cellNo=528
rlabel pdiffusion 997 -376 997 -376 0 feedthrough
rlabel pdiffusion 1004 -376 1004 -376 0 feedthrough
rlabel pdiffusion 1011 -376 1011 -376 0 feedthrough
rlabel pdiffusion 1018 -376 1018 -376 0 cellNo=292
rlabel pdiffusion 1025 -376 1025 -376 0 cellNo=928
rlabel pdiffusion 1032 -376 1032 -376 0 feedthrough
rlabel pdiffusion 1039 -376 1039 -376 0 feedthrough
rlabel pdiffusion 1046 -376 1046 -376 0 feedthrough
rlabel pdiffusion 1053 -376 1053 -376 0 feedthrough
rlabel pdiffusion 1060 -376 1060 -376 0 feedthrough
rlabel pdiffusion 1067 -376 1067 -376 0 feedthrough
rlabel pdiffusion 1074 -376 1074 -376 0 cellNo=164
rlabel pdiffusion 1081 -376 1081 -376 0 cellNo=210
rlabel pdiffusion 1088 -376 1088 -376 0 feedthrough
rlabel pdiffusion 1095 -376 1095 -376 0 feedthrough
rlabel pdiffusion 1102 -376 1102 -376 0 cellNo=508
rlabel pdiffusion 1109 -376 1109 -376 0 feedthrough
rlabel pdiffusion 1116 -376 1116 -376 0 feedthrough
rlabel pdiffusion 1123 -376 1123 -376 0 feedthrough
rlabel pdiffusion 1130 -376 1130 -376 0 feedthrough
rlabel pdiffusion 1137 -376 1137 -376 0 feedthrough
rlabel pdiffusion 1144 -376 1144 -376 0 feedthrough
rlabel pdiffusion 1151 -376 1151 -376 0 feedthrough
rlabel pdiffusion 1158 -376 1158 -376 0 feedthrough
rlabel pdiffusion 1165 -376 1165 -376 0 feedthrough
rlabel pdiffusion 1172 -376 1172 -376 0 feedthrough
rlabel pdiffusion 1179 -376 1179 -376 0 cellNo=530
rlabel pdiffusion 1186 -376 1186 -376 0 feedthrough
rlabel pdiffusion 1193 -376 1193 -376 0 feedthrough
rlabel pdiffusion 1200 -376 1200 -376 0 feedthrough
rlabel pdiffusion 1207 -376 1207 -376 0 feedthrough
rlabel pdiffusion 1214 -376 1214 -376 0 feedthrough
rlabel pdiffusion 1221 -376 1221 -376 0 feedthrough
rlabel pdiffusion 1228 -376 1228 -376 0 feedthrough
rlabel pdiffusion 1235 -376 1235 -376 0 feedthrough
rlabel pdiffusion 1242 -376 1242 -376 0 feedthrough
rlabel pdiffusion 1249 -376 1249 -376 0 feedthrough
rlabel pdiffusion 1256 -376 1256 -376 0 feedthrough
rlabel pdiffusion 1263 -376 1263 -376 0 feedthrough
rlabel pdiffusion 1270 -376 1270 -376 0 feedthrough
rlabel pdiffusion 1277 -376 1277 -376 0 feedthrough
rlabel pdiffusion 1284 -376 1284 -376 0 feedthrough
rlabel pdiffusion 1291 -376 1291 -376 0 feedthrough
rlabel pdiffusion 1298 -376 1298 -376 0 feedthrough
rlabel pdiffusion 1305 -376 1305 -376 0 feedthrough
rlabel pdiffusion 1312 -376 1312 -376 0 feedthrough
rlabel pdiffusion 1319 -376 1319 -376 0 feedthrough
rlabel pdiffusion 1326 -376 1326 -376 0 cellNo=891
rlabel pdiffusion 1333 -376 1333 -376 0 feedthrough
rlabel pdiffusion 1340 -376 1340 -376 0 feedthrough
rlabel pdiffusion 1347 -376 1347 -376 0 feedthrough
rlabel pdiffusion 1354 -376 1354 -376 0 cellNo=118
rlabel pdiffusion 1361 -376 1361 -376 0 feedthrough
rlabel pdiffusion 1368 -376 1368 -376 0 feedthrough
rlabel pdiffusion 1375 -376 1375 -376 0 feedthrough
rlabel pdiffusion 1382 -376 1382 -376 0 feedthrough
rlabel pdiffusion 1389 -376 1389 -376 0 feedthrough
rlabel pdiffusion 1396 -376 1396 -376 0 feedthrough
rlabel pdiffusion 1403 -376 1403 -376 0 feedthrough
rlabel pdiffusion 1410 -376 1410 -376 0 feedthrough
rlabel pdiffusion 1417 -376 1417 -376 0 feedthrough
rlabel pdiffusion 1424 -376 1424 -376 0 feedthrough
rlabel pdiffusion 1431 -376 1431 -376 0 feedthrough
rlabel pdiffusion 1438 -376 1438 -376 0 feedthrough
rlabel pdiffusion 1445 -376 1445 -376 0 feedthrough
rlabel pdiffusion 1452 -376 1452 -376 0 feedthrough
rlabel pdiffusion 1459 -376 1459 -376 0 feedthrough
rlabel pdiffusion 1466 -376 1466 -376 0 feedthrough
rlabel pdiffusion 1473 -376 1473 -376 0 feedthrough
rlabel pdiffusion 1480 -376 1480 -376 0 feedthrough
rlabel pdiffusion 1487 -376 1487 -376 0 feedthrough
rlabel pdiffusion 1494 -376 1494 -376 0 feedthrough
rlabel pdiffusion 1501 -376 1501 -376 0 feedthrough
rlabel pdiffusion 1508 -376 1508 -376 0 feedthrough
rlabel pdiffusion 1515 -376 1515 -376 0 feedthrough
rlabel pdiffusion 1522 -376 1522 -376 0 feedthrough
rlabel pdiffusion 1529 -376 1529 -376 0 feedthrough
rlabel pdiffusion 1536 -376 1536 -376 0 feedthrough
rlabel pdiffusion 1543 -376 1543 -376 0 feedthrough
rlabel pdiffusion 1550 -376 1550 -376 0 feedthrough
rlabel pdiffusion 1557 -376 1557 -376 0 feedthrough
rlabel pdiffusion 1564 -376 1564 -376 0 feedthrough
rlabel pdiffusion 1571 -376 1571 -376 0 feedthrough
rlabel pdiffusion 1578 -376 1578 -376 0 feedthrough
rlabel pdiffusion 1585 -376 1585 -376 0 feedthrough
rlabel pdiffusion 1592 -376 1592 -376 0 feedthrough
rlabel pdiffusion 1599 -376 1599 -376 0 feedthrough
rlabel pdiffusion 1606 -376 1606 -376 0 feedthrough
rlabel pdiffusion 1613 -376 1613 -376 0 cellNo=302
rlabel pdiffusion 1620 -376 1620 -376 0 feedthrough
rlabel pdiffusion 1627 -376 1627 -376 0 feedthrough
rlabel pdiffusion 1634 -376 1634 -376 0 feedthrough
rlabel pdiffusion 1641 -376 1641 -376 0 feedthrough
rlabel pdiffusion 1648 -376 1648 -376 0 feedthrough
rlabel pdiffusion 1655 -376 1655 -376 0 feedthrough
rlabel pdiffusion 1662 -376 1662 -376 0 feedthrough
rlabel pdiffusion 1669 -376 1669 -376 0 feedthrough
rlabel pdiffusion 1676 -376 1676 -376 0 feedthrough
rlabel pdiffusion 1683 -376 1683 -376 0 feedthrough
rlabel pdiffusion 1690 -376 1690 -376 0 feedthrough
rlabel pdiffusion 1697 -376 1697 -376 0 feedthrough
rlabel pdiffusion 1704 -376 1704 -376 0 feedthrough
rlabel pdiffusion 1711 -376 1711 -376 0 feedthrough
rlabel pdiffusion 1718 -376 1718 -376 0 feedthrough
rlabel pdiffusion 1725 -376 1725 -376 0 feedthrough
rlabel pdiffusion 1732 -376 1732 -376 0 feedthrough
rlabel pdiffusion 1739 -376 1739 -376 0 feedthrough
rlabel pdiffusion 1746 -376 1746 -376 0 feedthrough
rlabel pdiffusion 1753 -376 1753 -376 0 feedthrough
rlabel pdiffusion 1760 -376 1760 -376 0 feedthrough
rlabel pdiffusion 1767 -376 1767 -376 0 feedthrough
rlabel pdiffusion 1774 -376 1774 -376 0 feedthrough
rlabel pdiffusion 1781 -376 1781 -376 0 feedthrough
rlabel pdiffusion 1788 -376 1788 -376 0 feedthrough
rlabel pdiffusion 1795 -376 1795 -376 0 feedthrough
rlabel pdiffusion 1802 -376 1802 -376 0 feedthrough
rlabel pdiffusion 1809 -376 1809 -376 0 feedthrough
rlabel pdiffusion 1816 -376 1816 -376 0 feedthrough
rlabel pdiffusion 1823 -376 1823 -376 0 feedthrough
rlabel pdiffusion 1830 -376 1830 -376 0 feedthrough
rlabel pdiffusion 1837 -376 1837 -376 0 feedthrough
rlabel pdiffusion 1844 -376 1844 -376 0 feedthrough
rlabel pdiffusion 1928 -376 1928 -376 0 feedthrough
rlabel pdiffusion 1963 -376 1963 -376 0 cellNo=184
rlabel pdiffusion 1970 -376 1970 -376 0 feedthrough
rlabel pdiffusion 1984 -376 1984 -376 0 feedthrough
rlabel pdiffusion 2005 -376 2005 -376 0 feedthrough
rlabel pdiffusion 2194 -376 2194 -376 0 feedthrough
rlabel pdiffusion 3 -505 3 -505 0 feedthrough
rlabel pdiffusion 10 -505 10 -505 0 cellNo=234
rlabel pdiffusion 17 -505 17 -505 0 feedthrough
rlabel pdiffusion 24 -505 24 -505 0 feedthrough
rlabel pdiffusion 31 -505 31 -505 0 cellNo=1197
rlabel pdiffusion 38 -505 38 -505 0 cellNo=1034
rlabel pdiffusion 45 -505 45 -505 0 feedthrough
rlabel pdiffusion 52 -505 52 -505 0 feedthrough
rlabel pdiffusion 59 -505 59 -505 0 cellNo=555
rlabel pdiffusion 66 -505 66 -505 0 feedthrough
rlabel pdiffusion 73 -505 73 -505 0 feedthrough
rlabel pdiffusion 80 -505 80 -505 0 feedthrough
rlabel pdiffusion 87 -505 87 -505 0 feedthrough
rlabel pdiffusion 94 -505 94 -505 0 feedthrough
rlabel pdiffusion 101 -505 101 -505 0 feedthrough
rlabel pdiffusion 108 -505 108 -505 0 feedthrough
rlabel pdiffusion 115 -505 115 -505 0 cellNo=518
rlabel pdiffusion 122 -505 122 -505 0 feedthrough
rlabel pdiffusion 129 -505 129 -505 0 feedthrough
rlabel pdiffusion 136 -505 136 -505 0 feedthrough
rlabel pdiffusion 143 -505 143 -505 0 feedthrough
rlabel pdiffusion 150 -505 150 -505 0 feedthrough
rlabel pdiffusion 157 -505 157 -505 0 feedthrough
rlabel pdiffusion 164 -505 164 -505 0 cellNo=842
rlabel pdiffusion 171 -505 171 -505 0 cellNo=248
rlabel pdiffusion 178 -505 178 -505 0 feedthrough
rlabel pdiffusion 185 -505 185 -505 0 feedthrough
rlabel pdiffusion 192 -505 192 -505 0 feedthrough
rlabel pdiffusion 199 -505 199 -505 0 feedthrough
rlabel pdiffusion 206 -505 206 -505 0 feedthrough
rlabel pdiffusion 213 -505 213 -505 0 cellNo=45
rlabel pdiffusion 220 -505 220 -505 0 cellNo=461
rlabel pdiffusion 227 -505 227 -505 0 feedthrough
rlabel pdiffusion 234 -505 234 -505 0 cellNo=455
rlabel pdiffusion 241 -505 241 -505 0 feedthrough
rlabel pdiffusion 248 -505 248 -505 0 feedthrough
rlabel pdiffusion 255 -505 255 -505 0 feedthrough
rlabel pdiffusion 262 -505 262 -505 0 feedthrough
rlabel pdiffusion 269 -505 269 -505 0 feedthrough
rlabel pdiffusion 276 -505 276 -505 0 feedthrough
rlabel pdiffusion 283 -505 283 -505 0 feedthrough
rlabel pdiffusion 290 -505 290 -505 0 feedthrough
rlabel pdiffusion 297 -505 297 -505 0 feedthrough
rlabel pdiffusion 304 -505 304 -505 0 feedthrough
rlabel pdiffusion 311 -505 311 -505 0 feedthrough
rlabel pdiffusion 318 -505 318 -505 0 feedthrough
rlabel pdiffusion 325 -505 325 -505 0 feedthrough
rlabel pdiffusion 332 -505 332 -505 0 feedthrough
rlabel pdiffusion 339 -505 339 -505 0 feedthrough
rlabel pdiffusion 346 -505 346 -505 0 feedthrough
rlabel pdiffusion 353 -505 353 -505 0 feedthrough
rlabel pdiffusion 360 -505 360 -505 0 feedthrough
rlabel pdiffusion 367 -505 367 -505 0 feedthrough
rlabel pdiffusion 374 -505 374 -505 0 feedthrough
rlabel pdiffusion 381 -505 381 -505 0 feedthrough
rlabel pdiffusion 388 -505 388 -505 0 feedthrough
rlabel pdiffusion 395 -505 395 -505 0 feedthrough
rlabel pdiffusion 402 -505 402 -505 0 feedthrough
rlabel pdiffusion 409 -505 409 -505 0 feedthrough
rlabel pdiffusion 416 -505 416 -505 0 feedthrough
rlabel pdiffusion 423 -505 423 -505 0 feedthrough
rlabel pdiffusion 430 -505 430 -505 0 feedthrough
rlabel pdiffusion 437 -505 437 -505 0 feedthrough
rlabel pdiffusion 444 -505 444 -505 0 feedthrough
rlabel pdiffusion 451 -505 451 -505 0 feedthrough
rlabel pdiffusion 458 -505 458 -505 0 feedthrough
rlabel pdiffusion 465 -505 465 -505 0 feedthrough
rlabel pdiffusion 472 -505 472 -505 0 feedthrough
rlabel pdiffusion 479 -505 479 -505 0 feedthrough
rlabel pdiffusion 486 -505 486 -505 0 feedthrough
rlabel pdiffusion 493 -505 493 -505 0 cellNo=300
rlabel pdiffusion 500 -505 500 -505 0 feedthrough
rlabel pdiffusion 507 -505 507 -505 0 feedthrough
rlabel pdiffusion 514 -505 514 -505 0 feedthrough
rlabel pdiffusion 521 -505 521 -505 0 feedthrough
rlabel pdiffusion 528 -505 528 -505 0 feedthrough
rlabel pdiffusion 535 -505 535 -505 0 cellNo=77
rlabel pdiffusion 542 -505 542 -505 0 feedthrough
rlabel pdiffusion 549 -505 549 -505 0 feedthrough
rlabel pdiffusion 556 -505 556 -505 0 feedthrough
rlabel pdiffusion 563 -505 563 -505 0 feedthrough
rlabel pdiffusion 570 -505 570 -505 0 feedthrough
rlabel pdiffusion 577 -505 577 -505 0 feedthrough
rlabel pdiffusion 584 -505 584 -505 0 feedthrough
rlabel pdiffusion 591 -505 591 -505 0 feedthrough
rlabel pdiffusion 598 -505 598 -505 0 cellNo=564
rlabel pdiffusion 605 -505 605 -505 0 feedthrough
rlabel pdiffusion 612 -505 612 -505 0 feedthrough
rlabel pdiffusion 619 -505 619 -505 0 cellNo=287
rlabel pdiffusion 626 -505 626 -505 0 feedthrough
rlabel pdiffusion 633 -505 633 -505 0 cellNo=252
rlabel pdiffusion 640 -505 640 -505 0 feedthrough
rlabel pdiffusion 647 -505 647 -505 0 feedthrough
rlabel pdiffusion 654 -505 654 -505 0 cellNo=66
rlabel pdiffusion 661 -505 661 -505 0 feedthrough
rlabel pdiffusion 668 -505 668 -505 0 feedthrough
rlabel pdiffusion 675 -505 675 -505 0 feedthrough
rlabel pdiffusion 682 -505 682 -505 0 feedthrough
rlabel pdiffusion 689 -505 689 -505 0 feedthrough
rlabel pdiffusion 696 -505 696 -505 0 feedthrough
rlabel pdiffusion 703 -505 703 -505 0 feedthrough
rlabel pdiffusion 710 -505 710 -505 0 feedthrough
rlabel pdiffusion 717 -505 717 -505 0 cellNo=78
rlabel pdiffusion 724 -505 724 -505 0 cellNo=739
rlabel pdiffusion 731 -505 731 -505 0 feedthrough
rlabel pdiffusion 738 -505 738 -505 0 cellNo=398
rlabel pdiffusion 745 -505 745 -505 0 feedthrough
rlabel pdiffusion 752 -505 752 -505 0 feedthrough
rlabel pdiffusion 759 -505 759 -505 0 feedthrough
rlabel pdiffusion 766 -505 766 -505 0 feedthrough
rlabel pdiffusion 773 -505 773 -505 0 feedthrough
rlabel pdiffusion 780 -505 780 -505 0 feedthrough
rlabel pdiffusion 787 -505 787 -505 0 feedthrough
rlabel pdiffusion 794 -505 794 -505 0 feedthrough
rlabel pdiffusion 801 -505 801 -505 0 feedthrough
rlabel pdiffusion 808 -505 808 -505 0 feedthrough
rlabel pdiffusion 815 -505 815 -505 0 feedthrough
rlabel pdiffusion 822 -505 822 -505 0 feedthrough
rlabel pdiffusion 829 -505 829 -505 0 feedthrough
rlabel pdiffusion 836 -505 836 -505 0 feedthrough
rlabel pdiffusion 843 -505 843 -505 0 feedthrough
rlabel pdiffusion 850 -505 850 -505 0 cellNo=11
rlabel pdiffusion 857 -505 857 -505 0 feedthrough
rlabel pdiffusion 864 -505 864 -505 0 feedthrough
rlabel pdiffusion 871 -505 871 -505 0 feedthrough
rlabel pdiffusion 878 -505 878 -505 0 feedthrough
rlabel pdiffusion 885 -505 885 -505 0 cellNo=20
rlabel pdiffusion 892 -505 892 -505 0 feedthrough
rlabel pdiffusion 899 -505 899 -505 0 feedthrough
rlabel pdiffusion 906 -505 906 -505 0 feedthrough
rlabel pdiffusion 913 -505 913 -505 0 cellNo=124
rlabel pdiffusion 920 -505 920 -505 0 feedthrough
rlabel pdiffusion 927 -505 927 -505 0 feedthrough
rlabel pdiffusion 934 -505 934 -505 0 cellNo=787
rlabel pdiffusion 941 -505 941 -505 0 feedthrough
rlabel pdiffusion 948 -505 948 -505 0 feedthrough
rlabel pdiffusion 955 -505 955 -505 0 cellNo=271
rlabel pdiffusion 962 -505 962 -505 0 feedthrough
rlabel pdiffusion 969 -505 969 -505 0 cellNo=265
rlabel pdiffusion 976 -505 976 -505 0 cellNo=147
rlabel pdiffusion 983 -505 983 -505 0 cellNo=717
rlabel pdiffusion 990 -505 990 -505 0 cellNo=728
rlabel pdiffusion 997 -505 997 -505 0 feedthrough
rlabel pdiffusion 1004 -505 1004 -505 0 cellNo=847
rlabel pdiffusion 1011 -505 1011 -505 0 feedthrough
rlabel pdiffusion 1018 -505 1018 -505 0 feedthrough
rlabel pdiffusion 1025 -505 1025 -505 0 cellNo=167
rlabel pdiffusion 1032 -505 1032 -505 0 feedthrough
rlabel pdiffusion 1039 -505 1039 -505 0 feedthrough
rlabel pdiffusion 1046 -505 1046 -505 0 feedthrough
rlabel pdiffusion 1053 -505 1053 -505 0 feedthrough
rlabel pdiffusion 1060 -505 1060 -505 0 feedthrough
rlabel pdiffusion 1067 -505 1067 -505 0 feedthrough
rlabel pdiffusion 1074 -505 1074 -505 0 feedthrough
rlabel pdiffusion 1081 -505 1081 -505 0 cellNo=536
rlabel pdiffusion 1088 -505 1088 -505 0 feedthrough
rlabel pdiffusion 1095 -505 1095 -505 0 feedthrough
rlabel pdiffusion 1102 -505 1102 -505 0 feedthrough
rlabel pdiffusion 1109 -505 1109 -505 0 feedthrough
rlabel pdiffusion 1116 -505 1116 -505 0 feedthrough
rlabel pdiffusion 1123 -505 1123 -505 0 cellNo=603
rlabel pdiffusion 1130 -505 1130 -505 0 feedthrough
rlabel pdiffusion 1137 -505 1137 -505 0 feedthrough
rlabel pdiffusion 1144 -505 1144 -505 0 feedthrough
rlabel pdiffusion 1151 -505 1151 -505 0 feedthrough
rlabel pdiffusion 1158 -505 1158 -505 0 feedthrough
rlabel pdiffusion 1165 -505 1165 -505 0 cellNo=818
rlabel pdiffusion 1172 -505 1172 -505 0 feedthrough
rlabel pdiffusion 1179 -505 1179 -505 0 feedthrough
rlabel pdiffusion 1186 -505 1186 -505 0 feedthrough
rlabel pdiffusion 1193 -505 1193 -505 0 feedthrough
rlabel pdiffusion 1200 -505 1200 -505 0 feedthrough
rlabel pdiffusion 1207 -505 1207 -505 0 feedthrough
rlabel pdiffusion 1214 -505 1214 -505 0 feedthrough
rlabel pdiffusion 1221 -505 1221 -505 0 feedthrough
rlabel pdiffusion 1228 -505 1228 -505 0 feedthrough
rlabel pdiffusion 1235 -505 1235 -505 0 feedthrough
rlabel pdiffusion 1242 -505 1242 -505 0 feedthrough
rlabel pdiffusion 1249 -505 1249 -505 0 feedthrough
rlabel pdiffusion 1256 -505 1256 -505 0 feedthrough
rlabel pdiffusion 1263 -505 1263 -505 0 feedthrough
rlabel pdiffusion 1270 -505 1270 -505 0 feedthrough
rlabel pdiffusion 1277 -505 1277 -505 0 feedthrough
rlabel pdiffusion 1284 -505 1284 -505 0 feedthrough
rlabel pdiffusion 1291 -505 1291 -505 0 feedthrough
rlabel pdiffusion 1298 -505 1298 -505 0 feedthrough
rlabel pdiffusion 1305 -505 1305 -505 0 feedthrough
rlabel pdiffusion 1312 -505 1312 -505 0 feedthrough
rlabel pdiffusion 1319 -505 1319 -505 0 feedthrough
rlabel pdiffusion 1326 -505 1326 -505 0 feedthrough
rlabel pdiffusion 1333 -505 1333 -505 0 feedthrough
rlabel pdiffusion 1340 -505 1340 -505 0 feedthrough
rlabel pdiffusion 1347 -505 1347 -505 0 feedthrough
rlabel pdiffusion 1354 -505 1354 -505 0 feedthrough
rlabel pdiffusion 1361 -505 1361 -505 0 feedthrough
rlabel pdiffusion 1368 -505 1368 -505 0 feedthrough
rlabel pdiffusion 1375 -505 1375 -505 0 feedthrough
rlabel pdiffusion 1382 -505 1382 -505 0 feedthrough
rlabel pdiffusion 1389 -505 1389 -505 0 feedthrough
rlabel pdiffusion 1396 -505 1396 -505 0 feedthrough
rlabel pdiffusion 1403 -505 1403 -505 0 feedthrough
rlabel pdiffusion 1410 -505 1410 -505 0 feedthrough
rlabel pdiffusion 1417 -505 1417 -505 0 feedthrough
rlabel pdiffusion 1424 -505 1424 -505 0 feedthrough
rlabel pdiffusion 1431 -505 1431 -505 0 feedthrough
rlabel pdiffusion 1438 -505 1438 -505 0 cellNo=742
rlabel pdiffusion 1445 -505 1445 -505 0 feedthrough
rlabel pdiffusion 1452 -505 1452 -505 0 feedthrough
rlabel pdiffusion 1459 -505 1459 -505 0 feedthrough
rlabel pdiffusion 1466 -505 1466 -505 0 feedthrough
rlabel pdiffusion 1473 -505 1473 -505 0 feedthrough
rlabel pdiffusion 1480 -505 1480 -505 0 feedthrough
rlabel pdiffusion 1487 -505 1487 -505 0 feedthrough
rlabel pdiffusion 1494 -505 1494 -505 0 feedthrough
rlabel pdiffusion 1501 -505 1501 -505 0 feedthrough
rlabel pdiffusion 1508 -505 1508 -505 0 feedthrough
rlabel pdiffusion 1515 -505 1515 -505 0 feedthrough
rlabel pdiffusion 1522 -505 1522 -505 0 feedthrough
rlabel pdiffusion 1529 -505 1529 -505 0 feedthrough
rlabel pdiffusion 1536 -505 1536 -505 0 feedthrough
rlabel pdiffusion 1543 -505 1543 -505 0 feedthrough
rlabel pdiffusion 1550 -505 1550 -505 0 feedthrough
rlabel pdiffusion 1557 -505 1557 -505 0 feedthrough
rlabel pdiffusion 1564 -505 1564 -505 0 feedthrough
rlabel pdiffusion 1571 -505 1571 -505 0 feedthrough
rlabel pdiffusion 1578 -505 1578 -505 0 feedthrough
rlabel pdiffusion 1585 -505 1585 -505 0 feedthrough
rlabel pdiffusion 1592 -505 1592 -505 0 feedthrough
rlabel pdiffusion 1599 -505 1599 -505 0 feedthrough
rlabel pdiffusion 1606 -505 1606 -505 0 feedthrough
rlabel pdiffusion 1613 -505 1613 -505 0 feedthrough
rlabel pdiffusion 1620 -505 1620 -505 0 feedthrough
rlabel pdiffusion 1627 -505 1627 -505 0 feedthrough
rlabel pdiffusion 1634 -505 1634 -505 0 feedthrough
rlabel pdiffusion 1641 -505 1641 -505 0 feedthrough
rlabel pdiffusion 1648 -505 1648 -505 0 feedthrough
rlabel pdiffusion 1655 -505 1655 -505 0 feedthrough
rlabel pdiffusion 1662 -505 1662 -505 0 feedthrough
rlabel pdiffusion 1669 -505 1669 -505 0 feedthrough
rlabel pdiffusion 1676 -505 1676 -505 0 feedthrough
rlabel pdiffusion 1683 -505 1683 -505 0 feedthrough
rlabel pdiffusion 1690 -505 1690 -505 0 feedthrough
rlabel pdiffusion 1697 -505 1697 -505 0 feedthrough
rlabel pdiffusion 1704 -505 1704 -505 0 feedthrough
rlabel pdiffusion 1711 -505 1711 -505 0 feedthrough
rlabel pdiffusion 1718 -505 1718 -505 0 feedthrough
rlabel pdiffusion 1725 -505 1725 -505 0 feedthrough
rlabel pdiffusion 1732 -505 1732 -505 0 feedthrough
rlabel pdiffusion 1739 -505 1739 -505 0 feedthrough
rlabel pdiffusion 1746 -505 1746 -505 0 feedthrough
rlabel pdiffusion 1753 -505 1753 -505 0 feedthrough
rlabel pdiffusion 1760 -505 1760 -505 0 feedthrough
rlabel pdiffusion 1767 -505 1767 -505 0 feedthrough
rlabel pdiffusion 1774 -505 1774 -505 0 feedthrough
rlabel pdiffusion 1781 -505 1781 -505 0 feedthrough
rlabel pdiffusion 1788 -505 1788 -505 0 feedthrough
rlabel pdiffusion 1795 -505 1795 -505 0 feedthrough
rlabel pdiffusion 1802 -505 1802 -505 0 feedthrough
rlabel pdiffusion 1809 -505 1809 -505 0 feedthrough
rlabel pdiffusion 1816 -505 1816 -505 0 feedthrough
rlabel pdiffusion 1823 -505 1823 -505 0 feedthrough
rlabel pdiffusion 1830 -505 1830 -505 0 feedthrough
rlabel pdiffusion 1837 -505 1837 -505 0 feedthrough
rlabel pdiffusion 1844 -505 1844 -505 0 feedthrough
rlabel pdiffusion 1851 -505 1851 -505 0 feedthrough
rlabel pdiffusion 1858 -505 1858 -505 0 feedthrough
rlabel pdiffusion 1865 -505 1865 -505 0 feedthrough
rlabel pdiffusion 1872 -505 1872 -505 0 feedthrough
rlabel pdiffusion 1879 -505 1879 -505 0 feedthrough
rlabel pdiffusion 1886 -505 1886 -505 0 feedthrough
rlabel pdiffusion 1893 -505 1893 -505 0 feedthrough
rlabel pdiffusion 1900 -505 1900 -505 0 feedthrough
rlabel pdiffusion 1907 -505 1907 -505 0 feedthrough
rlabel pdiffusion 1914 -505 1914 -505 0 feedthrough
rlabel pdiffusion 1921 -505 1921 -505 0 feedthrough
rlabel pdiffusion 1928 -505 1928 -505 0 feedthrough
rlabel pdiffusion 1935 -505 1935 -505 0 feedthrough
rlabel pdiffusion 1942 -505 1942 -505 0 feedthrough
rlabel pdiffusion 1949 -505 1949 -505 0 feedthrough
rlabel pdiffusion 1956 -505 1956 -505 0 cellNo=259
rlabel pdiffusion 1963 -505 1963 -505 0 feedthrough
rlabel pdiffusion 1970 -505 1970 -505 0 feedthrough
rlabel pdiffusion 1977 -505 1977 -505 0 cellNo=305
rlabel pdiffusion 1984 -505 1984 -505 0 feedthrough
rlabel pdiffusion 1991 -505 1991 -505 0 feedthrough
rlabel pdiffusion 1998 -505 1998 -505 0 feedthrough
rlabel pdiffusion 2005 -505 2005 -505 0 cellNo=435
rlabel pdiffusion 2012 -505 2012 -505 0 cellNo=685
rlabel pdiffusion 2019 -505 2019 -505 0 cellNo=912
rlabel pdiffusion 2040 -505 2040 -505 0 feedthrough
rlabel pdiffusion 2089 -505 2089 -505 0 feedthrough
rlabel pdiffusion 2117 -505 2117 -505 0 feedthrough
rlabel pdiffusion 2145 -505 2145 -505 0 feedthrough
rlabel pdiffusion 2264 -505 2264 -505 0 feedthrough
rlabel pdiffusion 2285 -505 2285 -505 0 feedthrough
rlabel pdiffusion 3 -638 3 -638 0 cellNo=677
rlabel pdiffusion 10 -638 10 -638 0 feedthrough
rlabel pdiffusion 17 -638 17 -638 0 feedthrough
rlabel pdiffusion 24 -638 24 -638 0 feedthrough
rlabel pdiffusion 31 -638 31 -638 0 feedthrough
rlabel pdiffusion 38 -638 38 -638 0 feedthrough
rlabel pdiffusion 45 -638 45 -638 0 feedthrough
rlabel pdiffusion 52 -638 52 -638 0 feedthrough
rlabel pdiffusion 59 -638 59 -638 0 cellNo=860
rlabel pdiffusion 66 -638 66 -638 0 feedthrough
rlabel pdiffusion 73 -638 73 -638 0 cellNo=952
rlabel pdiffusion 80 -638 80 -638 0 feedthrough
rlabel pdiffusion 87 -638 87 -638 0 feedthrough
rlabel pdiffusion 94 -638 94 -638 0 feedthrough
rlabel pdiffusion 101 -638 101 -638 0 cellNo=373
rlabel pdiffusion 108 -638 108 -638 0 feedthrough
rlabel pdiffusion 115 -638 115 -638 0 feedthrough
rlabel pdiffusion 122 -638 122 -638 0 feedthrough
rlabel pdiffusion 129 -638 129 -638 0 feedthrough
rlabel pdiffusion 136 -638 136 -638 0 cellNo=241
rlabel pdiffusion 143 -638 143 -638 0 feedthrough
rlabel pdiffusion 150 -638 150 -638 0 feedthrough
rlabel pdiffusion 157 -638 157 -638 0 feedthrough
rlabel pdiffusion 164 -638 164 -638 0 feedthrough
rlabel pdiffusion 171 -638 171 -638 0 cellNo=713
rlabel pdiffusion 178 -638 178 -638 0 feedthrough
rlabel pdiffusion 185 -638 185 -638 0 feedthrough
rlabel pdiffusion 192 -638 192 -638 0 feedthrough
rlabel pdiffusion 199 -638 199 -638 0 feedthrough
rlabel pdiffusion 206 -638 206 -638 0 cellNo=283
rlabel pdiffusion 213 -638 213 -638 0 feedthrough
rlabel pdiffusion 220 -638 220 -638 0 feedthrough
rlabel pdiffusion 227 -638 227 -638 0 feedthrough
rlabel pdiffusion 234 -638 234 -638 0 feedthrough
rlabel pdiffusion 241 -638 241 -638 0 feedthrough
rlabel pdiffusion 248 -638 248 -638 0 cellNo=738
rlabel pdiffusion 255 -638 255 -638 0 feedthrough
rlabel pdiffusion 262 -638 262 -638 0 feedthrough
rlabel pdiffusion 269 -638 269 -638 0 cellNo=209
rlabel pdiffusion 276 -638 276 -638 0 feedthrough
rlabel pdiffusion 283 -638 283 -638 0 feedthrough
rlabel pdiffusion 290 -638 290 -638 0 feedthrough
rlabel pdiffusion 297 -638 297 -638 0 feedthrough
rlabel pdiffusion 304 -638 304 -638 0 feedthrough
rlabel pdiffusion 311 -638 311 -638 0 feedthrough
rlabel pdiffusion 318 -638 318 -638 0 feedthrough
rlabel pdiffusion 325 -638 325 -638 0 feedthrough
rlabel pdiffusion 332 -638 332 -638 0 feedthrough
rlabel pdiffusion 339 -638 339 -638 0 feedthrough
rlabel pdiffusion 346 -638 346 -638 0 feedthrough
rlabel pdiffusion 353 -638 353 -638 0 feedthrough
rlabel pdiffusion 360 -638 360 -638 0 feedthrough
rlabel pdiffusion 367 -638 367 -638 0 feedthrough
rlabel pdiffusion 374 -638 374 -638 0 feedthrough
rlabel pdiffusion 381 -638 381 -638 0 feedthrough
rlabel pdiffusion 388 -638 388 -638 0 feedthrough
rlabel pdiffusion 395 -638 395 -638 0 feedthrough
rlabel pdiffusion 402 -638 402 -638 0 feedthrough
rlabel pdiffusion 409 -638 409 -638 0 feedthrough
rlabel pdiffusion 416 -638 416 -638 0 feedthrough
rlabel pdiffusion 423 -638 423 -638 0 feedthrough
rlabel pdiffusion 430 -638 430 -638 0 cellNo=754
rlabel pdiffusion 437 -638 437 -638 0 feedthrough
rlabel pdiffusion 444 -638 444 -638 0 feedthrough
rlabel pdiffusion 451 -638 451 -638 0 feedthrough
rlabel pdiffusion 458 -638 458 -638 0 feedthrough
rlabel pdiffusion 465 -638 465 -638 0 feedthrough
rlabel pdiffusion 472 -638 472 -638 0 feedthrough
rlabel pdiffusion 479 -638 479 -638 0 feedthrough
rlabel pdiffusion 486 -638 486 -638 0 feedthrough
rlabel pdiffusion 493 -638 493 -638 0 feedthrough
rlabel pdiffusion 500 -638 500 -638 0 feedthrough
rlabel pdiffusion 507 -638 507 -638 0 feedthrough
rlabel pdiffusion 514 -638 514 -638 0 feedthrough
rlabel pdiffusion 521 -638 521 -638 0 feedthrough
rlabel pdiffusion 528 -638 528 -638 0 feedthrough
rlabel pdiffusion 535 -638 535 -638 0 cellNo=573
rlabel pdiffusion 542 -638 542 -638 0 feedthrough
rlabel pdiffusion 549 -638 549 -638 0 feedthrough
rlabel pdiffusion 556 -638 556 -638 0 feedthrough
rlabel pdiffusion 563 -638 563 -638 0 cellNo=406
rlabel pdiffusion 570 -638 570 -638 0 feedthrough
rlabel pdiffusion 577 -638 577 -638 0 feedthrough
rlabel pdiffusion 584 -638 584 -638 0 cellNo=74
rlabel pdiffusion 591 -638 591 -638 0 cellNo=117
rlabel pdiffusion 598 -638 598 -638 0 feedthrough
rlabel pdiffusion 605 -638 605 -638 0 feedthrough
rlabel pdiffusion 612 -638 612 -638 0 feedthrough
rlabel pdiffusion 619 -638 619 -638 0 feedthrough
rlabel pdiffusion 626 -638 626 -638 0 feedthrough
rlabel pdiffusion 633 -638 633 -638 0 feedthrough
rlabel pdiffusion 640 -638 640 -638 0 feedthrough
rlabel pdiffusion 647 -638 647 -638 0 cellNo=579
rlabel pdiffusion 654 -638 654 -638 0 feedthrough
rlabel pdiffusion 661 -638 661 -638 0 cellNo=355
rlabel pdiffusion 668 -638 668 -638 0 feedthrough
rlabel pdiffusion 675 -638 675 -638 0 feedthrough
rlabel pdiffusion 682 -638 682 -638 0 feedthrough
rlabel pdiffusion 689 -638 689 -638 0 feedthrough
rlabel pdiffusion 696 -638 696 -638 0 feedthrough
rlabel pdiffusion 703 -638 703 -638 0 feedthrough
rlabel pdiffusion 710 -638 710 -638 0 feedthrough
rlabel pdiffusion 717 -638 717 -638 0 feedthrough
rlabel pdiffusion 724 -638 724 -638 0 feedthrough
rlabel pdiffusion 731 -638 731 -638 0 cellNo=687
rlabel pdiffusion 738 -638 738 -638 0 feedthrough
rlabel pdiffusion 745 -638 745 -638 0 cellNo=13
rlabel pdiffusion 752 -638 752 -638 0 feedthrough
rlabel pdiffusion 759 -638 759 -638 0 feedthrough
rlabel pdiffusion 766 -638 766 -638 0 feedthrough
rlabel pdiffusion 773 -638 773 -638 0 feedthrough
rlabel pdiffusion 780 -638 780 -638 0 feedthrough
rlabel pdiffusion 787 -638 787 -638 0 cellNo=116
rlabel pdiffusion 794 -638 794 -638 0 feedthrough
rlabel pdiffusion 801 -638 801 -638 0 feedthrough
rlabel pdiffusion 808 -638 808 -638 0 cellNo=158
rlabel pdiffusion 815 -638 815 -638 0 feedthrough
rlabel pdiffusion 822 -638 822 -638 0 cellNo=186
rlabel pdiffusion 829 -638 829 -638 0 feedthrough
rlabel pdiffusion 836 -638 836 -638 0 feedthrough
rlabel pdiffusion 843 -638 843 -638 0 feedthrough
rlabel pdiffusion 850 -638 850 -638 0 cellNo=138
rlabel pdiffusion 857 -638 857 -638 0 feedthrough
rlabel pdiffusion 864 -638 864 -638 0 feedthrough
rlabel pdiffusion 871 -638 871 -638 0 feedthrough
rlabel pdiffusion 878 -638 878 -638 0 feedthrough
rlabel pdiffusion 885 -638 885 -638 0 feedthrough
rlabel pdiffusion 892 -638 892 -638 0 feedthrough
rlabel pdiffusion 899 -638 899 -638 0 feedthrough
rlabel pdiffusion 906 -638 906 -638 0 feedthrough
rlabel pdiffusion 913 -638 913 -638 0 feedthrough
rlabel pdiffusion 920 -638 920 -638 0 feedthrough
rlabel pdiffusion 927 -638 927 -638 0 cellNo=692
rlabel pdiffusion 934 -638 934 -638 0 feedthrough
rlabel pdiffusion 941 -638 941 -638 0 cellNo=841
rlabel pdiffusion 948 -638 948 -638 0 feedthrough
rlabel pdiffusion 955 -638 955 -638 0 feedthrough
rlabel pdiffusion 962 -638 962 -638 0 feedthrough
rlabel pdiffusion 969 -638 969 -638 0 feedthrough
rlabel pdiffusion 976 -638 976 -638 0 feedthrough
rlabel pdiffusion 983 -638 983 -638 0 cellNo=71
rlabel pdiffusion 990 -638 990 -638 0 feedthrough
rlabel pdiffusion 997 -638 997 -638 0 feedthrough
rlabel pdiffusion 1004 -638 1004 -638 0 feedthrough
rlabel pdiffusion 1011 -638 1011 -638 0 cellNo=554
rlabel pdiffusion 1018 -638 1018 -638 0 feedthrough
rlabel pdiffusion 1025 -638 1025 -638 0 feedthrough
rlabel pdiffusion 1032 -638 1032 -638 0 cellNo=566
rlabel pdiffusion 1039 -638 1039 -638 0 feedthrough
rlabel pdiffusion 1046 -638 1046 -638 0 feedthrough
rlabel pdiffusion 1053 -638 1053 -638 0 feedthrough
rlabel pdiffusion 1060 -638 1060 -638 0 cellNo=54
rlabel pdiffusion 1067 -638 1067 -638 0 feedthrough
rlabel pdiffusion 1074 -638 1074 -638 0 feedthrough
rlabel pdiffusion 1081 -638 1081 -638 0 cellNo=43
rlabel pdiffusion 1088 -638 1088 -638 0 feedthrough
rlabel pdiffusion 1095 -638 1095 -638 0 cellNo=445
rlabel pdiffusion 1102 -638 1102 -638 0 feedthrough
rlabel pdiffusion 1109 -638 1109 -638 0 feedthrough
rlabel pdiffusion 1116 -638 1116 -638 0 feedthrough
rlabel pdiffusion 1123 -638 1123 -638 0 feedthrough
rlabel pdiffusion 1130 -638 1130 -638 0 feedthrough
rlabel pdiffusion 1137 -638 1137 -638 0 feedthrough
rlabel pdiffusion 1144 -638 1144 -638 0 cellNo=83
rlabel pdiffusion 1151 -638 1151 -638 0 cellNo=611
rlabel pdiffusion 1158 -638 1158 -638 0 feedthrough
rlabel pdiffusion 1165 -638 1165 -638 0 feedthrough
rlabel pdiffusion 1172 -638 1172 -638 0 feedthrough
rlabel pdiffusion 1179 -638 1179 -638 0 feedthrough
rlabel pdiffusion 1186 -638 1186 -638 0 feedthrough
rlabel pdiffusion 1193 -638 1193 -638 0 feedthrough
rlabel pdiffusion 1200 -638 1200 -638 0 cellNo=401
rlabel pdiffusion 1207 -638 1207 -638 0 feedthrough
rlabel pdiffusion 1214 -638 1214 -638 0 cellNo=63
rlabel pdiffusion 1221 -638 1221 -638 0 feedthrough
rlabel pdiffusion 1228 -638 1228 -638 0 feedthrough
rlabel pdiffusion 1235 -638 1235 -638 0 feedthrough
rlabel pdiffusion 1242 -638 1242 -638 0 feedthrough
rlabel pdiffusion 1249 -638 1249 -638 0 feedthrough
rlabel pdiffusion 1256 -638 1256 -638 0 feedthrough
rlabel pdiffusion 1263 -638 1263 -638 0 feedthrough
rlabel pdiffusion 1270 -638 1270 -638 0 feedthrough
rlabel pdiffusion 1277 -638 1277 -638 0 feedthrough
rlabel pdiffusion 1284 -638 1284 -638 0 feedthrough
rlabel pdiffusion 1291 -638 1291 -638 0 feedthrough
rlabel pdiffusion 1298 -638 1298 -638 0 cellNo=179
rlabel pdiffusion 1305 -638 1305 -638 0 feedthrough
rlabel pdiffusion 1312 -638 1312 -638 0 feedthrough
rlabel pdiffusion 1319 -638 1319 -638 0 feedthrough
rlabel pdiffusion 1326 -638 1326 -638 0 feedthrough
rlabel pdiffusion 1333 -638 1333 -638 0 feedthrough
rlabel pdiffusion 1340 -638 1340 -638 0 feedthrough
rlabel pdiffusion 1347 -638 1347 -638 0 feedthrough
rlabel pdiffusion 1354 -638 1354 -638 0 feedthrough
rlabel pdiffusion 1361 -638 1361 -638 0 feedthrough
rlabel pdiffusion 1368 -638 1368 -638 0 feedthrough
rlabel pdiffusion 1375 -638 1375 -638 0 feedthrough
rlabel pdiffusion 1382 -638 1382 -638 0 feedthrough
rlabel pdiffusion 1389 -638 1389 -638 0 feedthrough
rlabel pdiffusion 1396 -638 1396 -638 0 feedthrough
rlabel pdiffusion 1403 -638 1403 -638 0 feedthrough
rlabel pdiffusion 1410 -638 1410 -638 0 feedthrough
rlabel pdiffusion 1417 -638 1417 -638 0 feedthrough
rlabel pdiffusion 1424 -638 1424 -638 0 feedthrough
rlabel pdiffusion 1431 -638 1431 -638 0 feedthrough
rlabel pdiffusion 1438 -638 1438 -638 0 feedthrough
rlabel pdiffusion 1445 -638 1445 -638 0 feedthrough
rlabel pdiffusion 1452 -638 1452 -638 0 feedthrough
rlabel pdiffusion 1459 -638 1459 -638 0 feedthrough
rlabel pdiffusion 1466 -638 1466 -638 0 feedthrough
rlabel pdiffusion 1473 -638 1473 -638 0 feedthrough
rlabel pdiffusion 1480 -638 1480 -638 0 feedthrough
rlabel pdiffusion 1487 -638 1487 -638 0 cellNo=92
rlabel pdiffusion 1494 -638 1494 -638 0 feedthrough
rlabel pdiffusion 1501 -638 1501 -638 0 feedthrough
rlabel pdiffusion 1508 -638 1508 -638 0 feedthrough
rlabel pdiffusion 1515 -638 1515 -638 0 feedthrough
rlabel pdiffusion 1522 -638 1522 -638 0 feedthrough
rlabel pdiffusion 1529 -638 1529 -638 0 feedthrough
rlabel pdiffusion 1536 -638 1536 -638 0 feedthrough
rlabel pdiffusion 1543 -638 1543 -638 0 feedthrough
rlabel pdiffusion 1550 -638 1550 -638 0 feedthrough
rlabel pdiffusion 1557 -638 1557 -638 0 feedthrough
rlabel pdiffusion 1564 -638 1564 -638 0 feedthrough
rlabel pdiffusion 1571 -638 1571 -638 0 feedthrough
rlabel pdiffusion 1578 -638 1578 -638 0 feedthrough
rlabel pdiffusion 1585 -638 1585 -638 0 feedthrough
rlabel pdiffusion 1592 -638 1592 -638 0 feedthrough
rlabel pdiffusion 1599 -638 1599 -638 0 feedthrough
rlabel pdiffusion 1606 -638 1606 -638 0 feedthrough
rlabel pdiffusion 1613 -638 1613 -638 0 feedthrough
rlabel pdiffusion 1620 -638 1620 -638 0 feedthrough
rlabel pdiffusion 1627 -638 1627 -638 0 feedthrough
rlabel pdiffusion 1634 -638 1634 -638 0 feedthrough
rlabel pdiffusion 1641 -638 1641 -638 0 feedthrough
rlabel pdiffusion 1648 -638 1648 -638 0 feedthrough
rlabel pdiffusion 1655 -638 1655 -638 0 feedthrough
rlabel pdiffusion 1662 -638 1662 -638 0 feedthrough
rlabel pdiffusion 1669 -638 1669 -638 0 feedthrough
rlabel pdiffusion 1676 -638 1676 -638 0 feedthrough
rlabel pdiffusion 1683 -638 1683 -638 0 feedthrough
rlabel pdiffusion 1690 -638 1690 -638 0 feedthrough
rlabel pdiffusion 1697 -638 1697 -638 0 feedthrough
rlabel pdiffusion 1704 -638 1704 -638 0 feedthrough
rlabel pdiffusion 1711 -638 1711 -638 0 feedthrough
rlabel pdiffusion 1718 -638 1718 -638 0 feedthrough
rlabel pdiffusion 1725 -638 1725 -638 0 feedthrough
rlabel pdiffusion 1732 -638 1732 -638 0 feedthrough
rlabel pdiffusion 1739 -638 1739 -638 0 feedthrough
rlabel pdiffusion 1746 -638 1746 -638 0 feedthrough
rlabel pdiffusion 1753 -638 1753 -638 0 feedthrough
rlabel pdiffusion 1760 -638 1760 -638 0 feedthrough
rlabel pdiffusion 1767 -638 1767 -638 0 feedthrough
rlabel pdiffusion 1774 -638 1774 -638 0 feedthrough
rlabel pdiffusion 1781 -638 1781 -638 0 feedthrough
rlabel pdiffusion 1788 -638 1788 -638 0 feedthrough
rlabel pdiffusion 1795 -638 1795 -638 0 feedthrough
rlabel pdiffusion 1802 -638 1802 -638 0 feedthrough
rlabel pdiffusion 1809 -638 1809 -638 0 feedthrough
rlabel pdiffusion 1816 -638 1816 -638 0 feedthrough
rlabel pdiffusion 1823 -638 1823 -638 0 feedthrough
rlabel pdiffusion 1830 -638 1830 -638 0 feedthrough
rlabel pdiffusion 1837 -638 1837 -638 0 feedthrough
rlabel pdiffusion 1844 -638 1844 -638 0 feedthrough
rlabel pdiffusion 1851 -638 1851 -638 0 feedthrough
rlabel pdiffusion 1858 -638 1858 -638 0 feedthrough
rlabel pdiffusion 1865 -638 1865 -638 0 feedthrough
rlabel pdiffusion 1872 -638 1872 -638 0 feedthrough
rlabel pdiffusion 1879 -638 1879 -638 0 feedthrough
rlabel pdiffusion 1886 -638 1886 -638 0 feedthrough
rlabel pdiffusion 1893 -638 1893 -638 0 feedthrough
rlabel pdiffusion 1900 -638 1900 -638 0 feedthrough
rlabel pdiffusion 1907 -638 1907 -638 0 feedthrough
rlabel pdiffusion 1914 -638 1914 -638 0 feedthrough
rlabel pdiffusion 1921 -638 1921 -638 0 feedthrough
rlabel pdiffusion 1928 -638 1928 -638 0 feedthrough
rlabel pdiffusion 1935 -638 1935 -638 0 feedthrough
rlabel pdiffusion 1942 -638 1942 -638 0 feedthrough
rlabel pdiffusion 1949 -638 1949 -638 0 feedthrough
rlabel pdiffusion 1956 -638 1956 -638 0 feedthrough
rlabel pdiffusion 1963 -638 1963 -638 0 feedthrough
rlabel pdiffusion 1970 -638 1970 -638 0 feedthrough
rlabel pdiffusion 1977 -638 1977 -638 0 feedthrough
rlabel pdiffusion 1984 -638 1984 -638 0 feedthrough
rlabel pdiffusion 1991 -638 1991 -638 0 feedthrough
rlabel pdiffusion 1998 -638 1998 -638 0 feedthrough
rlabel pdiffusion 2005 -638 2005 -638 0 feedthrough
rlabel pdiffusion 2012 -638 2012 -638 0 feedthrough
rlabel pdiffusion 2019 -638 2019 -638 0 feedthrough
rlabel pdiffusion 2026 -638 2026 -638 0 feedthrough
rlabel pdiffusion 2033 -638 2033 -638 0 feedthrough
rlabel pdiffusion 2040 -638 2040 -638 0 feedthrough
rlabel pdiffusion 2047 -638 2047 -638 0 feedthrough
rlabel pdiffusion 2054 -638 2054 -638 0 feedthrough
rlabel pdiffusion 2061 -638 2061 -638 0 feedthrough
rlabel pdiffusion 2068 -638 2068 -638 0 feedthrough
rlabel pdiffusion 2075 -638 2075 -638 0 feedthrough
rlabel pdiffusion 2082 -638 2082 -638 0 feedthrough
rlabel pdiffusion 2089 -638 2089 -638 0 feedthrough
rlabel pdiffusion 2096 -638 2096 -638 0 feedthrough
rlabel pdiffusion 2103 -638 2103 -638 0 feedthrough
rlabel pdiffusion 2110 -638 2110 -638 0 feedthrough
rlabel pdiffusion 2117 -638 2117 -638 0 feedthrough
rlabel pdiffusion 2124 -638 2124 -638 0 feedthrough
rlabel pdiffusion 2131 -638 2131 -638 0 feedthrough
rlabel pdiffusion 2138 -638 2138 -638 0 feedthrough
rlabel pdiffusion 2145 -638 2145 -638 0 feedthrough
rlabel pdiffusion 2152 -638 2152 -638 0 feedthrough
rlabel pdiffusion 2159 -638 2159 -638 0 feedthrough
rlabel pdiffusion 2166 -638 2166 -638 0 feedthrough
rlabel pdiffusion 2173 -638 2173 -638 0 feedthrough
rlabel pdiffusion 2180 -638 2180 -638 0 feedthrough
rlabel pdiffusion 2187 -638 2187 -638 0 feedthrough
rlabel pdiffusion 2194 -638 2194 -638 0 feedthrough
rlabel pdiffusion 2201 -638 2201 -638 0 feedthrough
rlabel pdiffusion 2208 -638 2208 -638 0 cellNo=339
rlabel pdiffusion 2215 -638 2215 -638 0 cellNo=151
rlabel pdiffusion 2222 -638 2222 -638 0 cellNo=344
rlabel pdiffusion 2292 -638 2292 -638 0 feedthrough
rlabel pdiffusion 2327 -638 2327 -638 0 feedthrough
rlabel pdiffusion 2362 -638 2362 -638 0 feedthrough
rlabel pdiffusion 3 -815 3 -815 0 feedthrough
rlabel pdiffusion 10 -815 10 -815 0 cellNo=821
rlabel pdiffusion 17 -815 17 -815 0 cellNo=947
rlabel pdiffusion 24 -815 24 -815 0 feedthrough
rlabel pdiffusion 31 -815 31 -815 0 feedthrough
rlabel pdiffusion 38 -815 38 -815 0 feedthrough
rlabel pdiffusion 45 -815 45 -815 0 cellNo=527
rlabel pdiffusion 52 -815 52 -815 0 feedthrough
rlabel pdiffusion 59 -815 59 -815 0 feedthrough
rlabel pdiffusion 66 -815 66 -815 0 cellNo=370
rlabel pdiffusion 73 -815 73 -815 0 feedthrough
rlabel pdiffusion 80 -815 80 -815 0 cellNo=307
rlabel pdiffusion 87 -815 87 -815 0 feedthrough
rlabel pdiffusion 94 -815 94 -815 0 feedthrough
rlabel pdiffusion 101 -815 101 -815 0 feedthrough
rlabel pdiffusion 108 -815 108 -815 0 feedthrough
rlabel pdiffusion 115 -815 115 -815 0 feedthrough
rlabel pdiffusion 122 -815 122 -815 0 cellNo=87
rlabel pdiffusion 129 -815 129 -815 0 cellNo=153
rlabel pdiffusion 136 -815 136 -815 0 feedthrough
rlabel pdiffusion 143 -815 143 -815 0 cellNo=225
rlabel pdiffusion 150 -815 150 -815 0 feedthrough
rlabel pdiffusion 157 -815 157 -815 0 feedthrough
rlabel pdiffusion 164 -815 164 -815 0 feedthrough
rlabel pdiffusion 171 -815 171 -815 0 feedthrough
rlabel pdiffusion 178 -815 178 -815 0 feedthrough
rlabel pdiffusion 185 -815 185 -815 0 cellNo=904
rlabel pdiffusion 192 -815 192 -815 0 feedthrough
rlabel pdiffusion 199 -815 199 -815 0 feedthrough
rlabel pdiffusion 206 -815 206 -815 0 cellNo=286
rlabel pdiffusion 213 -815 213 -815 0 feedthrough
rlabel pdiffusion 220 -815 220 -815 0 cellNo=656
rlabel pdiffusion 227 -815 227 -815 0 feedthrough
rlabel pdiffusion 234 -815 234 -815 0 cellNo=839
rlabel pdiffusion 241 -815 241 -815 0 feedthrough
rlabel pdiffusion 248 -815 248 -815 0 feedthrough
rlabel pdiffusion 255 -815 255 -815 0 feedthrough
rlabel pdiffusion 262 -815 262 -815 0 feedthrough
rlabel pdiffusion 269 -815 269 -815 0 feedthrough
rlabel pdiffusion 276 -815 276 -815 0 feedthrough
rlabel pdiffusion 283 -815 283 -815 0 feedthrough
rlabel pdiffusion 290 -815 290 -815 0 feedthrough
rlabel pdiffusion 297 -815 297 -815 0 feedthrough
rlabel pdiffusion 304 -815 304 -815 0 feedthrough
rlabel pdiffusion 311 -815 311 -815 0 feedthrough
rlabel pdiffusion 318 -815 318 -815 0 feedthrough
rlabel pdiffusion 325 -815 325 -815 0 feedthrough
rlabel pdiffusion 332 -815 332 -815 0 feedthrough
rlabel pdiffusion 339 -815 339 -815 0 feedthrough
rlabel pdiffusion 346 -815 346 -815 0 feedthrough
rlabel pdiffusion 353 -815 353 -815 0 feedthrough
rlabel pdiffusion 360 -815 360 -815 0 cellNo=1
rlabel pdiffusion 367 -815 367 -815 0 feedthrough
rlabel pdiffusion 374 -815 374 -815 0 feedthrough
rlabel pdiffusion 381 -815 381 -815 0 feedthrough
rlabel pdiffusion 388 -815 388 -815 0 feedthrough
rlabel pdiffusion 395 -815 395 -815 0 feedthrough
rlabel pdiffusion 402 -815 402 -815 0 feedthrough
rlabel pdiffusion 409 -815 409 -815 0 feedthrough
rlabel pdiffusion 416 -815 416 -815 0 feedthrough
rlabel pdiffusion 423 -815 423 -815 0 feedthrough
rlabel pdiffusion 430 -815 430 -815 0 feedthrough
rlabel pdiffusion 437 -815 437 -815 0 feedthrough
rlabel pdiffusion 444 -815 444 -815 0 feedthrough
rlabel pdiffusion 451 -815 451 -815 0 feedthrough
rlabel pdiffusion 458 -815 458 -815 0 feedthrough
rlabel pdiffusion 465 -815 465 -815 0 feedthrough
rlabel pdiffusion 472 -815 472 -815 0 feedthrough
rlabel pdiffusion 479 -815 479 -815 0 feedthrough
rlabel pdiffusion 486 -815 486 -815 0 feedthrough
rlabel pdiffusion 493 -815 493 -815 0 feedthrough
rlabel pdiffusion 500 -815 500 -815 0 feedthrough
rlabel pdiffusion 507 -815 507 -815 0 feedthrough
rlabel pdiffusion 514 -815 514 -815 0 feedthrough
rlabel pdiffusion 521 -815 521 -815 0 cellNo=898
rlabel pdiffusion 528 -815 528 -815 0 feedthrough
rlabel pdiffusion 535 -815 535 -815 0 feedthrough
rlabel pdiffusion 542 -815 542 -815 0 feedthrough
rlabel pdiffusion 549 -815 549 -815 0 feedthrough
rlabel pdiffusion 556 -815 556 -815 0 feedthrough
rlabel pdiffusion 563 -815 563 -815 0 feedthrough
rlabel pdiffusion 570 -815 570 -815 0 feedthrough
rlabel pdiffusion 577 -815 577 -815 0 feedthrough
rlabel pdiffusion 584 -815 584 -815 0 cellNo=366
rlabel pdiffusion 591 -815 591 -815 0 cellNo=199
rlabel pdiffusion 598 -815 598 -815 0 feedthrough
rlabel pdiffusion 605 -815 605 -815 0 feedthrough
rlabel pdiffusion 612 -815 612 -815 0 feedthrough
rlabel pdiffusion 619 -815 619 -815 0 feedthrough
rlabel pdiffusion 626 -815 626 -815 0 feedthrough
rlabel pdiffusion 633 -815 633 -815 0 feedthrough
rlabel pdiffusion 640 -815 640 -815 0 feedthrough
rlabel pdiffusion 647 -815 647 -815 0 feedthrough
rlabel pdiffusion 654 -815 654 -815 0 feedthrough
rlabel pdiffusion 661 -815 661 -815 0 feedthrough
rlabel pdiffusion 668 -815 668 -815 0 feedthrough
rlabel pdiffusion 675 -815 675 -815 0 feedthrough
rlabel pdiffusion 682 -815 682 -815 0 cellNo=522
rlabel pdiffusion 689 -815 689 -815 0 feedthrough
rlabel pdiffusion 696 -815 696 -815 0 cellNo=858
rlabel pdiffusion 703 -815 703 -815 0 feedthrough
rlabel pdiffusion 710 -815 710 -815 0 feedthrough
rlabel pdiffusion 717 -815 717 -815 0 feedthrough
rlabel pdiffusion 724 -815 724 -815 0 cellNo=107
rlabel pdiffusion 731 -815 731 -815 0 feedthrough
rlabel pdiffusion 738 -815 738 -815 0 feedthrough
rlabel pdiffusion 745 -815 745 -815 0 cellNo=541
rlabel pdiffusion 752 -815 752 -815 0 cellNo=817
rlabel pdiffusion 759 -815 759 -815 0 feedthrough
rlabel pdiffusion 766 -815 766 -815 0 feedthrough
rlabel pdiffusion 773 -815 773 -815 0 feedthrough
rlabel pdiffusion 780 -815 780 -815 0 feedthrough
rlabel pdiffusion 787 -815 787 -815 0 feedthrough
rlabel pdiffusion 794 -815 794 -815 0 feedthrough
rlabel pdiffusion 801 -815 801 -815 0 feedthrough
rlabel pdiffusion 808 -815 808 -815 0 feedthrough
rlabel pdiffusion 815 -815 815 -815 0 feedthrough
rlabel pdiffusion 822 -815 822 -815 0 feedthrough
rlabel pdiffusion 829 -815 829 -815 0 cellNo=273
rlabel pdiffusion 836 -815 836 -815 0 feedthrough
rlabel pdiffusion 843 -815 843 -815 0 feedthrough
rlabel pdiffusion 850 -815 850 -815 0 feedthrough
rlabel pdiffusion 857 -815 857 -815 0 feedthrough
rlabel pdiffusion 864 -815 864 -815 0 feedthrough
rlabel pdiffusion 871 -815 871 -815 0 feedthrough
rlabel pdiffusion 878 -815 878 -815 0 cellNo=752
rlabel pdiffusion 885 -815 885 -815 0 feedthrough
rlabel pdiffusion 892 -815 892 -815 0 feedthrough
rlabel pdiffusion 899 -815 899 -815 0 feedthrough
rlabel pdiffusion 906 -815 906 -815 0 feedthrough
rlabel pdiffusion 913 -815 913 -815 0 feedthrough
rlabel pdiffusion 920 -815 920 -815 0 feedthrough
rlabel pdiffusion 927 -815 927 -815 0 feedthrough
rlabel pdiffusion 934 -815 934 -815 0 feedthrough
rlabel pdiffusion 941 -815 941 -815 0 feedthrough
rlabel pdiffusion 948 -815 948 -815 0 feedthrough
rlabel pdiffusion 955 -815 955 -815 0 cellNo=295
rlabel pdiffusion 962 -815 962 -815 0 feedthrough
rlabel pdiffusion 969 -815 969 -815 0 feedthrough
rlabel pdiffusion 976 -815 976 -815 0 feedthrough
rlabel pdiffusion 983 -815 983 -815 0 feedthrough
rlabel pdiffusion 990 -815 990 -815 0 feedthrough
rlabel pdiffusion 997 -815 997 -815 0 feedthrough
rlabel pdiffusion 1004 -815 1004 -815 0 feedthrough
rlabel pdiffusion 1011 -815 1011 -815 0 cellNo=613
rlabel pdiffusion 1018 -815 1018 -815 0 feedthrough
rlabel pdiffusion 1025 -815 1025 -815 0 feedthrough
rlabel pdiffusion 1032 -815 1032 -815 0 feedthrough
rlabel pdiffusion 1039 -815 1039 -815 0 feedthrough
rlabel pdiffusion 1046 -815 1046 -815 0 feedthrough
rlabel pdiffusion 1053 -815 1053 -815 0 feedthrough
rlabel pdiffusion 1060 -815 1060 -815 0 feedthrough
rlabel pdiffusion 1067 -815 1067 -815 0 feedthrough
rlabel pdiffusion 1074 -815 1074 -815 0 feedthrough
rlabel pdiffusion 1081 -815 1081 -815 0 feedthrough
rlabel pdiffusion 1088 -815 1088 -815 0 feedthrough
rlabel pdiffusion 1095 -815 1095 -815 0 cellNo=427
rlabel pdiffusion 1102 -815 1102 -815 0 feedthrough
rlabel pdiffusion 1109 -815 1109 -815 0 cellNo=383
rlabel pdiffusion 1116 -815 1116 -815 0 feedthrough
rlabel pdiffusion 1123 -815 1123 -815 0 feedthrough
rlabel pdiffusion 1130 -815 1130 -815 0 cellNo=657
rlabel pdiffusion 1137 -815 1137 -815 0 cellNo=111
rlabel pdiffusion 1144 -815 1144 -815 0 cellNo=349
rlabel pdiffusion 1151 -815 1151 -815 0 feedthrough
rlabel pdiffusion 1158 -815 1158 -815 0 cellNo=550
rlabel pdiffusion 1165 -815 1165 -815 0 feedthrough
rlabel pdiffusion 1172 -815 1172 -815 0 cellNo=298
rlabel pdiffusion 1179 -815 1179 -815 0 feedthrough
rlabel pdiffusion 1186 -815 1186 -815 0 feedthrough
rlabel pdiffusion 1193 -815 1193 -815 0 feedthrough
rlabel pdiffusion 1200 -815 1200 -815 0 feedthrough
rlabel pdiffusion 1207 -815 1207 -815 0 cellNo=221
rlabel pdiffusion 1214 -815 1214 -815 0 cellNo=4
rlabel pdiffusion 1221 -815 1221 -815 0 cellNo=214
rlabel pdiffusion 1228 -815 1228 -815 0 feedthrough
rlabel pdiffusion 1235 -815 1235 -815 0 feedthrough
rlabel pdiffusion 1242 -815 1242 -815 0 feedthrough
rlabel pdiffusion 1249 -815 1249 -815 0 feedthrough
rlabel pdiffusion 1256 -815 1256 -815 0 feedthrough
rlabel pdiffusion 1263 -815 1263 -815 0 feedthrough
rlabel pdiffusion 1270 -815 1270 -815 0 feedthrough
rlabel pdiffusion 1277 -815 1277 -815 0 feedthrough
rlabel pdiffusion 1284 -815 1284 -815 0 feedthrough
rlabel pdiffusion 1291 -815 1291 -815 0 feedthrough
rlabel pdiffusion 1298 -815 1298 -815 0 feedthrough
rlabel pdiffusion 1305 -815 1305 -815 0 feedthrough
rlabel pdiffusion 1312 -815 1312 -815 0 feedthrough
rlabel pdiffusion 1319 -815 1319 -815 0 feedthrough
rlabel pdiffusion 1326 -815 1326 -815 0 feedthrough
rlabel pdiffusion 1333 -815 1333 -815 0 cellNo=545
rlabel pdiffusion 1340 -815 1340 -815 0 feedthrough
rlabel pdiffusion 1347 -815 1347 -815 0 feedthrough
rlabel pdiffusion 1354 -815 1354 -815 0 feedthrough
rlabel pdiffusion 1361 -815 1361 -815 0 cellNo=35
rlabel pdiffusion 1368 -815 1368 -815 0 cellNo=477
rlabel pdiffusion 1375 -815 1375 -815 0 feedthrough
rlabel pdiffusion 1382 -815 1382 -815 0 feedthrough
rlabel pdiffusion 1389 -815 1389 -815 0 feedthrough
rlabel pdiffusion 1396 -815 1396 -815 0 feedthrough
rlabel pdiffusion 1403 -815 1403 -815 0 feedthrough
rlabel pdiffusion 1410 -815 1410 -815 0 feedthrough
rlabel pdiffusion 1417 -815 1417 -815 0 feedthrough
rlabel pdiffusion 1424 -815 1424 -815 0 feedthrough
rlabel pdiffusion 1431 -815 1431 -815 0 feedthrough
rlabel pdiffusion 1438 -815 1438 -815 0 feedthrough
rlabel pdiffusion 1445 -815 1445 -815 0 feedthrough
rlabel pdiffusion 1452 -815 1452 -815 0 feedthrough
rlabel pdiffusion 1459 -815 1459 -815 0 feedthrough
rlabel pdiffusion 1466 -815 1466 -815 0 feedthrough
rlabel pdiffusion 1473 -815 1473 -815 0 feedthrough
rlabel pdiffusion 1480 -815 1480 -815 0 feedthrough
rlabel pdiffusion 1487 -815 1487 -815 0 feedthrough
rlabel pdiffusion 1494 -815 1494 -815 0 feedthrough
rlabel pdiffusion 1501 -815 1501 -815 0 feedthrough
rlabel pdiffusion 1508 -815 1508 -815 0 feedthrough
rlabel pdiffusion 1515 -815 1515 -815 0 feedthrough
rlabel pdiffusion 1522 -815 1522 -815 0 feedthrough
rlabel pdiffusion 1529 -815 1529 -815 0 feedthrough
rlabel pdiffusion 1536 -815 1536 -815 0 cellNo=980
rlabel pdiffusion 1543 -815 1543 -815 0 feedthrough
rlabel pdiffusion 1550 -815 1550 -815 0 feedthrough
rlabel pdiffusion 1557 -815 1557 -815 0 feedthrough
rlabel pdiffusion 1564 -815 1564 -815 0 feedthrough
rlabel pdiffusion 1571 -815 1571 -815 0 feedthrough
rlabel pdiffusion 1578 -815 1578 -815 0 feedthrough
rlabel pdiffusion 1585 -815 1585 -815 0 feedthrough
rlabel pdiffusion 1592 -815 1592 -815 0 feedthrough
rlabel pdiffusion 1599 -815 1599 -815 0 feedthrough
rlabel pdiffusion 1606 -815 1606 -815 0 feedthrough
rlabel pdiffusion 1613 -815 1613 -815 0 feedthrough
rlabel pdiffusion 1620 -815 1620 -815 0 feedthrough
rlabel pdiffusion 1627 -815 1627 -815 0 feedthrough
rlabel pdiffusion 1634 -815 1634 -815 0 feedthrough
rlabel pdiffusion 1641 -815 1641 -815 0 feedthrough
rlabel pdiffusion 1648 -815 1648 -815 0 feedthrough
rlabel pdiffusion 1655 -815 1655 -815 0 feedthrough
rlabel pdiffusion 1662 -815 1662 -815 0 feedthrough
rlabel pdiffusion 1669 -815 1669 -815 0 feedthrough
rlabel pdiffusion 1676 -815 1676 -815 0 feedthrough
rlabel pdiffusion 1683 -815 1683 -815 0 feedthrough
rlabel pdiffusion 1690 -815 1690 -815 0 feedthrough
rlabel pdiffusion 1697 -815 1697 -815 0 feedthrough
rlabel pdiffusion 1704 -815 1704 -815 0 feedthrough
rlabel pdiffusion 1711 -815 1711 -815 0 feedthrough
rlabel pdiffusion 1718 -815 1718 -815 0 feedthrough
rlabel pdiffusion 1725 -815 1725 -815 0 feedthrough
rlabel pdiffusion 1732 -815 1732 -815 0 feedthrough
rlabel pdiffusion 1739 -815 1739 -815 0 feedthrough
rlabel pdiffusion 1746 -815 1746 -815 0 feedthrough
rlabel pdiffusion 1753 -815 1753 -815 0 feedthrough
rlabel pdiffusion 1760 -815 1760 -815 0 feedthrough
rlabel pdiffusion 1767 -815 1767 -815 0 feedthrough
rlabel pdiffusion 1774 -815 1774 -815 0 feedthrough
rlabel pdiffusion 1781 -815 1781 -815 0 feedthrough
rlabel pdiffusion 1788 -815 1788 -815 0 feedthrough
rlabel pdiffusion 1795 -815 1795 -815 0 feedthrough
rlabel pdiffusion 1802 -815 1802 -815 0 feedthrough
rlabel pdiffusion 1809 -815 1809 -815 0 feedthrough
rlabel pdiffusion 1816 -815 1816 -815 0 feedthrough
rlabel pdiffusion 1823 -815 1823 -815 0 feedthrough
rlabel pdiffusion 1830 -815 1830 -815 0 feedthrough
rlabel pdiffusion 1837 -815 1837 -815 0 feedthrough
rlabel pdiffusion 1844 -815 1844 -815 0 feedthrough
rlabel pdiffusion 1851 -815 1851 -815 0 feedthrough
rlabel pdiffusion 1858 -815 1858 -815 0 feedthrough
rlabel pdiffusion 1865 -815 1865 -815 0 feedthrough
rlabel pdiffusion 1872 -815 1872 -815 0 feedthrough
rlabel pdiffusion 1879 -815 1879 -815 0 feedthrough
rlabel pdiffusion 1886 -815 1886 -815 0 feedthrough
rlabel pdiffusion 1893 -815 1893 -815 0 feedthrough
rlabel pdiffusion 1900 -815 1900 -815 0 feedthrough
rlabel pdiffusion 1907 -815 1907 -815 0 feedthrough
rlabel pdiffusion 1914 -815 1914 -815 0 feedthrough
rlabel pdiffusion 1921 -815 1921 -815 0 feedthrough
rlabel pdiffusion 1928 -815 1928 -815 0 feedthrough
rlabel pdiffusion 1935 -815 1935 -815 0 feedthrough
rlabel pdiffusion 1942 -815 1942 -815 0 feedthrough
rlabel pdiffusion 1949 -815 1949 -815 0 feedthrough
rlabel pdiffusion 1956 -815 1956 -815 0 feedthrough
rlabel pdiffusion 1963 -815 1963 -815 0 feedthrough
rlabel pdiffusion 1970 -815 1970 -815 0 feedthrough
rlabel pdiffusion 1977 -815 1977 -815 0 feedthrough
rlabel pdiffusion 1984 -815 1984 -815 0 feedthrough
rlabel pdiffusion 1991 -815 1991 -815 0 feedthrough
rlabel pdiffusion 1998 -815 1998 -815 0 feedthrough
rlabel pdiffusion 2005 -815 2005 -815 0 feedthrough
rlabel pdiffusion 2012 -815 2012 -815 0 feedthrough
rlabel pdiffusion 2019 -815 2019 -815 0 feedthrough
rlabel pdiffusion 2026 -815 2026 -815 0 feedthrough
rlabel pdiffusion 2033 -815 2033 -815 0 feedthrough
rlabel pdiffusion 2040 -815 2040 -815 0 feedthrough
rlabel pdiffusion 2047 -815 2047 -815 0 feedthrough
rlabel pdiffusion 2054 -815 2054 -815 0 feedthrough
rlabel pdiffusion 2061 -815 2061 -815 0 feedthrough
rlabel pdiffusion 2068 -815 2068 -815 0 feedthrough
rlabel pdiffusion 2075 -815 2075 -815 0 feedthrough
rlabel pdiffusion 2082 -815 2082 -815 0 feedthrough
rlabel pdiffusion 2089 -815 2089 -815 0 feedthrough
rlabel pdiffusion 2096 -815 2096 -815 0 feedthrough
rlabel pdiffusion 2103 -815 2103 -815 0 feedthrough
rlabel pdiffusion 2110 -815 2110 -815 0 feedthrough
rlabel pdiffusion 2117 -815 2117 -815 0 feedthrough
rlabel pdiffusion 2124 -815 2124 -815 0 feedthrough
rlabel pdiffusion 2131 -815 2131 -815 0 feedthrough
rlabel pdiffusion 2138 -815 2138 -815 0 feedthrough
rlabel pdiffusion 2145 -815 2145 -815 0 feedthrough
rlabel pdiffusion 2152 -815 2152 -815 0 feedthrough
rlabel pdiffusion 2159 -815 2159 -815 0 feedthrough
rlabel pdiffusion 2166 -815 2166 -815 0 feedthrough
rlabel pdiffusion 2173 -815 2173 -815 0 feedthrough
rlabel pdiffusion 2180 -815 2180 -815 0 feedthrough
rlabel pdiffusion 2187 -815 2187 -815 0 feedthrough
rlabel pdiffusion 2194 -815 2194 -815 0 feedthrough
rlabel pdiffusion 2201 -815 2201 -815 0 feedthrough
rlabel pdiffusion 2208 -815 2208 -815 0 feedthrough
rlabel pdiffusion 2215 -815 2215 -815 0 feedthrough
rlabel pdiffusion 2222 -815 2222 -815 0 feedthrough
rlabel pdiffusion 2229 -815 2229 -815 0 feedthrough
rlabel pdiffusion 2236 -815 2236 -815 0 feedthrough
rlabel pdiffusion 2243 -815 2243 -815 0 feedthrough
rlabel pdiffusion 2250 -815 2250 -815 0 feedthrough
rlabel pdiffusion 2257 -815 2257 -815 0 feedthrough
rlabel pdiffusion 2264 -815 2264 -815 0 feedthrough
rlabel pdiffusion 2271 -815 2271 -815 0 feedthrough
rlabel pdiffusion 2278 -815 2278 -815 0 feedthrough
rlabel pdiffusion 2285 -815 2285 -815 0 feedthrough
rlabel pdiffusion 2292 -815 2292 -815 0 feedthrough
rlabel pdiffusion 2299 -815 2299 -815 0 feedthrough
rlabel pdiffusion 2306 -815 2306 -815 0 feedthrough
rlabel pdiffusion 2313 -815 2313 -815 0 feedthrough
rlabel pdiffusion 2320 -815 2320 -815 0 feedthrough
rlabel pdiffusion 2327 -815 2327 -815 0 feedthrough
rlabel pdiffusion 2348 -815 2348 -815 0 feedthrough
rlabel pdiffusion 2404 -815 2404 -815 0 feedthrough
rlabel pdiffusion 3 -1004 3 -1004 0 feedthrough
rlabel pdiffusion 10 -1004 10 -1004 0 feedthrough
rlabel pdiffusion 17 -1004 17 -1004 0 feedthrough
rlabel pdiffusion 24 -1004 24 -1004 0 feedthrough
rlabel pdiffusion 31 -1004 31 -1004 0 feedthrough
rlabel pdiffusion 38 -1004 38 -1004 0 feedthrough
rlabel pdiffusion 45 -1004 45 -1004 0 feedthrough
rlabel pdiffusion 52 -1004 52 -1004 0 feedthrough
rlabel pdiffusion 59 -1004 59 -1004 0 feedthrough
rlabel pdiffusion 66 -1004 66 -1004 0 feedthrough
rlabel pdiffusion 73 -1004 73 -1004 0 feedthrough
rlabel pdiffusion 80 -1004 80 -1004 0 feedthrough
rlabel pdiffusion 87 -1004 87 -1004 0 feedthrough
rlabel pdiffusion 94 -1004 94 -1004 0 cellNo=163
rlabel pdiffusion 101 -1004 101 -1004 0 cellNo=933
rlabel pdiffusion 108 -1004 108 -1004 0 feedthrough
rlabel pdiffusion 115 -1004 115 -1004 0 feedthrough
rlabel pdiffusion 122 -1004 122 -1004 0 feedthrough
rlabel pdiffusion 129 -1004 129 -1004 0 feedthrough
rlabel pdiffusion 136 -1004 136 -1004 0 cellNo=127
rlabel pdiffusion 143 -1004 143 -1004 0 feedthrough
rlabel pdiffusion 150 -1004 150 -1004 0 feedthrough
rlabel pdiffusion 157 -1004 157 -1004 0 feedthrough
rlabel pdiffusion 164 -1004 164 -1004 0 feedthrough
rlabel pdiffusion 171 -1004 171 -1004 0 feedthrough
rlabel pdiffusion 178 -1004 178 -1004 0 cellNo=247
rlabel pdiffusion 185 -1004 185 -1004 0 cellNo=392
rlabel pdiffusion 192 -1004 192 -1004 0 feedthrough
rlabel pdiffusion 199 -1004 199 -1004 0 feedthrough
rlabel pdiffusion 206 -1004 206 -1004 0 feedthrough
rlabel pdiffusion 213 -1004 213 -1004 0 feedthrough
rlabel pdiffusion 220 -1004 220 -1004 0 cellNo=389
rlabel pdiffusion 227 -1004 227 -1004 0 feedthrough
rlabel pdiffusion 234 -1004 234 -1004 0 feedthrough
rlabel pdiffusion 241 -1004 241 -1004 0 feedthrough
rlabel pdiffusion 248 -1004 248 -1004 0 feedthrough
rlabel pdiffusion 255 -1004 255 -1004 0 feedthrough
rlabel pdiffusion 262 -1004 262 -1004 0 feedthrough
rlabel pdiffusion 269 -1004 269 -1004 0 cellNo=866
rlabel pdiffusion 276 -1004 276 -1004 0 feedthrough
rlabel pdiffusion 283 -1004 283 -1004 0 feedthrough
rlabel pdiffusion 290 -1004 290 -1004 0 feedthrough
rlabel pdiffusion 297 -1004 297 -1004 0 feedthrough
rlabel pdiffusion 304 -1004 304 -1004 0 feedthrough
rlabel pdiffusion 311 -1004 311 -1004 0 feedthrough
rlabel pdiffusion 318 -1004 318 -1004 0 feedthrough
rlabel pdiffusion 325 -1004 325 -1004 0 feedthrough
rlabel pdiffusion 332 -1004 332 -1004 0 feedthrough
rlabel pdiffusion 339 -1004 339 -1004 0 feedthrough
rlabel pdiffusion 346 -1004 346 -1004 0 feedthrough
rlabel pdiffusion 353 -1004 353 -1004 0 feedthrough
rlabel pdiffusion 360 -1004 360 -1004 0 feedthrough
rlabel pdiffusion 367 -1004 367 -1004 0 feedthrough
rlabel pdiffusion 374 -1004 374 -1004 0 cellNo=188
rlabel pdiffusion 381 -1004 381 -1004 0 feedthrough
rlabel pdiffusion 388 -1004 388 -1004 0 cellNo=361
rlabel pdiffusion 395 -1004 395 -1004 0 feedthrough
rlabel pdiffusion 402 -1004 402 -1004 0 feedthrough
rlabel pdiffusion 409 -1004 409 -1004 0 feedthrough
rlabel pdiffusion 416 -1004 416 -1004 0 feedthrough
rlabel pdiffusion 423 -1004 423 -1004 0 feedthrough
rlabel pdiffusion 430 -1004 430 -1004 0 feedthrough
rlabel pdiffusion 437 -1004 437 -1004 0 feedthrough
rlabel pdiffusion 444 -1004 444 -1004 0 feedthrough
rlabel pdiffusion 451 -1004 451 -1004 0 feedthrough
rlabel pdiffusion 458 -1004 458 -1004 0 feedthrough
rlabel pdiffusion 465 -1004 465 -1004 0 feedthrough
rlabel pdiffusion 472 -1004 472 -1004 0 feedthrough
rlabel pdiffusion 479 -1004 479 -1004 0 feedthrough
rlabel pdiffusion 486 -1004 486 -1004 0 feedthrough
rlabel pdiffusion 493 -1004 493 -1004 0 feedthrough
rlabel pdiffusion 500 -1004 500 -1004 0 feedthrough
rlabel pdiffusion 507 -1004 507 -1004 0 feedthrough
rlabel pdiffusion 514 -1004 514 -1004 0 feedthrough
rlabel pdiffusion 521 -1004 521 -1004 0 feedthrough
rlabel pdiffusion 528 -1004 528 -1004 0 cellNo=142
rlabel pdiffusion 535 -1004 535 -1004 0 feedthrough
rlabel pdiffusion 542 -1004 542 -1004 0 feedthrough
rlabel pdiffusion 549 -1004 549 -1004 0 feedthrough
rlabel pdiffusion 556 -1004 556 -1004 0 feedthrough
rlabel pdiffusion 563 -1004 563 -1004 0 feedthrough
rlabel pdiffusion 570 -1004 570 -1004 0 feedthrough
rlabel pdiffusion 577 -1004 577 -1004 0 feedthrough
rlabel pdiffusion 584 -1004 584 -1004 0 feedthrough
rlabel pdiffusion 591 -1004 591 -1004 0 feedthrough
rlabel pdiffusion 598 -1004 598 -1004 0 feedthrough
rlabel pdiffusion 605 -1004 605 -1004 0 feedthrough
rlabel pdiffusion 612 -1004 612 -1004 0 cellNo=79
rlabel pdiffusion 619 -1004 619 -1004 0 feedthrough
rlabel pdiffusion 626 -1004 626 -1004 0 cellNo=276
rlabel pdiffusion 633 -1004 633 -1004 0 cellNo=974
rlabel pdiffusion 640 -1004 640 -1004 0 feedthrough
rlabel pdiffusion 647 -1004 647 -1004 0 feedthrough
rlabel pdiffusion 654 -1004 654 -1004 0 feedthrough
rlabel pdiffusion 661 -1004 661 -1004 0 feedthrough
rlabel pdiffusion 668 -1004 668 -1004 0 feedthrough
rlabel pdiffusion 675 -1004 675 -1004 0 feedthrough
rlabel pdiffusion 682 -1004 682 -1004 0 feedthrough
rlabel pdiffusion 689 -1004 689 -1004 0 feedthrough
rlabel pdiffusion 696 -1004 696 -1004 0 feedthrough
rlabel pdiffusion 703 -1004 703 -1004 0 feedthrough
rlabel pdiffusion 710 -1004 710 -1004 0 feedthrough
rlabel pdiffusion 717 -1004 717 -1004 0 cellNo=495
rlabel pdiffusion 724 -1004 724 -1004 0 feedthrough
rlabel pdiffusion 731 -1004 731 -1004 0 feedthrough
rlabel pdiffusion 738 -1004 738 -1004 0 feedthrough
rlabel pdiffusion 745 -1004 745 -1004 0 feedthrough
rlabel pdiffusion 752 -1004 752 -1004 0 feedthrough
rlabel pdiffusion 759 -1004 759 -1004 0 feedthrough
rlabel pdiffusion 766 -1004 766 -1004 0 feedthrough
rlabel pdiffusion 773 -1004 773 -1004 0 cellNo=460
rlabel pdiffusion 780 -1004 780 -1004 0 cellNo=878
rlabel pdiffusion 787 -1004 787 -1004 0 feedthrough
rlabel pdiffusion 794 -1004 794 -1004 0 cellNo=402
rlabel pdiffusion 801 -1004 801 -1004 0 feedthrough
rlabel pdiffusion 808 -1004 808 -1004 0 feedthrough
rlabel pdiffusion 815 -1004 815 -1004 0 cellNo=658
rlabel pdiffusion 822 -1004 822 -1004 0 feedthrough
rlabel pdiffusion 829 -1004 829 -1004 0 cellNo=26
rlabel pdiffusion 836 -1004 836 -1004 0 feedthrough
rlabel pdiffusion 843 -1004 843 -1004 0 feedthrough
rlabel pdiffusion 850 -1004 850 -1004 0 feedthrough
rlabel pdiffusion 857 -1004 857 -1004 0 feedthrough
rlabel pdiffusion 864 -1004 864 -1004 0 feedthrough
rlabel pdiffusion 871 -1004 871 -1004 0 feedthrough
rlabel pdiffusion 878 -1004 878 -1004 0 feedthrough
rlabel pdiffusion 885 -1004 885 -1004 0 feedthrough
rlabel pdiffusion 892 -1004 892 -1004 0 feedthrough
rlabel pdiffusion 899 -1004 899 -1004 0 feedthrough
rlabel pdiffusion 906 -1004 906 -1004 0 feedthrough
rlabel pdiffusion 913 -1004 913 -1004 0 feedthrough
rlabel pdiffusion 920 -1004 920 -1004 0 feedthrough
rlabel pdiffusion 927 -1004 927 -1004 0 feedthrough
rlabel pdiffusion 934 -1004 934 -1004 0 cellNo=122
rlabel pdiffusion 941 -1004 941 -1004 0 feedthrough
rlabel pdiffusion 948 -1004 948 -1004 0 feedthrough
rlabel pdiffusion 955 -1004 955 -1004 0 cellNo=543
rlabel pdiffusion 962 -1004 962 -1004 0 feedthrough
rlabel pdiffusion 969 -1004 969 -1004 0 feedthrough
rlabel pdiffusion 976 -1004 976 -1004 0 feedthrough
rlabel pdiffusion 983 -1004 983 -1004 0 feedthrough
rlabel pdiffusion 990 -1004 990 -1004 0 feedthrough
rlabel pdiffusion 997 -1004 997 -1004 0 feedthrough
rlabel pdiffusion 1004 -1004 1004 -1004 0 feedthrough
rlabel pdiffusion 1011 -1004 1011 -1004 0 feedthrough
rlabel pdiffusion 1018 -1004 1018 -1004 0 cellNo=699
rlabel pdiffusion 1025 -1004 1025 -1004 0 feedthrough
rlabel pdiffusion 1032 -1004 1032 -1004 0 feedthrough
rlabel pdiffusion 1039 -1004 1039 -1004 0 cellNo=810
rlabel pdiffusion 1046 -1004 1046 -1004 0 feedthrough
rlabel pdiffusion 1053 -1004 1053 -1004 0 cellNo=176
rlabel pdiffusion 1060 -1004 1060 -1004 0 cellNo=39
rlabel pdiffusion 1067 -1004 1067 -1004 0 feedthrough
rlabel pdiffusion 1074 -1004 1074 -1004 0 feedthrough
rlabel pdiffusion 1081 -1004 1081 -1004 0 feedthrough
rlabel pdiffusion 1088 -1004 1088 -1004 0 feedthrough
rlabel pdiffusion 1095 -1004 1095 -1004 0 feedthrough
rlabel pdiffusion 1102 -1004 1102 -1004 0 feedthrough
rlabel pdiffusion 1109 -1004 1109 -1004 0 feedthrough
rlabel pdiffusion 1116 -1004 1116 -1004 0 feedthrough
rlabel pdiffusion 1123 -1004 1123 -1004 0 cellNo=191
rlabel pdiffusion 1130 -1004 1130 -1004 0 feedthrough
rlabel pdiffusion 1137 -1004 1137 -1004 0 feedthrough
rlabel pdiffusion 1144 -1004 1144 -1004 0 feedthrough
rlabel pdiffusion 1151 -1004 1151 -1004 0 feedthrough
rlabel pdiffusion 1158 -1004 1158 -1004 0 feedthrough
rlabel pdiffusion 1165 -1004 1165 -1004 0 feedthrough
rlabel pdiffusion 1172 -1004 1172 -1004 0 cellNo=679
rlabel pdiffusion 1179 -1004 1179 -1004 0 feedthrough
rlabel pdiffusion 1186 -1004 1186 -1004 0 feedthrough
rlabel pdiffusion 1193 -1004 1193 -1004 0 cellNo=494
rlabel pdiffusion 1200 -1004 1200 -1004 0 feedthrough
rlabel pdiffusion 1207 -1004 1207 -1004 0 feedthrough
rlabel pdiffusion 1214 -1004 1214 -1004 0 feedthrough
rlabel pdiffusion 1221 -1004 1221 -1004 0 feedthrough
rlabel pdiffusion 1228 -1004 1228 -1004 0 feedthrough
rlabel pdiffusion 1235 -1004 1235 -1004 0 feedthrough
rlabel pdiffusion 1242 -1004 1242 -1004 0 cellNo=684
rlabel pdiffusion 1249 -1004 1249 -1004 0 feedthrough
rlabel pdiffusion 1256 -1004 1256 -1004 0 feedthrough
rlabel pdiffusion 1263 -1004 1263 -1004 0 feedthrough
rlabel pdiffusion 1270 -1004 1270 -1004 0 cellNo=990
rlabel pdiffusion 1277 -1004 1277 -1004 0 feedthrough
rlabel pdiffusion 1284 -1004 1284 -1004 0 cellNo=652
rlabel pdiffusion 1291 -1004 1291 -1004 0 feedthrough
rlabel pdiffusion 1298 -1004 1298 -1004 0 feedthrough
rlabel pdiffusion 1305 -1004 1305 -1004 0 feedthrough
rlabel pdiffusion 1312 -1004 1312 -1004 0 cellNo=172
rlabel pdiffusion 1319 -1004 1319 -1004 0 feedthrough
rlabel pdiffusion 1326 -1004 1326 -1004 0 feedthrough
rlabel pdiffusion 1333 -1004 1333 -1004 0 feedthrough
rlabel pdiffusion 1340 -1004 1340 -1004 0 feedthrough
rlabel pdiffusion 1347 -1004 1347 -1004 0 feedthrough
rlabel pdiffusion 1354 -1004 1354 -1004 0 feedthrough
rlabel pdiffusion 1361 -1004 1361 -1004 0 feedthrough
rlabel pdiffusion 1368 -1004 1368 -1004 0 feedthrough
rlabel pdiffusion 1375 -1004 1375 -1004 0 feedthrough
rlabel pdiffusion 1382 -1004 1382 -1004 0 feedthrough
rlabel pdiffusion 1389 -1004 1389 -1004 0 feedthrough
rlabel pdiffusion 1396 -1004 1396 -1004 0 cellNo=219
rlabel pdiffusion 1403 -1004 1403 -1004 0 feedthrough
rlabel pdiffusion 1410 -1004 1410 -1004 0 feedthrough
rlabel pdiffusion 1417 -1004 1417 -1004 0 feedthrough
rlabel pdiffusion 1424 -1004 1424 -1004 0 feedthrough
rlabel pdiffusion 1431 -1004 1431 -1004 0 feedthrough
rlabel pdiffusion 1438 -1004 1438 -1004 0 feedthrough
rlabel pdiffusion 1445 -1004 1445 -1004 0 feedthrough
rlabel pdiffusion 1452 -1004 1452 -1004 0 feedthrough
rlabel pdiffusion 1459 -1004 1459 -1004 0 feedthrough
rlabel pdiffusion 1466 -1004 1466 -1004 0 feedthrough
rlabel pdiffusion 1473 -1004 1473 -1004 0 feedthrough
rlabel pdiffusion 1480 -1004 1480 -1004 0 feedthrough
rlabel pdiffusion 1487 -1004 1487 -1004 0 feedthrough
rlabel pdiffusion 1494 -1004 1494 -1004 0 feedthrough
rlabel pdiffusion 1501 -1004 1501 -1004 0 feedthrough
rlabel pdiffusion 1508 -1004 1508 -1004 0 feedthrough
rlabel pdiffusion 1515 -1004 1515 -1004 0 cellNo=103
rlabel pdiffusion 1522 -1004 1522 -1004 0 feedthrough
rlabel pdiffusion 1529 -1004 1529 -1004 0 feedthrough
rlabel pdiffusion 1536 -1004 1536 -1004 0 feedthrough
rlabel pdiffusion 1543 -1004 1543 -1004 0 feedthrough
rlabel pdiffusion 1550 -1004 1550 -1004 0 feedthrough
rlabel pdiffusion 1557 -1004 1557 -1004 0 feedthrough
rlabel pdiffusion 1564 -1004 1564 -1004 0 feedthrough
rlabel pdiffusion 1571 -1004 1571 -1004 0 cellNo=630
rlabel pdiffusion 1578 -1004 1578 -1004 0 cellNo=682
rlabel pdiffusion 1585 -1004 1585 -1004 0 feedthrough
rlabel pdiffusion 1592 -1004 1592 -1004 0 feedthrough
rlabel pdiffusion 1599 -1004 1599 -1004 0 feedthrough
rlabel pdiffusion 1606 -1004 1606 -1004 0 feedthrough
rlabel pdiffusion 1613 -1004 1613 -1004 0 feedthrough
rlabel pdiffusion 1620 -1004 1620 -1004 0 feedthrough
rlabel pdiffusion 1627 -1004 1627 -1004 0 feedthrough
rlabel pdiffusion 1634 -1004 1634 -1004 0 feedthrough
rlabel pdiffusion 1641 -1004 1641 -1004 0 feedthrough
rlabel pdiffusion 1648 -1004 1648 -1004 0 feedthrough
rlabel pdiffusion 1655 -1004 1655 -1004 0 feedthrough
rlabel pdiffusion 1662 -1004 1662 -1004 0 feedthrough
rlabel pdiffusion 1669 -1004 1669 -1004 0 feedthrough
rlabel pdiffusion 1676 -1004 1676 -1004 0 feedthrough
rlabel pdiffusion 1683 -1004 1683 -1004 0 feedthrough
rlabel pdiffusion 1690 -1004 1690 -1004 0 feedthrough
rlabel pdiffusion 1697 -1004 1697 -1004 0 feedthrough
rlabel pdiffusion 1704 -1004 1704 -1004 0 feedthrough
rlabel pdiffusion 1711 -1004 1711 -1004 0 feedthrough
rlabel pdiffusion 1718 -1004 1718 -1004 0 feedthrough
rlabel pdiffusion 1725 -1004 1725 -1004 0 feedthrough
rlabel pdiffusion 1732 -1004 1732 -1004 0 feedthrough
rlabel pdiffusion 1739 -1004 1739 -1004 0 feedthrough
rlabel pdiffusion 1746 -1004 1746 -1004 0 feedthrough
rlabel pdiffusion 1753 -1004 1753 -1004 0 feedthrough
rlabel pdiffusion 1760 -1004 1760 -1004 0 feedthrough
rlabel pdiffusion 1767 -1004 1767 -1004 0 feedthrough
rlabel pdiffusion 1774 -1004 1774 -1004 0 feedthrough
rlabel pdiffusion 1781 -1004 1781 -1004 0 feedthrough
rlabel pdiffusion 1788 -1004 1788 -1004 0 feedthrough
rlabel pdiffusion 1795 -1004 1795 -1004 0 feedthrough
rlabel pdiffusion 1802 -1004 1802 -1004 0 feedthrough
rlabel pdiffusion 1809 -1004 1809 -1004 0 feedthrough
rlabel pdiffusion 1816 -1004 1816 -1004 0 feedthrough
rlabel pdiffusion 1823 -1004 1823 -1004 0 feedthrough
rlabel pdiffusion 1830 -1004 1830 -1004 0 feedthrough
rlabel pdiffusion 1837 -1004 1837 -1004 0 feedthrough
rlabel pdiffusion 1844 -1004 1844 -1004 0 feedthrough
rlabel pdiffusion 1851 -1004 1851 -1004 0 feedthrough
rlabel pdiffusion 1858 -1004 1858 -1004 0 feedthrough
rlabel pdiffusion 1865 -1004 1865 -1004 0 feedthrough
rlabel pdiffusion 1872 -1004 1872 -1004 0 feedthrough
rlabel pdiffusion 1879 -1004 1879 -1004 0 feedthrough
rlabel pdiffusion 1886 -1004 1886 -1004 0 feedthrough
rlabel pdiffusion 1893 -1004 1893 -1004 0 feedthrough
rlabel pdiffusion 1900 -1004 1900 -1004 0 feedthrough
rlabel pdiffusion 1907 -1004 1907 -1004 0 feedthrough
rlabel pdiffusion 1914 -1004 1914 -1004 0 feedthrough
rlabel pdiffusion 1921 -1004 1921 -1004 0 feedthrough
rlabel pdiffusion 1928 -1004 1928 -1004 0 feedthrough
rlabel pdiffusion 1935 -1004 1935 -1004 0 feedthrough
rlabel pdiffusion 1942 -1004 1942 -1004 0 feedthrough
rlabel pdiffusion 1949 -1004 1949 -1004 0 feedthrough
rlabel pdiffusion 1956 -1004 1956 -1004 0 feedthrough
rlabel pdiffusion 1963 -1004 1963 -1004 0 feedthrough
rlabel pdiffusion 1970 -1004 1970 -1004 0 feedthrough
rlabel pdiffusion 1977 -1004 1977 -1004 0 feedthrough
rlabel pdiffusion 1984 -1004 1984 -1004 0 feedthrough
rlabel pdiffusion 1991 -1004 1991 -1004 0 feedthrough
rlabel pdiffusion 1998 -1004 1998 -1004 0 feedthrough
rlabel pdiffusion 2005 -1004 2005 -1004 0 feedthrough
rlabel pdiffusion 2012 -1004 2012 -1004 0 feedthrough
rlabel pdiffusion 2019 -1004 2019 -1004 0 feedthrough
rlabel pdiffusion 2026 -1004 2026 -1004 0 feedthrough
rlabel pdiffusion 2033 -1004 2033 -1004 0 feedthrough
rlabel pdiffusion 2040 -1004 2040 -1004 0 feedthrough
rlabel pdiffusion 2047 -1004 2047 -1004 0 feedthrough
rlabel pdiffusion 2054 -1004 2054 -1004 0 feedthrough
rlabel pdiffusion 2061 -1004 2061 -1004 0 feedthrough
rlabel pdiffusion 2068 -1004 2068 -1004 0 feedthrough
rlabel pdiffusion 2075 -1004 2075 -1004 0 feedthrough
rlabel pdiffusion 2082 -1004 2082 -1004 0 feedthrough
rlabel pdiffusion 2089 -1004 2089 -1004 0 feedthrough
rlabel pdiffusion 2096 -1004 2096 -1004 0 feedthrough
rlabel pdiffusion 2103 -1004 2103 -1004 0 feedthrough
rlabel pdiffusion 2110 -1004 2110 -1004 0 feedthrough
rlabel pdiffusion 2117 -1004 2117 -1004 0 feedthrough
rlabel pdiffusion 2124 -1004 2124 -1004 0 feedthrough
rlabel pdiffusion 2131 -1004 2131 -1004 0 feedthrough
rlabel pdiffusion 2138 -1004 2138 -1004 0 feedthrough
rlabel pdiffusion 2145 -1004 2145 -1004 0 feedthrough
rlabel pdiffusion 2152 -1004 2152 -1004 0 feedthrough
rlabel pdiffusion 2159 -1004 2159 -1004 0 feedthrough
rlabel pdiffusion 2166 -1004 2166 -1004 0 feedthrough
rlabel pdiffusion 2173 -1004 2173 -1004 0 feedthrough
rlabel pdiffusion 2180 -1004 2180 -1004 0 feedthrough
rlabel pdiffusion 2187 -1004 2187 -1004 0 feedthrough
rlabel pdiffusion 2194 -1004 2194 -1004 0 feedthrough
rlabel pdiffusion 2201 -1004 2201 -1004 0 feedthrough
rlabel pdiffusion 2208 -1004 2208 -1004 0 feedthrough
rlabel pdiffusion 2215 -1004 2215 -1004 0 feedthrough
rlabel pdiffusion 2222 -1004 2222 -1004 0 feedthrough
rlabel pdiffusion 2229 -1004 2229 -1004 0 feedthrough
rlabel pdiffusion 2236 -1004 2236 -1004 0 feedthrough
rlabel pdiffusion 2243 -1004 2243 -1004 0 feedthrough
rlabel pdiffusion 2250 -1004 2250 -1004 0 feedthrough
rlabel pdiffusion 2257 -1004 2257 -1004 0 feedthrough
rlabel pdiffusion 2264 -1004 2264 -1004 0 feedthrough
rlabel pdiffusion 2271 -1004 2271 -1004 0 feedthrough
rlabel pdiffusion 2278 -1004 2278 -1004 0 feedthrough
rlabel pdiffusion 2285 -1004 2285 -1004 0 feedthrough
rlabel pdiffusion 2292 -1004 2292 -1004 0 feedthrough
rlabel pdiffusion 2299 -1004 2299 -1004 0 feedthrough
rlabel pdiffusion 2306 -1004 2306 -1004 0 feedthrough
rlabel pdiffusion 2313 -1004 2313 -1004 0 feedthrough
rlabel pdiffusion 2320 -1004 2320 -1004 0 feedthrough
rlabel pdiffusion 2327 -1004 2327 -1004 0 feedthrough
rlabel pdiffusion 2334 -1004 2334 -1004 0 cellNo=908
rlabel pdiffusion 2341 -1004 2341 -1004 0 cellNo=232
rlabel pdiffusion 2348 -1004 2348 -1004 0 cellNo=540
rlabel pdiffusion 2355 -1004 2355 -1004 0 feedthrough
rlabel pdiffusion 2362 -1004 2362 -1004 0 feedthrough
rlabel pdiffusion 2369 -1004 2369 -1004 0 feedthrough
rlabel pdiffusion 2376 -1004 2376 -1004 0 feedthrough
rlabel pdiffusion 2404 -1004 2404 -1004 0 feedthrough
rlabel pdiffusion 2418 -1004 2418 -1004 0 feedthrough
rlabel pdiffusion 3 -1171 3 -1171 0 cellNo=1013
rlabel pdiffusion 10 -1171 10 -1171 0 feedthrough
rlabel pdiffusion 17 -1171 17 -1171 0 feedthrough
rlabel pdiffusion 24 -1171 24 -1171 0 feedthrough
rlabel pdiffusion 31 -1171 31 -1171 0 feedthrough
rlabel pdiffusion 38 -1171 38 -1171 0 feedthrough
rlabel pdiffusion 45 -1171 45 -1171 0 feedthrough
rlabel pdiffusion 52 -1171 52 -1171 0 feedthrough
rlabel pdiffusion 59 -1171 59 -1171 0 feedthrough
rlabel pdiffusion 66 -1171 66 -1171 0 feedthrough
rlabel pdiffusion 73 -1171 73 -1171 0 feedthrough
rlabel pdiffusion 80 -1171 80 -1171 0 feedthrough
rlabel pdiffusion 87 -1171 87 -1171 0 cellNo=507
rlabel pdiffusion 94 -1171 94 -1171 0 feedthrough
rlabel pdiffusion 101 -1171 101 -1171 0 feedthrough
rlabel pdiffusion 108 -1171 108 -1171 0 cellNo=606
rlabel pdiffusion 115 -1171 115 -1171 0 cellNo=382
rlabel pdiffusion 122 -1171 122 -1171 0 feedthrough
rlabel pdiffusion 129 -1171 129 -1171 0 feedthrough
rlabel pdiffusion 136 -1171 136 -1171 0 cellNo=421
rlabel pdiffusion 143 -1171 143 -1171 0 cellNo=362
rlabel pdiffusion 150 -1171 150 -1171 0 feedthrough
rlabel pdiffusion 157 -1171 157 -1171 0 feedthrough
rlabel pdiffusion 164 -1171 164 -1171 0 feedthrough
rlabel pdiffusion 171 -1171 171 -1171 0 feedthrough
rlabel pdiffusion 178 -1171 178 -1171 0 feedthrough
rlabel pdiffusion 185 -1171 185 -1171 0 feedthrough
rlabel pdiffusion 192 -1171 192 -1171 0 feedthrough
rlabel pdiffusion 199 -1171 199 -1171 0 feedthrough
rlabel pdiffusion 206 -1171 206 -1171 0 feedthrough
rlabel pdiffusion 213 -1171 213 -1171 0 feedthrough
rlabel pdiffusion 220 -1171 220 -1171 0 feedthrough
rlabel pdiffusion 227 -1171 227 -1171 0 feedthrough
rlabel pdiffusion 234 -1171 234 -1171 0 feedthrough
rlabel pdiffusion 241 -1171 241 -1171 0 cellNo=750
rlabel pdiffusion 248 -1171 248 -1171 0 feedthrough
rlabel pdiffusion 255 -1171 255 -1171 0 feedthrough
rlabel pdiffusion 262 -1171 262 -1171 0 feedthrough
rlabel pdiffusion 269 -1171 269 -1171 0 feedthrough
rlabel pdiffusion 276 -1171 276 -1171 0 feedthrough
rlabel pdiffusion 283 -1171 283 -1171 0 feedthrough
rlabel pdiffusion 290 -1171 290 -1171 0 feedthrough
rlabel pdiffusion 297 -1171 297 -1171 0 feedthrough
rlabel pdiffusion 304 -1171 304 -1171 0 feedthrough
rlabel pdiffusion 311 -1171 311 -1171 0 feedthrough
rlabel pdiffusion 318 -1171 318 -1171 0 feedthrough
rlabel pdiffusion 325 -1171 325 -1171 0 feedthrough
rlabel pdiffusion 332 -1171 332 -1171 0 feedthrough
rlabel pdiffusion 339 -1171 339 -1171 0 feedthrough
rlabel pdiffusion 346 -1171 346 -1171 0 feedthrough
rlabel pdiffusion 353 -1171 353 -1171 0 feedthrough
rlabel pdiffusion 360 -1171 360 -1171 0 feedthrough
rlabel pdiffusion 367 -1171 367 -1171 0 feedthrough
rlabel pdiffusion 374 -1171 374 -1171 0 feedthrough
rlabel pdiffusion 381 -1171 381 -1171 0 feedthrough
rlabel pdiffusion 388 -1171 388 -1171 0 feedthrough
rlabel pdiffusion 395 -1171 395 -1171 0 feedthrough
rlabel pdiffusion 402 -1171 402 -1171 0 feedthrough
rlabel pdiffusion 409 -1171 409 -1171 0 feedthrough
rlabel pdiffusion 416 -1171 416 -1171 0 feedthrough
rlabel pdiffusion 423 -1171 423 -1171 0 cellNo=439
rlabel pdiffusion 430 -1171 430 -1171 0 cellNo=245
rlabel pdiffusion 437 -1171 437 -1171 0 feedthrough
rlabel pdiffusion 444 -1171 444 -1171 0 feedthrough
rlabel pdiffusion 451 -1171 451 -1171 0 feedthrough
rlabel pdiffusion 458 -1171 458 -1171 0 feedthrough
rlabel pdiffusion 465 -1171 465 -1171 0 feedthrough
rlabel pdiffusion 472 -1171 472 -1171 0 feedthrough
rlabel pdiffusion 479 -1171 479 -1171 0 feedthrough
rlabel pdiffusion 486 -1171 486 -1171 0 feedthrough
rlabel pdiffusion 493 -1171 493 -1171 0 feedthrough
rlabel pdiffusion 500 -1171 500 -1171 0 feedthrough
rlabel pdiffusion 507 -1171 507 -1171 0 cellNo=831
rlabel pdiffusion 514 -1171 514 -1171 0 feedthrough
rlabel pdiffusion 521 -1171 521 -1171 0 feedthrough
rlabel pdiffusion 528 -1171 528 -1171 0 feedthrough
rlabel pdiffusion 535 -1171 535 -1171 0 feedthrough
rlabel pdiffusion 542 -1171 542 -1171 0 feedthrough
rlabel pdiffusion 549 -1171 549 -1171 0 feedthrough
rlabel pdiffusion 556 -1171 556 -1171 0 feedthrough
rlabel pdiffusion 563 -1171 563 -1171 0 feedthrough
rlabel pdiffusion 570 -1171 570 -1171 0 feedthrough
rlabel pdiffusion 577 -1171 577 -1171 0 feedthrough
rlabel pdiffusion 584 -1171 584 -1171 0 feedthrough
rlabel pdiffusion 591 -1171 591 -1171 0 cellNo=597
rlabel pdiffusion 598 -1171 598 -1171 0 feedthrough
rlabel pdiffusion 605 -1171 605 -1171 0 cellNo=110
rlabel pdiffusion 612 -1171 612 -1171 0 feedthrough
rlabel pdiffusion 619 -1171 619 -1171 0 feedthrough
rlabel pdiffusion 626 -1171 626 -1171 0 feedthrough
rlabel pdiffusion 633 -1171 633 -1171 0 feedthrough
rlabel pdiffusion 640 -1171 640 -1171 0 feedthrough
rlabel pdiffusion 647 -1171 647 -1171 0 feedthrough
rlabel pdiffusion 654 -1171 654 -1171 0 cellNo=70
rlabel pdiffusion 661 -1171 661 -1171 0 feedthrough
rlabel pdiffusion 668 -1171 668 -1171 0 feedthrough
rlabel pdiffusion 675 -1171 675 -1171 0 feedthrough
rlabel pdiffusion 682 -1171 682 -1171 0 feedthrough
rlabel pdiffusion 689 -1171 689 -1171 0 feedthrough
rlabel pdiffusion 696 -1171 696 -1171 0 feedthrough
rlabel pdiffusion 703 -1171 703 -1171 0 feedthrough
rlabel pdiffusion 710 -1171 710 -1171 0 feedthrough
rlabel pdiffusion 717 -1171 717 -1171 0 feedthrough
rlabel pdiffusion 724 -1171 724 -1171 0 feedthrough
rlabel pdiffusion 731 -1171 731 -1171 0 cellNo=101
rlabel pdiffusion 738 -1171 738 -1171 0 feedthrough
rlabel pdiffusion 745 -1171 745 -1171 0 feedthrough
rlabel pdiffusion 752 -1171 752 -1171 0 feedthrough
rlabel pdiffusion 759 -1171 759 -1171 0 cellNo=336
rlabel pdiffusion 766 -1171 766 -1171 0 feedthrough
rlabel pdiffusion 773 -1171 773 -1171 0 cellNo=450
rlabel pdiffusion 780 -1171 780 -1171 0 feedthrough
rlabel pdiffusion 787 -1171 787 -1171 0 feedthrough
rlabel pdiffusion 794 -1171 794 -1171 0 feedthrough
rlabel pdiffusion 801 -1171 801 -1171 0 feedthrough
rlabel pdiffusion 808 -1171 808 -1171 0 feedthrough
rlabel pdiffusion 815 -1171 815 -1171 0 feedthrough
rlabel pdiffusion 822 -1171 822 -1171 0 cellNo=294
rlabel pdiffusion 829 -1171 829 -1171 0 feedthrough
rlabel pdiffusion 836 -1171 836 -1171 0 feedthrough
rlabel pdiffusion 843 -1171 843 -1171 0 feedthrough
rlabel pdiffusion 850 -1171 850 -1171 0 cellNo=556
rlabel pdiffusion 857 -1171 857 -1171 0 feedthrough
rlabel pdiffusion 864 -1171 864 -1171 0 cellNo=638
rlabel pdiffusion 871 -1171 871 -1171 0 feedthrough
rlabel pdiffusion 878 -1171 878 -1171 0 cellNo=526
rlabel pdiffusion 885 -1171 885 -1171 0 feedthrough
rlabel pdiffusion 892 -1171 892 -1171 0 feedthrough
rlabel pdiffusion 899 -1171 899 -1171 0 feedthrough
rlabel pdiffusion 906 -1171 906 -1171 0 cellNo=129
rlabel pdiffusion 913 -1171 913 -1171 0 feedthrough
rlabel pdiffusion 920 -1171 920 -1171 0 feedthrough
rlabel pdiffusion 927 -1171 927 -1171 0 feedthrough
rlabel pdiffusion 934 -1171 934 -1171 0 feedthrough
rlabel pdiffusion 941 -1171 941 -1171 0 feedthrough
rlabel pdiffusion 948 -1171 948 -1171 0 cellNo=93
rlabel pdiffusion 955 -1171 955 -1171 0 cellNo=971
rlabel pdiffusion 962 -1171 962 -1171 0 cellNo=645
rlabel pdiffusion 969 -1171 969 -1171 0 feedthrough
rlabel pdiffusion 976 -1171 976 -1171 0 feedthrough
rlabel pdiffusion 983 -1171 983 -1171 0 feedthrough
rlabel pdiffusion 990 -1171 990 -1171 0 feedthrough
rlabel pdiffusion 997 -1171 997 -1171 0 feedthrough
rlabel pdiffusion 1004 -1171 1004 -1171 0 cellNo=174
rlabel pdiffusion 1011 -1171 1011 -1171 0 feedthrough
rlabel pdiffusion 1018 -1171 1018 -1171 0 feedthrough
rlabel pdiffusion 1025 -1171 1025 -1171 0 feedthrough
rlabel pdiffusion 1032 -1171 1032 -1171 0 feedthrough
rlabel pdiffusion 1039 -1171 1039 -1171 0 feedthrough
rlabel pdiffusion 1046 -1171 1046 -1171 0 cellNo=72
rlabel pdiffusion 1053 -1171 1053 -1171 0 feedthrough
rlabel pdiffusion 1060 -1171 1060 -1171 0 feedthrough
rlabel pdiffusion 1067 -1171 1067 -1171 0 feedthrough
rlabel pdiffusion 1074 -1171 1074 -1171 0 feedthrough
rlabel pdiffusion 1081 -1171 1081 -1171 0 feedthrough
rlabel pdiffusion 1088 -1171 1088 -1171 0 feedthrough
rlabel pdiffusion 1095 -1171 1095 -1171 0 feedthrough
rlabel pdiffusion 1102 -1171 1102 -1171 0 feedthrough
rlabel pdiffusion 1109 -1171 1109 -1171 0 feedthrough
rlabel pdiffusion 1116 -1171 1116 -1171 0 feedthrough
rlabel pdiffusion 1123 -1171 1123 -1171 0 feedthrough
rlabel pdiffusion 1130 -1171 1130 -1171 0 feedthrough
rlabel pdiffusion 1137 -1171 1137 -1171 0 feedthrough
rlabel pdiffusion 1144 -1171 1144 -1171 0 feedthrough
rlabel pdiffusion 1151 -1171 1151 -1171 0 feedthrough
rlabel pdiffusion 1158 -1171 1158 -1171 0 cellNo=141
rlabel pdiffusion 1165 -1171 1165 -1171 0 cellNo=89
rlabel pdiffusion 1172 -1171 1172 -1171 0 feedthrough
rlabel pdiffusion 1179 -1171 1179 -1171 0 cellNo=8
rlabel pdiffusion 1186 -1171 1186 -1171 0 feedthrough
rlabel pdiffusion 1193 -1171 1193 -1171 0 feedthrough
rlabel pdiffusion 1200 -1171 1200 -1171 0 cellNo=331
rlabel pdiffusion 1207 -1171 1207 -1171 0 feedthrough
rlabel pdiffusion 1214 -1171 1214 -1171 0 feedthrough
rlabel pdiffusion 1221 -1171 1221 -1171 0 cellNo=622
rlabel pdiffusion 1228 -1171 1228 -1171 0 feedthrough
rlabel pdiffusion 1235 -1171 1235 -1171 0 cellNo=560
rlabel pdiffusion 1242 -1171 1242 -1171 0 feedthrough
rlabel pdiffusion 1249 -1171 1249 -1171 0 feedthrough
rlabel pdiffusion 1256 -1171 1256 -1171 0 feedthrough
rlabel pdiffusion 1263 -1171 1263 -1171 0 feedthrough
rlabel pdiffusion 1270 -1171 1270 -1171 0 feedthrough
rlabel pdiffusion 1277 -1171 1277 -1171 0 feedthrough
rlabel pdiffusion 1284 -1171 1284 -1171 0 feedthrough
rlabel pdiffusion 1291 -1171 1291 -1171 0 feedthrough
rlabel pdiffusion 1298 -1171 1298 -1171 0 feedthrough
rlabel pdiffusion 1305 -1171 1305 -1171 0 cellNo=409
rlabel pdiffusion 1312 -1171 1312 -1171 0 feedthrough
rlabel pdiffusion 1319 -1171 1319 -1171 0 feedthrough
rlabel pdiffusion 1326 -1171 1326 -1171 0 feedthrough
rlabel pdiffusion 1333 -1171 1333 -1171 0 cellNo=464
rlabel pdiffusion 1340 -1171 1340 -1171 0 feedthrough
rlabel pdiffusion 1347 -1171 1347 -1171 0 feedthrough
rlabel pdiffusion 1354 -1171 1354 -1171 0 feedthrough
rlabel pdiffusion 1361 -1171 1361 -1171 0 feedthrough
rlabel pdiffusion 1368 -1171 1368 -1171 0 feedthrough
rlabel pdiffusion 1375 -1171 1375 -1171 0 feedthrough
rlabel pdiffusion 1382 -1171 1382 -1171 0 feedthrough
rlabel pdiffusion 1389 -1171 1389 -1171 0 feedthrough
rlabel pdiffusion 1396 -1171 1396 -1171 0 feedthrough
rlabel pdiffusion 1403 -1171 1403 -1171 0 feedthrough
rlabel pdiffusion 1410 -1171 1410 -1171 0 feedthrough
rlabel pdiffusion 1417 -1171 1417 -1171 0 feedthrough
rlabel pdiffusion 1424 -1171 1424 -1171 0 feedthrough
rlabel pdiffusion 1431 -1171 1431 -1171 0 feedthrough
rlabel pdiffusion 1438 -1171 1438 -1171 0 feedthrough
rlabel pdiffusion 1445 -1171 1445 -1171 0 cellNo=462
rlabel pdiffusion 1452 -1171 1452 -1171 0 feedthrough
rlabel pdiffusion 1459 -1171 1459 -1171 0 feedthrough
rlabel pdiffusion 1466 -1171 1466 -1171 0 feedthrough
rlabel pdiffusion 1473 -1171 1473 -1171 0 feedthrough
rlabel pdiffusion 1480 -1171 1480 -1171 0 feedthrough
rlabel pdiffusion 1487 -1171 1487 -1171 0 feedthrough
rlabel pdiffusion 1494 -1171 1494 -1171 0 feedthrough
rlabel pdiffusion 1501 -1171 1501 -1171 0 feedthrough
rlabel pdiffusion 1508 -1171 1508 -1171 0 feedthrough
rlabel pdiffusion 1515 -1171 1515 -1171 0 feedthrough
rlabel pdiffusion 1522 -1171 1522 -1171 0 feedthrough
rlabel pdiffusion 1529 -1171 1529 -1171 0 feedthrough
rlabel pdiffusion 1536 -1171 1536 -1171 0 feedthrough
rlabel pdiffusion 1543 -1171 1543 -1171 0 feedthrough
rlabel pdiffusion 1550 -1171 1550 -1171 0 cellNo=780
rlabel pdiffusion 1557 -1171 1557 -1171 0 feedthrough
rlabel pdiffusion 1564 -1171 1564 -1171 0 feedthrough
rlabel pdiffusion 1571 -1171 1571 -1171 0 feedthrough
rlabel pdiffusion 1578 -1171 1578 -1171 0 feedthrough
rlabel pdiffusion 1585 -1171 1585 -1171 0 feedthrough
rlabel pdiffusion 1592 -1171 1592 -1171 0 feedthrough
rlabel pdiffusion 1599 -1171 1599 -1171 0 feedthrough
rlabel pdiffusion 1606 -1171 1606 -1171 0 feedthrough
rlabel pdiffusion 1613 -1171 1613 -1171 0 feedthrough
rlabel pdiffusion 1620 -1171 1620 -1171 0 feedthrough
rlabel pdiffusion 1627 -1171 1627 -1171 0 feedthrough
rlabel pdiffusion 1634 -1171 1634 -1171 0 feedthrough
rlabel pdiffusion 1641 -1171 1641 -1171 0 feedthrough
rlabel pdiffusion 1648 -1171 1648 -1171 0 feedthrough
rlabel pdiffusion 1655 -1171 1655 -1171 0 feedthrough
rlabel pdiffusion 1662 -1171 1662 -1171 0 feedthrough
rlabel pdiffusion 1669 -1171 1669 -1171 0 feedthrough
rlabel pdiffusion 1676 -1171 1676 -1171 0 feedthrough
rlabel pdiffusion 1683 -1171 1683 -1171 0 feedthrough
rlabel pdiffusion 1690 -1171 1690 -1171 0 feedthrough
rlabel pdiffusion 1697 -1171 1697 -1171 0 feedthrough
rlabel pdiffusion 1704 -1171 1704 -1171 0 feedthrough
rlabel pdiffusion 1711 -1171 1711 -1171 0 feedthrough
rlabel pdiffusion 1718 -1171 1718 -1171 0 feedthrough
rlabel pdiffusion 1725 -1171 1725 -1171 0 feedthrough
rlabel pdiffusion 1732 -1171 1732 -1171 0 feedthrough
rlabel pdiffusion 1739 -1171 1739 -1171 0 cellNo=538
rlabel pdiffusion 1746 -1171 1746 -1171 0 feedthrough
rlabel pdiffusion 1753 -1171 1753 -1171 0 feedthrough
rlabel pdiffusion 1760 -1171 1760 -1171 0 feedthrough
rlabel pdiffusion 1767 -1171 1767 -1171 0 feedthrough
rlabel pdiffusion 1774 -1171 1774 -1171 0 feedthrough
rlabel pdiffusion 1781 -1171 1781 -1171 0 feedthrough
rlabel pdiffusion 1788 -1171 1788 -1171 0 feedthrough
rlabel pdiffusion 1795 -1171 1795 -1171 0 feedthrough
rlabel pdiffusion 1802 -1171 1802 -1171 0 feedthrough
rlabel pdiffusion 1809 -1171 1809 -1171 0 feedthrough
rlabel pdiffusion 1816 -1171 1816 -1171 0 feedthrough
rlabel pdiffusion 1823 -1171 1823 -1171 0 feedthrough
rlabel pdiffusion 1830 -1171 1830 -1171 0 feedthrough
rlabel pdiffusion 1837 -1171 1837 -1171 0 feedthrough
rlabel pdiffusion 1844 -1171 1844 -1171 0 feedthrough
rlabel pdiffusion 1851 -1171 1851 -1171 0 feedthrough
rlabel pdiffusion 1858 -1171 1858 -1171 0 feedthrough
rlabel pdiffusion 1865 -1171 1865 -1171 0 feedthrough
rlabel pdiffusion 1872 -1171 1872 -1171 0 feedthrough
rlabel pdiffusion 1879 -1171 1879 -1171 0 feedthrough
rlabel pdiffusion 1886 -1171 1886 -1171 0 feedthrough
rlabel pdiffusion 1893 -1171 1893 -1171 0 feedthrough
rlabel pdiffusion 1900 -1171 1900 -1171 0 feedthrough
rlabel pdiffusion 1907 -1171 1907 -1171 0 feedthrough
rlabel pdiffusion 1914 -1171 1914 -1171 0 feedthrough
rlabel pdiffusion 1921 -1171 1921 -1171 0 feedthrough
rlabel pdiffusion 1928 -1171 1928 -1171 0 feedthrough
rlabel pdiffusion 1935 -1171 1935 -1171 0 feedthrough
rlabel pdiffusion 1942 -1171 1942 -1171 0 feedthrough
rlabel pdiffusion 1949 -1171 1949 -1171 0 feedthrough
rlabel pdiffusion 1956 -1171 1956 -1171 0 feedthrough
rlabel pdiffusion 1963 -1171 1963 -1171 0 feedthrough
rlabel pdiffusion 1970 -1171 1970 -1171 0 feedthrough
rlabel pdiffusion 1977 -1171 1977 -1171 0 feedthrough
rlabel pdiffusion 1984 -1171 1984 -1171 0 feedthrough
rlabel pdiffusion 1991 -1171 1991 -1171 0 feedthrough
rlabel pdiffusion 1998 -1171 1998 -1171 0 feedthrough
rlabel pdiffusion 2005 -1171 2005 -1171 0 feedthrough
rlabel pdiffusion 2012 -1171 2012 -1171 0 feedthrough
rlabel pdiffusion 2019 -1171 2019 -1171 0 feedthrough
rlabel pdiffusion 2026 -1171 2026 -1171 0 feedthrough
rlabel pdiffusion 2033 -1171 2033 -1171 0 feedthrough
rlabel pdiffusion 2040 -1171 2040 -1171 0 feedthrough
rlabel pdiffusion 2047 -1171 2047 -1171 0 feedthrough
rlabel pdiffusion 2054 -1171 2054 -1171 0 feedthrough
rlabel pdiffusion 2061 -1171 2061 -1171 0 feedthrough
rlabel pdiffusion 2068 -1171 2068 -1171 0 feedthrough
rlabel pdiffusion 2075 -1171 2075 -1171 0 feedthrough
rlabel pdiffusion 2082 -1171 2082 -1171 0 feedthrough
rlabel pdiffusion 2089 -1171 2089 -1171 0 feedthrough
rlabel pdiffusion 2096 -1171 2096 -1171 0 feedthrough
rlabel pdiffusion 2103 -1171 2103 -1171 0 feedthrough
rlabel pdiffusion 2110 -1171 2110 -1171 0 feedthrough
rlabel pdiffusion 2117 -1171 2117 -1171 0 feedthrough
rlabel pdiffusion 2124 -1171 2124 -1171 0 feedthrough
rlabel pdiffusion 2131 -1171 2131 -1171 0 feedthrough
rlabel pdiffusion 2138 -1171 2138 -1171 0 feedthrough
rlabel pdiffusion 2145 -1171 2145 -1171 0 feedthrough
rlabel pdiffusion 2152 -1171 2152 -1171 0 feedthrough
rlabel pdiffusion 2159 -1171 2159 -1171 0 feedthrough
rlabel pdiffusion 2166 -1171 2166 -1171 0 feedthrough
rlabel pdiffusion 2173 -1171 2173 -1171 0 feedthrough
rlabel pdiffusion 2180 -1171 2180 -1171 0 feedthrough
rlabel pdiffusion 2187 -1171 2187 -1171 0 feedthrough
rlabel pdiffusion 2194 -1171 2194 -1171 0 feedthrough
rlabel pdiffusion 2201 -1171 2201 -1171 0 feedthrough
rlabel pdiffusion 2208 -1171 2208 -1171 0 feedthrough
rlabel pdiffusion 2215 -1171 2215 -1171 0 feedthrough
rlabel pdiffusion 2222 -1171 2222 -1171 0 feedthrough
rlabel pdiffusion 2229 -1171 2229 -1171 0 feedthrough
rlabel pdiffusion 2236 -1171 2236 -1171 0 feedthrough
rlabel pdiffusion 2243 -1171 2243 -1171 0 feedthrough
rlabel pdiffusion 2250 -1171 2250 -1171 0 feedthrough
rlabel pdiffusion 2257 -1171 2257 -1171 0 feedthrough
rlabel pdiffusion 2264 -1171 2264 -1171 0 feedthrough
rlabel pdiffusion 2271 -1171 2271 -1171 0 feedthrough
rlabel pdiffusion 2278 -1171 2278 -1171 0 feedthrough
rlabel pdiffusion 2285 -1171 2285 -1171 0 feedthrough
rlabel pdiffusion 2292 -1171 2292 -1171 0 feedthrough
rlabel pdiffusion 2299 -1171 2299 -1171 0 feedthrough
rlabel pdiffusion 2306 -1171 2306 -1171 0 feedthrough
rlabel pdiffusion 2313 -1171 2313 -1171 0 feedthrough
rlabel pdiffusion 2320 -1171 2320 -1171 0 feedthrough
rlabel pdiffusion 2327 -1171 2327 -1171 0 feedthrough
rlabel pdiffusion 2334 -1171 2334 -1171 0 feedthrough
rlabel pdiffusion 2341 -1171 2341 -1171 0 feedthrough
rlabel pdiffusion 2348 -1171 2348 -1171 0 feedthrough
rlabel pdiffusion 2355 -1171 2355 -1171 0 feedthrough
rlabel pdiffusion 2362 -1171 2362 -1171 0 feedthrough
rlabel pdiffusion 2369 -1171 2369 -1171 0 feedthrough
rlabel pdiffusion 2376 -1171 2376 -1171 0 feedthrough
rlabel pdiffusion 2383 -1171 2383 -1171 0 feedthrough
rlabel pdiffusion 2390 -1171 2390 -1171 0 cellNo=434
rlabel pdiffusion 2397 -1171 2397 -1171 0 cellNo=269
rlabel pdiffusion 2404 -1171 2404 -1171 0 feedthrough
rlabel pdiffusion 2425 -1171 2425 -1171 0 feedthrough
rlabel pdiffusion 2432 -1171 2432 -1171 0 feedthrough
rlabel pdiffusion 2439 -1171 2439 -1171 0 feedthrough
rlabel pdiffusion 3 -1354 3 -1354 0 cellNo=470
rlabel pdiffusion 10 -1354 10 -1354 0 feedthrough
rlabel pdiffusion 17 -1354 17 -1354 0 cellNo=231
rlabel pdiffusion 24 -1354 24 -1354 0 feedthrough
rlabel pdiffusion 31 -1354 31 -1354 0 feedthrough
rlabel pdiffusion 38 -1354 38 -1354 0 feedthrough
rlabel pdiffusion 45 -1354 45 -1354 0 feedthrough
rlabel pdiffusion 52 -1354 52 -1354 0 feedthrough
rlabel pdiffusion 59 -1354 59 -1354 0 feedthrough
rlabel pdiffusion 66 -1354 66 -1354 0 feedthrough
rlabel pdiffusion 73 -1354 73 -1354 0 feedthrough
rlabel pdiffusion 80 -1354 80 -1354 0 cellNo=743
rlabel pdiffusion 87 -1354 87 -1354 0 feedthrough
rlabel pdiffusion 94 -1354 94 -1354 0 feedthrough
rlabel pdiffusion 101 -1354 101 -1354 0 feedthrough
rlabel pdiffusion 108 -1354 108 -1354 0 feedthrough
rlabel pdiffusion 115 -1354 115 -1354 0 feedthrough
rlabel pdiffusion 122 -1354 122 -1354 0 cellNo=580
rlabel pdiffusion 129 -1354 129 -1354 0 feedthrough
rlabel pdiffusion 136 -1354 136 -1354 0 feedthrough
rlabel pdiffusion 143 -1354 143 -1354 0 feedthrough
rlabel pdiffusion 150 -1354 150 -1354 0 feedthrough
rlabel pdiffusion 157 -1354 157 -1354 0 feedthrough
rlabel pdiffusion 164 -1354 164 -1354 0 feedthrough
rlabel pdiffusion 171 -1354 171 -1354 0 feedthrough
rlabel pdiffusion 178 -1354 178 -1354 0 feedthrough
rlabel pdiffusion 185 -1354 185 -1354 0 feedthrough
rlabel pdiffusion 192 -1354 192 -1354 0 feedthrough
rlabel pdiffusion 199 -1354 199 -1354 0 feedthrough
rlabel pdiffusion 206 -1354 206 -1354 0 cellNo=806
rlabel pdiffusion 213 -1354 213 -1354 0 feedthrough
rlabel pdiffusion 220 -1354 220 -1354 0 feedthrough
rlabel pdiffusion 227 -1354 227 -1354 0 cellNo=490
rlabel pdiffusion 234 -1354 234 -1354 0 feedthrough
rlabel pdiffusion 241 -1354 241 -1354 0 feedthrough
rlabel pdiffusion 248 -1354 248 -1354 0 cellNo=396
rlabel pdiffusion 255 -1354 255 -1354 0 cellNo=374
rlabel pdiffusion 262 -1354 262 -1354 0 feedthrough
rlabel pdiffusion 269 -1354 269 -1354 0 cellNo=808
rlabel pdiffusion 276 -1354 276 -1354 0 feedthrough
rlabel pdiffusion 283 -1354 283 -1354 0 feedthrough
rlabel pdiffusion 290 -1354 290 -1354 0 feedthrough
rlabel pdiffusion 297 -1354 297 -1354 0 feedthrough
rlabel pdiffusion 304 -1354 304 -1354 0 feedthrough
rlabel pdiffusion 311 -1354 311 -1354 0 feedthrough
rlabel pdiffusion 318 -1354 318 -1354 0 feedthrough
rlabel pdiffusion 325 -1354 325 -1354 0 feedthrough
rlabel pdiffusion 332 -1354 332 -1354 0 feedthrough
rlabel pdiffusion 339 -1354 339 -1354 0 feedthrough
rlabel pdiffusion 346 -1354 346 -1354 0 feedthrough
rlabel pdiffusion 353 -1354 353 -1354 0 feedthrough
rlabel pdiffusion 360 -1354 360 -1354 0 feedthrough
rlabel pdiffusion 367 -1354 367 -1354 0 feedthrough
rlabel pdiffusion 374 -1354 374 -1354 0 feedthrough
rlabel pdiffusion 381 -1354 381 -1354 0 feedthrough
rlabel pdiffusion 388 -1354 388 -1354 0 feedthrough
rlabel pdiffusion 395 -1354 395 -1354 0 feedthrough
rlabel pdiffusion 402 -1354 402 -1354 0 feedthrough
rlabel pdiffusion 409 -1354 409 -1354 0 feedthrough
rlabel pdiffusion 416 -1354 416 -1354 0 feedthrough
rlabel pdiffusion 423 -1354 423 -1354 0 feedthrough
rlabel pdiffusion 430 -1354 430 -1354 0 feedthrough
rlabel pdiffusion 437 -1354 437 -1354 0 feedthrough
rlabel pdiffusion 444 -1354 444 -1354 0 feedthrough
rlabel pdiffusion 451 -1354 451 -1354 0 feedthrough
rlabel pdiffusion 458 -1354 458 -1354 0 feedthrough
rlabel pdiffusion 465 -1354 465 -1354 0 feedthrough
rlabel pdiffusion 472 -1354 472 -1354 0 feedthrough
rlabel pdiffusion 479 -1354 479 -1354 0 feedthrough
rlabel pdiffusion 486 -1354 486 -1354 0 feedthrough
rlabel pdiffusion 493 -1354 493 -1354 0 feedthrough
rlabel pdiffusion 500 -1354 500 -1354 0 feedthrough
rlabel pdiffusion 507 -1354 507 -1354 0 feedthrough
rlabel pdiffusion 514 -1354 514 -1354 0 feedthrough
rlabel pdiffusion 521 -1354 521 -1354 0 feedthrough
rlabel pdiffusion 528 -1354 528 -1354 0 feedthrough
rlabel pdiffusion 535 -1354 535 -1354 0 feedthrough
rlabel pdiffusion 542 -1354 542 -1354 0 feedthrough
rlabel pdiffusion 549 -1354 549 -1354 0 feedthrough
rlabel pdiffusion 556 -1354 556 -1354 0 feedthrough
rlabel pdiffusion 563 -1354 563 -1354 0 feedthrough
rlabel pdiffusion 570 -1354 570 -1354 0 feedthrough
rlabel pdiffusion 577 -1354 577 -1354 0 feedthrough
rlabel pdiffusion 584 -1354 584 -1354 0 feedthrough
rlabel pdiffusion 591 -1354 591 -1354 0 feedthrough
rlabel pdiffusion 598 -1354 598 -1354 0 feedthrough
rlabel pdiffusion 605 -1354 605 -1354 0 cellNo=794
rlabel pdiffusion 612 -1354 612 -1354 0 feedthrough
rlabel pdiffusion 619 -1354 619 -1354 0 feedthrough
rlabel pdiffusion 626 -1354 626 -1354 0 feedthrough
rlabel pdiffusion 633 -1354 633 -1354 0 feedthrough
rlabel pdiffusion 640 -1354 640 -1354 0 cellNo=720
rlabel pdiffusion 647 -1354 647 -1354 0 feedthrough
rlabel pdiffusion 654 -1354 654 -1354 0 feedthrough
rlabel pdiffusion 661 -1354 661 -1354 0 feedthrough
rlabel pdiffusion 668 -1354 668 -1354 0 feedthrough
rlabel pdiffusion 675 -1354 675 -1354 0 cellNo=60
rlabel pdiffusion 682 -1354 682 -1354 0 feedthrough
rlabel pdiffusion 689 -1354 689 -1354 0 feedthrough
rlabel pdiffusion 696 -1354 696 -1354 0 feedthrough
rlabel pdiffusion 703 -1354 703 -1354 0 feedthrough
rlabel pdiffusion 710 -1354 710 -1354 0 feedthrough
rlabel pdiffusion 717 -1354 717 -1354 0 feedthrough
rlabel pdiffusion 724 -1354 724 -1354 0 cellNo=542
rlabel pdiffusion 731 -1354 731 -1354 0 feedthrough
rlabel pdiffusion 738 -1354 738 -1354 0 feedthrough
rlabel pdiffusion 745 -1354 745 -1354 0 feedthrough
rlabel pdiffusion 752 -1354 752 -1354 0 feedthrough
rlabel pdiffusion 759 -1354 759 -1354 0 feedthrough
rlabel pdiffusion 766 -1354 766 -1354 0 feedthrough
rlabel pdiffusion 773 -1354 773 -1354 0 feedthrough
rlabel pdiffusion 780 -1354 780 -1354 0 cellNo=65
rlabel pdiffusion 787 -1354 787 -1354 0 cellNo=637
rlabel pdiffusion 794 -1354 794 -1354 0 cellNo=41
rlabel pdiffusion 801 -1354 801 -1354 0 feedthrough
rlabel pdiffusion 808 -1354 808 -1354 0 feedthrough
rlabel pdiffusion 815 -1354 815 -1354 0 feedthrough
rlabel pdiffusion 822 -1354 822 -1354 0 feedthrough
rlabel pdiffusion 829 -1354 829 -1354 0 cellNo=552
rlabel pdiffusion 836 -1354 836 -1354 0 cellNo=551
rlabel pdiffusion 843 -1354 843 -1354 0 feedthrough
rlabel pdiffusion 850 -1354 850 -1354 0 feedthrough
rlabel pdiffusion 857 -1354 857 -1354 0 feedthrough
rlabel pdiffusion 864 -1354 864 -1354 0 cellNo=451
rlabel pdiffusion 871 -1354 871 -1354 0 feedthrough
rlabel pdiffusion 878 -1354 878 -1354 0 cellNo=166
rlabel pdiffusion 885 -1354 885 -1354 0 feedthrough
rlabel pdiffusion 892 -1354 892 -1354 0 cellNo=139
rlabel pdiffusion 899 -1354 899 -1354 0 feedthrough
rlabel pdiffusion 906 -1354 906 -1354 0 feedthrough
rlabel pdiffusion 913 -1354 913 -1354 0 feedthrough
rlabel pdiffusion 920 -1354 920 -1354 0 feedthrough
rlabel pdiffusion 927 -1354 927 -1354 0 feedthrough
rlabel pdiffusion 934 -1354 934 -1354 0 feedthrough
rlabel pdiffusion 941 -1354 941 -1354 0 feedthrough
rlabel pdiffusion 948 -1354 948 -1354 0 feedthrough
rlabel pdiffusion 955 -1354 955 -1354 0 cellNo=313
rlabel pdiffusion 962 -1354 962 -1354 0 feedthrough
rlabel pdiffusion 969 -1354 969 -1354 0 feedthrough
rlabel pdiffusion 976 -1354 976 -1354 0 feedthrough
rlabel pdiffusion 983 -1354 983 -1354 0 cellNo=944
rlabel pdiffusion 990 -1354 990 -1354 0 cellNo=256
rlabel pdiffusion 997 -1354 997 -1354 0 cellNo=852
rlabel pdiffusion 1004 -1354 1004 -1354 0 cellNo=58
rlabel pdiffusion 1011 -1354 1011 -1354 0 cellNo=740
rlabel pdiffusion 1018 -1354 1018 -1354 0 feedthrough
rlabel pdiffusion 1025 -1354 1025 -1354 0 feedthrough
rlabel pdiffusion 1032 -1354 1032 -1354 0 feedthrough
rlabel pdiffusion 1039 -1354 1039 -1354 0 cellNo=504
rlabel pdiffusion 1046 -1354 1046 -1354 0 feedthrough
rlabel pdiffusion 1053 -1354 1053 -1354 0 feedthrough
rlabel pdiffusion 1060 -1354 1060 -1354 0 feedthrough
rlabel pdiffusion 1067 -1354 1067 -1354 0 feedthrough
rlabel pdiffusion 1074 -1354 1074 -1354 0 feedthrough
rlabel pdiffusion 1081 -1354 1081 -1354 0 feedthrough
rlabel pdiffusion 1088 -1354 1088 -1354 0 feedthrough
rlabel pdiffusion 1095 -1354 1095 -1354 0 feedthrough
rlabel pdiffusion 1102 -1354 1102 -1354 0 cellNo=113
rlabel pdiffusion 1109 -1354 1109 -1354 0 feedthrough
rlabel pdiffusion 1116 -1354 1116 -1354 0 feedthrough
rlabel pdiffusion 1123 -1354 1123 -1354 0 feedthrough
rlabel pdiffusion 1130 -1354 1130 -1354 0 feedthrough
rlabel pdiffusion 1137 -1354 1137 -1354 0 feedthrough
rlabel pdiffusion 1144 -1354 1144 -1354 0 feedthrough
rlabel pdiffusion 1151 -1354 1151 -1354 0 cellNo=165
rlabel pdiffusion 1158 -1354 1158 -1354 0 feedthrough
rlabel pdiffusion 1165 -1354 1165 -1354 0 feedthrough
rlabel pdiffusion 1172 -1354 1172 -1354 0 feedthrough
rlabel pdiffusion 1179 -1354 1179 -1354 0 feedthrough
rlabel pdiffusion 1186 -1354 1186 -1354 0 feedthrough
rlabel pdiffusion 1193 -1354 1193 -1354 0 feedthrough
rlabel pdiffusion 1200 -1354 1200 -1354 0 feedthrough
rlabel pdiffusion 1207 -1354 1207 -1354 0 feedthrough
rlabel pdiffusion 1214 -1354 1214 -1354 0 cellNo=805
rlabel pdiffusion 1221 -1354 1221 -1354 0 feedthrough
rlabel pdiffusion 1228 -1354 1228 -1354 0 feedthrough
rlabel pdiffusion 1235 -1354 1235 -1354 0 feedthrough
rlabel pdiffusion 1242 -1354 1242 -1354 0 feedthrough
rlabel pdiffusion 1249 -1354 1249 -1354 0 feedthrough
rlabel pdiffusion 1256 -1354 1256 -1354 0 feedthrough
rlabel pdiffusion 1263 -1354 1263 -1354 0 feedthrough
rlabel pdiffusion 1270 -1354 1270 -1354 0 feedthrough
rlabel pdiffusion 1277 -1354 1277 -1354 0 feedthrough
rlabel pdiffusion 1284 -1354 1284 -1354 0 feedthrough
rlabel pdiffusion 1291 -1354 1291 -1354 0 feedthrough
rlabel pdiffusion 1298 -1354 1298 -1354 0 feedthrough
rlabel pdiffusion 1305 -1354 1305 -1354 0 feedthrough
rlabel pdiffusion 1312 -1354 1312 -1354 0 feedthrough
rlabel pdiffusion 1319 -1354 1319 -1354 0 feedthrough
rlabel pdiffusion 1326 -1354 1326 -1354 0 feedthrough
rlabel pdiffusion 1333 -1354 1333 -1354 0 feedthrough
rlabel pdiffusion 1340 -1354 1340 -1354 0 feedthrough
rlabel pdiffusion 1347 -1354 1347 -1354 0 feedthrough
rlabel pdiffusion 1354 -1354 1354 -1354 0 feedthrough
rlabel pdiffusion 1361 -1354 1361 -1354 0 feedthrough
rlabel pdiffusion 1368 -1354 1368 -1354 0 cellNo=762
rlabel pdiffusion 1375 -1354 1375 -1354 0 feedthrough
rlabel pdiffusion 1382 -1354 1382 -1354 0 cellNo=285
rlabel pdiffusion 1389 -1354 1389 -1354 0 feedthrough
rlabel pdiffusion 1396 -1354 1396 -1354 0 feedthrough
rlabel pdiffusion 1403 -1354 1403 -1354 0 feedthrough
rlabel pdiffusion 1410 -1354 1410 -1354 0 feedthrough
rlabel pdiffusion 1417 -1354 1417 -1354 0 cellNo=19
rlabel pdiffusion 1424 -1354 1424 -1354 0 feedthrough
rlabel pdiffusion 1431 -1354 1431 -1354 0 cellNo=472
rlabel pdiffusion 1438 -1354 1438 -1354 0 feedthrough
rlabel pdiffusion 1445 -1354 1445 -1354 0 cellNo=546
rlabel pdiffusion 1452 -1354 1452 -1354 0 feedthrough
rlabel pdiffusion 1459 -1354 1459 -1354 0 feedthrough
rlabel pdiffusion 1466 -1354 1466 -1354 0 feedthrough
rlabel pdiffusion 1473 -1354 1473 -1354 0 feedthrough
rlabel pdiffusion 1480 -1354 1480 -1354 0 feedthrough
rlabel pdiffusion 1487 -1354 1487 -1354 0 feedthrough
rlabel pdiffusion 1494 -1354 1494 -1354 0 feedthrough
rlabel pdiffusion 1501 -1354 1501 -1354 0 feedthrough
rlabel pdiffusion 1508 -1354 1508 -1354 0 cellNo=190
rlabel pdiffusion 1515 -1354 1515 -1354 0 feedthrough
rlabel pdiffusion 1522 -1354 1522 -1354 0 feedthrough
rlabel pdiffusion 1529 -1354 1529 -1354 0 feedthrough
rlabel pdiffusion 1536 -1354 1536 -1354 0 feedthrough
rlabel pdiffusion 1543 -1354 1543 -1354 0 feedthrough
rlabel pdiffusion 1550 -1354 1550 -1354 0 feedthrough
rlabel pdiffusion 1557 -1354 1557 -1354 0 feedthrough
rlabel pdiffusion 1564 -1354 1564 -1354 0 feedthrough
rlabel pdiffusion 1571 -1354 1571 -1354 0 feedthrough
rlabel pdiffusion 1578 -1354 1578 -1354 0 feedthrough
rlabel pdiffusion 1585 -1354 1585 -1354 0 feedthrough
rlabel pdiffusion 1592 -1354 1592 -1354 0 feedthrough
rlabel pdiffusion 1599 -1354 1599 -1354 0 feedthrough
rlabel pdiffusion 1606 -1354 1606 -1354 0 feedthrough
rlabel pdiffusion 1613 -1354 1613 -1354 0 feedthrough
rlabel pdiffusion 1620 -1354 1620 -1354 0 feedthrough
rlabel pdiffusion 1627 -1354 1627 -1354 0 feedthrough
rlabel pdiffusion 1634 -1354 1634 -1354 0 feedthrough
rlabel pdiffusion 1641 -1354 1641 -1354 0 feedthrough
rlabel pdiffusion 1648 -1354 1648 -1354 0 feedthrough
rlabel pdiffusion 1655 -1354 1655 -1354 0 feedthrough
rlabel pdiffusion 1662 -1354 1662 -1354 0 feedthrough
rlabel pdiffusion 1669 -1354 1669 -1354 0 feedthrough
rlabel pdiffusion 1676 -1354 1676 -1354 0 cellNo=196
rlabel pdiffusion 1683 -1354 1683 -1354 0 feedthrough
rlabel pdiffusion 1690 -1354 1690 -1354 0 feedthrough
rlabel pdiffusion 1697 -1354 1697 -1354 0 feedthrough
rlabel pdiffusion 1704 -1354 1704 -1354 0 feedthrough
rlabel pdiffusion 1711 -1354 1711 -1354 0 feedthrough
rlabel pdiffusion 1718 -1354 1718 -1354 0 feedthrough
rlabel pdiffusion 1725 -1354 1725 -1354 0 feedthrough
rlabel pdiffusion 1732 -1354 1732 -1354 0 feedthrough
rlabel pdiffusion 1739 -1354 1739 -1354 0 feedthrough
rlabel pdiffusion 1746 -1354 1746 -1354 0 feedthrough
rlabel pdiffusion 1753 -1354 1753 -1354 0 feedthrough
rlabel pdiffusion 1760 -1354 1760 -1354 0 feedthrough
rlabel pdiffusion 1767 -1354 1767 -1354 0 feedthrough
rlabel pdiffusion 1774 -1354 1774 -1354 0 feedthrough
rlabel pdiffusion 1781 -1354 1781 -1354 0 feedthrough
rlabel pdiffusion 1788 -1354 1788 -1354 0 feedthrough
rlabel pdiffusion 1795 -1354 1795 -1354 0 feedthrough
rlabel pdiffusion 1802 -1354 1802 -1354 0 feedthrough
rlabel pdiffusion 1809 -1354 1809 -1354 0 feedthrough
rlabel pdiffusion 1816 -1354 1816 -1354 0 feedthrough
rlabel pdiffusion 1823 -1354 1823 -1354 0 feedthrough
rlabel pdiffusion 1830 -1354 1830 -1354 0 feedthrough
rlabel pdiffusion 1837 -1354 1837 -1354 0 feedthrough
rlabel pdiffusion 1844 -1354 1844 -1354 0 feedthrough
rlabel pdiffusion 1851 -1354 1851 -1354 0 feedthrough
rlabel pdiffusion 1858 -1354 1858 -1354 0 feedthrough
rlabel pdiffusion 1865 -1354 1865 -1354 0 feedthrough
rlabel pdiffusion 1872 -1354 1872 -1354 0 feedthrough
rlabel pdiffusion 1879 -1354 1879 -1354 0 feedthrough
rlabel pdiffusion 1886 -1354 1886 -1354 0 feedthrough
rlabel pdiffusion 1893 -1354 1893 -1354 0 feedthrough
rlabel pdiffusion 1900 -1354 1900 -1354 0 feedthrough
rlabel pdiffusion 1907 -1354 1907 -1354 0 feedthrough
rlabel pdiffusion 1914 -1354 1914 -1354 0 feedthrough
rlabel pdiffusion 1921 -1354 1921 -1354 0 feedthrough
rlabel pdiffusion 1928 -1354 1928 -1354 0 feedthrough
rlabel pdiffusion 1935 -1354 1935 -1354 0 feedthrough
rlabel pdiffusion 1942 -1354 1942 -1354 0 feedthrough
rlabel pdiffusion 1949 -1354 1949 -1354 0 feedthrough
rlabel pdiffusion 1956 -1354 1956 -1354 0 feedthrough
rlabel pdiffusion 1963 -1354 1963 -1354 0 feedthrough
rlabel pdiffusion 1970 -1354 1970 -1354 0 feedthrough
rlabel pdiffusion 1977 -1354 1977 -1354 0 feedthrough
rlabel pdiffusion 1984 -1354 1984 -1354 0 feedthrough
rlabel pdiffusion 1991 -1354 1991 -1354 0 feedthrough
rlabel pdiffusion 1998 -1354 1998 -1354 0 feedthrough
rlabel pdiffusion 2005 -1354 2005 -1354 0 feedthrough
rlabel pdiffusion 2012 -1354 2012 -1354 0 feedthrough
rlabel pdiffusion 2019 -1354 2019 -1354 0 feedthrough
rlabel pdiffusion 2026 -1354 2026 -1354 0 feedthrough
rlabel pdiffusion 2033 -1354 2033 -1354 0 feedthrough
rlabel pdiffusion 2040 -1354 2040 -1354 0 feedthrough
rlabel pdiffusion 2047 -1354 2047 -1354 0 feedthrough
rlabel pdiffusion 2054 -1354 2054 -1354 0 feedthrough
rlabel pdiffusion 2061 -1354 2061 -1354 0 feedthrough
rlabel pdiffusion 2068 -1354 2068 -1354 0 feedthrough
rlabel pdiffusion 2075 -1354 2075 -1354 0 feedthrough
rlabel pdiffusion 2082 -1354 2082 -1354 0 feedthrough
rlabel pdiffusion 2089 -1354 2089 -1354 0 feedthrough
rlabel pdiffusion 2096 -1354 2096 -1354 0 feedthrough
rlabel pdiffusion 2103 -1354 2103 -1354 0 feedthrough
rlabel pdiffusion 2110 -1354 2110 -1354 0 feedthrough
rlabel pdiffusion 2117 -1354 2117 -1354 0 feedthrough
rlabel pdiffusion 2124 -1354 2124 -1354 0 feedthrough
rlabel pdiffusion 2131 -1354 2131 -1354 0 feedthrough
rlabel pdiffusion 2138 -1354 2138 -1354 0 feedthrough
rlabel pdiffusion 2145 -1354 2145 -1354 0 feedthrough
rlabel pdiffusion 2152 -1354 2152 -1354 0 feedthrough
rlabel pdiffusion 2159 -1354 2159 -1354 0 feedthrough
rlabel pdiffusion 2166 -1354 2166 -1354 0 feedthrough
rlabel pdiffusion 2173 -1354 2173 -1354 0 feedthrough
rlabel pdiffusion 2180 -1354 2180 -1354 0 feedthrough
rlabel pdiffusion 2187 -1354 2187 -1354 0 feedthrough
rlabel pdiffusion 2194 -1354 2194 -1354 0 feedthrough
rlabel pdiffusion 2201 -1354 2201 -1354 0 feedthrough
rlabel pdiffusion 2208 -1354 2208 -1354 0 feedthrough
rlabel pdiffusion 2215 -1354 2215 -1354 0 feedthrough
rlabel pdiffusion 2222 -1354 2222 -1354 0 feedthrough
rlabel pdiffusion 2229 -1354 2229 -1354 0 feedthrough
rlabel pdiffusion 2236 -1354 2236 -1354 0 feedthrough
rlabel pdiffusion 2243 -1354 2243 -1354 0 feedthrough
rlabel pdiffusion 2250 -1354 2250 -1354 0 feedthrough
rlabel pdiffusion 2257 -1354 2257 -1354 0 feedthrough
rlabel pdiffusion 2264 -1354 2264 -1354 0 feedthrough
rlabel pdiffusion 2271 -1354 2271 -1354 0 feedthrough
rlabel pdiffusion 2278 -1354 2278 -1354 0 feedthrough
rlabel pdiffusion 2285 -1354 2285 -1354 0 feedthrough
rlabel pdiffusion 2292 -1354 2292 -1354 0 feedthrough
rlabel pdiffusion 2299 -1354 2299 -1354 0 feedthrough
rlabel pdiffusion 2306 -1354 2306 -1354 0 feedthrough
rlabel pdiffusion 2313 -1354 2313 -1354 0 feedthrough
rlabel pdiffusion 2320 -1354 2320 -1354 0 feedthrough
rlabel pdiffusion 2327 -1354 2327 -1354 0 feedthrough
rlabel pdiffusion 2334 -1354 2334 -1354 0 feedthrough
rlabel pdiffusion 2341 -1354 2341 -1354 0 cellNo=105
rlabel pdiffusion 2348 -1354 2348 -1354 0 feedthrough
rlabel pdiffusion 2355 -1354 2355 -1354 0 feedthrough
rlabel pdiffusion 2362 -1354 2362 -1354 0 feedthrough
rlabel pdiffusion 2369 -1354 2369 -1354 0 feedthrough
rlabel pdiffusion 2376 -1354 2376 -1354 0 feedthrough
rlabel pdiffusion 2383 -1354 2383 -1354 0 feedthrough
rlabel pdiffusion 2390 -1354 2390 -1354 0 feedthrough
rlabel pdiffusion 2397 -1354 2397 -1354 0 feedthrough
rlabel pdiffusion 2404 -1354 2404 -1354 0 feedthrough
rlabel pdiffusion 2411 -1354 2411 -1354 0 feedthrough
rlabel pdiffusion 2418 -1354 2418 -1354 0 feedthrough
rlabel pdiffusion 2425 -1354 2425 -1354 0 feedthrough
rlabel pdiffusion 2432 -1354 2432 -1354 0 feedthrough
rlabel pdiffusion 2439 -1354 2439 -1354 0 feedthrough
rlabel pdiffusion 2446 -1354 2446 -1354 0 feedthrough
rlabel pdiffusion 2453 -1354 2453 -1354 0 feedthrough
rlabel pdiffusion 2460 -1354 2460 -1354 0 feedthrough
rlabel pdiffusion 2467 -1354 2467 -1354 0 feedthrough
rlabel pdiffusion 2474 -1354 2474 -1354 0 feedthrough
rlabel pdiffusion 2481 -1354 2481 -1354 0 feedthrough
rlabel pdiffusion 2488 -1354 2488 -1354 0 feedthrough
rlabel pdiffusion 2495 -1354 2495 -1354 0 feedthrough
rlabel pdiffusion 2502 -1354 2502 -1354 0 feedthrough
rlabel pdiffusion 2509 -1354 2509 -1354 0 feedthrough
rlabel pdiffusion 2516 -1354 2516 -1354 0 feedthrough
rlabel pdiffusion 2523 -1354 2523 -1354 0 feedthrough
rlabel pdiffusion 2530 -1354 2530 -1354 0 feedthrough
rlabel pdiffusion 2537 -1354 2537 -1354 0 feedthrough
rlabel pdiffusion 2544 -1354 2544 -1354 0 feedthrough
rlabel pdiffusion 2551 -1354 2551 -1354 0 feedthrough
rlabel pdiffusion 2558 -1354 2558 -1354 0 feedthrough
rlabel pdiffusion 2565 -1354 2565 -1354 0 feedthrough
rlabel pdiffusion 2572 -1354 2572 -1354 0 feedthrough
rlabel pdiffusion 2579 -1354 2579 -1354 0 feedthrough
rlabel pdiffusion 3 -1531 3 -1531 0 feedthrough
rlabel pdiffusion 10 -1531 10 -1531 0 feedthrough
rlabel pdiffusion 17 -1531 17 -1531 0 cellNo=772
rlabel pdiffusion 24 -1531 24 -1531 0 cellNo=95
rlabel pdiffusion 31 -1531 31 -1531 0 feedthrough
rlabel pdiffusion 38 -1531 38 -1531 0 cellNo=731
rlabel pdiffusion 45 -1531 45 -1531 0 cellNo=917
rlabel pdiffusion 52 -1531 52 -1531 0 cellNo=437
rlabel pdiffusion 59 -1531 59 -1531 0 feedthrough
rlabel pdiffusion 66 -1531 66 -1531 0 feedthrough
rlabel pdiffusion 73 -1531 73 -1531 0 feedthrough
rlabel pdiffusion 80 -1531 80 -1531 0 feedthrough
rlabel pdiffusion 87 -1531 87 -1531 0 cellNo=532
rlabel pdiffusion 94 -1531 94 -1531 0 feedthrough
rlabel pdiffusion 101 -1531 101 -1531 0 feedthrough
rlabel pdiffusion 108 -1531 108 -1531 0 cellNo=126
rlabel pdiffusion 115 -1531 115 -1531 0 cellNo=378
rlabel pdiffusion 122 -1531 122 -1531 0 feedthrough
rlabel pdiffusion 129 -1531 129 -1531 0 feedthrough
rlabel pdiffusion 136 -1531 136 -1531 0 feedthrough
rlabel pdiffusion 143 -1531 143 -1531 0 feedthrough
rlabel pdiffusion 150 -1531 150 -1531 0 feedthrough
rlabel pdiffusion 157 -1531 157 -1531 0 feedthrough
rlabel pdiffusion 164 -1531 164 -1531 0 feedthrough
rlabel pdiffusion 171 -1531 171 -1531 0 feedthrough
rlabel pdiffusion 178 -1531 178 -1531 0 feedthrough
rlabel pdiffusion 185 -1531 185 -1531 0 feedthrough
rlabel pdiffusion 192 -1531 192 -1531 0 feedthrough
rlabel pdiffusion 199 -1531 199 -1531 0 cellNo=722
rlabel pdiffusion 206 -1531 206 -1531 0 cellNo=483
rlabel pdiffusion 213 -1531 213 -1531 0 feedthrough
rlabel pdiffusion 220 -1531 220 -1531 0 feedthrough
rlabel pdiffusion 227 -1531 227 -1531 0 feedthrough
rlabel pdiffusion 234 -1531 234 -1531 0 cellNo=686
rlabel pdiffusion 241 -1531 241 -1531 0 feedthrough
rlabel pdiffusion 248 -1531 248 -1531 0 feedthrough
rlabel pdiffusion 255 -1531 255 -1531 0 feedthrough
rlabel pdiffusion 262 -1531 262 -1531 0 feedthrough
rlabel pdiffusion 269 -1531 269 -1531 0 feedthrough
rlabel pdiffusion 276 -1531 276 -1531 0 feedthrough
rlabel pdiffusion 283 -1531 283 -1531 0 feedthrough
rlabel pdiffusion 290 -1531 290 -1531 0 feedthrough
rlabel pdiffusion 297 -1531 297 -1531 0 feedthrough
rlabel pdiffusion 304 -1531 304 -1531 0 feedthrough
rlabel pdiffusion 311 -1531 311 -1531 0 feedthrough
rlabel pdiffusion 318 -1531 318 -1531 0 feedthrough
rlabel pdiffusion 325 -1531 325 -1531 0 feedthrough
rlabel pdiffusion 332 -1531 332 -1531 0 feedthrough
rlabel pdiffusion 339 -1531 339 -1531 0 feedthrough
rlabel pdiffusion 346 -1531 346 -1531 0 feedthrough
rlabel pdiffusion 353 -1531 353 -1531 0 feedthrough
rlabel pdiffusion 360 -1531 360 -1531 0 feedthrough
rlabel pdiffusion 367 -1531 367 -1531 0 feedthrough
rlabel pdiffusion 374 -1531 374 -1531 0 feedthrough
rlabel pdiffusion 381 -1531 381 -1531 0 feedthrough
rlabel pdiffusion 388 -1531 388 -1531 0 feedthrough
rlabel pdiffusion 395 -1531 395 -1531 0 feedthrough
rlabel pdiffusion 402 -1531 402 -1531 0 feedthrough
rlabel pdiffusion 409 -1531 409 -1531 0 feedthrough
rlabel pdiffusion 416 -1531 416 -1531 0 feedthrough
rlabel pdiffusion 423 -1531 423 -1531 0 feedthrough
rlabel pdiffusion 430 -1531 430 -1531 0 feedthrough
rlabel pdiffusion 437 -1531 437 -1531 0 feedthrough
rlabel pdiffusion 444 -1531 444 -1531 0 feedthrough
rlabel pdiffusion 451 -1531 451 -1531 0 feedthrough
rlabel pdiffusion 458 -1531 458 -1531 0 feedthrough
rlabel pdiffusion 465 -1531 465 -1531 0 feedthrough
rlabel pdiffusion 472 -1531 472 -1531 0 feedthrough
rlabel pdiffusion 479 -1531 479 -1531 0 feedthrough
rlabel pdiffusion 486 -1531 486 -1531 0 feedthrough
rlabel pdiffusion 493 -1531 493 -1531 0 feedthrough
rlabel pdiffusion 500 -1531 500 -1531 0 feedthrough
rlabel pdiffusion 507 -1531 507 -1531 0 feedthrough
rlabel pdiffusion 514 -1531 514 -1531 0 cellNo=395
rlabel pdiffusion 521 -1531 521 -1531 0 feedthrough
rlabel pdiffusion 528 -1531 528 -1531 0 feedthrough
rlabel pdiffusion 535 -1531 535 -1531 0 feedthrough
rlabel pdiffusion 542 -1531 542 -1531 0 feedthrough
rlabel pdiffusion 549 -1531 549 -1531 0 feedthrough
rlabel pdiffusion 556 -1531 556 -1531 0 feedthrough
rlabel pdiffusion 563 -1531 563 -1531 0 feedthrough
rlabel pdiffusion 570 -1531 570 -1531 0 feedthrough
rlabel pdiffusion 577 -1531 577 -1531 0 feedthrough
rlabel pdiffusion 584 -1531 584 -1531 0 feedthrough
rlabel pdiffusion 591 -1531 591 -1531 0 cellNo=161
rlabel pdiffusion 598 -1531 598 -1531 0 feedthrough
rlabel pdiffusion 605 -1531 605 -1531 0 feedthrough
rlabel pdiffusion 612 -1531 612 -1531 0 feedthrough
rlabel pdiffusion 619 -1531 619 -1531 0 feedthrough
rlabel pdiffusion 626 -1531 626 -1531 0 cellNo=634
rlabel pdiffusion 633 -1531 633 -1531 0 feedthrough
rlabel pdiffusion 640 -1531 640 -1531 0 cellNo=55
rlabel pdiffusion 647 -1531 647 -1531 0 feedthrough
rlabel pdiffusion 654 -1531 654 -1531 0 feedthrough
rlabel pdiffusion 661 -1531 661 -1531 0 feedthrough
rlabel pdiffusion 668 -1531 668 -1531 0 feedthrough
rlabel pdiffusion 675 -1531 675 -1531 0 feedthrough
rlabel pdiffusion 682 -1531 682 -1531 0 feedthrough
rlabel pdiffusion 689 -1531 689 -1531 0 cellNo=623
rlabel pdiffusion 696 -1531 696 -1531 0 feedthrough
rlabel pdiffusion 703 -1531 703 -1531 0 feedthrough
rlabel pdiffusion 710 -1531 710 -1531 0 feedthrough
rlabel pdiffusion 717 -1531 717 -1531 0 feedthrough
rlabel pdiffusion 724 -1531 724 -1531 0 feedthrough
rlabel pdiffusion 731 -1531 731 -1531 0 feedthrough
rlabel pdiffusion 738 -1531 738 -1531 0 cellNo=424
rlabel pdiffusion 745 -1531 745 -1531 0 feedthrough
rlabel pdiffusion 752 -1531 752 -1531 0 feedthrough
rlabel pdiffusion 759 -1531 759 -1531 0 feedthrough
rlabel pdiffusion 766 -1531 766 -1531 0 feedthrough
rlabel pdiffusion 773 -1531 773 -1531 0 feedthrough
rlabel pdiffusion 780 -1531 780 -1531 0 feedthrough
rlabel pdiffusion 787 -1531 787 -1531 0 feedthrough
rlabel pdiffusion 794 -1531 794 -1531 0 cellNo=123
rlabel pdiffusion 801 -1531 801 -1531 0 feedthrough
rlabel pdiffusion 808 -1531 808 -1531 0 cellNo=799
rlabel pdiffusion 815 -1531 815 -1531 0 feedthrough
rlabel pdiffusion 822 -1531 822 -1531 0 cellNo=372
rlabel pdiffusion 829 -1531 829 -1531 0 feedthrough
rlabel pdiffusion 836 -1531 836 -1531 0 feedthrough
rlabel pdiffusion 843 -1531 843 -1531 0 feedthrough
rlabel pdiffusion 850 -1531 850 -1531 0 feedthrough
rlabel pdiffusion 857 -1531 857 -1531 0 feedthrough
rlabel pdiffusion 864 -1531 864 -1531 0 cellNo=29
rlabel pdiffusion 871 -1531 871 -1531 0 feedthrough
rlabel pdiffusion 878 -1531 878 -1531 0 cellNo=627
rlabel pdiffusion 885 -1531 885 -1531 0 cellNo=641
rlabel pdiffusion 892 -1531 892 -1531 0 feedthrough
rlabel pdiffusion 899 -1531 899 -1531 0 feedthrough
rlabel pdiffusion 906 -1531 906 -1531 0 cellNo=569
rlabel pdiffusion 913 -1531 913 -1531 0 feedthrough
rlabel pdiffusion 920 -1531 920 -1531 0 feedthrough
rlabel pdiffusion 927 -1531 927 -1531 0 feedthrough
rlabel pdiffusion 934 -1531 934 -1531 0 feedthrough
rlabel pdiffusion 941 -1531 941 -1531 0 cellNo=680
rlabel pdiffusion 948 -1531 948 -1531 0 feedthrough
rlabel pdiffusion 955 -1531 955 -1531 0 feedthrough
rlabel pdiffusion 962 -1531 962 -1531 0 cellNo=155
rlabel pdiffusion 969 -1531 969 -1531 0 feedthrough
rlabel pdiffusion 976 -1531 976 -1531 0 feedthrough
rlabel pdiffusion 983 -1531 983 -1531 0 feedthrough
rlabel pdiffusion 990 -1531 990 -1531 0 feedthrough
rlabel pdiffusion 997 -1531 997 -1531 0 feedthrough
rlabel pdiffusion 1004 -1531 1004 -1531 0 feedthrough
rlabel pdiffusion 1011 -1531 1011 -1531 0 feedthrough
rlabel pdiffusion 1018 -1531 1018 -1531 0 cellNo=422
rlabel pdiffusion 1025 -1531 1025 -1531 0 feedthrough
rlabel pdiffusion 1032 -1531 1032 -1531 0 feedthrough
rlabel pdiffusion 1039 -1531 1039 -1531 0 feedthrough
rlabel pdiffusion 1046 -1531 1046 -1531 0 feedthrough
rlabel pdiffusion 1053 -1531 1053 -1531 0 feedthrough
rlabel pdiffusion 1060 -1531 1060 -1531 0 feedthrough
rlabel pdiffusion 1067 -1531 1067 -1531 0 feedthrough
rlabel pdiffusion 1074 -1531 1074 -1531 0 feedthrough
rlabel pdiffusion 1081 -1531 1081 -1531 0 feedthrough
rlabel pdiffusion 1088 -1531 1088 -1531 0 cellNo=220
rlabel pdiffusion 1095 -1531 1095 -1531 0 feedthrough
rlabel pdiffusion 1102 -1531 1102 -1531 0 feedthrough
rlabel pdiffusion 1109 -1531 1109 -1531 0 feedthrough
rlabel pdiffusion 1116 -1531 1116 -1531 0 feedthrough
rlabel pdiffusion 1123 -1531 1123 -1531 0 feedthrough
rlabel pdiffusion 1130 -1531 1130 -1531 0 feedthrough
rlabel pdiffusion 1137 -1531 1137 -1531 0 feedthrough
rlabel pdiffusion 1144 -1531 1144 -1531 0 feedthrough
rlabel pdiffusion 1151 -1531 1151 -1531 0 cellNo=609
rlabel pdiffusion 1158 -1531 1158 -1531 0 cellNo=896
rlabel pdiffusion 1165 -1531 1165 -1531 0 feedthrough
rlabel pdiffusion 1172 -1531 1172 -1531 0 feedthrough
rlabel pdiffusion 1179 -1531 1179 -1531 0 feedthrough
rlabel pdiffusion 1186 -1531 1186 -1531 0 feedthrough
rlabel pdiffusion 1193 -1531 1193 -1531 0 feedthrough
rlabel pdiffusion 1200 -1531 1200 -1531 0 feedthrough
rlabel pdiffusion 1207 -1531 1207 -1531 0 feedthrough
rlabel pdiffusion 1214 -1531 1214 -1531 0 feedthrough
rlabel pdiffusion 1221 -1531 1221 -1531 0 feedthrough
rlabel pdiffusion 1228 -1531 1228 -1531 0 feedthrough
rlabel pdiffusion 1235 -1531 1235 -1531 0 feedthrough
rlabel pdiffusion 1242 -1531 1242 -1531 0 feedthrough
rlabel pdiffusion 1249 -1531 1249 -1531 0 cellNo=771
rlabel pdiffusion 1256 -1531 1256 -1531 0 cellNo=360
rlabel pdiffusion 1263 -1531 1263 -1531 0 cellNo=53
rlabel pdiffusion 1270 -1531 1270 -1531 0 feedthrough
rlabel pdiffusion 1277 -1531 1277 -1531 0 feedthrough
rlabel pdiffusion 1284 -1531 1284 -1531 0 cellNo=189
rlabel pdiffusion 1291 -1531 1291 -1531 0 feedthrough
rlabel pdiffusion 1298 -1531 1298 -1531 0 feedthrough
rlabel pdiffusion 1305 -1531 1305 -1531 0 feedthrough
rlabel pdiffusion 1312 -1531 1312 -1531 0 feedthrough
rlabel pdiffusion 1319 -1531 1319 -1531 0 feedthrough
rlabel pdiffusion 1326 -1531 1326 -1531 0 feedthrough
rlabel pdiffusion 1333 -1531 1333 -1531 0 feedthrough
rlabel pdiffusion 1340 -1531 1340 -1531 0 feedthrough
rlabel pdiffusion 1347 -1531 1347 -1531 0 cellNo=254
rlabel pdiffusion 1354 -1531 1354 -1531 0 feedthrough
rlabel pdiffusion 1361 -1531 1361 -1531 0 feedthrough
rlabel pdiffusion 1368 -1531 1368 -1531 0 feedthrough
rlabel pdiffusion 1375 -1531 1375 -1531 0 feedthrough
rlabel pdiffusion 1382 -1531 1382 -1531 0 feedthrough
rlabel pdiffusion 1389 -1531 1389 -1531 0 feedthrough
rlabel pdiffusion 1396 -1531 1396 -1531 0 feedthrough
rlabel pdiffusion 1403 -1531 1403 -1531 0 feedthrough
rlabel pdiffusion 1410 -1531 1410 -1531 0 feedthrough
rlabel pdiffusion 1417 -1531 1417 -1531 0 feedthrough
rlabel pdiffusion 1424 -1531 1424 -1531 0 cellNo=807
rlabel pdiffusion 1431 -1531 1431 -1531 0 feedthrough
rlabel pdiffusion 1438 -1531 1438 -1531 0 feedthrough
rlabel pdiffusion 1445 -1531 1445 -1531 0 feedthrough
rlabel pdiffusion 1452 -1531 1452 -1531 0 feedthrough
rlabel pdiffusion 1459 -1531 1459 -1531 0 feedthrough
rlabel pdiffusion 1466 -1531 1466 -1531 0 feedthrough
rlabel pdiffusion 1473 -1531 1473 -1531 0 feedthrough
rlabel pdiffusion 1480 -1531 1480 -1531 0 cellNo=614
rlabel pdiffusion 1487 -1531 1487 -1531 0 cellNo=329
rlabel pdiffusion 1494 -1531 1494 -1531 0 feedthrough
rlabel pdiffusion 1501 -1531 1501 -1531 0 cellNo=595
rlabel pdiffusion 1508 -1531 1508 -1531 0 feedthrough
rlabel pdiffusion 1515 -1531 1515 -1531 0 feedthrough
rlabel pdiffusion 1522 -1531 1522 -1531 0 feedthrough
rlabel pdiffusion 1529 -1531 1529 -1531 0 feedthrough
rlabel pdiffusion 1536 -1531 1536 -1531 0 feedthrough
rlabel pdiffusion 1543 -1531 1543 -1531 0 feedthrough
rlabel pdiffusion 1550 -1531 1550 -1531 0 feedthrough
rlabel pdiffusion 1557 -1531 1557 -1531 0 feedthrough
rlabel pdiffusion 1564 -1531 1564 -1531 0 feedthrough
rlabel pdiffusion 1571 -1531 1571 -1531 0 feedthrough
rlabel pdiffusion 1578 -1531 1578 -1531 0 feedthrough
rlabel pdiffusion 1585 -1531 1585 -1531 0 feedthrough
rlabel pdiffusion 1592 -1531 1592 -1531 0 feedthrough
rlabel pdiffusion 1599 -1531 1599 -1531 0 feedthrough
rlabel pdiffusion 1606 -1531 1606 -1531 0 feedthrough
rlabel pdiffusion 1613 -1531 1613 -1531 0 feedthrough
rlabel pdiffusion 1620 -1531 1620 -1531 0 feedthrough
rlabel pdiffusion 1627 -1531 1627 -1531 0 feedthrough
rlabel pdiffusion 1634 -1531 1634 -1531 0 feedthrough
rlabel pdiffusion 1641 -1531 1641 -1531 0 feedthrough
rlabel pdiffusion 1648 -1531 1648 -1531 0 feedthrough
rlabel pdiffusion 1655 -1531 1655 -1531 0 feedthrough
rlabel pdiffusion 1662 -1531 1662 -1531 0 feedthrough
rlabel pdiffusion 1669 -1531 1669 -1531 0 feedthrough
rlabel pdiffusion 1676 -1531 1676 -1531 0 feedthrough
rlabel pdiffusion 1683 -1531 1683 -1531 0 feedthrough
rlabel pdiffusion 1690 -1531 1690 -1531 0 feedthrough
rlabel pdiffusion 1697 -1531 1697 -1531 0 feedthrough
rlabel pdiffusion 1704 -1531 1704 -1531 0 feedthrough
rlabel pdiffusion 1711 -1531 1711 -1531 0 feedthrough
rlabel pdiffusion 1718 -1531 1718 -1531 0 feedthrough
rlabel pdiffusion 1725 -1531 1725 -1531 0 feedthrough
rlabel pdiffusion 1732 -1531 1732 -1531 0 feedthrough
rlabel pdiffusion 1739 -1531 1739 -1531 0 feedthrough
rlabel pdiffusion 1746 -1531 1746 -1531 0 feedthrough
rlabel pdiffusion 1753 -1531 1753 -1531 0 feedthrough
rlabel pdiffusion 1760 -1531 1760 -1531 0 feedthrough
rlabel pdiffusion 1767 -1531 1767 -1531 0 feedthrough
rlabel pdiffusion 1774 -1531 1774 -1531 0 feedthrough
rlabel pdiffusion 1781 -1531 1781 -1531 0 feedthrough
rlabel pdiffusion 1788 -1531 1788 -1531 0 feedthrough
rlabel pdiffusion 1795 -1531 1795 -1531 0 feedthrough
rlabel pdiffusion 1802 -1531 1802 -1531 0 feedthrough
rlabel pdiffusion 1809 -1531 1809 -1531 0 feedthrough
rlabel pdiffusion 1816 -1531 1816 -1531 0 feedthrough
rlabel pdiffusion 1823 -1531 1823 -1531 0 feedthrough
rlabel pdiffusion 1830 -1531 1830 -1531 0 feedthrough
rlabel pdiffusion 1837 -1531 1837 -1531 0 feedthrough
rlabel pdiffusion 1844 -1531 1844 -1531 0 feedthrough
rlabel pdiffusion 1851 -1531 1851 -1531 0 feedthrough
rlabel pdiffusion 1858 -1531 1858 -1531 0 feedthrough
rlabel pdiffusion 1865 -1531 1865 -1531 0 feedthrough
rlabel pdiffusion 1872 -1531 1872 -1531 0 feedthrough
rlabel pdiffusion 1879 -1531 1879 -1531 0 feedthrough
rlabel pdiffusion 1886 -1531 1886 -1531 0 feedthrough
rlabel pdiffusion 1893 -1531 1893 -1531 0 feedthrough
rlabel pdiffusion 1900 -1531 1900 -1531 0 feedthrough
rlabel pdiffusion 1907 -1531 1907 -1531 0 feedthrough
rlabel pdiffusion 1914 -1531 1914 -1531 0 feedthrough
rlabel pdiffusion 1921 -1531 1921 -1531 0 feedthrough
rlabel pdiffusion 1928 -1531 1928 -1531 0 feedthrough
rlabel pdiffusion 1935 -1531 1935 -1531 0 feedthrough
rlabel pdiffusion 1942 -1531 1942 -1531 0 feedthrough
rlabel pdiffusion 1949 -1531 1949 -1531 0 feedthrough
rlabel pdiffusion 1956 -1531 1956 -1531 0 feedthrough
rlabel pdiffusion 1963 -1531 1963 -1531 0 feedthrough
rlabel pdiffusion 1970 -1531 1970 -1531 0 feedthrough
rlabel pdiffusion 1977 -1531 1977 -1531 0 feedthrough
rlabel pdiffusion 1984 -1531 1984 -1531 0 feedthrough
rlabel pdiffusion 1991 -1531 1991 -1531 0 feedthrough
rlabel pdiffusion 1998 -1531 1998 -1531 0 feedthrough
rlabel pdiffusion 2005 -1531 2005 -1531 0 feedthrough
rlabel pdiffusion 2012 -1531 2012 -1531 0 feedthrough
rlabel pdiffusion 2019 -1531 2019 -1531 0 feedthrough
rlabel pdiffusion 2026 -1531 2026 -1531 0 feedthrough
rlabel pdiffusion 2033 -1531 2033 -1531 0 feedthrough
rlabel pdiffusion 2040 -1531 2040 -1531 0 feedthrough
rlabel pdiffusion 2047 -1531 2047 -1531 0 feedthrough
rlabel pdiffusion 2054 -1531 2054 -1531 0 feedthrough
rlabel pdiffusion 2061 -1531 2061 -1531 0 feedthrough
rlabel pdiffusion 2068 -1531 2068 -1531 0 feedthrough
rlabel pdiffusion 2075 -1531 2075 -1531 0 feedthrough
rlabel pdiffusion 2082 -1531 2082 -1531 0 feedthrough
rlabel pdiffusion 2089 -1531 2089 -1531 0 feedthrough
rlabel pdiffusion 2096 -1531 2096 -1531 0 feedthrough
rlabel pdiffusion 2103 -1531 2103 -1531 0 feedthrough
rlabel pdiffusion 2110 -1531 2110 -1531 0 feedthrough
rlabel pdiffusion 2117 -1531 2117 -1531 0 feedthrough
rlabel pdiffusion 2124 -1531 2124 -1531 0 feedthrough
rlabel pdiffusion 2131 -1531 2131 -1531 0 feedthrough
rlabel pdiffusion 2138 -1531 2138 -1531 0 feedthrough
rlabel pdiffusion 2145 -1531 2145 -1531 0 feedthrough
rlabel pdiffusion 2152 -1531 2152 -1531 0 feedthrough
rlabel pdiffusion 2159 -1531 2159 -1531 0 feedthrough
rlabel pdiffusion 2166 -1531 2166 -1531 0 feedthrough
rlabel pdiffusion 2173 -1531 2173 -1531 0 feedthrough
rlabel pdiffusion 2180 -1531 2180 -1531 0 feedthrough
rlabel pdiffusion 2187 -1531 2187 -1531 0 feedthrough
rlabel pdiffusion 2194 -1531 2194 -1531 0 feedthrough
rlabel pdiffusion 2201 -1531 2201 -1531 0 feedthrough
rlabel pdiffusion 2208 -1531 2208 -1531 0 feedthrough
rlabel pdiffusion 2215 -1531 2215 -1531 0 feedthrough
rlabel pdiffusion 2222 -1531 2222 -1531 0 feedthrough
rlabel pdiffusion 2229 -1531 2229 -1531 0 feedthrough
rlabel pdiffusion 2236 -1531 2236 -1531 0 feedthrough
rlabel pdiffusion 2243 -1531 2243 -1531 0 feedthrough
rlabel pdiffusion 2250 -1531 2250 -1531 0 feedthrough
rlabel pdiffusion 2257 -1531 2257 -1531 0 feedthrough
rlabel pdiffusion 2264 -1531 2264 -1531 0 feedthrough
rlabel pdiffusion 2271 -1531 2271 -1531 0 feedthrough
rlabel pdiffusion 2278 -1531 2278 -1531 0 feedthrough
rlabel pdiffusion 2285 -1531 2285 -1531 0 feedthrough
rlabel pdiffusion 2292 -1531 2292 -1531 0 feedthrough
rlabel pdiffusion 2299 -1531 2299 -1531 0 feedthrough
rlabel pdiffusion 2306 -1531 2306 -1531 0 feedthrough
rlabel pdiffusion 2313 -1531 2313 -1531 0 feedthrough
rlabel pdiffusion 2320 -1531 2320 -1531 0 feedthrough
rlabel pdiffusion 2327 -1531 2327 -1531 0 feedthrough
rlabel pdiffusion 2334 -1531 2334 -1531 0 feedthrough
rlabel pdiffusion 2341 -1531 2341 -1531 0 feedthrough
rlabel pdiffusion 2348 -1531 2348 -1531 0 feedthrough
rlabel pdiffusion 2355 -1531 2355 -1531 0 feedthrough
rlabel pdiffusion 2362 -1531 2362 -1531 0 feedthrough
rlabel pdiffusion 2369 -1531 2369 -1531 0 feedthrough
rlabel pdiffusion 2376 -1531 2376 -1531 0 feedthrough
rlabel pdiffusion 2383 -1531 2383 -1531 0 feedthrough
rlabel pdiffusion 2390 -1531 2390 -1531 0 feedthrough
rlabel pdiffusion 2397 -1531 2397 -1531 0 feedthrough
rlabel pdiffusion 2404 -1531 2404 -1531 0 feedthrough
rlabel pdiffusion 2411 -1531 2411 -1531 0 feedthrough
rlabel pdiffusion 2418 -1531 2418 -1531 0 feedthrough
rlabel pdiffusion 2425 -1531 2425 -1531 0 feedthrough
rlabel pdiffusion 2432 -1531 2432 -1531 0 feedthrough
rlabel pdiffusion 2439 -1531 2439 -1531 0 feedthrough
rlabel pdiffusion 2446 -1531 2446 -1531 0 feedthrough
rlabel pdiffusion 2453 -1531 2453 -1531 0 feedthrough
rlabel pdiffusion 2460 -1531 2460 -1531 0 feedthrough
rlabel pdiffusion 2467 -1531 2467 -1531 0 feedthrough
rlabel pdiffusion 2474 -1531 2474 -1531 0 feedthrough
rlabel pdiffusion 2481 -1531 2481 -1531 0 feedthrough
rlabel pdiffusion 2488 -1531 2488 -1531 0 feedthrough
rlabel pdiffusion 2495 -1531 2495 -1531 0 feedthrough
rlabel pdiffusion 2502 -1531 2502 -1531 0 feedthrough
rlabel pdiffusion 2509 -1531 2509 -1531 0 feedthrough
rlabel pdiffusion 2516 -1531 2516 -1531 0 feedthrough
rlabel pdiffusion 2523 -1531 2523 -1531 0 feedthrough
rlabel pdiffusion 2530 -1531 2530 -1531 0 feedthrough
rlabel pdiffusion 2537 -1531 2537 -1531 0 feedthrough
rlabel pdiffusion 2544 -1531 2544 -1531 0 feedthrough
rlabel pdiffusion 2551 -1531 2551 -1531 0 feedthrough
rlabel pdiffusion 2558 -1531 2558 -1531 0 feedthrough
rlabel pdiffusion 3 -1704 3 -1704 0 cellNo=1046
rlabel pdiffusion 10 -1704 10 -1704 0 cellNo=1156
rlabel pdiffusion 17 -1704 17 -1704 0 feedthrough
rlabel pdiffusion 24 -1704 24 -1704 0 feedthrough
rlabel pdiffusion 31 -1704 31 -1704 0 feedthrough
rlabel pdiffusion 38 -1704 38 -1704 0 feedthrough
rlabel pdiffusion 45 -1704 45 -1704 0 feedthrough
rlabel pdiffusion 52 -1704 52 -1704 0 feedthrough
rlabel pdiffusion 59 -1704 59 -1704 0 feedthrough
rlabel pdiffusion 66 -1704 66 -1704 0 feedthrough
rlabel pdiffusion 73 -1704 73 -1704 0 feedthrough
rlabel pdiffusion 80 -1704 80 -1704 0 feedthrough
rlabel pdiffusion 87 -1704 87 -1704 0 feedthrough
rlabel pdiffusion 94 -1704 94 -1704 0 cellNo=869
rlabel pdiffusion 101 -1704 101 -1704 0 feedthrough
rlabel pdiffusion 108 -1704 108 -1704 0 feedthrough
rlabel pdiffusion 115 -1704 115 -1704 0 feedthrough
rlabel pdiffusion 122 -1704 122 -1704 0 feedthrough
rlabel pdiffusion 129 -1704 129 -1704 0 feedthrough
rlabel pdiffusion 136 -1704 136 -1704 0 feedthrough
rlabel pdiffusion 143 -1704 143 -1704 0 feedthrough
rlabel pdiffusion 150 -1704 150 -1704 0 feedthrough
rlabel pdiffusion 157 -1704 157 -1704 0 feedthrough
rlabel pdiffusion 164 -1704 164 -1704 0 feedthrough
rlabel pdiffusion 171 -1704 171 -1704 0 feedthrough
rlabel pdiffusion 178 -1704 178 -1704 0 cellNo=119
rlabel pdiffusion 185 -1704 185 -1704 0 feedthrough
rlabel pdiffusion 192 -1704 192 -1704 0 cellNo=299
rlabel pdiffusion 199 -1704 199 -1704 0 feedthrough
rlabel pdiffusion 206 -1704 206 -1704 0 feedthrough
rlabel pdiffusion 213 -1704 213 -1704 0 cellNo=700
rlabel pdiffusion 220 -1704 220 -1704 0 feedthrough
rlabel pdiffusion 227 -1704 227 -1704 0 cellNo=959
rlabel pdiffusion 234 -1704 234 -1704 0 cellNo=31
rlabel pdiffusion 241 -1704 241 -1704 0 feedthrough
rlabel pdiffusion 248 -1704 248 -1704 0 cellNo=10
rlabel pdiffusion 255 -1704 255 -1704 0 feedthrough
rlabel pdiffusion 262 -1704 262 -1704 0 feedthrough
rlabel pdiffusion 269 -1704 269 -1704 0 feedthrough
rlabel pdiffusion 276 -1704 276 -1704 0 feedthrough
rlabel pdiffusion 283 -1704 283 -1704 0 feedthrough
rlabel pdiffusion 290 -1704 290 -1704 0 feedthrough
rlabel pdiffusion 297 -1704 297 -1704 0 feedthrough
rlabel pdiffusion 304 -1704 304 -1704 0 feedthrough
rlabel pdiffusion 311 -1704 311 -1704 0 feedthrough
rlabel pdiffusion 318 -1704 318 -1704 0 feedthrough
rlabel pdiffusion 325 -1704 325 -1704 0 feedthrough
rlabel pdiffusion 332 -1704 332 -1704 0 feedthrough
rlabel pdiffusion 339 -1704 339 -1704 0 feedthrough
rlabel pdiffusion 346 -1704 346 -1704 0 feedthrough
rlabel pdiffusion 353 -1704 353 -1704 0 feedthrough
rlabel pdiffusion 360 -1704 360 -1704 0 feedthrough
rlabel pdiffusion 367 -1704 367 -1704 0 feedthrough
rlabel pdiffusion 374 -1704 374 -1704 0 feedthrough
rlabel pdiffusion 381 -1704 381 -1704 0 feedthrough
rlabel pdiffusion 388 -1704 388 -1704 0 feedthrough
rlabel pdiffusion 395 -1704 395 -1704 0 feedthrough
rlabel pdiffusion 402 -1704 402 -1704 0 feedthrough
rlabel pdiffusion 409 -1704 409 -1704 0 feedthrough
rlabel pdiffusion 416 -1704 416 -1704 0 feedthrough
rlabel pdiffusion 423 -1704 423 -1704 0 feedthrough
rlabel pdiffusion 430 -1704 430 -1704 0 feedthrough
rlabel pdiffusion 437 -1704 437 -1704 0 feedthrough
rlabel pdiffusion 444 -1704 444 -1704 0 feedthrough
rlabel pdiffusion 451 -1704 451 -1704 0 cellNo=236
rlabel pdiffusion 458 -1704 458 -1704 0 cellNo=693
rlabel pdiffusion 465 -1704 465 -1704 0 feedthrough
rlabel pdiffusion 472 -1704 472 -1704 0 feedthrough
rlabel pdiffusion 479 -1704 479 -1704 0 cellNo=910
rlabel pdiffusion 486 -1704 486 -1704 0 feedthrough
rlabel pdiffusion 493 -1704 493 -1704 0 feedthrough
rlabel pdiffusion 500 -1704 500 -1704 0 feedthrough
rlabel pdiffusion 507 -1704 507 -1704 0 feedthrough
rlabel pdiffusion 514 -1704 514 -1704 0 feedthrough
rlabel pdiffusion 521 -1704 521 -1704 0 feedthrough
rlabel pdiffusion 528 -1704 528 -1704 0 feedthrough
rlabel pdiffusion 535 -1704 535 -1704 0 feedthrough
rlabel pdiffusion 542 -1704 542 -1704 0 feedthrough
rlabel pdiffusion 549 -1704 549 -1704 0 feedthrough
rlabel pdiffusion 556 -1704 556 -1704 0 feedthrough
rlabel pdiffusion 563 -1704 563 -1704 0 feedthrough
rlabel pdiffusion 570 -1704 570 -1704 0 feedthrough
rlabel pdiffusion 577 -1704 577 -1704 0 cellNo=469
rlabel pdiffusion 584 -1704 584 -1704 0 feedthrough
rlabel pdiffusion 591 -1704 591 -1704 0 feedthrough
rlabel pdiffusion 598 -1704 598 -1704 0 feedthrough
rlabel pdiffusion 605 -1704 605 -1704 0 feedthrough
rlabel pdiffusion 612 -1704 612 -1704 0 feedthrough
rlabel pdiffusion 619 -1704 619 -1704 0 feedthrough
rlabel pdiffusion 626 -1704 626 -1704 0 feedthrough
rlabel pdiffusion 633 -1704 633 -1704 0 feedthrough
rlabel pdiffusion 640 -1704 640 -1704 0 cellNo=785
rlabel pdiffusion 647 -1704 647 -1704 0 feedthrough
rlabel pdiffusion 654 -1704 654 -1704 0 feedthrough
rlabel pdiffusion 661 -1704 661 -1704 0 feedthrough
rlabel pdiffusion 668 -1704 668 -1704 0 feedthrough
rlabel pdiffusion 675 -1704 675 -1704 0 feedthrough
rlabel pdiffusion 682 -1704 682 -1704 0 feedthrough
rlabel pdiffusion 689 -1704 689 -1704 0 feedthrough
rlabel pdiffusion 696 -1704 696 -1704 0 cellNo=447
rlabel pdiffusion 703 -1704 703 -1704 0 feedthrough
rlabel pdiffusion 710 -1704 710 -1704 0 feedthrough
rlabel pdiffusion 717 -1704 717 -1704 0 cellNo=828
rlabel pdiffusion 724 -1704 724 -1704 0 feedthrough
rlabel pdiffusion 731 -1704 731 -1704 0 feedthrough
rlabel pdiffusion 738 -1704 738 -1704 0 feedthrough
rlabel pdiffusion 745 -1704 745 -1704 0 feedthrough
rlabel pdiffusion 752 -1704 752 -1704 0 feedthrough
rlabel pdiffusion 759 -1704 759 -1704 0 feedthrough
rlabel pdiffusion 766 -1704 766 -1704 0 feedthrough
rlabel pdiffusion 773 -1704 773 -1704 0 feedthrough
rlabel pdiffusion 780 -1704 780 -1704 0 feedthrough
rlabel pdiffusion 787 -1704 787 -1704 0 feedthrough
rlabel pdiffusion 794 -1704 794 -1704 0 feedthrough
rlabel pdiffusion 801 -1704 801 -1704 0 feedthrough
rlabel pdiffusion 808 -1704 808 -1704 0 feedthrough
rlabel pdiffusion 815 -1704 815 -1704 0 feedthrough
rlabel pdiffusion 822 -1704 822 -1704 0 feedthrough
rlabel pdiffusion 829 -1704 829 -1704 0 feedthrough
rlabel pdiffusion 836 -1704 836 -1704 0 feedthrough
rlabel pdiffusion 843 -1704 843 -1704 0 feedthrough
rlabel pdiffusion 850 -1704 850 -1704 0 feedthrough
rlabel pdiffusion 857 -1704 857 -1704 0 cellNo=567
rlabel pdiffusion 864 -1704 864 -1704 0 feedthrough
rlabel pdiffusion 871 -1704 871 -1704 0 feedthrough
rlabel pdiffusion 878 -1704 878 -1704 0 feedthrough
rlabel pdiffusion 885 -1704 885 -1704 0 feedthrough
rlabel pdiffusion 892 -1704 892 -1704 0 feedthrough
rlabel pdiffusion 899 -1704 899 -1704 0 feedthrough
rlabel pdiffusion 906 -1704 906 -1704 0 feedthrough
rlabel pdiffusion 913 -1704 913 -1704 0 feedthrough
rlabel pdiffusion 920 -1704 920 -1704 0 feedthrough
rlabel pdiffusion 927 -1704 927 -1704 0 feedthrough
rlabel pdiffusion 934 -1704 934 -1704 0 cellNo=577
rlabel pdiffusion 941 -1704 941 -1704 0 feedthrough
rlabel pdiffusion 948 -1704 948 -1704 0 feedthrough
rlabel pdiffusion 955 -1704 955 -1704 0 feedthrough
rlabel pdiffusion 962 -1704 962 -1704 0 feedthrough
rlabel pdiffusion 969 -1704 969 -1704 0 cellNo=689
rlabel pdiffusion 976 -1704 976 -1704 0 feedthrough
rlabel pdiffusion 983 -1704 983 -1704 0 feedthrough
rlabel pdiffusion 990 -1704 990 -1704 0 feedthrough
rlabel pdiffusion 997 -1704 997 -1704 0 feedthrough
rlabel pdiffusion 1004 -1704 1004 -1704 0 feedthrough
rlabel pdiffusion 1011 -1704 1011 -1704 0 feedthrough
rlabel pdiffusion 1018 -1704 1018 -1704 0 cellNo=475
rlabel pdiffusion 1025 -1704 1025 -1704 0 feedthrough
rlabel pdiffusion 1032 -1704 1032 -1704 0 cellNo=46
rlabel pdiffusion 1039 -1704 1039 -1704 0 feedthrough
rlabel pdiffusion 1046 -1704 1046 -1704 0 feedthrough
rlabel pdiffusion 1053 -1704 1053 -1704 0 feedthrough
rlabel pdiffusion 1060 -1704 1060 -1704 0 feedthrough
rlabel pdiffusion 1067 -1704 1067 -1704 0 feedthrough
rlabel pdiffusion 1074 -1704 1074 -1704 0 cellNo=607
rlabel pdiffusion 1081 -1704 1081 -1704 0 feedthrough
rlabel pdiffusion 1088 -1704 1088 -1704 0 feedthrough
rlabel pdiffusion 1095 -1704 1095 -1704 0 feedthrough
rlabel pdiffusion 1102 -1704 1102 -1704 0 feedthrough
rlabel pdiffusion 1109 -1704 1109 -1704 0 cellNo=149
rlabel pdiffusion 1116 -1704 1116 -1704 0 feedthrough
rlabel pdiffusion 1123 -1704 1123 -1704 0 feedthrough
rlabel pdiffusion 1130 -1704 1130 -1704 0 feedthrough
rlabel pdiffusion 1137 -1704 1137 -1704 0 feedthrough
rlabel pdiffusion 1144 -1704 1144 -1704 0 feedthrough
rlabel pdiffusion 1151 -1704 1151 -1704 0 cellNo=230
rlabel pdiffusion 1158 -1704 1158 -1704 0 feedthrough
rlabel pdiffusion 1165 -1704 1165 -1704 0 feedthrough
rlabel pdiffusion 1172 -1704 1172 -1704 0 feedthrough
rlabel pdiffusion 1179 -1704 1179 -1704 0 feedthrough
rlabel pdiffusion 1186 -1704 1186 -1704 0 feedthrough
rlabel pdiffusion 1193 -1704 1193 -1704 0 feedthrough
rlabel pdiffusion 1200 -1704 1200 -1704 0 feedthrough
rlabel pdiffusion 1207 -1704 1207 -1704 0 feedthrough
rlabel pdiffusion 1214 -1704 1214 -1704 0 feedthrough
rlabel pdiffusion 1221 -1704 1221 -1704 0 feedthrough
rlabel pdiffusion 1228 -1704 1228 -1704 0 feedthrough
rlabel pdiffusion 1235 -1704 1235 -1704 0 feedthrough
rlabel pdiffusion 1242 -1704 1242 -1704 0 feedthrough
rlabel pdiffusion 1249 -1704 1249 -1704 0 feedthrough
rlabel pdiffusion 1256 -1704 1256 -1704 0 feedthrough
rlabel pdiffusion 1263 -1704 1263 -1704 0 cellNo=206
rlabel pdiffusion 1270 -1704 1270 -1704 0 feedthrough
rlabel pdiffusion 1277 -1704 1277 -1704 0 cellNo=882
rlabel pdiffusion 1284 -1704 1284 -1704 0 feedthrough
rlabel pdiffusion 1291 -1704 1291 -1704 0 cellNo=791
rlabel pdiffusion 1298 -1704 1298 -1704 0 feedthrough
rlabel pdiffusion 1305 -1704 1305 -1704 0 feedthrough
rlabel pdiffusion 1312 -1704 1312 -1704 0 feedthrough
rlabel pdiffusion 1319 -1704 1319 -1704 0 feedthrough
rlabel pdiffusion 1326 -1704 1326 -1704 0 feedthrough
rlabel pdiffusion 1333 -1704 1333 -1704 0 feedthrough
rlabel pdiffusion 1340 -1704 1340 -1704 0 feedthrough
rlabel pdiffusion 1347 -1704 1347 -1704 0 feedthrough
rlabel pdiffusion 1354 -1704 1354 -1704 0 feedthrough
rlabel pdiffusion 1361 -1704 1361 -1704 0 cellNo=756
rlabel pdiffusion 1368 -1704 1368 -1704 0 feedthrough
rlabel pdiffusion 1375 -1704 1375 -1704 0 feedthrough
rlabel pdiffusion 1382 -1704 1382 -1704 0 feedthrough
rlabel pdiffusion 1389 -1704 1389 -1704 0 feedthrough
rlabel pdiffusion 1396 -1704 1396 -1704 0 feedthrough
rlabel pdiffusion 1403 -1704 1403 -1704 0 feedthrough
rlabel pdiffusion 1410 -1704 1410 -1704 0 feedthrough
rlabel pdiffusion 1417 -1704 1417 -1704 0 feedthrough
rlabel pdiffusion 1424 -1704 1424 -1704 0 feedthrough
rlabel pdiffusion 1431 -1704 1431 -1704 0 feedthrough
rlabel pdiffusion 1438 -1704 1438 -1704 0 cellNo=674
rlabel pdiffusion 1445 -1704 1445 -1704 0 feedthrough
rlabel pdiffusion 1452 -1704 1452 -1704 0 feedthrough
rlabel pdiffusion 1459 -1704 1459 -1704 0 feedthrough
rlabel pdiffusion 1466 -1704 1466 -1704 0 cellNo=436
rlabel pdiffusion 1473 -1704 1473 -1704 0 feedthrough
rlabel pdiffusion 1480 -1704 1480 -1704 0 feedthrough
rlabel pdiffusion 1487 -1704 1487 -1704 0 feedthrough
rlabel pdiffusion 1494 -1704 1494 -1704 0 cellNo=68
rlabel pdiffusion 1501 -1704 1501 -1704 0 feedthrough
rlabel pdiffusion 1508 -1704 1508 -1704 0 cellNo=664
rlabel pdiffusion 1515 -1704 1515 -1704 0 feedthrough
rlabel pdiffusion 1522 -1704 1522 -1704 0 feedthrough
rlabel pdiffusion 1529 -1704 1529 -1704 0 cellNo=106
rlabel pdiffusion 1536 -1704 1536 -1704 0 cellNo=593
rlabel pdiffusion 1543 -1704 1543 -1704 0 feedthrough
rlabel pdiffusion 1550 -1704 1550 -1704 0 feedthrough
rlabel pdiffusion 1557 -1704 1557 -1704 0 feedthrough
rlabel pdiffusion 1564 -1704 1564 -1704 0 feedthrough
rlabel pdiffusion 1571 -1704 1571 -1704 0 feedthrough
rlabel pdiffusion 1578 -1704 1578 -1704 0 feedthrough
rlabel pdiffusion 1585 -1704 1585 -1704 0 feedthrough
rlabel pdiffusion 1592 -1704 1592 -1704 0 feedthrough
rlabel pdiffusion 1599 -1704 1599 -1704 0 feedthrough
rlabel pdiffusion 1606 -1704 1606 -1704 0 feedthrough
rlabel pdiffusion 1613 -1704 1613 -1704 0 feedthrough
rlabel pdiffusion 1620 -1704 1620 -1704 0 feedthrough
rlabel pdiffusion 1627 -1704 1627 -1704 0 feedthrough
rlabel pdiffusion 1634 -1704 1634 -1704 0 feedthrough
rlabel pdiffusion 1641 -1704 1641 -1704 0 feedthrough
rlabel pdiffusion 1648 -1704 1648 -1704 0 feedthrough
rlabel pdiffusion 1655 -1704 1655 -1704 0 feedthrough
rlabel pdiffusion 1662 -1704 1662 -1704 0 feedthrough
rlabel pdiffusion 1669 -1704 1669 -1704 0 feedthrough
rlabel pdiffusion 1676 -1704 1676 -1704 0 feedthrough
rlabel pdiffusion 1683 -1704 1683 -1704 0 feedthrough
rlabel pdiffusion 1690 -1704 1690 -1704 0 feedthrough
rlabel pdiffusion 1697 -1704 1697 -1704 0 feedthrough
rlabel pdiffusion 1704 -1704 1704 -1704 0 cellNo=440
rlabel pdiffusion 1711 -1704 1711 -1704 0 feedthrough
rlabel pdiffusion 1718 -1704 1718 -1704 0 feedthrough
rlabel pdiffusion 1725 -1704 1725 -1704 0 feedthrough
rlabel pdiffusion 1732 -1704 1732 -1704 0 feedthrough
rlabel pdiffusion 1739 -1704 1739 -1704 0 feedthrough
rlabel pdiffusion 1746 -1704 1746 -1704 0 feedthrough
rlabel pdiffusion 1753 -1704 1753 -1704 0 feedthrough
rlabel pdiffusion 1760 -1704 1760 -1704 0 feedthrough
rlabel pdiffusion 1767 -1704 1767 -1704 0 feedthrough
rlabel pdiffusion 1774 -1704 1774 -1704 0 feedthrough
rlabel pdiffusion 1781 -1704 1781 -1704 0 feedthrough
rlabel pdiffusion 1788 -1704 1788 -1704 0 feedthrough
rlabel pdiffusion 1795 -1704 1795 -1704 0 feedthrough
rlabel pdiffusion 1802 -1704 1802 -1704 0 feedthrough
rlabel pdiffusion 1809 -1704 1809 -1704 0 cellNo=194
rlabel pdiffusion 1816 -1704 1816 -1704 0 feedthrough
rlabel pdiffusion 1823 -1704 1823 -1704 0 feedthrough
rlabel pdiffusion 1830 -1704 1830 -1704 0 feedthrough
rlabel pdiffusion 1837 -1704 1837 -1704 0 feedthrough
rlabel pdiffusion 1844 -1704 1844 -1704 0 feedthrough
rlabel pdiffusion 1851 -1704 1851 -1704 0 feedthrough
rlabel pdiffusion 1858 -1704 1858 -1704 0 feedthrough
rlabel pdiffusion 1865 -1704 1865 -1704 0 feedthrough
rlabel pdiffusion 1872 -1704 1872 -1704 0 feedthrough
rlabel pdiffusion 1879 -1704 1879 -1704 0 feedthrough
rlabel pdiffusion 1886 -1704 1886 -1704 0 feedthrough
rlabel pdiffusion 1893 -1704 1893 -1704 0 feedthrough
rlabel pdiffusion 1900 -1704 1900 -1704 0 feedthrough
rlabel pdiffusion 1907 -1704 1907 -1704 0 feedthrough
rlabel pdiffusion 1914 -1704 1914 -1704 0 feedthrough
rlabel pdiffusion 1921 -1704 1921 -1704 0 feedthrough
rlabel pdiffusion 1928 -1704 1928 -1704 0 feedthrough
rlabel pdiffusion 1935 -1704 1935 -1704 0 feedthrough
rlabel pdiffusion 1942 -1704 1942 -1704 0 feedthrough
rlabel pdiffusion 1949 -1704 1949 -1704 0 feedthrough
rlabel pdiffusion 1956 -1704 1956 -1704 0 feedthrough
rlabel pdiffusion 1963 -1704 1963 -1704 0 feedthrough
rlabel pdiffusion 1970 -1704 1970 -1704 0 feedthrough
rlabel pdiffusion 1977 -1704 1977 -1704 0 feedthrough
rlabel pdiffusion 1984 -1704 1984 -1704 0 feedthrough
rlabel pdiffusion 1991 -1704 1991 -1704 0 feedthrough
rlabel pdiffusion 1998 -1704 1998 -1704 0 feedthrough
rlabel pdiffusion 2005 -1704 2005 -1704 0 feedthrough
rlabel pdiffusion 2012 -1704 2012 -1704 0 feedthrough
rlabel pdiffusion 2019 -1704 2019 -1704 0 feedthrough
rlabel pdiffusion 2026 -1704 2026 -1704 0 feedthrough
rlabel pdiffusion 2033 -1704 2033 -1704 0 feedthrough
rlabel pdiffusion 2040 -1704 2040 -1704 0 feedthrough
rlabel pdiffusion 2047 -1704 2047 -1704 0 feedthrough
rlabel pdiffusion 2054 -1704 2054 -1704 0 feedthrough
rlabel pdiffusion 2061 -1704 2061 -1704 0 feedthrough
rlabel pdiffusion 2068 -1704 2068 -1704 0 feedthrough
rlabel pdiffusion 2075 -1704 2075 -1704 0 feedthrough
rlabel pdiffusion 2082 -1704 2082 -1704 0 feedthrough
rlabel pdiffusion 2089 -1704 2089 -1704 0 feedthrough
rlabel pdiffusion 2096 -1704 2096 -1704 0 feedthrough
rlabel pdiffusion 2103 -1704 2103 -1704 0 feedthrough
rlabel pdiffusion 2110 -1704 2110 -1704 0 feedthrough
rlabel pdiffusion 2117 -1704 2117 -1704 0 feedthrough
rlabel pdiffusion 2124 -1704 2124 -1704 0 feedthrough
rlabel pdiffusion 2131 -1704 2131 -1704 0 feedthrough
rlabel pdiffusion 2138 -1704 2138 -1704 0 feedthrough
rlabel pdiffusion 2145 -1704 2145 -1704 0 feedthrough
rlabel pdiffusion 2152 -1704 2152 -1704 0 feedthrough
rlabel pdiffusion 2159 -1704 2159 -1704 0 feedthrough
rlabel pdiffusion 2166 -1704 2166 -1704 0 feedthrough
rlabel pdiffusion 2173 -1704 2173 -1704 0 feedthrough
rlabel pdiffusion 2180 -1704 2180 -1704 0 feedthrough
rlabel pdiffusion 2187 -1704 2187 -1704 0 feedthrough
rlabel pdiffusion 2194 -1704 2194 -1704 0 feedthrough
rlabel pdiffusion 2201 -1704 2201 -1704 0 feedthrough
rlabel pdiffusion 2208 -1704 2208 -1704 0 feedthrough
rlabel pdiffusion 2215 -1704 2215 -1704 0 feedthrough
rlabel pdiffusion 2222 -1704 2222 -1704 0 feedthrough
rlabel pdiffusion 2229 -1704 2229 -1704 0 feedthrough
rlabel pdiffusion 2236 -1704 2236 -1704 0 feedthrough
rlabel pdiffusion 2243 -1704 2243 -1704 0 feedthrough
rlabel pdiffusion 2250 -1704 2250 -1704 0 feedthrough
rlabel pdiffusion 2257 -1704 2257 -1704 0 feedthrough
rlabel pdiffusion 2264 -1704 2264 -1704 0 feedthrough
rlabel pdiffusion 2271 -1704 2271 -1704 0 feedthrough
rlabel pdiffusion 2278 -1704 2278 -1704 0 feedthrough
rlabel pdiffusion 2285 -1704 2285 -1704 0 feedthrough
rlabel pdiffusion 2292 -1704 2292 -1704 0 feedthrough
rlabel pdiffusion 2299 -1704 2299 -1704 0 feedthrough
rlabel pdiffusion 2306 -1704 2306 -1704 0 feedthrough
rlabel pdiffusion 2313 -1704 2313 -1704 0 feedthrough
rlabel pdiffusion 2320 -1704 2320 -1704 0 feedthrough
rlabel pdiffusion 2327 -1704 2327 -1704 0 feedthrough
rlabel pdiffusion 2334 -1704 2334 -1704 0 feedthrough
rlabel pdiffusion 2341 -1704 2341 -1704 0 feedthrough
rlabel pdiffusion 2348 -1704 2348 -1704 0 feedthrough
rlabel pdiffusion 2355 -1704 2355 -1704 0 feedthrough
rlabel pdiffusion 2362 -1704 2362 -1704 0 feedthrough
rlabel pdiffusion 2369 -1704 2369 -1704 0 feedthrough
rlabel pdiffusion 2376 -1704 2376 -1704 0 feedthrough
rlabel pdiffusion 2383 -1704 2383 -1704 0 feedthrough
rlabel pdiffusion 2390 -1704 2390 -1704 0 feedthrough
rlabel pdiffusion 2397 -1704 2397 -1704 0 feedthrough
rlabel pdiffusion 2404 -1704 2404 -1704 0 feedthrough
rlabel pdiffusion 2411 -1704 2411 -1704 0 feedthrough
rlabel pdiffusion 2418 -1704 2418 -1704 0 feedthrough
rlabel pdiffusion 2425 -1704 2425 -1704 0 cellNo=707
rlabel pdiffusion 2432 -1704 2432 -1704 0 cellNo=282
rlabel pdiffusion 2439 -1704 2439 -1704 0 cellNo=516
rlabel pdiffusion 2446 -1704 2446 -1704 0 feedthrough
rlabel pdiffusion 2453 -1704 2453 -1704 0 feedthrough
rlabel pdiffusion 2495 -1704 2495 -1704 0 feedthrough
rlabel pdiffusion 3 -1855 3 -1855 0 feedthrough
rlabel pdiffusion 10 -1855 10 -1855 0 feedthrough
rlabel pdiffusion 17 -1855 17 -1855 0 feedthrough
rlabel pdiffusion 24 -1855 24 -1855 0 feedthrough
rlabel pdiffusion 31 -1855 31 -1855 0 feedthrough
rlabel pdiffusion 38 -1855 38 -1855 0 feedthrough
rlabel pdiffusion 45 -1855 45 -1855 0 cellNo=479
rlabel pdiffusion 52 -1855 52 -1855 0 feedthrough
rlabel pdiffusion 59 -1855 59 -1855 0 feedthrough
rlabel pdiffusion 66 -1855 66 -1855 0 feedthrough
rlabel pdiffusion 73 -1855 73 -1855 0 feedthrough
rlabel pdiffusion 80 -1855 80 -1855 0 feedthrough
rlabel pdiffusion 87 -1855 87 -1855 0 feedthrough
rlabel pdiffusion 94 -1855 94 -1855 0 feedthrough
rlabel pdiffusion 101 -1855 101 -1855 0 feedthrough
rlabel pdiffusion 108 -1855 108 -1855 0 feedthrough
rlabel pdiffusion 115 -1855 115 -1855 0 feedthrough
rlabel pdiffusion 122 -1855 122 -1855 0 cellNo=958
rlabel pdiffusion 129 -1855 129 -1855 0 feedthrough
rlabel pdiffusion 136 -1855 136 -1855 0 feedthrough
rlabel pdiffusion 143 -1855 143 -1855 0 feedthrough
rlabel pdiffusion 150 -1855 150 -1855 0 feedthrough
rlabel pdiffusion 157 -1855 157 -1855 0 cellNo=452
rlabel pdiffusion 164 -1855 164 -1855 0 feedthrough
rlabel pdiffusion 171 -1855 171 -1855 0 feedthrough
rlabel pdiffusion 178 -1855 178 -1855 0 feedthrough
rlabel pdiffusion 185 -1855 185 -1855 0 cellNo=338
rlabel pdiffusion 192 -1855 192 -1855 0 feedthrough
rlabel pdiffusion 199 -1855 199 -1855 0 cellNo=416
rlabel pdiffusion 206 -1855 206 -1855 0 feedthrough
rlabel pdiffusion 213 -1855 213 -1855 0 feedthrough
rlabel pdiffusion 220 -1855 220 -1855 0 feedthrough
rlabel pdiffusion 227 -1855 227 -1855 0 cellNo=561
rlabel pdiffusion 234 -1855 234 -1855 0 cellNo=883
rlabel pdiffusion 241 -1855 241 -1855 0 feedthrough
rlabel pdiffusion 248 -1855 248 -1855 0 cellNo=920
rlabel pdiffusion 255 -1855 255 -1855 0 feedthrough
rlabel pdiffusion 262 -1855 262 -1855 0 feedthrough
rlabel pdiffusion 269 -1855 269 -1855 0 feedthrough
rlabel pdiffusion 276 -1855 276 -1855 0 feedthrough
rlabel pdiffusion 283 -1855 283 -1855 0 feedthrough
rlabel pdiffusion 290 -1855 290 -1855 0 feedthrough
rlabel pdiffusion 297 -1855 297 -1855 0 feedthrough
rlabel pdiffusion 304 -1855 304 -1855 0 feedthrough
rlabel pdiffusion 311 -1855 311 -1855 0 feedthrough
rlabel pdiffusion 318 -1855 318 -1855 0 feedthrough
rlabel pdiffusion 325 -1855 325 -1855 0 feedthrough
rlabel pdiffusion 332 -1855 332 -1855 0 feedthrough
rlabel pdiffusion 339 -1855 339 -1855 0 feedthrough
rlabel pdiffusion 346 -1855 346 -1855 0 feedthrough
rlabel pdiffusion 353 -1855 353 -1855 0 feedthrough
rlabel pdiffusion 360 -1855 360 -1855 0 feedthrough
rlabel pdiffusion 367 -1855 367 -1855 0 feedthrough
rlabel pdiffusion 374 -1855 374 -1855 0 feedthrough
rlabel pdiffusion 381 -1855 381 -1855 0 feedthrough
rlabel pdiffusion 388 -1855 388 -1855 0 feedthrough
rlabel pdiffusion 395 -1855 395 -1855 0 feedthrough
rlabel pdiffusion 402 -1855 402 -1855 0 feedthrough
rlabel pdiffusion 409 -1855 409 -1855 0 feedthrough
rlabel pdiffusion 416 -1855 416 -1855 0 feedthrough
rlabel pdiffusion 423 -1855 423 -1855 0 feedthrough
rlabel pdiffusion 430 -1855 430 -1855 0 cellNo=17
rlabel pdiffusion 437 -1855 437 -1855 0 feedthrough
rlabel pdiffusion 444 -1855 444 -1855 0 cellNo=443
rlabel pdiffusion 451 -1855 451 -1855 0 feedthrough
rlabel pdiffusion 458 -1855 458 -1855 0 feedthrough
rlabel pdiffusion 465 -1855 465 -1855 0 feedthrough
rlabel pdiffusion 472 -1855 472 -1855 0 feedthrough
rlabel pdiffusion 479 -1855 479 -1855 0 feedthrough
rlabel pdiffusion 486 -1855 486 -1855 0 feedthrough
rlabel pdiffusion 493 -1855 493 -1855 0 feedthrough
rlabel pdiffusion 500 -1855 500 -1855 0 feedthrough
rlabel pdiffusion 507 -1855 507 -1855 0 feedthrough
rlabel pdiffusion 514 -1855 514 -1855 0 cellNo=877
rlabel pdiffusion 521 -1855 521 -1855 0 feedthrough
rlabel pdiffusion 528 -1855 528 -1855 0 feedthrough
rlabel pdiffusion 535 -1855 535 -1855 0 feedthrough
rlabel pdiffusion 542 -1855 542 -1855 0 feedthrough
rlabel pdiffusion 549 -1855 549 -1855 0 feedthrough
rlabel pdiffusion 556 -1855 556 -1855 0 feedthrough
rlabel pdiffusion 563 -1855 563 -1855 0 cellNo=491
rlabel pdiffusion 570 -1855 570 -1855 0 feedthrough
rlabel pdiffusion 577 -1855 577 -1855 0 feedthrough
rlabel pdiffusion 584 -1855 584 -1855 0 feedthrough
rlabel pdiffusion 591 -1855 591 -1855 0 feedthrough
rlabel pdiffusion 598 -1855 598 -1855 0 feedthrough
rlabel pdiffusion 605 -1855 605 -1855 0 feedthrough
rlabel pdiffusion 612 -1855 612 -1855 0 cellNo=310
rlabel pdiffusion 619 -1855 619 -1855 0 feedthrough
rlabel pdiffusion 626 -1855 626 -1855 0 feedthrough
rlabel pdiffusion 633 -1855 633 -1855 0 cellNo=180
rlabel pdiffusion 640 -1855 640 -1855 0 feedthrough
rlabel pdiffusion 647 -1855 647 -1855 0 cellNo=998
rlabel pdiffusion 654 -1855 654 -1855 0 feedthrough
rlabel pdiffusion 661 -1855 661 -1855 0 feedthrough
rlabel pdiffusion 668 -1855 668 -1855 0 feedthrough
rlabel pdiffusion 675 -1855 675 -1855 0 feedthrough
rlabel pdiffusion 682 -1855 682 -1855 0 feedthrough
rlabel pdiffusion 689 -1855 689 -1855 0 feedthrough
rlabel pdiffusion 696 -1855 696 -1855 0 feedthrough
rlabel pdiffusion 703 -1855 703 -1855 0 feedthrough
rlabel pdiffusion 710 -1855 710 -1855 0 feedthrough
rlabel pdiffusion 717 -1855 717 -1855 0 feedthrough
rlabel pdiffusion 724 -1855 724 -1855 0 cellNo=843
rlabel pdiffusion 731 -1855 731 -1855 0 cellNo=94
rlabel pdiffusion 738 -1855 738 -1855 0 cellNo=955
rlabel pdiffusion 745 -1855 745 -1855 0 feedthrough
rlabel pdiffusion 752 -1855 752 -1855 0 feedthrough
rlabel pdiffusion 759 -1855 759 -1855 0 feedthrough
rlabel pdiffusion 766 -1855 766 -1855 0 feedthrough
rlabel pdiffusion 773 -1855 773 -1855 0 feedthrough
rlabel pdiffusion 780 -1855 780 -1855 0 feedthrough
rlabel pdiffusion 787 -1855 787 -1855 0 feedthrough
rlabel pdiffusion 794 -1855 794 -1855 0 feedthrough
rlabel pdiffusion 801 -1855 801 -1855 0 cellNo=459
rlabel pdiffusion 808 -1855 808 -1855 0 feedthrough
rlabel pdiffusion 815 -1855 815 -1855 0 feedthrough
rlabel pdiffusion 822 -1855 822 -1855 0 feedthrough
rlabel pdiffusion 829 -1855 829 -1855 0 feedthrough
rlabel pdiffusion 836 -1855 836 -1855 0 feedthrough
rlabel pdiffusion 843 -1855 843 -1855 0 feedthrough
rlabel pdiffusion 850 -1855 850 -1855 0 cellNo=311
rlabel pdiffusion 857 -1855 857 -1855 0 feedthrough
rlabel pdiffusion 864 -1855 864 -1855 0 feedthrough
rlabel pdiffusion 871 -1855 871 -1855 0 feedthrough
rlabel pdiffusion 878 -1855 878 -1855 0 feedthrough
rlabel pdiffusion 885 -1855 885 -1855 0 feedthrough
rlabel pdiffusion 892 -1855 892 -1855 0 cellNo=258
rlabel pdiffusion 899 -1855 899 -1855 0 feedthrough
rlabel pdiffusion 906 -1855 906 -1855 0 cellNo=25
rlabel pdiffusion 913 -1855 913 -1855 0 feedthrough
rlabel pdiffusion 920 -1855 920 -1855 0 feedthrough
rlabel pdiffusion 927 -1855 927 -1855 0 feedthrough
rlabel pdiffusion 934 -1855 934 -1855 0 feedthrough
rlabel pdiffusion 941 -1855 941 -1855 0 cellNo=351
rlabel pdiffusion 948 -1855 948 -1855 0 feedthrough
rlabel pdiffusion 955 -1855 955 -1855 0 cellNo=723
rlabel pdiffusion 962 -1855 962 -1855 0 feedthrough
rlabel pdiffusion 969 -1855 969 -1855 0 feedthrough
rlabel pdiffusion 976 -1855 976 -1855 0 feedthrough
rlabel pdiffusion 983 -1855 983 -1855 0 feedthrough
rlabel pdiffusion 990 -1855 990 -1855 0 feedthrough
rlabel pdiffusion 997 -1855 997 -1855 0 feedthrough
rlabel pdiffusion 1004 -1855 1004 -1855 0 feedthrough
rlabel pdiffusion 1011 -1855 1011 -1855 0 feedthrough
rlabel pdiffusion 1018 -1855 1018 -1855 0 feedthrough
rlabel pdiffusion 1025 -1855 1025 -1855 0 feedthrough
rlabel pdiffusion 1032 -1855 1032 -1855 0 feedthrough
rlabel pdiffusion 1039 -1855 1039 -1855 0 feedthrough
rlabel pdiffusion 1046 -1855 1046 -1855 0 feedthrough
rlabel pdiffusion 1053 -1855 1053 -1855 0 feedthrough
rlabel pdiffusion 1060 -1855 1060 -1855 0 feedthrough
rlabel pdiffusion 1067 -1855 1067 -1855 0 feedthrough
rlabel pdiffusion 1074 -1855 1074 -1855 0 feedthrough
rlabel pdiffusion 1081 -1855 1081 -1855 0 feedthrough
rlabel pdiffusion 1088 -1855 1088 -1855 0 feedthrough
rlabel pdiffusion 1095 -1855 1095 -1855 0 feedthrough
rlabel pdiffusion 1102 -1855 1102 -1855 0 feedthrough
rlabel pdiffusion 1109 -1855 1109 -1855 0 feedthrough
rlabel pdiffusion 1116 -1855 1116 -1855 0 feedthrough
rlabel pdiffusion 1123 -1855 1123 -1855 0 feedthrough
rlabel pdiffusion 1130 -1855 1130 -1855 0 feedthrough
rlabel pdiffusion 1137 -1855 1137 -1855 0 cellNo=6
rlabel pdiffusion 1144 -1855 1144 -1855 0 feedthrough
rlabel pdiffusion 1151 -1855 1151 -1855 0 feedthrough
rlabel pdiffusion 1158 -1855 1158 -1855 0 feedthrough
rlabel pdiffusion 1165 -1855 1165 -1855 0 feedthrough
rlabel pdiffusion 1172 -1855 1172 -1855 0 feedthrough
rlabel pdiffusion 1179 -1855 1179 -1855 0 cellNo=471
rlabel pdiffusion 1186 -1855 1186 -1855 0 feedthrough
rlabel pdiffusion 1193 -1855 1193 -1855 0 feedthrough
rlabel pdiffusion 1200 -1855 1200 -1855 0 feedthrough
rlabel pdiffusion 1207 -1855 1207 -1855 0 cellNo=951
rlabel pdiffusion 1214 -1855 1214 -1855 0 feedthrough
rlabel pdiffusion 1221 -1855 1221 -1855 0 feedthrough
rlabel pdiffusion 1228 -1855 1228 -1855 0 feedthrough
rlabel pdiffusion 1235 -1855 1235 -1855 0 feedthrough
rlabel pdiffusion 1242 -1855 1242 -1855 0 feedthrough
rlabel pdiffusion 1249 -1855 1249 -1855 0 feedthrough
rlabel pdiffusion 1256 -1855 1256 -1855 0 feedthrough
rlabel pdiffusion 1263 -1855 1263 -1855 0 feedthrough
rlabel pdiffusion 1270 -1855 1270 -1855 0 feedthrough
rlabel pdiffusion 1277 -1855 1277 -1855 0 cellNo=829
rlabel pdiffusion 1284 -1855 1284 -1855 0 feedthrough
rlabel pdiffusion 1291 -1855 1291 -1855 0 cellNo=511
rlabel pdiffusion 1298 -1855 1298 -1855 0 feedthrough
rlabel pdiffusion 1305 -1855 1305 -1855 0 cellNo=662
rlabel pdiffusion 1312 -1855 1312 -1855 0 feedthrough
rlabel pdiffusion 1319 -1855 1319 -1855 0 feedthrough
rlabel pdiffusion 1326 -1855 1326 -1855 0 feedthrough
rlabel pdiffusion 1333 -1855 1333 -1855 0 feedthrough
rlabel pdiffusion 1340 -1855 1340 -1855 0 feedthrough
rlabel pdiffusion 1347 -1855 1347 -1855 0 feedthrough
rlabel pdiffusion 1354 -1855 1354 -1855 0 feedthrough
rlabel pdiffusion 1361 -1855 1361 -1855 0 feedthrough
rlabel pdiffusion 1368 -1855 1368 -1855 0 feedthrough
rlabel pdiffusion 1375 -1855 1375 -1855 0 feedthrough
rlabel pdiffusion 1382 -1855 1382 -1855 0 feedthrough
rlabel pdiffusion 1389 -1855 1389 -1855 0 feedthrough
rlabel pdiffusion 1396 -1855 1396 -1855 0 feedthrough
rlabel pdiffusion 1403 -1855 1403 -1855 0 feedthrough
rlabel pdiffusion 1410 -1855 1410 -1855 0 feedthrough
rlabel pdiffusion 1417 -1855 1417 -1855 0 feedthrough
rlabel pdiffusion 1424 -1855 1424 -1855 0 feedthrough
rlabel pdiffusion 1431 -1855 1431 -1855 0 feedthrough
rlabel pdiffusion 1438 -1855 1438 -1855 0 cellNo=377
rlabel pdiffusion 1445 -1855 1445 -1855 0 feedthrough
rlabel pdiffusion 1452 -1855 1452 -1855 0 feedthrough
rlabel pdiffusion 1459 -1855 1459 -1855 0 feedthrough
rlabel pdiffusion 1466 -1855 1466 -1855 0 cellNo=337
rlabel pdiffusion 1473 -1855 1473 -1855 0 feedthrough
rlabel pdiffusion 1480 -1855 1480 -1855 0 feedthrough
rlabel pdiffusion 1487 -1855 1487 -1855 0 feedthrough
rlabel pdiffusion 1494 -1855 1494 -1855 0 feedthrough
rlabel pdiffusion 1501 -1855 1501 -1855 0 feedthrough
rlabel pdiffusion 1508 -1855 1508 -1855 0 cellNo=217
rlabel pdiffusion 1515 -1855 1515 -1855 0 feedthrough
rlabel pdiffusion 1522 -1855 1522 -1855 0 feedthrough
rlabel pdiffusion 1529 -1855 1529 -1855 0 feedthrough
rlabel pdiffusion 1536 -1855 1536 -1855 0 feedthrough
rlabel pdiffusion 1543 -1855 1543 -1855 0 feedthrough
rlabel pdiffusion 1550 -1855 1550 -1855 0 feedthrough
rlabel pdiffusion 1557 -1855 1557 -1855 0 feedthrough
rlabel pdiffusion 1564 -1855 1564 -1855 0 feedthrough
rlabel pdiffusion 1571 -1855 1571 -1855 0 feedthrough
rlabel pdiffusion 1578 -1855 1578 -1855 0 feedthrough
rlabel pdiffusion 1585 -1855 1585 -1855 0 feedthrough
rlabel pdiffusion 1592 -1855 1592 -1855 0 feedthrough
rlabel pdiffusion 1599 -1855 1599 -1855 0 feedthrough
rlabel pdiffusion 1606 -1855 1606 -1855 0 feedthrough
rlabel pdiffusion 1613 -1855 1613 -1855 0 feedthrough
rlabel pdiffusion 1620 -1855 1620 -1855 0 feedthrough
rlabel pdiffusion 1627 -1855 1627 -1855 0 cellNo=363
rlabel pdiffusion 1634 -1855 1634 -1855 0 feedthrough
rlabel pdiffusion 1641 -1855 1641 -1855 0 feedthrough
rlabel pdiffusion 1648 -1855 1648 -1855 0 feedthrough
rlabel pdiffusion 1655 -1855 1655 -1855 0 feedthrough
rlabel pdiffusion 1662 -1855 1662 -1855 0 cellNo=824
rlabel pdiffusion 1669 -1855 1669 -1855 0 feedthrough
rlabel pdiffusion 1676 -1855 1676 -1855 0 feedthrough
rlabel pdiffusion 1683 -1855 1683 -1855 0 feedthrough
rlabel pdiffusion 1690 -1855 1690 -1855 0 feedthrough
rlabel pdiffusion 1697 -1855 1697 -1855 0 feedthrough
rlabel pdiffusion 1704 -1855 1704 -1855 0 feedthrough
rlabel pdiffusion 1711 -1855 1711 -1855 0 feedthrough
rlabel pdiffusion 1718 -1855 1718 -1855 0 feedthrough
rlabel pdiffusion 1725 -1855 1725 -1855 0 feedthrough
rlabel pdiffusion 1732 -1855 1732 -1855 0 feedthrough
rlabel pdiffusion 1739 -1855 1739 -1855 0 feedthrough
rlabel pdiffusion 1746 -1855 1746 -1855 0 feedthrough
rlabel pdiffusion 1753 -1855 1753 -1855 0 feedthrough
rlabel pdiffusion 1760 -1855 1760 -1855 0 feedthrough
rlabel pdiffusion 1767 -1855 1767 -1855 0 feedthrough
rlabel pdiffusion 1774 -1855 1774 -1855 0 feedthrough
rlabel pdiffusion 1781 -1855 1781 -1855 0 feedthrough
rlabel pdiffusion 1788 -1855 1788 -1855 0 feedthrough
rlabel pdiffusion 1795 -1855 1795 -1855 0 feedthrough
rlabel pdiffusion 1802 -1855 1802 -1855 0 feedthrough
rlabel pdiffusion 1809 -1855 1809 -1855 0 feedthrough
rlabel pdiffusion 1816 -1855 1816 -1855 0 feedthrough
rlabel pdiffusion 1823 -1855 1823 -1855 0 feedthrough
rlabel pdiffusion 1830 -1855 1830 -1855 0 feedthrough
rlabel pdiffusion 1837 -1855 1837 -1855 0 feedthrough
rlabel pdiffusion 1844 -1855 1844 -1855 0 feedthrough
rlabel pdiffusion 1851 -1855 1851 -1855 0 cellNo=748
rlabel pdiffusion 1858 -1855 1858 -1855 0 feedthrough
rlabel pdiffusion 1865 -1855 1865 -1855 0 cellNo=262
rlabel pdiffusion 1872 -1855 1872 -1855 0 feedthrough
rlabel pdiffusion 1879 -1855 1879 -1855 0 feedthrough
rlabel pdiffusion 1886 -1855 1886 -1855 0 feedthrough
rlabel pdiffusion 1893 -1855 1893 -1855 0 feedthrough
rlabel pdiffusion 1900 -1855 1900 -1855 0 feedthrough
rlabel pdiffusion 1907 -1855 1907 -1855 0 feedthrough
rlabel pdiffusion 1914 -1855 1914 -1855 0 feedthrough
rlabel pdiffusion 1921 -1855 1921 -1855 0 feedthrough
rlabel pdiffusion 1928 -1855 1928 -1855 0 feedthrough
rlabel pdiffusion 1935 -1855 1935 -1855 0 feedthrough
rlabel pdiffusion 1942 -1855 1942 -1855 0 feedthrough
rlabel pdiffusion 1949 -1855 1949 -1855 0 feedthrough
rlabel pdiffusion 1956 -1855 1956 -1855 0 feedthrough
rlabel pdiffusion 1963 -1855 1963 -1855 0 feedthrough
rlabel pdiffusion 1970 -1855 1970 -1855 0 feedthrough
rlabel pdiffusion 1977 -1855 1977 -1855 0 feedthrough
rlabel pdiffusion 1984 -1855 1984 -1855 0 feedthrough
rlabel pdiffusion 1991 -1855 1991 -1855 0 feedthrough
rlabel pdiffusion 1998 -1855 1998 -1855 0 feedthrough
rlabel pdiffusion 2005 -1855 2005 -1855 0 feedthrough
rlabel pdiffusion 2012 -1855 2012 -1855 0 feedthrough
rlabel pdiffusion 2019 -1855 2019 -1855 0 feedthrough
rlabel pdiffusion 2026 -1855 2026 -1855 0 feedthrough
rlabel pdiffusion 2033 -1855 2033 -1855 0 feedthrough
rlabel pdiffusion 2040 -1855 2040 -1855 0 feedthrough
rlabel pdiffusion 2047 -1855 2047 -1855 0 feedthrough
rlabel pdiffusion 2054 -1855 2054 -1855 0 feedthrough
rlabel pdiffusion 2061 -1855 2061 -1855 0 feedthrough
rlabel pdiffusion 2068 -1855 2068 -1855 0 feedthrough
rlabel pdiffusion 2075 -1855 2075 -1855 0 feedthrough
rlabel pdiffusion 2082 -1855 2082 -1855 0 feedthrough
rlabel pdiffusion 2089 -1855 2089 -1855 0 feedthrough
rlabel pdiffusion 2096 -1855 2096 -1855 0 feedthrough
rlabel pdiffusion 2103 -1855 2103 -1855 0 feedthrough
rlabel pdiffusion 2110 -1855 2110 -1855 0 feedthrough
rlabel pdiffusion 2117 -1855 2117 -1855 0 feedthrough
rlabel pdiffusion 2124 -1855 2124 -1855 0 feedthrough
rlabel pdiffusion 2131 -1855 2131 -1855 0 feedthrough
rlabel pdiffusion 2138 -1855 2138 -1855 0 feedthrough
rlabel pdiffusion 2145 -1855 2145 -1855 0 feedthrough
rlabel pdiffusion 2152 -1855 2152 -1855 0 feedthrough
rlabel pdiffusion 2159 -1855 2159 -1855 0 feedthrough
rlabel pdiffusion 2166 -1855 2166 -1855 0 feedthrough
rlabel pdiffusion 2173 -1855 2173 -1855 0 feedthrough
rlabel pdiffusion 2180 -1855 2180 -1855 0 feedthrough
rlabel pdiffusion 2187 -1855 2187 -1855 0 feedthrough
rlabel pdiffusion 2194 -1855 2194 -1855 0 feedthrough
rlabel pdiffusion 2201 -1855 2201 -1855 0 feedthrough
rlabel pdiffusion 2208 -1855 2208 -1855 0 feedthrough
rlabel pdiffusion 2215 -1855 2215 -1855 0 feedthrough
rlabel pdiffusion 2222 -1855 2222 -1855 0 feedthrough
rlabel pdiffusion 2229 -1855 2229 -1855 0 feedthrough
rlabel pdiffusion 2236 -1855 2236 -1855 0 feedthrough
rlabel pdiffusion 2243 -1855 2243 -1855 0 feedthrough
rlabel pdiffusion 2250 -1855 2250 -1855 0 feedthrough
rlabel pdiffusion 2257 -1855 2257 -1855 0 feedthrough
rlabel pdiffusion 2264 -1855 2264 -1855 0 feedthrough
rlabel pdiffusion 2271 -1855 2271 -1855 0 feedthrough
rlabel pdiffusion 2278 -1855 2278 -1855 0 feedthrough
rlabel pdiffusion 2285 -1855 2285 -1855 0 feedthrough
rlabel pdiffusion 2292 -1855 2292 -1855 0 feedthrough
rlabel pdiffusion 2299 -1855 2299 -1855 0 feedthrough
rlabel pdiffusion 2306 -1855 2306 -1855 0 feedthrough
rlabel pdiffusion 2313 -1855 2313 -1855 0 feedthrough
rlabel pdiffusion 2320 -1855 2320 -1855 0 feedthrough
rlabel pdiffusion 2327 -1855 2327 -1855 0 feedthrough
rlabel pdiffusion 2334 -1855 2334 -1855 0 feedthrough
rlabel pdiffusion 2341 -1855 2341 -1855 0 feedthrough
rlabel pdiffusion 2348 -1855 2348 -1855 0 feedthrough
rlabel pdiffusion 2355 -1855 2355 -1855 0 feedthrough
rlabel pdiffusion 2362 -1855 2362 -1855 0 feedthrough
rlabel pdiffusion 2369 -1855 2369 -1855 0 feedthrough
rlabel pdiffusion 2376 -1855 2376 -1855 0 feedthrough
rlabel pdiffusion 2383 -1855 2383 -1855 0 feedthrough
rlabel pdiffusion 2390 -1855 2390 -1855 0 feedthrough
rlabel pdiffusion 2397 -1855 2397 -1855 0 feedthrough
rlabel pdiffusion 2404 -1855 2404 -1855 0 feedthrough
rlabel pdiffusion 2411 -1855 2411 -1855 0 feedthrough
rlabel pdiffusion 2418 -1855 2418 -1855 0 feedthrough
rlabel pdiffusion 2425 -1855 2425 -1855 0 feedthrough
rlabel pdiffusion 2432 -1855 2432 -1855 0 feedthrough
rlabel pdiffusion 2439 -1855 2439 -1855 0 feedthrough
rlabel pdiffusion 2446 -1855 2446 -1855 0 feedthrough
rlabel pdiffusion 2453 -1855 2453 -1855 0 feedthrough
rlabel pdiffusion 2460 -1855 2460 -1855 0 feedthrough
rlabel pdiffusion 2467 -1855 2467 -1855 0 cellNo=280
rlabel pdiffusion 2474 -1855 2474 -1855 0 cellNo=571
rlabel pdiffusion 3 -2030 3 -2030 0 feedthrough
rlabel pdiffusion 10 -2030 10 -2030 0 feedthrough
rlabel pdiffusion 17 -2030 17 -2030 0 feedthrough
rlabel pdiffusion 24 -2030 24 -2030 0 feedthrough
rlabel pdiffusion 31 -2030 31 -2030 0 feedthrough
rlabel pdiffusion 38 -2030 38 -2030 0 feedthrough
rlabel pdiffusion 45 -2030 45 -2030 0 feedthrough
rlabel pdiffusion 52 -2030 52 -2030 0 cellNo=239
rlabel pdiffusion 59 -2030 59 -2030 0 feedthrough
rlabel pdiffusion 66 -2030 66 -2030 0 feedthrough
rlabel pdiffusion 73 -2030 73 -2030 0 feedthrough
rlabel pdiffusion 80 -2030 80 -2030 0 feedthrough
rlabel pdiffusion 87 -2030 87 -2030 0 cellNo=335
rlabel pdiffusion 94 -2030 94 -2030 0 feedthrough
rlabel pdiffusion 101 -2030 101 -2030 0 cellNo=154
rlabel pdiffusion 108 -2030 108 -2030 0 feedthrough
rlabel pdiffusion 115 -2030 115 -2030 0 feedthrough
rlabel pdiffusion 122 -2030 122 -2030 0 feedthrough
rlabel pdiffusion 129 -2030 129 -2030 0 cellNo=37
rlabel pdiffusion 136 -2030 136 -2030 0 feedthrough
rlabel pdiffusion 143 -2030 143 -2030 0 feedthrough
rlabel pdiffusion 150 -2030 150 -2030 0 feedthrough
rlabel pdiffusion 157 -2030 157 -2030 0 cellNo=32
rlabel pdiffusion 164 -2030 164 -2030 0 feedthrough
rlabel pdiffusion 171 -2030 171 -2030 0 cellNo=796
rlabel pdiffusion 178 -2030 178 -2030 0 feedthrough
rlabel pdiffusion 185 -2030 185 -2030 0 feedthrough
rlabel pdiffusion 192 -2030 192 -2030 0 cellNo=741
rlabel pdiffusion 199 -2030 199 -2030 0 feedthrough
rlabel pdiffusion 206 -2030 206 -2030 0 feedthrough
rlabel pdiffusion 213 -2030 213 -2030 0 cellNo=130
rlabel pdiffusion 220 -2030 220 -2030 0 feedthrough
rlabel pdiffusion 227 -2030 227 -2030 0 feedthrough
rlabel pdiffusion 234 -2030 234 -2030 0 feedthrough
rlabel pdiffusion 241 -2030 241 -2030 0 feedthrough
rlabel pdiffusion 248 -2030 248 -2030 0 feedthrough
rlabel pdiffusion 255 -2030 255 -2030 0 feedthrough
rlabel pdiffusion 262 -2030 262 -2030 0 feedthrough
rlabel pdiffusion 269 -2030 269 -2030 0 feedthrough
rlabel pdiffusion 276 -2030 276 -2030 0 feedthrough
rlabel pdiffusion 283 -2030 283 -2030 0 feedthrough
rlabel pdiffusion 290 -2030 290 -2030 0 feedthrough
rlabel pdiffusion 297 -2030 297 -2030 0 feedthrough
rlabel pdiffusion 304 -2030 304 -2030 0 feedthrough
rlabel pdiffusion 311 -2030 311 -2030 0 feedthrough
rlabel pdiffusion 318 -2030 318 -2030 0 feedthrough
rlabel pdiffusion 325 -2030 325 -2030 0 feedthrough
rlabel pdiffusion 332 -2030 332 -2030 0 feedthrough
rlabel pdiffusion 339 -2030 339 -2030 0 feedthrough
rlabel pdiffusion 346 -2030 346 -2030 0 feedthrough
rlabel pdiffusion 353 -2030 353 -2030 0 feedthrough
rlabel pdiffusion 360 -2030 360 -2030 0 feedthrough
rlabel pdiffusion 367 -2030 367 -2030 0 feedthrough
rlabel pdiffusion 374 -2030 374 -2030 0 feedthrough
rlabel pdiffusion 381 -2030 381 -2030 0 feedthrough
rlabel pdiffusion 388 -2030 388 -2030 0 feedthrough
rlabel pdiffusion 395 -2030 395 -2030 0 feedthrough
rlabel pdiffusion 402 -2030 402 -2030 0 feedthrough
rlabel pdiffusion 409 -2030 409 -2030 0 feedthrough
rlabel pdiffusion 416 -2030 416 -2030 0 feedthrough
rlabel pdiffusion 423 -2030 423 -2030 0 feedthrough
rlabel pdiffusion 430 -2030 430 -2030 0 feedthrough
rlabel pdiffusion 437 -2030 437 -2030 0 feedthrough
rlabel pdiffusion 444 -2030 444 -2030 0 feedthrough
rlabel pdiffusion 451 -2030 451 -2030 0 feedthrough
rlabel pdiffusion 458 -2030 458 -2030 0 feedthrough
rlabel pdiffusion 465 -2030 465 -2030 0 feedthrough
rlabel pdiffusion 472 -2030 472 -2030 0 feedthrough
rlabel pdiffusion 479 -2030 479 -2030 0 feedthrough
rlabel pdiffusion 486 -2030 486 -2030 0 feedthrough
rlabel pdiffusion 493 -2030 493 -2030 0 feedthrough
rlabel pdiffusion 500 -2030 500 -2030 0 feedthrough
rlabel pdiffusion 507 -2030 507 -2030 0 feedthrough
rlabel pdiffusion 514 -2030 514 -2030 0 feedthrough
rlabel pdiffusion 521 -2030 521 -2030 0 feedthrough
rlabel pdiffusion 528 -2030 528 -2030 0 feedthrough
rlabel pdiffusion 535 -2030 535 -2030 0 feedthrough
rlabel pdiffusion 542 -2030 542 -2030 0 cellNo=906
rlabel pdiffusion 549 -2030 549 -2030 0 feedthrough
rlabel pdiffusion 556 -2030 556 -2030 0 feedthrough
rlabel pdiffusion 563 -2030 563 -2030 0 feedthrough
rlabel pdiffusion 570 -2030 570 -2030 0 feedthrough
rlabel pdiffusion 577 -2030 577 -2030 0 feedthrough
rlabel pdiffusion 584 -2030 584 -2030 0 cellNo=150
rlabel pdiffusion 591 -2030 591 -2030 0 feedthrough
rlabel pdiffusion 598 -2030 598 -2030 0 feedthrough
rlabel pdiffusion 605 -2030 605 -2030 0 feedthrough
rlabel pdiffusion 612 -2030 612 -2030 0 feedthrough
rlabel pdiffusion 619 -2030 619 -2030 0 feedthrough
rlabel pdiffusion 626 -2030 626 -2030 0 feedthrough
rlabel pdiffusion 633 -2030 633 -2030 0 cellNo=24
rlabel pdiffusion 640 -2030 640 -2030 0 feedthrough
rlabel pdiffusion 647 -2030 647 -2030 0 feedthrough
rlabel pdiffusion 654 -2030 654 -2030 0 feedthrough
rlabel pdiffusion 661 -2030 661 -2030 0 feedthrough
rlabel pdiffusion 668 -2030 668 -2030 0 feedthrough
rlabel pdiffusion 675 -2030 675 -2030 0 feedthrough
rlabel pdiffusion 682 -2030 682 -2030 0 feedthrough
rlabel pdiffusion 689 -2030 689 -2030 0 feedthrough
rlabel pdiffusion 696 -2030 696 -2030 0 feedthrough
rlabel pdiffusion 703 -2030 703 -2030 0 feedthrough
rlabel pdiffusion 710 -2030 710 -2030 0 feedthrough
rlabel pdiffusion 717 -2030 717 -2030 0 feedthrough
rlabel pdiffusion 724 -2030 724 -2030 0 feedthrough
rlabel pdiffusion 731 -2030 731 -2030 0 feedthrough
rlabel pdiffusion 738 -2030 738 -2030 0 cellNo=7
rlabel pdiffusion 745 -2030 745 -2030 0 feedthrough
rlabel pdiffusion 752 -2030 752 -2030 0 feedthrough
rlabel pdiffusion 759 -2030 759 -2030 0 feedthrough
rlabel pdiffusion 766 -2030 766 -2030 0 feedthrough
rlabel pdiffusion 773 -2030 773 -2030 0 feedthrough
rlabel pdiffusion 780 -2030 780 -2030 0 cellNo=586
rlabel pdiffusion 787 -2030 787 -2030 0 feedthrough
rlabel pdiffusion 794 -2030 794 -2030 0 feedthrough
rlabel pdiffusion 801 -2030 801 -2030 0 cellNo=930
rlabel pdiffusion 808 -2030 808 -2030 0 feedthrough
rlabel pdiffusion 815 -2030 815 -2030 0 feedthrough
rlabel pdiffusion 822 -2030 822 -2030 0 feedthrough
rlabel pdiffusion 829 -2030 829 -2030 0 cellNo=760
rlabel pdiffusion 836 -2030 836 -2030 0 feedthrough
rlabel pdiffusion 843 -2030 843 -2030 0 feedthrough
rlabel pdiffusion 850 -2030 850 -2030 0 feedthrough
rlabel pdiffusion 857 -2030 857 -2030 0 feedthrough
rlabel pdiffusion 864 -2030 864 -2030 0 feedthrough
rlabel pdiffusion 871 -2030 871 -2030 0 feedthrough
rlabel pdiffusion 878 -2030 878 -2030 0 feedthrough
rlabel pdiffusion 885 -2030 885 -2030 0 feedthrough
rlabel pdiffusion 892 -2030 892 -2030 0 feedthrough
rlabel pdiffusion 899 -2030 899 -2030 0 feedthrough
rlabel pdiffusion 906 -2030 906 -2030 0 feedthrough
rlabel pdiffusion 913 -2030 913 -2030 0 feedthrough
rlabel pdiffusion 920 -2030 920 -2030 0 cellNo=708
rlabel pdiffusion 927 -2030 927 -2030 0 feedthrough
rlabel pdiffusion 934 -2030 934 -2030 0 feedthrough
rlabel pdiffusion 941 -2030 941 -2030 0 feedthrough
rlabel pdiffusion 948 -2030 948 -2030 0 feedthrough
rlabel pdiffusion 955 -2030 955 -2030 0 cellNo=654
rlabel pdiffusion 962 -2030 962 -2030 0 feedthrough
rlabel pdiffusion 969 -2030 969 -2030 0 feedthrough
rlabel pdiffusion 976 -2030 976 -2030 0 cellNo=598
rlabel pdiffusion 983 -2030 983 -2030 0 feedthrough
rlabel pdiffusion 990 -2030 990 -2030 0 feedthrough
rlabel pdiffusion 997 -2030 997 -2030 0 feedthrough
rlabel pdiffusion 1004 -2030 1004 -2030 0 feedthrough
rlabel pdiffusion 1011 -2030 1011 -2030 0 feedthrough
rlabel pdiffusion 1018 -2030 1018 -2030 0 feedthrough
rlabel pdiffusion 1025 -2030 1025 -2030 0 feedthrough
rlabel pdiffusion 1032 -2030 1032 -2030 0 feedthrough
rlabel pdiffusion 1039 -2030 1039 -2030 0 feedthrough
rlabel pdiffusion 1046 -2030 1046 -2030 0 feedthrough
rlabel pdiffusion 1053 -2030 1053 -2030 0 feedthrough
rlabel pdiffusion 1060 -2030 1060 -2030 0 cellNo=999
rlabel pdiffusion 1067 -2030 1067 -2030 0 feedthrough
rlabel pdiffusion 1074 -2030 1074 -2030 0 feedthrough
rlabel pdiffusion 1081 -2030 1081 -2030 0 feedthrough
rlabel pdiffusion 1088 -2030 1088 -2030 0 feedthrough
rlabel pdiffusion 1095 -2030 1095 -2030 0 feedthrough
rlabel pdiffusion 1102 -2030 1102 -2030 0 feedthrough
rlabel pdiffusion 1109 -2030 1109 -2030 0 cellNo=649
rlabel pdiffusion 1116 -2030 1116 -2030 0 feedthrough
rlabel pdiffusion 1123 -2030 1123 -2030 0 cellNo=228
rlabel pdiffusion 1130 -2030 1130 -2030 0 feedthrough
rlabel pdiffusion 1137 -2030 1137 -2030 0 feedthrough
rlabel pdiffusion 1144 -2030 1144 -2030 0 feedthrough
rlabel pdiffusion 1151 -2030 1151 -2030 0 cellNo=467
rlabel pdiffusion 1158 -2030 1158 -2030 0 feedthrough
rlabel pdiffusion 1165 -2030 1165 -2030 0 cellNo=12
rlabel pdiffusion 1172 -2030 1172 -2030 0 feedthrough
rlabel pdiffusion 1179 -2030 1179 -2030 0 feedthrough
rlabel pdiffusion 1186 -2030 1186 -2030 0 cellNo=201
rlabel pdiffusion 1193 -2030 1193 -2030 0 feedthrough
rlabel pdiffusion 1200 -2030 1200 -2030 0 feedthrough
rlabel pdiffusion 1207 -2030 1207 -2030 0 feedthrough
rlabel pdiffusion 1214 -2030 1214 -2030 0 feedthrough
rlabel pdiffusion 1221 -2030 1221 -2030 0 feedthrough
rlabel pdiffusion 1228 -2030 1228 -2030 0 cellNo=753
rlabel pdiffusion 1235 -2030 1235 -2030 0 feedthrough
rlabel pdiffusion 1242 -2030 1242 -2030 0 feedthrough
rlabel pdiffusion 1249 -2030 1249 -2030 0 feedthrough
rlabel pdiffusion 1256 -2030 1256 -2030 0 feedthrough
rlabel pdiffusion 1263 -2030 1263 -2030 0 feedthrough
rlabel pdiffusion 1270 -2030 1270 -2030 0 feedthrough
rlabel pdiffusion 1277 -2030 1277 -2030 0 feedthrough
rlabel pdiffusion 1284 -2030 1284 -2030 0 feedthrough
rlabel pdiffusion 1291 -2030 1291 -2030 0 feedthrough
rlabel pdiffusion 1298 -2030 1298 -2030 0 cellNo=861
rlabel pdiffusion 1305 -2030 1305 -2030 0 feedthrough
rlabel pdiffusion 1312 -2030 1312 -2030 0 feedthrough
rlabel pdiffusion 1319 -2030 1319 -2030 0 feedthrough
rlabel pdiffusion 1326 -2030 1326 -2030 0 feedthrough
rlabel pdiffusion 1333 -2030 1333 -2030 0 feedthrough
rlabel pdiffusion 1340 -2030 1340 -2030 0 feedthrough
rlabel pdiffusion 1347 -2030 1347 -2030 0 feedthrough
rlabel pdiffusion 1354 -2030 1354 -2030 0 feedthrough
rlabel pdiffusion 1361 -2030 1361 -2030 0 cellNo=890
rlabel pdiffusion 1368 -2030 1368 -2030 0 feedthrough
rlabel pdiffusion 1375 -2030 1375 -2030 0 feedthrough
rlabel pdiffusion 1382 -2030 1382 -2030 0 feedthrough
rlabel pdiffusion 1389 -2030 1389 -2030 0 feedthrough
rlabel pdiffusion 1396 -2030 1396 -2030 0 feedthrough
rlabel pdiffusion 1403 -2030 1403 -2030 0 feedthrough
rlabel pdiffusion 1410 -2030 1410 -2030 0 feedthrough
rlabel pdiffusion 1417 -2030 1417 -2030 0 feedthrough
rlabel pdiffusion 1424 -2030 1424 -2030 0 feedthrough
rlabel pdiffusion 1431 -2030 1431 -2030 0 feedthrough
rlabel pdiffusion 1438 -2030 1438 -2030 0 cellNo=833
rlabel pdiffusion 1445 -2030 1445 -2030 0 feedthrough
rlabel pdiffusion 1452 -2030 1452 -2030 0 feedthrough
rlabel pdiffusion 1459 -2030 1459 -2030 0 feedthrough
rlabel pdiffusion 1466 -2030 1466 -2030 0 feedthrough
rlabel pdiffusion 1473 -2030 1473 -2030 0 cellNo=585
rlabel pdiffusion 1480 -2030 1480 -2030 0 feedthrough
rlabel pdiffusion 1487 -2030 1487 -2030 0 cellNo=505
rlabel pdiffusion 1494 -2030 1494 -2030 0 cellNo=274
rlabel pdiffusion 1501 -2030 1501 -2030 0 feedthrough
rlabel pdiffusion 1508 -2030 1508 -2030 0 feedthrough
rlabel pdiffusion 1515 -2030 1515 -2030 0 feedthrough
rlabel pdiffusion 1522 -2030 1522 -2030 0 cellNo=934
rlabel pdiffusion 1529 -2030 1529 -2030 0 feedthrough
rlabel pdiffusion 1536 -2030 1536 -2030 0 cellNo=104
rlabel pdiffusion 1543 -2030 1543 -2030 0 feedthrough
rlabel pdiffusion 1550 -2030 1550 -2030 0 cellNo=454
rlabel pdiffusion 1557 -2030 1557 -2030 0 feedthrough
rlabel pdiffusion 1564 -2030 1564 -2030 0 feedthrough
rlabel pdiffusion 1571 -2030 1571 -2030 0 feedthrough
rlabel pdiffusion 1578 -2030 1578 -2030 0 feedthrough
rlabel pdiffusion 1585 -2030 1585 -2030 0 feedthrough
rlabel pdiffusion 1592 -2030 1592 -2030 0 feedthrough
rlabel pdiffusion 1599 -2030 1599 -2030 0 feedthrough
rlabel pdiffusion 1606 -2030 1606 -2030 0 feedthrough
rlabel pdiffusion 1613 -2030 1613 -2030 0 feedthrough
rlabel pdiffusion 1620 -2030 1620 -2030 0 cellNo=529
rlabel pdiffusion 1627 -2030 1627 -2030 0 feedthrough
rlabel pdiffusion 1634 -2030 1634 -2030 0 cellNo=316
rlabel pdiffusion 1641 -2030 1641 -2030 0 feedthrough
rlabel pdiffusion 1648 -2030 1648 -2030 0 feedthrough
rlabel pdiffusion 1655 -2030 1655 -2030 0 feedthrough
rlabel pdiffusion 1662 -2030 1662 -2030 0 cellNo=413
rlabel pdiffusion 1669 -2030 1669 -2030 0 feedthrough
rlabel pdiffusion 1676 -2030 1676 -2030 0 feedthrough
rlabel pdiffusion 1683 -2030 1683 -2030 0 feedthrough
rlabel pdiffusion 1690 -2030 1690 -2030 0 feedthrough
rlabel pdiffusion 1697 -2030 1697 -2030 0 feedthrough
rlabel pdiffusion 1704 -2030 1704 -2030 0 feedthrough
rlabel pdiffusion 1711 -2030 1711 -2030 0 feedthrough
rlabel pdiffusion 1718 -2030 1718 -2030 0 feedthrough
rlabel pdiffusion 1725 -2030 1725 -2030 0 feedthrough
rlabel pdiffusion 1732 -2030 1732 -2030 0 cellNo=865
rlabel pdiffusion 1739 -2030 1739 -2030 0 feedthrough
rlabel pdiffusion 1746 -2030 1746 -2030 0 feedthrough
rlabel pdiffusion 1753 -2030 1753 -2030 0 feedthrough
rlabel pdiffusion 1760 -2030 1760 -2030 0 feedthrough
rlabel pdiffusion 1767 -2030 1767 -2030 0 feedthrough
rlabel pdiffusion 1774 -2030 1774 -2030 0 feedthrough
rlabel pdiffusion 1781 -2030 1781 -2030 0 feedthrough
rlabel pdiffusion 1788 -2030 1788 -2030 0 feedthrough
rlabel pdiffusion 1795 -2030 1795 -2030 0 feedthrough
rlabel pdiffusion 1802 -2030 1802 -2030 0 feedthrough
rlabel pdiffusion 1809 -2030 1809 -2030 0 feedthrough
rlabel pdiffusion 1816 -2030 1816 -2030 0 feedthrough
rlabel pdiffusion 1823 -2030 1823 -2030 0 feedthrough
rlabel pdiffusion 1830 -2030 1830 -2030 0 feedthrough
rlabel pdiffusion 1837 -2030 1837 -2030 0 feedthrough
rlabel pdiffusion 1844 -2030 1844 -2030 0 feedthrough
rlabel pdiffusion 1851 -2030 1851 -2030 0 feedthrough
rlabel pdiffusion 1858 -2030 1858 -2030 0 feedthrough
rlabel pdiffusion 1865 -2030 1865 -2030 0 feedthrough
rlabel pdiffusion 1872 -2030 1872 -2030 0 feedthrough
rlabel pdiffusion 1879 -2030 1879 -2030 0 feedthrough
rlabel pdiffusion 1886 -2030 1886 -2030 0 feedthrough
rlabel pdiffusion 1893 -2030 1893 -2030 0 feedthrough
rlabel pdiffusion 1900 -2030 1900 -2030 0 feedthrough
rlabel pdiffusion 1907 -2030 1907 -2030 0 feedthrough
rlabel pdiffusion 1914 -2030 1914 -2030 0 feedthrough
rlabel pdiffusion 1921 -2030 1921 -2030 0 feedthrough
rlabel pdiffusion 1928 -2030 1928 -2030 0 feedthrough
rlabel pdiffusion 1935 -2030 1935 -2030 0 feedthrough
rlabel pdiffusion 1942 -2030 1942 -2030 0 feedthrough
rlabel pdiffusion 1949 -2030 1949 -2030 0 feedthrough
rlabel pdiffusion 1956 -2030 1956 -2030 0 feedthrough
rlabel pdiffusion 1963 -2030 1963 -2030 0 feedthrough
rlabel pdiffusion 1970 -2030 1970 -2030 0 feedthrough
rlabel pdiffusion 1977 -2030 1977 -2030 0 feedthrough
rlabel pdiffusion 1984 -2030 1984 -2030 0 feedthrough
rlabel pdiffusion 1991 -2030 1991 -2030 0 feedthrough
rlabel pdiffusion 1998 -2030 1998 -2030 0 feedthrough
rlabel pdiffusion 2005 -2030 2005 -2030 0 feedthrough
rlabel pdiffusion 2012 -2030 2012 -2030 0 feedthrough
rlabel pdiffusion 2019 -2030 2019 -2030 0 feedthrough
rlabel pdiffusion 2026 -2030 2026 -2030 0 feedthrough
rlabel pdiffusion 2033 -2030 2033 -2030 0 feedthrough
rlabel pdiffusion 2040 -2030 2040 -2030 0 feedthrough
rlabel pdiffusion 2047 -2030 2047 -2030 0 feedthrough
rlabel pdiffusion 2054 -2030 2054 -2030 0 feedthrough
rlabel pdiffusion 2061 -2030 2061 -2030 0 feedthrough
rlabel pdiffusion 2068 -2030 2068 -2030 0 feedthrough
rlabel pdiffusion 2075 -2030 2075 -2030 0 feedthrough
rlabel pdiffusion 2082 -2030 2082 -2030 0 feedthrough
rlabel pdiffusion 2089 -2030 2089 -2030 0 feedthrough
rlabel pdiffusion 2096 -2030 2096 -2030 0 feedthrough
rlabel pdiffusion 2103 -2030 2103 -2030 0 feedthrough
rlabel pdiffusion 2110 -2030 2110 -2030 0 feedthrough
rlabel pdiffusion 2117 -2030 2117 -2030 0 feedthrough
rlabel pdiffusion 2124 -2030 2124 -2030 0 feedthrough
rlabel pdiffusion 2131 -2030 2131 -2030 0 feedthrough
rlabel pdiffusion 2138 -2030 2138 -2030 0 feedthrough
rlabel pdiffusion 2145 -2030 2145 -2030 0 feedthrough
rlabel pdiffusion 2152 -2030 2152 -2030 0 feedthrough
rlabel pdiffusion 2159 -2030 2159 -2030 0 feedthrough
rlabel pdiffusion 2166 -2030 2166 -2030 0 feedthrough
rlabel pdiffusion 2173 -2030 2173 -2030 0 feedthrough
rlabel pdiffusion 2180 -2030 2180 -2030 0 feedthrough
rlabel pdiffusion 2187 -2030 2187 -2030 0 feedthrough
rlabel pdiffusion 2194 -2030 2194 -2030 0 feedthrough
rlabel pdiffusion 2201 -2030 2201 -2030 0 feedthrough
rlabel pdiffusion 2208 -2030 2208 -2030 0 feedthrough
rlabel pdiffusion 2215 -2030 2215 -2030 0 feedthrough
rlabel pdiffusion 2222 -2030 2222 -2030 0 feedthrough
rlabel pdiffusion 2229 -2030 2229 -2030 0 feedthrough
rlabel pdiffusion 2236 -2030 2236 -2030 0 feedthrough
rlabel pdiffusion 2243 -2030 2243 -2030 0 feedthrough
rlabel pdiffusion 2250 -2030 2250 -2030 0 feedthrough
rlabel pdiffusion 2257 -2030 2257 -2030 0 feedthrough
rlabel pdiffusion 2264 -2030 2264 -2030 0 feedthrough
rlabel pdiffusion 2271 -2030 2271 -2030 0 feedthrough
rlabel pdiffusion 2278 -2030 2278 -2030 0 feedthrough
rlabel pdiffusion 2285 -2030 2285 -2030 0 feedthrough
rlabel pdiffusion 2292 -2030 2292 -2030 0 feedthrough
rlabel pdiffusion 2299 -2030 2299 -2030 0 feedthrough
rlabel pdiffusion 2306 -2030 2306 -2030 0 feedthrough
rlabel pdiffusion 2313 -2030 2313 -2030 0 feedthrough
rlabel pdiffusion 2320 -2030 2320 -2030 0 feedthrough
rlabel pdiffusion 2327 -2030 2327 -2030 0 feedthrough
rlabel pdiffusion 2334 -2030 2334 -2030 0 feedthrough
rlabel pdiffusion 2341 -2030 2341 -2030 0 feedthrough
rlabel pdiffusion 2348 -2030 2348 -2030 0 feedthrough
rlabel pdiffusion 2355 -2030 2355 -2030 0 feedthrough
rlabel pdiffusion 2362 -2030 2362 -2030 0 feedthrough
rlabel pdiffusion 2369 -2030 2369 -2030 0 feedthrough
rlabel pdiffusion 2376 -2030 2376 -2030 0 feedthrough
rlabel pdiffusion 2383 -2030 2383 -2030 0 feedthrough
rlabel pdiffusion 2390 -2030 2390 -2030 0 feedthrough
rlabel pdiffusion 2397 -2030 2397 -2030 0 feedthrough
rlabel pdiffusion 2404 -2030 2404 -2030 0 feedthrough
rlabel pdiffusion 2411 -2030 2411 -2030 0 feedthrough
rlabel pdiffusion 2418 -2030 2418 -2030 0 cellNo=501
rlabel pdiffusion 2425 -2030 2425 -2030 0 feedthrough
rlabel pdiffusion 3 -2181 3 -2181 0 cellNo=1014
rlabel pdiffusion 10 -2181 10 -2181 0 feedthrough
rlabel pdiffusion 17 -2181 17 -2181 0 feedthrough
rlabel pdiffusion 24 -2181 24 -2181 0 feedthrough
rlabel pdiffusion 31 -2181 31 -2181 0 feedthrough
rlabel pdiffusion 38 -2181 38 -2181 0 cellNo=27
rlabel pdiffusion 45 -2181 45 -2181 0 feedthrough
rlabel pdiffusion 52 -2181 52 -2181 0 cellNo=367
rlabel pdiffusion 59 -2181 59 -2181 0 feedthrough
rlabel pdiffusion 66 -2181 66 -2181 0 feedthrough
rlabel pdiffusion 73 -2181 73 -2181 0 feedthrough
rlabel pdiffusion 80 -2181 80 -2181 0 feedthrough
rlabel pdiffusion 87 -2181 87 -2181 0 feedthrough
rlabel pdiffusion 94 -2181 94 -2181 0 cellNo=48
rlabel pdiffusion 101 -2181 101 -2181 0 feedthrough
rlabel pdiffusion 108 -2181 108 -2181 0 feedthrough
rlabel pdiffusion 115 -2181 115 -2181 0 feedthrough
rlabel pdiffusion 122 -2181 122 -2181 0 cellNo=909
rlabel pdiffusion 129 -2181 129 -2181 0 cellNo=61
rlabel pdiffusion 136 -2181 136 -2181 0 cellNo=463
rlabel pdiffusion 143 -2181 143 -2181 0 feedthrough
rlabel pdiffusion 150 -2181 150 -2181 0 feedthrough
rlabel pdiffusion 157 -2181 157 -2181 0 feedthrough
rlabel pdiffusion 164 -2181 164 -2181 0 feedthrough
rlabel pdiffusion 171 -2181 171 -2181 0 feedthrough
rlabel pdiffusion 178 -2181 178 -2181 0 feedthrough
rlabel pdiffusion 185 -2181 185 -2181 0 feedthrough
rlabel pdiffusion 192 -2181 192 -2181 0 feedthrough
rlabel pdiffusion 199 -2181 199 -2181 0 feedthrough
rlabel pdiffusion 206 -2181 206 -2181 0 feedthrough
rlabel pdiffusion 213 -2181 213 -2181 0 feedthrough
rlabel pdiffusion 220 -2181 220 -2181 0 feedthrough
rlabel pdiffusion 227 -2181 227 -2181 0 feedthrough
rlabel pdiffusion 234 -2181 234 -2181 0 cellNo=749
rlabel pdiffusion 241 -2181 241 -2181 0 cellNo=835
rlabel pdiffusion 248 -2181 248 -2181 0 feedthrough
rlabel pdiffusion 255 -2181 255 -2181 0 cellNo=480
rlabel pdiffusion 262 -2181 262 -2181 0 feedthrough
rlabel pdiffusion 269 -2181 269 -2181 0 feedthrough
rlabel pdiffusion 276 -2181 276 -2181 0 feedthrough
rlabel pdiffusion 283 -2181 283 -2181 0 feedthrough
rlabel pdiffusion 290 -2181 290 -2181 0 feedthrough
rlabel pdiffusion 297 -2181 297 -2181 0 feedthrough
rlabel pdiffusion 304 -2181 304 -2181 0 feedthrough
rlabel pdiffusion 311 -2181 311 -2181 0 feedthrough
rlabel pdiffusion 318 -2181 318 -2181 0 feedthrough
rlabel pdiffusion 325 -2181 325 -2181 0 feedthrough
rlabel pdiffusion 332 -2181 332 -2181 0 feedthrough
rlabel pdiffusion 339 -2181 339 -2181 0 feedthrough
rlabel pdiffusion 346 -2181 346 -2181 0 feedthrough
rlabel pdiffusion 353 -2181 353 -2181 0 feedthrough
rlabel pdiffusion 360 -2181 360 -2181 0 feedthrough
rlabel pdiffusion 367 -2181 367 -2181 0 feedthrough
rlabel pdiffusion 374 -2181 374 -2181 0 feedthrough
rlabel pdiffusion 381 -2181 381 -2181 0 feedthrough
rlabel pdiffusion 388 -2181 388 -2181 0 feedthrough
rlabel pdiffusion 395 -2181 395 -2181 0 feedthrough
rlabel pdiffusion 402 -2181 402 -2181 0 cellNo=984
rlabel pdiffusion 409 -2181 409 -2181 0 feedthrough
rlabel pdiffusion 416 -2181 416 -2181 0 feedthrough
rlabel pdiffusion 423 -2181 423 -2181 0 feedthrough
rlabel pdiffusion 430 -2181 430 -2181 0 feedthrough
rlabel pdiffusion 437 -2181 437 -2181 0 feedthrough
rlabel pdiffusion 444 -2181 444 -2181 0 feedthrough
rlabel pdiffusion 451 -2181 451 -2181 0 feedthrough
rlabel pdiffusion 458 -2181 458 -2181 0 feedthrough
rlabel pdiffusion 465 -2181 465 -2181 0 feedthrough
rlabel pdiffusion 472 -2181 472 -2181 0 feedthrough
rlabel pdiffusion 479 -2181 479 -2181 0 feedthrough
rlabel pdiffusion 486 -2181 486 -2181 0 feedthrough
rlabel pdiffusion 493 -2181 493 -2181 0 cellNo=330
rlabel pdiffusion 500 -2181 500 -2181 0 feedthrough
rlabel pdiffusion 507 -2181 507 -2181 0 feedthrough
rlabel pdiffusion 514 -2181 514 -2181 0 cellNo=145
rlabel pdiffusion 521 -2181 521 -2181 0 feedthrough
rlabel pdiffusion 528 -2181 528 -2181 0 feedthrough
rlabel pdiffusion 535 -2181 535 -2181 0 feedthrough
rlabel pdiffusion 542 -2181 542 -2181 0 feedthrough
rlabel pdiffusion 549 -2181 549 -2181 0 feedthrough
rlabel pdiffusion 556 -2181 556 -2181 0 feedthrough
rlabel pdiffusion 563 -2181 563 -2181 0 feedthrough
rlabel pdiffusion 570 -2181 570 -2181 0 feedthrough
rlabel pdiffusion 577 -2181 577 -2181 0 feedthrough
rlabel pdiffusion 584 -2181 584 -2181 0 feedthrough
rlabel pdiffusion 591 -2181 591 -2181 0 feedthrough
rlabel pdiffusion 598 -2181 598 -2181 0 feedthrough
rlabel pdiffusion 605 -2181 605 -2181 0 feedthrough
rlabel pdiffusion 612 -2181 612 -2181 0 feedthrough
rlabel pdiffusion 619 -2181 619 -2181 0 feedthrough
rlabel pdiffusion 626 -2181 626 -2181 0 feedthrough
rlabel pdiffusion 633 -2181 633 -2181 0 feedthrough
rlabel pdiffusion 640 -2181 640 -2181 0 feedthrough
rlabel pdiffusion 647 -2181 647 -2181 0 feedthrough
rlabel pdiffusion 654 -2181 654 -2181 0 cellNo=940
rlabel pdiffusion 661 -2181 661 -2181 0 feedthrough
rlabel pdiffusion 668 -2181 668 -2181 0 cellNo=18
rlabel pdiffusion 675 -2181 675 -2181 0 feedthrough
rlabel pdiffusion 682 -2181 682 -2181 0 feedthrough
rlabel pdiffusion 689 -2181 689 -2181 0 feedthrough
rlabel pdiffusion 696 -2181 696 -2181 0 feedthrough
rlabel pdiffusion 703 -2181 703 -2181 0 feedthrough
rlabel pdiffusion 710 -2181 710 -2181 0 feedthrough
rlabel pdiffusion 717 -2181 717 -2181 0 feedthrough
rlabel pdiffusion 724 -2181 724 -2181 0 feedthrough
rlabel pdiffusion 731 -2181 731 -2181 0 feedthrough
rlabel pdiffusion 738 -2181 738 -2181 0 feedthrough
rlabel pdiffusion 745 -2181 745 -2181 0 cellNo=850
rlabel pdiffusion 752 -2181 752 -2181 0 feedthrough
rlabel pdiffusion 759 -2181 759 -2181 0 cellNo=695
rlabel pdiffusion 766 -2181 766 -2181 0 feedthrough
rlabel pdiffusion 773 -2181 773 -2181 0 feedthrough
rlabel pdiffusion 780 -2181 780 -2181 0 feedthrough
rlabel pdiffusion 787 -2181 787 -2181 0 cellNo=517
rlabel pdiffusion 794 -2181 794 -2181 0 feedthrough
rlabel pdiffusion 801 -2181 801 -2181 0 feedthrough
rlabel pdiffusion 808 -2181 808 -2181 0 feedthrough
rlabel pdiffusion 815 -2181 815 -2181 0 feedthrough
rlabel pdiffusion 822 -2181 822 -2181 0 feedthrough
rlabel pdiffusion 829 -2181 829 -2181 0 feedthrough
rlabel pdiffusion 836 -2181 836 -2181 0 feedthrough
rlabel pdiffusion 843 -2181 843 -2181 0 feedthrough
rlabel pdiffusion 850 -2181 850 -2181 0 feedthrough
rlabel pdiffusion 857 -2181 857 -2181 0 feedthrough
rlabel pdiffusion 864 -2181 864 -2181 0 feedthrough
rlabel pdiffusion 871 -2181 871 -2181 0 feedthrough
rlabel pdiffusion 878 -2181 878 -2181 0 feedthrough
rlabel pdiffusion 885 -2181 885 -2181 0 feedthrough
rlabel pdiffusion 892 -2181 892 -2181 0 feedthrough
rlabel pdiffusion 899 -2181 899 -2181 0 feedthrough
rlabel pdiffusion 906 -2181 906 -2181 0 feedthrough
rlabel pdiffusion 913 -2181 913 -2181 0 feedthrough
rlabel pdiffusion 920 -2181 920 -2181 0 feedthrough
rlabel pdiffusion 927 -2181 927 -2181 0 feedthrough
rlabel pdiffusion 934 -2181 934 -2181 0 feedthrough
rlabel pdiffusion 941 -2181 941 -2181 0 feedthrough
rlabel pdiffusion 948 -2181 948 -2181 0 feedthrough
rlabel pdiffusion 955 -2181 955 -2181 0 feedthrough
rlabel pdiffusion 962 -2181 962 -2181 0 feedthrough
rlabel pdiffusion 969 -2181 969 -2181 0 feedthrough
rlabel pdiffusion 976 -2181 976 -2181 0 cellNo=301
rlabel pdiffusion 983 -2181 983 -2181 0 feedthrough
rlabel pdiffusion 990 -2181 990 -2181 0 feedthrough
rlabel pdiffusion 997 -2181 997 -2181 0 feedthrough
rlabel pdiffusion 1004 -2181 1004 -2181 0 feedthrough
rlabel pdiffusion 1011 -2181 1011 -2181 0 feedthrough
rlabel pdiffusion 1018 -2181 1018 -2181 0 feedthrough
rlabel pdiffusion 1025 -2181 1025 -2181 0 feedthrough
rlabel pdiffusion 1032 -2181 1032 -2181 0 feedthrough
rlabel pdiffusion 1039 -2181 1039 -2181 0 feedthrough
rlabel pdiffusion 1046 -2181 1046 -2181 0 feedthrough
rlabel pdiffusion 1053 -2181 1053 -2181 0 cellNo=423
rlabel pdiffusion 1060 -2181 1060 -2181 0 feedthrough
rlabel pdiffusion 1067 -2181 1067 -2181 0 feedthrough
rlabel pdiffusion 1074 -2181 1074 -2181 0 feedthrough
rlabel pdiffusion 1081 -2181 1081 -2181 0 feedthrough
rlabel pdiffusion 1088 -2181 1088 -2181 0 feedthrough
rlabel pdiffusion 1095 -2181 1095 -2181 0 feedthrough
rlabel pdiffusion 1102 -2181 1102 -2181 0 feedthrough
rlabel pdiffusion 1109 -2181 1109 -2181 0 feedthrough
rlabel pdiffusion 1116 -2181 1116 -2181 0 feedthrough
rlabel pdiffusion 1123 -2181 1123 -2181 0 feedthrough
rlabel pdiffusion 1130 -2181 1130 -2181 0 feedthrough
rlabel pdiffusion 1137 -2181 1137 -2181 0 feedthrough
rlabel pdiffusion 1144 -2181 1144 -2181 0 feedthrough
rlabel pdiffusion 1151 -2181 1151 -2181 0 cellNo=356
rlabel pdiffusion 1158 -2181 1158 -2181 0 feedthrough
rlabel pdiffusion 1165 -2181 1165 -2181 0 feedthrough
rlabel pdiffusion 1172 -2181 1172 -2181 0 feedthrough
rlabel pdiffusion 1179 -2181 1179 -2181 0 feedthrough
rlabel pdiffusion 1186 -2181 1186 -2181 0 cellNo=379
rlabel pdiffusion 1193 -2181 1193 -2181 0 feedthrough
rlabel pdiffusion 1200 -2181 1200 -2181 0 cellNo=140
rlabel pdiffusion 1207 -2181 1207 -2181 0 feedthrough
rlabel pdiffusion 1214 -2181 1214 -2181 0 feedthrough
rlabel pdiffusion 1221 -2181 1221 -2181 0 cellNo=156
rlabel pdiffusion 1228 -2181 1228 -2181 0 cellNo=576
rlabel pdiffusion 1235 -2181 1235 -2181 0 feedthrough
rlabel pdiffusion 1242 -2181 1242 -2181 0 feedthrough
rlabel pdiffusion 1249 -2181 1249 -2181 0 feedthrough
rlabel pdiffusion 1256 -2181 1256 -2181 0 cellNo=182
rlabel pdiffusion 1263 -2181 1263 -2181 0 feedthrough
rlabel pdiffusion 1270 -2181 1270 -2181 0 feedthrough
rlabel pdiffusion 1277 -2181 1277 -2181 0 feedthrough
rlabel pdiffusion 1284 -2181 1284 -2181 0 feedthrough
rlabel pdiffusion 1291 -2181 1291 -2181 0 feedthrough
rlabel pdiffusion 1298 -2181 1298 -2181 0 feedthrough
rlabel pdiffusion 1305 -2181 1305 -2181 0 cellNo=668
rlabel pdiffusion 1312 -2181 1312 -2181 0 feedthrough
rlabel pdiffusion 1319 -2181 1319 -2181 0 feedthrough
rlabel pdiffusion 1326 -2181 1326 -2181 0 feedthrough
rlabel pdiffusion 1333 -2181 1333 -2181 0 cellNo=986
rlabel pdiffusion 1340 -2181 1340 -2181 0 cellNo=314
rlabel pdiffusion 1347 -2181 1347 -2181 0 feedthrough
rlabel pdiffusion 1354 -2181 1354 -2181 0 feedthrough
rlabel pdiffusion 1361 -2181 1361 -2181 0 feedthrough
rlabel pdiffusion 1368 -2181 1368 -2181 0 cellNo=114
rlabel pdiffusion 1375 -2181 1375 -2181 0 feedthrough
rlabel pdiffusion 1382 -2181 1382 -2181 0 cellNo=768
rlabel pdiffusion 1389 -2181 1389 -2181 0 feedthrough
rlabel pdiffusion 1396 -2181 1396 -2181 0 feedthrough
rlabel pdiffusion 1403 -2181 1403 -2181 0 cellNo=324
rlabel pdiffusion 1410 -2181 1410 -2181 0 feedthrough
rlabel pdiffusion 1417 -2181 1417 -2181 0 feedthrough
rlabel pdiffusion 1424 -2181 1424 -2181 0 feedthrough
rlabel pdiffusion 1431 -2181 1431 -2181 0 feedthrough
rlabel pdiffusion 1438 -2181 1438 -2181 0 feedthrough
rlabel pdiffusion 1445 -2181 1445 -2181 0 feedthrough
rlabel pdiffusion 1452 -2181 1452 -2181 0 feedthrough
rlabel pdiffusion 1459 -2181 1459 -2181 0 feedthrough
rlabel pdiffusion 1466 -2181 1466 -2181 0 feedthrough
rlabel pdiffusion 1473 -2181 1473 -2181 0 feedthrough
rlabel pdiffusion 1480 -2181 1480 -2181 0 feedthrough
rlabel pdiffusion 1487 -2181 1487 -2181 0 cellNo=226
rlabel pdiffusion 1494 -2181 1494 -2181 0 feedthrough
rlabel pdiffusion 1501 -2181 1501 -2181 0 feedthrough
rlabel pdiffusion 1508 -2181 1508 -2181 0 feedthrough
rlabel pdiffusion 1515 -2181 1515 -2181 0 feedthrough
rlabel pdiffusion 1522 -2181 1522 -2181 0 feedthrough
rlabel pdiffusion 1529 -2181 1529 -2181 0 feedthrough
rlabel pdiffusion 1536 -2181 1536 -2181 0 feedthrough
rlabel pdiffusion 1543 -2181 1543 -2181 0 feedthrough
rlabel pdiffusion 1550 -2181 1550 -2181 0 feedthrough
rlabel pdiffusion 1557 -2181 1557 -2181 0 feedthrough
rlabel pdiffusion 1564 -2181 1564 -2181 0 feedthrough
rlabel pdiffusion 1571 -2181 1571 -2181 0 feedthrough
rlabel pdiffusion 1578 -2181 1578 -2181 0 cellNo=193
rlabel pdiffusion 1585 -2181 1585 -2181 0 feedthrough
rlabel pdiffusion 1592 -2181 1592 -2181 0 feedthrough
rlabel pdiffusion 1599 -2181 1599 -2181 0 feedthrough
rlabel pdiffusion 1606 -2181 1606 -2181 0 feedthrough
rlabel pdiffusion 1613 -2181 1613 -2181 0 feedthrough
rlabel pdiffusion 1620 -2181 1620 -2181 0 feedthrough
rlabel pdiffusion 1627 -2181 1627 -2181 0 feedthrough
rlabel pdiffusion 1634 -2181 1634 -2181 0 feedthrough
rlabel pdiffusion 1641 -2181 1641 -2181 0 feedthrough
rlabel pdiffusion 1648 -2181 1648 -2181 0 cellNo=98
rlabel pdiffusion 1655 -2181 1655 -2181 0 feedthrough
rlabel pdiffusion 1662 -2181 1662 -2181 0 feedthrough
rlabel pdiffusion 1669 -2181 1669 -2181 0 feedthrough
rlabel pdiffusion 1676 -2181 1676 -2181 0 feedthrough
rlabel pdiffusion 1683 -2181 1683 -2181 0 feedthrough
rlabel pdiffusion 1690 -2181 1690 -2181 0 feedthrough
rlabel pdiffusion 1697 -2181 1697 -2181 0 feedthrough
rlabel pdiffusion 1704 -2181 1704 -2181 0 feedthrough
rlabel pdiffusion 1711 -2181 1711 -2181 0 cellNo=558
rlabel pdiffusion 1718 -2181 1718 -2181 0 feedthrough
rlabel pdiffusion 1725 -2181 1725 -2181 0 feedthrough
rlabel pdiffusion 1732 -2181 1732 -2181 0 feedthrough
rlabel pdiffusion 1739 -2181 1739 -2181 0 feedthrough
rlabel pdiffusion 1746 -2181 1746 -2181 0 feedthrough
rlabel pdiffusion 1753 -2181 1753 -2181 0 feedthrough
rlabel pdiffusion 1760 -2181 1760 -2181 0 feedthrough
rlabel pdiffusion 1767 -2181 1767 -2181 0 feedthrough
rlabel pdiffusion 1774 -2181 1774 -2181 0 feedthrough
rlabel pdiffusion 1781 -2181 1781 -2181 0 feedthrough
rlabel pdiffusion 1788 -2181 1788 -2181 0 feedthrough
rlabel pdiffusion 1795 -2181 1795 -2181 0 feedthrough
rlabel pdiffusion 1802 -2181 1802 -2181 0 feedthrough
rlabel pdiffusion 1809 -2181 1809 -2181 0 feedthrough
rlabel pdiffusion 1816 -2181 1816 -2181 0 feedthrough
rlabel pdiffusion 1823 -2181 1823 -2181 0 feedthrough
rlabel pdiffusion 1830 -2181 1830 -2181 0 feedthrough
rlabel pdiffusion 1837 -2181 1837 -2181 0 cellNo=626
rlabel pdiffusion 1844 -2181 1844 -2181 0 feedthrough
rlabel pdiffusion 1851 -2181 1851 -2181 0 feedthrough
rlabel pdiffusion 1858 -2181 1858 -2181 0 cellNo=242
rlabel pdiffusion 1865 -2181 1865 -2181 0 feedthrough
rlabel pdiffusion 1872 -2181 1872 -2181 0 feedthrough
rlabel pdiffusion 1879 -2181 1879 -2181 0 feedthrough
rlabel pdiffusion 1886 -2181 1886 -2181 0 feedthrough
rlabel pdiffusion 1893 -2181 1893 -2181 0 feedthrough
rlabel pdiffusion 1900 -2181 1900 -2181 0 feedthrough
rlabel pdiffusion 1907 -2181 1907 -2181 0 feedthrough
rlabel pdiffusion 1914 -2181 1914 -2181 0 feedthrough
rlabel pdiffusion 1921 -2181 1921 -2181 0 feedthrough
rlabel pdiffusion 1928 -2181 1928 -2181 0 feedthrough
rlabel pdiffusion 1935 -2181 1935 -2181 0 feedthrough
rlabel pdiffusion 1942 -2181 1942 -2181 0 feedthrough
rlabel pdiffusion 1949 -2181 1949 -2181 0 feedthrough
rlabel pdiffusion 1956 -2181 1956 -2181 0 cellNo=62
rlabel pdiffusion 1963 -2181 1963 -2181 0 feedthrough
rlabel pdiffusion 1970 -2181 1970 -2181 0 feedthrough
rlabel pdiffusion 1977 -2181 1977 -2181 0 feedthrough
rlabel pdiffusion 1984 -2181 1984 -2181 0 feedthrough
rlabel pdiffusion 1991 -2181 1991 -2181 0 feedthrough
rlabel pdiffusion 1998 -2181 1998 -2181 0 feedthrough
rlabel pdiffusion 2005 -2181 2005 -2181 0 feedthrough
rlabel pdiffusion 2012 -2181 2012 -2181 0 feedthrough
rlabel pdiffusion 2019 -2181 2019 -2181 0 feedthrough
rlabel pdiffusion 2026 -2181 2026 -2181 0 feedthrough
rlabel pdiffusion 2033 -2181 2033 -2181 0 feedthrough
rlabel pdiffusion 2040 -2181 2040 -2181 0 feedthrough
rlabel pdiffusion 2047 -2181 2047 -2181 0 feedthrough
rlabel pdiffusion 2054 -2181 2054 -2181 0 feedthrough
rlabel pdiffusion 2061 -2181 2061 -2181 0 feedthrough
rlabel pdiffusion 2068 -2181 2068 -2181 0 feedthrough
rlabel pdiffusion 2075 -2181 2075 -2181 0 feedthrough
rlabel pdiffusion 2082 -2181 2082 -2181 0 feedthrough
rlabel pdiffusion 2089 -2181 2089 -2181 0 feedthrough
rlabel pdiffusion 2096 -2181 2096 -2181 0 feedthrough
rlabel pdiffusion 2103 -2181 2103 -2181 0 feedthrough
rlabel pdiffusion 2110 -2181 2110 -2181 0 feedthrough
rlabel pdiffusion 2117 -2181 2117 -2181 0 feedthrough
rlabel pdiffusion 2124 -2181 2124 -2181 0 feedthrough
rlabel pdiffusion 2131 -2181 2131 -2181 0 feedthrough
rlabel pdiffusion 2138 -2181 2138 -2181 0 feedthrough
rlabel pdiffusion 2145 -2181 2145 -2181 0 feedthrough
rlabel pdiffusion 2152 -2181 2152 -2181 0 feedthrough
rlabel pdiffusion 2159 -2181 2159 -2181 0 feedthrough
rlabel pdiffusion 2166 -2181 2166 -2181 0 feedthrough
rlabel pdiffusion 2173 -2181 2173 -2181 0 feedthrough
rlabel pdiffusion 2180 -2181 2180 -2181 0 feedthrough
rlabel pdiffusion 2187 -2181 2187 -2181 0 feedthrough
rlabel pdiffusion 2194 -2181 2194 -2181 0 feedthrough
rlabel pdiffusion 2201 -2181 2201 -2181 0 feedthrough
rlabel pdiffusion 2208 -2181 2208 -2181 0 feedthrough
rlabel pdiffusion 2215 -2181 2215 -2181 0 feedthrough
rlabel pdiffusion 2222 -2181 2222 -2181 0 feedthrough
rlabel pdiffusion 2229 -2181 2229 -2181 0 feedthrough
rlabel pdiffusion 2236 -2181 2236 -2181 0 feedthrough
rlabel pdiffusion 2243 -2181 2243 -2181 0 feedthrough
rlabel pdiffusion 2250 -2181 2250 -2181 0 feedthrough
rlabel pdiffusion 2257 -2181 2257 -2181 0 feedthrough
rlabel pdiffusion 2264 -2181 2264 -2181 0 feedthrough
rlabel pdiffusion 2271 -2181 2271 -2181 0 feedthrough
rlabel pdiffusion 2278 -2181 2278 -2181 0 feedthrough
rlabel pdiffusion 2285 -2181 2285 -2181 0 feedthrough
rlabel pdiffusion 2292 -2181 2292 -2181 0 feedthrough
rlabel pdiffusion 2299 -2181 2299 -2181 0 feedthrough
rlabel pdiffusion 2306 -2181 2306 -2181 0 feedthrough
rlabel pdiffusion 2313 -2181 2313 -2181 0 feedthrough
rlabel pdiffusion 2320 -2181 2320 -2181 0 feedthrough
rlabel pdiffusion 2327 -2181 2327 -2181 0 feedthrough
rlabel pdiffusion 2334 -2181 2334 -2181 0 feedthrough
rlabel pdiffusion 2341 -2181 2341 -2181 0 feedthrough
rlabel pdiffusion 2348 -2181 2348 -2181 0 feedthrough
rlabel pdiffusion 2355 -2181 2355 -2181 0 feedthrough
rlabel pdiffusion 2362 -2181 2362 -2181 0 feedthrough
rlabel pdiffusion 2369 -2181 2369 -2181 0 feedthrough
rlabel pdiffusion 2376 -2181 2376 -2181 0 feedthrough
rlabel pdiffusion 2383 -2181 2383 -2181 0 feedthrough
rlabel pdiffusion 2390 -2181 2390 -2181 0 feedthrough
rlabel pdiffusion 2397 -2181 2397 -2181 0 feedthrough
rlabel pdiffusion 2404 -2181 2404 -2181 0 feedthrough
rlabel pdiffusion 2411 -2181 2411 -2181 0 feedthrough
rlabel pdiffusion 2418 -2181 2418 -2181 0 feedthrough
rlabel pdiffusion 2425 -2181 2425 -2181 0 feedthrough
rlabel pdiffusion 3 -2330 3 -2330 0 feedthrough
rlabel pdiffusion 10 -2330 10 -2330 0 cellNo=1003
rlabel pdiffusion 17 -2330 17 -2330 0 feedthrough
rlabel pdiffusion 24 -2330 24 -2330 0 feedthrough
rlabel pdiffusion 31 -2330 31 -2330 0 cellNo=639
rlabel pdiffusion 38 -2330 38 -2330 0 feedthrough
rlabel pdiffusion 45 -2330 45 -2330 0 feedthrough
rlabel pdiffusion 52 -2330 52 -2330 0 feedthrough
rlabel pdiffusion 59 -2330 59 -2330 0 feedthrough
rlabel pdiffusion 66 -2330 66 -2330 0 feedthrough
rlabel pdiffusion 73 -2330 73 -2330 0 feedthrough
rlabel pdiffusion 80 -2330 80 -2330 0 feedthrough
rlabel pdiffusion 87 -2330 87 -2330 0 feedthrough
rlabel pdiffusion 94 -2330 94 -2330 0 cellNo=348
rlabel pdiffusion 101 -2330 101 -2330 0 feedthrough
rlabel pdiffusion 108 -2330 108 -2330 0 feedthrough
rlabel pdiffusion 115 -2330 115 -2330 0 feedthrough
rlabel pdiffusion 122 -2330 122 -2330 0 feedthrough
rlabel pdiffusion 129 -2330 129 -2330 0 feedthrough
rlabel pdiffusion 136 -2330 136 -2330 0 feedthrough
rlabel pdiffusion 143 -2330 143 -2330 0 cellNo=466
rlabel pdiffusion 150 -2330 150 -2330 0 feedthrough
rlabel pdiffusion 157 -2330 157 -2330 0 feedthrough
rlabel pdiffusion 164 -2330 164 -2330 0 cellNo=653
rlabel pdiffusion 171 -2330 171 -2330 0 feedthrough
rlabel pdiffusion 178 -2330 178 -2330 0 feedthrough
rlabel pdiffusion 185 -2330 185 -2330 0 feedthrough
rlabel pdiffusion 192 -2330 192 -2330 0 feedthrough
rlabel pdiffusion 199 -2330 199 -2330 0 feedthrough
rlabel pdiffusion 206 -2330 206 -2330 0 feedthrough
rlabel pdiffusion 213 -2330 213 -2330 0 feedthrough
rlabel pdiffusion 220 -2330 220 -2330 0 feedthrough
rlabel pdiffusion 227 -2330 227 -2330 0 feedthrough
rlabel pdiffusion 234 -2330 234 -2330 0 feedthrough
rlabel pdiffusion 241 -2330 241 -2330 0 cellNo=223
rlabel pdiffusion 248 -2330 248 -2330 0 cellNo=306
rlabel pdiffusion 255 -2330 255 -2330 0 feedthrough
rlabel pdiffusion 262 -2330 262 -2330 0 feedthrough
rlabel pdiffusion 269 -2330 269 -2330 0 feedthrough
rlabel pdiffusion 276 -2330 276 -2330 0 feedthrough
rlabel pdiffusion 283 -2330 283 -2330 0 feedthrough
rlabel pdiffusion 290 -2330 290 -2330 0 feedthrough
rlabel pdiffusion 297 -2330 297 -2330 0 feedthrough
rlabel pdiffusion 304 -2330 304 -2330 0 feedthrough
rlabel pdiffusion 311 -2330 311 -2330 0 feedthrough
rlabel pdiffusion 318 -2330 318 -2330 0 feedthrough
rlabel pdiffusion 325 -2330 325 -2330 0 feedthrough
rlabel pdiffusion 332 -2330 332 -2330 0 feedthrough
rlabel pdiffusion 339 -2330 339 -2330 0 feedthrough
rlabel pdiffusion 346 -2330 346 -2330 0 feedthrough
rlabel pdiffusion 353 -2330 353 -2330 0 feedthrough
rlabel pdiffusion 360 -2330 360 -2330 0 feedthrough
rlabel pdiffusion 367 -2330 367 -2330 0 feedthrough
rlabel pdiffusion 374 -2330 374 -2330 0 feedthrough
rlabel pdiffusion 381 -2330 381 -2330 0 feedthrough
rlabel pdiffusion 388 -2330 388 -2330 0 feedthrough
rlabel pdiffusion 395 -2330 395 -2330 0 feedthrough
rlabel pdiffusion 402 -2330 402 -2330 0 feedthrough
rlabel pdiffusion 409 -2330 409 -2330 0 feedthrough
rlabel pdiffusion 416 -2330 416 -2330 0 feedthrough
rlabel pdiffusion 423 -2330 423 -2330 0 feedthrough
rlabel pdiffusion 430 -2330 430 -2330 0 cellNo=848
rlabel pdiffusion 437 -2330 437 -2330 0 feedthrough
rlabel pdiffusion 444 -2330 444 -2330 0 feedthrough
rlabel pdiffusion 451 -2330 451 -2330 0 feedthrough
rlabel pdiffusion 458 -2330 458 -2330 0 feedthrough
rlabel pdiffusion 465 -2330 465 -2330 0 feedthrough
rlabel pdiffusion 472 -2330 472 -2330 0 feedthrough
rlabel pdiffusion 479 -2330 479 -2330 0 feedthrough
rlabel pdiffusion 486 -2330 486 -2330 0 feedthrough
rlabel pdiffusion 493 -2330 493 -2330 0 feedthrough
rlabel pdiffusion 500 -2330 500 -2330 0 feedthrough
rlabel pdiffusion 507 -2330 507 -2330 0 feedthrough
rlabel pdiffusion 514 -2330 514 -2330 0 feedthrough
rlabel pdiffusion 521 -2330 521 -2330 0 feedthrough
rlabel pdiffusion 528 -2330 528 -2330 0 feedthrough
rlabel pdiffusion 535 -2330 535 -2330 0 feedthrough
rlabel pdiffusion 542 -2330 542 -2330 0 feedthrough
rlabel pdiffusion 549 -2330 549 -2330 0 feedthrough
rlabel pdiffusion 556 -2330 556 -2330 0 feedthrough
rlabel pdiffusion 563 -2330 563 -2330 0 feedthrough
rlabel pdiffusion 570 -2330 570 -2330 0 feedthrough
rlabel pdiffusion 577 -2330 577 -2330 0 feedthrough
rlabel pdiffusion 584 -2330 584 -2330 0 feedthrough
rlabel pdiffusion 591 -2330 591 -2330 0 cellNo=2
rlabel pdiffusion 598 -2330 598 -2330 0 feedthrough
rlabel pdiffusion 605 -2330 605 -2330 0 feedthrough
rlabel pdiffusion 612 -2330 612 -2330 0 feedthrough
rlabel pdiffusion 619 -2330 619 -2330 0 cellNo=213
rlabel pdiffusion 626 -2330 626 -2330 0 cellNo=761
rlabel pdiffusion 633 -2330 633 -2330 0 feedthrough
rlabel pdiffusion 640 -2330 640 -2330 0 feedthrough
rlabel pdiffusion 647 -2330 647 -2330 0 feedthrough
rlabel pdiffusion 654 -2330 654 -2330 0 feedthrough
rlabel pdiffusion 661 -2330 661 -2330 0 cellNo=549
rlabel pdiffusion 668 -2330 668 -2330 0 cellNo=510
rlabel pdiffusion 675 -2330 675 -2330 0 feedthrough
rlabel pdiffusion 682 -2330 682 -2330 0 feedthrough
rlabel pdiffusion 689 -2330 689 -2330 0 feedthrough
rlabel pdiffusion 696 -2330 696 -2330 0 feedthrough
rlabel pdiffusion 703 -2330 703 -2330 0 cellNo=410
rlabel pdiffusion 710 -2330 710 -2330 0 feedthrough
rlabel pdiffusion 717 -2330 717 -2330 0 feedthrough
rlabel pdiffusion 724 -2330 724 -2330 0 cellNo=444
rlabel pdiffusion 731 -2330 731 -2330 0 feedthrough
rlabel pdiffusion 738 -2330 738 -2330 0 feedthrough
rlabel pdiffusion 745 -2330 745 -2330 0 feedthrough
rlabel pdiffusion 752 -2330 752 -2330 0 feedthrough
rlabel pdiffusion 759 -2330 759 -2330 0 feedthrough
rlabel pdiffusion 766 -2330 766 -2330 0 cellNo=333
rlabel pdiffusion 773 -2330 773 -2330 0 feedthrough
rlabel pdiffusion 780 -2330 780 -2330 0 cellNo=418
rlabel pdiffusion 787 -2330 787 -2330 0 feedthrough
rlabel pdiffusion 794 -2330 794 -2330 0 feedthrough
rlabel pdiffusion 801 -2330 801 -2330 0 feedthrough
rlabel pdiffusion 808 -2330 808 -2330 0 feedthrough
rlabel pdiffusion 815 -2330 815 -2330 0 feedthrough
rlabel pdiffusion 822 -2330 822 -2330 0 feedthrough
rlabel pdiffusion 829 -2330 829 -2330 0 feedthrough
rlabel pdiffusion 836 -2330 836 -2330 0 feedthrough
rlabel pdiffusion 843 -2330 843 -2330 0 feedthrough
rlabel pdiffusion 850 -2330 850 -2330 0 feedthrough
rlabel pdiffusion 857 -2330 857 -2330 0 cellNo=773
rlabel pdiffusion 864 -2330 864 -2330 0 feedthrough
rlabel pdiffusion 871 -2330 871 -2330 0 feedthrough
rlabel pdiffusion 878 -2330 878 -2330 0 feedthrough
rlabel pdiffusion 885 -2330 885 -2330 0 feedthrough
rlabel pdiffusion 892 -2330 892 -2330 0 feedthrough
rlabel pdiffusion 899 -2330 899 -2330 0 feedthrough
rlabel pdiffusion 906 -2330 906 -2330 0 feedthrough
rlabel pdiffusion 913 -2330 913 -2330 0 feedthrough
rlabel pdiffusion 920 -2330 920 -2330 0 cellNo=683
rlabel pdiffusion 927 -2330 927 -2330 0 feedthrough
rlabel pdiffusion 934 -2330 934 -2330 0 cellNo=59
rlabel pdiffusion 941 -2330 941 -2330 0 feedthrough
rlabel pdiffusion 948 -2330 948 -2330 0 feedthrough
rlabel pdiffusion 955 -2330 955 -2330 0 feedthrough
rlabel pdiffusion 962 -2330 962 -2330 0 feedthrough
rlabel pdiffusion 969 -2330 969 -2330 0 feedthrough
rlabel pdiffusion 976 -2330 976 -2330 0 cellNo=790
rlabel pdiffusion 983 -2330 983 -2330 0 feedthrough
rlabel pdiffusion 990 -2330 990 -2330 0 cellNo=243
rlabel pdiffusion 997 -2330 997 -2330 0 feedthrough
rlabel pdiffusion 1004 -2330 1004 -2330 0 feedthrough
rlabel pdiffusion 1011 -2330 1011 -2330 0 feedthrough
rlabel pdiffusion 1018 -2330 1018 -2330 0 feedthrough
rlabel pdiffusion 1025 -2330 1025 -2330 0 feedthrough
rlabel pdiffusion 1032 -2330 1032 -2330 0 feedthrough
rlabel pdiffusion 1039 -2330 1039 -2330 0 cellNo=672
rlabel pdiffusion 1046 -2330 1046 -2330 0 feedthrough
rlabel pdiffusion 1053 -2330 1053 -2330 0 feedthrough
rlabel pdiffusion 1060 -2330 1060 -2330 0 feedthrough
rlabel pdiffusion 1067 -2330 1067 -2330 0 feedthrough
rlabel pdiffusion 1074 -2330 1074 -2330 0 feedthrough
rlabel pdiffusion 1081 -2330 1081 -2330 0 feedthrough
rlabel pdiffusion 1088 -2330 1088 -2330 0 feedthrough
rlabel pdiffusion 1095 -2330 1095 -2330 0 feedthrough
rlabel pdiffusion 1102 -2330 1102 -2330 0 feedthrough
rlabel pdiffusion 1109 -2330 1109 -2330 0 feedthrough
rlabel pdiffusion 1116 -2330 1116 -2330 0 feedthrough
rlabel pdiffusion 1123 -2330 1123 -2330 0 feedthrough
rlabel pdiffusion 1130 -2330 1130 -2330 0 feedthrough
rlabel pdiffusion 1137 -2330 1137 -2330 0 cellNo=962
rlabel pdiffusion 1144 -2330 1144 -2330 0 feedthrough
rlabel pdiffusion 1151 -2330 1151 -2330 0 feedthrough
rlabel pdiffusion 1158 -2330 1158 -2330 0 feedthrough
rlabel pdiffusion 1165 -2330 1165 -2330 0 feedthrough
rlabel pdiffusion 1172 -2330 1172 -2330 0 feedthrough
rlabel pdiffusion 1179 -2330 1179 -2330 0 feedthrough
rlabel pdiffusion 1186 -2330 1186 -2330 0 feedthrough
rlabel pdiffusion 1193 -2330 1193 -2330 0 feedthrough
rlabel pdiffusion 1200 -2330 1200 -2330 0 feedthrough
rlabel pdiffusion 1207 -2330 1207 -2330 0 feedthrough
rlabel pdiffusion 1214 -2330 1214 -2330 0 feedthrough
rlabel pdiffusion 1221 -2330 1221 -2330 0 feedthrough
rlabel pdiffusion 1228 -2330 1228 -2330 0 feedthrough
rlabel pdiffusion 1235 -2330 1235 -2330 0 feedthrough
rlabel pdiffusion 1242 -2330 1242 -2330 0 feedthrough
rlabel pdiffusion 1249 -2330 1249 -2330 0 cellNo=647
rlabel pdiffusion 1256 -2330 1256 -2330 0 feedthrough
rlabel pdiffusion 1263 -2330 1263 -2330 0 feedthrough
rlabel pdiffusion 1270 -2330 1270 -2330 0 feedthrough
rlabel pdiffusion 1277 -2330 1277 -2330 0 feedthrough
rlabel pdiffusion 1284 -2330 1284 -2330 0 feedthrough
rlabel pdiffusion 1291 -2330 1291 -2330 0 cellNo=803
rlabel pdiffusion 1298 -2330 1298 -2330 0 feedthrough
rlabel pdiffusion 1305 -2330 1305 -2330 0 feedthrough
rlabel pdiffusion 1312 -2330 1312 -2330 0 feedthrough
rlabel pdiffusion 1319 -2330 1319 -2330 0 cellNo=457
rlabel pdiffusion 1326 -2330 1326 -2330 0 feedthrough
rlabel pdiffusion 1333 -2330 1333 -2330 0 feedthrough
rlabel pdiffusion 1340 -2330 1340 -2330 0 feedthrough
rlabel pdiffusion 1347 -2330 1347 -2330 0 feedthrough
rlabel pdiffusion 1354 -2330 1354 -2330 0 feedthrough
rlabel pdiffusion 1361 -2330 1361 -2330 0 feedthrough
rlabel pdiffusion 1368 -2330 1368 -2330 0 feedthrough
rlabel pdiffusion 1375 -2330 1375 -2330 0 feedthrough
rlabel pdiffusion 1382 -2330 1382 -2330 0 feedthrough
rlabel pdiffusion 1389 -2330 1389 -2330 0 feedthrough
rlabel pdiffusion 1396 -2330 1396 -2330 0 cellNo=212
rlabel pdiffusion 1403 -2330 1403 -2330 0 feedthrough
rlabel pdiffusion 1410 -2330 1410 -2330 0 feedthrough
rlabel pdiffusion 1417 -2330 1417 -2330 0 feedthrough
rlabel pdiffusion 1424 -2330 1424 -2330 0 feedthrough
rlabel pdiffusion 1431 -2330 1431 -2330 0 feedthrough
rlabel pdiffusion 1438 -2330 1438 -2330 0 feedthrough
rlabel pdiffusion 1445 -2330 1445 -2330 0 feedthrough
rlabel pdiffusion 1452 -2330 1452 -2330 0 feedthrough
rlabel pdiffusion 1459 -2330 1459 -2330 0 feedthrough
rlabel pdiffusion 1466 -2330 1466 -2330 0 feedthrough
rlabel pdiffusion 1473 -2330 1473 -2330 0 feedthrough
rlabel pdiffusion 1480 -2330 1480 -2330 0 feedthrough
rlabel pdiffusion 1487 -2330 1487 -2330 0 feedthrough
rlabel pdiffusion 1494 -2330 1494 -2330 0 cellNo=328
rlabel pdiffusion 1501 -2330 1501 -2330 0 cellNo=249
rlabel pdiffusion 1508 -2330 1508 -2330 0 feedthrough
rlabel pdiffusion 1515 -2330 1515 -2330 0 cellNo=855
rlabel pdiffusion 1522 -2330 1522 -2330 0 feedthrough
rlabel pdiffusion 1529 -2330 1529 -2330 0 feedthrough
rlabel pdiffusion 1536 -2330 1536 -2330 0 feedthrough
rlabel pdiffusion 1543 -2330 1543 -2330 0 cellNo=913
rlabel pdiffusion 1550 -2330 1550 -2330 0 feedthrough
rlabel pdiffusion 1557 -2330 1557 -2330 0 feedthrough
rlabel pdiffusion 1564 -2330 1564 -2330 0 feedthrough
rlabel pdiffusion 1571 -2330 1571 -2330 0 feedthrough
rlabel pdiffusion 1578 -2330 1578 -2330 0 feedthrough
rlabel pdiffusion 1585 -2330 1585 -2330 0 feedthrough
rlabel pdiffusion 1592 -2330 1592 -2330 0 feedthrough
rlabel pdiffusion 1599 -2330 1599 -2330 0 feedthrough
rlabel pdiffusion 1606 -2330 1606 -2330 0 feedthrough
rlabel pdiffusion 1613 -2330 1613 -2330 0 feedthrough
rlabel pdiffusion 1620 -2330 1620 -2330 0 feedthrough
rlabel pdiffusion 1627 -2330 1627 -2330 0 cellNo=907
rlabel pdiffusion 1634 -2330 1634 -2330 0 feedthrough
rlabel pdiffusion 1641 -2330 1641 -2330 0 feedthrough
rlabel pdiffusion 1648 -2330 1648 -2330 0 feedthrough
rlabel pdiffusion 1655 -2330 1655 -2330 0 feedthrough
rlabel pdiffusion 1662 -2330 1662 -2330 0 feedthrough
rlabel pdiffusion 1669 -2330 1669 -2330 0 feedthrough
rlabel pdiffusion 1676 -2330 1676 -2330 0 feedthrough
rlabel pdiffusion 1683 -2330 1683 -2330 0 cellNo=489
rlabel pdiffusion 1690 -2330 1690 -2330 0 feedthrough
rlabel pdiffusion 1697 -2330 1697 -2330 0 feedthrough
rlabel pdiffusion 1704 -2330 1704 -2330 0 feedthrough
rlabel pdiffusion 1711 -2330 1711 -2330 0 feedthrough
rlabel pdiffusion 1718 -2330 1718 -2330 0 feedthrough
rlabel pdiffusion 1725 -2330 1725 -2330 0 feedthrough
rlabel pdiffusion 1732 -2330 1732 -2330 0 feedthrough
rlabel pdiffusion 1739 -2330 1739 -2330 0 feedthrough
rlabel pdiffusion 1746 -2330 1746 -2330 0 feedthrough
rlabel pdiffusion 1753 -2330 1753 -2330 0 feedthrough
rlabel pdiffusion 1760 -2330 1760 -2330 0 feedthrough
rlabel pdiffusion 1767 -2330 1767 -2330 0 feedthrough
rlabel pdiffusion 1774 -2330 1774 -2330 0 feedthrough
rlabel pdiffusion 1781 -2330 1781 -2330 0 feedthrough
rlabel pdiffusion 1788 -2330 1788 -2330 0 feedthrough
rlabel pdiffusion 1795 -2330 1795 -2330 0 feedthrough
rlabel pdiffusion 1802 -2330 1802 -2330 0 feedthrough
rlabel pdiffusion 1809 -2330 1809 -2330 0 feedthrough
rlabel pdiffusion 1816 -2330 1816 -2330 0 feedthrough
rlabel pdiffusion 1823 -2330 1823 -2330 0 feedthrough
rlabel pdiffusion 1830 -2330 1830 -2330 0 feedthrough
rlabel pdiffusion 1837 -2330 1837 -2330 0 feedthrough
rlabel pdiffusion 1844 -2330 1844 -2330 0 feedthrough
rlabel pdiffusion 1851 -2330 1851 -2330 0 feedthrough
rlabel pdiffusion 1858 -2330 1858 -2330 0 feedthrough
rlabel pdiffusion 1865 -2330 1865 -2330 0 feedthrough
rlabel pdiffusion 1872 -2330 1872 -2330 0 feedthrough
rlabel pdiffusion 1879 -2330 1879 -2330 0 feedthrough
rlabel pdiffusion 1886 -2330 1886 -2330 0 feedthrough
rlabel pdiffusion 1893 -2330 1893 -2330 0 cellNo=465
rlabel pdiffusion 1900 -2330 1900 -2330 0 feedthrough
rlabel pdiffusion 1907 -2330 1907 -2330 0 feedthrough
rlabel pdiffusion 1914 -2330 1914 -2330 0 feedthrough
rlabel pdiffusion 1921 -2330 1921 -2330 0 feedthrough
rlabel pdiffusion 1928 -2330 1928 -2330 0 feedthrough
rlabel pdiffusion 1935 -2330 1935 -2330 0 cellNo=945
rlabel pdiffusion 1942 -2330 1942 -2330 0 feedthrough
rlabel pdiffusion 1949 -2330 1949 -2330 0 feedthrough
rlabel pdiffusion 1956 -2330 1956 -2330 0 feedthrough
rlabel pdiffusion 1963 -2330 1963 -2330 0 feedthrough
rlabel pdiffusion 1970 -2330 1970 -2330 0 feedthrough
rlabel pdiffusion 1977 -2330 1977 -2330 0 cellNo=56
rlabel pdiffusion 1984 -2330 1984 -2330 0 feedthrough
rlabel pdiffusion 1991 -2330 1991 -2330 0 feedthrough
rlabel pdiffusion 1998 -2330 1998 -2330 0 feedthrough
rlabel pdiffusion 2005 -2330 2005 -2330 0 feedthrough
rlabel pdiffusion 2012 -2330 2012 -2330 0 feedthrough
rlabel pdiffusion 2019 -2330 2019 -2330 0 feedthrough
rlabel pdiffusion 2026 -2330 2026 -2330 0 feedthrough
rlabel pdiffusion 2033 -2330 2033 -2330 0 feedthrough
rlabel pdiffusion 2040 -2330 2040 -2330 0 feedthrough
rlabel pdiffusion 2047 -2330 2047 -2330 0 feedthrough
rlabel pdiffusion 2054 -2330 2054 -2330 0 feedthrough
rlabel pdiffusion 2061 -2330 2061 -2330 0 feedthrough
rlabel pdiffusion 2068 -2330 2068 -2330 0 feedthrough
rlabel pdiffusion 2075 -2330 2075 -2330 0 feedthrough
rlabel pdiffusion 2082 -2330 2082 -2330 0 feedthrough
rlabel pdiffusion 2089 -2330 2089 -2330 0 feedthrough
rlabel pdiffusion 2096 -2330 2096 -2330 0 feedthrough
rlabel pdiffusion 2103 -2330 2103 -2330 0 feedthrough
rlabel pdiffusion 2110 -2330 2110 -2330 0 feedthrough
rlabel pdiffusion 2117 -2330 2117 -2330 0 feedthrough
rlabel pdiffusion 2124 -2330 2124 -2330 0 feedthrough
rlabel pdiffusion 2131 -2330 2131 -2330 0 feedthrough
rlabel pdiffusion 2138 -2330 2138 -2330 0 feedthrough
rlabel pdiffusion 2145 -2330 2145 -2330 0 feedthrough
rlabel pdiffusion 2152 -2330 2152 -2330 0 feedthrough
rlabel pdiffusion 2159 -2330 2159 -2330 0 feedthrough
rlabel pdiffusion 2166 -2330 2166 -2330 0 feedthrough
rlabel pdiffusion 2173 -2330 2173 -2330 0 feedthrough
rlabel pdiffusion 2180 -2330 2180 -2330 0 feedthrough
rlabel pdiffusion 2187 -2330 2187 -2330 0 feedthrough
rlabel pdiffusion 2194 -2330 2194 -2330 0 feedthrough
rlabel pdiffusion 2201 -2330 2201 -2330 0 feedthrough
rlabel pdiffusion 2208 -2330 2208 -2330 0 feedthrough
rlabel pdiffusion 2215 -2330 2215 -2330 0 feedthrough
rlabel pdiffusion 2222 -2330 2222 -2330 0 feedthrough
rlabel pdiffusion 2229 -2330 2229 -2330 0 feedthrough
rlabel pdiffusion 2236 -2330 2236 -2330 0 feedthrough
rlabel pdiffusion 2243 -2330 2243 -2330 0 feedthrough
rlabel pdiffusion 2250 -2330 2250 -2330 0 feedthrough
rlabel pdiffusion 2257 -2330 2257 -2330 0 feedthrough
rlabel pdiffusion 2264 -2330 2264 -2330 0 feedthrough
rlabel pdiffusion 2271 -2330 2271 -2330 0 feedthrough
rlabel pdiffusion 2278 -2330 2278 -2330 0 feedthrough
rlabel pdiffusion 2285 -2330 2285 -2330 0 feedthrough
rlabel pdiffusion 2292 -2330 2292 -2330 0 feedthrough
rlabel pdiffusion 2299 -2330 2299 -2330 0 feedthrough
rlabel pdiffusion 2306 -2330 2306 -2330 0 feedthrough
rlabel pdiffusion 2313 -2330 2313 -2330 0 feedthrough
rlabel pdiffusion 2320 -2330 2320 -2330 0 feedthrough
rlabel pdiffusion 2327 -2330 2327 -2330 0 feedthrough
rlabel pdiffusion 2334 -2330 2334 -2330 0 cellNo=99
rlabel pdiffusion 2341 -2330 2341 -2330 0 cellNo=960
rlabel pdiffusion 2348 -2330 2348 -2330 0 feedthrough
rlabel pdiffusion 3 -2503 3 -2503 0 cellNo=619
rlabel pdiffusion 10 -2503 10 -2503 0 cellNo=900
rlabel pdiffusion 17 -2503 17 -2503 0 cellNo=859
rlabel pdiffusion 24 -2503 24 -2503 0 feedthrough
rlabel pdiffusion 31 -2503 31 -2503 0 cellNo=751
rlabel pdiffusion 38 -2503 38 -2503 0 cellNo=862
rlabel pdiffusion 45 -2503 45 -2503 0 feedthrough
rlabel pdiffusion 52 -2503 52 -2503 0 feedthrough
rlabel pdiffusion 59 -2503 59 -2503 0 cellNo=978
rlabel pdiffusion 66 -2503 66 -2503 0 feedthrough
rlabel pdiffusion 73 -2503 73 -2503 0 feedthrough
rlabel pdiffusion 80 -2503 80 -2503 0 feedthrough
rlabel pdiffusion 87 -2503 87 -2503 0 feedthrough
rlabel pdiffusion 94 -2503 94 -2503 0 cellNo=397
rlabel pdiffusion 101 -2503 101 -2503 0 feedthrough
rlabel pdiffusion 108 -2503 108 -2503 0 cellNo=430
rlabel pdiffusion 115 -2503 115 -2503 0 feedthrough
rlabel pdiffusion 122 -2503 122 -2503 0 feedthrough
rlabel pdiffusion 129 -2503 129 -2503 0 feedthrough
rlabel pdiffusion 136 -2503 136 -2503 0 feedthrough
rlabel pdiffusion 143 -2503 143 -2503 0 feedthrough
rlabel pdiffusion 150 -2503 150 -2503 0 feedthrough
rlabel pdiffusion 157 -2503 157 -2503 0 feedthrough
rlabel pdiffusion 164 -2503 164 -2503 0 cellNo=438
rlabel pdiffusion 171 -2503 171 -2503 0 feedthrough
rlabel pdiffusion 178 -2503 178 -2503 0 feedthrough
rlabel pdiffusion 185 -2503 185 -2503 0 feedthrough
rlabel pdiffusion 192 -2503 192 -2503 0 feedthrough
rlabel pdiffusion 199 -2503 199 -2503 0 feedthrough
rlabel pdiffusion 206 -2503 206 -2503 0 feedthrough
rlabel pdiffusion 213 -2503 213 -2503 0 feedthrough
rlabel pdiffusion 220 -2503 220 -2503 0 feedthrough
rlabel pdiffusion 227 -2503 227 -2503 0 feedthrough
rlabel pdiffusion 234 -2503 234 -2503 0 feedthrough
rlabel pdiffusion 241 -2503 241 -2503 0 feedthrough
rlabel pdiffusion 248 -2503 248 -2503 0 feedthrough
rlabel pdiffusion 255 -2503 255 -2503 0 feedthrough
rlabel pdiffusion 262 -2503 262 -2503 0 feedthrough
rlabel pdiffusion 269 -2503 269 -2503 0 feedthrough
rlabel pdiffusion 276 -2503 276 -2503 0 feedthrough
rlabel pdiffusion 283 -2503 283 -2503 0 feedthrough
rlabel pdiffusion 290 -2503 290 -2503 0 feedthrough
rlabel pdiffusion 297 -2503 297 -2503 0 feedthrough
rlabel pdiffusion 304 -2503 304 -2503 0 feedthrough
rlabel pdiffusion 311 -2503 311 -2503 0 feedthrough
rlabel pdiffusion 318 -2503 318 -2503 0 feedthrough
rlabel pdiffusion 325 -2503 325 -2503 0 feedthrough
rlabel pdiffusion 332 -2503 332 -2503 0 feedthrough
rlabel pdiffusion 339 -2503 339 -2503 0 feedthrough
rlabel pdiffusion 346 -2503 346 -2503 0 feedthrough
rlabel pdiffusion 353 -2503 353 -2503 0 feedthrough
rlabel pdiffusion 360 -2503 360 -2503 0 feedthrough
rlabel pdiffusion 367 -2503 367 -2503 0 feedthrough
rlabel pdiffusion 374 -2503 374 -2503 0 feedthrough
rlabel pdiffusion 381 -2503 381 -2503 0 feedthrough
rlabel pdiffusion 388 -2503 388 -2503 0 feedthrough
rlabel pdiffusion 395 -2503 395 -2503 0 feedthrough
rlabel pdiffusion 402 -2503 402 -2503 0 feedthrough
rlabel pdiffusion 409 -2503 409 -2503 0 feedthrough
rlabel pdiffusion 416 -2503 416 -2503 0 feedthrough
rlabel pdiffusion 423 -2503 423 -2503 0 feedthrough
rlabel pdiffusion 430 -2503 430 -2503 0 feedthrough
rlabel pdiffusion 437 -2503 437 -2503 0 feedthrough
rlabel pdiffusion 444 -2503 444 -2503 0 feedthrough
rlabel pdiffusion 451 -2503 451 -2503 0 feedthrough
rlabel pdiffusion 458 -2503 458 -2503 0 feedthrough
rlabel pdiffusion 465 -2503 465 -2503 0 feedthrough
rlabel pdiffusion 472 -2503 472 -2503 0 feedthrough
rlabel pdiffusion 479 -2503 479 -2503 0 cellNo=849
rlabel pdiffusion 486 -2503 486 -2503 0 feedthrough
rlabel pdiffusion 493 -2503 493 -2503 0 feedthrough
rlabel pdiffusion 500 -2503 500 -2503 0 feedthrough
rlabel pdiffusion 507 -2503 507 -2503 0 feedthrough
rlabel pdiffusion 514 -2503 514 -2503 0 feedthrough
rlabel pdiffusion 521 -2503 521 -2503 0 feedthrough
rlabel pdiffusion 528 -2503 528 -2503 0 feedthrough
rlabel pdiffusion 535 -2503 535 -2503 0 feedthrough
rlabel pdiffusion 542 -2503 542 -2503 0 feedthrough
rlabel pdiffusion 549 -2503 549 -2503 0 feedthrough
rlabel pdiffusion 556 -2503 556 -2503 0 feedthrough
rlabel pdiffusion 563 -2503 563 -2503 0 feedthrough
rlabel pdiffusion 570 -2503 570 -2503 0 feedthrough
rlabel pdiffusion 577 -2503 577 -2503 0 feedthrough
rlabel pdiffusion 584 -2503 584 -2503 0 feedthrough
rlabel pdiffusion 591 -2503 591 -2503 0 feedthrough
rlabel pdiffusion 598 -2503 598 -2503 0 feedthrough
rlabel pdiffusion 605 -2503 605 -2503 0 cellNo=133
rlabel pdiffusion 612 -2503 612 -2503 0 feedthrough
rlabel pdiffusion 619 -2503 619 -2503 0 feedthrough
rlabel pdiffusion 626 -2503 626 -2503 0 feedthrough
rlabel pdiffusion 633 -2503 633 -2503 0 feedthrough
rlabel pdiffusion 640 -2503 640 -2503 0 feedthrough
rlabel pdiffusion 647 -2503 647 -2503 0 feedthrough
rlabel pdiffusion 654 -2503 654 -2503 0 feedthrough
rlabel pdiffusion 661 -2503 661 -2503 0 feedthrough
rlabel pdiffusion 668 -2503 668 -2503 0 cellNo=16
rlabel pdiffusion 675 -2503 675 -2503 0 feedthrough
rlabel pdiffusion 682 -2503 682 -2503 0 feedthrough
rlabel pdiffusion 689 -2503 689 -2503 0 feedthrough
rlabel pdiffusion 696 -2503 696 -2503 0 feedthrough
rlabel pdiffusion 703 -2503 703 -2503 0 feedthrough
rlabel pdiffusion 710 -2503 710 -2503 0 feedthrough
rlabel pdiffusion 717 -2503 717 -2503 0 feedthrough
rlabel pdiffusion 724 -2503 724 -2503 0 feedthrough
rlabel pdiffusion 731 -2503 731 -2503 0 feedthrough
rlabel pdiffusion 738 -2503 738 -2503 0 cellNo=1000
rlabel pdiffusion 745 -2503 745 -2503 0 feedthrough
rlabel pdiffusion 752 -2503 752 -2503 0 feedthrough
rlabel pdiffusion 759 -2503 759 -2503 0 feedthrough
rlabel pdiffusion 766 -2503 766 -2503 0 feedthrough
rlabel pdiffusion 773 -2503 773 -2503 0 cellNo=625
rlabel pdiffusion 780 -2503 780 -2503 0 feedthrough
rlabel pdiffusion 787 -2503 787 -2503 0 feedthrough
rlabel pdiffusion 794 -2503 794 -2503 0 cellNo=886
rlabel pdiffusion 801 -2503 801 -2503 0 feedthrough
rlabel pdiffusion 808 -2503 808 -2503 0 feedthrough
rlabel pdiffusion 815 -2503 815 -2503 0 feedthrough
rlabel pdiffusion 822 -2503 822 -2503 0 feedthrough
rlabel pdiffusion 829 -2503 829 -2503 0 feedthrough
rlabel pdiffusion 836 -2503 836 -2503 0 feedthrough
rlabel pdiffusion 843 -2503 843 -2503 0 feedthrough
rlabel pdiffusion 850 -2503 850 -2503 0 feedthrough
rlabel pdiffusion 857 -2503 857 -2503 0 cellNo=825
rlabel pdiffusion 864 -2503 864 -2503 0 feedthrough
rlabel pdiffusion 871 -2503 871 -2503 0 cellNo=736
rlabel pdiffusion 878 -2503 878 -2503 0 feedthrough
rlabel pdiffusion 885 -2503 885 -2503 0 feedthrough
rlabel pdiffusion 892 -2503 892 -2503 0 feedthrough
rlabel pdiffusion 899 -2503 899 -2503 0 feedthrough
rlabel pdiffusion 906 -2503 906 -2503 0 feedthrough
rlabel pdiffusion 913 -2503 913 -2503 0 feedthrough
rlabel pdiffusion 920 -2503 920 -2503 0 cellNo=33
rlabel pdiffusion 927 -2503 927 -2503 0 feedthrough
rlabel pdiffusion 934 -2503 934 -2503 0 feedthrough
rlabel pdiffusion 941 -2503 941 -2503 0 feedthrough
rlabel pdiffusion 948 -2503 948 -2503 0 feedthrough
rlabel pdiffusion 955 -2503 955 -2503 0 cellNo=583
rlabel pdiffusion 962 -2503 962 -2503 0 feedthrough
rlabel pdiffusion 969 -2503 969 -2503 0 feedthrough
rlabel pdiffusion 976 -2503 976 -2503 0 cellNo=815
rlabel pdiffusion 983 -2503 983 -2503 0 feedthrough
rlabel pdiffusion 990 -2503 990 -2503 0 cellNo=624
rlabel pdiffusion 997 -2503 997 -2503 0 feedthrough
rlabel pdiffusion 1004 -2503 1004 -2503 0 feedthrough
rlabel pdiffusion 1011 -2503 1011 -2503 0 cellNo=972
rlabel pdiffusion 1018 -2503 1018 -2503 0 cellNo=380
rlabel pdiffusion 1025 -2503 1025 -2503 0 feedthrough
rlabel pdiffusion 1032 -2503 1032 -2503 0 feedthrough
rlabel pdiffusion 1039 -2503 1039 -2503 0 feedthrough
rlabel pdiffusion 1046 -2503 1046 -2503 0 feedthrough
rlabel pdiffusion 1053 -2503 1053 -2503 0 cellNo=500
rlabel pdiffusion 1060 -2503 1060 -2503 0 feedthrough
rlabel pdiffusion 1067 -2503 1067 -2503 0 feedthrough
rlabel pdiffusion 1074 -2503 1074 -2503 0 cellNo=936
rlabel pdiffusion 1081 -2503 1081 -2503 0 cellNo=428
rlabel pdiffusion 1088 -2503 1088 -2503 0 feedthrough
rlabel pdiffusion 1095 -2503 1095 -2503 0 feedthrough
rlabel pdiffusion 1102 -2503 1102 -2503 0 feedthrough
rlabel pdiffusion 1109 -2503 1109 -2503 0 feedthrough
rlabel pdiffusion 1116 -2503 1116 -2503 0 feedthrough
rlabel pdiffusion 1123 -2503 1123 -2503 0 feedthrough
rlabel pdiffusion 1130 -2503 1130 -2503 0 feedthrough
rlabel pdiffusion 1137 -2503 1137 -2503 0 feedthrough
rlabel pdiffusion 1144 -2503 1144 -2503 0 feedthrough
rlabel pdiffusion 1151 -2503 1151 -2503 0 feedthrough
rlabel pdiffusion 1158 -2503 1158 -2503 0 feedthrough
rlabel pdiffusion 1165 -2503 1165 -2503 0 feedthrough
rlabel pdiffusion 1172 -2503 1172 -2503 0 cellNo=47
rlabel pdiffusion 1179 -2503 1179 -2503 0 feedthrough
rlabel pdiffusion 1186 -2503 1186 -2503 0 feedthrough
rlabel pdiffusion 1193 -2503 1193 -2503 0 feedthrough
rlabel pdiffusion 1200 -2503 1200 -2503 0 feedthrough
rlabel pdiffusion 1207 -2503 1207 -2503 0 feedthrough
rlabel pdiffusion 1214 -2503 1214 -2503 0 cellNo=88
rlabel pdiffusion 1221 -2503 1221 -2503 0 feedthrough
rlabel pdiffusion 1228 -2503 1228 -2503 0 feedthrough
rlabel pdiffusion 1235 -2503 1235 -2503 0 feedthrough
rlabel pdiffusion 1242 -2503 1242 -2503 0 feedthrough
rlabel pdiffusion 1249 -2503 1249 -2503 0 feedthrough
rlabel pdiffusion 1256 -2503 1256 -2503 0 feedthrough
rlabel pdiffusion 1263 -2503 1263 -2503 0 feedthrough
rlabel pdiffusion 1270 -2503 1270 -2503 0 cellNo=198
rlabel pdiffusion 1277 -2503 1277 -2503 0 feedthrough
rlabel pdiffusion 1284 -2503 1284 -2503 0 feedthrough
rlabel pdiffusion 1291 -2503 1291 -2503 0 cellNo=970
rlabel pdiffusion 1298 -2503 1298 -2503 0 feedthrough
rlabel pdiffusion 1305 -2503 1305 -2503 0 feedthrough
rlabel pdiffusion 1312 -2503 1312 -2503 0 feedthrough
rlabel pdiffusion 1319 -2503 1319 -2503 0 feedthrough
rlabel pdiffusion 1326 -2503 1326 -2503 0 feedthrough
rlabel pdiffusion 1333 -2503 1333 -2503 0 cellNo=734
rlabel pdiffusion 1340 -2503 1340 -2503 0 feedthrough
rlabel pdiffusion 1347 -2503 1347 -2503 0 feedthrough
rlabel pdiffusion 1354 -2503 1354 -2503 0 cellNo=481
rlabel pdiffusion 1361 -2503 1361 -2503 0 cellNo=605
rlabel pdiffusion 1368 -2503 1368 -2503 0 feedthrough
rlabel pdiffusion 1375 -2503 1375 -2503 0 cellNo=192
rlabel pdiffusion 1382 -2503 1382 -2503 0 feedthrough
rlabel pdiffusion 1389 -2503 1389 -2503 0 feedthrough
rlabel pdiffusion 1396 -2503 1396 -2503 0 feedthrough
rlabel pdiffusion 1403 -2503 1403 -2503 0 feedthrough
rlabel pdiffusion 1410 -2503 1410 -2503 0 feedthrough
rlabel pdiffusion 1417 -2503 1417 -2503 0 feedthrough
rlabel pdiffusion 1424 -2503 1424 -2503 0 feedthrough
rlabel pdiffusion 1431 -2503 1431 -2503 0 feedthrough
rlabel pdiffusion 1438 -2503 1438 -2503 0 feedthrough
rlabel pdiffusion 1445 -2503 1445 -2503 0 feedthrough
rlabel pdiffusion 1452 -2503 1452 -2503 0 feedthrough
rlabel pdiffusion 1459 -2503 1459 -2503 0 feedthrough
rlabel pdiffusion 1466 -2503 1466 -2503 0 feedthrough
rlabel pdiffusion 1473 -2503 1473 -2503 0 feedthrough
rlabel pdiffusion 1480 -2503 1480 -2503 0 feedthrough
rlabel pdiffusion 1487 -2503 1487 -2503 0 feedthrough
rlabel pdiffusion 1494 -2503 1494 -2503 0 feedthrough
rlabel pdiffusion 1501 -2503 1501 -2503 0 feedthrough
rlabel pdiffusion 1508 -2503 1508 -2503 0 feedthrough
rlabel pdiffusion 1515 -2503 1515 -2503 0 feedthrough
rlabel pdiffusion 1522 -2503 1522 -2503 0 feedthrough
rlabel pdiffusion 1529 -2503 1529 -2503 0 feedthrough
rlabel pdiffusion 1536 -2503 1536 -2503 0 feedthrough
rlabel pdiffusion 1543 -2503 1543 -2503 0 feedthrough
rlabel pdiffusion 1550 -2503 1550 -2503 0 feedthrough
rlabel pdiffusion 1557 -2503 1557 -2503 0 feedthrough
rlabel pdiffusion 1564 -2503 1564 -2503 0 feedthrough
rlabel pdiffusion 1571 -2503 1571 -2503 0 feedthrough
rlabel pdiffusion 1578 -2503 1578 -2503 0 cellNo=923
rlabel pdiffusion 1585 -2503 1585 -2503 0 feedthrough
rlabel pdiffusion 1592 -2503 1592 -2503 0 feedthrough
rlabel pdiffusion 1599 -2503 1599 -2503 0 cellNo=881
rlabel pdiffusion 1606 -2503 1606 -2503 0 feedthrough
rlabel pdiffusion 1613 -2503 1613 -2503 0 feedthrough
rlabel pdiffusion 1620 -2503 1620 -2503 0 feedthrough
rlabel pdiffusion 1627 -2503 1627 -2503 0 feedthrough
rlabel pdiffusion 1634 -2503 1634 -2503 0 feedthrough
rlabel pdiffusion 1641 -2503 1641 -2503 0 feedthrough
rlabel pdiffusion 1648 -2503 1648 -2503 0 feedthrough
rlabel pdiffusion 1655 -2503 1655 -2503 0 feedthrough
rlabel pdiffusion 1662 -2503 1662 -2503 0 feedthrough
rlabel pdiffusion 1669 -2503 1669 -2503 0 feedthrough
rlabel pdiffusion 1676 -2503 1676 -2503 0 cellNo=341
rlabel pdiffusion 1683 -2503 1683 -2503 0 feedthrough
rlabel pdiffusion 1690 -2503 1690 -2503 0 feedthrough
rlabel pdiffusion 1697 -2503 1697 -2503 0 feedthrough
rlabel pdiffusion 1704 -2503 1704 -2503 0 feedthrough
rlabel pdiffusion 1711 -2503 1711 -2503 0 feedthrough
rlabel pdiffusion 1718 -2503 1718 -2503 0 feedthrough
rlabel pdiffusion 1725 -2503 1725 -2503 0 feedthrough
rlabel pdiffusion 1732 -2503 1732 -2503 0 feedthrough
rlabel pdiffusion 1739 -2503 1739 -2503 0 feedthrough
rlabel pdiffusion 1746 -2503 1746 -2503 0 feedthrough
rlabel pdiffusion 1753 -2503 1753 -2503 0 feedthrough
rlabel pdiffusion 1760 -2503 1760 -2503 0 feedthrough
rlabel pdiffusion 1767 -2503 1767 -2503 0 feedthrough
rlabel pdiffusion 1774 -2503 1774 -2503 0 feedthrough
rlabel pdiffusion 1781 -2503 1781 -2503 0 feedthrough
rlabel pdiffusion 1788 -2503 1788 -2503 0 feedthrough
rlabel pdiffusion 1795 -2503 1795 -2503 0 feedthrough
rlabel pdiffusion 1802 -2503 1802 -2503 0 cellNo=399
rlabel pdiffusion 1809 -2503 1809 -2503 0 feedthrough
rlabel pdiffusion 1816 -2503 1816 -2503 0 feedthrough
rlabel pdiffusion 1823 -2503 1823 -2503 0 feedthrough
rlabel pdiffusion 1830 -2503 1830 -2503 0 feedthrough
rlabel pdiffusion 1837 -2503 1837 -2503 0 feedthrough
rlabel pdiffusion 1844 -2503 1844 -2503 0 feedthrough
rlabel pdiffusion 1851 -2503 1851 -2503 0 feedthrough
rlabel pdiffusion 1858 -2503 1858 -2503 0 feedthrough
rlabel pdiffusion 1865 -2503 1865 -2503 0 feedthrough
rlabel pdiffusion 1872 -2503 1872 -2503 0 feedthrough
rlabel pdiffusion 1879 -2503 1879 -2503 0 feedthrough
rlabel pdiffusion 1886 -2503 1886 -2503 0 feedthrough
rlabel pdiffusion 1893 -2503 1893 -2503 0 feedthrough
rlabel pdiffusion 1900 -2503 1900 -2503 0 feedthrough
rlabel pdiffusion 1907 -2503 1907 -2503 0 feedthrough
rlabel pdiffusion 1914 -2503 1914 -2503 0 feedthrough
rlabel pdiffusion 1921 -2503 1921 -2503 0 feedthrough
rlabel pdiffusion 1928 -2503 1928 -2503 0 feedthrough
rlabel pdiffusion 1935 -2503 1935 -2503 0 feedthrough
rlabel pdiffusion 1942 -2503 1942 -2503 0 feedthrough
rlabel pdiffusion 1949 -2503 1949 -2503 0 feedthrough
rlabel pdiffusion 1956 -2503 1956 -2503 0 feedthrough
rlabel pdiffusion 1963 -2503 1963 -2503 0 feedthrough
rlabel pdiffusion 1970 -2503 1970 -2503 0 feedthrough
rlabel pdiffusion 1977 -2503 1977 -2503 0 feedthrough
rlabel pdiffusion 1984 -2503 1984 -2503 0 feedthrough
rlabel pdiffusion 1991 -2503 1991 -2503 0 feedthrough
rlabel pdiffusion 1998 -2503 1998 -2503 0 feedthrough
rlabel pdiffusion 2005 -2503 2005 -2503 0 feedthrough
rlabel pdiffusion 2012 -2503 2012 -2503 0 feedthrough
rlabel pdiffusion 2019 -2503 2019 -2503 0 feedthrough
rlabel pdiffusion 2026 -2503 2026 -2503 0 feedthrough
rlabel pdiffusion 2033 -2503 2033 -2503 0 feedthrough
rlabel pdiffusion 2040 -2503 2040 -2503 0 feedthrough
rlabel pdiffusion 2047 -2503 2047 -2503 0 feedthrough
rlabel pdiffusion 2054 -2503 2054 -2503 0 feedthrough
rlabel pdiffusion 2061 -2503 2061 -2503 0 feedthrough
rlabel pdiffusion 2068 -2503 2068 -2503 0 feedthrough
rlabel pdiffusion 2075 -2503 2075 -2503 0 feedthrough
rlabel pdiffusion 2082 -2503 2082 -2503 0 feedthrough
rlabel pdiffusion 2089 -2503 2089 -2503 0 feedthrough
rlabel pdiffusion 2096 -2503 2096 -2503 0 feedthrough
rlabel pdiffusion 2103 -2503 2103 -2503 0 feedthrough
rlabel pdiffusion 2110 -2503 2110 -2503 0 feedthrough
rlabel pdiffusion 2117 -2503 2117 -2503 0 feedthrough
rlabel pdiffusion 2124 -2503 2124 -2503 0 feedthrough
rlabel pdiffusion 2131 -2503 2131 -2503 0 feedthrough
rlabel pdiffusion 2138 -2503 2138 -2503 0 feedthrough
rlabel pdiffusion 2145 -2503 2145 -2503 0 feedthrough
rlabel pdiffusion 2152 -2503 2152 -2503 0 feedthrough
rlabel pdiffusion 2159 -2503 2159 -2503 0 feedthrough
rlabel pdiffusion 2166 -2503 2166 -2503 0 feedthrough
rlabel pdiffusion 2173 -2503 2173 -2503 0 feedthrough
rlabel pdiffusion 2180 -2503 2180 -2503 0 feedthrough
rlabel pdiffusion 2187 -2503 2187 -2503 0 feedthrough
rlabel pdiffusion 2194 -2503 2194 -2503 0 feedthrough
rlabel pdiffusion 2201 -2503 2201 -2503 0 feedthrough
rlabel pdiffusion 2208 -2503 2208 -2503 0 feedthrough
rlabel pdiffusion 2215 -2503 2215 -2503 0 feedthrough
rlabel pdiffusion 2222 -2503 2222 -2503 0 feedthrough
rlabel pdiffusion 2229 -2503 2229 -2503 0 feedthrough
rlabel pdiffusion 2236 -2503 2236 -2503 0 feedthrough
rlabel pdiffusion 2243 -2503 2243 -2503 0 feedthrough
rlabel pdiffusion 2250 -2503 2250 -2503 0 feedthrough
rlabel pdiffusion 2257 -2503 2257 -2503 0 feedthrough
rlabel pdiffusion 2264 -2503 2264 -2503 0 feedthrough
rlabel pdiffusion 2271 -2503 2271 -2503 0 feedthrough
rlabel pdiffusion 2278 -2503 2278 -2503 0 cellNo=340
rlabel pdiffusion 2285 -2503 2285 -2503 0 feedthrough
rlabel pdiffusion 2292 -2503 2292 -2503 0 feedthrough
rlabel pdiffusion 2299 -2503 2299 -2503 0 feedthrough
rlabel pdiffusion 2306 -2503 2306 -2503 0 feedthrough
rlabel pdiffusion 2313 -2503 2313 -2503 0 feedthrough
rlabel pdiffusion 3 -2676 3 -2676 0 cellNo=1072
rlabel pdiffusion 10 -2676 10 -2676 0 feedthrough
rlabel pdiffusion 17 -2676 17 -2676 0 feedthrough
rlabel pdiffusion 24 -2676 24 -2676 0 cellNo=476
rlabel pdiffusion 31 -2676 31 -2676 0 feedthrough
rlabel pdiffusion 38 -2676 38 -2676 0 feedthrough
rlabel pdiffusion 45 -2676 45 -2676 0 feedthrough
rlabel pdiffusion 52 -2676 52 -2676 0 cellNo=535
rlabel pdiffusion 59 -2676 59 -2676 0 feedthrough
rlabel pdiffusion 66 -2676 66 -2676 0 cellNo=321
rlabel pdiffusion 73 -2676 73 -2676 0 cellNo=69
rlabel pdiffusion 80 -2676 80 -2676 0 feedthrough
rlabel pdiffusion 87 -2676 87 -2676 0 feedthrough
rlabel pdiffusion 94 -2676 94 -2676 0 feedthrough
rlabel pdiffusion 101 -2676 101 -2676 0 cellNo=343
rlabel pdiffusion 108 -2676 108 -2676 0 feedthrough
rlabel pdiffusion 115 -2676 115 -2676 0 feedthrough
rlabel pdiffusion 122 -2676 122 -2676 0 feedthrough
rlabel pdiffusion 129 -2676 129 -2676 0 cellNo=358
rlabel pdiffusion 136 -2676 136 -2676 0 feedthrough
rlabel pdiffusion 143 -2676 143 -2676 0 feedthrough
rlabel pdiffusion 150 -2676 150 -2676 0 feedthrough
rlabel pdiffusion 157 -2676 157 -2676 0 feedthrough
rlabel pdiffusion 164 -2676 164 -2676 0 feedthrough
rlabel pdiffusion 171 -2676 171 -2676 0 feedthrough
rlabel pdiffusion 178 -2676 178 -2676 0 feedthrough
rlabel pdiffusion 185 -2676 185 -2676 0 feedthrough
rlabel pdiffusion 192 -2676 192 -2676 0 feedthrough
rlabel pdiffusion 199 -2676 199 -2676 0 cellNo=173
rlabel pdiffusion 206 -2676 206 -2676 0 feedthrough
rlabel pdiffusion 213 -2676 213 -2676 0 feedthrough
rlabel pdiffusion 220 -2676 220 -2676 0 feedthrough
rlabel pdiffusion 227 -2676 227 -2676 0 feedthrough
rlabel pdiffusion 234 -2676 234 -2676 0 feedthrough
rlabel pdiffusion 241 -2676 241 -2676 0 cellNo=873
rlabel pdiffusion 248 -2676 248 -2676 0 feedthrough
rlabel pdiffusion 255 -2676 255 -2676 0 feedthrough
rlabel pdiffusion 262 -2676 262 -2676 0 feedthrough
rlabel pdiffusion 269 -2676 269 -2676 0 feedthrough
rlabel pdiffusion 276 -2676 276 -2676 0 feedthrough
rlabel pdiffusion 283 -2676 283 -2676 0 feedthrough
rlabel pdiffusion 290 -2676 290 -2676 0 feedthrough
rlabel pdiffusion 297 -2676 297 -2676 0 feedthrough
rlabel pdiffusion 304 -2676 304 -2676 0 feedthrough
rlabel pdiffusion 311 -2676 311 -2676 0 feedthrough
rlabel pdiffusion 318 -2676 318 -2676 0 feedthrough
rlabel pdiffusion 325 -2676 325 -2676 0 feedthrough
rlabel pdiffusion 332 -2676 332 -2676 0 feedthrough
rlabel pdiffusion 339 -2676 339 -2676 0 feedthrough
rlabel pdiffusion 346 -2676 346 -2676 0 feedthrough
rlabel pdiffusion 353 -2676 353 -2676 0 feedthrough
rlabel pdiffusion 360 -2676 360 -2676 0 feedthrough
rlabel pdiffusion 367 -2676 367 -2676 0 feedthrough
rlabel pdiffusion 374 -2676 374 -2676 0 feedthrough
rlabel pdiffusion 381 -2676 381 -2676 0 feedthrough
rlabel pdiffusion 388 -2676 388 -2676 0 feedthrough
rlabel pdiffusion 395 -2676 395 -2676 0 feedthrough
rlabel pdiffusion 402 -2676 402 -2676 0 feedthrough
rlabel pdiffusion 409 -2676 409 -2676 0 cellNo=350
rlabel pdiffusion 416 -2676 416 -2676 0 feedthrough
rlabel pdiffusion 423 -2676 423 -2676 0 feedthrough
rlabel pdiffusion 430 -2676 430 -2676 0 feedthrough
rlabel pdiffusion 437 -2676 437 -2676 0 feedthrough
rlabel pdiffusion 444 -2676 444 -2676 0 feedthrough
rlabel pdiffusion 451 -2676 451 -2676 0 feedthrough
rlabel pdiffusion 458 -2676 458 -2676 0 feedthrough
rlabel pdiffusion 465 -2676 465 -2676 0 feedthrough
rlabel pdiffusion 472 -2676 472 -2676 0 feedthrough
rlabel pdiffusion 479 -2676 479 -2676 0 feedthrough
rlabel pdiffusion 486 -2676 486 -2676 0 feedthrough
rlabel pdiffusion 493 -2676 493 -2676 0 feedthrough
rlabel pdiffusion 500 -2676 500 -2676 0 feedthrough
rlabel pdiffusion 507 -2676 507 -2676 0 feedthrough
rlabel pdiffusion 514 -2676 514 -2676 0 feedthrough
rlabel pdiffusion 521 -2676 521 -2676 0 feedthrough
rlabel pdiffusion 528 -2676 528 -2676 0 feedthrough
rlabel pdiffusion 535 -2676 535 -2676 0 feedthrough
rlabel pdiffusion 542 -2676 542 -2676 0 feedthrough
rlabel pdiffusion 549 -2676 549 -2676 0 feedthrough
rlabel pdiffusion 556 -2676 556 -2676 0 cellNo=814
rlabel pdiffusion 563 -2676 563 -2676 0 feedthrough
rlabel pdiffusion 570 -2676 570 -2676 0 feedthrough
rlabel pdiffusion 577 -2676 577 -2676 0 feedthrough
rlabel pdiffusion 584 -2676 584 -2676 0 feedthrough
rlabel pdiffusion 591 -2676 591 -2676 0 feedthrough
rlabel pdiffusion 598 -2676 598 -2676 0 feedthrough
rlabel pdiffusion 605 -2676 605 -2676 0 feedthrough
rlabel pdiffusion 612 -2676 612 -2676 0 feedthrough
rlabel pdiffusion 619 -2676 619 -2676 0 feedthrough
rlabel pdiffusion 626 -2676 626 -2676 0 feedthrough
rlabel pdiffusion 633 -2676 633 -2676 0 feedthrough
rlabel pdiffusion 640 -2676 640 -2676 0 feedthrough
rlabel pdiffusion 647 -2676 647 -2676 0 feedthrough
rlabel pdiffusion 654 -2676 654 -2676 0 feedthrough
rlabel pdiffusion 661 -2676 661 -2676 0 feedthrough
rlabel pdiffusion 668 -2676 668 -2676 0 feedthrough
rlabel pdiffusion 675 -2676 675 -2676 0 feedthrough
rlabel pdiffusion 682 -2676 682 -2676 0 feedthrough
rlabel pdiffusion 689 -2676 689 -2676 0 feedthrough
rlabel pdiffusion 696 -2676 696 -2676 0 feedthrough
rlabel pdiffusion 703 -2676 703 -2676 0 feedthrough
rlabel pdiffusion 710 -2676 710 -2676 0 feedthrough
rlabel pdiffusion 717 -2676 717 -2676 0 feedthrough
rlabel pdiffusion 724 -2676 724 -2676 0 cellNo=548
rlabel pdiffusion 731 -2676 731 -2676 0 feedthrough
rlabel pdiffusion 738 -2676 738 -2676 0 feedthrough
rlabel pdiffusion 745 -2676 745 -2676 0 feedthrough
rlabel pdiffusion 752 -2676 752 -2676 0 feedthrough
rlabel pdiffusion 759 -2676 759 -2676 0 feedthrough
rlabel pdiffusion 766 -2676 766 -2676 0 feedthrough
rlabel pdiffusion 773 -2676 773 -2676 0 feedthrough
rlabel pdiffusion 780 -2676 780 -2676 0 feedthrough
rlabel pdiffusion 787 -2676 787 -2676 0 cellNo=729
rlabel pdiffusion 794 -2676 794 -2676 0 feedthrough
rlabel pdiffusion 801 -2676 801 -2676 0 feedthrough
rlabel pdiffusion 808 -2676 808 -2676 0 cellNo=519
rlabel pdiffusion 815 -2676 815 -2676 0 cellNo=899
rlabel pdiffusion 822 -2676 822 -2676 0 cellNo=207
rlabel pdiffusion 829 -2676 829 -2676 0 feedthrough
rlabel pdiffusion 836 -2676 836 -2676 0 feedthrough
rlabel pdiffusion 843 -2676 843 -2676 0 feedthrough
rlabel pdiffusion 850 -2676 850 -2676 0 feedthrough
rlabel pdiffusion 857 -2676 857 -2676 0 feedthrough
rlabel pdiffusion 864 -2676 864 -2676 0 feedthrough
rlabel pdiffusion 871 -2676 871 -2676 0 feedthrough
rlabel pdiffusion 878 -2676 878 -2676 0 feedthrough
rlabel pdiffusion 885 -2676 885 -2676 0 feedthrough
rlabel pdiffusion 892 -2676 892 -2676 0 cellNo=288
rlabel pdiffusion 899 -2676 899 -2676 0 feedthrough
rlabel pdiffusion 906 -2676 906 -2676 0 feedthrough
rlabel pdiffusion 913 -2676 913 -2676 0 feedthrough
rlabel pdiffusion 920 -2676 920 -2676 0 cellNo=650
rlabel pdiffusion 927 -2676 927 -2676 0 feedthrough
rlabel pdiffusion 934 -2676 934 -2676 0 feedthrough
rlabel pdiffusion 941 -2676 941 -2676 0 feedthrough
rlabel pdiffusion 948 -2676 948 -2676 0 cellNo=322
rlabel pdiffusion 955 -2676 955 -2676 0 cellNo=134
rlabel pdiffusion 962 -2676 962 -2676 0 feedthrough
rlabel pdiffusion 969 -2676 969 -2676 0 feedthrough
rlabel pdiffusion 976 -2676 976 -2676 0 feedthrough
rlabel pdiffusion 983 -2676 983 -2676 0 feedthrough
rlabel pdiffusion 990 -2676 990 -2676 0 feedthrough
rlabel pdiffusion 997 -2676 997 -2676 0 feedthrough
rlabel pdiffusion 1004 -2676 1004 -2676 0 cellNo=804
rlabel pdiffusion 1011 -2676 1011 -2676 0 cellNo=364
rlabel pdiffusion 1018 -2676 1018 -2676 0 feedthrough
rlabel pdiffusion 1025 -2676 1025 -2676 0 feedthrough
rlabel pdiffusion 1032 -2676 1032 -2676 0 feedthrough
rlabel pdiffusion 1039 -2676 1039 -2676 0 cellNo=473
rlabel pdiffusion 1046 -2676 1046 -2676 0 feedthrough
rlabel pdiffusion 1053 -2676 1053 -2676 0 feedthrough
rlabel pdiffusion 1060 -2676 1060 -2676 0 feedthrough
rlabel pdiffusion 1067 -2676 1067 -2676 0 feedthrough
rlabel pdiffusion 1074 -2676 1074 -2676 0 feedthrough
rlabel pdiffusion 1081 -2676 1081 -2676 0 feedthrough
rlabel pdiffusion 1088 -2676 1088 -2676 0 feedthrough
rlabel pdiffusion 1095 -2676 1095 -2676 0 feedthrough
rlabel pdiffusion 1102 -2676 1102 -2676 0 feedthrough
rlabel pdiffusion 1109 -2676 1109 -2676 0 feedthrough
rlabel pdiffusion 1116 -2676 1116 -2676 0 feedthrough
rlabel pdiffusion 1123 -2676 1123 -2676 0 cellNo=240
rlabel pdiffusion 1130 -2676 1130 -2676 0 feedthrough
rlabel pdiffusion 1137 -2676 1137 -2676 0 cellNo=798
rlabel pdiffusion 1144 -2676 1144 -2676 0 feedthrough
rlabel pdiffusion 1151 -2676 1151 -2676 0 feedthrough
rlabel pdiffusion 1158 -2676 1158 -2676 0 feedthrough
rlabel pdiffusion 1165 -2676 1165 -2676 0 feedthrough
rlabel pdiffusion 1172 -2676 1172 -2676 0 feedthrough
rlabel pdiffusion 1179 -2676 1179 -2676 0 feedthrough
rlabel pdiffusion 1186 -2676 1186 -2676 0 cellNo=975
rlabel pdiffusion 1193 -2676 1193 -2676 0 cellNo=270
rlabel pdiffusion 1200 -2676 1200 -2676 0 feedthrough
rlabel pdiffusion 1207 -2676 1207 -2676 0 feedthrough
rlabel pdiffusion 1214 -2676 1214 -2676 0 feedthrough
rlabel pdiffusion 1221 -2676 1221 -2676 0 feedthrough
rlabel pdiffusion 1228 -2676 1228 -2676 0 feedthrough
rlabel pdiffusion 1235 -2676 1235 -2676 0 cellNo=400
rlabel pdiffusion 1242 -2676 1242 -2676 0 cellNo=889
rlabel pdiffusion 1249 -2676 1249 -2676 0 feedthrough
rlabel pdiffusion 1256 -2676 1256 -2676 0 feedthrough
rlabel pdiffusion 1263 -2676 1263 -2676 0 feedthrough
rlabel pdiffusion 1270 -2676 1270 -2676 0 feedthrough
rlabel pdiffusion 1277 -2676 1277 -2676 0 feedthrough
rlabel pdiffusion 1284 -2676 1284 -2676 0 feedthrough
rlabel pdiffusion 1291 -2676 1291 -2676 0 feedthrough
rlabel pdiffusion 1298 -2676 1298 -2676 0 feedthrough
rlabel pdiffusion 1305 -2676 1305 -2676 0 feedthrough
rlabel pdiffusion 1312 -2676 1312 -2676 0 cellNo=49
rlabel pdiffusion 1319 -2676 1319 -2676 0 feedthrough
rlabel pdiffusion 1326 -2676 1326 -2676 0 cellNo=431
rlabel pdiffusion 1333 -2676 1333 -2676 0 feedthrough
rlabel pdiffusion 1340 -2676 1340 -2676 0 feedthrough
rlabel pdiffusion 1347 -2676 1347 -2676 0 feedthrough
rlabel pdiffusion 1354 -2676 1354 -2676 0 feedthrough
rlabel pdiffusion 1361 -2676 1361 -2676 0 feedthrough
rlabel pdiffusion 1368 -2676 1368 -2676 0 feedthrough
rlabel pdiffusion 1375 -2676 1375 -2676 0 feedthrough
rlabel pdiffusion 1382 -2676 1382 -2676 0 feedthrough
rlabel pdiffusion 1389 -2676 1389 -2676 0 feedthrough
rlabel pdiffusion 1396 -2676 1396 -2676 0 cellNo=171
rlabel pdiffusion 1403 -2676 1403 -2676 0 feedthrough
rlabel pdiffusion 1410 -2676 1410 -2676 0 cellNo=108
rlabel pdiffusion 1417 -2676 1417 -2676 0 feedthrough
rlabel pdiffusion 1424 -2676 1424 -2676 0 feedthrough
rlabel pdiffusion 1431 -2676 1431 -2676 0 cellNo=716
rlabel pdiffusion 1438 -2676 1438 -2676 0 cellNo=376
rlabel pdiffusion 1445 -2676 1445 -2676 0 cellNo=935
rlabel pdiffusion 1452 -2676 1452 -2676 0 feedthrough
rlabel pdiffusion 1459 -2676 1459 -2676 0 feedthrough
rlabel pdiffusion 1466 -2676 1466 -2676 0 feedthrough
rlabel pdiffusion 1473 -2676 1473 -2676 0 feedthrough
rlabel pdiffusion 1480 -2676 1480 -2676 0 feedthrough
rlabel pdiffusion 1487 -2676 1487 -2676 0 feedthrough
rlabel pdiffusion 1494 -2676 1494 -2676 0 feedthrough
rlabel pdiffusion 1501 -2676 1501 -2676 0 feedthrough
rlabel pdiffusion 1508 -2676 1508 -2676 0 cellNo=809
rlabel pdiffusion 1515 -2676 1515 -2676 0 feedthrough
rlabel pdiffusion 1522 -2676 1522 -2676 0 feedthrough
rlabel pdiffusion 1529 -2676 1529 -2676 0 feedthrough
rlabel pdiffusion 1536 -2676 1536 -2676 0 feedthrough
rlabel pdiffusion 1543 -2676 1543 -2676 0 feedthrough
rlabel pdiffusion 1550 -2676 1550 -2676 0 feedthrough
rlabel pdiffusion 1557 -2676 1557 -2676 0 feedthrough
rlabel pdiffusion 1564 -2676 1564 -2676 0 feedthrough
rlabel pdiffusion 1571 -2676 1571 -2676 0 feedthrough
rlabel pdiffusion 1578 -2676 1578 -2676 0 cellNo=994
rlabel pdiffusion 1585 -2676 1585 -2676 0 feedthrough
rlabel pdiffusion 1592 -2676 1592 -2676 0 feedthrough
rlabel pdiffusion 1599 -2676 1599 -2676 0 feedthrough
rlabel pdiffusion 1606 -2676 1606 -2676 0 feedthrough
rlabel pdiffusion 1613 -2676 1613 -2676 0 feedthrough
rlabel pdiffusion 1620 -2676 1620 -2676 0 feedthrough
rlabel pdiffusion 1627 -2676 1627 -2676 0 feedthrough
rlabel pdiffusion 1634 -2676 1634 -2676 0 feedthrough
rlabel pdiffusion 1641 -2676 1641 -2676 0 feedthrough
rlabel pdiffusion 1648 -2676 1648 -2676 0 feedthrough
rlabel pdiffusion 1655 -2676 1655 -2676 0 feedthrough
rlabel pdiffusion 1662 -2676 1662 -2676 0 feedthrough
rlabel pdiffusion 1669 -2676 1669 -2676 0 feedthrough
rlabel pdiffusion 1676 -2676 1676 -2676 0 feedthrough
rlabel pdiffusion 1683 -2676 1683 -2676 0 feedthrough
rlabel pdiffusion 1690 -2676 1690 -2676 0 feedthrough
rlabel pdiffusion 1697 -2676 1697 -2676 0 feedthrough
rlabel pdiffusion 1704 -2676 1704 -2676 0 feedthrough
rlabel pdiffusion 1711 -2676 1711 -2676 0 feedthrough
rlabel pdiffusion 1718 -2676 1718 -2676 0 feedthrough
rlabel pdiffusion 1725 -2676 1725 -2676 0 feedthrough
rlabel pdiffusion 1732 -2676 1732 -2676 0 feedthrough
rlabel pdiffusion 1739 -2676 1739 -2676 0 feedthrough
rlabel pdiffusion 1746 -2676 1746 -2676 0 feedthrough
rlabel pdiffusion 1753 -2676 1753 -2676 0 cellNo=162
rlabel pdiffusion 1760 -2676 1760 -2676 0 feedthrough
rlabel pdiffusion 1767 -2676 1767 -2676 0 feedthrough
rlabel pdiffusion 1774 -2676 1774 -2676 0 feedthrough
rlabel pdiffusion 1781 -2676 1781 -2676 0 feedthrough
rlabel pdiffusion 1788 -2676 1788 -2676 0 feedthrough
rlabel pdiffusion 1795 -2676 1795 -2676 0 feedthrough
rlabel pdiffusion 1802 -2676 1802 -2676 0 feedthrough
rlabel pdiffusion 1809 -2676 1809 -2676 0 feedthrough
rlabel pdiffusion 1816 -2676 1816 -2676 0 feedthrough
rlabel pdiffusion 1823 -2676 1823 -2676 0 feedthrough
rlabel pdiffusion 1830 -2676 1830 -2676 0 feedthrough
rlabel pdiffusion 1837 -2676 1837 -2676 0 feedthrough
rlabel pdiffusion 1844 -2676 1844 -2676 0 feedthrough
rlabel pdiffusion 1851 -2676 1851 -2676 0 feedthrough
rlabel pdiffusion 1858 -2676 1858 -2676 0 feedthrough
rlabel pdiffusion 1865 -2676 1865 -2676 0 feedthrough
rlabel pdiffusion 1872 -2676 1872 -2676 0 feedthrough
rlabel pdiffusion 1879 -2676 1879 -2676 0 feedthrough
rlabel pdiffusion 1886 -2676 1886 -2676 0 feedthrough
rlabel pdiffusion 1893 -2676 1893 -2676 0 feedthrough
rlabel pdiffusion 1900 -2676 1900 -2676 0 feedthrough
rlabel pdiffusion 1907 -2676 1907 -2676 0 feedthrough
rlabel pdiffusion 1914 -2676 1914 -2676 0 feedthrough
rlabel pdiffusion 1921 -2676 1921 -2676 0 feedthrough
rlabel pdiffusion 1928 -2676 1928 -2676 0 feedthrough
rlabel pdiffusion 1935 -2676 1935 -2676 0 feedthrough
rlabel pdiffusion 1942 -2676 1942 -2676 0 feedthrough
rlabel pdiffusion 1949 -2676 1949 -2676 0 feedthrough
rlabel pdiffusion 1956 -2676 1956 -2676 0 feedthrough
rlabel pdiffusion 1963 -2676 1963 -2676 0 feedthrough
rlabel pdiffusion 1970 -2676 1970 -2676 0 feedthrough
rlabel pdiffusion 1977 -2676 1977 -2676 0 feedthrough
rlabel pdiffusion 1984 -2676 1984 -2676 0 feedthrough
rlabel pdiffusion 1991 -2676 1991 -2676 0 feedthrough
rlabel pdiffusion 1998 -2676 1998 -2676 0 feedthrough
rlabel pdiffusion 2005 -2676 2005 -2676 0 feedthrough
rlabel pdiffusion 2012 -2676 2012 -2676 0 feedthrough
rlabel pdiffusion 2019 -2676 2019 -2676 0 feedthrough
rlabel pdiffusion 2026 -2676 2026 -2676 0 feedthrough
rlabel pdiffusion 2033 -2676 2033 -2676 0 feedthrough
rlabel pdiffusion 2040 -2676 2040 -2676 0 feedthrough
rlabel pdiffusion 2047 -2676 2047 -2676 0 feedthrough
rlabel pdiffusion 2054 -2676 2054 -2676 0 feedthrough
rlabel pdiffusion 2061 -2676 2061 -2676 0 feedthrough
rlabel pdiffusion 2068 -2676 2068 -2676 0 feedthrough
rlabel pdiffusion 2075 -2676 2075 -2676 0 feedthrough
rlabel pdiffusion 2082 -2676 2082 -2676 0 feedthrough
rlabel pdiffusion 2089 -2676 2089 -2676 0 feedthrough
rlabel pdiffusion 2096 -2676 2096 -2676 0 feedthrough
rlabel pdiffusion 2103 -2676 2103 -2676 0 feedthrough
rlabel pdiffusion 2110 -2676 2110 -2676 0 feedthrough
rlabel pdiffusion 2117 -2676 2117 -2676 0 feedthrough
rlabel pdiffusion 2124 -2676 2124 -2676 0 feedthrough
rlabel pdiffusion 2131 -2676 2131 -2676 0 feedthrough
rlabel pdiffusion 2138 -2676 2138 -2676 0 feedthrough
rlabel pdiffusion 2145 -2676 2145 -2676 0 feedthrough
rlabel pdiffusion 2152 -2676 2152 -2676 0 feedthrough
rlabel pdiffusion 2159 -2676 2159 -2676 0 feedthrough
rlabel pdiffusion 2166 -2676 2166 -2676 0 feedthrough
rlabel pdiffusion 2173 -2676 2173 -2676 0 feedthrough
rlabel pdiffusion 2180 -2676 2180 -2676 0 feedthrough
rlabel pdiffusion 2187 -2676 2187 -2676 0 feedthrough
rlabel pdiffusion 2194 -2676 2194 -2676 0 feedthrough
rlabel pdiffusion 2201 -2676 2201 -2676 0 feedthrough
rlabel pdiffusion 2208 -2676 2208 -2676 0 feedthrough
rlabel pdiffusion 2215 -2676 2215 -2676 0 feedthrough
rlabel pdiffusion 2222 -2676 2222 -2676 0 feedthrough
rlabel pdiffusion 2229 -2676 2229 -2676 0 feedthrough
rlabel pdiffusion 2236 -2676 2236 -2676 0 feedthrough
rlabel pdiffusion 2243 -2676 2243 -2676 0 feedthrough
rlabel pdiffusion 2264 -2676 2264 -2676 0 feedthrough
rlabel pdiffusion 2271 -2676 2271 -2676 0 feedthrough
rlabel pdiffusion 3 -2839 3 -2839 0 feedthrough
rlabel pdiffusion 10 -2839 10 -2839 0 feedthrough
rlabel pdiffusion 17 -2839 17 -2839 0 feedthrough
rlabel pdiffusion 24 -2839 24 -2839 0 feedthrough
rlabel pdiffusion 31 -2839 31 -2839 0 feedthrough
rlabel pdiffusion 38 -2839 38 -2839 0 feedthrough
rlabel pdiffusion 45 -2839 45 -2839 0 feedthrough
rlabel pdiffusion 52 -2839 52 -2839 0 cellNo=769
rlabel pdiffusion 59 -2839 59 -2839 0 feedthrough
rlabel pdiffusion 66 -2839 66 -2839 0 feedthrough
rlabel pdiffusion 73 -2839 73 -2839 0 feedthrough
rlabel pdiffusion 80 -2839 80 -2839 0 cellNo=327
rlabel pdiffusion 87 -2839 87 -2839 0 feedthrough
rlabel pdiffusion 94 -2839 94 -2839 0 feedthrough
rlabel pdiffusion 101 -2839 101 -2839 0 feedthrough
rlabel pdiffusion 108 -2839 108 -2839 0 cellNo=925
rlabel pdiffusion 115 -2839 115 -2839 0 feedthrough
rlabel pdiffusion 122 -2839 122 -2839 0 feedthrough
rlabel pdiffusion 129 -2839 129 -2839 0 feedthrough
rlabel pdiffusion 136 -2839 136 -2839 0 feedthrough
rlabel pdiffusion 143 -2839 143 -2839 0 feedthrough
rlabel pdiffusion 150 -2839 150 -2839 0 feedthrough
rlabel pdiffusion 157 -2839 157 -2839 0 feedthrough
rlabel pdiffusion 164 -2839 164 -2839 0 feedthrough
rlabel pdiffusion 171 -2839 171 -2839 0 feedthrough
rlabel pdiffusion 178 -2839 178 -2839 0 feedthrough
rlabel pdiffusion 185 -2839 185 -2839 0 feedthrough
rlabel pdiffusion 192 -2839 192 -2839 0 feedthrough
rlabel pdiffusion 199 -2839 199 -2839 0 feedthrough
rlabel pdiffusion 206 -2839 206 -2839 0 feedthrough
rlabel pdiffusion 213 -2839 213 -2839 0 feedthrough
rlabel pdiffusion 220 -2839 220 -2839 0 cellNo=929
rlabel pdiffusion 227 -2839 227 -2839 0 feedthrough
rlabel pdiffusion 234 -2839 234 -2839 0 cellNo=204
rlabel pdiffusion 241 -2839 241 -2839 0 feedthrough
rlabel pdiffusion 248 -2839 248 -2839 0 cellNo=827
rlabel pdiffusion 255 -2839 255 -2839 0 feedthrough
rlabel pdiffusion 262 -2839 262 -2839 0 feedthrough
rlabel pdiffusion 269 -2839 269 -2839 0 feedthrough
rlabel pdiffusion 276 -2839 276 -2839 0 feedthrough
rlabel pdiffusion 283 -2839 283 -2839 0 feedthrough
rlabel pdiffusion 290 -2839 290 -2839 0 feedthrough
rlabel pdiffusion 297 -2839 297 -2839 0 feedthrough
rlabel pdiffusion 304 -2839 304 -2839 0 feedthrough
rlabel pdiffusion 311 -2839 311 -2839 0 feedthrough
rlabel pdiffusion 318 -2839 318 -2839 0 feedthrough
rlabel pdiffusion 325 -2839 325 -2839 0 feedthrough
rlabel pdiffusion 332 -2839 332 -2839 0 feedthrough
rlabel pdiffusion 339 -2839 339 -2839 0 feedthrough
rlabel pdiffusion 346 -2839 346 -2839 0 feedthrough
rlabel pdiffusion 353 -2839 353 -2839 0 feedthrough
rlabel pdiffusion 360 -2839 360 -2839 0 feedthrough
rlabel pdiffusion 367 -2839 367 -2839 0 feedthrough
rlabel pdiffusion 374 -2839 374 -2839 0 feedthrough
rlabel pdiffusion 381 -2839 381 -2839 0 feedthrough
rlabel pdiffusion 388 -2839 388 -2839 0 feedthrough
rlabel pdiffusion 395 -2839 395 -2839 0 feedthrough
rlabel pdiffusion 402 -2839 402 -2839 0 feedthrough
rlabel pdiffusion 409 -2839 409 -2839 0 feedthrough
rlabel pdiffusion 416 -2839 416 -2839 0 feedthrough
rlabel pdiffusion 423 -2839 423 -2839 0 feedthrough
rlabel pdiffusion 430 -2839 430 -2839 0 cellNo=75
rlabel pdiffusion 437 -2839 437 -2839 0 feedthrough
rlabel pdiffusion 444 -2839 444 -2839 0 feedthrough
rlabel pdiffusion 451 -2839 451 -2839 0 feedthrough
rlabel pdiffusion 458 -2839 458 -2839 0 cellNo=727
rlabel pdiffusion 465 -2839 465 -2839 0 feedthrough
rlabel pdiffusion 472 -2839 472 -2839 0 feedthrough
rlabel pdiffusion 479 -2839 479 -2839 0 feedthrough
rlabel pdiffusion 486 -2839 486 -2839 0 feedthrough
rlabel pdiffusion 493 -2839 493 -2839 0 feedthrough
rlabel pdiffusion 500 -2839 500 -2839 0 feedthrough
rlabel pdiffusion 507 -2839 507 -2839 0 feedthrough
rlabel pdiffusion 514 -2839 514 -2839 0 feedthrough
rlabel pdiffusion 521 -2839 521 -2839 0 feedthrough
rlabel pdiffusion 528 -2839 528 -2839 0 feedthrough
rlabel pdiffusion 535 -2839 535 -2839 0 feedthrough
rlabel pdiffusion 542 -2839 542 -2839 0 cellNo=533
rlabel pdiffusion 549 -2839 549 -2839 0 feedthrough
rlabel pdiffusion 556 -2839 556 -2839 0 feedthrough
rlabel pdiffusion 563 -2839 563 -2839 0 feedthrough
rlabel pdiffusion 570 -2839 570 -2839 0 feedthrough
rlabel pdiffusion 577 -2839 577 -2839 0 feedthrough
rlabel pdiffusion 584 -2839 584 -2839 0 feedthrough
rlabel pdiffusion 591 -2839 591 -2839 0 feedthrough
rlabel pdiffusion 598 -2839 598 -2839 0 feedthrough
rlabel pdiffusion 605 -2839 605 -2839 0 feedthrough
rlabel pdiffusion 612 -2839 612 -2839 0 feedthrough
rlabel pdiffusion 619 -2839 619 -2839 0 cellNo=655
rlabel pdiffusion 626 -2839 626 -2839 0 feedthrough
rlabel pdiffusion 633 -2839 633 -2839 0 feedthrough
rlabel pdiffusion 640 -2839 640 -2839 0 feedthrough
rlabel pdiffusion 647 -2839 647 -2839 0 feedthrough
rlabel pdiffusion 654 -2839 654 -2839 0 feedthrough
rlabel pdiffusion 661 -2839 661 -2839 0 cellNo=266
rlabel pdiffusion 668 -2839 668 -2839 0 feedthrough
rlabel pdiffusion 675 -2839 675 -2839 0 feedthrough
rlabel pdiffusion 682 -2839 682 -2839 0 feedthrough
rlabel pdiffusion 689 -2839 689 -2839 0 feedthrough
rlabel pdiffusion 696 -2839 696 -2839 0 feedthrough
rlabel pdiffusion 703 -2839 703 -2839 0 cellNo=290
rlabel pdiffusion 710 -2839 710 -2839 0 feedthrough
rlabel pdiffusion 717 -2839 717 -2839 0 feedthrough
rlabel pdiffusion 724 -2839 724 -2839 0 feedthrough
rlabel pdiffusion 731 -2839 731 -2839 0 cellNo=50
rlabel pdiffusion 738 -2839 738 -2839 0 feedthrough
rlabel pdiffusion 745 -2839 745 -2839 0 cellNo=419
rlabel pdiffusion 752 -2839 752 -2839 0 feedthrough
rlabel pdiffusion 759 -2839 759 -2839 0 feedthrough
rlabel pdiffusion 766 -2839 766 -2839 0 feedthrough
rlabel pdiffusion 773 -2839 773 -2839 0 feedthrough
rlabel pdiffusion 780 -2839 780 -2839 0 feedthrough
rlabel pdiffusion 787 -2839 787 -2839 0 cellNo=767
rlabel pdiffusion 794 -2839 794 -2839 0 feedthrough
rlabel pdiffusion 801 -2839 801 -2839 0 feedthrough
rlabel pdiffusion 808 -2839 808 -2839 0 feedthrough
rlabel pdiffusion 815 -2839 815 -2839 0 feedthrough
rlabel pdiffusion 822 -2839 822 -2839 0 feedthrough
rlabel pdiffusion 829 -2839 829 -2839 0 feedthrough
rlabel pdiffusion 836 -2839 836 -2839 0 cellNo=931
rlabel pdiffusion 843 -2839 843 -2839 0 feedthrough
rlabel pdiffusion 850 -2839 850 -2839 0 feedthrough
rlabel pdiffusion 857 -2839 857 -2839 0 feedthrough
rlabel pdiffusion 864 -2839 864 -2839 0 cellNo=915
rlabel pdiffusion 871 -2839 871 -2839 0 feedthrough
rlabel pdiffusion 878 -2839 878 -2839 0 feedthrough
rlabel pdiffusion 885 -2839 885 -2839 0 feedthrough
rlabel pdiffusion 892 -2839 892 -2839 0 feedthrough
rlabel pdiffusion 899 -2839 899 -2839 0 feedthrough
rlabel pdiffusion 906 -2839 906 -2839 0 feedthrough
rlabel pdiffusion 913 -2839 913 -2839 0 cellNo=838
rlabel pdiffusion 920 -2839 920 -2839 0 feedthrough
rlabel pdiffusion 927 -2839 927 -2839 0 feedthrough
rlabel pdiffusion 934 -2839 934 -2839 0 feedthrough
rlabel pdiffusion 941 -2839 941 -2839 0 cellNo=961
rlabel pdiffusion 948 -2839 948 -2839 0 feedthrough
rlabel pdiffusion 955 -2839 955 -2839 0 feedthrough
rlabel pdiffusion 962 -2839 962 -2839 0 cellNo=34
rlabel pdiffusion 969 -2839 969 -2839 0 feedthrough
rlabel pdiffusion 976 -2839 976 -2839 0 cellNo=429
rlabel pdiffusion 983 -2839 983 -2839 0 feedthrough
rlabel pdiffusion 990 -2839 990 -2839 0 feedthrough
rlabel pdiffusion 997 -2839 997 -2839 0 feedthrough
rlabel pdiffusion 1004 -2839 1004 -2839 0 feedthrough
rlabel pdiffusion 1011 -2839 1011 -2839 0 feedthrough
rlabel pdiffusion 1018 -2839 1018 -2839 0 feedthrough
rlabel pdiffusion 1025 -2839 1025 -2839 0 feedthrough
rlabel pdiffusion 1032 -2839 1032 -2839 0 feedthrough
rlabel pdiffusion 1039 -2839 1039 -2839 0 feedthrough
rlabel pdiffusion 1046 -2839 1046 -2839 0 feedthrough
rlabel pdiffusion 1053 -2839 1053 -2839 0 cellNo=704
rlabel pdiffusion 1060 -2839 1060 -2839 0 cellNo=868
rlabel pdiffusion 1067 -2839 1067 -2839 0 feedthrough
rlabel pdiffusion 1074 -2839 1074 -2839 0 feedthrough
rlabel pdiffusion 1081 -2839 1081 -2839 0 feedthrough
rlabel pdiffusion 1088 -2839 1088 -2839 0 feedthrough
rlabel pdiffusion 1095 -2839 1095 -2839 0 cellNo=388
rlabel pdiffusion 1102 -2839 1102 -2839 0 feedthrough
rlabel pdiffusion 1109 -2839 1109 -2839 0 feedthrough
rlabel pdiffusion 1116 -2839 1116 -2839 0 feedthrough
rlabel pdiffusion 1123 -2839 1123 -2839 0 feedthrough
rlabel pdiffusion 1130 -2839 1130 -2839 0 feedthrough
rlabel pdiffusion 1137 -2839 1137 -2839 0 feedthrough
rlabel pdiffusion 1144 -2839 1144 -2839 0 feedthrough
rlabel pdiffusion 1151 -2839 1151 -2839 0 feedthrough
rlabel pdiffusion 1158 -2839 1158 -2839 0 feedthrough
rlabel pdiffusion 1165 -2839 1165 -2839 0 feedthrough
rlabel pdiffusion 1172 -2839 1172 -2839 0 feedthrough
rlabel pdiffusion 1179 -2839 1179 -2839 0 feedthrough
rlabel pdiffusion 1186 -2839 1186 -2839 0 feedthrough
rlabel pdiffusion 1193 -2839 1193 -2839 0 feedthrough
rlabel pdiffusion 1200 -2839 1200 -2839 0 feedthrough
rlabel pdiffusion 1207 -2839 1207 -2839 0 feedthrough
rlabel pdiffusion 1214 -2839 1214 -2839 0 feedthrough
rlabel pdiffusion 1221 -2839 1221 -2839 0 feedthrough
rlabel pdiffusion 1228 -2839 1228 -2839 0 feedthrough
rlabel pdiffusion 1235 -2839 1235 -2839 0 feedthrough
rlabel pdiffusion 1242 -2839 1242 -2839 0 feedthrough
rlabel pdiffusion 1249 -2839 1249 -2839 0 feedthrough
rlabel pdiffusion 1256 -2839 1256 -2839 0 cellNo=131
rlabel pdiffusion 1263 -2839 1263 -2839 0 feedthrough
rlabel pdiffusion 1270 -2839 1270 -2839 0 feedthrough
rlabel pdiffusion 1277 -2839 1277 -2839 0 feedthrough
rlabel pdiffusion 1284 -2839 1284 -2839 0 cellNo=983
rlabel pdiffusion 1291 -2839 1291 -2839 0 feedthrough
rlabel pdiffusion 1298 -2839 1298 -2839 0 feedthrough
rlabel pdiffusion 1305 -2839 1305 -2839 0 feedthrough
rlabel pdiffusion 1312 -2839 1312 -2839 0 cellNo=227
rlabel pdiffusion 1319 -2839 1319 -2839 0 feedthrough
rlabel pdiffusion 1326 -2839 1326 -2839 0 feedthrough
rlabel pdiffusion 1333 -2839 1333 -2839 0 feedthrough
rlabel pdiffusion 1340 -2839 1340 -2839 0 feedthrough
rlabel pdiffusion 1347 -2839 1347 -2839 0 cellNo=488
rlabel pdiffusion 1354 -2839 1354 -2839 0 feedthrough
rlabel pdiffusion 1361 -2839 1361 -2839 0 feedthrough
rlabel pdiffusion 1368 -2839 1368 -2839 0 feedthrough
rlabel pdiffusion 1375 -2839 1375 -2839 0 feedthrough
rlabel pdiffusion 1382 -2839 1382 -2839 0 feedthrough
rlabel pdiffusion 1389 -2839 1389 -2839 0 cellNo=222
rlabel pdiffusion 1396 -2839 1396 -2839 0 feedthrough
rlabel pdiffusion 1403 -2839 1403 -2839 0 feedthrough
rlabel pdiffusion 1410 -2839 1410 -2839 0 feedthrough
rlabel pdiffusion 1417 -2839 1417 -2839 0 feedthrough
rlabel pdiffusion 1424 -2839 1424 -2839 0 feedthrough
rlabel pdiffusion 1431 -2839 1431 -2839 0 cellNo=325
rlabel pdiffusion 1438 -2839 1438 -2839 0 feedthrough
rlabel pdiffusion 1445 -2839 1445 -2839 0 feedthrough
rlabel pdiffusion 1452 -2839 1452 -2839 0 cellNo=297
rlabel pdiffusion 1459 -2839 1459 -2839 0 feedthrough
rlabel pdiffusion 1466 -2839 1466 -2839 0 feedthrough
rlabel pdiffusion 1473 -2839 1473 -2839 0 feedthrough
rlabel pdiffusion 1480 -2839 1480 -2839 0 feedthrough
rlabel pdiffusion 1487 -2839 1487 -2839 0 cellNo=255
rlabel pdiffusion 1494 -2839 1494 -2839 0 cellNo=570
rlabel pdiffusion 1501 -2839 1501 -2839 0 feedthrough
rlabel pdiffusion 1508 -2839 1508 -2839 0 feedthrough
rlabel pdiffusion 1515 -2839 1515 -2839 0 feedthrough
rlabel pdiffusion 1522 -2839 1522 -2839 0 feedthrough
rlabel pdiffusion 1529 -2839 1529 -2839 0 feedthrough
rlabel pdiffusion 1536 -2839 1536 -2839 0 feedthrough
rlabel pdiffusion 1543 -2839 1543 -2839 0 feedthrough
rlabel pdiffusion 1550 -2839 1550 -2839 0 feedthrough
rlabel pdiffusion 1557 -2839 1557 -2839 0 feedthrough
rlabel pdiffusion 1564 -2839 1564 -2839 0 cellNo=544
rlabel pdiffusion 1571 -2839 1571 -2839 0 feedthrough
rlabel pdiffusion 1578 -2839 1578 -2839 0 feedthrough
rlabel pdiffusion 1585 -2839 1585 -2839 0 feedthrough
rlabel pdiffusion 1592 -2839 1592 -2839 0 feedthrough
rlabel pdiffusion 1599 -2839 1599 -2839 0 feedthrough
rlabel pdiffusion 1606 -2839 1606 -2839 0 feedthrough
rlabel pdiffusion 1613 -2839 1613 -2839 0 feedthrough
rlabel pdiffusion 1620 -2839 1620 -2839 0 feedthrough
rlabel pdiffusion 1627 -2839 1627 -2839 0 feedthrough
rlabel pdiffusion 1634 -2839 1634 -2839 0 feedthrough
rlabel pdiffusion 1641 -2839 1641 -2839 0 feedthrough
rlabel pdiffusion 1648 -2839 1648 -2839 0 feedthrough
rlabel pdiffusion 1655 -2839 1655 -2839 0 feedthrough
rlabel pdiffusion 1662 -2839 1662 -2839 0 feedthrough
rlabel pdiffusion 1669 -2839 1669 -2839 0 feedthrough
rlabel pdiffusion 1676 -2839 1676 -2839 0 feedthrough
rlabel pdiffusion 1683 -2839 1683 -2839 0 cellNo=319
rlabel pdiffusion 1690 -2839 1690 -2839 0 feedthrough
rlabel pdiffusion 1697 -2839 1697 -2839 0 feedthrough
rlabel pdiffusion 1704 -2839 1704 -2839 0 cellNo=660
rlabel pdiffusion 1711 -2839 1711 -2839 0 feedthrough
rlabel pdiffusion 1718 -2839 1718 -2839 0 feedthrough
rlabel pdiffusion 1725 -2839 1725 -2839 0 feedthrough
rlabel pdiffusion 1732 -2839 1732 -2839 0 feedthrough
rlabel pdiffusion 1739 -2839 1739 -2839 0 feedthrough
rlabel pdiffusion 1746 -2839 1746 -2839 0 feedthrough
rlabel pdiffusion 1753 -2839 1753 -2839 0 cellNo=905
rlabel pdiffusion 1760 -2839 1760 -2839 0 feedthrough
rlabel pdiffusion 1767 -2839 1767 -2839 0 feedthrough
rlabel pdiffusion 1774 -2839 1774 -2839 0 feedthrough
rlabel pdiffusion 1781 -2839 1781 -2839 0 feedthrough
rlabel pdiffusion 1788 -2839 1788 -2839 0 feedthrough
rlabel pdiffusion 1795 -2839 1795 -2839 0 feedthrough
rlabel pdiffusion 1802 -2839 1802 -2839 0 feedthrough
rlabel pdiffusion 1809 -2839 1809 -2839 0 feedthrough
rlabel pdiffusion 1816 -2839 1816 -2839 0 feedthrough
rlabel pdiffusion 1823 -2839 1823 -2839 0 feedthrough
rlabel pdiffusion 1830 -2839 1830 -2839 0 feedthrough
rlabel pdiffusion 1837 -2839 1837 -2839 0 feedthrough
rlabel pdiffusion 1844 -2839 1844 -2839 0 feedthrough
rlabel pdiffusion 1851 -2839 1851 -2839 0 feedthrough
rlabel pdiffusion 1858 -2839 1858 -2839 0 feedthrough
rlabel pdiffusion 1865 -2839 1865 -2839 0 feedthrough
rlabel pdiffusion 1872 -2839 1872 -2839 0 feedthrough
rlabel pdiffusion 1879 -2839 1879 -2839 0 feedthrough
rlabel pdiffusion 1886 -2839 1886 -2839 0 feedthrough
rlabel pdiffusion 1893 -2839 1893 -2839 0 feedthrough
rlabel pdiffusion 1900 -2839 1900 -2839 0 feedthrough
rlabel pdiffusion 1907 -2839 1907 -2839 0 feedthrough
rlabel pdiffusion 1914 -2839 1914 -2839 0 feedthrough
rlabel pdiffusion 1921 -2839 1921 -2839 0 feedthrough
rlabel pdiffusion 1928 -2839 1928 -2839 0 feedthrough
rlabel pdiffusion 1935 -2839 1935 -2839 0 feedthrough
rlabel pdiffusion 1942 -2839 1942 -2839 0 feedthrough
rlabel pdiffusion 1949 -2839 1949 -2839 0 feedthrough
rlabel pdiffusion 1956 -2839 1956 -2839 0 feedthrough
rlabel pdiffusion 1963 -2839 1963 -2839 0 feedthrough
rlabel pdiffusion 1970 -2839 1970 -2839 0 feedthrough
rlabel pdiffusion 1977 -2839 1977 -2839 0 feedthrough
rlabel pdiffusion 1984 -2839 1984 -2839 0 feedthrough
rlabel pdiffusion 1991 -2839 1991 -2839 0 feedthrough
rlabel pdiffusion 1998 -2839 1998 -2839 0 feedthrough
rlabel pdiffusion 2005 -2839 2005 -2839 0 feedthrough
rlabel pdiffusion 2012 -2839 2012 -2839 0 feedthrough
rlabel pdiffusion 2019 -2839 2019 -2839 0 feedthrough
rlabel pdiffusion 2026 -2839 2026 -2839 0 feedthrough
rlabel pdiffusion 2033 -2839 2033 -2839 0 feedthrough
rlabel pdiffusion 2040 -2839 2040 -2839 0 feedthrough
rlabel pdiffusion 2047 -2839 2047 -2839 0 feedthrough
rlabel pdiffusion 2054 -2839 2054 -2839 0 feedthrough
rlabel pdiffusion 2061 -2839 2061 -2839 0 feedthrough
rlabel pdiffusion 2068 -2839 2068 -2839 0 feedthrough
rlabel pdiffusion 2075 -2839 2075 -2839 0 feedthrough
rlabel pdiffusion 2082 -2839 2082 -2839 0 feedthrough
rlabel pdiffusion 2089 -2839 2089 -2839 0 feedthrough
rlabel pdiffusion 2096 -2839 2096 -2839 0 feedthrough
rlabel pdiffusion 2103 -2839 2103 -2839 0 feedthrough
rlabel pdiffusion 2110 -2839 2110 -2839 0 feedthrough
rlabel pdiffusion 2117 -2839 2117 -2839 0 feedthrough
rlabel pdiffusion 2124 -2839 2124 -2839 0 feedthrough
rlabel pdiffusion 2131 -2839 2131 -2839 0 feedthrough
rlabel pdiffusion 2138 -2839 2138 -2839 0 feedthrough
rlabel pdiffusion 2145 -2839 2145 -2839 0 feedthrough
rlabel pdiffusion 2152 -2839 2152 -2839 0 feedthrough
rlabel pdiffusion 2159 -2839 2159 -2839 0 feedthrough
rlabel pdiffusion 2166 -2839 2166 -2839 0 feedthrough
rlabel pdiffusion 2173 -2839 2173 -2839 0 feedthrough
rlabel pdiffusion 2180 -2839 2180 -2839 0 feedthrough
rlabel pdiffusion 2187 -2839 2187 -2839 0 feedthrough
rlabel pdiffusion 2194 -2839 2194 -2839 0 feedthrough
rlabel pdiffusion 2201 -2839 2201 -2839 0 feedthrough
rlabel pdiffusion 2208 -2839 2208 -2839 0 feedthrough
rlabel pdiffusion 2215 -2839 2215 -2839 0 feedthrough
rlabel pdiffusion 2222 -2839 2222 -2839 0 cellNo=534
rlabel pdiffusion 2229 -2839 2229 -2839 0 feedthrough
rlabel pdiffusion 2236 -2839 2236 -2839 0 feedthrough
rlabel pdiffusion 2243 -2839 2243 -2839 0 feedthrough
rlabel pdiffusion 2250 -2839 2250 -2839 0 feedthrough
rlabel pdiffusion 2257 -2839 2257 -2839 0 cellNo=737
rlabel pdiffusion 2264 -2839 2264 -2839 0 feedthrough
rlabel pdiffusion 2271 -2839 2271 -2839 0 feedthrough
rlabel pdiffusion 3 -2984 3 -2984 0 cellNo=1087
rlabel pdiffusion 10 -2984 10 -2984 0 cellNo=1110
rlabel pdiffusion 17 -2984 17 -2984 0 feedthrough
rlabel pdiffusion 24 -2984 24 -2984 0 feedthrough
rlabel pdiffusion 31 -2984 31 -2984 0 feedthrough
rlabel pdiffusion 38 -2984 38 -2984 0 feedthrough
rlabel pdiffusion 45 -2984 45 -2984 0 feedthrough
rlabel pdiffusion 52 -2984 52 -2984 0 cellNo=487
rlabel pdiffusion 59 -2984 59 -2984 0 feedthrough
rlabel pdiffusion 66 -2984 66 -2984 0 feedthrough
rlabel pdiffusion 73 -2984 73 -2984 0 feedthrough
rlabel pdiffusion 80 -2984 80 -2984 0 feedthrough
rlabel pdiffusion 87 -2984 87 -2984 0 feedthrough
rlabel pdiffusion 94 -2984 94 -2984 0 feedthrough
rlabel pdiffusion 101 -2984 101 -2984 0 cellNo=334
rlabel pdiffusion 108 -2984 108 -2984 0 cellNo=433
rlabel pdiffusion 115 -2984 115 -2984 0 cellNo=618
rlabel pdiffusion 122 -2984 122 -2984 0 cellNo=289
rlabel pdiffusion 129 -2984 129 -2984 0 feedthrough
rlabel pdiffusion 136 -2984 136 -2984 0 feedthrough
rlabel pdiffusion 143 -2984 143 -2984 0 feedthrough
rlabel pdiffusion 150 -2984 150 -2984 0 feedthrough
rlabel pdiffusion 157 -2984 157 -2984 0 cellNo=403
rlabel pdiffusion 164 -2984 164 -2984 0 feedthrough
rlabel pdiffusion 171 -2984 171 -2984 0 feedthrough
rlabel pdiffusion 178 -2984 178 -2984 0 feedthrough
rlabel pdiffusion 185 -2984 185 -2984 0 feedthrough
rlabel pdiffusion 192 -2984 192 -2984 0 feedthrough
rlabel pdiffusion 199 -2984 199 -2984 0 feedthrough
rlabel pdiffusion 206 -2984 206 -2984 0 feedthrough
rlabel pdiffusion 213 -2984 213 -2984 0 cellNo=989
rlabel pdiffusion 220 -2984 220 -2984 0 feedthrough
rlabel pdiffusion 227 -2984 227 -2984 0 feedthrough
rlabel pdiffusion 234 -2984 234 -2984 0 feedthrough
rlabel pdiffusion 241 -2984 241 -2984 0 feedthrough
rlabel pdiffusion 248 -2984 248 -2984 0 feedthrough
rlabel pdiffusion 255 -2984 255 -2984 0 cellNo=870
rlabel pdiffusion 262 -2984 262 -2984 0 feedthrough
rlabel pdiffusion 269 -2984 269 -2984 0 feedthrough
rlabel pdiffusion 276 -2984 276 -2984 0 feedthrough
rlabel pdiffusion 283 -2984 283 -2984 0 feedthrough
rlabel pdiffusion 290 -2984 290 -2984 0 feedthrough
rlabel pdiffusion 297 -2984 297 -2984 0 feedthrough
rlabel pdiffusion 304 -2984 304 -2984 0 feedthrough
rlabel pdiffusion 311 -2984 311 -2984 0 feedthrough
rlabel pdiffusion 318 -2984 318 -2984 0 feedthrough
rlabel pdiffusion 325 -2984 325 -2984 0 feedthrough
rlabel pdiffusion 332 -2984 332 -2984 0 feedthrough
rlabel pdiffusion 339 -2984 339 -2984 0 feedthrough
rlabel pdiffusion 346 -2984 346 -2984 0 feedthrough
rlabel pdiffusion 353 -2984 353 -2984 0 feedthrough
rlabel pdiffusion 360 -2984 360 -2984 0 feedthrough
rlabel pdiffusion 367 -2984 367 -2984 0 feedthrough
rlabel pdiffusion 374 -2984 374 -2984 0 feedthrough
rlabel pdiffusion 381 -2984 381 -2984 0 feedthrough
rlabel pdiffusion 388 -2984 388 -2984 0 feedthrough
rlabel pdiffusion 395 -2984 395 -2984 0 feedthrough
rlabel pdiffusion 402 -2984 402 -2984 0 feedthrough
rlabel pdiffusion 409 -2984 409 -2984 0 feedthrough
rlabel pdiffusion 416 -2984 416 -2984 0 feedthrough
rlabel pdiffusion 423 -2984 423 -2984 0 feedthrough
rlabel pdiffusion 430 -2984 430 -2984 0 feedthrough
rlabel pdiffusion 437 -2984 437 -2984 0 feedthrough
rlabel pdiffusion 444 -2984 444 -2984 0 feedthrough
rlabel pdiffusion 451 -2984 451 -2984 0 feedthrough
rlabel pdiffusion 458 -2984 458 -2984 0 feedthrough
rlabel pdiffusion 465 -2984 465 -2984 0 cellNo=22
rlabel pdiffusion 472 -2984 472 -2984 0 feedthrough
rlabel pdiffusion 479 -2984 479 -2984 0 feedthrough
rlabel pdiffusion 486 -2984 486 -2984 0 feedthrough
rlabel pdiffusion 493 -2984 493 -2984 0 feedthrough
rlabel pdiffusion 500 -2984 500 -2984 0 feedthrough
rlabel pdiffusion 507 -2984 507 -2984 0 feedthrough
rlabel pdiffusion 514 -2984 514 -2984 0 feedthrough
rlabel pdiffusion 521 -2984 521 -2984 0 feedthrough
rlabel pdiffusion 528 -2984 528 -2984 0 feedthrough
rlabel pdiffusion 535 -2984 535 -2984 0 feedthrough
rlabel pdiffusion 542 -2984 542 -2984 0 cellNo=851
rlabel pdiffusion 549 -2984 549 -2984 0 feedthrough
rlabel pdiffusion 556 -2984 556 -2984 0 feedthrough
rlabel pdiffusion 563 -2984 563 -2984 0 cellNo=872
rlabel pdiffusion 570 -2984 570 -2984 0 cellNo=432
rlabel pdiffusion 577 -2984 577 -2984 0 feedthrough
rlabel pdiffusion 584 -2984 584 -2984 0 feedthrough
rlabel pdiffusion 591 -2984 591 -2984 0 feedthrough
rlabel pdiffusion 598 -2984 598 -2984 0 feedthrough
rlabel pdiffusion 605 -2984 605 -2984 0 feedthrough
rlabel pdiffusion 612 -2984 612 -2984 0 feedthrough
rlabel pdiffusion 619 -2984 619 -2984 0 feedthrough
rlabel pdiffusion 626 -2984 626 -2984 0 feedthrough
rlabel pdiffusion 633 -2984 633 -2984 0 feedthrough
rlabel pdiffusion 640 -2984 640 -2984 0 cellNo=599
rlabel pdiffusion 647 -2984 647 -2984 0 feedthrough
rlabel pdiffusion 654 -2984 654 -2984 0 feedthrough
rlabel pdiffusion 661 -2984 661 -2984 0 cellNo=963
rlabel pdiffusion 668 -2984 668 -2984 0 feedthrough
rlabel pdiffusion 675 -2984 675 -2984 0 feedthrough
rlabel pdiffusion 682 -2984 682 -2984 0 feedthrough
rlabel pdiffusion 689 -2984 689 -2984 0 feedthrough
rlabel pdiffusion 696 -2984 696 -2984 0 feedthrough
rlabel pdiffusion 703 -2984 703 -2984 0 feedthrough
rlabel pdiffusion 710 -2984 710 -2984 0 feedthrough
rlabel pdiffusion 717 -2984 717 -2984 0 feedthrough
rlabel pdiffusion 724 -2984 724 -2984 0 feedthrough
rlabel pdiffusion 731 -2984 731 -2984 0 feedthrough
rlabel pdiffusion 738 -2984 738 -2984 0 cellNo=82
rlabel pdiffusion 745 -2984 745 -2984 0 feedthrough
rlabel pdiffusion 752 -2984 752 -2984 0 feedthrough
rlabel pdiffusion 759 -2984 759 -2984 0 feedthrough
rlabel pdiffusion 766 -2984 766 -2984 0 feedthrough
rlabel pdiffusion 773 -2984 773 -2984 0 feedthrough
rlabel pdiffusion 780 -2984 780 -2984 0 feedthrough
rlabel pdiffusion 787 -2984 787 -2984 0 feedthrough
rlabel pdiffusion 794 -2984 794 -2984 0 feedthrough
rlabel pdiffusion 801 -2984 801 -2984 0 feedthrough
rlabel pdiffusion 808 -2984 808 -2984 0 feedthrough
rlabel pdiffusion 815 -2984 815 -2984 0 feedthrough
rlabel pdiffusion 822 -2984 822 -2984 0 feedthrough
rlabel pdiffusion 829 -2984 829 -2984 0 feedthrough
rlabel pdiffusion 836 -2984 836 -2984 0 feedthrough
rlabel pdiffusion 843 -2984 843 -2984 0 feedthrough
rlabel pdiffusion 850 -2984 850 -2984 0 feedthrough
rlabel pdiffusion 857 -2984 857 -2984 0 feedthrough
rlabel pdiffusion 864 -2984 864 -2984 0 feedthrough
rlabel pdiffusion 871 -2984 871 -2984 0 feedthrough
rlabel pdiffusion 878 -2984 878 -2984 0 cellNo=705
rlabel pdiffusion 885 -2984 885 -2984 0 feedthrough
rlabel pdiffusion 892 -2984 892 -2984 0 feedthrough
rlabel pdiffusion 899 -2984 899 -2984 0 feedthrough
rlabel pdiffusion 906 -2984 906 -2984 0 feedthrough
rlabel pdiffusion 913 -2984 913 -2984 0 cellNo=857
rlabel pdiffusion 920 -2984 920 -2984 0 cellNo=417
rlabel pdiffusion 927 -2984 927 -2984 0 feedthrough
rlabel pdiffusion 934 -2984 934 -2984 0 feedthrough
rlabel pdiffusion 941 -2984 941 -2984 0 feedthrough
rlabel pdiffusion 948 -2984 948 -2984 0 feedthrough
rlabel pdiffusion 955 -2984 955 -2984 0 feedthrough
rlabel pdiffusion 962 -2984 962 -2984 0 cellNo=408
rlabel pdiffusion 969 -2984 969 -2984 0 feedthrough
rlabel pdiffusion 976 -2984 976 -2984 0 feedthrough
rlabel pdiffusion 983 -2984 983 -2984 0 cellNo=786
rlabel pdiffusion 990 -2984 990 -2984 0 feedthrough
rlabel pdiffusion 997 -2984 997 -2984 0 feedthrough
rlabel pdiffusion 1004 -2984 1004 -2984 0 feedthrough
rlabel pdiffusion 1011 -2984 1011 -2984 0 feedthrough
rlabel pdiffusion 1018 -2984 1018 -2984 0 feedthrough
rlabel pdiffusion 1025 -2984 1025 -2984 0 feedthrough
rlabel pdiffusion 1032 -2984 1032 -2984 0 cellNo=592
rlabel pdiffusion 1039 -2984 1039 -2984 0 cellNo=296
rlabel pdiffusion 1046 -2984 1046 -2984 0 feedthrough
rlabel pdiffusion 1053 -2984 1053 -2984 0 cellNo=995
rlabel pdiffusion 1060 -2984 1060 -2984 0 cellNo=426
rlabel pdiffusion 1067 -2984 1067 -2984 0 cellNo=946
rlabel pdiffusion 1074 -2984 1074 -2984 0 feedthrough
rlabel pdiffusion 1081 -2984 1081 -2984 0 feedthrough
rlabel pdiffusion 1088 -2984 1088 -2984 0 feedthrough
rlabel pdiffusion 1095 -2984 1095 -2984 0 cellNo=730
rlabel pdiffusion 1102 -2984 1102 -2984 0 feedthrough
rlabel pdiffusion 1109 -2984 1109 -2984 0 feedthrough
rlabel pdiffusion 1116 -2984 1116 -2984 0 feedthrough
rlabel pdiffusion 1123 -2984 1123 -2984 0 cellNo=353
rlabel pdiffusion 1130 -2984 1130 -2984 0 feedthrough
rlabel pdiffusion 1137 -2984 1137 -2984 0 cellNo=867
rlabel pdiffusion 1144 -2984 1144 -2984 0 feedthrough
rlabel pdiffusion 1151 -2984 1151 -2984 0 feedthrough
rlabel pdiffusion 1158 -2984 1158 -2984 0 cellNo=797
rlabel pdiffusion 1165 -2984 1165 -2984 0 feedthrough
rlabel pdiffusion 1172 -2984 1172 -2984 0 feedthrough
rlabel pdiffusion 1179 -2984 1179 -2984 0 feedthrough
rlabel pdiffusion 1186 -2984 1186 -2984 0 feedthrough
rlabel pdiffusion 1193 -2984 1193 -2984 0 feedthrough
rlabel pdiffusion 1200 -2984 1200 -2984 0 cellNo=368
rlabel pdiffusion 1207 -2984 1207 -2984 0 cellNo=250
rlabel pdiffusion 1214 -2984 1214 -2984 0 feedthrough
rlabel pdiffusion 1221 -2984 1221 -2984 0 feedthrough
rlabel pdiffusion 1228 -2984 1228 -2984 0 feedthrough
rlabel pdiffusion 1235 -2984 1235 -2984 0 feedthrough
rlabel pdiffusion 1242 -2984 1242 -2984 0 feedthrough
rlabel pdiffusion 1249 -2984 1249 -2984 0 feedthrough
rlabel pdiffusion 1256 -2984 1256 -2984 0 feedthrough
rlabel pdiffusion 1263 -2984 1263 -2984 0 feedthrough
rlabel pdiffusion 1270 -2984 1270 -2984 0 feedthrough
rlabel pdiffusion 1277 -2984 1277 -2984 0 feedthrough
rlabel pdiffusion 1284 -2984 1284 -2984 0 feedthrough
rlabel pdiffusion 1291 -2984 1291 -2984 0 feedthrough
rlabel pdiffusion 1298 -2984 1298 -2984 0 feedthrough
rlabel pdiffusion 1305 -2984 1305 -2984 0 feedthrough
rlabel pdiffusion 1312 -2984 1312 -2984 0 cellNo=629
rlabel pdiffusion 1319 -2984 1319 -2984 0 feedthrough
rlabel pdiffusion 1326 -2984 1326 -2984 0 feedthrough
rlabel pdiffusion 1333 -2984 1333 -2984 0 feedthrough
rlabel pdiffusion 1340 -2984 1340 -2984 0 feedthrough
rlabel pdiffusion 1347 -2984 1347 -2984 0 feedthrough
rlabel pdiffusion 1354 -2984 1354 -2984 0 feedthrough
rlabel pdiffusion 1361 -2984 1361 -2984 0 cellNo=547
rlabel pdiffusion 1368 -2984 1368 -2984 0 feedthrough
rlabel pdiffusion 1375 -2984 1375 -2984 0 feedthrough
rlabel pdiffusion 1382 -2984 1382 -2984 0 feedthrough
rlabel pdiffusion 1389 -2984 1389 -2984 0 feedthrough
rlabel pdiffusion 1396 -2984 1396 -2984 0 feedthrough
rlabel pdiffusion 1403 -2984 1403 -2984 0 feedthrough
rlabel pdiffusion 1410 -2984 1410 -2984 0 feedthrough
rlabel pdiffusion 1417 -2984 1417 -2984 0 cellNo=830
rlabel pdiffusion 1424 -2984 1424 -2984 0 feedthrough
rlabel pdiffusion 1431 -2984 1431 -2984 0 feedthrough
rlabel pdiffusion 1438 -2984 1438 -2984 0 feedthrough
rlabel pdiffusion 1445 -2984 1445 -2984 0 feedthrough
rlabel pdiffusion 1452 -2984 1452 -2984 0 feedthrough
rlabel pdiffusion 1459 -2984 1459 -2984 0 feedthrough
rlabel pdiffusion 1466 -2984 1466 -2984 0 feedthrough
rlabel pdiffusion 1473 -2984 1473 -2984 0 feedthrough
rlabel pdiffusion 1480 -2984 1480 -2984 0 feedthrough
rlabel pdiffusion 1487 -2984 1487 -2984 0 feedthrough
rlabel pdiffusion 1494 -2984 1494 -2984 0 feedthrough
rlabel pdiffusion 1501 -2984 1501 -2984 0 feedthrough
rlabel pdiffusion 1508 -2984 1508 -2984 0 feedthrough
rlabel pdiffusion 1515 -2984 1515 -2984 0 feedthrough
rlabel pdiffusion 1522 -2984 1522 -2984 0 feedthrough
rlabel pdiffusion 1529 -2984 1529 -2984 0 feedthrough
rlabel pdiffusion 1536 -2984 1536 -2984 0 feedthrough
rlabel pdiffusion 1543 -2984 1543 -2984 0 feedthrough
rlabel pdiffusion 1550 -2984 1550 -2984 0 feedthrough
rlabel pdiffusion 1557 -2984 1557 -2984 0 feedthrough
rlabel pdiffusion 1564 -2984 1564 -2984 0 feedthrough
rlabel pdiffusion 1571 -2984 1571 -2984 0 cellNo=502
rlabel pdiffusion 1578 -2984 1578 -2984 0 feedthrough
rlabel pdiffusion 1585 -2984 1585 -2984 0 feedthrough
rlabel pdiffusion 1592 -2984 1592 -2984 0 feedthrough
rlabel pdiffusion 1599 -2984 1599 -2984 0 feedthrough
rlabel pdiffusion 1606 -2984 1606 -2984 0 feedthrough
rlabel pdiffusion 1613 -2984 1613 -2984 0 feedthrough
rlabel pdiffusion 1620 -2984 1620 -2984 0 feedthrough
rlabel pdiffusion 1627 -2984 1627 -2984 0 feedthrough
rlabel pdiffusion 1634 -2984 1634 -2984 0 feedthrough
rlabel pdiffusion 1641 -2984 1641 -2984 0 feedthrough
rlabel pdiffusion 1648 -2984 1648 -2984 0 feedthrough
rlabel pdiffusion 1655 -2984 1655 -2984 0 feedthrough
rlabel pdiffusion 1662 -2984 1662 -2984 0 feedthrough
rlabel pdiffusion 1669 -2984 1669 -2984 0 feedthrough
rlabel pdiffusion 1676 -2984 1676 -2984 0 feedthrough
rlabel pdiffusion 1683 -2984 1683 -2984 0 feedthrough
rlabel pdiffusion 1690 -2984 1690 -2984 0 feedthrough
rlabel pdiffusion 1697 -2984 1697 -2984 0 feedthrough
rlabel pdiffusion 1704 -2984 1704 -2984 0 feedthrough
rlabel pdiffusion 1711 -2984 1711 -2984 0 feedthrough
rlabel pdiffusion 1718 -2984 1718 -2984 0 feedthrough
rlabel pdiffusion 1725 -2984 1725 -2984 0 feedthrough
rlabel pdiffusion 1732 -2984 1732 -2984 0 feedthrough
rlabel pdiffusion 1739 -2984 1739 -2984 0 feedthrough
rlabel pdiffusion 1746 -2984 1746 -2984 0 feedthrough
rlabel pdiffusion 1753 -2984 1753 -2984 0 feedthrough
rlabel pdiffusion 1760 -2984 1760 -2984 0 feedthrough
rlabel pdiffusion 1767 -2984 1767 -2984 0 cellNo=235
rlabel pdiffusion 1774 -2984 1774 -2984 0 feedthrough
rlabel pdiffusion 1781 -2984 1781 -2984 0 feedthrough
rlabel pdiffusion 1788 -2984 1788 -2984 0 feedthrough
rlabel pdiffusion 1795 -2984 1795 -2984 0 feedthrough
rlabel pdiffusion 1802 -2984 1802 -2984 0 feedthrough
rlabel pdiffusion 1809 -2984 1809 -2984 0 feedthrough
rlabel pdiffusion 1816 -2984 1816 -2984 0 feedthrough
rlabel pdiffusion 1823 -2984 1823 -2984 0 feedthrough
rlabel pdiffusion 1830 -2984 1830 -2984 0 feedthrough
rlabel pdiffusion 1837 -2984 1837 -2984 0 feedthrough
rlabel pdiffusion 1844 -2984 1844 -2984 0 feedthrough
rlabel pdiffusion 1851 -2984 1851 -2984 0 feedthrough
rlabel pdiffusion 1858 -2984 1858 -2984 0 feedthrough
rlabel pdiffusion 1865 -2984 1865 -2984 0 feedthrough
rlabel pdiffusion 1872 -2984 1872 -2984 0 feedthrough
rlabel pdiffusion 1879 -2984 1879 -2984 0 feedthrough
rlabel pdiffusion 1886 -2984 1886 -2984 0 feedthrough
rlabel pdiffusion 1893 -2984 1893 -2984 0 feedthrough
rlabel pdiffusion 1900 -2984 1900 -2984 0 feedthrough
rlabel pdiffusion 1907 -2984 1907 -2984 0 feedthrough
rlabel pdiffusion 1914 -2984 1914 -2984 0 feedthrough
rlabel pdiffusion 1921 -2984 1921 -2984 0 feedthrough
rlabel pdiffusion 1928 -2984 1928 -2984 0 feedthrough
rlabel pdiffusion 1935 -2984 1935 -2984 0 feedthrough
rlabel pdiffusion 1942 -2984 1942 -2984 0 feedthrough
rlabel pdiffusion 1949 -2984 1949 -2984 0 feedthrough
rlabel pdiffusion 1956 -2984 1956 -2984 0 feedthrough
rlabel pdiffusion 1963 -2984 1963 -2984 0 feedthrough
rlabel pdiffusion 1970 -2984 1970 -2984 0 feedthrough
rlabel pdiffusion 1977 -2984 1977 -2984 0 feedthrough
rlabel pdiffusion 1984 -2984 1984 -2984 0 feedthrough
rlabel pdiffusion 1991 -2984 1991 -2984 0 feedthrough
rlabel pdiffusion 1998 -2984 1998 -2984 0 feedthrough
rlabel pdiffusion 2005 -2984 2005 -2984 0 feedthrough
rlabel pdiffusion 2012 -2984 2012 -2984 0 feedthrough
rlabel pdiffusion 2019 -2984 2019 -2984 0 feedthrough
rlabel pdiffusion 2026 -2984 2026 -2984 0 feedthrough
rlabel pdiffusion 2033 -2984 2033 -2984 0 feedthrough
rlabel pdiffusion 2040 -2984 2040 -2984 0 feedthrough
rlabel pdiffusion 2047 -2984 2047 -2984 0 feedthrough
rlabel pdiffusion 2054 -2984 2054 -2984 0 feedthrough
rlabel pdiffusion 2061 -2984 2061 -2984 0 feedthrough
rlabel pdiffusion 2068 -2984 2068 -2984 0 feedthrough
rlabel pdiffusion 2075 -2984 2075 -2984 0 feedthrough
rlabel pdiffusion 2082 -2984 2082 -2984 0 feedthrough
rlabel pdiffusion 2089 -2984 2089 -2984 0 feedthrough
rlabel pdiffusion 2096 -2984 2096 -2984 0 cellNo=177
rlabel pdiffusion 2103 -2984 2103 -2984 0 feedthrough
rlabel pdiffusion 2110 -2984 2110 -2984 0 feedthrough
rlabel pdiffusion 2117 -2984 2117 -2984 0 feedthrough
rlabel pdiffusion 2124 -2984 2124 -2984 0 feedthrough
rlabel pdiffusion 2131 -2984 2131 -2984 0 feedthrough
rlabel pdiffusion 2138 -2984 2138 -2984 0 feedthrough
rlabel pdiffusion 2145 -2984 2145 -2984 0 feedthrough
rlabel pdiffusion 2152 -2984 2152 -2984 0 feedthrough
rlabel pdiffusion 3 -3099 3 -3099 0 cellNo=1004
rlabel pdiffusion 10 -3099 10 -3099 0 cellNo=1038
rlabel pdiffusion 17 -3099 17 -3099 0 cellNo=1048
rlabel pdiffusion 24 -3099 24 -3099 0 feedthrough
rlabel pdiffusion 31 -3099 31 -3099 0 feedthrough
rlabel pdiffusion 38 -3099 38 -3099 0 feedthrough
rlabel pdiffusion 45 -3099 45 -3099 0 cellNo=1086
rlabel pdiffusion 52 -3099 52 -3099 0 cellNo=1076
rlabel pdiffusion 59 -3099 59 -3099 0 feedthrough
rlabel pdiffusion 66 -3099 66 -3099 0 feedthrough
rlabel pdiffusion 73 -3099 73 -3099 0 feedthrough
rlabel pdiffusion 80 -3099 80 -3099 0 cellNo=574
rlabel pdiffusion 87 -3099 87 -3099 0 feedthrough
rlabel pdiffusion 94 -3099 94 -3099 0 cellNo=52
rlabel pdiffusion 101 -3099 101 -3099 0 feedthrough
rlabel pdiffusion 108 -3099 108 -3099 0 feedthrough
rlabel pdiffusion 115 -3099 115 -3099 0 feedthrough
rlabel pdiffusion 122 -3099 122 -3099 0 feedthrough
rlabel pdiffusion 129 -3099 129 -3099 0 cellNo=559
rlabel pdiffusion 136 -3099 136 -3099 0 cellNo=381
rlabel pdiffusion 143 -3099 143 -3099 0 feedthrough
rlabel pdiffusion 150 -3099 150 -3099 0 feedthrough
rlabel pdiffusion 157 -3099 157 -3099 0 feedthrough
rlabel pdiffusion 164 -3099 164 -3099 0 cellNo=977
rlabel pdiffusion 171 -3099 171 -3099 0 cellNo=244
rlabel pdiffusion 178 -3099 178 -3099 0 feedthrough
rlabel pdiffusion 185 -3099 185 -3099 0 feedthrough
rlabel pdiffusion 192 -3099 192 -3099 0 feedthrough
rlabel pdiffusion 199 -3099 199 -3099 0 feedthrough
rlabel pdiffusion 206 -3099 206 -3099 0 cellNo=407
rlabel pdiffusion 213 -3099 213 -3099 0 feedthrough
rlabel pdiffusion 220 -3099 220 -3099 0 feedthrough
rlabel pdiffusion 227 -3099 227 -3099 0 feedthrough
rlabel pdiffusion 234 -3099 234 -3099 0 cellNo=967
rlabel pdiffusion 241 -3099 241 -3099 0 feedthrough
rlabel pdiffusion 248 -3099 248 -3099 0 feedthrough
rlabel pdiffusion 255 -3099 255 -3099 0 feedthrough
rlabel pdiffusion 262 -3099 262 -3099 0 feedthrough
rlabel pdiffusion 269 -3099 269 -3099 0 feedthrough
rlabel pdiffusion 276 -3099 276 -3099 0 feedthrough
rlabel pdiffusion 283 -3099 283 -3099 0 feedthrough
rlabel pdiffusion 290 -3099 290 -3099 0 feedthrough
rlabel pdiffusion 297 -3099 297 -3099 0 feedthrough
rlabel pdiffusion 304 -3099 304 -3099 0 feedthrough
rlabel pdiffusion 311 -3099 311 -3099 0 feedthrough
rlabel pdiffusion 318 -3099 318 -3099 0 feedthrough
rlabel pdiffusion 325 -3099 325 -3099 0 feedthrough
rlabel pdiffusion 332 -3099 332 -3099 0 feedthrough
rlabel pdiffusion 339 -3099 339 -3099 0 feedthrough
rlabel pdiffusion 346 -3099 346 -3099 0 feedthrough
rlabel pdiffusion 353 -3099 353 -3099 0 feedthrough
rlabel pdiffusion 360 -3099 360 -3099 0 feedthrough
rlabel pdiffusion 367 -3099 367 -3099 0 feedthrough
rlabel pdiffusion 374 -3099 374 -3099 0 feedthrough
rlabel pdiffusion 381 -3099 381 -3099 0 feedthrough
rlabel pdiffusion 388 -3099 388 -3099 0 feedthrough
rlabel pdiffusion 395 -3099 395 -3099 0 feedthrough
rlabel pdiffusion 402 -3099 402 -3099 0 feedthrough
rlabel pdiffusion 409 -3099 409 -3099 0 feedthrough
rlabel pdiffusion 416 -3099 416 -3099 0 feedthrough
rlabel pdiffusion 423 -3099 423 -3099 0 feedthrough
rlabel pdiffusion 430 -3099 430 -3099 0 feedthrough
rlabel pdiffusion 437 -3099 437 -3099 0 feedthrough
rlabel pdiffusion 444 -3099 444 -3099 0 feedthrough
rlabel pdiffusion 451 -3099 451 -3099 0 feedthrough
rlabel pdiffusion 458 -3099 458 -3099 0 cellNo=715
rlabel pdiffusion 465 -3099 465 -3099 0 feedthrough
rlabel pdiffusion 472 -3099 472 -3099 0 feedthrough
rlabel pdiffusion 479 -3099 479 -3099 0 feedthrough
rlabel pdiffusion 486 -3099 486 -3099 0 feedthrough
rlabel pdiffusion 493 -3099 493 -3099 0 feedthrough
rlabel pdiffusion 500 -3099 500 -3099 0 feedthrough
rlabel pdiffusion 507 -3099 507 -3099 0 feedthrough
rlabel pdiffusion 514 -3099 514 -3099 0 feedthrough
rlabel pdiffusion 521 -3099 521 -3099 0 feedthrough
rlabel pdiffusion 528 -3099 528 -3099 0 cellNo=642
rlabel pdiffusion 535 -3099 535 -3099 0 feedthrough
rlabel pdiffusion 542 -3099 542 -3099 0 feedthrough
rlabel pdiffusion 549 -3099 549 -3099 0 feedthrough
rlabel pdiffusion 556 -3099 556 -3099 0 feedthrough
rlabel pdiffusion 563 -3099 563 -3099 0 feedthrough
rlabel pdiffusion 570 -3099 570 -3099 0 feedthrough
rlabel pdiffusion 577 -3099 577 -3099 0 feedthrough
rlabel pdiffusion 584 -3099 584 -3099 0 feedthrough
rlabel pdiffusion 591 -3099 591 -3099 0 feedthrough
rlabel pdiffusion 598 -3099 598 -3099 0 feedthrough
rlabel pdiffusion 605 -3099 605 -3099 0 feedthrough
rlabel pdiffusion 612 -3099 612 -3099 0 cellNo=346
rlabel pdiffusion 619 -3099 619 -3099 0 feedthrough
rlabel pdiffusion 626 -3099 626 -3099 0 feedthrough
rlabel pdiffusion 633 -3099 633 -3099 0 feedthrough
rlabel pdiffusion 640 -3099 640 -3099 0 feedthrough
rlabel pdiffusion 647 -3099 647 -3099 0 feedthrough
rlabel pdiffusion 654 -3099 654 -3099 0 feedthrough
rlabel pdiffusion 661 -3099 661 -3099 0 feedthrough
rlabel pdiffusion 668 -3099 668 -3099 0 feedthrough
rlabel pdiffusion 675 -3099 675 -3099 0 feedthrough
rlabel pdiffusion 682 -3099 682 -3099 0 feedthrough
rlabel pdiffusion 689 -3099 689 -3099 0 feedthrough
rlabel pdiffusion 696 -3099 696 -3099 0 feedthrough
rlabel pdiffusion 703 -3099 703 -3099 0 feedthrough
rlabel pdiffusion 710 -3099 710 -3099 0 feedthrough
rlabel pdiffusion 717 -3099 717 -3099 0 feedthrough
rlabel pdiffusion 724 -3099 724 -3099 0 feedthrough
rlabel pdiffusion 731 -3099 731 -3099 0 feedthrough
rlabel pdiffusion 738 -3099 738 -3099 0 feedthrough
rlabel pdiffusion 745 -3099 745 -3099 0 feedthrough
rlabel pdiffusion 752 -3099 752 -3099 0 feedthrough
rlabel pdiffusion 759 -3099 759 -3099 0 feedthrough
rlabel pdiffusion 766 -3099 766 -3099 0 feedthrough
rlabel pdiffusion 773 -3099 773 -3099 0 feedthrough
rlabel pdiffusion 780 -3099 780 -3099 0 feedthrough
rlabel pdiffusion 787 -3099 787 -3099 0 feedthrough
rlabel pdiffusion 794 -3099 794 -3099 0 feedthrough
rlabel pdiffusion 801 -3099 801 -3099 0 feedthrough
rlabel pdiffusion 808 -3099 808 -3099 0 feedthrough
rlabel pdiffusion 815 -3099 815 -3099 0 cellNo=777
rlabel pdiffusion 822 -3099 822 -3099 0 feedthrough
rlabel pdiffusion 829 -3099 829 -3099 0 feedthrough
rlabel pdiffusion 836 -3099 836 -3099 0 feedthrough
rlabel pdiffusion 843 -3099 843 -3099 0 feedthrough
rlabel pdiffusion 850 -3099 850 -3099 0 feedthrough
rlabel pdiffusion 857 -3099 857 -3099 0 feedthrough
rlabel pdiffusion 864 -3099 864 -3099 0 cellNo=391
rlabel pdiffusion 871 -3099 871 -3099 0 feedthrough
rlabel pdiffusion 878 -3099 878 -3099 0 cellNo=844
rlabel pdiffusion 885 -3099 885 -3099 0 feedthrough
rlabel pdiffusion 892 -3099 892 -3099 0 cellNo=257
rlabel pdiffusion 899 -3099 899 -3099 0 feedthrough
rlabel pdiffusion 906 -3099 906 -3099 0 feedthrough
rlabel pdiffusion 913 -3099 913 -3099 0 cellNo=813
rlabel pdiffusion 920 -3099 920 -3099 0 feedthrough
rlabel pdiffusion 927 -3099 927 -3099 0 feedthrough
rlabel pdiffusion 934 -3099 934 -3099 0 feedthrough
rlabel pdiffusion 941 -3099 941 -3099 0 feedthrough
rlabel pdiffusion 948 -3099 948 -3099 0 feedthrough
rlabel pdiffusion 955 -3099 955 -3099 0 feedthrough
rlabel pdiffusion 962 -3099 962 -3099 0 feedthrough
rlabel pdiffusion 969 -3099 969 -3099 0 feedthrough
rlabel pdiffusion 976 -3099 976 -3099 0 feedthrough
rlabel pdiffusion 983 -3099 983 -3099 0 feedthrough
rlabel pdiffusion 990 -3099 990 -3099 0 feedthrough
rlabel pdiffusion 997 -3099 997 -3099 0 feedthrough
rlabel pdiffusion 1004 -3099 1004 -3099 0 feedthrough
rlabel pdiffusion 1011 -3099 1011 -3099 0 feedthrough
rlabel pdiffusion 1018 -3099 1018 -3099 0 feedthrough
rlabel pdiffusion 1025 -3099 1025 -3099 0 feedthrough
rlabel pdiffusion 1032 -3099 1032 -3099 0 feedthrough
rlabel pdiffusion 1039 -3099 1039 -3099 0 feedthrough
rlabel pdiffusion 1046 -3099 1046 -3099 0 feedthrough
rlabel pdiffusion 1053 -3099 1053 -3099 0 cellNo=788
rlabel pdiffusion 1060 -3099 1060 -3099 0 feedthrough
rlabel pdiffusion 1067 -3099 1067 -3099 0 feedthrough
rlabel pdiffusion 1074 -3099 1074 -3099 0 cellNo=557
rlabel pdiffusion 1081 -3099 1081 -3099 0 cellNo=136
rlabel pdiffusion 1088 -3099 1088 -3099 0 feedthrough
rlabel pdiffusion 1095 -3099 1095 -3099 0 feedthrough
rlabel pdiffusion 1102 -3099 1102 -3099 0 feedthrough
rlabel pdiffusion 1109 -3099 1109 -3099 0 feedthrough
rlabel pdiffusion 1116 -3099 1116 -3099 0 feedthrough
rlabel pdiffusion 1123 -3099 1123 -3099 0 cellNo=197
rlabel pdiffusion 1130 -3099 1130 -3099 0 feedthrough
rlabel pdiffusion 1137 -3099 1137 -3099 0 feedthrough
rlabel pdiffusion 1144 -3099 1144 -3099 0 feedthrough
rlabel pdiffusion 1151 -3099 1151 -3099 0 feedthrough
rlabel pdiffusion 1158 -3099 1158 -3099 0 cellNo=267
rlabel pdiffusion 1165 -3099 1165 -3099 0 feedthrough
rlabel pdiffusion 1172 -3099 1172 -3099 0 feedthrough
rlabel pdiffusion 1179 -3099 1179 -3099 0 feedthrough
rlabel pdiffusion 1186 -3099 1186 -3099 0 feedthrough
rlabel pdiffusion 1193 -3099 1193 -3099 0 feedthrough
rlabel pdiffusion 1200 -3099 1200 -3099 0 feedthrough
rlabel pdiffusion 1207 -3099 1207 -3099 0 feedthrough
rlabel pdiffusion 1214 -3099 1214 -3099 0 cellNo=954
rlabel pdiffusion 1221 -3099 1221 -3099 0 feedthrough
rlabel pdiffusion 1228 -3099 1228 -3099 0 feedthrough
rlabel pdiffusion 1235 -3099 1235 -3099 0 cellNo=261
rlabel pdiffusion 1242 -3099 1242 -3099 0 feedthrough
rlabel pdiffusion 1249 -3099 1249 -3099 0 cellNo=393
rlabel pdiffusion 1256 -3099 1256 -3099 0 feedthrough
rlabel pdiffusion 1263 -3099 1263 -3099 0 feedthrough
rlabel pdiffusion 1270 -3099 1270 -3099 0 feedthrough
rlabel pdiffusion 1277 -3099 1277 -3099 0 cellNo=969
rlabel pdiffusion 1284 -3099 1284 -3099 0 feedthrough
rlabel pdiffusion 1291 -3099 1291 -3099 0 feedthrough
rlabel pdiffusion 1298 -3099 1298 -3099 0 feedthrough
rlabel pdiffusion 1305 -3099 1305 -3099 0 feedthrough
rlabel pdiffusion 1312 -3099 1312 -3099 0 cellNo=584
rlabel pdiffusion 1319 -3099 1319 -3099 0 feedthrough
rlabel pdiffusion 1326 -3099 1326 -3099 0 feedthrough
rlabel pdiffusion 1333 -3099 1333 -3099 0 feedthrough
rlabel pdiffusion 1340 -3099 1340 -3099 0 feedthrough
rlabel pdiffusion 1347 -3099 1347 -3099 0 feedthrough
rlabel pdiffusion 1354 -3099 1354 -3099 0 feedthrough
rlabel pdiffusion 1361 -3099 1361 -3099 0 feedthrough
rlabel pdiffusion 1368 -3099 1368 -3099 0 feedthrough
rlabel pdiffusion 1375 -3099 1375 -3099 0 feedthrough
rlabel pdiffusion 1382 -3099 1382 -3099 0 feedthrough
rlabel pdiffusion 1389 -3099 1389 -3099 0 feedthrough
rlabel pdiffusion 1396 -3099 1396 -3099 0 cellNo=375
rlabel pdiffusion 1403 -3099 1403 -3099 0 cellNo=224
rlabel pdiffusion 1410 -3099 1410 -3099 0 feedthrough
rlabel pdiffusion 1417 -3099 1417 -3099 0 feedthrough
rlabel pdiffusion 1424 -3099 1424 -3099 0 feedthrough
rlabel pdiffusion 1431 -3099 1431 -3099 0 feedthrough
rlabel pdiffusion 1438 -3099 1438 -3099 0 feedthrough
rlabel pdiffusion 1445 -3099 1445 -3099 0 cellNo=894
rlabel pdiffusion 1452 -3099 1452 -3099 0 feedthrough
rlabel pdiffusion 1459 -3099 1459 -3099 0 feedthrough
rlabel pdiffusion 1466 -3099 1466 -3099 0 feedthrough
rlabel pdiffusion 1473 -3099 1473 -3099 0 feedthrough
rlabel pdiffusion 1480 -3099 1480 -3099 0 feedthrough
rlabel pdiffusion 1487 -3099 1487 -3099 0 feedthrough
rlabel pdiffusion 1494 -3099 1494 -3099 0 feedthrough
rlabel pdiffusion 1501 -3099 1501 -3099 0 feedthrough
rlabel pdiffusion 1508 -3099 1508 -3099 0 feedthrough
rlabel pdiffusion 1515 -3099 1515 -3099 0 feedthrough
rlabel pdiffusion 1522 -3099 1522 -3099 0 feedthrough
rlabel pdiffusion 1529 -3099 1529 -3099 0 feedthrough
rlabel pdiffusion 1536 -3099 1536 -3099 0 feedthrough
rlabel pdiffusion 1543 -3099 1543 -3099 0 feedthrough
rlabel pdiffusion 1550 -3099 1550 -3099 0 feedthrough
rlabel pdiffusion 1557 -3099 1557 -3099 0 cellNo=456
rlabel pdiffusion 1564 -3099 1564 -3099 0 cellNo=152
rlabel pdiffusion 1571 -3099 1571 -3099 0 feedthrough
rlabel pdiffusion 1578 -3099 1578 -3099 0 feedthrough
rlabel pdiffusion 1585 -3099 1585 -3099 0 feedthrough
rlabel pdiffusion 1592 -3099 1592 -3099 0 feedthrough
rlabel pdiffusion 1599 -3099 1599 -3099 0 feedthrough
rlabel pdiffusion 1606 -3099 1606 -3099 0 feedthrough
rlabel pdiffusion 1613 -3099 1613 -3099 0 feedthrough
rlabel pdiffusion 1620 -3099 1620 -3099 0 feedthrough
rlabel pdiffusion 1627 -3099 1627 -3099 0 feedthrough
rlabel pdiffusion 1634 -3099 1634 -3099 0 feedthrough
rlabel pdiffusion 1641 -3099 1641 -3099 0 feedthrough
rlabel pdiffusion 1648 -3099 1648 -3099 0 feedthrough
rlabel pdiffusion 1655 -3099 1655 -3099 0 feedthrough
rlabel pdiffusion 1662 -3099 1662 -3099 0 feedthrough
rlabel pdiffusion 1669 -3099 1669 -3099 0 feedthrough
rlabel pdiffusion 1676 -3099 1676 -3099 0 feedthrough
rlabel pdiffusion 1683 -3099 1683 -3099 0 cellNo=503
rlabel pdiffusion 1690 -3099 1690 -3099 0 feedthrough
rlabel pdiffusion 1697 -3099 1697 -3099 0 feedthrough
rlabel pdiffusion 1704 -3099 1704 -3099 0 feedthrough
rlabel pdiffusion 1711 -3099 1711 -3099 0 feedthrough
rlabel pdiffusion 1718 -3099 1718 -3099 0 feedthrough
rlabel pdiffusion 1725 -3099 1725 -3099 0 feedthrough
rlabel pdiffusion 1732 -3099 1732 -3099 0 feedthrough
rlabel pdiffusion 1739 -3099 1739 -3099 0 feedthrough
rlabel pdiffusion 1746 -3099 1746 -3099 0 feedthrough
rlabel pdiffusion 1753 -3099 1753 -3099 0 feedthrough
rlabel pdiffusion 1760 -3099 1760 -3099 0 feedthrough
rlabel pdiffusion 1767 -3099 1767 -3099 0 feedthrough
rlabel pdiffusion 1774 -3099 1774 -3099 0 feedthrough
rlabel pdiffusion 1781 -3099 1781 -3099 0 feedthrough
rlabel pdiffusion 1788 -3099 1788 -3099 0 feedthrough
rlabel pdiffusion 1795 -3099 1795 -3099 0 feedthrough
rlabel pdiffusion 1802 -3099 1802 -3099 0 feedthrough
rlabel pdiffusion 1809 -3099 1809 -3099 0 feedthrough
rlabel pdiffusion 1816 -3099 1816 -3099 0 feedthrough
rlabel pdiffusion 1823 -3099 1823 -3099 0 feedthrough
rlabel pdiffusion 1830 -3099 1830 -3099 0 feedthrough
rlabel pdiffusion 1837 -3099 1837 -3099 0 feedthrough
rlabel pdiffusion 1844 -3099 1844 -3099 0 feedthrough
rlabel pdiffusion 1851 -3099 1851 -3099 0 feedthrough
rlabel pdiffusion 1858 -3099 1858 -3099 0 feedthrough
rlabel pdiffusion 1865 -3099 1865 -3099 0 feedthrough
rlabel pdiffusion 1872 -3099 1872 -3099 0 feedthrough
rlabel pdiffusion 1879 -3099 1879 -3099 0 cellNo=96
rlabel pdiffusion 1886 -3099 1886 -3099 0 feedthrough
rlabel pdiffusion 1893 -3099 1893 -3099 0 feedthrough
rlabel pdiffusion 1900 -3099 1900 -3099 0 feedthrough
rlabel pdiffusion 1907 -3099 1907 -3099 0 feedthrough
rlabel pdiffusion 1914 -3099 1914 -3099 0 feedthrough
rlabel pdiffusion 1921 -3099 1921 -3099 0 feedthrough
rlabel pdiffusion 1928 -3099 1928 -3099 0 feedthrough
rlabel pdiffusion 1935 -3099 1935 -3099 0 feedthrough
rlabel pdiffusion 1942 -3099 1942 -3099 0 feedthrough
rlabel pdiffusion 1949 -3099 1949 -3099 0 feedthrough
rlabel pdiffusion 1956 -3099 1956 -3099 0 feedthrough
rlabel pdiffusion 1963 -3099 1963 -3099 0 cellNo=922
rlabel pdiffusion 1970 -3099 1970 -3099 0 feedthrough
rlabel pdiffusion 1977 -3099 1977 -3099 0 feedthrough
rlabel pdiffusion 1984 -3099 1984 -3099 0 feedthrough
rlabel pdiffusion 1991 -3099 1991 -3099 0 feedthrough
rlabel pdiffusion 1998 -3099 1998 -3099 0 feedthrough
rlabel pdiffusion 2005 -3099 2005 -3099 0 feedthrough
rlabel pdiffusion 2033 -3099 2033 -3099 0 feedthrough
rlabel pdiffusion 2047 -3099 2047 -3099 0 feedthrough
rlabel pdiffusion 2075 -3099 2075 -3099 0 feedthrough
rlabel pdiffusion 3 -3230 3 -3230 0 cellNo=1039
rlabel pdiffusion 10 -3230 10 -3230 0 cellNo=1351
rlabel pdiffusion 17 -3230 17 -3230 0 cellNo=1069
rlabel pdiffusion 94 -3230 94 -3230 0 feedthrough
rlabel pdiffusion 101 -3230 101 -3230 0 feedthrough
rlabel pdiffusion 108 -3230 108 -3230 0 feedthrough
rlabel pdiffusion 115 -3230 115 -3230 0 cellNo=863
rlabel pdiffusion 122 -3230 122 -3230 0 feedthrough
rlabel pdiffusion 129 -3230 129 -3230 0 feedthrough
rlabel pdiffusion 136 -3230 136 -3230 0 feedthrough
rlabel pdiffusion 143 -3230 143 -3230 0 feedthrough
rlabel pdiffusion 150 -3230 150 -3230 0 feedthrough
rlabel pdiffusion 157 -3230 157 -3230 0 feedthrough
rlabel pdiffusion 164 -3230 164 -3230 0 feedthrough
rlabel pdiffusion 171 -3230 171 -3230 0 cellNo=836
rlabel pdiffusion 178 -3230 178 -3230 0 feedthrough
rlabel pdiffusion 185 -3230 185 -3230 0 cellNo=755
rlabel pdiffusion 192 -3230 192 -3230 0 cellNo=589
rlabel pdiffusion 199 -3230 199 -3230 0 feedthrough
rlabel pdiffusion 206 -3230 206 -3230 0 cellNo=976
rlabel pdiffusion 213 -3230 213 -3230 0 feedthrough
rlabel pdiffusion 220 -3230 220 -3230 0 feedthrough
rlabel pdiffusion 227 -3230 227 -3230 0 feedthrough
rlabel pdiffusion 234 -3230 234 -3230 0 feedthrough
rlabel pdiffusion 241 -3230 241 -3230 0 feedthrough
rlabel pdiffusion 248 -3230 248 -3230 0 feedthrough
rlabel pdiffusion 255 -3230 255 -3230 0 feedthrough
rlabel pdiffusion 262 -3230 262 -3230 0 feedthrough
rlabel pdiffusion 269 -3230 269 -3230 0 feedthrough
rlabel pdiffusion 276 -3230 276 -3230 0 feedthrough
rlabel pdiffusion 283 -3230 283 -3230 0 feedthrough
rlabel pdiffusion 290 -3230 290 -3230 0 feedthrough
rlabel pdiffusion 297 -3230 297 -3230 0 feedthrough
rlabel pdiffusion 304 -3230 304 -3230 0 feedthrough
rlabel pdiffusion 311 -3230 311 -3230 0 feedthrough
rlabel pdiffusion 318 -3230 318 -3230 0 feedthrough
rlabel pdiffusion 325 -3230 325 -3230 0 feedthrough
rlabel pdiffusion 332 -3230 332 -3230 0 feedthrough
rlabel pdiffusion 339 -3230 339 -3230 0 feedthrough
rlabel pdiffusion 346 -3230 346 -3230 0 feedthrough
rlabel pdiffusion 353 -3230 353 -3230 0 feedthrough
rlabel pdiffusion 360 -3230 360 -3230 0 feedthrough
rlabel pdiffusion 367 -3230 367 -3230 0 feedthrough
rlabel pdiffusion 374 -3230 374 -3230 0 feedthrough
rlabel pdiffusion 381 -3230 381 -3230 0 feedthrough
rlabel pdiffusion 388 -3230 388 -3230 0 feedthrough
rlabel pdiffusion 395 -3230 395 -3230 0 feedthrough
rlabel pdiffusion 402 -3230 402 -3230 0 cellNo=572
rlabel pdiffusion 409 -3230 409 -3230 0 feedthrough
rlabel pdiffusion 416 -3230 416 -3230 0 cellNo=293
rlabel pdiffusion 423 -3230 423 -3230 0 cellNo=412
rlabel pdiffusion 430 -3230 430 -3230 0 feedthrough
rlabel pdiffusion 437 -3230 437 -3230 0 feedthrough
rlabel pdiffusion 444 -3230 444 -3230 0 feedthrough
rlabel pdiffusion 451 -3230 451 -3230 0 feedthrough
rlabel pdiffusion 458 -3230 458 -3230 0 feedthrough
rlabel pdiffusion 465 -3230 465 -3230 0 feedthrough
rlabel pdiffusion 472 -3230 472 -3230 0 feedthrough
rlabel pdiffusion 479 -3230 479 -3230 0 feedthrough
rlabel pdiffusion 486 -3230 486 -3230 0 feedthrough
rlabel pdiffusion 493 -3230 493 -3230 0 cellNo=617
rlabel pdiffusion 500 -3230 500 -3230 0 feedthrough
rlabel pdiffusion 507 -3230 507 -3230 0 feedthrough
rlabel pdiffusion 514 -3230 514 -3230 0 feedthrough
rlabel pdiffusion 521 -3230 521 -3230 0 feedthrough
rlabel pdiffusion 528 -3230 528 -3230 0 feedthrough
rlabel pdiffusion 535 -3230 535 -3230 0 feedthrough
rlabel pdiffusion 542 -3230 542 -3230 0 feedthrough
rlabel pdiffusion 549 -3230 549 -3230 0 feedthrough
rlabel pdiffusion 556 -3230 556 -3230 0 feedthrough
rlabel pdiffusion 563 -3230 563 -3230 0 feedthrough
rlabel pdiffusion 570 -3230 570 -3230 0 feedthrough
rlabel pdiffusion 577 -3230 577 -3230 0 cellNo=537
rlabel pdiffusion 584 -3230 584 -3230 0 feedthrough
rlabel pdiffusion 591 -3230 591 -3230 0 feedthrough
rlabel pdiffusion 598 -3230 598 -3230 0 feedthrough
rlabel pdiffusion 605 -3230 605 -3230 0 feedthrough
rlabel pdiffusion 612 -3230 612 -3230 0 cellNo=939
rlabel pdiffusion 619 -3230 619 -3230 0 feedthrough
rlabel pdiffusion 626 -3230 626 -3230 0 feedthrough
rlabel pdiffusion 633 -3230 633 -3230 0 feedthrough
rlabel pdiffusion 640 -3230 640 -3230 0 feedthrough
rlabel pdiffusion 647 -3230 647 -3230 0 feedthrough
rlabel pdiffusion 654 -3230 654 -3230 0 feedthrough
rlabel pdiffusion 661 -3230 661 -3230 0 feedthrough
rlabel pdiffusion 668 -3230 668 -3230 0 feedthrough
rlabel pdiffusion 675 -3230 675 -3230 0 cellNo=943
rlabel pdiffusion 682 -3230 682 -3230 0 feedthrough
rlabel pdiffusion 689 -3230 689 -3230 0 feedthrough
rlabel pdiffusion 696 -3230 696 -3230 0 feedthrough
rlabel pdiffusion 703 -3230 703 -3230 0 feedthrough
rlabel pdiffusion 710 -3230 710 -3230 0 feedthrough
rlabel pdiffusion 717 -3230 717 -3230 0 cellNo=385
rlabel pdiffusion 724 -3230 724 -3230 0 feedthrough
rlabel pdiffusion 731 -3230 731 -3230 0 feedthrough
rlabel pdiffusion 738 -3230 738 -3230 0 feedthrough
rlabel pdiffusion 745 -3230 745 -3230 0 cellNo=588
rlabel pdiffusion 752 -3230 752 -3230 0 feedthrough
rlabel pdiffusion 759 -3230 759 -3230 0 feedthrough
rlabel pdiffusion 766 -3230 766 -3230 0 cellNo=30
rlabel pdiffusion 773 -3230 773 -3230 0 feedthrough
rlabel pdiffusion 780 -3230 780 -3230 0 feedthrough
rlabel pdiffusion 787 -3230 787 -3230 0 feedthrough
rlabel pdiffusion 794 -3230 794 -3230 0 feedthrough
rlabel pdiffusion 801 -3230 801 -3230 0 cellNo=594
rlabel pdiffusion 808 -3230 808 -3230 0 feedthrough
rlabel pdiffusion 815 -3230 815 -3230 0 cellNo=203
rlabel pdiffusion 822 -3230 822 -3230 0 feedthrough
rlabel pdiffusion 829 -3230 829 -3230 0 feedthrough
rlabel pdiffusion 836 -3230 836 -3230 0 feedthrough
rlabel pdiffusion 843 -3230 843 -3230 0 feedthrough
rlabel pdiffusion 850 -3230 850 -3230 0 feedthrough
rlabel pdiffusion 857 -3230 857 -3230 0 feedthrough
rlabel pdiffusion 864 -3230 864 -3230 0 feedthrough
rlabel pdiffusion 871 -3230 871 -3230 0 cellNo=776
rlabel pdiffusion 878 -3230 878 -3230 0 feedthrough
rlabel pdiffusion 885 -3230 885 -3230 0 feedthrough
rlabel pdiffusion 892 -3230 892 -3230 0 feedthrough
rlabel pdiffusion 899 -3230 899 -3230 0 feedthrough
rlabel pdiffusion 906 -3230 906 -3230 0 feedthrough
rlabel pdiffusion 913 -3230 913 -3230 0 feedthrough
rlabel pdiffusion 920 -3230 920 -3230 0 feedthrough
rlabel pdiffusion 927 -3230 927 -3230 0 feedthrough
rlabel pdiffusion 934 -3230 934 -3230 0 feedthrough
rlabel pdiffusion 941 -3230 941 -3230 0 cellNo=326
rlabel pdiffusion 948 -3230 948 -3230 0 feedthrough
rlabel pdiffusion 955 -3230 955 -3230 0 cellNo=512
rlabel pdiffusion 962 -3230 962 -3230 0 feedthrough
rlabel pdiffusion 969 -3230 969 -3230 0 feedthrough
rlabel pdiffusion 976 -3230 976 -3230 0 feedthrough
rlabel pdiffusion 983 -3230 983 -3230 0 cellNo=880
rlabel pdiffusion 990 -3230 990 -3230 0 feedthrough
rlabel pdiffusion 997 -3230 997 -3230 0 feedthrough
rlabel pdiffusion 1004 -3230 1004 -3230 0 feedthrough
rlabel pdiffusion 1011 -3230 1011 -3230 0 feedthrough
rlabel pdiffusion 1018 -3230 1018 -3230 0 feedthrough
rlabel pdiffusion 1025 -3230 1025 -3230 0 feedthrough
rlabel pdiffusion 1032 -3230 1032 -3230 0 feedthrough
rlabel pdiffusion 1039 -3230 1039 -3230 0 feedthrough
rlabel pdiffusion 1046 -3230 1046 -3230 0 feedthrough
rlabel pdiffusion 1053 -3230 1053 -3230 0 feedthrough
rlabel pdiffusion 1060 -3230 1060 -3230 0 feedthrough
rlabel pdiffusion 1067 -3230 1067 -3230 0 feedthrough
rlabel pdiffusion 1074 -3230 1074 -3230 0 feedthrough
rlabel pdiffusion 1081 -3230 1081 -3230 0 feedthrough
rlabel pdiffusion 1088 -3230 1088 -3230 0 feedthrough
rlabel pdiffusion 1095 -3230 1095 -3230 0 feedthrough
rlabel pdiffusion 1102 -3230 1102 -3230 0 feedthrough
rlabel pdiffusion 1109 -3230 1109 -3230 0 cellNo=644
rlabel pdiffusion 1116 -3230 1116 -3230 0 feedthrough
rlabel pdiffusion 1123 -3230 1123 -3230 0 feedthrough
rlabel pdiffusion 1130 -3230 1130 -3230 0 feedthrough
rlabel pdiffusion 1137 -3230 1137 -3230 0 feedthrough
rlabel pdiffusion 1144 -3230 1144 -3230 0 feedthrough
rlabel pdiffusion 1151 -3230 1151 -3230 0 feedthrough
rlabel pdiffusion 1158 -3230 1158 -3230 0 feedthrough
rlabel pdiffusion 1165 -3230 1165 -3230 0 cellNo=448
rlabel pdiffusion 1172 -3230 1172 -3230 0 feedthrough
rlabel pdiffusion 1179 -3230 1179 -3230 0 feedthrough
rlabel pdiffusion 1186 -3230 1186 -3230 0 feedthrough
rlabel pdiffusion 1193 -3230 1193 -3230 0 feedthrough
rlabel pdiffusion 1200 -3230 1200 -3230 0 feedthrough
rlabel pdiffusion 1207 -3230 1207 -3230 0 feedthrough
rlabel pdiffusion 1214 -3230 1214 -3230 0 cellNo=390
rlabel pdiffusion 1221 -3230 1221 -3230 0 feedthrough
rlabel pdiffusion 1228 -3230 1228 -3230 0 feedthrough
rlabel pdiffusion 1235 -3230 1235 -3230 0 cellNo=845
rlabel pdiffusion 1242 -3230 1242 -3230 0 feedthrough
rlabel pdiffusion 1249 -3230 1249 -3230 0 feedthrough
rlabel pdiffusion 1256 -3230 1256 -3230 0 cellNo=582
rlabel pdiffusion 1263 -3230 1263 -3230 0 feedthrough
rlabel pdiffusion 1270 -3230 1270 -3230 0 feedthrough
rlabel pdiffusion 1277 -3230 1277 -3230 0 feedthrough
rlabel pdiffusion 1284 -3230 1284 -3230 0 feedthrough
rlabel pdiffusion 1291 -3230 1291 -3230 0 feedthrough
rlabel pdiffusion 1298 -3230 1298 -3230 0 feedthrough
rlabel pdiffusion 1305 -3230 1305 -3230 0 feedthrough
rlabel pdiffusion 1312 -3230 1312 -3230 0 feedthrough
rlabel pdiffusion 1319 -3230 1319 -3230 0 feedthrough
rlabel pdiffusion 1326 -3230 1326 -3230 0 feedthrough
rlabel pdiffusion 1333 -3230 1333 -3230 0 feedthrough
rlabel pdiffusion 1340 -3230 1340 -3230 0 feedthrough
rlabel pdiffusion 1347 -3230 1347 -3230 0 feedthrough
rlabel pdiffusion 1354 -3230 1354 -3230 0 cellNo=513
rlabel pdiffusion 1361 -3230 1361 -3230 0 feedthrough
rlabel pdiffusion 1368 -3230 1368 -3230 0 feedthrough
rlabel pdiffusion 1375 -3230 1375 -3230 0 feedthrough
rlabel pdiffusion 1382 -3230 1382 -3230 0 feedthrough
rlabel pdiffusion 1389 -3230 1389 -3230 0 feedthrough
rlabel pdiffusion 1396 -3230 1396 -3230 0 feedthrough
rlabel pdiffusion 1403 -3230 1403 -3230 0 feedthrough
rlabel pdiffusion 1410 -3230 1410 -3230 0 feedthrough
rlabel pdiffusion 1417 -3230 1417 -3230 0 feedthrough
rlabel pdiffusion 1424 -3230 1424 -3230 0 feedthrough
rlabel pdiffusion 1431 -3230 1431 -3230 0 feedthrough
rlabel pdiffusion 1438 -3230 1438 -3230 0 feedthrough
rlabel pdiffusion 1445 -3230 1445 -3230 0 feedthrough
rlabel pdiffusion 1452 -3230 1452 -3230 0 feedthrough
rlabel pdiffusion 1459 -3230 1459 -3230 0 cellNo=901
rlabel pdiffusion 1466 -3230 1466 -3230 0 feedthrough
rlabel pdiffusion 1473 -3230 1473 -3230 0 feedthrough
rlabel pdiffusion 1480 -3230 1480 -3230 0 feedthrough
rlabel pdiffusion 1487 -3230 1487 -3230 0 feedthrough
rlabel pdiffusion 1494 -3230 1494 -3230 0 feedthrough
rlabel pdiffusion 1501 -3230 1501 -3230 0 feedthrough
rlabel pdiffusion 1508 -3230 1508 -3230 0 feedthrough
rlabel pdiffusion 1515 -3230 1515 -3230 0 feedthrough
rlabel pdiffusion 1522 -3230 1522 -3230 0 feedthrough
rlabel pdiffusion 1529 -3230 1529 -3230 0 feedthrough
rlabel pdiffusion 1536 -3230 1536 -3230 0 feedthrough
rlabel pdiffusion 1543 -3230 1543 -3230 0 feedthrough
rlabel pdiffusion 1550 -3230 1550 -3230 0 feedthrough
rlabel pdiffusion 1557 -3230 1557 -3230 0 feedthrough
rlabel pdiffusion 1564 -3230 1564 -3230 0 feedthrough
rlabel pdiffusion 1571 -3230 1571 -3230 0 feedthrough
rlabel pdiffusion 1578 -3230 1578 -3230 0 cellNo=610
rlabel pdiffusion 1585 -3230 1585 -3230 0 feedthrough
rlabel pdiffusion 1592 -3230 1592 -3230 0 feedthrough
rlabel pdiffusion 1599 -3230 1599 -3230 0 feedthrough
rlabel pdiffusion 1606 -3230 1606 -3230 0 feedthrough
rlabel pdiffusion 1613 -3230 1613 -3230 0 feedthrough
rlabel pdiffusion 1620 -3230 1620 -3230 0 feedthrough
rlabel pdiffusion 1627 -3230 1627 -3230 0 feedthrough
rlabel pdiffusion 1634 -3230 1634 -3230 0 feedthrough
rlabel pdiffusion 1641 -3230 1641 -3230 0 cellNo=757
rlabel pdiffusion 1648 -3230 1648 -3230 0 cellNo=90
rlabel pdiffusion 1655 -3230 1655 -3230 0 cellNo=168
rlabel pdiffusion 1662 -3230 1662 -3230 0 feedthrough
rlabel pdiffusion 1669 -3230 1669 -3230 0 cellNo=938
rlabel pdiffusion 1676 -3230 1676 -3230 0 feedthrough
rlabel pdiffusion 1683 -3230 1683 -3230 0 cellNo=442
rlabel pdiffusion 1690 -3230 1690 -3230 0 feedthrough
rlabel pdiffusion 1697 -3230 1697 -3230 0 feedthrough
rlabel pdiffusion 1704 -3230 1704 -3230 0 feedthrough
rlabel pdiffusion 1711 -3230 1711 -3230 0 feedthrough
rlabel pdiffusion 1718 -3230 1718 -3230 0 feedthrough
rlabel pdiffusion 1725 -3230 1725 -3230 0 feedthrough
rlabel pdiffusion 1732 -3230 1732 -3230 0 feedthrough
rlabel pdiffusion 1739 -3230 1739 -3230 0 feedthrough
rlabel pdiffusion 1746 -3230 1746 -3230 0 feedthrough
rlabel pdiffusion 1753 -3230 1753 -3230 0 feedthrough
rlabel pdiffusion 1760 -3230 1760 -3230 0 feedthrough
rlabel pdiffusion 1767 -3230 1767 -3230 0 feedthrough
rlabel pdiffusion 1774 -3230 1774 -3230 0 feedthrough
rlabel pdiffusion 1781 -3230 1781 -3230 0 feedthrough
rlabel pdiffusion 1809 -3230 1809 -3230 0 feedthrough
rlabel pdiffusion 1816 -3230 1816 -3230 0 feedthrough
rlabel pdiffusion 1823 -3230 1823 -3230 0 feedthrough
rlabel pdiffusion 1851 -3230 1851 -3230 0 cellNo=315
rlabel pdiffusion 1858 -3230 1858 -3230 0 feedthrough
rlabel pdiffusion 1865 -3230 1865 -3230 0 feedthrough
rlabel pdiffusion 1879 -3230 1879 -3230 0 feedthrough
rlabel pdiffusion 1886 -3230 1886 -3230 0 feedthrough
rlabel pdiffusion 1893 -3230 1893 -3230 0 feedthrough
rlabel pdiffusion 1907 -3230 1907 -3230 0 feedthrough
rlabel pdiffusion 1921 -3230 1921 -3230 0 feedthrough
rlabel pdiffusion 1963 -3230 1963 -3230 0 cellNo=710
rlabel pdiffusion 1970 -3230 1970 -3230 0 feedthrough
rlabel pdiffusion 1977 -3230 1977 -3230 0 feedthrough
rlabel pdiffusion 1984 -3230 1984 -3230 0 feedthrough
rlabel pdiffusion 2019 -3230 2019 -3230 0 feedthrough
rlabel pdiffusion 2047 -3230 2047 -3230 0 feedthrough
rlabel pdiffusion 3 -3333 3 -3333 0 cellNo=1029
rlabel pdiffusion 10 -3333 10 -3333 0 cellNo=1091
rlabel pdiffusion 17 -3333 17 -3333 0 cellNo=1047
rlabel pdiffusion 24 -3333 24 -3333 0 cellNo=1053
rlabel pdiffusion 31 -3333 31 -3333 0 cellNo=1120
rlabel pdiffusion 38 -3333 38 -3333 0 cellNo=1240
rlabel pdiffusion 143 -3333 143 -3333 0 feedthrough
rlabel pdiffusion 164 -3333 164 -3333 0 feedthrough
rlabel pdiffusion 171 -3333 171 -3333 0 feedthrough
rlabel pdiffusion 178 -3333 178 -3333 0 feedthrough
rlabel pdiffusion 185 -3333 185 -3333 0 feedthrough
rlabel pdiffusion 192 -3333 192 -3333 0 feedthrough
rlabel pdiffusion 199 -3333 199 -3333 0 feedthrough
rlabel pdiffusion 206 -3333 206 -3333 0 feedthrough
rlabel pdiffusion 213 -3333 213 -3333 0 cellNo=853
rlabel pdiffusion 220 -3333 220 -3333 0 feedthrough
rlabel pdiffusion 227 -3333 227 -3333 0 cellNo=246
rlabel pdiffusion 234 -3333 234 -3333 0 cellNo=211
rlabel pdiffusion 241 -3333 241 -3333 0 feedthrough
rlabel pdiffusion 248 -3333 248 -3333 0 feedthrough
rlabel pdiffusion 255 -3333 255 -3333 0 cellNo=892
rlabel pdiffusion 262 -3333 262 -3333 0 feedthrough
rlabel pdiffusion 269 -3333 269 -3333 0 feedthrough
rlabel pdiffusion 276 -3333 276 -3333 0 feedthrough
rlabel pdiffusion 283 -3333 283 -3333 0 feedthrough
rlabel pdiffusion 290 -3333 290 -3333 0 feedthrough
rlabel pdiffusion 297 -3333 297 -3333 0 feedthrough
rlabel pdiffusion 304 -3333 304 -3333 0 feedthrough
rlabel pdiffusion 311 -3333 311 -3333 0 feedthrough
rlabel pdiffusion 318 -3333 318 -3333 0 feedthrough
rlabel pdiffusion 325 -3333 325 -3333 0 feedthrough
rlabel pdiffusion 332 -3333 332 -3333 0 feedthrough
rlabel pdiffusion 339 -3333 339 -3333 0 feedthrough
rlabel pdiffusion 346 -3333 346 -3333 0 feedthrough
rlabel pdiffusion 353 -3333 353 -3333 0 feedthrough
rlabel pdiffusion 360 -3333 360 -3333 0 feedthrough
rlabel pdiffusion 367 -3333 367 -3333 0 feedthrough
rlabel pdiffusion 374 -3333 374 -3333 0 feedthrough
rlabel pdiffusion 381 -3333 381 -3333 0 cellNo=676
rlabel pdiffusion 388 -3333 388 -3333 0 feedthrough
rlabel pdiffusion 395 -3333 395 -3333 0 feedthrough
rlabel pdiffusion 402 -3333 402 -3333 0 feedthrough
rlabel pdiffusion 409 -3333 409 -3333 0 feedthrough
rlabel pdiffusion 416 -3333 416 -3333 0 cellNo=359
rlabel pdiffusion 423 -3333 423 -3333 0 feedthrough
rlabel pdiffusion 430 -3333 430 -3333 0 feedthrough
rlabel pdiffusion 437 -3333 437 -3333 0 feedthrough
rlabel pdiffusion 444 -3333 444 -3333 0 feedthrough
rlabel pdiffusion 451 -3333 451 -3333 0 feedthrough
rlabel pdiffusion 458 -3333 458 -3333 0 feedthrough
rlabel pdiffusion 465 -3333 465 -3333 0 feedthrough
rlabel pdiffusion 472 -3333 472 -3333 0 feedthrough
rlabel pdiffusion 479 -3333 479 -3333 0 feedthrough
rlabel pdiffusion 486 -3333 486 -3333 0 feedthrough
rlabel pdiffusion 493 -3333 493 -3333 0 feedthrough
rlabel pdiffusion 500 -3333 500 -3333 0 feedthrough
rlabel pdiffusion 507 -3333 507 -3333 0 feedthrough
rlabel pdiffusion 514 -3333 514 -3333 0 feedthrough
rlabel pdiffusion 521 -3333 521 -3333 0 feedthrough
rlabel pdiffusion 528 -3333 528 -3333 0 feedthrough
rlabel pdiffusion 535 -3333 535 -3333 0 cellNo=496
rlabel pdiffusion 542 -3333 542 -3333 0 feedthrough
rlabel pdiffusion 549 -3333 549 -3333 0 feedthrough
rlabel pdiffusion 556 -3333 556 -3333 0 feedthrough
rlabel pdiffusion 563 -3333 563 -3333 0 feedthrough
rlabel pdiffusion 570 -3333 570 -3333 0 feedthrough
rlabel pdiffusion 577 -3333 577 -3333 0 feedthrough
rlabel pdiffusion 584 -3333 584 -3333 0 feedthrough
rlabel pdiffusion 591 -3333 591 -3333 0 feedthrough
rlabel pdiffusion 598 -3333 598 -3333 0 cellNo=44
rlabel pdiffusion 605 -3333 605 -3333 0 feedthrough
rlabel pdiffusion 612 -3333 612 -3333 0 feedthrough
rlabel pdiffusion 619 -3333 619 -3333 0 feedthrough
rlabel pdiffusion 626 -3333 626 -3333 0 feedthrough
rlabel pdiffusion 633 -3333 633 -3333 0 feedthrough
rlabel pdiffusion 640 -3333 640 -3333 0 cellNo=789
rlabel pdiffusion 647 -3333 647 -3333 0 feedthrough
rlabel pdiffusion 654 -3333 654 -3333 0 feedthrough
rlabel pdiffusion 661 -3333 661 -3333 0 feedthrough
rlabel pdiffusion 668 -3333 668 -3333 0 feedthrough
rlabel pdiffusion 675 -3333 675 -3333 0 feedthrough
rlabel pdiffusion 682 -3333 682 -3333 0 feedthrough
rlabel pdiffusion 689 -3333 689 -3333 0 feedthrough
rlabel pdiffusion 696 -3333 696 -3333 0 feedthrough
rlabel pdiffusion 703 -3333 703 -3333 0 feedthrough
rlabel pdiffusion 710 -3333 710 -3333 0 feedthrough
rlabel pdiffusion 717 -3333 717 -3333 0 feedthrough
rlabel pdiffusion 724 -3333 724 -3333 0 cellNo=832
rlabel pdiffusion 731 -3333 731 -3333 0 cellNo=942
rlabel pdiffusion 738 -3333 738 -3333 0 feedthrough
rlabel pdiffusion 745 -3333 745 -3333 0 feedthrough
rlabel pdiffusion 752 -3333 752 -3333 0 feedthrough
rlabel pdiffusion 759 -3333 759 -3333 0 feedthrough
rlabel pdiffusion 766 -3333 766 -3333 0 feedthrough
rlabel pdiffusion 773 -3333 773 -3333 0 feedthrough
rlabel pdiffusion 780 -3333 780 -3333 0 cellNo=903
rlabel pdiffusion 787 -3333 787 -3333 0 feedthrough
rlabel pdiffusion 794 -3333 794 -3333 0 feedthrough
rlabel pdiffusion 801 -3333 801 -3333 0 feedthrough
rlabel pdiffusion 808 -3333 808 -3333 0 feedthrough
rlabel pdiffusion 815 -3333 815 -3333 0 feedthrough
rlabel pdiffusion 822 -3333 822 -3333 0 feedthrough
rlabel pdiffusion 829 -3333 829 -3333 0 feedthrough
rlabel pdiffusion 836 -3333 836 -3333 0 feedthrough
rlabel pdiffusion 843 -3333 843 -3333 0 feedthrough
rlabel pdiffusion 850 -3333 850 -3333 0 cellNo=956
rlabel pdiffusion 857 -3333 857 -3333 0 feedthrough
rlabel pdiffusion 864 -3333 864 -3333 0 feedthrough
rlabel pdiffusion 871 -3333 871 -3333 0 feedthrough
rlabel pdiffusion 878 -3333 878 -3333 0 feedthrough
rlabel pdiffusion 885 -3333 885 -3333 0 feedthrough
rlabel pdiffusion 892 -3333 892 -3333 0 feedthrough
rlabel pdiffusion 899 -3333 899 -3333 0 feedthrough
rlabel pdiffusion 906 -3333 906 -3333 0 feedthrough
rlabel pdiffusion 913 -3333 913 -3333 0 feedthrough
rlabel pdiffusion 920 -3333 920 -3333 0 feedthrough
rlabel pdiffusion 927 -3333 927 -3333 0 cellNo=669
rlabel pdiffusion 934 -3333 934 -3333 0 feedthrough
rlabel pdiffusion 941 -3333 941 -3333 0 feedthrough
rlabel pdiffusion 948 -3333 948 -3333 0 feedthrough
rlabel pdiffusion 955 -3333 955 -3333 0 cellNo=238
rlabel pdiffusion 962 -3333 962 -3333 0 feedthrough
rlabel pdiffusion 969 -3333 969 -3333 0 cellNo=697
rlabel pdiffusion 976 -3333 976 -3333 0 cellNo=616
rlabel pdiffusion 983 -3333 983 -3333 0 feedthrough
rlabel pdiffusion 990 -3333 990 -3333 0 cellNo=121
rlabel pdiffusion 997 -3333 997 -3333 0 feedthrough
rlabel pdiffusion 1004 -3333 1004 -3333 0 feedthrough
rlabel pdiffusion 1011 -3333 1011 -3333 0 feedthrough
rlabel pdiffusion 1018 -3333 1018 -3333 0 feedthrough
rlabel pdiffusion 1025 -3333 1025 -3333 0 feedthrough
rlabel pdiffusion 1032 -3333 1032 -3333 0 feedthrough
rlabel pdiffusion 1039 -3333 1039 -3333 0 feedthrough
rlabel pdiffusion 1046 -3333 1046 -3333 0 feedthrough
rlabel pdiffusion 1053 -3333 1053 -3333 0 feedthrough
rlabel pdiffusion 1060 -3333 1060 -3333 0 feedthrough
rlabel pdiffusion 1067 -3333 1067 -3333 0 cellNo=681
rlabel pdiffusion 1074 -3333 1074 -3333 0 feedthrough
rlabel pdiffusion 1081 -3333 1081 -3333 0 cellNo=185
rlabel pdiffusion 1088 -3333 1088 -3333 0 feedthrough
rlabel pdiffusion 1095 -3333 1095 -3333 0 cellNo=774
rlabel pdiffusion 1102 -3333 1102 -3333 0 cellNo=384
rlabel pdiffusion 1109 -3333 1109 -3333 0 feedthrough
rlabel pdiffusion 1116 -3333 1116 -3333 0 feedthrough
rlabel pdiffusion 1123 -3333 1123 -3333 0 feedthrough
rlabel pdiffusion 1130 -3333 1130 -3333 0 feedthrough
rlabel pdiffusion 1137 -3333 1137 -3333 0 feedthrough
rlabel pdiffusion 1144 -3333 1144 -3333 0 feedthrough
rlabel pdiffusion 1151 -3333 1151 -3333 0 feedthrough
rlabel pdiffusion 1158 -3333 1158 -3333 0 feedthrough
rlabel pdiffusion 1165 -3333 1165 -3333 0 feedthrough
rlabel pdiffusion 1172 -3333 1172 -3333 0 feedthrough
rlabel pdiffusion 1179 -3333 1179 -3333 0 feedthrough
rlabel pdiffusion 1186 -3333 1186 -3333 0 feedthrough
rlabel pdiffusion 1193 -3333 1193 -3333 0 feedthrough
rlabel pdiffusion 1200 -3333 1200 -3333 0 feedthrough
rlabel pdiffusion 1207 -3333 1207 -3333 0 feedthrough
rlabel pdiffusion 1214 -3333 1214 -3333 0 cellNo=932
rlabel pdiffusion 1221 -3333 1221 -3333 0 feedthrough
rlabel pdiffusion 1228 -3333 1228 -3333 0 feedthrough
rlabel pdiffusion 1235 -3333 1235 -3333 0 cellNo=759
rlabel pdiffusion 1242 -3333 1242 -3333 0 feedthrough
rlabel pdiffusion 1249 -3333 1249 -3333 0 feedthrough
rlabel pdiffusion 1256 -3333 1256 -3333 0 feedthrough
rlabel pdiffusion 1263 -3333 1263 -3333 0 feedthrough
rlabel pdiffusion 1270 -3333 1270 -3333 0 cellNo=816
rlabel pdiffusion 1277 -3333 1277 -3333 0 feedthrough
rlabel pdiffusion 1284 -3333 1284 -3333 0 feedthrough
rlabel pdiffusion 1291 -3333 1291 -3333 0 feedthrough
rlabel pdiffusion 1298 -3333 1298 -3333 0 feedthrough
rlabel pdiffusion 1305 -3333 1305 -3333 0 feedthrough
rlabel pdiffusion 1312 -3333 1312 -3333 0 feedthrough
rlabel pdiffusion 1319 -3333 1319 -3333 0 feedthrough
rlabel pdiffusion 1326 -3333 1326 -3333 0 feedthrough
rlabel pdiffusion 1333 -3333 1333 -3333 0 feedthrough
rlabel pdiffusion 1340 -3333 1340 -3333 0 cellNo=332
rlabel pdiffusion 1347 -3333 1347 -3333 0 feedthrough
rlabel pdiffusion 1354 -3333 1354 -3333 0 feedthrough
rlabel pdiffusion 1361 -3333 1361 -3333 0 feedthrough
rlabel pdiffusion 1368 -3333 1368 -3333 0 cellNo=525
rlabel pdiffusion 1375 -3333 1375 -3333 0 feedthrough
rlabel pdiffusion 1382 -3333 1382 -3333 0 cellNo=747
rlabel pdiffusion 1389 -3333 1389 -3333 0 feedthrough
rlabel pdiffusion 1396 -3333 1396 -3333 0 feedthrough
rlabel pdiffusion 1403 -3333 1403 -3333 0 feedthrough
rlabel pdiffusion 1410 -3333 1410 -3333 0 feedthrough
rlabel pdiffusion 1417 -3333 1417 -3333 0 cellNo=982
rlabel pdiffusion 1424 -3333 1424 -3333 0 feedthrough
rlabel pdiffusion 1431 -3333 1431 -3333 0 feedthrough
rlabel pdiffusion 1438 -3333 1438 -3333 0 feedthrough
rlabel pdiffusion 1445 -3333 1445 -3333 0 feedthrough
rlabel pdiffusion 1452 -3333 1452 -3333 0 feedthrough
rlabel pdiffusion 1459 -3333 1459 -3333 0 feedthrough
rlabel pdiffusion 1466 -3333 1466 -3333 0 feedthrough
rlabel pdiffusion 1473 -3333 1473 -3333 0 feedthrough
rlabel pdiffusion 1480 -3333 1480 -3333 0 feedthrough
rlabel pdiffusion 1487 -3333 1487 -3333 0 feedthrough
rlabel pdiffusion 1494 -3333 1494 -3333 0 feedthrough
rlabel pdiffusion 1501 -3333 1501 -3333 0 feedthrough
rlabel pdiffusion 1508 -3333 1508 -3333 0 feedthrough
rlabel pdiffusion 1515 -3333 1515 -3333 0 feedthrough
rlabel pdiffusion 1522 -3333 1522 -3333 0 feedthrough
rlabel pdiffusion 1529 -3333 1529 -3333 0 feedthrough
rlabel pdiffusion 1557 -3333 1557 -3333 0 feedthrough
rlabel pdiffusion 1564 -3333 1564 -3333 0 feedthrough
rlabel pdiffusion 1592 -3333 1592 -3333 0 feedthrough
rlabel pdiffusion 1599 -3333 1599 -3333 0 feedthrough
rlabel pdiffusion 1606 -3333 1606 -3333 0 cellNo=725
rlabel pdiffusion 1627 -3333 1627 -3333 0 feedthrough
rlabel pdiffusion 1655 -3333 1655 -3333 0 feedthrough
rlabel pdiffusion 1662 -3333 1662 -3333 0 feedthrough
rlabel pdiffusion 1669 -3333 1669 -3333 0 feedthrough
rlabel pdiffusion 1718 -3333 1718 -3333 0 feedthrough
rlabel pdiffusion 1725 -3333 1725 -3333 0 cellNo=691
rlabel pdiffusion 1732 -3333 1732 -3333 0 feedthrough
rlabel pdiffusion 1739 -3333 1739 -3333 0 feedthrough
rlabel pdiffusion 1746 -3333 1746 -3333 0 feedthrough
rlabel pdiffusion 1753 -3333 1753 -3333 0 feedthrough
rlabel pdiffusion 1767 -3333 1767 -3333 0 feedthrough
rlabel pdiffusion 1781 -3333 1781 -3333 0 feedthrough
rlabel pdiffusion 1788 -3333 1788 -3333 0 feedthrough
rlabel pdiffusion 1795 -3333 1795 -3333 0 feedthrough
rlabel pdiffusion 1802 -3333 1802 -3333 0 feedthrough
rlabel pdiffusion 1816 -3333 1816 -3333 0 feedthrough
rlabel pdiffusion 1837 -3333 1837 -3333 0 feedthrough
rlabel pdiffusion 1844 -3333 1844 -3333 0 feedthrough
rlabel pdiffusion 1851 -3333 1851 -3333 0 cellNo=953
rlabel pdiffusion 1858 -3333 1858 -3333 0 feedthrough
rlabel pdiffusion 1865 -3333 1865 -3333 0 feedthrough
rlabel pdiffusion 1872 -3333 1872 -3333 0 feedthrough
rlabel pdiffusion 1879 -3333 1879 -3333 0 feedthrough
rlabel pdiffusion 1886 -3333 1886 -3333 0 cellNo=320
rlabel pdiffusion 1893 -3333 1893 -3333 0 feedthrough
rlabel pdiffusion 1907 -3333 1907 -3333 0 feedthrough
rlabel pdiffusion 1963 -3333 1963 -3333 0 feedthrough
rlabel pdiffusion 1970 -3333 1970 -3333 0 feedthrough
rlabel pdiffusion 2026 -3333 2026 -3333 0 feedthrough
rlabel pdiffusion 2033 -3333 2033 -3333 0 feedthrough
rlabel pdiffusion 3 -3420 3 -3420 0 cellNo=1005
rlabel pdiffusion 10 -3420 10 -3420 0 cellNo=1170
rlabel pdiffusion 17 -3420 17 -3420 0 cellNo=1050
rlabel pdiffusion 24 -3420 24 -3420 0 cellNo=1073
rlabel pdiffusion 31 -3420 31 -3420 0 cellNo=1112
rlabel pdiffusion 38 -3420 38 -3420 0 cellNo=1122
rlabel pdiffusion 45 -3420 45 -3420 0 cellNo=1126
rlabel pdiffusion 52 -3420 52 -3420 0 cellNo=1085
rlabel pdiffusion 171 -3420 171 -3420 0 cellNo=621
rlabel pdiffusion 178 -3420 178 -3420 0 cellNo=21
rlabel pdiffusion 297 -3420 297 -3420 0 feedthrough
rlabel pdiffusion 311 -3420 311 -3420 0 feedthrough
rlabel pdiffusion 318 -3420 318 -3420 0 cellNo=874
rlabel pdiffusion 332 -3420 332 -3420 0 feedthrough
rlabel pdiffusion 339 -3420 339 -3420 0 feedthrough
rlabel pdiffusion 346 -3420 346 -3420 0 feedthrough
rlabel pdiffusion 360 -3420 360 -3420 0 feedthrough
rlabel pdiffusion 374 -3420 374 -3420 0 feedthrough
rlabel pdiffusion 381 -3420 381 -3420 0 feedthrough
rlabel pdiffusion 388 -3420 388 -3420 0 cellNo=701
rlabel pdiffusion 395 -3420 395 -3420 0 feedthrough
rlabel pdiffusion 402 -3420 402 -3420 0 cellNo=23
rlabel pdiffusion 409 -3420 409 -3420 0 feedthrough
rlabel pdiffusion 423 -3420 423 -3420 0 feedthrough
rlabel pdiffusion 430 -3420 430 -3420 0 feedthrough
rlabel pdiffusion 437 -3420 437 -3420 0 cellNo=100
rlabel pdiffusion 444 -3420 444 -3420 0 feedthrough
rlabel pdiffusion 451 -3420 451 -3420 0 feedthrough
rlabel pdiffusion 458 -3420 458 -3420 0 feedthrough
rlabel pdiffusion 465 -3420 465 -3420 0 feedthrough
rlabel pdiffusion 472 -3420 472 -3420 0 cellNo=800
rlabel pdiffusion 479 -3420 479 -3420 0 feedthrough
rlabel pdiffusion 486 -3420 486 -3420 0 cellNo=670
rlabel pdiffusion 493 -3420 493 -3420 0 feedthrough
rlabel pdiffusion 500 -3420 500 -3420 0 feedthrough
rlabel pdiffusion 507 -3420 507 -3420 0 feedthrough
rlabel pdiffusion 514 -3420 514 -3420 0 feedthrough
rlabel pdiffusion 521 -3420 521 -3420 0 feedthrough
rlabel pdiffusion 528 -3420 528 -3420 0 feedthrough
rlabel pdiffusion 535 -3420 535 -3420 0 feedthrough
rlabel pdiffusion 542 -3420 542 -3420 0 feedthrough
rlabel pdiffusion 549 -3420 549 -3420 0 feedthrough
rlabel pdiffusion 556 -3420 556 -3420 0 cellNo=600
rlabel pdiffusion 563 -3420 563 -3420 0 feedthrough
rlabel pdiffusion 570 -3420 570 -3420 0 feedthrough
rlabel pdiffusion 577 -3420 577 -3420 0 feedthrough
rlabel pdiffusion 584 -3420 584 -3420 0 feedthrough
rlabel pdiffusion 591 -3420 591 -3420 0 feedthrough
rlabel pdiffusion 598 -3420 598 -3420 0 feedthrough
rlabel pdiffusion 605 -3420 605 -3420 0 feedthrough
rlabel pdiffusion 612 -3420 612 -3420 0 feedthrough
rlabel pdiffusion 619 -3420 619 -3420 0 feedthrough
rlabel pdiffusion 626 -3420 626 -3420 0 feedthrough
rlabel pdiffusion 633 -3420 633 -3420 0 feedthrough
rlabel pdiffusion 640 -3420 640 -3420 0 feedthrough
rlabel pdiffusion 647 -3420 647 -3420 0 feedthrough
rlabel pdiffusion 654 -3420 654 -3420 0 feedthrough
rlabel pdiffusion 661 -3420 661 -3420 0 feedthrough
rlabel pdiffusion 668 -3420 668 -3420 0 cellNo=712
rlabel pdiffusion 675 -3420 675 -3420 0 feedthrough
rlabel pdiffusion 682 -3420 682 -3420 0 feedthrough
rlabel pdiffusion 689 -3420 689 -3420 0 feedthrough
rlabel pdiffusion 696 -3420 696 -3420 0 feedthrough
rlabel pdiffusion 703 -3420 703 -3420 0 feedthrough
rlabel pdiffusion 710 -3420 710 -3420 0 feedthrough
rlabel pdiffusion 717 -3420 717 -3420 0 feedthrough
rlabel pdiffusion 724 -3420 724 -3420 0 cellNo=499
rlabel pdiffusion 731 -3420 731 -3420 0 feedthrough
rlabel pdiffusion 738 -3420 738 -3420 0 feedthrough
rlabel pdiffusion 745 -3420 745 -3420 0 feedthrough
rlabel pdiffusion 752 -3420 752 -3420 0 feedthrough
rlabel pdiffusion 759 -3420 759 -3420 0 feedthrough
rlabel pdiffusion 766 -3420 766 -3420 0 feedthrough
rlabel pdiffusion 773 -3420 773 -3420 0 feedthrough
rlabel pdiffusion 780 -3420 780 -3420 0 feedthrough
rlabel pdiffusion 787 -3420 787 -3420 0 feedthrough
rlabel pdiffusion 794 -3420 794 -3420 0 feedthrough
rlabel pdiffusion 801 -3420 801 -3420 0 cellNo=968
rlabel pdiffusion 808 -3420 808 -3420 0 feedthrough
rlabel pdiffusion 815 -3420 815 -3420 0 feedthrough
rlabel pdiffusion 822 -3420 822 -3420 0 feedthrough
rlabel pdiffusion 829 -3420 829 -3420 0 feedthrough
rlabel pdiffusion 836 -3420 836 -3420 0 feedthrough
rlabel pdiffusion 843 -3420 843 -3420 0 cellNo=996
rlabel pdiffusion 850 -3420 850 -3420 0 feedthrough
rlabel pdiffusion 857 -3420 857 -3420 0 cellNo=279
rlabel pdiffusion 864 -3420 864 -3420 0 feedthrough
rlabel pdiffusion 871 -3420 871 -3420 0 feedthrough
rlabel pdiffusion 878 -3420 878 -3420 0 feedthrough
rlabel pdiffusion 885 -3420 885 -3420 0 feedthrough
rlabel pdiffusion 892 -3420 892 -3420 0 feedthrough
rlabel pdiffusion 899 -3420 899 -3420 0 cellNo=411
rlabel pdiffusion 906 -3420 906 -3420 0 feedthrough
rlabel pdiffusion 913 -3420 913 -3420 0 feedthrough
rlabel pdiffusion 920 -3420 920 -3420 0 cellNo=979
rlabel pdiffusion 927 -3420 927 -3420 0 feedthrough
rlabel pdiffusion 934 -3420 934 -3420 0 cellNo=146
rlabel pdiffusion 941 -3420 941 -3420 0 feedthrough
rlabel pdiffusion 948 -3420 948 -3420 0 feedthrough
rlabel pdiffusion 955 -3420 955 -3420 0 feedthrough
rlabel pdiffusion 962 -3420 962 -3420 0 feedthrough
rlabel pdiffusion 969 -3420 969 -3420 0 feedthrough
rlabel pdiffusion 976 -3420 976 -3420 0 feedthrough
rlabel pdiffusion 983 -3420 983 -3420 0 feedthrough
rlabel pdiffusion 990 -3420 990 -3420 0 cellNo=135
rlabel pdiffusion 997 -3420 997 -3420 0 feedthrough
rlabel pdiffusion 1004 -3420 1004 -3420 0 feedthrough
rlabel pdiffusion 1011 -3420 1011 -3420 0 feedthrough
rlabel pdiffusion 1018 -3420 1018 -3420 0 feedthrough
rlabel pdiffusion 1025 -3420 1025 -3420 0 cellNo=745
rlabel pdiffusion 1032 -3420 1032 -3420 0 cellNo=927
rlabel pdiffusion 1039 -3420 1039 -3420 0 feedthrough
rlabel pdiffusion 1046 -3420 1046 -3420 0 feedthrough
rlabel pdiffusion 1053 -3420 1053 -3420 0 feedthrough
rlabel pdiffusion 1060 -3420 1060 -3420 0 feedthrough
rlabel pdiffusion 1067 -3420 1067 -3420 0 cellNo=764
rlabel pdiffusion 1074 -3420 1074 -3420 0 feedthrough
rlabel pdiffusion 1081 -3420 1081 -3420 0 feedthrough
rlabel pdiffusion 1088 -3420 1088 -3420 0 feedthrough
rlabel pdiffusion 1095 -3420 1095 -3420 0 feedthrough
rlabel pdiffusion 1102 -3420 1102 -3420 0 feedthrough
rlabel pdiffusion 1109 -3420 1109 -3420 0 feedthrough
rlabel pdiffusion 1116 -3420 1116 -3420 0 feedthrough
rlabel pdiffusion 1123 -3420 1123 -3420 0 cellNo=202
rlabel pdiffusion 1137 -3420 1137 -3420 0 feedthrough
rlabel pdiffusion 1144 -3420 1144 -3420 0 feedthrough
rlabel pdiffusion 1158 -3420 1158 -3420 0 cellNo=721
rlabel pdiffusion 1172 -3420 1172 -3420 0 feedthrough
rlabel pdiffusion 1179 -3420 1179 -3420 0 feedthrough
rlabel pdiffusion 1186 -3420 1186 -3420 0 feedthrough
rlabel pdiffusion 1193 -3420 1193 -3420 0 feedthrough
rlabel pdiffusion 1200 -3420 1200 -3420 0 feedthrough
rlabel pdiffusion 1207 -3420 1207 -3420 0 cellNo=531
rlabel pdiffusion 1214 -3420 1214 -3420 0 feedthrough
rlabel pdiffusion 1221 -3420 1221 -3420 0 feedthrough
rlabel pdiffusion 1228 -3420 1228 -3420 0 feedthrough
rlabel pdiffusion 1235 -3420 1235 -3420 0 feedthrough
rlabel pdiffusion 1242 -3420 1242 -3420 0 feedthrough
rlabel pdiffusion 1249 -3420 1249 -3420 0 feedthrough
rlabel pdiffusion 1256 -3420 1256 -3420 0 feedthrough
rlabel pdiffusion 1263 -3420 1263 -3420 0 feedthrough
rlabel pdiffusion 1270 -3420 1270 -3420 0 feedthrough
rlabel pdiffusion 1277 -3420 1277 -3420 0 cellNo=992
rlabel pdiffusion 1284 -3420 1284 -3420 0 feedthrough
rlabel pdiffusion 1291 -3420 1291 -3420 0 feedthrough
rlabel pdiffusion 1298 -3420 1298 -3420 0 feedthrough
rlabel pdiffusion 1305 -3420 1305 -3420 0 cellNo=515
rlabel pdiffusion 1333 -3420 1333 -3420 0 feedthrough
rlabel pdiffusion 1347 -3420 1347 -3420 0 feedthrough
rlabel pdiffusion 1361 -3420 1361 -3420 0 feedthrough
rlabel pdiffusion 1368 -3420 1368 -3420 0 feedthrough
rlabel pdiffusion 1375 -3420 1375 -3420 0 cellNo=260
rlabel pdiffusion 1382 -3420 1382 -3420 0 feedthrough
rlabel pdiffusion 1452 -3420 1452 -3420 0 feedthrough
rlabel pdiffusion 1459 -3420 1459 -3420 0 feedthrough
rlabel pdiffusion 1466 -3420 1466 -3420 0 feedthrough
rlabel pdiffusion 1473 -3420 1473 -3420 0 feedthrough
rlabel pdiffusion 1501 -3420 1501 -3420 0 feedthrough
rlabel pdiffusion 1522 -3420 1522 -3420 0 feedthrough
rlabel pdiffusion 1529 -3420 1529 -3420 0 feedthrough
rlabel pdiffusion 1550 -3420 1550 -3420 0 cellNo=318
rlabel pdiffusion 1585 -3420 1585 -3420 0 cellNo=596
rlabel pdiffusion 1613 -3420 1613 -3420 0 feedthrough
rlabel pdiffusion 1648 -3420 1648 -3420 0 feedthrough
rlabel pdiffusion 1655 -3420 1655 -3420 0 feedthrough
rlabel pdiffusion 1725 -3420 1725 -3420 0 feedthrough
rlabel pdiffusion 1732 -3420 1732 -3420 0 feedthrough
rlabel pdiffusion 1739 -3420 1739 -3420 0 feedthrough
rlabel pdiffusion 1760 -3420 1760 -3420 0 feedthrough
rlabel pdiffusion 1767 -3420 1767 -3420 0 cellNo=42
rlabel pdiffusion 1781 -3420 1781 -3420 0 feedthrough
rlabel pdiffusion 1788 -3420 1788 -3420 0 feedthrough
rlabel pdiffusion 1802 -3420 1802 -3420 0 feedthrough
rlabel pdiffusion 1809 -3420 1809 -3420 0 cellNo=916
rlabel pdiffusion 1823 -3420 1823 -3420 0 feedthrough
rlabel pdiffusion 1830 -3420 1830 -3420 0 feedthrough
rlabel pdiffusion 1837 -3420 1837 -3420 0 feedthrough
rlabel pdiffusion 1844 -3420 1844 -3420 0 feedthrough
rlabel pdiffusion 1851 -3420 1851 -3420 0 feedthrough
rlabel pdiffusion 1858 -3420 1858 -3420 0 feedthrough
rlabel pdiffusion 1865 -3420 1865 -3420 0 feedthrough
rlabel pdiffusion 1872 -3420 1872 -3420 0 feedthrough
rlabel pdiffusion 1956 -3420 1956 -3420 0 feedthrough
rlabel pdiffusion 1963 -3420 1963 -3420 0 feedthrough
rlabel pdiffusion 2026 -3420 2026 -3420 0 feedthrough
rlabel pdiffusion 2033 -3420 2033 -3420 0 feedthrough
rlabel pdiffusion 3 -3465 3 -3465 0 cellNo=1008
rlabel pdiffusion 10 -3465 10 -3465 0 cellNo=1200
rlabel pdiffusion 17 -3465 17 -3465 0 cellNo=1131
rlabel pdiffusion 24 -3465 24 -3465 0 cellNo=1030
rlabel pdiffusion 31 -3465 31 -3465 0 cellNo=1119
rlabel pdiffusion 38 -3465 38 -3465 0 cellNo=1127
rlabel pdiffusion 45 -3465 45 -3465 0 cellNo=1169
rlabel pdiffusion 52 -3465 52 -3465 0 cellNo=1036
rlabel pdiffusion 59 -3465 59 -3465 0 cellNo=1049
rlabel pdiffusion 66 -3465 66 -3465 0 cellNo=1243
rlabel pdiffusion 73 -3465 73 -3465 0 cellNo=1191
rlabel pdiffusion 171 -3465 171 -3465 0 cellNo=354
rlabel pdiffusion 269 -3465 269 -3465 0 cellNo=562
rlabel pdiffusion 325 -3465 325 -3465 0 feedthrough
rlabel pdiffusion 381 -3465 381 -3465 0 feedthrough
rlabel pdiffusion 416 -3465 416 -3465 0 feedthrough
rlabel pdiffusion 423 -3465 423 -3465 0 feedthrough
rlabel pdiffusion 437 -3465 437 -3465 0 cellNo=702
rlabel pdiffusion 444 -3465 444 -3465 0 feedthrough
rlabel pdiffusion 458 -3465 458 -3465 0 feedthrough
rlabel pdiffusion 465 -3465 465 -3465 0 cellNo=834
rlabel pdiffusion 486 -3465 486 -3465 0 feedthrough
rlabel pdiffusion 493 -3465 493 -3465 0 feedthrough
rlabel pdiffusion 500 -3465 500 -3465 0 feedthrough
rlabel pdiffusion 507 -3465 507 -3465 0 feedthrough
rlabel pdiffusion 514 -3465 514 -3465 0 feedthrough
rlabel pdiffusion 521 -3465 521 -3465 0 cellNo=187
rlabel pdiffusion 535 -3465 535 -3465 0 feedthrough
rlabel pdiffusion 542 -3465 542 -3465 0 feedthrough
rlabel pdiffusion 549 -3465 549 -3465 0 cellNo=498
rlabel pdiffusion 556 -3465 556 -3465 0 feedthrough
rlabel pdiffusion 563 -3465 563 -3465 0 feedthrough
rlabel pdiffusion 570 -3465 570 -3465 0 feedthrough
rlabel pdiffusion 577 -3465 577 -3465 0 cellNo=765
rlabel pdiffusion 584 -3465 584 -3465 0 feedthrough
rlabel pdiffusion 591 -3465 591 -3465 0 cellNo=879
rlabel pdiffusion 598 -3465 598 -3465 0 feedthrough
rlabel pdiffusion 605 -3465 605 -3465 0 feedthrough
rlabel pdiffusion 612 -3465 612 -3465 0 feedthrough
rlabel pdiffusion 619 -3465 619 -3465 0 cellNo=277
rlabel pdiffusion 626 -3465 626 -3465 0 cellNo=792
rlabel pdiffusion 633 -3465 633 -3465 0 feedthrough
rlabel pdiffusion 640 -3465 640 -3465 0 cellNo=744
rlabel pdiffusion 647 -3465 647 -3465 0 feedthrough
rlabel pdiffusion 654 -3465 654 -3465 0 feedthrough
rlabel pdiffusion 661 -3465 661 -3465 0 feedthrough
rlabel pdiffusion 668 -3465 668 -3465 0 feedthrough
rlabel pdiffusion 675 -3465 675 -3465 0 feedthrough
rlabel pdiffusion 682 -3465 682 -3465 0 cellNo=802
rlabel pdiffusion 689 -3465 689 -3465 0 feedthrough
rlabel pdiffusion 696 -3465 696 -3465 0 feedthrough
rlabel pdiffusion 703 -3465 703 -3465 0 cellNo=506
rlabel pdiffusion 710 -3465 710 -3465 0 feedthrough
rlabel pdiffusion 717 -3465 717 -3465 0 feedthrough
rlabel pdiffusion 724 -3465 724 -3465 0 feedthrough
rlabel pdiffusion 731 -3465 731 -3465 0 cellNo=14
rlabel pdiffusion 738 -3465 738 -3465 0 feedthrough
rlabel pdiffusion 745 -3465 745 -3465 0 feedthrough
rlabel pdiffusion 752 -3465 752 -3465 0 feedthrough
rlabel pdiffusion 759 -3465 759 -3465 0 feedthrough
rlabel pdiffusion 780 -3465 780 -3465 0 feedthrough
rlabel pdiffusion 794 -3465 794 -3465 0 feedthrough
rlabel pdiffusion 801 -3465 801 -3465 0 feedthrough
rlabel pdiffusion 808 -3465 808 -3465 0 feedthrough
rlabel pdiffusion 815 -3465 815 -3465 0 feedthrough
rlabel pdiffusion 822 -3465 822 -3465 0 feedthrough
rlabel pdiffusion 829 -3465 829 -3465 0 feedthrough
rlabel pdiffusion 836 -3465 836 -3465 0 feedthrough
rlabel pdiffusion 843 -3465 843 -3465 0 feedthrough
rlabel pdiffusion 850 -3465 850 -3465 0 feedthrough
rlabel pdiffusion 878 -3465 878 -3465 0 feedthrough
rlabel pdiffusion 885 -3465 885 -3465 0 feedthrough
rlabel pdiffusion 913 -3465 913 -3465 0 cellNo=987
rlabel pdiffusion 920 -3465 920 -3465 0 cellNo=781
rlabel pdiffusion 955 -3465 955 -3465 0 feedthrough
rlabel pdiffusion 976 -3465 976 -3465 0 feedthrough
rlabel pdiffusion 997 -3465 997 -3465 0 feedthrough
rlabel pdiffusion 1004 -3465 1004 -3465 0 feedthrough
rlabel pdiffusion 1011 -3465 1011 -3465 0 feedthrough
rlabel pdiffusion 1018 -3465 1018 -3465 0 feedthrough
rlabel pdiffusion 1025 -3465 1025 -3465 0 feedthrough
rlabel pdiffusion 1032 -3465 1032 -3465 0 feedthrough
rlabel pdiffusion 1039 -3465 1039 -3465 0 feedthrough
rlabel pdiffusion 1046 -3465 1046 -3465 0 feedthrough
rlabel pdiffusion 1053 -3465 1053 -3465 0 feedthrough
rlabel pdiffusion 1060 -3465 1060 -3465 0 cellNo=673
rlabel pdiffusion 1067 -3465 1067 -3465 0 feedthrough
rlabel pdiffusion 1074 -3465 1074 -3465 0 feedthrough
rlabel pdiffusion 1081 -3465 1081 -3465 0 cellNo=565
rlabel pdiffusion 1088 -3465 1088 -3465 0 feedthrough
rlabel pdiffusion 1095 -3465 1095 -3465 0 feedthrough
rlabel pdiffusion 1102 -3465 1102 -3465 0 feedthrough
rlabel pdiffusion 1109 -3465 1109 -3465 0 feedthrough
rlabel pdiffusion 1123 -3465 1123 -3465 0 cellNo=871
rlabel pdiffusion 1130 -3465 1130 -3465 0 feedthrough
rlabel pdiffusion 1158 -3465 1158 -3465 0 feedthrough
rlabel pdiffusion 1165 -3465 1165 -3465 0 feedthrough
rlabel pdiffusion 1172 -3465 1172 -3465 0 feedthrough
rlabel pdiffusion 1179 -3465 1179 -3465 0 cellNo=918
rlabel pdiffusion 1186 -3465 1186 -3465 0 feedthrough
rlabel pdiffusion 1193 -3465 1193 -3465 0 feedthrough
rlabel pdiffusion 1200 -3465 1200 -3465 0 feedthrough
rlabel pdiffusion 1207 -3465 1207 -3465 0 feedthrough
rlabel pdiffusion 1214 -3465 1214 -3465 0 feedthrough
rlabel pdiffusion 1221 -3465 1221 -3465 0 feedthrough
rlabel pdiffusion 1228 -3465 1228 -3465 0 feedthrough
rlabel pdiffusion 1235 -3465 1235 -3465 0 feedthrough
rlabel pdiffusion 1242 -3465 1242 -3465 0 feedthrough
rlabel pdiffusion 1249 -3465 1249 -3465 0 feedthrough
rlabel pdiffusion 1284 -3465 1284 -3465 0 cellNo=719
rlabel pdiffusion 1291 -3465 1291 -3465 0 feedthrough
rlabel pdiffusion 1305 -3465 1305 -3465 0 cellNo=304
rlabel pdiffusion 1312 -3465 1312 -3465 0 feedthrough
rlabel pdiffusion 1319 -3465 1319 -3465 0 cellNo=895
rlabel pdiffusion 1326 -3465 1326 -3465 0 feedthrough
rlabel pdiffusion 1333 -3465 1333 -3465 0 feedthrough
rlabel pdiffusion 1361 -3465 1361 -3465 0 feedthrough
rlabel pdiffusion 1438 -3465 1438 -3465 0 feedthrough
rlabel pdiffusion 1445 -3465 1445 -3465 0 feedthrough
rlabel pdiffusion 1452 -3465 1452 -3465 0 feedthrough
rlabel pdiffusion 1459 -3465 1459 -3465 0 cellNo=229
rlabel pdiffusion 1466 -3465 1466 -3465 0 feedthrough
rlabel pdiffusion 1494 -3465 1494 -3465 0 feedthrough
rlabel pdiffusion 1501 -3465 1501 -3465 0 feedthrough
rlabel pdiffusion 1515 -3465 1515 -3465 0 feedthrough
rlabel pdiffusion 1522 -3465 1522 -3465 0 feedthrough
rlabel pdiffusion 1627 -3465 1627 -3465 0 cellNo=941
rlabel pdiffusion 1641 -3465 1641 -3465 0 feedthrough
rlabel pdiffusion 1725 -3465 1725 -3465 0 feedthrough
rlabel pdiffusion 1732 -3465 1732 -3465 0 feedthrough
rlabel pdiffusion 1746 -3465 1746 -3465 0 cellNo=846
rlabel pdiffusion 1767 -3465 1767 -3465 0 feedthrough
rlabel pdiffusion 1781 -3465 1781 -3465 0 feedthrough
rlabel pdiffusion 1795 -3465 1795 -3465 0 feedthrough
rlabel pdiffusion 1823 -3465 1823 -3465 0 feedthrough
rlabel pdiffusion 1830 -3465 1830 -3465 0 feedthrough
rlabel pdiffusion 1837 -3465 1837 -3465 0 cellNo=703
rlabel pdiffusion 1844 -3465 1844 -3465 0 feedthrough
rlabel pdiffusion 1851 -3465 1851 -3465 0 feedthrough
rlabel pdiffusion 1858 -3465 1858 -3465 0 cellNo=784
rlabel pdiffusion 1865 -3465 1865 -3465 0 feedthrough
rlabel pdiffusion 1872 -3465 1872 -3465 0 feedthrough
rlabel pdiffusion 1956 -3465 1956 -3465 0 feedthrough
rlabel pdiffusion 1963 -3465 1963 -3465 0 feedthrough
rlabel pdiffusion 2026 -3465 2026 -3465 0 feedthrough
rlabel pdiffusion 2033 -3465 2033 -3465 0 feedthrough
rlabel pdiffusion 3 -3494 3 -3494 0 cellNo=1015
rlabel pdiffusion 10 -3494 10 -3494 0 cellNo=1016
rlabel pdiffusion 17 -3494 17 -3494 0 cellNo=1017
rlabel pdiffusion 24 -3494 24 -3494 0 cellNo=1018
rlabel pdiffusion 31 -3494 31 -3494 0 cellNo=1019
rlabel pdiffusion 38 -3494 38 -3494 0 cellNo=1020
rlabel pdiffusion 45 -3494 45 -3494 0 cellNo=1021
rlabel pdiffusion 52 -3494 52 -3494 0 cellNo=1022
rlabel pdiffusion 59 -3494 59 -3494 0 cellNo=1023
rlabel pdiffusion 66 -3494 66 -3494 0 cellNo=1024
rlabel pdiffusion 73 -3494 73 -3494 0 cellNo=1025
rlabel pdiffusion 80 -3494 80 -3494 0 cellNo=1027
rlabel pdiffusion 87 -3494 87 -3494 0 cellNo=1031
rlabel pdiffusion 94 -3494 94 -3494 0 cellNo=1032
rlabel pdiffusion 101 -3494 101 -3494 0 cellNo=1078
rlabel pdiffusion 108 -3494 108 -3494 0 cellNo=1199
rlabel pdiffusion 115 -3494 115 -3494 0 cellNo=1089
rlabel pdiffusion 122 -3494 122 -3494 0 cellNo=1090
rlabel pdiffusion 129 -3494 129 -3494 0 cellNo=1130
rlabel pdiffusion 136 -3494 136 -3494 0 cellNo=1168
rlabel pdiffusion 143 -3494 143 -3494 0 cellNo=1238
rlabel pdiffusion 150 -3494 150 -3494 0 cellNo=1283
rlabel pdiffusion 332 -3494 332 -3494 0 feedthrough
rlabel pdiffusion 367 -3494 367 -3494 0 cellNo=415
rlabel pdiffusion 388 -3494 388 -3494 0 feedthrough
rlabel pdiffusion 395 -3494 395 -3494 0 feedthrough
rlabel pdiffusion 430 -3494 430 -3494 0 cellNo=957
rlabel pdiffusion 465 -3494 465 -3494 0 feedthrough
rlabel pdiffusion 472 -3494 472 -3494 0 feedthrough
rlabel pdiffusion 479 -3494 479 -3494 0 feedthrough
rlabel pdiffusion 486 -3494 486 -3494 0 feedthrough
rlabel pdiffusion 521 -3494 521 -3494 0 cellNo=887
rlabel pdiffusion 535 -3494 535 -3494 0 feedthrough
rlabel pdiffusion 542 -3494 542 -3494 0 feedthrough
rlabel pdiffusion 570 -3494 570 -3494 0 feedthrough
rlabel pdiffusion 584 -3494 584 -3494 0 feedthrough
rlabel pdiffusion 591 -3494 591 -3494 0 feedthrough
rlabel pdiffusion 605 -3494 605 -3494 0 feedthrough
rlabel pdiffusion 612 -3494 612 -3494 0 feedthrough
rlabel pdiffusion 619 -3494 619 -3494 0 feedthrough
rlabel pdiffusion 633 -3494 633 -3494 0 feedthrough
rlabel pdiffusion 640 -3494 640 -3494 0 feedthrough
rlabel pdiffusion 647 -3494 647 -3494 0 feedthrough
rlabel pdiffusion 654 -3494 654 -3494 0 cellNo=875
rlabel pdiffusion 682 -3494 682 -3494 0 feedthrough
rlabel pdiffusion 717 -3494 717 -3494 0 feedthrough
rlabel pdiffusion 738 -3494 738 -3494 0 feedthrough
rlabel pdiffusion 745 -3494 745 -3494 0 feedthrough
rlabel pdiffusion 752 -3494 752 -3494 0 feedthrough
rlabel pdiffusion 759 -3494 759 -3494 0 feedthrough
rlabel pdiffusion 766 -3494 766 -3494 0 feedthrough
rlabel pdiffusion 773 -3494 773 -3494 0 feedthrough
rlabel pdiffusion 780 -3494 780 -3494 0 feedthrough
rlabel pdiffusion 787 -3494 787 -3494 0 cellNo=837
rlabel pdiffusion 794 -3494 794 -3494 0 feedthrough
rlabel pdiffusion 815 -3494 815 -3494 0 feedthrough
rlabel pdiffusion 829 -3494 829 -3494 0 feedthrough
rlabel pdiffusion 843 -3494 843 -3494 0 feedthrough
rlabel pdiffusion 864 -3494 864 -3494 0 cellNo=919
rlabel pdiffusion 871 -3494 871 -3494 0 feedthrough
rlabel pdiffusion 885 -3494 885 -3494 0 cellNo=733
rlabel pdiffusion 899 -3494 899 -3494 0 feedthrough
rlabel pdiffusion 976 -3494 976 -3494 0 feedthrough
rlabel pdiffusion 997 -3494 997 -3494 0 feedthrough
rlabel pdiffusion 1011 -3494 1011 -3494 0 feedthrough
rlabel pdiffusion 1018 -3494 1018 -3494 0 feedthrough
rlabel pdiffusion 1025 -3494 1025 -3494 0 feedthrough
rlabel pdiffusion 1032 -3494 1032 -3494 0 feedthrough
rlabel pdiffusion 1039 -3494 1039 -3494 0 feedthrough
rlabel pdiffusion 1046 -3494 1046 -3494 0 feedthrough
rlabel pdiffusion 1053 -3494 1053 -3494 0 feedthrough
rlabel pdiffusion 1060 -3494 1060 -3494 0 feedthrough
rlabel pdiffusion 1067 -3494 1067 -3494 0 feedthrough
rlabel pdiffusion 1081 -3494 1081 -3494 0 feedthrough
rlabel pdiffusion 1144 -3494 1144 -3494 0 feedthrough
rlabel pdiffusion 1179 -3494 1179 -3494 0 feedthrough
rlabel pdiffusion 1193 -3494 1193 -3494 0 feedthrough
rlabel pdiffusion 1235 -3494 1235 -3494 0 feedthrough
rlabel pdiffusion 1242 -3494 1242 -3494 0 feedthrough
rlabel pdiffusion 1249 -3494 1249 -3494 0 cellNo=726
rlabel pdiffusion 1256 -3494 1256 -3494 0 feedthrough
rlabel pdiffusion 1263 -3494 1263 -3494 0 cellNo=949
rlabel pdiffusion 1270 -3494 1270 -3494 0 cellNo=40
rlabel pdiffusion 1277 -3494 1277 -3494 0 feedthrough
rlabel pdiffusion 1284 -3494 1284 -3494 0 cellNo=988
rlabel pdiffusion 1291 -3494 1291 -3494 0 feedthrough
rlabel pdiffusion 1305 -3494 1305 -3494 0 feedthrough
rlabel pdiffusion 1312 -3494 1312 -3494 0 cellNo=73
rlabel pdiffusion 1361 -3494 1361 -3494 0 feedthrough
rlabel pdiffusion 1431 -3494 1431 -3494 0 cellNo=985
rlabel pdiffusion 1438 -3494 1438 -3494 0 feedthrough
rlabel pdiffusion 1494 -3494 1494 -3494 0 feedthrough
rlabel pdiffusion 1501 -3494 1501 -3494 0 cellNo=763
rlabel pdiffusion 1508 -3494 1508 -3494 0 feedthrough
rlabel pdiffusion 1515 -3494 1515 -3494 0 feedthrough
rlabel pdiffusion 1522 -3494 1522 -3494 0 feedthrough
rlabel pdiffusion 1571 -3494 1571 -3494 0 feedthrough
rlabel pdiffusion 1641 -3494 1641 -3494 0 feedthrough
rlabel pdiffusion 1725 -3494 1725 -3494 0 cellNo=981
rlabel pdiffusion 1732 -3494 1732 -3494 0 feedthrough
rlabel pdiffusion 1781 -3494 1781 -3494 0 feedthrough
rlabel pdiffusion 1788 -3494 1788 -3494 0 cellNo=826
rlabel pdiffusion 1844 -3494 1844 -3494 0 feedthrough
rlabel pdiffusion 1851 -3494 1851 -3494 0 feedthrough
rlabel pdiffusion 1865 -3494 1865 -3494 0 feedthrough
rlabel pdiffusion 1956 -3494 1956 -3494 0 cellNo=819
rlabel pdiffusion 2026 -3494 2026 -3494 0 feedthrough
rlabel pdiffusion 2033 -3494 2033 -3494 0 feedthrough
rlabel pdiffusion 3 -3517 3 -3517 0 cellNo=1033
rlabel pdiffusion 10 -3517 10 -3517 0 cellNo=1055
rlabel pdiffusion 17 -3517 17 -3517 0 cellNo=1056
rlabel pdiffusion 24 -3517 24 -3517 0 cellNo=1057
rlabel pdiffusion 31 -3517 31 -3517 0 cellNo=1058
rlabel pdiffusion 38 -3517 38 -3517 0 cellNo=1059
rlabel pdiffusion 45 -3517 45 -3517 0 cellNo=1060
rlabel pdiffusion 52 -3517 52 -3517 0 cellNo=1061
rlabel pdiffusion 59 -3517 59 -3517 0 cellNo=1062
rlabel pdiffusion 66 -3517 66 -3517 0 cellNo=1063
rlabel pdiffusion 73 -3517 73 -3517 0 cellNo=1064
rlabel pdiffusion 80 -3517 80 -3517 0 cellNo=1065
rlabel pdiffusion 87 -3517 87 -3517 0 cellNo=1066
rlabel pdiffusion 94 -3517 94 -3517 0 cellNo=1054
rlabel pdiffusion 101 -3517 101 -3517 0 cellNo=1067
rlabel pdiffusion 108 -3517 108 -3517 0 cellNo=1070
rlabel pdiffusion 115 -3517 115 -3517 0 cellNo=1071
rlabel pdiffusion 122 -3517 122 -3517 0 cellNo=1079
rlabel pdiffusion 129 -3517 129 -3517 0 cellNo=1081
rlabel pdiffusion 136 -3517 136 -3517 0 cellNo=1082
rlabel pdiffusion 143 -3517 143 -3517 0 cellNo=1151
rlabel pdiffusion 150 -3517 150 -3517 0 cellNo=1088
rlabel pdiffusion 157 -3517 157 -3517 0 cellNo=1092
rlabel pdiffusion 164 -3517 164 -3517 0 cellNo=1123
rlabel pdiffusion 171 -3517 171 -3517 0 cellNo=1129
rlabel pdiffusion 178 -3517 178 -3517 0 cellNo=1186
rlabel pdiffusion 185 -3517 185 -3517 0 cellNo=1160
rlabel pdiffusion 192 -3517 192 -3517 0 cellNo=1167
rlabel pdiffusion 199 -3517 199 -3517 0 cellNo=1208
rlabel pdiffusion 206 -3517 206 -3517 0 cellNo=1282
rlabel pdiffusion 213 -3517 213 -3517 0 cellNo=1323
rlabel pdiffusion 339 -3517 339 -3517 0 cellNo=696
rlabel pdiffusion 395 -3517 395 -3517 0 feedthrough
rlabel pdiffusion 430 -3517 430 -3517 0 feedthrough
rlabel pdiffusion 465 -3517 465 -3517 0 feedthrough
rlabel pdiffusion 479 -3517 479 -3517 0 feedthrough
rlabel pdiffusion 542 -3517 542 -3517 0 feedthrough
rlabel pdiffusion 549 -3517 549 -3517 0 feedthrough
rlabel pdiffusion 577 -3517 577 -3517 0 feedthrough
rlabel pdiffusion 584 -3517 584 -3517 0 feedthrough
rlabel pdiffusion 605 -3517 605 -3517 0 feedthrough
rlabel pdiffusion 612 -3517 612 -3517 0 feedthrough
rlabel pdiffusion 619 -3517 619 -3517 0 feedthrough
rlabel pdiffusion 626 -3517 626 -3517 0 feedthrough
rlabel pdiffusion 633 -3517 633 -3517 0 feedthrough
rlabel pdiffusion 640 -3517 640 -3517 0 feedthrough
rlabel pdiffusion 710 -3517 710 -3517 0 feedthrough
rlabel pdiffusion 731 -3517 731 -3517 0 feedthrough
rlabel pdiffusion 738 -3517 738 -3517 0 feedthrough
rlabel pdiffusion 745 -3517 745 -3517 0 feedthrough
rlabel pdiffusion 752 -3517 752 -3517 0 feedthrough
rlabel pdiffusion 759 -3517 759 -3517 0 feedthrough
rlabel pdiffusion 766 -3517 766 -3517 0 feedthrough
rlabel pdiffusion 773 -3517 773 -3517 0 cellNo=539
rlabel pdiffusion 780 -3517 780 -3517 0 feedthrough
rlabel pdiffusion 787 -3517 787 -3517 0 cellNo=812
rlabel pdiffusion 794 -3517 794 -3517 0 feedthrough
rlabel pdiffusion 801 -3517 801 -3517 0 feedthrough
rlabel pdiffusion 808 -3517 808 -3517 0 cellNo=924
rlabel pdiffusion 892 -3517 892 -3517 0 feedthrough
rlabel pdiffusion 969 -3517 969 -3517 0 feedthrough
rlabel pdiffusion 1004 -3517 1004 -3517 0 feedthrough
rlabel pdiffusion 1011 -3517 1011 -3517 0 feedthrough
rlabel pdiffusion 1018 -3517 1018 -3517 0 feedthrough
rlabel pdiffusion 1025 -3517 1025 -3517 0 feedthrough
rlabel pdiffusion 1032 -3517 1032 -3517 0 feedthrough
rlabel pdiffusion 1039 -3517 1039 -3517 0 feedthrough
rlabel pdiffusion 1046 -3517 1046 -3517 0 feedthrough
rlabel pdiffusion 1053 -3517 1053 -3517 0 feedthrough
rlabel pdiffusion 1060 -3517 1060 -3517 0 cellNo=914
rlabel pdiffusion 1067 -3517 1067 -3517 0 feedthrough
rlabel pdiffusion 1123 -3517 1123 -3517 0 feedthrough
rlabel pdiffusion 1151 -3517 1151 -3517 0 feedthrough
rlabel pdiffusion 1158 -3517 1158 -3517 0 cellNo=973
rlabel pdiffusion 1207 -3517 1207 -3517 0 feedthrough
rlabel pdiffusion 1235 -3517 1235 -3517 0 feedthrough
rlabel pdiffusion 1361 -3517 1361 -3517 0 feedthrough
rlabel pdiffusion 1368 -3517 1368 -3517 0 cellNo=888
rlabel pdiffusion 1508 -3517 1508 -3517 0 feedthrough
rlabel pdiffusion 1515 -3517 1515 -3517 0 feedthrough
rlabel pdiffusion 1522 -3517 1522 -3517 0 feedthrough
rlabel pdiffusion 1613 -3517 1613 -3517 0 feedthrough
rlabel pdiffusion 1641 -3517 1641 -3517 0 feedthrough
rlabel pdiffusion 1851 -3517 1851 -3517 0 feedthrough
rlabel pdiffusion 1858 -3517 1858 -3517 0 cellNo=520
rlabel pdiffusion 2026 -3517 2026 -3517 0 feedthrough
rlabel pdiffusion 2033 -3517 2033 -3517 0 feedthrough
rlabel pdiffusion 3 -3536 3 -3536 0 cellNo=1028
rlabel pdiffusion 10 -3536 10 -3536 0 cellNo=1094
rlabel pdiffusion 17 -3536 17 -3536 0 cellNo=1095
rlabel pdiffusion 24 -3536 24 -3536 0 cellNo=1096
rlabel pdiffusion 31 -3536 31 -3536 0 cellNo=1097
rlabel pdiffusion 38 -3536 38 -3536 0 cellNo=1098
rlabel pdiffusion 45 -3536 45 -3536 0 cellNo=1099
rlabel pdiffusion 52 -3536 52 -3536 0 cellNo=1100
rlabel pdiffusion 59 -3536 59 -3536 0 cellNo=1101
rlabel pdiffusion 66 -3536 66 -3536 0 cellNo=1102
rlabel pdiffusion 73 -3536 73 -3536 0 cellNo=1103
rlabel pdiffusion 80 -3536 80 -3536 0 cellNo=1104
rlabel pdiffusion 87 -3536 87 -3536 0 cellNo=1105
rlabel pdiffusion 94 -3536 94 -3536 0 cellNo=1106
rlabel pdiffusion 101 -3536 101 -3536 0 cellNo=1107
rlabel pdiffusion 108 -3536 108 -3536 0 cellNo=1108
rlabel pdiffusion 115 -3536 115 -3536 0 cellNo=1068
rlabel pdiffusion 122 -3536 122 -3536 0 cellNo=1093
rlabel pdiffusion 129 -3536 129 -3536 0 cellNo=1075
rlabel pdiffusion 136 -3536 136 -3536 0 cellNo=1084
rlabel pdiffusion 143 -3536 143 -3536 0 cellNo=1115
rlabel pdiffusion 150 -3536 150 -3536 0 cellNo=1116
rlabel pdiffusion 157 -3536 157 -3536 0 cellNo=1121
rlabel pdiffusion 164 -3536 164 -3536 0 cellNo=1124
rlabel pdiffusion 171 -3536 171 -3536 0 cellNo=1125
rlabel pdiffusion 178 -3536 178 -3536 0 cellNo=1128
rlabel pdiffusion 185 -3536 185 -3536 0 cellNo=1203
rlabel pdiffusion 192 -3536 192 -3536 0 cellNo=1207
rlabel pdiffusion 199 -3536 199 -3536 0 cellNo=1248
rlabel pdiffusion 206 -3536 206 -3536 0 cellNo=1322
rlabel pdiffusion 213 -3536 213 -3536 0 cellNo=1362
rlabel pdiffusion 395 -3536 395 -3536 0 feedthrough
rlabel pdiffusion 409 -3536 409 -3536 0 feedthrough
rlabel pdiffusion 465 -3536 465 -3536 0 feedthrough
rlabel pdiffusion 472 -3536 472 -3536 0 cellNo=633
rlabel pdiffusion 479 -3536 479 -3536 0 feedthrough
rlabel pdiffusion 542 -3536 542 -3536 0 feedthrough
rlabel pdiffusion 549 -3536 549 -3536 0 feedthrough
rlabel pdiffusion 577 -3536 577 -3536 0 feedthrough
rlabel pdiffusion 584 -3536 584 -3536 0 feedthrough
rlabel pdiffusion 605 -3536 605 -3536 0 feedthrough
rlabel pdiffusion 612 -3536 612 -3536 0 feedthrough
rlabel pdiffusion 619 -3536 619 -3536 0 feedthrough
rlabel pdiffusion 626 -3536 626 -3536 0 cellNo=648
rlabel pdiffusion 633 -3536 633 -3536 0 cellNo=921
rlabel pdiffusion 640 -3536 640 -3536 0 feedthrough
rlabel pdiffusion 647 -3536 647 -3536 0 feedthrough
rlabel pdiffusion 710 -3536 710 -3536 0 feedthrough
rlabel pdiffusion 717 -3536 717 -3536 0 feedthrough
rlabel pdiffusion 724 -3536 724 -3536 0 feedthrough
rlabel pdiffusion 731 -3536 731 -3536 0 feedthrough
rlabel pdiffusion 738 -3536 738 -3536 0 cellNo=523
rlabel pdiffusion 745 -3536 745 -3536 0 feedthrough
rlabel pdiffusion 766 -3536 766 -3536 0 feedthrough
rlabel pdiffusion 787 -3536 787 -3536 0 feedthrough
rlabel pdiffusion 794 -3536 794 -3536 0 feedthrough
rlabel pdiffusion 927 -3536 927 -3536 0 feedthrough
rlabel pdiffusion 969 -3536 969 -3536 0 cellNo=779
rlabel pdiffusion 1011 -3536 1011 -3536 0 feedthrough
rlabel pdiffusion 1025 -3536 1025 -3536 0 cellNo=840
rlabel pdiffusion 1032 -3536 1032 -3536 0 feedthrough
rlabel pdiffusion 1039 -3536 1039 -3536 0 cellNo=178
rlabel pdiffusion 1046 -3536 1046 -3536 0 feedthrough
rlabel pdiffusion 1060 -3536 1060 -3536 0 feedthrough
rlabel pdiffusion 1067 -3536 1067 -3536 0 feedthrough
rlabel pdiffusion 1214 -3536 1214 -3536 0 feedthrough
rlabel pdiffusion 1221 -3536 1221 -3536 0 cellNo=937
rlabel pdiffusion 1508 -3536 1508 -3536 0 feedthrough
rlabel pdiffusion 1515 -3536 1515 -3536 0 feedthrough
rlabel pdiffusion 1522 -3536 1522 -3536 0 feedthrough
rlabel pdiffusion 1634 -3536 1634 -3536 0 feedthrough
rlabel pdiffusion 1641 -3536 1641 -3536 0 feedthrough
rlabel pdiffusion 2026 -3536 2026 -3536 0 feedthrough
rlabel pdiffusion 2033 -3536 2033 -3536 0 feedthrough
rlabel pdiffusion 3 -3551 3 -3551 0 cellNo=1083
rlabel pdiffusion 10 -3551 10 -3551 0 cellNo=1133
rlabel pdiffusion 17 -3551 17 -3551 0 cellNo=1134
rlabel pdiffusion 24 -3551 24 -3551 0 cellNo=1135
rlabel pdiffusion 31 -3551 31 -3551 0 cellNo=1136
rlabel pdiffusion 38 -3551 38 -3551 0 cellNo=1137
rlabel pdiffusion 45 -3551 45 -3551 0 cellNo=1138
rlabel pdiffusion 52 -3551 52 -3551 0 cellNo=1139
rlabel pdiffusion 59 -3551 59 -3551 0 cellNo=1140
rlabel pdiffusion 66 -3551 66 -3551 0 cellNo=1141
rlabel pdiffusion 73 -3551 73 -3551 0 cellNo=1142
rlabel pdiffusion 80 -3551 80 -3551 0 cellNo=1143
rlabel pdiffusion 87 -3551 87 -3551 0 cellNo=1144
rlabel pdiffusion 94 -3551 94 -3551 0 cellNo=1145
rlabel pdiffusion 101 -3551 101 -3551 0 cellNo=1146
rlabel pdiffusion 108 -3551 108 -3551 0 cellNo=1147
rlabel pdiffusion 115 -3551 115 -3551 0 cellNo=1148
rlabel pdiffusion 122 -3551 122 -3551 0 cellNo=1149
rlabel pdiffusion 129 -3551 129 -3551 0 cellNo=1117
rlabel pdiffusion 136 -3551 136 -3551 0 cellNo=1190
rlabel pdiffusion 143 -3551 143 -3551 0 cellNo=1132
rlabel pdiffusion 150 -3551 150 -3551 0 cellNo=1153
rlabel pdiffusion 157 -3551 157 -3551 0 cellNo=1118
rlabel pdiffusion 164 -3551 164 -3551 0 cellNo=1155
rlabel pdiffusion 171 -3551 171 -3551 0 cellNo=1392
rlabel pdiffusion 178 -3551 178 -3551 0 cellNo=1152
rlabel pdiffusion 185 -3551 185 -3551 0 cellNo=1163
rlabel pdiffusion 192 -3551 192 -3551 0 cellNo=1164
rlabel pdiffusion 199 -3551 199 -3551 0 cellNo=1166
rlabel pdiffusion 206 -3551 206 -3551 0 cellNo=1201
rlabel pdiffusion 213 -3551 213 -3551 0 cellNo=1206
rlabel pdiffusion 220 -3551 220 -3551 0 cellNo=1247
rlabel pdiffusion 227 -3551 227 -3551 0 cellNo=1321
rlabel pdiffusion 234 -3551 234 -3551 0 cellNo=1361
rlabel pdiffusion 241 -3551 241 -3551 0 cellNo=1400
rlabel pdiffusion 402 -3551 402 -3551 0 feedthrough
rlabel pdiffusion 409 -3551 409 -3551 0 feedthrough
rlabel pdiffusion 542 -3551 542 -3551 0 feedthrough
rlabel pdiffusion 549 -3551 549 -3551 0 cellNo=659
rlabel pdiffusion 556 -3551 556 -3551 0 feedthrough
rlabel pdiffusion 584 -3551 584 -3551 0 cellNo=486
rlabel pdiffusion 591 -3551 591 -3551 0 feedthrough
rlabel pdiffusion 605 -3551 605 -3551 0 feedthrough
rlabel pdiffusion 612 -3551 612 -3551 0 feedthrough
rlabel pdiffusion 619 -3551 619 -3551 0 feedthrough
rlabel pdiffusion 647 -3551 647 -3551 0 feedthrough
rlabel pdiffusion 703 -3551 703 -3551 0 feedthrough
rlabel pdiffusion 717 -3551 717 -3551 0 feedthrough
rlabel pdiffusion 724 -3551 724 -3551 0 feedthrough
rlabel pdiffusion 731 -3551 731 -3551 0 feedthrough
rlabel pdiffusion 759 -3551 759 -3551 0 feedthrough
rlabel pdiffusion 787 -3551 787 -3551 0 cellNo=698
rlabel pdiffusion 794 -3551 794 -3551 0 feedthrough
rlabel pdiffusion 1018 -3551 1018 -3551 0 cellNo=718
rlabel pdiffusion 1039 -3551 1039 -3551 0 feedthrough
rlabel pdiffusion 1060 -3551 1060 -3551 0 feedthrough
rlabel pdiffusion 1508 -3551 1508 -3551 0 feedthrough
rlabel pdiffusion 1515 -3551 1515 -3551 0 feedthrough
rlabel pdiffusion 1522 -3551 1522 -3551 0 feedthrough
rlabel pdiffusion 1641 -3551 1641 -3551 0 feedthrough
rlabel pdiffusion 1648 -3551 1648 -3551 0 feedthrough
rlabel pdiffusion 2026 -3551 2026 -3551 0 feedthrough
rlabel pdiffusion 2033 -3551 2033 -3551 0 feedthrough
rlabel pdiffusion 3 -3566 3 -3566 0 cellNo=1044
rlabel pdiffusion 10 -3566 10 -3566 0 cellNo=1172
rlabel pdiffusion 17 -3566 17 -3566 0 cellNo=1173
rlabel pdiffusion 24 -3566 24 -3566 0 cellNo=1174
rlabel pdiffusion 31 -3566 31 -3566 0 cellNo=1175
rlabel pdiffusion 38 -3566 38 -3566 0 cellNo=1176
rlabel pdiffusion 45 -3566 45 -3566 0 cellNo=1177
rlabel pdiffusion 52 -3566 52 -3566 0 cellNo=1178
rlabel pdiffusion 59 -3566 59 -3566 0 cellNo=1179
rlabel pdiffusion 66 -3566 66 -3566 0 cellNo=1180
rlabel pdiffusion 73 -3566 73 -3566 0 cellNo=1181
rlabel pdiffusion 80 -3566 80 -3566 0 cellNo=1182
rlabel pdiffusion 87 -3566 87 -3566 0 cellNo=1183
rlabel pdiffusion 94 -3566 94 -3566 0 cellNo=1171
rlabel pdiffusion 101 -3566 101 -3566 0 cellNo=1185
rlabel pdiffusion 108 -3566 108 -3566 0 cellNo=1111
rlabel pdiffusion 115 -3566 115 -3566 0 cellNo=1187
rlabel pdiffusion 122 -3566 122 -3566 0 cellNo=1188
rlabel pdiffusion 129 -3566 129 -3566 0 cellNo=1113
rlabel pdiffusion 136 -3566 136 -3566 0 cellNo=1154
rlabel pdiffusion 143 -3566 143 -3566 0 cellNo=1157
rlabel pdiffusion 150 -3566 150 -3566 0 cellNo=1192
rlabel pdiffusion 157 -3566 157 -3566 0 cellNo=1159
rlabel pdiffusion 164 -3566 164 -3566 0 cellNo=1194
rlabel pdiffusion 171 -3566 171 -3566 0 cellNo=1195
rlabel pdiffusion 178 -3566 178 -3566 0 cellNo=1196
rlabel pdiffusion 185 -3566 185 -3566 0 cellNo=1162
rlabel pdiffusion 192 -3566 192 -3566 0 cellNo=1161
rlabel pdiffusion 199 -3566 199 -3566 0 cellNo=1202
rlabel pdiffusion 206 -3566 206 -3566 0 cellNo=1205
rlabel pdiffusion 213 -3566 213 -3566 0 cellNo=1246
rlabel pdiffusion 220 -3566 220 -3566 0 cellNo=1279
rlabel pdiffusion 227 -3566 227 -3566 0 cellNo=1287
rlabel pdiffusion 234 -3566 234 -3566 0 cellNo=1360
rlabel pdiffusion 241 -3566 241 -3566 0 cellNo=1399
rlabel pdiffusion 402 -3566 402 -3566 0 feedthrough
rlabel pdiffusion 409 -3566 409 -3566 0 feedthrough
rlabel pdiffusion 605 -3566 605 -3566 0 feedthrough
rlabel pdiffusion 612 -3566 612 -3566 0 feedthrough
rlabel pdiffusion 619 -3566 619 -3566 0 feedthrough
rlabel pdiffusion 647 -3566 647 -3566 0 cellNo=628
rlabel pdiffusion 703 -3566 703 -3566 0 feedthrough
rlabel pdiffusion 717 -3566 717 -3566 0 feedthrough
rlabel pdiffusion 724 -3566 724 -3566 0 feedthrough
rlabel pdiffusion 731 -3566 731 -3566 0 feedthrough
rlabel pdiffusion 759 -3566 759 -3566 0 feedthrough
rlabel pdiffusion 1060 -3566 1060 -3566 0 cellNo=578
rlabel pdiffusion 1067 -3566 1067 -3566 0 feedthrough
rlabel pdiffusion 1515 -3566 1515 -3566 0 cellNo=897
rlabel pdiffusion 1522 -3566 1522 -3566 0 feedthrough
rlabel pdiffusion 1641 -3566 1641 -3566 0 feedthrough
rlabel pdiffusion 1648 -3566 1648 -3566 0 feedthrough
rlabel pdiffusion 2026 -3566 2026 -3566 0 cellNo=601
rlabel pdiffusion 3 -3581 3 -3581 0 cellNo=1043
rlabel pdiffusion 10 -3581 10 -3581 0 cellNo=1211
rlabel pdiffusion 17 -3581 17 -3581 0 cellNo=1212
rlabel pdiffusion 24 -3581 24 -3581 0 cellNo=1213
rlabel pdiffusion 31 -3581 31 -3581 0 cellNo=1214
rlabel pdiffusion 38 -3581 38 -3581 0 cellNo=1215
rlabel pdiffusion 45 -3581 45 -3581 0 cellNo=1216
rlabel pdiffusion 52 -3581 52 -3581 0 cellNo=1217
rlabel pdiffusion 59 -3581 59 -3581 0 cellNo=1218
rlabel pdiffusion 66 -3581 66 -3581 0 cellNo=1219
rlabel pdiffusion 73 -3581 73 -3581 0 cellNo=1220
rlabel pdiffusion 80 -3581 80 -3581 0 cellNo=1221
rlabel pdiffusion 87 -3581 87 -3581 0 cellNo=1222
rlabel pdiffusion 94 -3581 94 -3581 0 cellNo=1223
rlabel pdiffusion 101 -3581 101 -3581 0 cellNo=1224
rlabel pdiffusion 108 -3581 108 -3581 0 cellNo=1225
rlabel pdiffusion 115 -3581 115 -3581 0 cellNo=1226
rlabel pdiffusion 122 -3581 122 -3581 0 cellNo=1227
rlabel pdiffusion 129 -3581 129 -3581 0 cellNo=1228
rlabel pdiffusion 136 -3581 136 -3581 0 cellNo=1229
rlabel pdiffusion 143 -3581 143 -3581 0 cellNo=1230
rlabel pdiffusion 150 -3581 150 -3581 0 cellNo=1231
rlabel pdiffusion 157 -3581 157 -3581 0 cellNo=1232
rlabel pdiffusion 164 -3581 164 -3581 0 cellNo=1233
rlabel pdiffusion 171 -3581 171 -3581 0 cellNo=1234
rlabel pdiffusion 178 -3581 178 -3581 0 cellNo=1235
rlabel pdiffusion 185 -3581 185 -3581 0 cellNo=1236
rlabel pdiffusion 192 -3581 192 -3581 0 cellNo=1237
rlabel pdiffusion 199 -3581 199 -3581 0 cellNo=1158
rlabel pdiffusion 206 -3581 206 -3581 0 cellNo=1239
rlabel pdiffusion 213 -3581 213 -3581 0 cellNo=1278
rlabel pdiffusion 220 -3581 220 -3581 0 cellNo=1241
rlabel pdiffusion 227 -3581 227 -3581 0 cellNo=1242
rlabel pdiffusion 234 -3581 234 -3581 0 cellNo=1245
rlabel pdiffusion 241 -3581 241 -3581 0 cellNo=1286
rlabel pdiffusion 248 -3581 248 -3581 0 cellNo=1352
rlabel pdiffusion 255 -3581 255 -3581 0 cellNo=1210
rlabel pdiffusion 262 -3581 262 -3581 0 cellNo=1438
rlabel pdiffusion 269 -3581 269 -3581 0 cellNo=1443
rlabel pdiffusion 402 -3581 402 -3581 0 feedthrough
rlabel pdiffusion 409 -3581 409 -3581 0 feedthrough
rlabel pdiffusion 605 -3581 605 -3581 0 feedthrough
rlabel pdiffusion 612 -3581 612 -3581 0 feedthrough
rlabel pdiffusion 619 -3581 619 -3581 0 feedthrough
rlabel pdiffusion 703 -3581 703 -3581 0 feedthrough
rlabel pdiffusion 717 -3581 717 -3581 0 feedthrough
rlabel pdiffusion 724 -3581 724 -3581 0 feedthrough
rlabel pdiffusion 731 -3581 731 -3581 0 feedthrough
rlabel pdiffusion 759 -3581 759 -3581 0 feedthrough
rlabel pdiffusion 1641 -3581 1641 -3581 0 feedthrough
rlabel pdiffusion 1648 -3581 1648 -3581 0 feedthrough
rlabel pdiffusion 3 -3594 3 -3594 0 cellNo=1249
rlabel pdiffusion 10 -3594 10 -3594 0 cellNo=1250
rlabel pdiffusion 17 -3594 17 -3594 0 cellNo=1251
rlabel pdiffusion 24 -3594 24 -3594 0 cellNo=1252
rlabel pdiffusion 31 -3594 31 -3594 0 cellNo=1253
rlabel pdiffusion 38 -3594 38 -3594 0 cellNo=1254
rlabel pdiffusion 45 -3594 45 -3594 0 cellNo=1255
rlabel pdiffusion 52 -3594 52 -3594 0 cellNo=1256
rlabel pdiffusion 59 -3594 59 -3594 0 cellNo=1257
rlabel pdiffusion 66 -3594 66 -3594 0 cellNo=1258
rlabel pdiffusion 73 -3594 73 -3594 0 cellNo=1259
rlabel pdiffusion 80 -3594 80 -3594 0 cellNo=1260
rlabel pdiffusion 87 -3594 87 -3594 0 cellNo=1261
rlabel pdiffusion 94 -3594 94 -3594 0 cellNo=1262
rlabel pdiffusion 101 -3594 101 -3594 0 cellNo=1263
rlabel pdiffusion 108 -3594 108 -3594 0 cellNo=1264
rlabel pdiffusion 115 -3594 115 -3594 0 cellNo=1265
rlabel pdiffusion 122 -3594 122 -3594 0 cellNo=1266
rlabel pdiffusion 129 -3594 129 -3594 0 cellNo=1267
rlabel pdiffusion 136 -3594 136 -3594 0 cellNo=1268
rlabel pdiffusion 143 -3594 143 -3594 0 cellNo=1269
rlabel pdiffusion 150 -3594 150 -3594 0 cellNo=1270
rlabel pdiffusion 157 -3594 157 -3594 0 cellNo=1271
rlabel pdiffusion 164 -3594 164 -3594 0 cellNo=1272
rlabel pdiffusion 171 -3594 171 -3594 0 cellNo=1273
rlabel pdiffusion 178 -3594 178 -3594 0 cellNo=1274
rlabel pdiffusion 185 -3594 185 -3594 0 cellNo=1275
rlabel pdiffusion 192 -3594 192 -3594 0 cellNo=1276
rlabel pdiffusion 199 -3594 199 -3594 0 cellNo=1277
rlabel pdiffusion 206 -3594 206 -3594 0 cellNo=1396
rlabel pdiffusion 213 -3594 213 -3594 0 cellNo=1317
rlabel pdiffusion 220 -3594 220 -3594 0 cellNo=1280
rlabel pdiffusion 227 -3594 227 -3594 0 cellNo=1281
rlabel pdiffusion 234 -3594 234 -3594 0 cellNo=1285
rlabel pdiffusion 241 -3594 241 -3594 0 cellNo=1326
rlabel pdiffusion 248 -3594 248 -3594 0 cellNo=1442
rlabel pdiffusion 395 -3594 395 -3594 0 feedthrough
rlabel pdiffusion 402 -3594 402 -3594 0 feedthrough
rlabel pdiffusion 605 -3594 605 -3594 0 feedthrough
rlabel pdiffusion 612 -3594 612 -3594 0 feedthrough
rlabel pdiffusion 619 -3594 619 -3594 0 cellNo=484
rlabel pdiffusion 703 -3594 703 -3594 0 feedthrough
rlabel pdiffusion 724 -3594 724 -3594 0 cellNo=964
rlabel pdiffusion 731 -3594 731 -3594 0 feedthrough
rlabel pdiffusion 759 -3594 759 -3594 0 feedthrough
rlabel pdiffusion 1641 -3594 1641 -3594 0 feedthrough
rlabel pdiffusion 1648 -3594 1648 -3594 0 feedthrough
rlabel pdiffusion 3 -3605 3 -3605 0 cellNo=1288
rlabel pdiffusion 10 -3605 10 -3605 0 cellNo=1289
rlabel pdiffusion 17 -3605 17 -3605 0 cellNo=1290
rlabel pdiffusion 24 -3605 24 -3605 0 cellNo=1291
rlabel pdiffusion 31 -3605 31 -3605 0 cellNo=1292
rlabel pdiffusion 38 -3605 38 -3605 0 cellNo=1293
rlabel pdiffusion 45 -3605 45 -3605 0 cellNo=1294
rlabel pdiffusion 52 -3605 52 -3605 0 cellNo=1295
rlabel pdiffusion 59 -3605 59 -3605 0 cellNo=1296
rlabel pdiffusion 66 -3605 66 -3605 0 cellNo=1297
rlabel pdiffusion 73 -3605 73 -3605 0 cellNo=1298
rlabel pdiffusion 80 -3605 80 -3605 0 cellNo=1299
rlabel pdiffusion 87 -3605 87 -3605 0 cellNo=1300
rlabel pdiffusion 94 -3605 94 -3605 0 cellNo=1301
rlabel pdiffusion 101 -3605 101 -3605 0 cellNo=1302
rlabel pdiffusion 108 -3605 108 -3605 0 cellNo=1303
rlabel pdiffusion 115 -3605 115 -3605 0 cellNo=1304
rlabel pdiffusion 122 -3605 122 -3605 0 cellNo=1305
rlabel pdiffusion 129 -3605 129 -3605 0 cellNo=1306
rlabel pdiffusion 136 -3605 136 -3605 0 cellNo=1307
rlabel pdiffusion 143 -3605 143 -3605 0 cellNo=1308
rlabel pdiffusion 150 -3605 150 -3605 0 cellNo=1309
rlabel pdiffusion 157 -3605 157 -3605 0 cellNo=1310
rlabel pdiffusion 164 -3605 164 -3605 0 cellNo=1311
rlabel pdiffusion 171 -3605 171 -3605 0 cellNo=1312
rlabel pdiffusion 178 -3605 178 -3605 0 cellNo=1313
rlabel pdiffusion 185 -3605 185 -3605 0 cellNo=1314
rlabel pdiffusion 192 -3605 192 -3605 0 cellNo=1315
rlabel pdiffusion 199 -3605 199 -3605 0 cellNo=1355
rlabel pdiffusion 206 -3605 206 -3605 0 cellNo=1318
rlabel pdiffusion 213 -3605 213 -3605 0 cellNo=1319
rlabel pdiffusion 220 -3605 220 -3605 0 cellNo=1320
rlabel pdiffusion 227 -3605 227 -3605 0 cellNo=1325
rlabel pdiffusion 234 -3605 234 -3605 0 cellNo=1365
rlabel pdiffusion 241 -3605 241 -3605 0 cellNo=1404
rlabel pdiffusion 248 -3605 248 -3605 0 cellNo=1441
rlabel pdiffusion 395 -3605 395 -3605 0 feedthrough
rlabel pdiffusion 402 -3605 402 -3605 0 feedthrough
rlabel pdiffusion 605 -3605 605 -3605 0 feedthrough
rlabel pdiffusion 612 -3605 612 -3605 0 feedthrough
rlabel pdiffusion 703 -3605 703 -3605 0 cellNo=665
rlabel pdiffusion 759 -3605 759 -3605 0 feedthrough
rlabel pdiffusion 1641 -3605 1641 -3605 0 feedthrough
rlabel pdiffusion 1648 -3605 1648 -3605 0 feedthrough
rlabel pdiffusion 3 -3616 3 -3616 0 cellNo=1042
rlabel pdiffusion 10 -3616 10 -3616 0 cellNo=1328
rlabel pdiffusion 17 -3616 17 -3616 0 cellNo=1329
rlabel pdiffusion 24 -3616 24 -3616 0 cellNo=1330
rlabel pdiffusion 31 -3616 31 -3616 0 cellNo=1331
rlabel pdiffusion 38 -3616 38 -3616 0 cellNo=1332
rlabel pdiffusion 45 -3616 45 -3616 0 cellNo=1333
rlabel pdiffusion 52 -3616 52 -3616 0 cellNo=1334
rlabel pdiffusion 59 -3616 59 -3616 0 cellNo=1335
rlabel pdiffusion 66 -3616 66 -3616 0 cellNo=1336
rlabel pdiffusion 73 -3616 73 -3616 0 cellNo=1337
rlabel pdiffusion 80 -3616 80 -3616 0 cellNo=1338
rlabel pdiffusion 87 -3616 87 -3616 0 cellNo=1339
rlabel pdiffusion 94 -3616 94 -3616 0 cellNo=1340
rlabel pdiffusion 101 -3616 101 -3616 0 cellNo=1341
rlabel pdiffusion 108 -3616 108 -3616 0 cellNo=1342
rlabel pdiffusion 115 -3616 115 -3616 0 cellNo=1343
rlabel pdiffusion 122 -3616 122 -3616 0 cellNo=1344
rlabel pdiffusion 129 -3616 129 -3616 0 cellNo=1345
rlabel pdiffusion 136 -3616 136 -3616 0 cellNo=1346
rlabel pdiffusion 143 -3616 143 -3616 0 cellNo=1347
rlabel pdiffusion 150 -3616 150 -3616 0 cellNo=1348
rlabel pdiffusion 157 -3616 157 -3616 0 cellNo=1349
rlabel pdiffusion 164 -3616 164 -3616 0 cellNo=1350
rlabel pdiffusion 171 -3616 171 -3616 0 cellNo=1327
rlabel pdiffusion 178 -3616 178 -3616 0 cellNo=1114
rlabel pdiffusion 185 -3616 185 -3616 0 cellNo=1353
rlabel pdiffusion 192 -3616 192 -3616 0 cellNo=1354
rlabel pdiffusion 199 -3616 199 -3616 0 cellNo=1316
rlabel pdiffusion 206 -3616 206 -3616 0 cellNo=1356
rlabel pdiffusion 213 -3616 213 -3616 0 cellNo=1358
rlabel pdiffusion 220 -3616 220 -3616 0 cellNo=1359
rlabel pdiffusion 227 -3616 227 -3616 0 cellNo=1364
rlabel pdiffusion 234 -3616 234 -3616 0 cellNo=1403
rlabel pdiffusion 241 -3616 241 -3616 0 cellNo=1440
rlabel pdiffusion 395 -3616 395 -3616 0 feedthrough
rlabel pdiffusion 402 -3616 402 -3616 0 feedthrough
rlabel pdiffusion 605 -3616 605 -3616 0 feedthrough
rlabel pdiffusion 612 -3616 612 -3616 0 feedthrough
rlabel pdiffusion 696 -3616 696 -3616 0 feedthrough
rlabel pdiffusion 759 -3616 759 -3616 0 feedthrough
rlabel pdiffusion 1641 -3616 1641 -3616 0 cellNo=997
rlabel pdiffusion 1648 -3616 1648 -3616 0 feedthrough
rlabel pdiffusion 3 -3627 3 -3627 0 cellNo=1366
rlabel pdiffusion 10 -3627 10 -3627 0 cellNo=1367
rlabel pdiffusion 17 -3627 17 -3627 0 cellNo=1368
rlabel pdiffusion 24 -3627 24 -3627 0 cellNo=1369
rlabel pdiffusion 31 -3627 31 -3627 0 cellNo=1370
rlabel pdiffusion 38 -3627 38 -3627 0 cellNo=1371
rlabel pdiffusion 45 -3627 45 -3627 0 cellNo=1372
rlabel pdiffusion 52 -3627 52 -3627 0 cellNo=1373
rlabel pdiffusion 59 -3627 59 -3627 0 cellNo=1374
rlabel pdiffusion 66 -3627 66 -3627 0 cellNo=1375
rlabel pdiffusion 73 -3627 73 -3627 0 cellNo=1376
rlabel pdiffusion 80 -3627 80 -3627 0 cellNo=1377
rlabel pdiffusion 87 -3627 87 -3627 0 cellNo=1378
rlabel pdiffusion 94 -3627 94 -3627 0 cellNo=1379
rlabel pdiffusion 101 -3627 101 -3627 0 cellNo=1380
rlabel pdiffusion 108 -3627 108 -3627 0 cellNo=1381
rlabel pdiffusion 115 -3627 115 -3627 0 cellNo=1382
rlabel pdiffusion 122 -3627 122 -3627 0 cellNo=1383
rlabel pdiffusion 129 -3627 129 -3627 0 cellNo=1384
rlabel pdiffusion 136 -3627 136 -3627 0 cellNo=1385
rlabel pdiffusion 143 -3627 143 -3627 0 cellNo=1386
rlabel pdiffusion 150 -3627 150 -3627 0 cellNo=1387
rlabel pdiffusion 157 -3627 157 -3627 0 cellNo=1388
rlabel pdiffusion 164 -3627 164 -3627 0 cellNo=1389
rlabel pdiffusion 171 -3627 171 -3627 0 cellNo=1390
rlabel pdiffusion 178 -3627 178 -3627 0 cellNo=1391
rlabel pdiffusion 185 -3627 185 -3627 0 cellNo=1432
rlabel pdiffusion 192 -3627 192 -3627 0 cellNo=1393
rlabel pdiffusion 199 -3627 199 -3627 0 cellNo=1394
rlabel pdiffusion 206 -3627 206 -3627 0 cellNo=1395
rlabel pdiffusion 213 -3627 213 -3627 0 cellNo=1435
rlabel pdiffusion 220 -3627 220 -3627 0 cellNo=1397
rlabel pdiffusion 227 -3627 227 -3627 0 cellNo=1398
rlabel pdiffusion 234 -3627 234 -3627 0 cellNo=1402
rlabel pdiffusion 395 -3627 395 -3627 0 feedthrough
rlabel pdiffusion 402 -3627 402 -3627 0 feedthrough
rlabel pdiffusion 605 -3627 605 -3627 0 feedthrough
rlabel pdiffusion 612 -3627 612 -3627 0 feedthrough
rlabel pdiffusion 696 -3627 696 -3627 0 feedthrough
rlabel pdiffusion 759 -3627 759 -3627 0 cellNo=876
rlabel pdiffusion 766 -3627 766 -3627 0 feedthrough
rlabel pdiffusion 3 -3638 3 -3638 0 cellNo=1204
rlabel pdiffusion 10 -3638 10 -3638 0 cellNo=1406
rlabel pdiffusion 17 -3638 17 -3638 0 cellNo=1407
rlabel pdiffusion 24 -3638 24 -3638 0 cellNo=1408
rlabel pdiffusion 31 -3638 31 -3638 0 cellNo=1409
rlabel pdiffusion 38 -3638 38 -3638 0 cellNo=1410
rlabel pdiffusion 45 -3638 45 -3638 0 cellNo=1411
rlabel pdiffusion 52 -3638 52 -3638 0 cellNo=1412
rlabel pdiffusion 59 -3638 59 -3638 0 cellNo=1413
rlabel pdiffusion 66 -3638 66 -3638 0 cellNo=1414
rlabel pdiffusion 73 -3638 73 -3638 0 cellNo=1415
rlabel pdiffusion 80 -3638 80 -3638 0 cellNo=1416
rlabel pdiffusion 87 -3638 87 -3638 0 cellNo=1417
rlabel pdiffusion 94 -3638 94 -3638 0 cellNo=1418
rlabel pdiffusion 101 -3638 101 -3638 0 cellNo=1419
rlabel pdiffusion 108 -3638 108 -3638 0 cellNo=1420
rlabel pdiffusion 115 -3638 115 -3638 0 cellNo=1421
rlabel pdiffusion 122 -3638 122 -3638 0 cellNo=1422
rlabel pdiffusion 129 -3638 129 -3638 0 cellNo=1423
rlabel pdiffusion 136 -3638 136 -3638 0 cellNo=1424
rlabel pdiffusion 143 -3638 143 -3638 0 cellNo=1425
rlabel pdiffusion 150 -3638 150 -3638 0 cellNo=1426
rlabel pdiffusion 157 -3638 157 -3638 0 cellNo=1427
rlabel pdiffusion 164 -3638 164 -3638 0 cellNo=1428
rlabel pdiffusion 171 -3638 171 -3638 0 cellNo=1429
rlabel pdiffusion 178 -3638 178 -3638 0 cellNo=1430
rlabel pdiffusion 185 -3638 185 -3638 0 cellNo=1431
rlabel pdiffusion 192 -3638 192 -3638 0 cellNo=1405
rlabel pdiffusion 199 -3638 199 -3638 0 cellNo=1433
rlabel pdiffusion 206 -3638 206 -3638 0 cellNo=1434
rlabel pdiffusion 213 -3638 213 -3638 0 cellNo=1357
rlabel pdiffusion 220 -3638 220 -3638 0 cellNo=1436
rlabel pdiffusion 227 -3638 227 -3638 0 cellNo=1437
rlabel pdiffusion 234 -3638 234 -3638 0 cellNo=1439
rlabel pdiffusion 395 -3638 395 -3638 0 feedthrough
rlabel pdiffusion 402 -3638 402 -3638 0 feedthrough
rlabel pdiffusion 605 -3638 605 -3638 0 feedthrough
rlabel pdiffusion 612 -3638 612 -3638 0 feedthrough
rlabel pdiffusion 696 -3638 696 -3638 0 feedthrough
rlabel pdiffusion 3 -3649 3 -3649 0 cellNo=1444
rlabel pdiffusion 10 -3649 10 -3649 0 cellNo=1445
rlabel pdiffusion 17 -3649 17 -3649 0 cellNo=1446
rlabel pdiffusion 24 -3649 24 -3649 0 cellNo=1447
rlabel pdiffusion 31 -3649 31 -3649 0 cellNo=1448
rlabel pdiffusion 38 -3649 38 -3649 0 cellNo=1449
rlabel pdiffusion 45 -3649 45 -3649 0 cellNo=1450
rlabel pdiffusion 52 -3649 52 -3649 0 cellNo=1451
rlabel pdiffusion 59 -3649 59 -3649 0 cellNo=1452
rlabel pdiffusion 66 -3649 66 -3649 0 cellNo=1453
rlabel pdiffusion 73 -3649 73 -3649 0 cellNo=1454
rlabel pdiffusion 80 -3649 80 -3649 0 cellNo=1455
rlabel pdiffusion 87 -3649 87 -3649 0 cellNo=1456
rlabel pdiffusion 94 -3649 94 -3649 0 cellNo=1457
rlabel pdiffusion 101 -3649 101 -3649 0 cellNo=1458
rlabel pdiffusion 108 -3649 108 -3649 0 cellNo=1459
rlabel pdiffusion 115 -3649 115 -3649 0 cellNo=1460
rlabel pdiffusion 122 -3649 122 -3649 0 cellNo=1461
rlabel pdiffusion 129 -3649 129 -3649 0 cellNo=1462
rlabel pdiffusion 136 -3649 136 -3649 0 cellNo=1463
rlabel pdiffusion 143 -3649 143 -3649 0 cellNo=1464
rlabel pdiffusion 150 -3649 150 -3649 0 cellNo=1465
rlabel pdiffusion 157 -3649 157 -3649 0 cellNo=1466
rlabel pdiffusion 164 -3649 164 -3649 0 cellNo=1467
rlabel pdiffusion 171 -3649 171 -3649 0 cellNo=1468
rlabel pdiffusion 178 -3649 178 -3649 0 cellNo=1469
rlabel pdiffusion 185 -3649 185 -3649 0 cellNo=1470
rlabel pdiffusion 192 -3649 192 -3649 0 cellNo=1471
rlabel pdiffusion 199 -3649 199 -3649 0 cellNo=1472
rlabel pdiffusion 206 -3649 206 -3649 0 cellNo=1473
rlabel pdiffusion 213 -3649 213 -3649 0 cellNo=1474
rlabel pdiffusion 220 -3649 220 -3649 0 cellNo=1475
rlabel pdiffusion 227 -3649 227 -3649 0 cellNo=1476
rlabel pdiffusion 234 -3649 234 -3649 0 cellNo=1477
rlabel pdiffusion 241 -3649 241 -3649 0 cellNo=1478
rlabel pdiffusion 248 -3649 248 -3649 0 cellNo=1479
rlabel pdiffusion 255 -3649 255 -3649 0 cellNo=1480
rlabel pdiffusion 262 -3649 262 -3649 0 cellNo=1481
rlabel pdiffusion 269 -3649 269 -3649 0 cellNo=1482
rlabel pdiffusion 395 -3649 395 -3649 0 feedthrough
rlabel pdiffusion 402 -3649 402 -3649 0 feedthrough
rlabel pdiffusion 605 -3649 605 -3649 0 feedthrough
rlabel pdiffusion 612 -3649 612 -3649 0 feedthrough
rlabel pdiffusion 696 -3649 696 -3649 0 feedthrough
rlabel pdiffusion 3 -3664 3 -3664 0 cellNo=1040
rlabel pdiffusion 10 -3664 10 -3664 0 cellNo=1484
rlabel pdiffusion 17 -3664 17 -3664 0 cellNo=1485
rlabel pdiffusion 24 -3664 24 -3664 0 cellNo=1486
rlabel pdiffusion 31 -3664 31 -3664 0 cellNo=1487
rlabel pdiffusion 38 -3664 38 -3664 0 cellNo=1488
rlabel pdiffusion 45 -3664 45 -3664 0 cellNo=1489
rlabel pdiffusion 52 -3664 52 -3664 0 cellNo=1490
rlabel pdiffusion 59 -3664 59 -3664 0 cellNo=1491
rlabel pdiffusion 66 -3664 66 -3664 0 cellNo=1492
rlabel pdiffusion 73 -3664 73 -3664 0 cellNo=1493
rlabel pdiffusion 80 -3664 80 -3664 0 cellNo=1494
rlabel pdiffusion 87 -3664 87 -3664 0 cellNo=1495
rlabel pdiffusion 94 -3664 94 -3664 0 cellNo=1496
rlabel pdiffusion 101 -3664 101 -3664 0 cellNo=1497
rlabel pdiffusion 108 -3664 108 -3664 0 cellNo=1498
rlabel pdiffusion 115 -3664 115 -3664 0 cellNo=1499
rlabel pdiffusion 122 -3664 122 -3664 0 cellNo=1500
rlabel pdiffusion 129 -3664 129 -3664 0 cellNo=1189
rlabel pdiffusion 136 -3664 136 -3664 0 cellNo=1483
rlabel pdiffusion 143 -3664 143 -3664 0 cellNo=1074
rlabel pdiffusion 150 -3664 150 -3664 0 cellNo=1051
rlabel pdiffusion 157 -3664 157 -3664 0 cellNo=1109
rlabel pdiffusion 164 -3664 164 -3664 0 cellNo=1165
rlabel pdiffusion 171 -3664 171 -3664 0 cellNo=1198
rlabel pdiffusion 178 -3664 178 -3664 0 cellNo=1244
rlabel pdiffusion 185 -3664 185 -3664 0 cellNo=1284
rlabel pdiffusion 192 -3664 192 -3664 0 cellNo=1324
rlabel pdiffusion 199 -3664 199 -3664 0 cellNo=1363
rlabel pdiffusion 206 -3664 206 -3664 0 cellNo=1401
rlabel pdiffusion 395 -3664 395 -3664 0 cellNo=822
rlabel pdiffusion 402 -3664 402 -3664 0 feedthrough
rlabel pdiffusion 605 -3664 605 -3664 0 feedthrough
rlabel pdiffusion 612 -3664 612 -3664 0 cellNo=524
rlabel pdiffusion 696 -3664 696 -3664 0 cellNo=893
rlabel polysilicon 212 -26 212 -26 0 3
rlabel polysilicon 254 -20 254 -20 0 1
rlabel polysilicon 254 -26 254 -26 0 3
rlabel polysilicon 352 -20 352 -20 0 1
rlabel polysilicon 352 -26 352 -26 0 3
rlabel polysilicon 397 -20 397 -20 0 2
rlabel polysilicon 397 -26 397 -26 0 4
rlabel polysilicon 415 -20 415 -20 0 1
rlabel polysilicon 422 -20 422 -20 0 1
rlabel polysilicon 422 -26 422 -26 0 3
rlabel polysilicon 432 -20 432 -20 0 2
rlabel polysilicon 432 -26 432 -26 0 4
rlabel polysilicon 446 -26 446 -26 0 4
rlabel polysilicon 485 -20 485 -20 0 1
rlabel polysilicon 485 -26 485 -26 0 3
rlabel polysilicon 548 -20 548 -20 0 1
rlabel polysilicon 548 -26 548 -26 0 3
rlabel polysilicon 555 -20 555 -20 0 1
rlabel polysilicon 572 -20 572 -20 0 2
rlabel polysilicon 569 -26 569 -26 0 3
rlabel polysilicon 572 -26 572 -26 0 4
rlabel polysilicon 576 -20 576 -20 0 1
rlabel polysilicon 576 -26 576 -26 0 3
rlabel polysilicon 583 -20 583 -20 0 1
rlabel polysilicon 583 -26 583 -26 0 3
rlabel polysilicon 604 -20 604 -20 0 1
rlabel polysilicon 604 -26 604 -26 0 3
rlabel polysilicon 611 -20 611 -20 0 1
rlabel polysilicon 611 -26 611 -26 0 3
rlabel polysilicon 618 -20 618 -20 0 1
rlabel polysilicon 618 -26 618 -26 0 3
rlabel polysilicon 625 -20 625 -20 0 1
rlabel polysilicon 625 -26 625 -26 0 3
rlabel polysilicon 632 -20 632 -20 0 1
rlabel polysilicon 635 -20 635 -20 0 2
rlabel polysilicon 639 -20 639 -20 0 1
rlabel polysilicon 639 -26 639 -26 0 3
rlabel polysilicon 646 -20 646 -20 0 1
rlabel polysilicon 646 -26 646 -26 0 3
rlabel polysilicon 653 -26 653 -26 0 3
rlabel polysilicon 656 -26 656 -26 0 4
rlabel polysilicon 663 -20 663 -20 0 2
rlabel polysilicon 660 -26 660 -26 0 3
rlabel polysilicon 681 -20 681 -20 0 1
rlabel polysilicon 681 -26 681 -26 0 3
rlabel polysilicon 688 -20 688 -20 0 1
rlabel polysilicon 688 -26 688 -26 0 3
rlabel polysilicon 705 -20 705 -20 0 2
rlabel polysilicon 702 -26 702 -26 0 3
rlabel polysilicon 709 -20 709 -20 0 1
rlabel polysilicon 709 -26 709 -26 0 3
rlabel polysilicon 716 -20 716 -20 0 1
rlabel polysilicon 716 -26 716 -26 0 3
rlabel polysilicon 730 -20 730 -20 0 1
rlabel polysilicon 730 -26 730 -26 0 3
rlabel polysilicon 765 -20 765 -20 0 1
rlabel polysilicon 768 -26 768 -26 0 4
rlabel polysilicon 772 -20 772 -20 0 1
rlabel polysilicon 772 -26 772 -26 0 3
rlabel polysilicon 796 -20 796 -20 0 2
rlabel polysilicon 800 -20 800 -20 0 1
rlabel polysilicon 803 -20 803 -20 0 2
rlabel polysilicon 810 -20 810 -20 0 2
rlabel polysilicon 807 -26 807 -26 0 3
rlabel polysilicon 810 -26 810 -26 0 4
rlabel polysilicon 814 -20 814 -20 0 1
rlabel polysilicon 814 -26 814 -26 0 3
rlabel polysilicon 821 -20 821 -20 0 1
rlabel polysilicon 824 -20 824 -20 0 2
rlabel polysilicon 828 -20 828 -20 0 1
rlabel polysilicon 828 -26 828 -26 0 3
rlabel polysilicon 835 -20 835 -20 0 1
rlabel polysilicon 835 -26 835 -26 0 3
rlabel polysilicon 842 -20 842 -20 0 1
rlabel polysilicon 845 -20 845 -20 0 2
rlabel polysilicon 842 -26 842 -26 0 3
rlabel polysilicon 852 -20 852 -20 0 2
rlabel polysilicon 849 -26 849 -26 0 3
rlabel polysilicon 859 -20 859 -20 0 2
rlabel polysilicon 863 -20 863 -20 0 1
rlabel polysilicon 863 -26 863 -26 0 3
rlabel polysilicon 870 -20 870 -20 0 1
rlabel polysilicon 870 -26 870 -26 0 3
rlabel polysilicon 884 -20 884 -20 0 1
rlabel polysilicon 887 -20 887 -20 0 2
rlabel polysilicon 887 -26 887 -26 0 4
rlabel polysilicon 891 -20 891 -20 0 1
rlabel polysilicon 891 -26 891 -26 0 3
rlabel polysilicon 898 -26 898 -26 0 3
rlabel polysilicon 915 -20 915 -20 0 2
rlabel polysilicon 912 -26 912 -26 0 3
rlabel polysilicon 915 -26 915 -26 0 4
rlabel polysilicon 919 -20 919 -20 0 1
rlabel polysilicon 919 -26 919 -26 0 3
rlabel polysilicon 961 -20 961 -20 0 1
rlabel polysilicon 961 -26 961 -26 0 3
rlabel polysilicon 968 -20 968 -20 0 1
rlabel polysilicon 968 -26 968 -26 0 3
rlabel polysilicon 978 -20 978 -20 0 2
rlabel polysilicon 978 -26 978 -26 0 4
rlabel polysilicon 982 -20 982 -20 0 1
rlabel polysilicon 982 -26 982 -26 0 3
rlabel polysilicon 989 -20 989 -20 0 1
rlabel polysilicon 989 -26 989 -26 0 3
rlabel polysilicon 1038 -20 1038 -20 0 1
rlabel polysilicon 1038 -26 1038 -26 0 3
rlabel polysilicon 1073 -20 1073 -20 0 1
rlabel polysilicon 1073 -26 1073 -26 0 3
rlabel polysilicon 1087 -20 1087 -20 0 1
rlabel polysilicon 1087 -26 1087 -26 0 3
rlabel polysilicon 1094 -20 1094 -20 0 1
rlabel polysilicon 1094 -26 1094 -26 0 3
rlabel polysilicon 1125 -20 1125 -20 0 2
rlabel polysilicon 1129 -20 1129 -20 0 1
rlabel polysilicon 1132 -26 1132 -26 0 4
rlabel polysilicon 1206 -20 1206 -20 0 1
rlabel polysilicon 1206 -26 1206 -26 0 3
rlabel polysilicon 1437 -20 1437 -20 0 1
rlabel polysilicon 1437 -26 1437 -26 0 3
rlabel polysilicon 1440 -26 1440 -26 0 4
rlabel polysilicon 1629 -26 1629 -26 0 4
rlabel polysilicon 184 -67 184 -67 0 1
rlabel polysilicon 184 -73 184 -73 0 3
rlabel polysilicon 198 -67 198 -67 0 1
rlabel polysilicon 198 -73 198 -73 0 3
rlabel polysilicon 240 -67 240 -67 0 1
rlabel polysilicon 240 -73 240 -73 0 3
rlabel polysilicon 275 -67 275 -67 0 1
rlabel polysilicon 275 -73 275 -73 0 3
rlabel polysilicon 296 -67 296 -67 0 1
rlabel polysilicon 296 -73 296 -73 0 3
rlabel polysilicon 313 -67 313 -67 0 2
rlabel polysilicon 310 -73 310 -73 0 3
rlabel polysilicon 317 -67 317 -67 0 1
rlabel polysilicon 317 -73 317 -73 0 3
rlabel polysilicon 355 -67 355 -67 0 2
rlabel polysilicon 352 -73 352 -73 0 3
rlabel polysilicon 394 -67 394 -67 0 1
rlabel polysilicon 394 -73 394 -73 0 3
rlabel polysilicon 404 -67 404 -67 0 2
rlabel polysilicon 401 -73 401 -73 0 3
rlabel polysilicon 404 -73 404 -73 0 4
rlabel polysilicon 408 -73 408 -73 0 3
rlabel polysilicon 411 -73 411 -73 0 4
rlabel polysilicon 415 -67 415 -67 0 1
rlabel polysilicon 415 -73 415 -73 0 3
rlabel polysilicon 422 -67 422 -67 0 1
rlabel polysilicon 422 -73 422 -73 0 3
rlabel polysilicon 464 -67 464 -67 0 1
rlabel polysilicon 464 -73 464 -73 0 3
rlabel polysilicon 471 -67 471 -67 0 1
rlabel polysilicon 471 -73 471 -73 0 3
rlabel polysilicon 478 -67 478 -67 0 1
rlabel polysilicon 478 -73 478 -73 0 3
rlabel polysilicon 485 -67 485 -67 0 1
rlabel polysilicon 485 -73 485 -73 0 3
rlabel polysilicon 492 -67 492 -67 0 1
rlabel polysilicon 492 -73 492 -73 0 3
rlabel polysilicon 499 -67 499 -67 0 1
rlabel polysilicon 499 -73 499 -73 0 3
rlabel polysilicon 506 -67 506 -67 0 1
rlabel polysilicon 506 -73 506 -73 0 3
rlabel polysilicon 520 -67 520 -67 0 1
rlabel polysilicon 520 -73 520 -73 0 3
rlabel polysilicon 534 -67 534 -67 0 1
rlabel polysilicon 534 -73 534 -73 0 3
rlabel polysilicon 541 -73 541 -73 0 3
rlabel polysilicon 544 -73 544 -73 0 4
rlabel polysilicon 548 -67 548 -67 0 1
rlabel polysilicon 548 -73 548 -73 0 3
rlabel polysilicon 565 -67 565 -67 0 2
rlabel polysilicon 565 -73 565 -73 0 4
rlabel polysilicon 569 -67 569 -67 0 1
rlabel polysilicon 569 -73 569 -73 0 3
rlabel polysilicon 583 -67 583 -67 0 1
rlabel polysilicon 583 -73 583 -73 0 3
rlabel polysilicon 590 -67 590 -67 0 1
rlabel polysilicon 590 -73 590 -73 0 3
rlabel polysilicon 597 -67 597 -67 0 1
rlabel polysilicon 597 -73 597 -73 0 3
rlabel polysilicon 604 -67 604 -67 0 1
rlabel polysilicon 604 -73 604 -73 0 3
rlabel polysilicon 611 -67 611 -67 0 1
rlabel polysilicon 611 -73 611 -73 0 3
rlabel polysilicon 618 -67 618 -67 0 1
rlabel polysilicon 618 -73 618 -73 0 3
rlabel polysilicon 639 -67 639 -67 0 1
rlabel polysilicon 639 -73 639 -73 0 3
rlabel polysilicon 646 -67 646 -67 0 1
rlabel polysilicon 646 -73 646 -73 0 3
rlabel polysilicon 653 -67 653 -67 0 1
rlabel polysilicon 656 -73 656 -73 0 4
rlabel polysilicon 660 -67 660 -67 0 1
rlabel polysilicon 660 -73 660 -73 0 3
rlabel polysilicon 667 -67 667 -67 0 1
rlabel polysilicon 667 -73 667 -73 0 3
rlabel polysilicon 674 -67 674 -67 0 1
rlabel polysilicon 677 -67 677 -67 0 2
rlabel polysilicon 677 -73 677 -73 0 4
rlabel polysilicon 681 -67 681 -67 0 1
rlabel polysilicon 681 -73 681 -73 0 3
rlabel polysilicon 688 -67 688 -67 0 1
rlabel polysilicon 688 -73 688 -73 0 3
rlabel polysilicon 695 -67 695 -67 0 1
rlabel polysilicon 702 -67 702 -67 0 1
rlabel polysilicon 702 -73 702 -73 0 3
rlabel polysilicon 709 -67 709 -67 0 1
rlabel polysilicon 709 -73 709 -73 0 3
rlabel polysilicon 716 -67 716 -67 0 1
rlabel polysilicon 716 -73 716 -73 0 3
rlabel polysilicon 723 -67 723 -67 0 1
rlabel polysilicon 723 -73 723 -73 0 3
rlabel polysilicon 730 -67 730 -67 0 1
rlabel polysilicon 730 -73 730 -73 0 3
rlabel polysilicon 737 -67 737 -67 0 1
rlabel polysilicon 740 -67 740 -67 0 2
rlabel polysilicon 744 -67 744 -67 0 1
rlabel polysilicon 744 -73 744 -73 0 3
rlabel polysilicon 751 -67 751 -67 0 1
rlabel polysilicon 751 -73 751 -73 0 3
rlabel polysilicon 758 -67 758 -67 0 1
rlabel polysilicon 758 -73 758 -73 0 3
rlabel polysilicon 765 -67 765 -67 0 1
rlabel polysilicon 765 -73 765 -73 0 3
rlabel polysilicon 772 -67 772 -67 0 1
rlabel polysilicon 772 -73 772 -73 0 3
rlabel polysilicon 779 -67 779 -67 0 1
rlabel polysilicon 779 -73 779 -73 0 3
rlabel polysilicon 789 -73 789 -73 0 4
rlabel polysilicon 793 -67 793 -67 0 1
rlabel polysilicon 793 -73 793 -73 0 3
rlabel polysilicon 800 -67 800 -67 0 1
rlabel polysilicon 803 -67 803 -67 0 2
rlabel polysilicon 800 -73 800 -73 0 3
rlabel polysilicon 807 -67 807 -67 0 1
rlabel polysilicon 807 -73 807 -73 0 3
rlabel polysilicon 814 -67 814 -67 0 1
rlabel polysilicon 814 -73 814 -73 0 3
rlabel polysilicon 821 -67 821 -67 0 1
rlabel polysilicon 821 -73 821 -73 0 3
rlabel polysilicon 828 -67 828 -67 0 1
rlabel polysilicon 828 -73 828 -73 0 3
rlabel polysilicon 835 -67 835 -67 0 1
rlabel polysilicon 835 -73 835 -73 0 3
rlabel polysilicon 842 -67 842 -67 0 1
rlabel polysilicon 842 -73 842 -73 0 3
rlabel polysilicon 849 -67 849 -67 0 1
rlabel polysilicon 852 -67 852 -67 0 2
rlabel polysilicon 852 -73 852 -73 0 4
rlabel polysilicon 856 -67 856 -67 0 1
rlabel polysilicon 856 -73 856 -73 0 3
rlabel polysilicon 859 -73 859 -73 0 4
rlabel polysilicon 863 -67 863 -67 0 1
rlabel polysilicon 863 -73 863 -73 0 3
rlabel polysilicon 870 -67 870 -67 0 1
rlabel polysilicon 870 -73 870 -73 0 3
rlabel polysilicon 877 -67 877 -67 0 1
rlabel polysilicon 877 -73 877 -73 0 3
rlabel polysilicon 884 -67 884 -67 0 1
rlabel polysilicon 887 -67 887 -67 0 2
rlabel polysilicon 891 -67 891 -67 0 1
rlabel polysilicon 891 -73 891 -73 0 3
rlabel polysilicon 901 -67 901 -67 0 2
rlabel polysilicon 898 -73 898 -73 0 3
rlabel polysilicon 908 -67 908 -67 0 2
rlabel polysilicon 908 -73 908 -73 0 4
rlabel polysilicon 912 -67 912 -67 0 1
rlabel polysilicon 912 -73 912 -73 0 3
rlabel polysilicon 919 -67 919 -67 0 1
rlabel polysilicon 919 -73 919 -73 0 3
rlabel polysilicon 926 -67 926 -67 0 1
rlabel polysilicon 926 -73 926 -73 0 3
rlabel polysilicon 933 -67 933 -67 0 1
rlabel polysilicon 933 -73 933 -73 0 3
rlabel polysilicon 940 -67 940 -67 0 1
rlabel polysilicon 943 -73 943 -73 0 4
rlabel polysilicon 947 -67 947 -67 0 1
rlabel polysilicon 947 -73 947 -73 0 3
rlabel polysilicon 954 -73 954 -73 0 3
rlabel polysilicon 957 -73 957 -73 0 4
rlabel polysilicon 961 -67 961 -67 0 1
rlabel polysilicon 961 -73 961 -73 0 3
rlabel polysilicon 968 -67 968 -67 0 1
rlabel polysilicon 968 -73 968 -73 0 3
rlabel polysilicon 975 -67 975 -67 0 1
rlabel polysilicon 975 -73 975 -73 0 3
rlabel polysilicon 982 -67 982 -67 0 1
rlabel polysilicon 982 -73 982 -73 0 3
rlabel polysilicon 989 -67 989 -67 0 1
rlabel polysilicon 989 -73 989 -73 0 3
rlabel polysilicon 996 -73 996 -73 0 3
rlabel polysilicon 999 -73 999 -73 0 4
rlabel polysilicon 1003 -67 1003 -67 0 1
rlabel polysilicon 1003 -73 1003 -73 0 3
rlabel polysilicon 1010 -67 1010 -67 0 1
rlabel polysilicon 1010 -73 1010 -73 0 3
rlabel polysilicon 1017 -67 1017 -67 0 1
rlabel polysilicon 1017 -73 1017 -73 0 3
rlabel polysilicon 1024 -67 1024 -67 0 1
rlabel polysilicon 1024 -73 1024 -73 0 3
rlabel polysilicon 1027 -73 1027 -73 0 4
rlabel polysilicon 1031 -67 1031 -67 0 1
rlabel polysilicon 1031 -73 1031 -73 0 3
rlabel polysilicon 1038 -67 1038 -67 0 1
rlabel polysilicon 1038 -73 1038 -73 0 3
rlabel polysilicon 1045 -67 1045 -67 0 1
rlabel polysilicon 1045 -73 1045 -73 0 3
rlabel polysilicon 1052 -67 1052 -67 0 1
rlabel polysilicon 1052 -73 1052 -73 0 3
rlabel polysilicon 1059 -67 1059 -67 0 1
rlabel polysilicon 1059 -73 1059 -73 0 3
rlabel polysilicon 1066 -67 1066 -67 0 1
rlabel polysilicon 1069 -67 1069 -67 0 2
rlabel polysilicon 1073 -67 1073 -67 0 1
rlabel polysilicon 1073 -73 1073 -73 0 3
rlabel polysilicon 1080 -67 1080 -67 0 1
rlabel polysilicon 1080 -73 1080 -73 0 3
rlabel polysilicon 1087 -67 1087 -67 0 1
rlabel polysilicon 1087 -73 1087 -73 0 3
rlabel polysilicon 1094 -67 1094 -67 0 1
rlabel polysilicon 1094 -73 1094 -73 0 3
rlabel polysilicon 1101 -67 1101 -67 0 1
rlabel polysilicon 1101 -73 1101 -73 0 3
rlabel polysilicon 1108 -67 1108 -67 0 1
rlabel polysilicon 1111 -73 1111 -73 0 4
rlabel polysilicon 1115 -67 1115 -67 0 1
rlabel polysilicon 1118 -73 1118 -73 0 4
rlabel polysilicon 1125 -67 1125 -67 0 2
rlabel polysilicon 1125 -73 1125 -73 0 4
rlabel polysilicon 1150 -67 1150 -67 0 1
rlabel polysilicon 1150 -73 1150 -73 0 3
rlabel polysilicon 1167 -73 1167 -73 0 4
rlabel polysilicon 1178 -67 1178 -67 0 1
rlabel polysilicon 1178 -73 1178 -73 0 3
rlabel polysilicon 1213 -67 1213 -67 0 1
rlabel polysilicon 1213 -73 1213 -73 0 3
rlabel polysilicon 1220 -67 1220 -67 0 1
rlabel polysilicon 1220 -73 1220 -73 0 3
rlabel polysilicon 1227 -73 1227 -73 0 3
rlabel polysilicon 1234 -67 1234 -67 0 1
rlabel polysilicon 1234 -73 1234 -73 0 3
rlabel polysilicon 1237 -73 1237 -73 0 4
rlabel polysilicon 1290 -67 1290 -67 0 1
rlabel polysilicon 1290 -73 1290 -73 0 3
rlabel polysilicon 1321 -67 1321 -67 0 2
rlabel polysilicon 1321 -73 1321 -73 0 4
rlabel polysilicon 1332 -67 1332 -67 0 1
rlabel polysilicon 1332 -73 1332 -73 0 3
rlabel polysilicon 1360 -67 1360 -67 0 1
rlabel polysilicon 1360 -73 1360 -73 0 3
rlabel polysilicon 1486 -67 1486 -67 0 1
rlabel polysilicon 1486 -73 1486 -73 0 3
rlabel polysilicon 1633 -67 1633 -67 0 1
rlabel polysilicon 1633 -73 1633 -73 0 3
rlabel polysilicon 1759 -67 1759 -67 0 1
rlabel polysilicon 1759 -73 1759 -73 0 3
rlabel polysilicon 58 -144 58 -144 0 1
rlabel polysilicon 58 -150 58 -150 0 3
rlabel polysilicon 65 -144 65 -144 0 1
rlabel polysilicon 65 -150 65 -150 0 3
rlabel polysilicon 72 -144 72 -144 0 1
rlabel polysilicon 72 -150 72 -150 0 3
rlabel polysilicon 79 -144 79 -144 0 1
rlabel polysilicon 79 -150 79 -150 0 3
rlabel polysilicon 86 -144 86 -144 0 1
rlabel polysilicon 86 -150 86 -150 0 3
rlabel polysilicon 93 -144 93 -144 0 1
rlabel polysilicon 93 -150 93 -150 0 3
rlabel polysilicon 100 -144 100 -144 0 1
rlabel polysilicon 100 -150 100 -150 0 3
rlabel polysilicon 107 -144 107 -144 0 1
rlabel polysilicon 107 -150 107 -150 0 3
rlabel polysilicon 114 -144 114 -144 0 1
rlabel polysilicon 114 -150 114 -150 0 3
rlabel polysilicon 121 -144 121 -144 0 1
rlabel polysilicon 124 -144 124 -144 0 2
rlabel polysilicon 124 -150 124 -150 0 4
rlabel polysilicon 128 -144 128 -144 0 1
rlabel polysilicon 128 -150 128 -150 0 3
rlabel polysilicon 135 -144 135 -144 0 1
rlabel polysilicon 135 -150 135 -150 0 3
rlabel polysilicon 142 -144 142 -144 0 1
rlabel polysilicon 145 -150 145 -150 0 4
rlabel polysilicon 149 -144 149 -144 0 1
rlabel polysilicon 152 -144 152 -144 0 2
rlabel polysilicon 152 -150 152 -150 0 4
rlabel polysilicon 156 -144 156 -144 0 1
rlabel polysilicon 156 -150 156 -150 0 3
rlabel polysilicon 163 -144 163 -144 0 1
rlabel polysilicon 163 -150 163 -150 0 3
rlabel polysilicon 170 -144 170 -144 0 1
rlabel polysilicon 170 -150 170 -150 0 3
rlabel polysilicon 177 -144 177 -144 0 1
rlabel polysilicon 177 -150 177 -150 0 3
rlabel polysilicon 184 -144 184 -144 0 1
rlabel polysilicon 184 -150 184 -150 0 3
rlabel polysilicon 191 -144 191 -144 0 1
rlabel polysilicon 191 -150 191 -150 0 3
rlabel polysilicon 198 -144 198 -144 0 1
rlabel polysilicon 198 -150 198 -150 0 3
rlabel polysilicon 205 -144 205 -144 0 1
rlabel polysilicon 205 -150 205 -150 0 3
rlabel polysilicon 212 -144 212 -144 0 1
rlabel polysilicon 212 -150 212 -150 0 3
rlabel polysilicon 219 -144 219 -144 0 1
rlabel polysilicon 219 -150 219 -150 0 3
rlabel polysilicon 226 -144 226 -144 0 1
rlabel polysilicon 229 -144 229 -144 0 2
rlabel polysilicon 226 -150 226 -150 0 3
rlabel polysilicon 233 -144 233 -144 0 1
rlabel polysilicon 236 -144 236 -144 0 2
rlabel polysilicon 240 -144 240 -144 0 1
rlabel polysilicon 240 -150 240 -150 0 3
rlabel polysilicon 247 -144 247 -144 0 1
rlabel polysilicon 247 -150 247 -150 0 3
rlabel polysilicon 254 -150 254 -150 0 3
rlabel polysilicon 257 -150 257 -150 0 4
rlabel polysilicon 261 -144 261 -144 0 1
rlabel polysilicon 264 -144 264 -144 0 2
rlabel polysilicon 261 -150 261 -150 0 3
rlabel polysilicon 268 -150 268 -150 0 3
rlabel polysilicon 275 -144 275 -144 0 1
rlabel polysilicon 275 -150 275 -150 0 3
rlabel polysilicon 282 -144 282 -144 0 1
rlabel polysilicon 282 -150 282 -150 0 3
rlabel polysilicon 289 -144 289 -144 0 1
rlabel polysilicon 289 -150 289 -150 0 3
rlabel polysilicon 296 -144 296 -144 0 1
rlabel polysilicon 296 -150 296 -150 0 3
rlabel polysilicon 303 -144 303 -144 0 1
rlabel polysilicon 303 -150 303 -150 0 3
rlabel polysilicon 310 -144 310 -144 0 1
rlabel polysilicon 310 -150 310 -150 0 3
rlabel polysilicon 317 -144 317 -144 0 1
rlabel polysilicon 317 -150 317 -150 0 3
rlabel polysilicon 324 -144 324 -144 0 1
rlabel polysilicon 324 -150 324 -150 0 3
rlabel polysilicon 331 -144 331 -144 0 1
rlabel polysilicon 331 -150 331 -150 0 3
rlabel polysilicon 338 -144 338 -144 0 1
rlabel polysilicon 338 -150 338 -150 0 3
rlabel polysilicon 345 -144 345 -144 0 1
rlabel polysilicon 345 -150 345 -150 0 3
rlabel polysilicon 352 -144 352 -144 0 1
rlabel polysilicon 352 -150 352 -150 0 3
rlabel polysilicon 359 -144 359 -144 0 1
rlabel polysilicon 359 -150 359 -150 0 3
rlabel polysilicon 366 -144 366 -144 0 1
rlabel polysilicon 366 -150 366 -150 0 3
rlabel polysilicon 373 -144 373 -144 0 1
rlabel polysilicon 373 -150 373 -150 0 3
rlabel polysilicon 380 -144 380 -144 0 1
rlabel polysilicon 380 -150 380 -150 0 3
rlabel polysilicon 387 -144 387 -144 0 1
rlabel polysilicon 390 -144 390 -144 0 2
rlabel polysilicon 390 -150 390 -150 0 4
rlabel polysilicon 394 -144 394 -144 0 1
rlabel polysilicon 394 -150 394 -150 0 3
rlabel polysilicon 401 -144 401 -144 0 1
rlabel polysilicon 401 -150 401 -150 0 3
rlabel polysilicon 408 -144 408 -144 0 1
rlabel polysilicon 408 -150 408 -150 0 3
rlabel polysilicon 415 -144 415 -144 0 1
rlabel polysilicon 415 -150 415 -150 0 3
rlabel polysilicon 422 -144 422 -144 0 1
rlabel polysilicon 422 -150 422 -150 0 3
rlabel polysilicon 429 -144 429 -144 0 1
rlabel polysilicon 429 -150 429 -150 0 3
rlabel polysilicon 436 -144 436 -144 0 1
rlabel polysilicon 436 -150 436 -150 0 3
rlabel polysilicon 443 -144 443 -144 0 1
rlabel polysilicon 446 -144 446 -144 0 2
rlabel polysilicon 450 -144 450 -144 0 1
rlabel polysilicon 450 -150 450 -150 0 3
rlabel polysilicon 457 -144 457 -144 0 1
rlabel polysilicon 460 -144 460 -144 0 2
rlabel polysilicon 460 -150 460 -150 0 4
rlabel polysilicon 467 -144 467 -144 0 2
rlabel polysilicon 467 -150 467 -150 0 4
rlabel polysilicon 471 -144 471 -144 0 1
rlabel polysilicon 474 -144 474 -144 0 2
rlabel polysilicon 478 -144 478 -144 0 1
rlabel polysilicon 478 -150 478 -150 0 3
rlabel polysilicon 485 -144 485 -144 0 1
rlabel polysilicon 485 -150 485 -150 0 3
rlabel polysilicon 492 -144 492 -144 0 1
rlabel polysilicon 492 -150 492 -150 0 3
rlabel polysilicon 499 -144 499 -144 0 1
rlabel polysilicon 499 -150 499 -150 0 3
rlabel polysilicon 506 -144 506 -144 0 1
rlabel polysilicon 506 -150 506 -150 0 3
rlabel polysilicon 513 -144 513 -144 0 1
rlabel polysilicon 513 -150 513 -150 0 3
rlabel polysilicon 523 -144 523 -144 0 2
rlabel polysilicon 520 -150 520 -150 0 3
rlabel polysilicon 523 -150 523 -150 0 4
rlabel polysilicon 527 -144 527 -144 0 1
rlabel polysilicon 530 -144 530 -144 0 2
rlabel polysilicon 527 -150 527 -150 0 3
rlabel polysilicon 530 -150 530 -150 0 4
rlabel polysilicon 534 -144 534 -144 0 1
rlabel polysilicon 534 -150 534 -150 0 3
rlabel polysilicon 541 -144 541 -144 0 1
rlabel polysilicon 541 -150 541 -150 0 3
rlabel polysilicon 548 -144 548 -144 0 1
rlabel polysilicon 548 -150 548 -150 0 3
rlabel polysilicon 555 -144 555 -144 0 1
rlabel polysilicon 555 -150 555 -150 0 3
rlabel polysilicon 562 -144 562 -144 0 1
rlabel polysilicon 565 -144 565 -144 0 2
rlabel polysilicon 565 -150 565 -150 0 4
rlabel polysilicon 569 -144 569 -144 0 1
rlabel polysilicon 569 -150 569 -150 0 3
rlabel polysilicon 576 -144 576 -144 0 1
rlabel polysilicon 576 -150 576 -150 0 3
rlabel polysilicon 583 -144 583 -144 0 1
rlabel polysilicon 583 -150 583 -150 0 3
rlabel polysilicon 590 -144 590 -144 0 1
rlabel polysilicon 590 -150 590 -150 0 3
rlabel polysilicon 597 -144 597 -144 0 1
rlabel polysilicon 600 -144 600 -144 0 2
rlabel polysilicon 600 -150 600 -150 0 4
rlabel polysilicon 604 -144 604 -144 0 1
rlabel polysilicon 604 -150 604 -150 0 3
rlabel polysilicon 611 -144 611 -144 0 1
rlabel polysilicon 611 -150 611 -150 0 3
rlabel polysilicon 618 -144 618 -144 0 1
rlabel polysilicon 618 -150 618 -150 0 3
rlabel polysilicon 625 -144 625 -144 0 1
rlabel polysilicon 625 -150 625 -150 0 3
rlabel polysilicon 632 -144 632 -144 0 1
rlabel polysilicon 632 -150 632 -150 0 3
rlabel polysilicon 639 -144 639 -144 0 1
rlabel polysilicon 639 -150 639 -150 0 3
rlabel polysilicon 649 -144 649 -144 0 2
rlabel polysilicon 649 -150 649 -150 0 4
rlabel polysilicon 653 -144 653 -144 0 1
rlabel polysilicon 653 -150 653 -150 0 3
rlabel polysilicon 660 -144 660 -144 0 1
rlabel polysilicon 660 -150 660 -150 0 3
rlabel polysilicon 667 -144 667 -144 0 1
rlabel polysilicon 667 -150 667 -150 0 3
rlabel polysilicon 674 -144 674 -144 0 1
rlabel polysilicon 674 -150 674 -150 0 3
rlabel polysilicon 681 -144 681 -144 0 1
rlabel polysilicon 684 -150 684 -150 0 4
rlabel polysilicon 688 -144 688 -144 0 1
rlabel polysilicon 688 -150 688 -150 0 3
rlabel polysilicon 698 -144 698 -144 0 2
rlabel polysilicon 695 -150 695 -150 0 3
rlabel polysilicon 698 -150 698 -150 0 4
rlabel polysilicon 702 -144 702 -144 0 1
rlabel polysilicon 702 -150 702 -150 0 3
rlabel polysilicon 709 -144 709 -144 0 1
rlabel polysilicon 709 -150 709 -150 0 3
rlabel polysilicon 716 -144 716 -144 0 1
rlabel polysilicon 716 -150 716 -150 0 3
rlabel polysilicon 723 -144 723 -144 0 1
rlabel polysilicon 723 -150 723 -150 0 3
rlabel polysilicon 730 -144 730 -144 0 1
rlabel polysilicon 733 -150 733 -150 0 4
rlabel polysilicon 737 -144 737 -144 0 1
rlabel polysilicon 740 -144 740 -144 0 2
rlabel polysilicon 737 -150 737 -150 0 3
rlabel polysilicon 744 -144 744 -144 0 1
rlabel polysilicon 744 -150 744 -150 0 3
rlabel polysilicon 751 -144 751 -144 0 1
rlabel polysilicon 751 -150 751 -150 0 3
rlabel polysilicon 758 -144 758 -144 0 1
rlabel polysilicon 758 -150 758 -150 0 3
rlabel polysilicon 765 -144 765 -144 0 1
rlabel polysilicon 765 -150 765 -150 0 3
rlabel polysilicon 768 -150 768 -150 0 4
rlabel polysilicon 772 -144 772 -144 0 1
rlabel polysilicon 772 -150 772 -150 0 3
rlabel polysilicon 779 -144 779 -144 0 1
rlabel polysilicon 779 -150 779 -150 0 3
rlabel polysilicon 786 -144 786 -144 0 1
rlabel polysilicon 786 -150 786 -150 0 3
rlabel polysilicon 793 -144 793 -144 0 1
rlabel polysilicon 793 -150 793 -150 0 3
rlabel polysilicon 803 -144 803 -144 0 2
rlabel polysilicon 800 -150 800 -150 0 3
rlabel polysilicon 803 -150 803 -150 0 4
rlabel polysilicon 807 -144 807 -144 0 1
rlabel polysilicon 807 -150 807 -150 0 3
rlabel polysilicon 814 -144 814 -144 0 1
rlabel polysilicon 814 -150 814 -150 0 3
rlabel polysilicon 821 -144 821 -144 0 1
rlabel polysilicon 821 -150 821 -150 0 3
rlabel polysilicon 828 -144 828 -144 0 1
rlabel polysilicon 828 -150 828 -150 0 3
rlabel polysilicon 835 -144 835 -144 0 1
rlabel polysilicon 835 -150 835 -150 0 3
rlabel polysilicon 838 -150 838 -150 0 4
rlabel polysilicon 842 -144 842 -144 0 1
rlabel polysilicon 842 -150 842 -150 0 3
rlabel polysilicon 849 -144 849 -144 0 1
rlabel polysilicon 849 -150 849 -150 0 3
rlabel polysilicon 856 -144 856 -144 0 1
rlabel polysilicon 856 -150 856 -150 0 3
rlabel polysilicon 863 -144 863 -144 0 1
rlabel polysilicon 863 -150 863 -150 0 3
rlabel polysilicon 870 -144 870 -144 0 1
rlabel polysilicon 870 -150 870 -150 0 3
rlabel polysilicon 877 -144 877 -144 0 1
rlabel polysilicon 877 -150 877 -150 0 3
rlabel polysilicon 884 -144 884 -144 0 1
rlabel polysilicon 884 -150 884 -150 0 3
rlabel polysilicon 891 -144 891 -144 0 1
rlabel polysilicon 891 -150 891 -150 0 3
rlabel polysilicon 898 -144 898 -144 0 1
rlabel polysilicon 898 -150 898 -150 0 3
rlabel polysilicon 905 -144 905 -144 0 1
rlabel polysilicon 905 -150 905 -150 0 3
rlabel polysilicon 912 -144 912 -144 0 1
rlabel polysilicon 912 -150 912 -150 0 3
rlabel polysilicon 919 -144 919 -144 0 1
rlabel polysilicon 919 -150 919 -150 0 3
rlabel polysilicon 929 -150 929 -150 0 4
rlabel polysilicon 933 -144 933 -144 0 1
rlabel polysilicon 936 -150 936 -150 0 4
rlabel polysilicon 940 -144 940 -144 0 1
rlabel polysilicon 940 -150 940 -150 0 3
rlabel polysilicon 947 -144 947 -144 0 1
rlabel polysilicon 947 -150 947 -150 0 3
rlabel polysilicon 950 -150 950 -150 0 4
rlabel polysilicon 954 -144 954 -144 0 1
rlabel polysilicon 954 -150 954 -150 0 3
rlabel polysilicon 961 -150 961 -150 0 3
rlabel polysilicon 968 -144 968 -144 0 1
rlabel polysilicon 968 -150 968 -150 0 3
rlabel polysilicon 975 -144 975 -144 0 1
rlabel polysilicon 975 -150 975 -150 0 3
rlabel polysilicon 982 -144 982 -144 0 1
rlabel polysilicon 982 -150 982 -150 0 3
rlabel polysilicon 989 -144 989 -144 0 1
rlabel polysilicon 989 -150 989 -150 0 3
rlabel polysilicon 996 -144 996 -144 0 1
rlabel polysilicon 996 -150 996 -150 0 3
rlabel polysilicon 1003 -144 1003 -144 0 1
rlabel polysilicon 1003 -150 1003 -150 0 3
rlabel polysilicon 1010 -144 1010 -144 0 1
rlabel polysilicon 1010 -150 1010 -150 0 3
rlabel polysilicon 1017 -144 1017 -144 0 1
rlabel polysilicon 1017 -150 1017 -150 0 3
rlabel polysilicon 1024 -144 1024 -144 0 1
rlabel polysilicon 1024 -150 1024 -150 0 3
rlabel polysilicon 1031 -144 1031 -144 0 1
rlabel polysilicon 1031 -150 1031 -150 0 3
rlabel polysilicon 1038 -144 1038 -144 0 1
rlabel polysilicon 1038 -150 1038 -150 0 3
rlabel polysilicon 1045 -144 1045 -144 0 1
rlabel polysilicon 1045 -150 1045 -150 0 3
rlabel polysilicon 1052 -144 1052 -144 0 1
rlabel polysilicon 1052 -150 1052 -150 0 3
rlabel polysilicon 1059 -144 1059 -144 0 1
rlabel polysilicon 1059 -150 1059 -150 0 3
rlabel polysilicon 1066 -144 1066 -144 0 1
rlabel polysilicon 1066 -150 1066 -150 0 3
rlabel polysilicon 1076 -144 1076 -144 0 2
rlabel polysilicon 1073 -150 1073 -150 0 3
rlabel polysilicon 1076 -150 1076 -150 0 4
rlabel polysilicon 1080 -144 1080 -144 0 1
rlabel polysilicon 1080 -150 1080 -150 0 3
rlabel polysilicon 1087 -144 1087 -144 0 1
rlabel polysilicon 1087 -150 1087 -150 0 3
rlabel polysilicon 1090 -150 1090 -150 0 4
rlabel polysilicon 1094 -144 1094 -144 0 1
rlabel polysilicon 1094 -150 1094 -150 0 3
rlabel polysilicon 1101 -144 1101 -144 0 1
rlabel polysilicon 1101 -150 1101 -150 0 3
rlabel polysilicon 1108 -144 1108 -144 0 1
rlabel polysilicon 1108 -150 1108 -150 0 3
rlabel polysilicon 1115 -144 1115 -144 0 1
rlabel polysilicon 1115 -150 1115 -150 0 3
rlabel polysilicon 1122 -144 1122 -144 0 1
rlabel polysilicon 1122 -150 1122 -150 0 3
rlabel polysilicon 1129 -144 1129 -144 0 1
rlabel polysilicon 1129 -150 1129 -150 0 3
rlabel polysilicon 1136 -144 1136 -144 0 1
rlabel polysilicon 1136 -150 1136 -150 0 3
rlabel polysilicon 1143 -144 1143 -144 0 1
rlabel polysilicon 1143 -150 1143 -150 0 3
rlabel polysilicon 1146 -150 1146 -150 0 4
rlabel polysilicon 1150 -144 1150 -144 0 1
rlabel polysilicon 1150 -150 1150 -150 0 3
rlabel polysilicon 1157 -144 1157 -144 0 1
rlabel polysilicon 1157 -150 1157 -150 0 3
rlabel polysilicon 1164 -144 1164 -144 0 1
rlabel polysilicon 1164 -150 1164 -150 0 3
rlabel polysilicon 1171 -144 1171 -144 0 1
rlabel polysilicon 1171 -150 1171 -150 0 3
rlabel polysilicon 1174 -150 1174 -150 0 4
rlabel polysilicon 1178 -144 1178 -144 0 1
rlabel polysilicon 1178 -150 1178 -150 0 3
rlabel polysilicon 1185 -144 1185 -144 0 1
rlabel polysilicon 1185 -150 1185 -150 0 3
rlabel polysilicon 1192 -144 1192 -144 0 1
rlabel polysilicon 1192 -150 1192 -150 0 3
rlabel polysilicon 1199 -144 1199 -144 0 1
rlabel polysilicon 1199 -150 1199 -150 0 3
rlabel polysilicon 1206 -144 1206 -144 0 1
rlabel polysilicon 1206 -150 1206 -150 0 3
rlabel polysilicon 1213 -144 1213 -144 0 1
rlabel polysilicon 1213 -150 1213 -150 0 3
rlabel polysilicon 1220 -144 1220 -144 0 1
rlabel polysilicon 1220 -150 1220 -150 0 3
rlabel polysilicon 1227 -144 1227 -144 0 1
rlabel polysilicon 1227 -150 1227 -150 0 3
rlabel polysilicon 1234 -144 1234 -144 0 1
rlabel polysilicon 1234 -150 1234 -150 0 3
rlabel polysilicon 1241 -144 1241 -144 0 1
rlabel polysilicon 1241 -150 1241 -150 0 3
rlabel polysilicon 1248 -144 1248 -144 0 1
rlabel polysilicon 1248 -150 1248 -150 0 3
rlabel polysilicon 1255 -144 1255 -144 0 1
rlabel polysilicon 1255 -150 1255 -150 0 3
rlabel polysilicon 1262 -150 1262 -150 0 3
rlabel polysilicon 1265 -150 1265 -150 0 4
rlabel polysilicon 1269 -144 1269 -144 0 1
rlabel polysilicon 1269 -150 1269 -150 0 3
rlabel polysilicon 1276 -144 1276 -144 0 1
rlabel polysilicon 1276 -150 1276 -150 0 3
rlabel polysilicon 1283 -144 1283 -144 0 1
rlabel polysilicon 1283 -150 1283 -150 0 3
rlabel polysilicon 1290 -144 1290 -144 0 1
rlabel polysilicon 1290 -150 1290 -150 0 3
rlabel polysilicon 1297 -144 1297 -144 0 1
rlabel polysilicon 1297 -150 1297 -150 0 3
rlabel polysilicon 1304 -144 1304 -144 0 1
rlabel polysilicon 1304 -150 1304 -150 0 3
rlabel polysilicon 1311 -144 1311 -144 0 1
rlabel polysilicon 1311 -150 1311 -150 0 3
rlabel polysilicon 1318 -144 1318 -144 0 1
rlabel polysilicon 1318 -150 1318 -150 0 3
rlabel polysilicon 1325 -144 1325 -144 0 1
rlabel polysilicon 1325 -150 1325 -150 0 3
rlabel polysilicon 1353 -144 1353 -144 0 1
rlabel polysilicon 1353 -150 1353 -150 0 3
rlabel polysilicon 1360 -144 1360 -144 0 1
rlabel polysilicon 1360 -150 1360 -150 0 3
rlabel polysilicon 1374 -144 1374 -144 0 1
rlabel polysilicon 1374 -150 1374 -150 0 3
rlabel polysilicon 1423 -144 1423 -144 0 1
rlabel polysilicon 1423 -150 1423 -150 0 3
rlabel polysilicon 1507 -144 1507 -144 0 1
rlabel polysilicon 1507 -150 1507 -150 0 3
rlabel polysilicon 1514 -144 1514 -144 0 1
rlabel polysilicon 1514 -150 1514 -150 0 3
rlabel polysilicon 1640 -144 1640 -144 0 1
rlabel polysilicon 1640 -150 1640 -150 0 3
rlabel polysilicon 1885 -144 1885 -144 0 1
rlabel polysilicon 1885 -150 1885 -150 0 3
rlabel polysilicon 16 -247 16 -247 0 1
rlabel polysilicon 16 -253 16 -253 0 3
rlabel polysilicon 23 -247 23 -247 0 1
rlabel polysilicon 23 -253 23 -253 0 3
rlabel polysilicon 30 -247 30 -247 0 1
rlabel polysilicon 30 -253 30 -253 0 3
rlabel polysilicon 37 -247 37 -247 0 1
rlabel polysilicon 37 -253 37 -253 0 3
rlabel polysilicon 44 -247 44 -247 0 1
rlabel polysilicon 44 -253 44 -253 0 3
rlabel polysilicon 51 -247 51 -247 0 1
rlabel polysilicon 51 -253 51 -253 0 3
rlabel polysilicon 58 -247 58 -247 0 1
rlabel polysilicon 58 -253 58 -253 0 3
rlabel polysilicon 72 -247 72 -247 0 1
rlabel polysilicon 72 -253 72 -253 0 3
rlabel polysilicon 79 -247 79 -247 0 1
rlabel polysilicon 79 -253 79 -253 0 3
rlabel polysilicon 89 -247 89 -247 0 2
rlabel polysilicon 89 -253 89 -253 0 4
rlabel polysilicon 93 -247 93 -247 0 1
rlabel polysilicon 93 -253 93 -253 0 3
rlabel polysilicon 100 -247 100 -247 0 1
rlabel polysilicon 100 -253 100 -253 0 3
rlabel polysilicon 107 -247 107 -247 0 1
rlabel polysilicon 107 -253 107 -253 0 3
rlabel polysilicon 117 -247 117 -247 0 2
rlabel polysilicon 117 -253 117 -253 0 4
rlabel polysilicon 121 -247 121 -247 0 1
rlabel polysilicon 121 -253 121 -253 0 3
rlabel polysilicon 128 -247 128 -247 0 1
rlabel polysilicon 128 -253 128 -253 0 3
rlabel polysilicon 135 -247 135 -247 0 1
rlabel polysilicon 135 -253 135 -253 0 3
rlabel polysilicon 138 -253 138 -253 0 4
rlabel polysilicon 142 -247 142 -247 0 1
rlabel polysilicon 142 -253 142 -253 0 3
rlabel polysilicon 149 -247 149 -247 0 1
rlabel polysilicon 149 -253 149 -253 0 3
rlabel polysilicon 156 -247 156 -247 0 1
rlabel polysilicon 159 -247 159 -247 0 2
rlabel polysilicon 156 -253 156 -253 0 3
rlabel polysilicon 163 -247 163 -247 0 1
rlabel polysilicon 163 -253 163 -253 0 3
rlabel polysilicon 170 -247 170 -247 0 1
rlabel polysilicon 170 -253 170 -253 0 3
rlabel polysilicon 177 -247 177 -247 0 1
rlabel polysilicon 177 -253 177 -253 0 3
rlabel polysilicon 184 -247 184 -247 0 1
rlabel polysilicon 184 -253 184 -253 0 3
rlabel polysilicon 194 -247 194 -247 0 2
rlabel polysilicon 194 -253 194 -253 0 4
rlabel polysilicon 198 -247 198 -247 0 1
rlabel polysilicon 201 -247 201 -247 0 2
rlabel polysilicon 205 -253 205 -253 0 3
rlabel polysilicon 208 -253 208 -253 0 4
rlabel polysilicon 212 -247 212 -247 0 1
rlabel polysilicon 212 -253 212 -253 0 3
rlabel polysilicon 219 -247 219 -247 0 1
rlabel polysilicon 219 -253 219 -253 0 3
rlabel polysilicon 226 -247 226 -247 0 1
rlabel polysilicon 226 -253 226 -253 0 3
rlabel polysilicon 233 -247 233 -247 0 1
rlabel polysilicon 233 -253 233 -253 0 3
rlabel polysilicon 240 -247 240 -247 0 1
rlabel polysilicon 243 -247 243 -247 0 2
rlabel polysilicon 240 -253 240 -253 0 3
rlabel polysilicon 247 -247 247 -247 0 1
rlabel polysilicon 247 -253 247 -253 0 3
rlabel polysilicon 254 -247 254 -247 0 1
rlabel polysilicon 254 -253 254 -253 0 3
rlabel polysilicon 261 -247 261 -247 0 1
rlabel polysilicon 261 -253 261 -253 0 3
rlabel polysilicon 271 -247 271 -247 0 2
rlabel polysilicon 268 -253 268 -253 0 3
rlabel polysilicon 271 -253 271 -253 0 4
rlabel polysilicon 275 -247 275 -247 0 1
rlabel polysilicon 275 -253 275 -253 0 3
rlabel polysilicon 282 -247 282 -247 0 1
rlabel polysilicon 282 -253 282 -253 0 3
rlabel polysilicon 289 -247 289 -247 0 1
rlabel polysilicon 289 -253 289 -253 0 3
rlabel polysilicon 296 -247 296 -247 0 1
rlabel polysilicon 299 -253 299 -253 0 4
rlabel polysilicon 303 -247 303 -247 0 1
rlabel polysilicon 303 -253 303 -253 0 3
rlabel polysilicon 310 -247 310 -247 0 1
rlabel polysilicon 310 -253 310 -253 0 3
rlabel polysilicon 313 -253 313 -253 0 4
rlabel polysilicon 317 -247 317 -247 0 1
rlabel polysilicon 317 -253 317 -253 0 3
rlabel polysilicon 324 -247 324 -247 0 1
rlabel polysilicon 324 -253 324 -253 0 3
rlabel polysilicon 331 -247 331 -247 0 1
rlabel polysilicon 331 -253 331 -253 0 3
rlabel polysilicon 338 -247 338 -247 0 1
rlabel polysilicon 338 -253 338 -253 0 3
rlabel polysilicon 345 -247 345 -247 0 1
rlabel polysilicon 345 -253 345 -253 0 3
rlabel polysilicon 352 -247 352 -247 0 1
rlabel polysilicon 352 -253 352 -253 0 3
rlabel polysilicon 359 -247 359 -247 0 1
rlabel polysilicon 359 -253 359 -253 0 3
rlabel polysilicon 366 -247 366 -247 0 1
rlabel polysilicon 366 -253 366 -253 0 3
rlabel polysilicon 373 -247 373 -247 0 1
rlabel polysilicon 373 -253 373 -253 0 3
rlabel polysilicon 380 -247 380 -247 0 1
rlabel polysilicon 380 -253 380 -253 0 3
rlabel polysilicon 387 -247 387 -247 0 1
rlabel polysilicon 387 -253 387 -253 0 3
rlabel polysilicon 394 -247 394 -247 0 1
rlabel polysilicon 394 -253 394 -253 0 3
rlabel polysilicon 401 -247 401 -247 0 1
rlabel polysilicon 401 -253 401 -253 0 3
rlabel polysilicon 408 -247 408 -247 0 1
rlabel polysilicon 408 -253 408 -253 0 3
rlabel polysilicon 415 -247 415 -247 0 1
rlabel polysilicon 415 -253 415 -253 0 3
rlabel polysilicon 422 -247 422 -247 0 1
rlabel polysilicon 422 -253 422 -253 0 3
rlabel polysilicon 429 -247 429 -247 0 1
rlabel polysilicon 429 -253 429 -253 0 3
rlabel polysilicon 436 -247 436 -247 0 1
rlabel polysilicon 439 -247 439 -247 0 2
rlabel polysilicon 436 -253 436 -253 0 3
rlabel polysilicon 439 -253 439 -253 0 4
rlabel polysilicon 443 -247 443 -247 0 1
rlabel polysilicon 443 -253 443 -253 0 3
rlabel polysilicon 450 -247 450 -247 0 1
rlabel polysilicon 450 -253 450 -253 0 3
rlabel polysilicon 457 -247 457 -247 0 1
rlabel polysilicon 457 -253 457 -253 0 3
rlabel polysilicon 464 -253 464 -253 0 3
rlabel polysilicon 467 -253 467 -253 0 4
rlabel polysilicon 471 -247 471 -247 0 1
rlabel polysilicon 471 -253 471 -253 0 3
rlabel polysilicon 478 -247 478 -247 0 1
rlabel polysilicon 478 -253 478 -253 0 3
rlabel polysilicon 485 -247 485 -247 0 1
rlabel polysilicon 485 -253 485 -253 0 3
rlabel polysilicon 492 -247 492 -247 0 1
rlabel polysilicon 492 -253 492 -253 0 3
rlabel polysilicon 499 -247 499 -247 0 1
rlabel polysilicon 499 -253 499 -253 0 3
rlabel polysilicon 506 -247 506 -247 0 1
rlabel polysilicon 506 -253 506 -253 0 3
rlabel polysilicon 513 -247 513 -247 0 1
rlabel polysilicon 513 -253 513 -253 0 3
rlabel polysilicon 520 -247 520 -247 0 1
rlabel polysilicon 523 -247 523 -247 0 2
rlabel polysilicon 523 -253 523 -253 0 4
rlabel polysilicon 527 -247 527 -247 0 1
rlabel polysilicon 527 -253 527 -253 0 3
rlabel polysilicon 534 -247 534 -247 0 1
rlabel polysilicon 537 -247 537 -247 0 2
rlabel polysilicon 534 -253 534 -253 0 3
rlabel polysilicon 537 -253 537 -253 0 4
rlabel polysilicon 541 -247 541 -247 0 1
rlabel polysilicon 541 -253 541 -253 0 3
rlabel polysilicon 548 -247 548 -247 0 1
rlabel polysilicon 548 -253 548 -253 0 3
rlabel polysilicon 555 -247 555 -247 0 1
rlabel polysilicon 555 -253 555 -253 0 3
rlabel polysilicon 562 -247 562 -247 0 1
rlabel polysilicon 562 -253 562 -253 0 3
rlabel polysilicon 569 -247 569 -247 0 1
rlabel polysilicon 569 -253 569 -253 0 3
rlabel polysilicon 576 -247 576 -247 0 1
rlabel polysilicon 576 -253 576 -253 0 3
rlabel polysilicon 583 -247 583 -247 0 1
rlabel polysilicon 583 -253 583 -253 0 3
rlabel polysilicon 593 -247 593 -247 0 2
rlabel polysilicon 590 -253 590 -253 0 3
rlabel polysilicon 597 -247 597 -247 0 1
rlabel polysilicon 597 -253 597 -253 0 3
rlabel polysilicon 604 -247 604 -247 0 1
rlabel polysilicon 604 -253 604 -253 0 3
rlabel polysilicon 611 -247 611 -247 0 1
rlabel polysilicon 611 -253 611 -253 0 3
rlabel polysilicon 621 -247 621 -247 0 2
rlabel polysilicon 618 -253 618 -253 0 3
rlabel polysilicon 621 -253 621 -253 0 4
rlabel polysilicon 625 -247 625 -247 0 1
rlabel polysilicon 625 -253 625 -253 0 3
rlabel polysilicon 632 -247 632 -247 0 1
rlabel polysilicon 632 -253 632 -253 0 3
rlabel polysilicon 639 -247 639 -247 0 1
rlabel polysilicon 639 -253 639 -253 0 3
rlabel polysilicon 646 -247 646 -247 0 1
rlabel polysilicon 646 -253 646 -253 0 3
rlabel polysilicon 653 -247 653 -247 0 1
rlabel polysilicon 653 -253 653 -253 0 3
rlabel polysilicon 660 -247 660 -247 0 1
rlabel polysilicon 660 -253 660 -253 0 3
rlabel polysilicon 667 -247 667 -247 0 1
rlabel polysilicon 667 -253 667 -253 0 3
rlabel polysilicon 674 -247 674 -247 0 1
rlabel polysilicon 674 -253 674 -253 0 3
rlabel polysilicon 681 -247 681 -247 0 1
rlabel polysilicon 681 -253 681 -253 0 3
rlabel polysilicon 688 -247 688 -247 0 1
rlabel polysilicon 688 -253 688 -253 0 3
rlabel polysilicon 695 -247 695 -247 0 1
rlabel polysilicon 695 -253 695 -253 0 3
rlabel polysilicon 705 -247 705 -247 0 2
rlabel polysilicon 702 -253 702 -253 0 3
rlabel polysilicon 705 -253 705 -253 0 4
rlabel polysilicon 709 -247 709 -247 0 1
rlabel polysilicon 712 -247 712 -247 0 2
rlabel polysilicon 709 -253 709 -253 0 3
rlabel polysilicon 712 -253 712 -253 0 4
rlabel polysilicon 716 -247 716 -247 0 1
rlabel polysilicon 716 -253 716 -253 0 3
rlabel polysilicon 723 -247 723 -247 0 1
rlabel polysilicon 723 -253 723 -253 0 3
rlabel polysilicon 730 -247 730 -247 0 1
rlabel polysilicon 730 -253 730 -253 0 3
rlabel polysilicon 737 -247 737 -247 0 1
rlabel polysilicon 737 -253 737 -253 0 3
rlabel polysilicon 744 -247 744 -247 0 1
rlabel polysilicon 744 -253 744 -253 0 3
rlabel polysilicon 751 -247 751 -247 0 1
rlabel polysilicon 751 -253 751 -253 0 3
rlabel polysilicon 758 -247 758 -247 0 1
rlabel polysilicon 758 -253 758 -253 0 3
rlabel polysilicon 765 -247 765 -247 0 1
rlabel polysilicon 765 -253 765 -253 0 3
rlabel polysilicon 772 -247 772 -247 0 1
rlabel polysilicon 772 -253 772 -253 0 3
rlabel polysilicon 779 -247 779 -247 0 1
rlabel polysilicon 779 -253 779 -253 0 3
rlabel polysilicon 786 -247 786 -247 0 1
rlabel polysilicon 786 -253 786 -253 0 3
rlabel polysilicon 793 -247 793 -247 0 1
rlabel polysilicon 793 -253 793 -253 0 3
rlabel polysilicon 800 -247 800 -247 0 1
rlabel polysilicon 800 -253 800 -253 0 3
rlabel polysilicon 807 -247 807 -247 0 1
rlabel polysilicon 807 -253 807 -253 0 3
rlabel polysilicon 814 -247 814 -247 0 1
rlabel polysilicon 814 -253 814 -253 0 3
rlabel polysilicon 821 -247 821 -247 0 1
rlabel polysilicon 821 -253 821 -253 0 3
rlabel polysilicon 828 -247 828 -247 0 1
rlabel polysilicon 828 -253 828 -253 0 3
rlabel polysilicon 835 -247 835 -247 0 1
rlabel polysilicon 835 -253 835 -253 0 3
rlabel polysilicon 842 -247 842 -247 0 1
rlabel polysilicon 842 -253 842 -253 0 3
rlabel polysilicon 849 -247 849 -247 0 1
rlabel polysilicon 849 -253 849 -253 0 3
rlabel polysilicon 856 -247 856 -247 0 1
rlabel polysilicon 856 -253 856 -253 0 3
rlabel polysilicon 863 -247 863 -247 0 1
rlabel polysilicon 863 -253 863 -253 0 3
rlabel polysilicon 870 -247 870 -247 0 1
rlabel polysilicon 870 -253 870 -253 0 3
rlabel polysilicon 877 -247 877 -247 0 1
rlabel polysilicon 877 -253 877 -253 0 3
rlabel polysilicon 884 -247 884 -247 0 1
rlabel polysilicon 887 -247 887 -247 0 2
rlabel polysilicon 887 -253 887 -253 0 4
rlabel polysilicon 894 -247 894 -247 0 2
rlabel polysilicon 894 -253 894 -253 0 4
rlabel polysilicon 898 -247 898 -247 0 1
rlabel polysilicon 898 -253 898 -253 0 3
rlabel polysilicon 905 -247 905 -247 0 1
rlabel polysilicon 905 -253 905 -253 0 3
rlabel polysilicon 915 -247 915 -247 0 2
rlabel polysilicon 912 -253 912 -253 0 3
rlabel polysilicon 915 -253 915 -253 0 4
rlabel polysilicon 919 -247 919 -247 0 1
rlabel polysilicon 919 -253 919 -253 0 3
rlabel polysilicon 926 -247 926 -247 0 1
rlabel polysilicon 926 -253 926 -253 0 3
rlabel polysilicon 933 -247 933 -247 0 1
rlabel polysilicon 933 -253 933 -253 0 3
rlabel polysilicon 940 -247 940 -247 0 1
rlabel polysilicon 940 -253 940 -253 0 3
rlabel polysilicon 947 -247 947 -247 0 1
rlabel polysilicon 947 -253 947 -253 0 3
rlabel polysilicon 954 -247 954 -247 0 1
rlabel polysilicon 954 -253 954 -253 0 3
rlabel polysilicon 961 -247 961 -247 0 1
rlabel polysilicon 961 -253 961 -253 0 3
rlabel polysilicon 968 -247 968 -247 0 1
rlabel polysilicon 968 -253 968 -253 0 3
rlabel polysilicon 975 -247 975 -247 0 1
rlabel polysilicon 975 -253 975 -253 0 3
rlabel polysilicon 982 -247 982 -247 0 1
rlabel polysilicon 982 -253 982 -253 0 3
rlabel polysilicon 989 -247 989 -247 0 1
rlabel polysilicon 992 -253 992 -253 0 4
rlabel polysilicon 999 -247 999 -247 0 2
rlabel polysilicon 996 -253 996 -253 0 3
rlabel polysilicon 1003 -247 1003 -247 0 1
rlabel polysilicon 1003 -253 1003 -253 0 3
rlabel polysilicon 1010 -247 1010 -247 0 1
rlabel polysilicon 1013 -247 1013 -247 0 2
rlabel polysilicon 1010 -253 1010 -253 0 3
rlabel polysilicon 1017 -247 1017 -247 0 1
rlabel polysilicon 1017 -253 1017 -253 0 3
rlabel polysilicon 1024 -247 1024 -247 0 1
rlabel polysilicon 1024 -253 1024 -253 0 3
rlabel polysilicon 1031 -247 1031 -247 0 1
rlabel polysilicon 1031 -253 1031 -253 0 3
rlabel polysilicon 1038 -247 1038 -247 0 1
rlabel polysilicon 1038 -253 1038 -253 0 3
rlabel polysilicon 1045 -247 1045 -247 0 1
rlabel polysilicon 1045 -253 1045 -253 0 3
rlabel polysilicon 1052 -247 1052 -247 0 1
rlabel polysilicon 1052 -253 1052 -253 0 3
rlabel polysilicon 1059 -247 1059 -247 0 1
rlabel polysilicon 1059 -253 1059 -253 0 3
rlabel polysilicon 1066 -247 1066 -247 0 1
rlabel polysilicon 1066 -253 1066 -253 0 3
rlabel polysilicon 1073 -247 1073 -247 0 1
rlabel polysilicon 1073 -253 1073 -253 0 3
rlabel polysilicon 1080 -247 1080 -247 0 1
rlabel polysilicon 1080 -253 1080 -253 0 3
rlabel polysilicon 1087 -247 1087 -247 0 1
rlabel polysilicon 1087 -253 1087 -253 0 3
rlabel polysilicon 1094 -247 1094 -247 0 1
rlabel polysilicon 1094 -253 1094 -253 0 3
rlabel polysilicon 1101 -247 1101 -247 0 1
rlabel polysilicon 1101 -253 1101 -253 0 3
rlabel polysilicon 1108 -247 1108 -247 0 1
rlabel polysilicon 1108 -253 1108 -253 0 3
rlabel polysilicon 1115 -247 1115 -247 0 1
rlabel polysilicon 1115 -253 1115 -253 0 3
rlabel polysilicon 1122 -247 1122 -247 0 1
rlabel polysilicon 1122 -253 1122 -253 0 3
rlabel polysilicon 1129 -247 1129 -247 0 1
rlabel polysilicon 1129 -253 1129 -253 0 3
rlabel polysilicon 1136 -247 1136 -247 0 1
rlabel polysilicon 1136 -253 1136 -253 0 3
rlabel polysilicon 1143 -247 1143 -247 0 1
rlabel polysilicon 1143 -253 1143 -253 0 3
rlabel polysilicon 1150 -247 1150 -247 0 1
rlabel polysilicon 1150 -253 1150 -253 0 3
rlabel polysilicon 1153 -253 1153 -253 0 4
rlabel polysilicon 1157 -247 1157 -247 0 1
rlabel polysilicon 1157 -253 1157 -253 0 3
rlabel polysilicon 1164 -247 1164 -247 0 1
rlabel polysilicon 1164 -253 1164 -253 0 3
rlabel polysilicon 1171 -247 1171 -247 0 1
rlabel polysilicon 1171 -253 1171 -253 0 3
rlabel polysilicon 1178 -247 1178 -247 0 1
rlabel polysilicon 1178 -253 1178 -253 0 3
rlabel polysilicon 1185 -247 1185 -247 0 1
rlabel polysilicon 1185 -253 1185 -253 0 3
rlabel polysilicon 1192 -247 1192 -247 0 1
rlabel polysilicon 1192 -253 1192 -253 0 3
rlabel polysilicon 1199 -247 1199 -247 0 1
rlabel polysilicon 1202 -247 1202 -247 0 2
rlabel polysilicon 1206 -247 1206 -247 0 1
rlabel polysilicon 1206 -253 1206 -253 0 3
rlabel polysilicon 1213 -247 1213 -247 0 1
rlabel polysilicon 1216 -247 1216 -247 0 2
rlabel polysilicon 1213 -253 1213 -253 0 3
rlabel polysilicon 1220 -247 1220 -247 0 1
rlabel polysilicon 1220 -253 1220 -253 0 3
rlabel polysilicon 1227 -247 1227 -247 0 1
rlabel polysilicon 1227 -253 1227 -253 0 3
rlabel polysilicon 1234 -247 1234 -247 0 1
rlabel polysilicon 1234 -253 1234 -253 0 3
rlabel polysilicon 1241 -247 1241 -247 0 1
rlabel polysilicon 1241 -253 1241 -253 0 3
rlabel polysilicon 1248 -247 1248 -247 0 1
rlabel polysilicon 1248 -253 1248 -253 0 3
rlabel polysilicon 1255 -247 1255 -247 0 1
rlabel polysilicon 1255 -253 1255 -253 0 3
rlabel polysilicon 1262 -247 1262 -247 0 1
rlabel polysilicon 1262 -253 1262 -253 0 3
rlabel polysilicon 1269 -247 1269 -247 0 1
rlabel polysilicon 1269 -253 1269 -253 0 3
rlabel polysilicon 1276 -247 1276 -247 0 1
rlabel polysilicon 1276 -253 1276 -253 0 3
rlabel polysilicon 1283 -247 1283 -247 0 1
rlabel polysilicon 1283 -253 1283 -253 0 3
rlabel polysilicon 1290 -247 1290 -247 0 1
rlabel polysilicon 1290 -253 1290 -253 0 3
rlabel polysilicon 1297 -247 1297 -247 0 1
rlabel polysilicon 1297 -253 1297 -253 0 3
rlabel polysilicon 1304 -247 1304 -247 0 1
rlabel polysilicon 1304 -253 1304 -253 0 3
rlabel polysilicon 1311 -247 1311 -247 0 1
rlabel polysilicon 1311 -253 1311 -253 0 3
rlabel polysilicon 1318 -247 1318 -247 0 1
rlabel polysilicon 1318 -253 1318 -253 0 3
rlabel polysilicon 1325 -247 1325 -247 0 1
rlabel polysilicon 1328 -247 1328 -247 0 2
rlabel polysilicon 1332 -247 1332 -247 0 1
rlabel polysilicon 1332 -253 1332 -253 0 3
rlabel polysilicon 1339 -247 1339 -247 0 1
rlabel polysilicon 1339 -253 1339 -253 0 3
rlabel polysilicon 1346 -247 1346 -247 0 1
rlabel polysilicon 1346 -253 1346 -253 0 3
rlabel polysilicon 1353 -247 1353 -247 0 1
rlabel polysilicon 1353 -253 1353 -253 0 3
rlabel polysilicon 1360 -247 1360 -247 0 1
rlabel polysilicon 1360 -253 1360 -253 0 3
rlabel polysilicon 1367 -247 1367 -247 0 1
rlabel polysilicon 1367 -253 1367 -253 0 3
rlabel polysilicon 1374 -247 1374 -247 0 1
rlabel polysilicon 1374 -253 1374 -253 0 3
rlabel polysilicon 1381 -247 1381 -247 0 1
rlabel polysilicon 1381 -253 1381 -253 0 3
rlabel polysilicon 1388 -247 1388 -247 0 1
rlabel polysilicon 1388 -253 1388 -253 0 3
rlabel polysilicon 1395 -247 1395 -247 0 1
rlabel polysilicon 1395 -253 1395 -253 0 3
rlabel polysilicon 1402 -247 1402 -247 0 1
rlabel polysilicon 1402 -253 1402 -253 0 3
rlabel polysilicon 1409 -247 1409 -247 0 1
rlabel polysilicon 1409 -253 1409 -253 0 3
rlabel polysilicon 1416 -247 1416 -247 0 1
rlabel polysilicon 1416 -253 1416 -253 0 3
rlabel polysilicon 1423 -247 1423 -247 0 1
rlabel polysilicon 1423 -253 1423 -253 0 3
rlabel polysilicon 1430 -247 1430 -247 0 1
rlabel polysilicon 1430 -253 1430 -253 0 3
rlabel polysilicon 1437 -247 1437 -247 0 1
rlabel polysilicon 1437 -253 1437 -253 0 3
rlabel polysilicon 1444 -247 1444 -247 0 1
rlabel polysilicon 1444 -253 1444 -253 0 3
rlabel polysilicon 1451 -247 1451 -247 0 1
rlabel polysilicon 1451 -253 1451 -253 0 3
rlabel polysilicon 1458 -247 1458 -247 0 1
rlabel polysilicon 1458 -253 1458 -253 0 3
rlabel polysilicon 1465 -247 1465 -247 0 1
rlabel polysilicon 1465 -253 1465 -253 0 3
rlabel polysilicon 1472 -247 1472 -247 0 1
rlabel polysilicon 1472 -253 1472 -253 0 3
rlabel polysilicon 1479 -247 1479 -247 0 1
rlabel polysilicon 1479 -253 1479 -253 0 3
rlabel polysilicon 1486 -247 1486 -247 0 1
rlabel polysilicon 1486 -253 1486 -253 0 3
rlabel polysilicon 1493 -247 1493 -247 0 1
rlabel polysilicon 1493 -253 1493 -253 0 3
rlabel polysilicon 1500 -247 1500 -247 0 1
rlabel polysilicon 1500 -253 1500 -253 0 3
rlabel polysilicon 1507 -247 1507 -247 0 1
rlabel polysilicon 1507 -253 1507 -253 0 3
rlabel polysilicon 1514 -247 1514 -247 0 1
rlabel polysilicon 1514 -253 1514 -253 0 3
rlabel polysilicon 1521 -247 1521 -247 0 1
rlabel polysilicon 1521 -253 1521 -253 0 3
rlabel polysilicon 1528 -247 1528 -247 0 1
rlabel polysilicon 1528 -253 1528 -253 0 3
rlabel polysilicon 1535 -247 1535 -247 0 1
rlabel polysilicon 1535 -253 1535 -253 0 3
rlabel polysilicon 1542 -247 1542 -247 0 1
rlabel polysilicon 1542 -253 1542 -253 0 3
rlabel polysilicon 1545 -253 1545 -253 0 4
rlabel polysilicon 1549 -247 1549 -247 0 1
rlabel polysilicon 1552 -253 1552 -253 0 4
rlabel polysilicon 1556 -247 1556 -247 0 1
rlabel polysilicon 1556 -253 1556 -253 0 3
rlabel polysilicon 1566 -247 1566 -247 0 2
rlabel polysilicon 1563 -253 1563 -253 0 3
rlabel polysilicon 1570 -247 1570 -247 0 1
rlabel polysilicon 1570 -253 1570 -253 0 3
rlabel polysilicon 1577 -247 1577 -247 0 1
rlabel polysilicon 1577 -253 1577 -253 0 3
rlabel polysilicon 1584 -247 1584 -247 0 1
rlabel polysilicon 1584 -253 1584 -253 0 3
rlabel polysilicon 1591 -247 1591 -247 0 1
rlabel polysilicon 1591 -253 1591 -253 0 3
rlabel polysilicon 1612 -247 1612 -247 0 1
rlabel polysilicon 1615 -247 1615 -247 0 2
rlabel polysilicon 1612 -253 1612 -253 0 3
rlabel polysilicon 1626 -247 1626 -247 0 1
rlabel polysilicon 1626 -253 1626 -253 0 3
rlabel polysilicon 1633 -247 1633 -247 0 1
rlabel polysilicon 1633 -253 1633 -253 0 3
rlabel polysilicon 1668 -247 1668 -247 0 1
rlabel polysilicon 1668 -253 1668 -253 0 3
rlabel polysilicon 1815 -247 1815 -247 0 1
rlabel polysilicon 1815 -253 1815 -253 0 3
rlabel polysilicon 1941 -247 1941 -247 0 1
rlabel polysilicon 1941 -253 1941 -253 0 3
rlabel polysilicon 16 -372 16 -372 0 1
rlabel polysilicon 16 -378 16 -378 0 3
rlabel polysilicon 23 -372 23 -372 0 1
rlabel polysilicon 23 -378 23 -378 0 3
rlabel polysilicon 30 -372 30 -372 0 1
rlabel polysilicon 30 -378 30 -378 0 3
rlabel polysilicon 37 -372 37 -372 0 1
rlabel polysilicon 37 -378 37 -378 0 3
rlabel polysilicon 47 -372 47 -372 0 2
rlabel polysilicon 44 -378 44 -378 0 3
rlabel polysilicon 51 -372 51 -372 0 1
rlabel polysilicon 54 -372 54 -372 0 2
rlabel polysilicon 54 -378 54 -378 0 4
rlabel polysilicon 58 -372 58 -372 0 1
rlabel polysilicon 58 -378 58 -378 0 3
rlabel polysilicon 65 -372 65 -372 0 1
rlabel polysilicon 65 -378 65 -378 0 3
rlabel polysilicon 72 -372 72 -372 0 1
rlabel polysilicon 72 -378 72 -378 0 3
rlabel polysilicon 79 -372 79 -372 0 1
rlabel polysilicon 79 -378 79 -378 0 3
rlabel polysilicon 86 -372 86 -372 0 1
rlabel polysilicon 86 -378 86 -378 0 3
rlabel polysilicon 93 -372 93 -372 0 1
rlabel polysilicon 93 -378 93 -378 0 3
rlabel polysilicon 96 -378 96 -378 0 4
rlabel polysilicon 100 -372 100 -372 0 1
rlabel polysilicon 100 -378 100 -378 0 3
rlabel polysilicon 107 -372 107 -372 0 1
rlabel polysilicon 107 -378 107 -378 0 3
rlabel polysilicon 114 -372 114 -372 0 1
rlabel polysilicon 114 -378 114 -378 0 3
rlabel polysilicon 121 -372 121 -372 0 1
rlabel polysilicon 121 -378 121 -378 0 3
rlabel polysilicon 128 -372 128 -372 0 1
rlabel polysilicon 128 -378 128 -378 0 3
rlabel polysilicon 135 -372 135 -372 0 1
rlabel polysilicon 138 -372 138 -372 0 2
rlabel polysilicon 142 -372 142 -372 0 1
rlabel polysilicon 142 -378 142 -378 0 3
rlabel polysilicon 149 -372 149 -372 0 1
rlabel polysilicon 149 -378 149 -378 0 3
rlabel polysilicon 156 -372 156 -372 0 1
rlabel polysilicon 156 -378 156 -378 0 3
rlabel polysilicon 163 -372 163 -372 0 1
rlabel polysilicon 166 -372 166 -372 0 2
rlabel polysilicon 163 -378 163 -378 0 3
rlabel polysilicon 166 -378 166 -378 0 4
rlabel polysilicon 170 -372 170 -372 0 1
rlabel polysilicon 170 -378 170 -378 0 3
rlabel polysilicon 177 -372 177 -372 0 1
rlabel polysilicon 177 -378 177 -378 0 3
rlabel polysilicon 187 -372 187 -372 0 2
rlabel polysilicon 184 -378 184 -378 0 3
rlabel polysilicon 187 -378 187 -378 0 4
rlabel polysilicon 191 -372 191 -372 0 1
rlabel polysilicon 191 -378 191 -378 0 3
rlabel polysilicon 198 -372 198 -372 0 1
rlabel polysilicon 198 -378 198 -378 0 3
rlabel polysilicon 205 -372 205 -372 0 1
rlabel polysilicon 205 -378 205 -378 0 3
rlabel polysilicon 212 -372 212 -372 0 1
rlabel polysilicon 212 -378 212 -378 0 3
rlabel polysilicon 219 -372 219 -372 0 1
rlabel polysilicon 219 -378 219 -378 0 3
rlabel polysilicon 226 -372 226 -372 0 1
rlabel polysilicon 226 -378 226 -378 0 3
rlabel polysilicon 233 -372 233 -372 0 1
rlabel polysilicon 233 -378 233 -378 0 3
rlabel polysilicon 240 -372 240 -372 0 1
rlabel polysilicon 243 -372 243 -372 0 2
rlabel polysilicon 240 -378 240 -378 0 3
rlabel polysilicon 247 -372 247 -372 0 1
rlabel polysilicon 247 -378 247 -378 0 3
rlabel polysilicon 254 -372 254 -372 0 1
rlabel polysilicon 254 -378 254 -378 0 3
rlabel polysilicon 261 -372 261 -372 0 1
rlabel polysilicon 261 -378 261 -378 0 3
rlabel polysilicon 268 -372 268 -372 0 1
rlabel polysilicon 268 -378 268 -378 0 3
rlabel polysilicon 275 -372 275 -372 0 1
rlabel polysilicon 275 -378 275 -378 0 3
rlabel polysilicon 282 -372 282 -372 0 1
rlabel polysilicon 282 -378 282 -378 0 3
rlabel polysilicon 289 -372 289 -372 0 1
rlabel polysilicon 289 -378 289 -378 0 3
rlabel polysilicon 296 -372 296 -372 0 1
rlabel polysilicon 296 -378 296 -378 0 3
rlabel polysilicon 303 -372 303 -372 0 1
rlabel polysilicon 303 -378 303 -378 0 3
rlabel polysilicon 310 -372 310 -372 0 1
rlabel polysilicon 310 -378 310 -378 0 3
rlabel polysilicon 317 -372 317 -372 0 1
rlabel polysilicon 317 -378 317 -378 0 3
rlabel polysilicon 324 -372 324 -372 0 1
rlabel polysilicon 324 -378 324 -378 0 3
rlabel polysilicon 331 -372 331 -372 0 1
rlabel polysilicon 331 -378 331 -378 0 3
rlabel polysilicon 338 -372 338 -372 0 1
rlabel polysilicon 338 -378 338 -378 0 3
rlabel polysilicon 345 -372 345 -372 0 1
rlabel polysilicon 345 -378 345 -378 0 3
rlabel polysilicon 352 -372 352 -372 0 1
rlabel polysilicon 352 -378 352 -378 0 3
rlabel polysilicon 359 -372 359 -372 0 1
rlabel polysilicon 359 -378 359 -378 0 3
rlabel polysilicon 366 -372 366 -372 0 1
rlabel polysilicon 366 -378 366 -378 0 3
rlabel polysilicon 373 -372 373 -372 0 1
rlabel polysilicon 373 -378 373 -378 0 3
rlabel polysilicon 380 -372 380 -372 0 1
rlabel polysilicon 380 -378 380 -378 0 3
rlabel polysilicon 387 -372 387 -372 0 1
rlabel polysilicon 387 -378 387 -378 0 3
rlabel polysilicon 394 -372 394 -372 0 1
rlabel polysilicon 394 -378 394 -378 0 3
rlabel polysilicon 401 -372 401 -372 0 1
rlabel polysilicon 404 -372 404 -372 0 2
rlabel polysilicon 401 -378 401 -378 0 3
rlabel polysilicon 408 -372 408 -372 0 1
rlabel polysilicon 408 -378 408 -378 0 3
rlabel polysilicon 415 -372 415 -372 0 1
rlabel polysilicon 415 -378 415 -378 0 3
rlabel polysilicon 422 -372 422 -372 0 1
rlabel polysilicon 422 -378 422 -378 0 3
rlabel polysilicon 432 -372 432 -372 0 2
rlabel polysilicon 429 -378 429 -378 0 3
rlabel polysilicon 432 -378 432 -378 0 4
rlabel polysilicon 436 -372 436 -372 0 1
rlabel polysilicon 436 -378 436 -378 0 3
rlabel polysilicon 443 -372 443 -372 0 1
rlabel polysilicon 443 -378 443 -378 0 3
rlabel polysilicon 446 -378 446 -378 0 4
rlabel polysilicon 450 -372 450 -372 0 1
rlabel polysilicon 450 -378 450 -378 0 3
rlabel polysilicon 457 -372 457 -372 0 1
rlabel polysilicon 457 -378 457 -378 0 3
rlabel polysilicon 464 -372 464 -372 0 1
rlabel polysilicon 464 -378 464 -378 0 3
rlabel polysilicon 471 -372 471 -372 0 1
rlabel polysilicon 471 -378 471 -378 0 3
rlabel polysilicon 478 -372 478 -372 0 1
rlabel polysilicon 481 -372 481 -372 0 2
rlabel polysilicon 478 -378 478 -378 0 3
rlabel polysilicon 481 -378 481 -378 0 4
rlabel polysilicon 485 -372 485 -372 0 1
rlabel polysilicon 485 -378 485 -378 0 3
rlabel polysilicon 492 -372 492 -372 0 1
rlabel polysilicon 492 -378 492 -378 0 3
rlabel polysilicon 499 -372 499 -372 0 1
rlabel polysilicon 499 -378 499 -378 0 3
rlabel polysilicon 506 -372 506 -372 0 1
rlabel polysilicon 506 -378 506 -378 0 3
rlabel polysilicon 513 -372 513 -372 0 1
rlabel polysilicon 513 -378 513 -378 0 3
rlabel polysilicon 520 -372 520 -372 0 1
rlabel polysilicon 520 -378 520 -378 0 3
rlabel polysilicon 527 -372 527 -372 0 1
rlabel polysilicon 527 -378 527 -378 0 3
rlabel polysilicon 534 -372 534 -372 0 1
rlabel polysilicon 534 -378 534 -378 0 3
rlabel polysilicon 541 -372 541 -372 0 1
rlabel polysilicon 541 -378 541 -378 0 3
rlabel polysilicon 548 -372 548 -372 0 1
rlabel polysilicon 548 -378 548 -378 0 3
rlabel polysilicon 555 -372 555 -372 0 1
rlabel polysilicon 555 -378 555 -378 0 3
rlabel polysilicon 562 -372 562 -372 0 1
rlabel polysilicon 562 -378 562 -378 0 3
rlabel polysilicon 569 -372 569 -372 0 1
rlabel polysilicon 569 -378 569 -378 0 3
rlabel polysilicon 576 -372 576 -372 0 1
rlabel polysilicon 576 -378 576 -378 0 3
rlabel polysilicon 583 -372 583 -372 0 1
rlabel polysilicon 583 -378 583 -378 0 3
rlabel polysilicon 590 -372 590 -372 0 1
rlabel polysilicon 590 -378 590 -378 0 3
rlabel polysilicon 597 -372 597 -372 0 1
rlabel polysilicon 597 -378 597 -378 0 3
rlabel polysilicon 604 -372 604 -372 0 1
rlabel polysilicon 604 -378 604 -378 0 3
rlabel polysilicon 611 -372 611 -372 0 1
rlabel polysilicon 611 -378 611 -378 0 3
rlabel polysilicon 618 -372 618 -372 0 1
rlabel polysilicon 618 -378 618 -378 0 3
rlabel polysilicon 625 -372 625 -372 0 1
rlabel polysilicon 628 -372 628 -372 0 2
rlabel polysilicon 625 -378 625 -378 0 3
rlabel polysilicon 632 -372 632 -372 0 1
rlabel polysilicon 632 -378 632 -378 0 3
rlabel polysilicon 635 -378 635 -378 0 4
rlabel polysilicon 639 -372 639 -372 0 1
rlabel polysilicon 639 -378 639 -378 0 3
rlabel polysilicon 646 -372 646 -372 0 1
rlabel polysilicon 649 -378 649 -378 0 4
rlabel polysilicon 653 -372 653 -372 0 1
rlabel polysilicon 653 -378 653 -378 0 3
rlabel polysilicon 660 -372 660 -372 0 1
rlabel polysilicon 660 -378 660 -378 0 3
rlabel polysilicon 667 -372 667 -372 0 1
rlabel polysilicon 667 -378 667 -378 0 3
rlabel polysilicon 674 -372 674 -372 0 1
rlabel polysilicon 674 -378 674 -378 0 3
rlabel polysilicon 681 -372 681 -372 0 1
rlabel polysilicon 681 -378 681 -378 0 3
rlabel polysilicon 688 -372 688 -372 0 1
rlabel polysilicon 688 -378 688 -378 0 3
rlabel polysilicon 695 -372 695 -372 0 1
rlabel polysilicon 695 -378 695 -378 0 3
rlabel polysilicon 702 -372 702 -372 0 1
rlabel polysilicon 702 -378 702 -378 0 3
rlabel polysilicon 709 -372 709 -372 0 1
rlabel polysilicon 709 -378 709 -378 0 3
rlabel polysilicon 716 -372 716 -372 0 1
rlabel polysilicon 716 -378 716 -378 0 3
rlabel polysilicon 723 -372 723 -372 0 1
rlabel polysilicon 723 -378 723 -378 0 3
rlabel polysilicon 730 -372 730 -372 0 1
rlabel polysilicon 730 -378 730 -378 0 3
rlabel polysilicon 737 -372 737 -372 0 1
rlabel polysilicon 737 -378 737 -378 0 3
rlabel polysilicon 747 -372 747 -372 0 2
rlabel polysilicon 744 -378 744 -378 0 3
rlabel polysilicon 747 -378 747 -378 0 4
rlabel polysilicon 751 -372 751 -372 0 1
rlabel polysilicon 751 -378 751 -378 0 3
rlabel polysilicon 761 -372 761 -372 0 2
rlabel polysilicon 758 -378 758 -378 0 3
rlabel polysilicon 761 -378 761 -378 0 4
rlabel polysilicon 765 -372 765 -372 0 1
rlabel polysilicon 765 -378 765 -378 0 3
rlabel polysilicon 772 -372 772 -372 0 1
rlabel polysilicon 772 -378 772 -378 0 3
rlabel polysilicon 775 -378 775 -378 0 4
rlabel polysilicon 779 -372 779 -372 0 1
rlabel polysilicon 779 -378 779 -378 0 3
rlabel polysilicon 786 -372 786 -372 0 1
rlabel polysilicon 786 -378 786 -378 0 3
rlabel polysilicon 793 -372 793 -372 0 1
rlabel polysilicon 796 -372 796 -372 0 2
rlabel polysilicon 793 -378 793 -378 0 3
rlabel polysilicon 796 -378 796 -378 0 4
rlabel polysilicon 800 -372 800 -372 0 1
rlabel polysilicon 803 -378 803 -378 0 4
rlabel polysilicon 810 -372 810 -372 0 2
rlabel polysilicon 807 -378 807 -378 0 3
rlabel polysilicon 810 -378 810 -378 0 4
rlabel polysilicon 814 -372 814 -372 0 1
rlabel polysilicon 814 -378 814 -378 0 3
rlabel polysilicon 821 -372 821 -372 0 1
rlabel polysilicon 821 -378 821 -378 0 3
rlabel polysilicon 828 -372 828 -372 0 1
rlabel polysilicon 828 -378 828 -378 0 3
rlabel polysilicon 835 -372 835 -372 0 1
rlabel polysilicon 838 -372 838 -372 0 2
rlabel polysilicon 835 -378 835 -378 0 3
rlabel polysilicon 842 -372 842 -372 0 1
rlabel polysilicon 845 -372 845 -372 0 2
rlabel polysilicon 842 -378 842 -378 0 3
rlabel polysilicon 845 -378 845 -378 0 4
rlabel polysilicon 849 -372 849 -372 0 1
rlabel polysilicon 849 -378 849 -378 0 3
rlabel polysilicon 856 -372 856 -372 0 1
rlabel polysilicon 856 -378 856 -378 0 3
rlabel polysilicon 863 -372 863 -372 0 1
rlabel polysilicon 863 -378 863 -378 0 3
rlabel polysilicon 870 -372 870 -372 0 1
rlabel polysilicon 870 -378 870 -378 0 3
rlabel polysilicon 877 -372 877 -372 0 1
rlabel polysilicon 880 -372 880 -372 0 2
rlabel polysilicon 877 -378 877 -378 0 3
rlabel polysilicon 884 -372 884 -372 0 1
rlabel polysilicon 884 -378 884 -378 0 3
rlabel polysilicon 891 -372 891 -372 0 1
rlabel polysilicon 894 -372 894 -372 0 2
rlabel polysilicon 891 -378 891 -378 0 3
rlabel polysilicon 898 -372 898 -372 0 1
rlabel polysilicon 898 -378 898 -378 0 3
rlabel polysilicon 905 -372 905 -372 0 1
rlabel polysilicon 905 -378 905 -378 0 3
rlabel polysilicon 912 -372 912 -372 0 1
rlabel polysilicon 912 -378 912 -378 0 3
rlabel polysilicon 919 -372 919 -372 0 1
rlabel polysilicon 919 -378 919 -378 0 3
rlabel polysilicon 926 -372 926 -372 0 1
rlabel polysilicon 926 -378 926 -378 0 3
rlabel polysilicon 933 -372 933 -372 0 1
rlabel polysilicon 933 -378 933 -378 0 3
rlabel polysilicon 940 -372 940 -372 0 1
rlabel polysilicon 940 -378 940 -378 0 3
rlabel polysilicon 947 -372 947 -372 0 1
rlabel polysilicon 947 -378 947 -378 0 3
rlabel polysilicon 954 -372 954 -372 0 1
rlabel polysilicon 954 -378 954 -378 0 3
rlabel polysilicon 961 -372 961 -372 0 1
rlabel polysilicon 961 -378 961 -378 0 3
rlabel polysilicon 968 -372 968 -372 0 1
rlabel polysilicon 968 -378 968 -378 0 3
rlabel polysilicon 975 -378 975 -378 0 3
rlabel polysilicon 978 -378 978 -378 0 4
rlabel polysilicon 982 -372 982 -372 0 1
rlabel polysilicon 982 -378 982 -378 0 3
rlabel polysilicon 989 -372 989 -372 0 1
rlabel polysilicon 989 -378 989 -378 0 3
rlabel polysilicon 992 -378 992 -378 0 4
rlabel polysilicon 996 -372 996 -372 0 1
rlabel polysilicon 996 -378 996 -378 0 3
rlabel polysilicon 1003 -372 1003 -372 0 1
rlabel polysilicon 1003 -378 1003 -378 0 3
rlabel polysilicon 1010 -372 1010 -372 0 1
rlabel polysilicon 1010 -378 1010 -378 0 3
rlabel polysilicon 1017 -372 1017 -372 0 1
rlabel polysilicon 1020 -372 1020 -372 0 2
rlabel polysilicon 1017 -378 1017 -378 0 3
rlabel polysilicon 1020 -378 1020 -378 0 4
rlabel polysilicon 1024 -372 1024 -372 0 1
rlabel polysilicon 1027 -372 1027 -372 0 2
rlabel polysilicon 1027 -378 1027 -378 0 4
rlabel polysilicon 1031 -372 1031 -372 0 1
rlabel polysilicon 1031 -378 1031 -378 0 3
rlabel polysilicon 1038 -372 1038 -372 0 1
rlabel polysilicon 1038 -378 1038 -378 0 3
rlabel polysilicon 1045 -372 1045 -372 0 1
rlabel polysilicon 1045 -378 1045 -378 0 3
rlabel polysilicon 1052 -372 1052 -372 0 1
rlabel polysilicon 1052 -378 1052 -378 0 3
rlabel polysilicon 1059 -372 1059 -372 0 1
rlabel polysilicon 1059 -378 1059 -378 0 3
rlabel polysilicon 1066 -372 1066 -372 0 1
rlabel polysilicon 1066 -378 1066 -378 0 3
rlabel polysilicon 1073 -372 1073 -372 0 1
rlabel polysilicon 1076 -372 1076 -372 0 2
rlabel polysilicon 1073 -378 1073 -378 0 3
rlabel polysilicon 1076 -378 1076 -378 0 4
rlabel polysilicon 1083 -372 1083 -372 0 2
rlabel polysilicon 1080 -378 1080 -378 0 3
rlabel polysilicon 1083 -378 1083 -378 0 4
rlabel polysilicon 1087 -372 1087 -372 0 1
rlabel polysilicon 1087 -378 1087 -378 0 3
rlabel polysilicon 1094 -372 1094 -372 0 1
rlabel polysilicon 1094 -378 1094 -378 0 3
rlabel polysilicon 1104 -372 1104 -372 0 2
rlabel polysilicon 1101 -378 1101 -378 0 3
rlabel polysilicon 1104 -378 1104 -378 0 4
rlabel polysilicon 1108 -372 1108 -372 0 1
rlabel polysilicon 1108 -378 1108 -378 0 3
rlabel polysilicon 1115 -372 1115 -372 0 1
rlabel polysilicon 1115 -378 1115 -378 0 3
rlabel polysilicon 1122 -372 1122 -372 0 1
rlabel polysilicon 1122 -378 1122 -378 0 3
rlabel polysilicon 1129 -372 1129 -372 0 1
rlabel polysilicon 1129 -378 1129 -378 0 3
rlabel polysilicon 1136 -372 1136 -372 0 1
rlabel polysilicon 1136 -378 1136 -378 0 3
rlabel polysilicon 1143 -372 1143 -372 0 1
rlabel polysilicon 1143 -378 1143 -378 0 3
rlabel polysilicon 1150 -372 1150 -372 0 1
rlabel polysilicon 1150 -378 1150 -378 0 3
rlabel polysilicon 1157 -372 1157 -372 0 1
rlabel polysilicon 1157 -378 1157 -378 0 3
rlabel polysilicon 1164 -372 1164 -372 0 1
rlabel polysilicon 1164 -378 1164 -378 0 3
rlabel polysilicon 1171 -372 1171 -372 0 1
rlabel polysilicon 1171 -378 1171 -378 0 3
rlabel polysilicon 1181 -372 1181 -372 0 2
rlabel polysilicon 1178 -378 1178 -378 0 3
rlabel polysilicon 1181 -378 1181 -378 0 4
rlabel polysilicon 1185 -372 1185 -372 0 1
rlabel polysilicon 1185 -378 1185 -378 0 3
rlabel polysilicon 1192 -372 1192 -372 0 1
rlabel polysilicon 1192 -378 1192 -378 0 3
rlabel polysilicon 1199 -372 1199 -372 0 1
rlabel polysilicon 1199 -378 1199 -378 0 3
rlabel polysilicon 1206 -372 1206 -372 0 1
rlabel polysilicon 1206 -378 1206 -378 0 3
rlabel polysilicon 1213 -372 1213 -372 0 1
rlabel polysilicon 1213 -378 1213 -378 0 3
rlabel polysilicon 1220 -372 1220 -372 0 1
rlabel polysilicon 1220 -378 1220 -378 0 3
rlabel polysilicon 1227 -372 1227 -372 0 1
rlabel polysilicon 1227 -378 1227 -378 0 3
rlabel polysilicon 1234 -372 1234 -372 0 1
rlabel polysilicon 1234 -378 1234 -378 0 3
rlabel polysilicon 1241 -372 1241 -372 0 1
rlabel polysilicon 1241 -378 1241 -378 0 3
rlabel polysilicon 1248 -372 1248 -372 0 1
rlabel polysilicon 1248 -378 1248 -378 0 3
rlabel polysilicon 1255 -372 1255 -372 0 1
rlabel polysilicon 1255 -378 1255 -378 0 3
rlabel polysilicon 1262 -372 1262 -372 0 1
rlabel polysilicon 1262 -378 1262 -378 0 3
rlabel polysilicon 1269 -372 1269 -372 0 1
rlabel polysilicon 1269 -378 1269 -378 0 3
rlabel polysilicon 1276 -372 1276 -372 0 1
rlabel polysilicon 1276 -378 1276 -378 0 3
rlabel polysilicon 1283 -372 1283 -372 0 1
rlabel polysilicon 1283 -378 1283 -378 0 3
rlabel polysilicon 1290 -372 1290 -372 0 1
rlabel polysilicon 1290 -378 1290 -378 0 3
rlabel polysilicon 1297 -372 1297 -372 0 1
rlabel polysilicon 1297 -378 1297 -378 0 3
rlabel polysilicon 1304 -372 1304 -372 0 1
rlabel polysilicon 1304 -378 1304 -378 0 3
rlabel polysilicon 1311 -372 1311 -372 0 1
rlabel polysilicon 1311 -378 1311 -378 0 3
rlabel polysilicon 1318 -372 1318 -372 0 1
rlabel polysilicon 1318 -378 1318 -378 0 3
rlabel polysilicon 1325 -372 1325 -372 0 1
rlabel polysilicon 1328 -372 1328 -372 0 2
rlabel polysilicon 1328 -378 1328 -378 0 4
rlabel polysilicon 1332 -372 1332 -372 0 1
rlabel polysilicon 1332 -378 1332 -378 0 3
rlabel polysilicon 1339 -372 1339 -372 0 1
rlabel polysilicon 1339 -378 1339 -378 0 3
rlabel polysilicon 1346 -372 1346 -372 0 1
rlabel polysilicon 1346 -378 1346 -378 0 3
rlabel polysilicon 1353 -378 1353 -378 0 3
rlabel polysilicon 1356 -378 1356 -378 0 4
rlabel polysilicon 1360 -372 1360 -372 0 1
rlabel polysilicon 1360 -378 1360 -378 0 3
rlabel polysilicon 1367 -372 1367 -372 0 1
rlabel polysilicon 1367 -378 1367 -378 0 3
rlabel polysilicon 1374 -372 1374 -372 0 1
rlabel polysilicon 1374 -378 1374 -378 0 3
rlabel polysilicon 1381 -372 1381 -372 0 1
rlabel polysilicon 1381 -378 1381 -378 0 3
rlabel polysilicon 1388 -372 1388 -372 0 1
rlabel polysilicon 1388 -378 1388 -378 0 3
rlabel polysilicon 1395 -372 1395 -372 0 1
rlabel polysilicon 1395 -378 1395 -378 0 3
rlabel polysilicon 1402 -372 1402 -372 0 1
rlabel polysilicon 1402 -378 1402 -378 0 3
rlabel polysilicon 1409 -372 1409 -372 0 1
rlabel polysilicon 1409 -378 1409 -378 0 3
rlabel polysilicon 1416 -372 1416 -372 0 1
rlabel polysilicon 1416 -378 1416 -378 0 3
rlabel polysilicon 1423 -372 1423 -372 0 1
rlabel polysilicon 1423 -378 1423 -378 0 3
rlabel polysilicon 1430 -372 1430 -372 0 1
rlabel polysilicon 1430 -378 1430 -378 0 3
rlabel polysilicon 1437 -372 1437 -372 0 1
rlabel polysilicon 1437 -378 1437 -378 0 3
rlabel polysilicon 1444 -372 1444 -372 0 1
rlabel polysilicon 1444 -378 1444 -378 0 3
rlabel polysilicon 1451 -372 1451 -372 0 1
rlabel polysilicon 1451 -378 1451 -378 0 3
rlabel polysilicon 1458 -372 1458 -372 0 1
rlabel polysilicon 1458 -378 1458 -378 0 3
rlabel polysilicon 1465 -372 1465 -372 0 1
rlabel polysilicon 1465 -378 1465 -378 0 3
rlabel polysilicon 1472 -372 1472 -372 0 1
rlabel polysilicon 1472 -378 1472 -378 0 3
rlabel polysilicon 1479 -372 1479 -372 0 1
rlabel polysilicon 1479 -378 1479 -378 0 3
rlabel polysilicon 1486 -372 1486 -372 0 1
rlabel polysilicon 1486 -378 1486 -378 0 3
rlabel polysilicon 1493 -372 1493 -372 0 1
rlabel polysilicon 1493 -378 1493 -378 0 3
rlabel polysilicon 1500 -372 1500 -372 0 1
rlabel polysilicon 1500 -378 1500 -378 0 3
rlabel polysilicon 1507 -372 1507 -372 0 1
rlabel polysilicon 1507 -378 1507 -378 0 3
rlabel polysilicon 1514 -372 1514 -372 0 1
rlabel polysilicon 1514 -378 1514 -378 0 3
rlabel polysilicon 1521 -372 1521 -372 0 1
rlabel polysilicon 1521 -378 1521 -378 0 3
rlabel polysilicon 1528 -372 1528 -372 0 1
rlabel polysilicon 1528 -378 1528 -378 0 3
rlabel polysilicon 1535 -372 1535 -372 0 1
rlabel polysilicon 1535 -378 1535 -378 0 3
rlabel polysilicon 1542 -372 1542 -372 0 1
rlabel polysilicon 1542 -378 1542 -378 0 3
rlabel polysilicon 1549 -372 1549 -372 0 1
rlabel polysilicon 1549 -378 1549 -378 0 3
rlabel polysilicon 1556 -372 1556 -372 0 1
rlabel polysilicon 1556 -378 1556 -378 0 3
rlabel polysilicon 1563 -372 1563 -372 0 1
rlabel polysilicon 1563 -378 1563 -378 0 3
rlabel polysilicon 1570 -372 1570 -372 0 1
rlabel polysilicon 1570 -378 1570 -378 0 3
rlabel polysilicon 1577 -372 1577 -372 0 1
rlabel polysilicon 1577 -378 1577 -378 0 3
rlabel polysilicon 1584 -372 1584 -372 0 1
rlabel polysilicon 1584 -378 1584 -378 0 3
rlabel polysilicon 1591 -372 1591 -372 0 1
rlabel polysilicon 1591 -378 1591 -378 0 3
rlabel polysilicon 1598 -372 1598 -372 0 1
rlabel polysilicon 1598 -378 1598 -378 0 3
rlabel polysilicon 1605 -372 1605 -372 0 1
rlabel polysilicon 1605 -378 1605 -378 0 3
rlabel polysilicon 1612 -372 1612 -372 0 1
rlabel polysilicon 1615 -372 1615 -372 0 2
rlabel polysilicon 1612 -378 1612 -378 0 3
rlabel polysilicon 1619 -372 1619 -372 0 1
rlabel polysilicon 1619 -378 1619 -378 0 3
rlabel polysilicon 1626 -372 1626 -372 0 1
rlabel polysilicon 1626 -378 1626 -378 0 3
rlabel polysilicon 1633 -372 1633 -372 0 1
rlabel polysilicon 1633 -378 1633 -378 0 3
rlabel polysilicon 1640 -372 1640 -372 0 1
rlabel polysilicon 1640 -378 1640 -378 0 3
rlabel polysilicon 1647 -372 1647 -372 0 1
rlabel polysilicon 1647 -378 1647 -378 0 3
rlabel polysilicon 1654 -372 1654 -372 0 1
rlabel polysilicon 1654 -378 1654 -378 0 3
rlabel polysilicon 1661 -372 1661 -372 0 1
rlabel polysilicon 1661 -378 1661 -378 0 3
rlabel polysilicon 1668 -372 1668 -372 0 1
rlabel polysilicon 1668 -378 1668 -378 0 3
rlabel polysilicon 1675 -372 1675 -372 0 1
rlabel polysilicon 1675 -378 1675 -378 0 3
rlabel polysilicon 1682 -372 1682 -372 0 1
rlabel polysilicon 1682 -378 1682 -378 0 3
rlabel polysilicon 1689 -372 1689 -372 0 1
rlabel polysilicon 1689 -378 1689 -378 0 3
rlabel polysilicon 1696 -372 1696 -372 0 1
rlabel polysilicon 1696 -378 1696 -378 0 3
rlabel polysilicon 1703 -372 1703 -372 0 1
rlabel polysilicon 1703 -378 1703 -378 0 3
rlabel polysilicon 1710 -372 1710 -372 0 1
rlabel polysilicon 1710 -378 1710 -378 0 3
rlabel polysilicon 1717 -372 1717 -372 0 1
rlabel polysilicon 1717 -378 1717 -378 0 3
rlabel polysilicon 1724 -372 1724 -372 0 1
rlabel polysilicon 1724 -378 1724 -378 0 3
rlabel polysilicon 1731 -372 1731 -372 0 1
rlabel polysilicon 1731 -378 1731 -378 0 3
rlabel polysilicon 1738 -372 1738 -372 0 1
rlabel polysilicon 1738 -378 1738 -378 0 3
rlabel polysilicon 1745 -372 1745 -372 0 1
rlabel polysilicon 1745 -378 1745 -378 0 3
rlabel polysilicon 1752 -372 1752 -372 0 1
rlabel polysilicon 1752 -378 1752 -378 0 3
rlabel polysilicon 1759 -372 1759 -372 0 1
rlabel polysilicon 1759 -378 1759 -378 0 3
rlabel polysilicon 1766 -372 1766 -372 0 1
rlabel polysilicon 1766 -378 1766 -378 0 3
rlabel polysilicon 1773 -372 1773 -372 0 1
rlabel polysilicon 1773 -378 1773 -378 0 3
rlabel polysilicon 1780 -372 1780 -372 0 1
rlabel polysilicon 1780 -378 1780 -378 0 3
rlabel polysilicon 1787 -372 1787 -372 0 1
rlabel polysilicon 1787 -378 1787 -378 0 3
rlabel polysilicon 1794 -372 1794 -372 0 1
rlabel polysilicon 1794 -378 1794 -378 0 3
rlabel polysilicon 1801 -372 1801 -372 0 1
rlabel polysilicon 1801 -378 1801 -378 0 3
rlabel polysilicon 1808 -372 1808 -372 0 1
rlabel polysilicon 1808 -378 1808 -378 0 3
rlabel polysilicon 1815 -372 1815 -372 0 1
rlabel polysilicon 1815 -378 1815 -378 0 3
rlabel polysilicon 1822 -372 1822 -372 0 1
rlabel polysilicon 1822 -378 1822 -378 0 3
rlabel polysilicon 1829 -372 1829 -372 0 1
rlabel polysilicon 1829 -378 1829 -378 0 3
rlabel polysilicon 1836 -372 1836 -372 0 1
rlabel polysilicon 1836 -378 1836 -378 0 3
rlabel polysilicon 1843 -372 1843 -372 0 1
rlabel polysilicon 1843 -378 1843 -378 0 3
rlabel polysilicon 1927 -372 1927 -372 0 1
rlabel polysilicon 1927 -378 1927 -378 0 3
rlabel polysilicon 1962 -372 1962 -372 0 1
rlabel polysilicon 1962 -378 1962 -378 0 3
rlabel polysilicon 1969 -372 1969 -372 0 1
rlabel polysilicon 1969 -378 1969 -378 0 3
rlabel polysilicon 1983 -372 1983 -372 0 1
rlabel polysilicon 1983 -378 1983 -378 0 3
rlabel polysilicon 2004 -372 2004 -372 0 1
rlabel polysilicon 2004 -378 2004 -378 0 3
rlabel polysilicon 2193 -372 2193 -372 0 1
rlabel polysilicon 2193 -378 2193 -378 0 3
rlabel polysilicon 2 -501 2 -501 0 1
rlabel polysilicon 2 -507 2 -507 0 3
rlabel polysilicon 9 -507 9 -507 0 3
rlabel polysilicon 16 -501 16 -501 0 1
rlabel polysilicon 16 -507 16 -507 0 3
rlabel polysilicon 23 -501 23 -501 0 1
rlabel polysilicon 23 -507 23 -507 0 3
rlabel polysilicon 44 -501 44 -501 0 1
rlabel polysilicon 44 -507 44 -507 0 3
rlabel polysilicon 51 -501 51 -501 0 1
rlabel polysilicon 51 -507 51 -507 0 3
rlabel polysilicon 61 -501 61 -501 0 2
rlabel polysilicon 61 -507 61 -507 0 4
rlabel polysilicon 65 -501 65 -501 0 1
rlabel polysilicon 65 -507 65 -507 0 3
rlabel polysilicon 72 -501 72 -501 0 1
rlabel polysilicon 72 -507 72 -507 0 3
rlabel polysilicon 79 -501 79 -501 0 1
rlabel polysilicon 79 -507 79 -507 0 3
rlabel polysilicon 86 -501 86 -501 0 1
rlabel polysilicon 86 -507 86 -507 0 3
rlabel polysilicon 93 -501 93 -501 0 1
rlabel polysilicon 93 -507 93 -507 0 3
rlabel polysilicon 100 -501 100 -501 0 1
rlabel polysilicon 100 -507 100 -507 0 3
rlabel polysilicon 107 -501 107 -501 0 1
rlabel polysilicon 107 -507 107 -507 0 3
rlabel polysilicon 114 -507 114 -507 0 3
rlabel polysilicon 117 -507 117 -507 0 4
rlabel polysilicon 121 -501 121 -501 0 1
rlabel polysilicon 121 -507 121 -507 0 3
rlabel polysilicon 128 -501 128 -501 0 1
rlabel polysilicon 128 -507 128 -507 0 3
rlabel polysilicon 135 -501 135 -501 0 1
rlabel polysilicon 135 -507 135 -507 0 3
rlabel polysilicon 142 -501 142 -501 0 1
rlabel polysilicon 142 -507 142 -507 0 3
rlabel polysilicon 149 -501 149 -501 0 1
rlabel polysilicon 149 -507 149 -507 0 3
rlabel polysilicon 156 -501 156 -501 0 1
rlabel polysilicon 156 -507 156 -507 0 3
rlabel polysilicon 163 -501 163 -501 0 1
rlabel polysilicon 166 -501 166 -501 0 2
rlabel polysilicon 166 -507 166 -507 0 4
rlabel polysilicon 173 -501 173 -501 0 2
rlabel polysilicon 170 -507 170 -507 0 3
rlabel polysilicon 173 -507 173 -507 0 4
rlabel polysilicon 177 -501 177 -501 0 1
rlabel polysilicon 177 -507 177 -507 0 3
rlabel polysilicon 184 -501 184 -501 0 1
rlabel polysilicon 184 -507 184 -507 0 3
rlabel polysilicon 191 -501 191 -501 0 1
rlabel polysilicon 191 -507 191 -507 0 3
rlabel polysilicon 198 -501 198 -501 0 1
rlabel polysilicon 198 -507 198 -507 0 3
rlabel polysilicon 205 -501 205 -501 0 1
rlabel polysilicon 205 -507 205 -507 0 3
rlabel polysilicon 212 -501 212 -501 0 1
rlabel polysilicon 215 -501 215 -501 0 2
rlabel polysilicon 215 -507 215 -507 0 4
rlabel polysilicon 219 -501 219 -501 0 1
rlabel polysilicon 222 -501 222 -501 0 2
rlabel polysilicon 219 -507 219 -507 0 3
rlabel polysilicon 222 -507 222 -507 0 4
rlabel polysilicon 226 -501 226 -501 0 1
rlabel polysilicon 226 -507 226 -507 0 3
rlabel polysilicon 233 -501 233 -501 0 1
rlabel polysilicon 233 -507 233 -507 0 3
rlabel polysilicon 236 -507 236 -507 0 4
rlabel polysilicon 240 -501 240 -501 0 1
rlabel polysilicon 240 -507 240 -507 0 3
rlabel polysilicon 247 -501 247 -501 0 1
rlabel polysilicon 247 -507 247 -507 0 3
rlabel polysilicon 254 -501 254 -501 0 1
rlabel polysilicon 254 -507 254 -507 0 3
rlabel polysilicon 261 -501 261 -501 0 1
rlabel polysilicon 261 -507 261 -507 0 3
rlabel polysilicon 268 -501 268 -501 0 1
rlabel polysilicon 268 -507 268 -507 0 3
rlabel polysilicon 275 -501 275 -501 0 1
rlabel polysilicon 275 -507 275 -507 0 3
rlabel polysilicon 282 -501 282 -501 0 1
rlabel polysilicon 282 -507 282 -507 0 3
rlabel polysilicon 289 -501 289 -501 0 1
rlabel polysilicon 289 -507 289 -507 0 3
rlabel polysilicon 296 -501 296 -501 0 1
rlabel polysilicon 296 -507 296 -507 0 3
rlabel polysilicon 303 -501 303 -501 0 1
rlabel polysilicon 303 -507 303 -507 0 3
rlabel polysilicon 310 -501 310 -501 0 1
rlabel polysilicon 310 -507 310 -507 0 3
rlabel polysilicon 317 -501 317 -501 0 1
rlabel polysilicon 317 -507 317 -507 0 3
rlabel polysilicon 324 -501 324 -501 0 1
rlabel polysilicon 324 -507 324 -507 0 3
rlabel polysilicon 331 -501 331 -501 0 1
rlabel polysilicon 331 -507 331 -507 0 3
rlabel polysilicon 338 -501 338 -501 0 1
rlabel polysilicon 338 -507 338 -507 0 3
rlabel polysilicon 345 -501 345 -501 0 1
rlabel polysilicon 345 -507 345 -507 0 3
rlabel polysilicon 352 -501 352 -501 0 1
rlabel polysilicon 352 -507 352 -507 0 3
rlabel polysilicon 359 -501 359 -501 0 1
rlabel polysilicon 359 -507 359 -507 0 3
rlabel polysilicon 366 -501 366 -501 0 1
rlabel polysilicon 366 -507 366 -507 0 3
rlabel polysilicon 373 -501 373 -501 0 1
rlabel polysilicon 373 -507 373 -507 0 3
rlabel polysilicon 380 -501 380 -501 0 1
rlabel polysilicon 380 -507 380 -507 0 3
rlabel polysilicon 387 -501 387 -501 0 1
rlabel polysilicon 387 -507 387 -507 0 3
rlabel polysilicon 394 -501 394 -501 0 1
rlabel polysilicon 394 -507 394 -507 0 3
rlabel polysilicon 401 -501 401 -501 0 1
rlabel polysilicon 401 -507 401 -507 0 3
rlabel polysilicon 408 -501 408 -501 0 1
rlabel polysilicon 408 -507 408 -507 0 3
rlabel polysilicon 415 -501 415 -501 0 1
rlabel polysilicon 415 -507 415 -507 0 3
rlabel polysilicon 422 -501 422 -501 0 1
rlabel polysilicon 422 -507 422 -507 0 3
rlabel polysilicon 429 -501 429 -501 0 1
rlabel polysilicon 429 -507 429 -507 0 3
rlabel polysilicon 436 -501 436 -501 0 1
rlabel polysilicon 436 -507 436 -507 0 3
rlabel polysilicon 443 -501 443 -501 0 1
rlabel polysilicon 443 -507 443 -507 0 3
rlabel polysilicon 450 -501 450 -501 0 1
rlabel polysilicon 450 -507 450 -507 0 3
rlabel polysilicon 457 -501 457 -501 0 1
rlabel polysilicon 457 -507 457 -507 0 3
rlabel polysilicon 464 -501 464 -501 0 1
rlabel polysilicon 464 -507 464 -507 0 3
rlabel polysilicon 471 -501 471 -501 0 1
rlabel polysilicon 471 -507 471 -507 0 3
rlabel polysilicon 478 -501 478 -501 0 1
rlabel polysilicon 478 -507 478 -507 0 3
rlabel polysilicon 485 -501 485 -501 0 1
rlabel polysilicon 485 -507 485 -507 0 3
rlabel polysilicon 492 -501 492 -501 0 1
rlabel polysilicon 495 -501 495 -501 0 2
rlabel polysilicon 492 -507 492 -507 0 3
rlabel polysilicon 495 -507 495 -507 0 4
rlabel polysilicon 499 -501 499 -501 0 1
rlabel polysilicon 499 -507 499 -507 0 3
rlabel polysilicon 506 -501 506 -501 0 1
rlabel polysilicon 506 -507 506 -507 0 3
rlabel polysilicon 513 -501 513 -501 0 1
rlabel polysilicon 513 -507 513 -507 0 3
rlabel polysilicon 520 -501 520 -501 0 1
rlabel polysilicon 520 -507 520 -507 0 3
rlabel polysilicon 527 -501 527 -501 0 1
rlabel polysilicon 527 -507 527 -507 0 3
rlabel polysilicon 534 -501 534 -501 0 1
rlabel polysilicon 534 -507 534 -507 0 3
rlabel polysilicon 537 -507 537 -507 0 4
rlabel polysilicon 541 -501 541 -501 0 1
rlabel polysilicon 541 -507 541 -507 0 3
rlabel polysilicon 548 -501 548 -501 0 1
rlabel polysilicon 548 -507 548 -507 0 3
rlabel polysilicon 555 -501 555 -501 0 1
rlabel polysilicon 555 -507 555 -507 0 3
rlabel polysilicon 562 -501 562 -501 0 1
rlabel polysilicon 562 -507 562 -507 0 3
rlabel polysilicon 569 -501 569 -501 0 1
rlabel polysilicon 569 -507 569 -507 0 3
rlabel polysilicon 576 -501 576 -501 0 1
rlabel polysilicon 576 -507 576 -507 0 3
rlabel polysilicon 583 -501 583 -501 0 1
rlabel polysilicon 583 -507 583 -507 0 3
rlabel polysilicon 590 -501 590 -501 0 1
rlabel polysilicon 590 -507 590 -507 0 3
rlabel polysilicon 597 -501 597 -501 0 1
rlabel polysilicon 600 -501 600 -501 0 2
rlabel polysilicon 600 -507 600 -507 0 4
rlabel polysilicon 604 -501 604 -501 0 1
rlabel polysilicon 604 -507 604 -507 0 3
rlabel polysilicon 611 -501 611 -501 0 1
rlabel polysilicon 611 -507 611 -507 0 3
rlabel polysilicon 618 -501 618 -501 0 1
rlabel polysilicon 621 -501 621 -501 0 2
rlabel polysilicon 618 -507 618 -507 0 3
rlabel polysilicon 621 -507 621 -507 0 4
rlabel polysilicon 625 -501 625 -501 0 1
rlabel polysilicon 625 -507 625 -507 0 3
rlabel polysilicon 632 -501 632 -501 0 1
rlabel polysilicon 635 -507 635 -507 0 4
rlabel polysilicon 639 -501 639 -501 0 1
rlabel polysilicon 639 -507 639 -507 0 3
rlabel polysilicon 646 -501 646 -501 0 1
rlabel polysilicon 646 -507 646 -507 0 3
rlabel polysilicon 653 -501 653 -501 0 1
rlabel polysilicon 653 -507 653 -507 0 3
rlabel polysilicon 656 -507 656 -507 0 4
rlabel polysilicon 660 -501 660 -501 0 1
rlabel polysilicon 660 -507 660 -507 0 3
rlabel polysilicon 667 -501 667 -501 0 1
rlabel polysilicon 667 -507 667 -507 0 3
rlabel polysilicon 674 -501 674 -501 0 1
rlabel polysilicon 674 -507 674 -507 0 3
rlabel polysilicon 681 -501 681 -501 0 1
rlabel polysilicon 681 -507 681 -507 0 3
rlabel polysilicon 688 -501 688 -501 0 1
rlabel polysilicon 688 -507 688 -507 0 3
rlabel polysilicon 695 -501 695 -501 0 1
rlabel polysilicon 695 -507 695 -507 0 3
rlabel polysilicon 702 -501 702 -501 0 1
rlabel polysilicon 702 -507 702 -507 0 3
rlabel polysilicon 709 -501 709 -501 0 1
rlabel polysilicon 709 -507 709 -507 0 3
rlabel polysilicon 716 -501 716 -501 0 1
rlabel polysilicon 719 -501 719 -501 0 2
rlabel polysilicon 716 -507 716 -507 0 3
rlabel polysilicon 723 -501 723 -501 0 1
rlabel polysilicon 726 -501 726 -501 0 2
rlabel polysilicon 723 -507 723 -507 0 3
rlabel polysilicon 726 -507 726 -507 0 4
rlabel polysilicon 730 -501 730 -501 0 1
rlabel polysilicon 730 -507 730 -507 0 3
rlabel polysilicon 737 -501 737 -501 0 1
rlabel polysilicon 740 -501 740 -501 0 2
rlabel polysilicon 737 -507 737 -507 0 3
rlabel polysilicon 740 -507 740 -507 0 4
rlabel polysilicon 744 -501 744 -501 0 1
rlabel polysilicon 744 -507 744 -507 0 3
rlabel polysilicon 751 -501 751 -501 0 1
rlabel polysilicon 751 -507 751 -507 0 3
rlabel polysilicon 758 -501 758 -501 0 1
rlabel polysilicon 758 -507 758 -507 0 3
rlabel polysilicon 765 -501 765 -501 0 1
rlabel polysilicon 765 -507 765 -507 0 3
rlabel polysilicon 772 -501 772 -501 0 1
rlabel polysilicon 772 -507 772 -507 0 3
rlabel polysilicon 779 -501 779 -501 0 1
rlabel polysilicon 779 -507 779 -507 0 3
rlabel polysilicon 786 -501 786 -501 0 1
rlabel polysilicon 786 -507 786 -507 0 3
rlabel polysilicon 793 -501 793 -501 0 1
rlabel polysilicon 793 -507 793 -507 0 3
rlabel polysilicon 800 -501 800 -501 0 1
rlabel polysilicon 800 -507 800 -507 0 3
rlabel polysilicon 807 -501 807 -501 0 1
rlabel polysilicon 807 -507 807 -507 0 3
rlabel polysilicon 814 -501 814 -501 0 1
rlabel polysilicon 814 -507 814 -507 0 3
rlabel polysilicon 821 -501 821 -501 0 1
rlabel polysilicon 821 -507 821 -507 0 3
rlabel polysilicon 828 -501 828 -501 0 1
rlabel polysilicon 828 -507 828 -507 0 3
rlabel polysilicon 835 -501 835 -501 0 1
rlabel polysilicon 835 -507 835 -507 0 3
rlabel polysilicon 842 -501 842 -501 0 1
rlabel polysilicon 842 -507 842 -507 0 3
rlabel polysilicon 849 -501 849 -501 0 1
rlabel polysilicon 852 -501 852 -501 0 2
rlabel polysilicon 849 -507 849 -507 0 3
rlabel polysilicon 856 -501 856 -501 0 1
rlabel polysilicon 856 -507 856 -507 0 3
rlabel polysilicon 863 -501 863 -501 0 1
rlabel polysilicon 863 -507 863 -507 0 3
rlabel polysilicon 870 -501 870 -501 0 1
rlabel polysilicon 870 -507 870 -507 0 3
rlabel polysilicon 877 -501 877 -501 0 1
rlabel polysilicon 877 -507 877 -507 0 3
rlabel polysilicon 887 -501 887 -501 0 2
rlabel polysilicon 887 -507 887 -507 0 4
rlabel polysilicon 891 -501 891 -501 0 1
rlabel polysilicon 891 -507 891 -507 0 3
rlabel polysilicon 898 -501 898 -501 0 1
rlabel polysilicon 898 -507 898 -507 0 3
rlabel polysilicon 905 -501 905 -501 0 1
rlabel polysilicon 905 -507 905 -507 0 3
rlabel polysilicon 912 -501 912 -501 0 1
rlabel polysilicon 912 -507 912 -507 0 3
rlabel polysilicon 915 -507 915 -507 0 4
rlabel polysilicon 919 -501 919 -501 0 1
rlabel polysilicon 919 -507 919 -507 0 3
rlabel polysilicon 926 -501 926 -501 0 1
rlabel polysilicon 926 -507 926 -507 0 3
rlabel polysilicon 933 -501 933 -501 0 1
rlabel polysilicon 933 -507 933 -507 0 3
rlabel polysilicon 936 -507 936 -507 0 4
rlabel polysilicon 940 -501 940 -501 0 1
rlabel polysilicon 940 -507 940 -507 0 3
rlabel polysilicon 947 -501 947 -501 0 1
rlabel polysilicon 947 -507 947 -507 0 3
rlabel polysilicon 954 -501 954 -501 0 1
rlabel polysilicon 957 -501 957 -501 0 2
rlabel polysilicon 954 -507 954 -507 0 3
rlabel polysilicon 961 -501 961 -501 0 1
rlabel polysilicon 961 -507 961 -507 0 3
rlabel polysilicon 968 -501 968 -501 0 1
rlabel polysilicon 971 -501 971 -501 0 2
rlabel polysilicon 968 -507 968 -507 0 3
rlabel polysilicon 971 -507 971 -507 0 4
rlabel polysilicon 978 -501 978 -501 0 2
rlabel polysilicon 975 -507 975 -507 0 3
rlabel polysilicon 978 -507 978 -507 0 4
rlabel polysilicon 982 -501 982 -501 0 1
rlabel polysilicon 985 -501 985 -501 0 2
rlabel polysilicon 982 -507 982 -507 0 3
rlabel polysilicon 985 -507 985 -507 0 4
rlabel polysilicon 989 -501 989 -501 0 1
rlabel polysilicon 989 -507 989 -507 0 3
rlabel polysilicon 992 -507 992 -507 0 4
rlabel polysilicon 996 -501 996 -501 0 1
rlabel polysilicon 996 -507 996 -507 0 3
rlabel polysilicon 1006 -501 1006 -501 0 2
rlabel polysilicon 1003 -507 1003 -507 0 3
rlabel polysilicon 1006 -507 1006 -507 0 4
rlabel polysilicon 1010 -501 1010 -501 0 1
rlabel polysilicon 1010 -507 1010 -507 0 3
rlabel polysilicon 1017 -501 1017 -501 0 1
rlabel polysilicon 1017 -507 1017 -507 0 3
rlabel polysilicon 1024 -501 1024 -501 0 1
rlabel polysilicon 1027 -501 1027 -501 0 2
rlabel polysilicon 1031 -501 1031 -501 0 1
rlabel polysilicon 1031 -507 1031 -507 0 3
rlabel polysilicon 1038 -501 1038 -501 0 1
rlabel polysilicon 1038 -507 1038 -507 0 3
rlabel polysilicon 1045 -501 1045 -501 0 1
rlabel polysilicon 1045 -507 1045 -507 0 3
rlabel polysilicon 1052 -501 1052 -501 0 1
rlabel polysilicon 1052 -507 1052 -507 0 3
rlabel polysilicon 1059 -501 1059 -501 0 1
rlabel polysilicon 1059 -507 1059 -507 0 3
rlabel polysilicon 1066 -501 1066 -501 0 1
rlabel polysilicon 1066 -507 1066 -507 0 3
rlabel polysilicon 1073 -501 1073 -501 0 1
rlabel polysilicon 1073 -507 1073 -507 0 3
rlabel polysilicon 1080 -501 1080 -501 0 1
rlabel polysilicon 1083 -501 1083 -501 0 2
rlabel polysilicon 1080 -507 1080 -507 0 3
rlabel polysilicon 1083 -507 1083 -507 0 4
rlabel polysilicon 1087 -501 1087 -501 0 1
rlabel polysilicon 1087 -507 1087 -507 0 3
rlabel polysilicon 1094 -501 1094 -501 0 1
rlabel polysilicon 1094 -507 1094 -507 0 3
rlabel polysilicon 1101 -501 1101 -501 0 1
rlabel polysilicon 1101 -507 1101 -507 0 3
rlabel polysilicon 1108 -501 1108 -501 0 1
rlabel polysilicon 1108 -507 1108 -507 0 3
rlabel polysilicon 1115 -501 1115 -501 0 1
rlabel polysilicon 1115 -507 1115 -507 0 3
rlabel polysilicon 1122 -501 1122 -501 0 1
rlabel polysilicon 1125 -501 1125 -501 0 2
rlabel polysilicon 1125 -507 1125 -507 0 4
rlabel polysilicon 1129 -501 1129 -501 0 1
rlabel polysilicon 1129 -507 1129 -507 0 3
rlabel polysilicon 1136 -501 1136 -501 0 1
rlabel polysilicon 1136 -507 1136 -507 0 3
rlabel polysilicon 1143 -501 1143 -501 0 1
rlabel polysilicon 1143 -507 1143 -507 0 3
rlabel polysilicon 1150 -501 1150 -501 0 1
rlabel polysilicon 1150 -507 1150 -507 0 3
rlabel polysilicon 1157 -501 1157 -501 0 1
rlabel polysilicon 1157 -507 1157 -507 0 3
rlabel polysilicon 1167 -501 1167 -501 0 2
rlabel polysilicon 1164 -507 1164 -507 0 3
rlabel polysilicon 1167 -507 1167 -507 0 4
rlabel polysilicon 1171 -501 1171 -501 0 1
rlabel polysilicon 1171 -507 1171 -507 0 3
rlabel polysilicon 1178 -501 1178 -501 0 1
rlabel polysilicon 1178 -507 1178 -507 0 3
rlabel polysilicon 1185 -501 1185 -501 0 1
rlabel polysilicon 1185 -507 1185 -507 0 3
rlabel polysilicon 1192 -501 1192 -501 0 1
rlabel polysilicon 1192 -507 1192 -507 0 3
rlabel polysilicon 1199 -501 1199 -501 0 1
rlabel polysilicon 1199 -507 1199 -507 0 3
rlabel polysilicon 1206 -501 1206 -501 0 1
rlabel polysilicon 1206 -507 1206 -507 0 3
rlabel polysilicon 1213 -501 1213 -501 0 1
rlabel polysilicon 1213 -507 1213 -507 0 3
rlabel polysilicon 1220 -501 1220 -501 0 1
rlabel polysilicon 1220 -507 1220 -507 0 3
rlabel polysilicon 1227 -501 1227 -501 0 1
rlabel polysilicon 1227 -507 1227 -507 0 3
rlabel polysilicon 1234 -501 1234 -501 0 1
rlabel polysilicon 1234 -507 1234 -507 0 3
rlabel polysilicon 1241 -501 1241 -501 0 1
rlabel polysilicon 1241 -507 1241 -507 0 3
rlabel polysilicon 1248 -501 1248 -501 0 1
rlabel polysilicon 1248 -507 1248 -507 0 3
rlabel polysilicon 1255 -501 1255 -501 0 1
rlabel polysilicon 1255 -507 1255 -507 0 3
rlabel polysilicon 1262 -501 1262 -501 0 1
rlabel polysilicon 1262 -507 1262 -507 0 3
rlabel polysilicon 1269 -501 1269 -501 0 1
rlabel polysilicon 1269 -507 1269 -507 0 3
rlabel polysilicon 1276 -501 1276 -501 0 1
rlabel polysilicon 1276 -507 1276 -507 0 3
rlabel polysilicon 1283 -501 1283 -501 0 1
rlabel polysilicon 1283 -507 1283 -507 0 3
rlabel polysilicon 1290 -501 1290 -501 0 1
rlabel polysilicon 1290 -507 1290 -507 0 3
rlabel polysilicon 1297 -501 1297 -501 0 1
rlabel polysilicon 1297 -507 1297 -507 0 3
rlabel polysilicon 1304 -501 1304 -501 0 1
rlabel polysilicon 1304 -507 1304 -507 0 3
rlabel polysilicon 1311 -501 1311 -501 0 1
rlabel polysilicon 1311 -507 1311 -507 0 3
rlabel polysilicon 1318 -501 1318 -501 0 1
rlabel polysilicon 1318 -507 1318 -507 0 3
rlabel polysilicon 1325 -501 1325 -501 0 1
rlabel polysilicon 1325 -507 1325 -507 0 3
rlabel polysilicon 1332 -501 1332 -501 0 1
rlabel polysilicon 1332 -507 1332 -507 0 3
rlabel polysilicon 1339 -501 1339 -501 0 1
rlabel polysilicon 1339 -507 1339 -507 0 3
rlabel polysilicon 1346 -501 1346 -501 0 1
rlabel polysilicon 1346 -507 1346 -507 0 3
rlabel polysilicon 1353 -501 1353 -501 0 1
rlabel polysilicon 1353 -507 1353 -507 0 3
rlabel polysilicon 1360 -501 1360 -501 0 1
rlabel polysilicon 1360 -507 1360 -507 0 3
rlabel polysilicon 1367 -501 1367 -501 0 1
rlabel polysilicon 1367 -507 1367 -507 0 3
rlabel polysilicon 1374 -501 1374 -501 0 1
rlabel polysilicon 1374 -507 1374 -507 0 3
rlabel polysilicon 1381 -501 1381 -501 0 1
rlabel polysilicon 1381 -507 1381 -507 0 3
rlabel polysilicon 1388 -501 1388 -501 0 1
rlabel polysilicon 1388 -507 1388 -507 0 3
rlabel polysilicon 1395 -501 1395 -501 0 1
rlabel polysilicon 1395 -507 1395 -507 0 3
rlabel polysilicon 1402 -501 1402 -501 0 1
rlabel polysilicon 1402 -507 1402 -507 0 3
rlabel polysilicon 1409 -501 1409 -501 0 1
rlabel polysilicon 1409 -507 1409 -507 0 3
rlabel polysilicon 1416 -501 1416 -501 0 1
rlabel polysilicon 1416 -507 1416 -507 0 3
rlabel polysilicon 1423 -501 1423 -501 0 1
rlabel polysilicon 1423 -507 1423 -507 0 3
rlabel polysilicon 1430 -501 1430 -501 0 1
rlabel polysilicon 1430 -507 1430 -507 0 3
rlabel polysilicon 1440 -501 1440 -501 0 2
rlabel polysilicon 1437 -507 1437 -507 0 3
rlabel polysilicon 1440 -507 1440 -507 0 4
rlabel polysilicon 1444 -501 1444 -501 0 1
rlabel polysilicon 1444 -507 1444 -507 0 3
rlabel polysilicon 1451 -501 1451 -501 0 1
rlabel polysilicon 1451 -507 1451 -507 0 3
rlabel polysilicon 1458 -501 1458 -501 0 1
rlabel polysilicon 1458 -507 1458 -507 0 3
rlabel polysilicon 1465 -501 1465 -501 0 1
rlabel polysilicon 1465 -507 1465 -507 0 3
rlabel polysilicon 1472 -501 1472 -501 0 1
rlabel polysilicon 1472 -507 1472 -507 0 3
rlabel polysilicon 1479 -501 1479 -501 0 1
rlabel polysilicon 1479 -507 1479 -507 0 3
rlabel polysilicon 1486 -501 1486 -501 0 1
rlabel polysilicon 1486 -507 1486 -507 0 3
rlabel polysilicon 1493 -501 1493 -501 0 1
rlabel polysilicon 1493 -507 1493 -507 0 3
rlabel polysilicon 1500 -501 1500 -501 0 1
rlabel polysilicon 1500 -507 1500 -507 0 3
rlabel polysilicon 1507 -501 1507 -501 0 1
rlabel polysilicon 1507 -507 1507 -507 0 3
rlabel polysilicon 1514 -501 1514 -501 0 1
rlabel polysilicon 1514 -507 1514 -507 0 3
rlabel polysilicon 1521 -501 1521 -501 0 1
rlabel polysilicon 1521 -507 1521 -507 0 3
rlabel polysilicon 1528 -501 1528 -501 0 1
rlabel polysilicon 1528 -507 1528 -507 0 3
rlabel polysilicon 1535 -501 1535 -501 0 1
rlabel polysilicon 1535 -507 1535 -507 0 3
rlabel polysilicon 1542 -501 1542 -501 0 1
rlabel polysilicon 1542 -507 1542 -507 0 3
rlabel polysilicon 1549 -501 1549 -501 0 1
rlabel polysilicon 1549 -507 1549 -507 0 3
rlabel polysilicon 1556 -501 1556 -501 0 1
rlabel polysilicon 1556 -507 1556 -507 0 3
rlabel polysilicon 1563 -501 1563 -501 0 1
rlabel polysilicon 1563 -507 1563 -507 0 3
rlabel polysilicon 1570 -501 1570 -501 0 1
rlabel polysilicon 1570 -507 1570 -507 0 3
rlabel polysilicon 1577 -501 1577 -501 0 1
rlabel polysilicon 1577 -507 1577 -507 0 3
rlabel polysilicon 1584 -501 1584 -501 0 1
rlabel polysilicon 1584 -507 1584 -507 0 3
rlabel polysilicon 1591 -501 1591 -501 0 1
rlabel polysilicon 1591 -507 1591 -507 0 3
rlabel polysilicon 1598 -501 1598 -501 0 1
rlabel polysilicon 1598 -507 1598 -507 0 3
rlabel polysilicon 1605 -501 1605 -501 0 1
rlabel polysilicon 1605 -507 1605 -507 0 3
rlabel polysilicon 1612 -501 1612 -501 0 1
rlabel polysilicon 1612 -507 1612 -507 0 3
rlabel polysilicon 1619 -501 1619 -501 0 1
rlabel polysilicon 1619 -507 1619 -507 0 3
rlabel polysilicon 1626 -501 1626 -501 0 1
rlabel polysilicon 1626 -507 1626 -507 0 3
rlabel polysilicon 1633 -501 1633 -501 0 1
rlabel polysilicon 1633 -507 1633 -507 0 3
rlabel polysilicon 1640 -501 1640 -501 0 1
rlabel polysilicon 1640 -507 1640 -507 0 3
rlabel polysilicon 1647 -501 1647 -501 0 1
rlabel polysilicon 1647 -507 1647 -507 0 3
rlabel polysilicon 1654 -501 1654 -501 0 1
rlabel polysilicon 1654 -507 1654 -507 0 3
rlabel polysilicon 1661 -501 1661 -501 0 1
rlabel polysilicon 1661 -507 1661 -507 0 3
rlabel polysilicon 1668 -501 1668 -501 0 1
rlabel polysilicon 1668 -507 1668 -507 0 3
rlabel polysilicon 1675 -501 1675 -501 0 1
rlabel polysilicon 1675 -507 1675 -507 0 3
rlabel polysilicon 1682 -501 1682 -501 0 1
rlabel polysilicon 1682 -507 1682 -507 0 3
rlabel polysilicon 1689 -501 1689 -501 0 1
rlabel polysilicon 1689 -507 1689 -507 0 3
rlabel polysilicon 1696 -501 1696 -501 0 1
rlabel polysilicon 1696 -507 1696 -507 0 3
rlabel polysilicon 1703 -501 1703 -501 0 1
rlabel polysilicon 1703 -507 1703 -507 0 3
rlabel polysilicon 1710 -501 1710 -501 0 1
rlabel polysilicon 1710 -507 1710 -507 0 3
rlabel polysilicon 1717 -501 1717 -501 0 1
rlabel polysilicon 1717 -507 1717 -507 0 3
rlabel polysilicon 1724 -501 1724 -501 0 1
rlabel polysilicon 1724 -507 1724 -507 0 3
rlabel polysilicon 1731 -501 1731 -501 0 1
rlabel polysilicon 1731 -507 1731 -507 0 3
rlabel polysilicon 1738 -501 1738 -501 0 1
rlabel polysilicon 1738 -507 1738 -507 0 3
rlabel polysilicon 1745 -501 1745 -501 0 1
rlabel polysilicon 1745 -507 1745 -507 0 3
rlabel polysilicon 1752 -501 1752 -501 0 1
rlabel polysilicon 1752 -507 1752 -507 0 3
rlabel polysilicon 1759 -501 1759 -501 0 1
rlabel polysilicon 1759 -507 1759 -507 0 3
rlabel polysilicon 1766 -501 1766 -501 0 1
rlabel polysilicon 1766 -507 1766 -507 0 3
rlabel polysilicon 1773 -501 1773 -501 0 1
rlabel polysilicon 1773 -507 1773 -507 0 3
rlabel polysilicon 1780 -501 1780 -501 0 1
rlabel polysilicon 1780 -507 1780 -507 0 3
rlabel polysilicon 1787 -501 1787 -501 0 1
rlabel polysilicon 1787 -507 1787 -507 0 3
rlabel polysilicon 1794 -501 1794 -501 0 1
rlabel polysilicon 1794 -507 1794 -507 0 3
rlabel polysilicon 1801 -501 1801 -501 0 1
rlabel polysilicon 1801 -507 1801 -507 0 3
rlabel polysilicon 1808 -501 1808 -501 0 1
rlabel polysilicon 1808 -507 1808 -507 0 3
rlabel polysilicon 1815 -501 1815 -501 0 1
rlabel polysilicon 1815 -507 1815 -507 0 3
rlabel polysilicon 1822 -501 1822 -501 0 1
rlabel polysilicon 1822 -507 1822 -507 0 3
rlabel polysilicon 1829 -501 1829 -501 0 1
rlabel polysilicon 1829 -507 1829 -507 0 3
rlabel polysilicon 1836 -501 1836 -501 0 1
rlabel polysilicon 1836 -507 1836 -507 0 3
rlabel polysilicon 1843 -501 1843 -501 0 1
rlabel polysilicon 1843 -507 1843 -507 0 3
rlabel polysilicon 1850 -501 1850 -501 0 1
rlabel polysilicon 1850 -507 1850 -507 0 3
rlabel polysilicon 1857 -501 1857 -501 0 1
rlabel polysilicon 1857 -507 1857 -507 0 3
rlabel polysilicon 1864 -501 1864 -501 0 1
rlabel polysilicon 1864 -507 1864 -507 0 3
rlabel polysilicon 1871 -501 1871 -501 0 1
rlabel polysilicon 1871 -507 1871 -507 0 3
rlabel polysilicon 1878 -501 1878 -501 0 1
rlabel polysilicon 1878 -507 1878 -507 0 3
rlabel polysilicon 1885 -501 1885 -501 0 1
rlabel polysilicon 1885 -507 1885 -507 0 3
rlabel polysilicon 1892 -501 1892 -501 0 1
rlabel polysilicon 1892 -507 1892 -507 0 3
rlabel polysilicon 1899 -501 1899 -501 0 1
rlabel polysilicon 1899 -507 1899 -507 0 3
rlabel polysilicon 1906 -501 1906 -501 0 1
rlabel polysilicon 1906 -507 1906 -507 0 3
rlabel polysilicon 1913 -501 1913 -501 0 1
rlabel polysilicon 1913 -507 1913 -507 0 3
rlabel polysilicon 1920 -501 1920 -501 0 1
rlabel polysilicon 1920 -507 1920 -507 0 3
rlabel polysilicon 1927 -501 1927 -501 0 1
rlabel polysilicon 1927 -507 1927 -507 0 3
rlabel polysilicon 1934 -501 1934 -501 0 1
rlabel polysilicon 1934 -507 1934 -507 0 3
rlabel polysilicon 1941 -501 1941 -501 0 1
rlabel polysilicon 1941 -507 1941 -507 0 3
rlabel polysilicon 1948 -501 1948 -501 0 1
rlabel polysilicon 1948 -507 1948 -507 0 3
rlabel polysilicon 1955 -501 1955 -501 0 1
rlabel polysilicon 1958 -501 1958 -501 0 2
rlabel polysilicon 1955 -507 1955 -507 0 3
rlabel polysilicon 1958 -507 1958 -507 0 4
rlabel polysilicon 1962 -501 1962 -501 0 1
rlabel polysilicon 1962 -507 1962 -507 0 3
rlabel polysilicon 1969 -501 1969 -501 0 1
rlabel polysilicon 1969 -507 1969 -507 0 3
rlabel polysilicon 1976 -501 1976 -501 0 1
rlabel polysilicon 1976 -507 1976 -507 0 3
rlabel polysilicon 1979 -507 1979 -507 0 4
rlabel polysilicon 1983 -501 1983 -501 0 1
rlabel polysilicon 1983 -507 1983 -507 0 3
rlabel polysilicon 1990 -501 1990 -501 0 1
rlabel polysilicon 1990 -507 1990 -507 0 3
rlabel polysilicon 1997 -501 1997 -501 0 1
rlabel polysilicon 1997 -507 1997 -507 0 3
rlabel polysilicon 2007 -507 2007 -507 0 4
rlabel polysilicon 2011 -501 2011 -501 0 1
rlabel polysilicon 2011 -507 2011 -507 0 3
rlabel polysilicon 2014 -507 2014 -507 0 4
rlabel polysilicon 2018 -507 2018 -507 0 3
rlabel polysilicon 2021 -507 2021 -507 0 4
rlabel polysilicon 2039 -501 2039 -501 0 1
rlabel polysilicon 2039 -507 2039 -507 0 3
rlabel polysilicon 2088 -501 2088 -501 0 1
rlabel polysilicon 2088 -507 2088 -507 0 3
rlabel polysilicon 2116 -501 2116 -501 0 1
rlabel polysilicon 2116 -507 2116 -507 0 3
rlabel polysilicon 2144 -501 2144 -501 0 1
rlabel polysilicon 2144 -507 2144 -507 0 3
rlabel polysilicon 2263 -501 2263 -501 0 1
rlabel polysilicon 2263 -507 2263 -507 0 3
rlabel polysilicon 2284 -501 2284 -501 0 1
rlabel polysilicon 2284 -507 2284 -507 0 3
rlabel polysilicon 5 -640 5 -640 0 4
rlabel polysilicon 9 -634 9 -634 0 1
rlabel polysilicon 9 -640 9 -640 0 3
rlabel polysilicon 16 -634 16 -634 0 1
rlabel polysilicon 16 -640 16 -640 0 3
rlabel polysilicon 23 -634 23 -634 0 1
rlabel polysilicon 23 -640 23 -640 0 3
rlabel polysilicon 30 -634 30 -634 0 1
rlabel polysilicon 30 -640 30 -640 0 3
rlabel polysilicon 37 -634 37 -634 0 1
rlabel polysilicon 37 -640 37 -640 0 3
rlabel polysilicon 44 -634 44 -634 0 1
rlabel polysilicon 44 -640 44 -640 0 3
rlabel polysilicon 51 -634 51 -634 0 1
rlabel polysilicon 51 -640 51 -640 0 3
rlabel polysilicon 58 -634 58 -634 0 1
rlabel polysilicon 61 -634 61 -634 0 2
rlabel polysilicon 58 -640 58 -640 0 3
rlabel polysilicon 65 -634 65 -634 0 1
rlabel polysilicon 65 -640 65 -640 0 3
rlabel polysilicon 72 -634 72 -634 0 1
rlabel polysilicon 75 -634 75 -634 0 2
rlabel polysilicon 72 -640 72 -640 0 3
rlabel polysilicon 75 -640 75 -640 0 4
rlabel polysilicon 79 -634 79 -634 0 1
rlabel polysilicon 79 -640 79 -640 0 3
rlabel polysilicon 86 -634 86 -634 0 1
rlabel polysilicon 86 -640 86 -640 0 3
rlabel polysilicon 93 -634 93 -634 0 1
rlabel polysilicon 93 -640 93 -640 0 3
rlabel polysilicon 100 -634 100 -634 0 1
rlabel polysilicon 103 -634 103 -634 0 2
rlabel polysilicon 100 -640 100 -640 0 3
rlabel polysilicon 107 -634 107 -634 0 1
rlabel polysilicon 107 -640 107 -640 0 3
rlabel polysilicon 114 -634 114 -634 0 1
rlabel polysilicon 114 -640 114 -640 0 3
rlabel polysilicon 121 -634 121 -634 0 1
rlabel polysilicon 121 -640 121 -640 0 3
rlabel polysilicon 128 -634 128 -634 0 1
rlabel polysilicon 128 -640 128 -640 0 3
rlabel polysilicon 135 -634 135 -634 0 1
rlabel polysilicon 138 -634 138 -634 0 2
rlabel polysilicon 135 -640 135 -640 0 3
rlabel polysilicon 142 -634 142 -634 0 1
rlabel polysilicon 142 -640 142 -640 0 3
rlabel polysilicon 149 -634 149 -634 0 1
rlabel polysilicon 149 -640 149 -640 0 3
rlabel polysilicon 156 -634 156 -634 0 1
rlabel polysilicon 156 -640 156 -640 0 3
rlabel polysilicon 163 -634 163 -634 0 1
rlabel polysilicon 163 -640 163 -640 0 3
rlabel polysilicon 173 -634 173 -634 0 2
rlabel polysilicon 173 -640 173 -640 0 4
rlabel polysilicon 177 -634 177 -634 0 1
rlabel polysilicon 177 -640 177 -640 0 3
rlabel polysilicon 184 -634 184 -634 0 1
rlabel polysilicon 184 -640 184 -640 0 3
rlabel polysilicon 191 -634 191 -634 0 1
rlabel polysilicon 191 -640 191 -640 0 3
rlabel polysilicon 198 -634 198 -634 0 1
rlabel polysilicon 198 -640 198 -640 0 3
rlabel polysilicon 205 -634 205 -634 0 1
rlabel polysilicon 205 -640 205 -640 0 3
rlabel polysilicon 208 -640 208 -640 0 4
rlabel polysilicon 212 -634 212 -634 0 1
rlabel polysilicon 212 -640 212 -640 0 3
rlabel polysilicon 219 -634 219 -634 0 1
rlabel polysilicon 219 -640 219 -640 0 3
rlabel polysilicon 226 -634 226 -634 0 1
rlabel polysilicon 226 -640 226 -640 0 3
rlabel polysilicon 233 -634 233 -634 0 1
rlabel polysilicon 233 -640 233 -640 0 3
rlabel polysilicon 240 -634 240 -634 0 1
rlabel polysilicon 240 -640 240 -640 0 3
rlabel polysilicon 247 -634 247 -634 0 1
rlabel polysilicon 250 -634 250 -634 0 2
rlabel polysilicon 250 -640 250 -640 0 4
rlabel polysilicon 254 -634 254 -634 0 1
rlabel polysilicon 254 -640 254 -640 0 3
rlabel polysilicon 261 -634 261 -634 0 1
rlabel polysilicon 261 -640 261 -640 0 3
rlabel polysilicon 268 -634 268 -634 0 1
rlabel polysilicon 268 -640 268 -640 0 3
rlabel polysilicon 275 -634 275 -634 0 1
rlabel polysilicon 275 -640 275 -640 0 3
rlabel polysilicon 282 -634 282 -634 0 1
rlabel polysilicon 282 -640 282 -640 0 3
rlabel polysilicon 289 -634 289 -634 0 1
rlabel polysilicon 289 -640 289 -640 0 3
rlabel polysilicon 296 -634 296 -634 0 1
rlabel polysilicon 296 -640 296 -640 0 3
rlabel polysilicon 303 -634 303 -634 0 1
rlabel polysilicon 303 -640 303 -640 0 3
rlabel polysilicon 310 -634 310 -634 0 1
rlabel polysilicon 310 -640 310 -640 0 3
rlabel polysilicon 317 -634 317 -634 0 1
rlabel polysilicon 317 -640 317 -640 0 3
rlabel polysilicon 324 -634 324 -634 0 1
rlabel polysilicon 324 -640 324 -640 0 3
rlabel polysilicon 331 -634 331 -634 0 1
rlabel polysilicon 331 -640 331 -640 0 3
rlabel polysilicon 338 -634 338 -634 0 1
rlabel polysilicon 338 -640 338 -640 0 3
rlabel polysilicon 345 -634 345 -634 0 1
rlabel polysilicon 345 -640 345 -640 0 3
rlabel polysilicon 352 -634 352 -634 0 1
rlabel polysilicon 352 -640 352 -640 0 3
rlabel polysilicon 359 -634 359 -634 0 1
rlabel polysilicon 359 -640 359 -640 0 3
rlabel polysilicon 366 -634 366 -634 0 1
rlabel polysilicon 366 -640 366 -640 0 3
rlabel polysilicon 373 -634 373 -634 0 1
rlabel polysilicon 373 -640 373 -640 0 3
rlabel polysilicon 380 -634 380 -634 0 1
rlabel polysilicon 380 -640 380 -640 0 3
rlabel polysilicon 387 -634 387 -634 0 1
rlabel polysilicon 387 -640 387 -640 0 3
rlabel polysilicon 394 -634 394 -634 0 1
rlabel polysilicon 394 -640 394 -640 0 3
rlabel polysilicon 401 -634 401 -634 0 1
rlabel polysilicon 401 -640 401 -640 0 3
rlabel polysilicon 408 -634 408 -634 0 1
rlabel polysilicon 408 -640 408 -640 0 3
rlabel polysilicon 415 -634 415 -634 0 1
rlabel polysilicon 415 -640 415 -640 0 3
rlabel polysilicon 422 -634 422 -634 0 1
rlabel polysilicon 422 -640 422 -640 0 3
rlabel polysilicon 429 -634 429 -634 0 1
rlabel polysilicon 432 -634 432 -634 0 2
rlabel polysilicon 429 -640 429 -640 0 3
rlabel polysilicon 432 -640 432 -640 0 4
rlabel polysilicon 436 -634 436 -634 0 1
rlabel polysilicon 436 -640 436 -640 0 3
rlabel polysilicon 443 -634 443 -634 0 1
rlabel polysilicon 443 -640 443 -640 0 3
rlabel polysilicon 450 -634 450 -634 0 1
rlabel polysilicon 450 -640 450 -640 0 3
rlabel polysilicon 457 -634 457 -634 0 1
rlabel polysilicon 457 -640 457 -640 0 3
rlabel polysilicon 464 -634 464 -634 0 1
rlabel polysilicon 464 -640 464 -640 0 3
rlabel polysilicon 471 -634 471 -634 0 1
rlabel polysilicon 471 -640 471 -640 0 3
rlabel polysilicon 478 -634 478 -634 0 1
rlabel polysilicon 478 -640 478 -640 0 3
rlabel polysilicon 485 -634 485 -634 0 1
rlabel polysilicon 485 -640 485 -640 0 3
rlabel polysilicon 492 -634 492 -634 0 1
rlabel polysilicon 492 -640 492 -640 0 3
rlabel polysilicon 499 -634 499 -634 0 1
rlabel polysilicon 499 -640 499 -640 0 3
rlabel polysilicon 506 -634 506 -634 0 1
rlabel polysilicon 506 -640 506 -640 0 3
rlabel polysilicon 513 -634 513 -634 0 1
rlabel polysilicon 513 -640 513 -640 0 3
rlabel polysilicon 520 -634 520 -634 0 1
rlabel polysilicon 520 -640 520 -640 0 3
rlabel polysilicon 527 -634 527 -634 0 1
rlabel polysilicon 527 -640 527 -640 0 3
rlabel polysilicon 537 -634 537 -634 0 2
rlabel polysilicon 534 -640 534 -640 0 3
rlabel polysilicon 537 -640 537 -640 0 4
rlabel polysilicon 541 -634 541 -634 0 1
rlabel polysilicon 541 -640 541 -640 0 3
rlabel polysilicon 548 -634 548 -634 0 1
rlabel polysilicon 548 -640 548 -640 0 3
rlabel polysilicon 555 -634 555 -634 0 1
rlabel polysilicon 555 -640 555 -640 0 3
rlabel polysilicon 562 -634 562 -634 0 1
rlabel polysilicon 565 -634 565 -634 0 2
rlabel polysilicon 562 -640 562 -640 0 3
rlabel polysilicon 565 -640 565 -640 0 4
rlabel polysilicon 569 -634 569 -634 0 1
rlabel polysilicon 569 -640 569 -640 0 3
rlabel polysilicon 576 -634 576 -634 0 1
rlabel polysilicon 576 -640 576 -640 0 3
rlabel polysilicon 583 -634 583 -634 0 1
rlabel polysilicon 586 -634 586 -634 0 2
rlabel polysilicon 583 -640 583 -640 0 3
rlabel polysilicon 586 -640 586 -640 0 4
rlabel polysilicon 590 -634 590 -634 0 1
rlabel polysilicon 593 -634 593 -634 0 2
rlabel polysilicon 590 -640 590 -640 0 3
rlabel polysilicon 597 -634 597 -634 0 1
rlabel polysilicon 597 -640 597 -640 0 3
rlabel polysilicon 604 -634 604 -634 0 1
rlabel polysilicon 604 -640 604 -640 0 3
rlabel polysilicon 611 -634 611 -634 0 1
rlabel polysilicon 611 -640 611 -640 0 3
rlabel polysilicon 618 -634 618 -634 0 1
rlabel polysilicon 618 -640 618 -640 0 3
rlabel polysilicon 625 -634 625 -634 0 1
rlabel polysilicon 625 -640 625 -640 0 3
rlabel polysilicon 632 -634 632 -634 0 1
rlabel polysilicon 632 -640 632 -640 0 3
rlabel polysilicon 639 -634 639 -634 0 1
rlabel polysilicon 639 -640 639 -640 0 3
rlabel polysilicon 649 -634 649 -634 0 2
rlabel polysilicon 646 -640 646 -640 0 3
rlabel polysilicon 649 -640 649 -640 0 4
rlabel polysilicon 653 -634 653 -634 0 1
rlabel polysilicon 653 -640 653 -640 0 3
rlabel polysilicon 660 -634 660 -634 0 1
rlabel polysilicon 663 -634 663 -634 0 2
rlabel polysilicon 660 -640 660 -640 0 3
rlabel polysilicon 663 -640 663 -640 0 4
rlabel polysilicon 667 -634 667 -634 0 1
rlabel polysilicon 667 -640 667 -640 0 3
rlabel polysilicon 674 -634 674 -634 0 1
rlabel polysilicon 674 -640 674 -640 0 3
rlabel polysilicon 681 -634 681 -634 0 1
rlabel polysilicon 681 -640 681 -640 0 3
rlabel polysilicon 688 -634 688 -634 0 1
rlabel polysilicon 688 -640 688 -640 0 3
rlabel polysilicon 695 -634 695 -634 0 1
rlabel polysilicon 695 -640 695 -640 0 3
rlabel polysilicon 702 -634 702 -634 0 1
rlabel polysilicon 702 -640 702 -640 0 3
rlabel polysilicon 709 -634 709 -634 0 1
rlabel polysilicon 709 -640 709 -640 0 3
rlabel polysilicon 716 -634 716 -634 0 1
rlabel polysilicon 716 -640 716 -640 0 3
rlabel polysilicon 723 -634 723 -634 0 1
rlabel polysilicon 723 -640 723 -640 0 3
rlabel polysilicon 730 -634 730 -634 0 1
rlabel polysilicon 733 -634 733 -634 0 2
rlabel polysilicon 730 -640 730 -640 0 3
rlabel polysilicon 733 -640 733 -640 0 4
rlabel polysilicon 737 -634 737 -634 0 1
rlabel polysilicon 737 -640 737 -640 0 3
rlabel polysilicon 744 -634 744 -634 0 1
rlabel polysilicon 744 -640 744 -640 0 3
rlabel polysilicon 747 -640 747 -640 0 4
rlabel polysilicon 751 -634 751 -634 0 1
rlabel polysilicon 751 -640 751 -640 0 3
rlabel polysilicon 758 -634 758 -634 0 1
rlabel polysilicon 758 -640 758 -640 0 3
rlabel polysilicon 765 -634 765 -634 0 1
rlabel polysilicon 765 -640 765 -640 0 3
rlabel polysilicon 772 -634 772 -634 0 1
rlabel polysilicon 772 -640 772 -640 0 3
rlabel polysilicon 779 -634 779 -634 0 1
rlabel polysilicon 779 -640 779 -640 0 3
rlabel polysilicon 786 -634 786 -634 0 1
rlabel polysilicon 789 -640 789 -640 0 4
rlabel polysilicon 793 -634 793 -634 0 1
rlabel polysilicon 793 -640 793 -640 0 3
rlabel polysilicon 800 -634 800 -634 0 1
rlabel polysilicon 800 -640 800 -640 0 3
rlabel polysilicon 810 -634 810 -634 0 2
rlabel polysilicon 807 -640 807 -640 0 3
rlabel polysilicon 810 -640 810 -640 0 4
rlabel polysilicon 814 -634 814 -634 0 1
rlabel polysilicon 814 -640 814 -640 0 3
rlabel polysilicon 821 -634 821 -634 0 1
rlabel polysilicon 824 -634 824 -634 0 2
rlabel polysilicon 821 -640 821 -640 0 3
rlabel polysilicon 824 -640 824 -640 0 4
rlabel polysilicon 828 -634 828 -634 0 1
rlabel polysilicon 828 -640 828 -640 0 3
rlabel polysilicon 835 -634 835 -634 0 1
rlabel polysilicon 835 -640 835 -640 0 3
rlabel polysilicon 842 -634 842 -634 0 1
rlabel polysilicon 842 -640 842 -640 0 3
rlabel polysilicon 849 -634 849 -634 0 1
rlabel polysilicon 852 -634 852 -634 0 2
rlabel polysilicon 849 -640 849 -640 0 3
rlabel polysilicon 852 -640 852 -640 0 4
rlabel polysilicon 856 -634 856 -634 0 1
rlabel polysilicon 856 -640 856 -640 0 3
rlabel polysilicon 863 -634 863 -634 0 1
rlabel polysilicon 863 -640 863 -640 0 3
rlabel polysilicon 870 -634 870 -634 0 1
rlabel polysilicon 870 -640 870 -640 0 3
rlabel polysilicon 877 -634 877 -634 0 1
rlabel polysilicon 877 -640 877 -640 0 3
rlabel polysilicon 884 -634 884 -634 0 1
rlabel polysilicon 884 -640 884 -640 0 3
rlabel polysilicon 891 -634 891 -634 0 1
rlabel polysilicon 891 -640 891 -640 0 3
rlabel polysilicon 898 -634 898 -634 0 1
rlabel polysilicon 898 -640 898 -640 0 3
rlabel polysilicon 905 -634 905 -634 0 1
rlabel polysilicon 905 -640 905 -640 0 3
rlabel polysilicon 912 -634 912 -634 0 1
rlabel polysilicon 912 -640 912 -640 0 3
rlabel polysilicon 919 -634 919 -634 0 1
rlabel polysilicon 919 -640 919 -640 0 3
rlabel polysilicon 926 -634 926 -634 0 1
rlabel polysilicon 929 -634 929 -634 0 2
rlabel polysilicon 926 -640 926 -640 0 3
rlabel polysilicon 929 -640 929 -640 0 4
rlabel polysilicon 933 -634 933 -634 0 1
rlabel polysilicon 933 -640 933 -640 0 3
rlabel polysilicon 940 -634 940 -634 0 1
rlabel polysilicon 940 -640 940 -640 0 3
rlabel polysilicon 943 -640 943 -640 0 4
rlabel polysilicon 947 -634 947 -634 0 1
rlabel polysilicon 947 -640 947 -640 0 3
rlabel polysilicon 954 -634 954 -634 0 1
rlabel polysilicon 954 -640 954 -640 0 3
rlabel polysilicon 961 -634 961 -634 0 1
rlabel polysilicon 961 -640 961 -640 0 3
rlabel polysilicon 968 -634 968 -634 0 1
rlabel polysilicon 968 -640 968 -640 0 3
rlabel polysilicon 975 -634 975 -634 0 1
rlabel polysilicon 975 -640 975 -640 0 3
rlabel polysilicon 985 -634 985 -634 0 2
rlabel polysilicon 985 -640 985 -640 0 4
rlabel polysilicon 989 -634 989 -634 0 1
rlabel polysilicon 989 -640 989 -640 0 3
rlabel polysilicon 996 -634 996 -634 0 1
rlabel polysilicon 996 -640 996 -640 0 3
rlabel polysilicon 1003 -634 1003 -634 0 1
rlabel polysilicon 1003 -640 1003 -640 0 3
rlabel polysilicon 1010 -634 1010 -634 0 1
rlabel polysilicon 1013 -634 1013 -634 0 2
rlabel polysilicon 1010 -640 1010 -640 0 3
rlabel polysilicon 1017 -634 1017 -634 0 1
rlabel polysilicon 1017 -640 1017 -640 0 3
rlabel polysilicon 1024 -634 1024 -634 0 1
rlabel polysilicon 1024 -640 1024 -640 0 3
rlabel polysilicon 1031 -634 1031 -634 0 1
rlabel polysilicon 1034 -634 1034 -634 0 2
rlabel polysilicon 1031 -640 1031 -640 0 3
rlabel polysilicon 1038 -634 1038 -634 0 1
rlabel polysilicon 1038 -640 1038 -640 0 3
rlabel polysilicon 1045 -634 1045 -634 0 1
rlabel polysilicon 1045 -640 1045 -640 0 3
rlabel polysilicon 1052 -634 1052 -634 0 1
rlabel polysilicon 1052 -640 1052 -640 0 3
rlabel polysilicon 1059 -634 1059 -634 0 1
rlabel polysilicon 1062 -634 1062 -634 0 2
rlabel polysilicon 1059 -640 1059 -640 0 3
rlabel polysilicon 1062 -640 1062 -640 0 4
rlabel polysilicon 1066 -634 1066 -634 0 1
rlabel polysilicon 1066 -640 1066 -640 0 3
rlabel polysilicon 1073 -634 1073 -634 0 1
rlabel polysilicon 1073 -640 1073 -640 0 3
rlabel polysilicon 1080 -634 1080 -634 0 1
rlabel polysilicon 1080 -640 1080 -640 0 3
rlabel polysilicon 1083 -640 1083 -640 0 4
rlabel polysilicon 1087 -634 1087 -634 0 1
rlabel polysilicon 1087 -640 1087 -640 0 3
rlabel polysilicon 1094 -634 1094 -634 0 1
rlabel polysilicon 1094 -640 1094 -640 0 3
rlabel polysilicon 1097 -640 1097 -640 0 4
rlabel polysilicon 1101 -634 1101 -634 0 1
rlabel polysilicon 1101 -640 1101 -640 0 3
rlabel polysilicon 1108 -634 1108 -634 0 1
rlabel polysilicon 1108 -640 1108 -640 0 3
rlabel polysilicon 1115 -634 1115 -634 0 1
rlabel polysilicon 1115 -640 1115 -640 0 3
rlabel polysilicon 1122 -634 1122 -634 0 1
rlabel polysilicon 1122 -640 1122 -640 0 3
rlabel polysilicon 1129 -634 1129 -634 0 1
rlabel polysilicon 1129 -640 1129 -640 0 3
rlabel polysilicon 1136 -634 1136 -634 0 1
rlabel polysilicon 1136 -640 1136 -640 0 3
rlabel polysilicon 1143 -634 1143 -634 0 1
rlabel polysilicon 1146 -634 1146 -634 0 2
rlabel polysilicon 1143 -640 1143 -640 0 3
rlabel polysilicon 1146 -640 1146 -640 0 4
rlabel polysilicon 1150 -634 1150 -634 0 1
rlabel polysilicon 1150 -640 1150 -640 0 3
rlabel polysilicon 1153 -640 1153 -640 0 4
rlabel polysilicon 1157 -634 1157 -634 0 1
rlabel polysilicon 1157 -640 1157 -640 0 3
rlabel polysilicon 1164 -634 1164 -634 0 1
rlabel polysilicon 1164 -640 1164 -640 0 3
rlabel polysilicon 1171 -634 1171 -634 0 1
rlabel polysilicon 1171 -640 1171 -640 0 3
rlabel polysilicon 1178 -634 1178 -634 0 1
rlabel polysilicon 1178 -640 1178 -640 0 3
rlabel polysilicon 1185 -634 1185 -634 0 1
rlabel polysilicon 1185 -640 1185 -640 0 3
rlabel polysilicon 1192 -634 1192 -634 0 1
rlabel polysilicon 1192 -640 1192 -640 0 3
rlabel polysilicon 1199 -634 1199 -634 0 1
rlabel polysilicon 1202 -634 1202 -634 0 2
rlabel polysilicon 1199 -640 1199 -640 0 3
rlabel polysilicon 1202 -640 1202 -640 0 4
rlabel polysilicon 1206 -634 1206 -634 0 1
rlabel polysilicon 1206 -640 1206 -640 0 3
rlabel polysilicon 1213 -634 1213 -634 0 1
rlabel polysilicon 1216 -634 1216 -634 0 2
rlabel polysilicon 1213 -640 1213 -640 0 3
rlabel polysilicon 1216 -640 1216 -640 0 4
rlabel polysilicon 1220 -634 1220 -634 0 1
rlabel polysilicon 1220 -640 1220 -640 0 3
rlabel polysilicon 1227 -634 1227 -634 0 1
rlabel polysilicon 1227 -640 1227 -640 0 3
rlabel polysilicon 1234 -634 1234 -634 0 1
rlabel polysilicon 1234 -640 1234 -640 0 3
rlabel polysilicon 1241 -634 1241 -634 0 1
rlabel polysilicon 1241 -640 1241 -640 0 3
rlabel polysilicon 1248 -634 1248 -634 0 1
rlabel polysilicon 1248 -640 1248 -640 0 3
rlabel polysilicon 1255 -634 1255 -634 0 1
rlabel polysilicon 1255 -640 1255 -640 0 3
rlabel polysilicon 1262 -634 1262 -634 0 1
rlabel polysilicon 1262 -640 1262 -640 0 3
rlabel polysilicon 1269 -634 1269 -634 0 1
rlabel polysilicon 1269 -640 1269 -640 0 3
rlabel polysilicon 1276 -634 1276 -634 0 1
rlabel polysilicon 1276 -640 1276 -640 0 3
rlabel polysilicon 1283 -634 1283 -634 0 1
rlabel polysilicon 1283 -640 1283 -640 0 3
rlabel polysilicon 1290 -634 1290 -634 0 1
rlabel polysilicon 1290 -640 1290 -640 0 3
rlabel polysilicon 1297 -634 1297 -634 0 1
rlabel polysilicon 1297 -640 1297 -640 0 3
rlabel polysilicon 1300 -640 1300 -640 0 4
rlabel polysilicon 1304 -634 1304 -634 0 1
rlabel polysilicon 1304 -640 1304 -640 0 3
rlabel polysilicon 1311 -634 1311 -634 0 1
rlabel polysilicon 1311 -640 1311 -640 0 3
rlabel polysilicon 1318 -634 1318 -634 0 1
rlabel polysilicon 1318 -640 1318 -640 0 3
rlabel polysilicon 1325 -634 1325 -634 0 1
rlabel polysilicon 1325 -640 1325 -640 0 3
rlabel polysilicon 1332 -634 1332 -634 0 1
rlabel polysilicon 1332 -640 1332 -640 0 3
rlabel polysilicon 1339 -634 1339 -634 0 1
rlabel polysilicon 1339 -640 1339 -640 0 3
rlabel polysilicon 1346 -634 1346 -634 0 1
rlabel polysilicon 1346 -640 1346 -640 0 3
rlabel polysilicon 1353 -634 1353 -634 0 1
rlabel polysilicon 1353 -640 1353 -640 0 3
rlabel polysilicon 1360 -634 1360 -634 0 1
rlabel polysilicon 1360 -640 1360 -640 0 3
rlabel polysilicon 1367 -634 1367 -634 0 1
rlabel polysilicon 1367 -640 1367 -640 0 3
rlabel polysilicon 1374 -634 1374 -634 0 1
rlabel polysilicon 1374 -640 1374 -640 0 3
rlabel polysilicon 1381 -634 1381 -634 0 1
rlabel polysilicon 1381 -640 1381 -640 0 3
rlabel polysilicon 1388 -634 1388 -634 0 1
rlabel polysilicon 1388 -640 1388 -640 0 3
rlabel polysilicon 1395 -634 1395 -634 0 1
rlabel polysilicon 1395 -640 1395 -640 0 3
rlabel polysilicon 1402 -634 1402 -634 0 1
rlabel polysilicon 1402 -640 1402 -640 0 3
rlabel polysilicon 1409 -634 1409 -634 0 1
rlabel polysilicon 1409 -640 1409 -640 0 3
rlabel polysilicon 1416 -634 1416 -634 0 1
rlabel polysilicon 1416 -640 1416 -640 0 3
rlabel polysilicon 1423 -634 1423 -634 0 1
rlabel polysilicon 1423 -640 1423 -640 0 3
rlabel polysilicon 1430 -634 1430 -634 0 1
rlabel polysilicon 1430 -640 1430 -640 0 3
rlabel polysilicon 1437 -634 1437 -634 0 1
rlabel polysilicon 1437 -640 1437 -640 0 3
rlabel polysilicon 1444 -634 1444 -634 0 1
rlabel polysilicon 1444 -640 1444 -640 0 3
rlabel polysilicon 1451 -634 1451 -634 0 1
rlabel polysilicon 1451 -640 1451 -640 0 3
rlabel polysilicon 1458 -634 1458 -634 0 1
rlabel polysilicon 1458 -640 1458 -640 0 3
rlabel polysilicon 1465 -634 1465 -634 0 1
rlabel polysilicon 1465 -640 1465 -640 0 3
rlabel polysilicon 1472 -634 1472 -634 0 1
rlabel polysilicon 1472 -640 1472 -640 0 3
rlabel polysilicon 1479 -634 1479 -634 0 1
rlabel polysilicon 1479 -640 1479 -640 0 3
rlabel polysilicon 1489 -634 1489 -634 0 2
rlabel polysilicon 1486 -640 1486 -640 0 3
rlabel polysilicon 1493 -634 1493 -634 0 1
rlabel polysilicon 1493 -640 1493 -640 0 3
rlabel polysilicon 1500 -634 1500 -634 0 1
rlabel polysilicon 1500 -640 1500 -640 0 3
rlabel polysilicon 1507 -634 1507 -634 0 1
rlabel polysilicon 1507 -640 1507 -640 0 3
rlabel polysilicon 1514 -634 1514 -634 0 1
rlabel polysilicon 1514 -640 1514 -640 0 3
rlabel polysilicon 1521 -634 1521 -634 0 1
rlabel polysilicon 1521 -640 1521 -640 0 3
rlabel polysilicon 1528 -634 1528 -634 0 1
rlabel polysilicon 1528 -640 1528 -640 0 3
rlabel polysilicon 1535 -634 1535 -634 0 1
rlabel polysilicon 1535 -640 1535 -640 0 3
rlabel polysilicon 1542 -634 1542 -634 0 1
rlabel polysilicon 1542 -640 1542 -640 0 3
rlabel polysilicon 1549 -634 1549 -634 0 1
rlabel polysilicon 1549 -640 1549 -640 0 3
rlabel polysilicon 1556 -634 1556 -634 0 1
rlabel polysilicon 1556 -640 1556 -640 0 3
rlabel polysilicon 1563 -634 1563 -634 0 1
rlabel polysilicon 1563 -640 1563 -640 0 3
rlabel polysilicon 1570 -634 1570 -634 0 1
rlabel polysilicon 1570 -640 1570 -640 0 3
rlabel polysilicon 1577 -634 1577 -634 0 1
rlabel polysilicon 1577 -640 1577 -640 0 3
rlabel polysilicon 1584 -634 1584 -634 0 1
rlabel polysilicon 1584 -640 1584 -640 0 3
rlabel polysilicon 1591 -634 1591 -634 0 1
rlabel polysilicon 1591 -640 1591 -640 0 3
rlabel polysilicon 1598 -634 1598 -634 0 1
rlabel polysilicon 1598 -640 1598 -640 0 3
rlabel polysilicon 1605 -634 1605 -634 0 1
rlabel polysilicon 1605 -640 1605 -640 0 3
rlabel polysilicon 1612 -634 1612 -634 0 1
rlabel polysilicon 1612 -640 1612 -640 0 3
rlabel polysilicon 1619 -634 1619 -634 0 1
rlabel polysilicon 1619 -640 1619 -640 0 3
rlabel polysilicon 1626 -634 1626 -634 0 1
rlabel polysilicon 1626 -640 1626 -640 0 3
rlabel polysilicon 1633 -634 1633 -634 0 1
rlabel polysilicon 1633 -640 1633 -640 0 3
rlabel polysilicon 1640 -634 1640 -634 0 1
rlabel polysilicon 1640 -640 1640 -640 0 3
rlabel polysilicon 1647 -634 1647 -634 0 1
rlabel polysilicon 1647 -640 1647 -640 0 3
rlabel polysilicon 1654 -634 1654 -634 0 1
rlabel polysilicon 1654 -640 1654 -640 0 3
rlabel polysilicon 1661 -634 1661 -634 0 1
rlabel polysilicon 1661 -640 1661 -640 0 3
rlabel polysilicon 1668 -634 1668 -634 0 1
rlabel polysilicon 1668 -640 1668 -640 0 3
rlabel polysilicon 1675 -634 1675 -634 0 1
rlabel polysilicon 1675 -640 1675 -640 0 3
rlabel polysilicon 1682 -634 1682 -634 0 1
rlabel polysilicon 1682 -640 1682 -640 0 3
rlabel polysilicon 1689 -634 1689 -634 0 1
rlabel polysilicon 1689 -640 1689 -640 0 3
rlabel polysilicon 1696 -634 1696 -634 0 1
rlabel polysilicon 1696 -640 1696 -640 0 3
rlabel polysilicon 1703 -634 1703 -634 0 1
rlabel polysilicon 1703 -640 1703 -640 0 3
rlabel polysilicon 1710 -634 1710 -634 0 1
rlabel polysilicon 1710 -640 1710 -640 0 3
rlabel polysilicon 1717 -634 1717 -634 0 1
rlabel polysilicon 1717 -640 1717 -640 0 3
rlabel polysilicon 1724 -634 1724 -634 0 1
rlabel polysilicon 1724 -640 1724 -640 0 3
rlabel polysilicon 1731 -634 1731 -634 0 1
rlabel polysilicon 1731 -640 1731 -640 0 3
rlabel polysilicon 1738 -634 1738 -634 0 1
rlabel polysilicon 1738 -640 1738 -640 0 3
rlabel polysilicon 1745 -634 1745 -634 0 1
rlabel polysilicon 1745 -640 1745 -640 0 3
rlabel polysilicon 1752 -634 1752 -634 0 1
rlabel polysilicon 1752 -640 1752 -640 0 3
rlabel polysilicon 1759 -634 1759 -634 0 1
rlabel polysilicon 1759 -640 1759 -640 0 3
rlabel polysilicon 1766 -634 1766 -634 0 1
rlabel polysilicon 1766 -640 1766 -640 0 3
rlabel polysilicon 1773 -634 1773 -634 0 1
rlabel polysilicon 1773 -640 1773 -640 0 3
rlabel polysilicon 1780 -634 1780 -634 0 1
rlabel polysilicon 1780 -640 1780 -640 0 3
rlabel polysilicon 1787 -634 1787 -634 0 1
rlabel polysilicon 1787 -640 1787 -640 0 3
rlabel polysilicon 1794 -634 1794 -634 0 1
rlabel polysilicon 1794 -640 1794 -640 0 3
rlabel polysilicon 1801 -634 1801 -634 0 1
rlabel polysilicon 1801 -640 1801 -640 0 3
rlabel polysilicon 1808 -634 1808 -634 0 1
rlabel polysilicon 1808 -640 1808 -640 0 3
rlabel polysilicon 1815 -634 1815 -634 0 1
rlabel polysilicon 1815 -640 1815 -640 0 3
rlabel polysilicon 1822 -634 1822 -634 0 1
rlabel polysilicon 1822 -640 1822 -640 0 3
rlabel polysilicon 1829 -634 1829 -634 0 1
rlabel polysilicon 1829 -640 1829 -640 0 3
rlabel polysilicon 1836 -634 1836 -634 0 1
rlabel polysilicon 1836 -640 1836 -640 0 3
rlabel polysilicon 1843 -634 1843 -634 0 1
rlabel polysilicon 1843 -640 1843 -640 0 3
rlabel polysilicon 1850 -634 1850 -634 0 1
rlabel polysilicon 1850 -640 1850 -640 0 3
rlabel polysilicon 1857 -634 1857 -634 0 1
rlabel polysilicon 1857 -640 1857 -640 0 3
rlabel polysilicon 1864 -634 1864 -634 0 1
rlabel polysilicon 1864 -640 1864 -640 0 3
rlabel polysilicon 1871 -634 1871 -634 0 1
rlabel polysilicon 1871 -640 1871 -640 0 3
rlabel polysilicon 1878 -634 1878 -634 0 1
rlabel polysilicon 1878 -640 1878 -640 0 3
rlabel polysilicon 1885 -634 1885 -634 0 1
rlabel polysilicon 1885 -640 1885 -640 0 3
rlabel polysilicon 1892 -634 1892 -634 0 1
rlabel polysilicon 1892 -640 1892 -640 0 3
rlabel polysilicon 1899 -634 1899 -634 0 1
rlabel polysilicon 1899 -640 1899 -640 0 3
rlabel polysilicon 1906 -634 1906 -634 0 1
rlabel polysilicon 1906 -640 1906 -640 0 3
rlabel polysilicon 1913 -634 1913 -634 0 1
rlabel polysilicon 1913 -640 1913 -640 0 3
rlabel polysilicon 1920 -634 1920 -634 0 1
rlabel polysilicon 1920 -640 1920 -640 0 3
rlabel polysilicon 1927 -634 1927 -634 0 1
rlabel polysilicon 1927 -640 1927 -640 0 3
rlabel polysilicon 1934 -634 1934 -634 0 1
rlabel polysilicon 1934 -640 1934 -640 0 3
rlabel polysilicon 1941 -634 1941 -634 0 1
rlabel polysilicon 1941 -640 1941 -640 0 3
rlabel polysilicon 1948 -634 1948 -634 0 1
rlabel polysilicon 1948 -640 1948 -640 0 3
rlabel polysilicon 1955 -634 1955 -634 0 1
rlabel polysilicon 1955 -640 1955 -640 0 3
rlabel polysilicon 1962 -634 1962 -634 0 1
rlabel polysilicon 1962 -640 1962 -640 0 3
rlabel polysilicon 1969 -634 1969 -634 0 1
rlabel polysilicon 1969 -640 1969 -640 0 3
rlabel polysilicon 1976 -634 1976 -634 0 1
rlabel polysilicon 1976 -640 1976 -640 0 3
rlabel polysilicon 1983 -634 1983 -634 0 1
rlabel polysilicon 1983 -640 1983 -640 0 3
rlabel polysilicon 1990 -634 1990 -634 0 1
rlabel polysilicon 1990 -640 1990 -640 0 3
rlabel polysilicon 1997 -634 1997 -634 0 1
rlabel polysilicon 1997 -640 1997 -640 0 3
rlabel polysilicon 2004 -634 2004 -634 0 1
rlabel polysilicon 2004 -640 2004 -640 0 3
rlabel polysilicon 2011 -634 2011 -634 0 1
rlabel polysilicon 2011 -640 2011 -640 0 3
rlabel polysilicon 2018 -634 2018 -634 0 1
rlabel polysilicon 2018 -640 2018 -640 0 3
rlabel polysilicon 2025 -634 2025 -634 0 1
rlabel polysilicon 2025 -640 2025 -640 0 3
rlabel polysilicon 2032 -634 2032 -634 0 1
rlabel polysilicon 2032 -640 2032 -640 0 3
rlabel polysilicon 2039 -634 2039 -634 0 1
rlabel polysilicon 2039 -640 2039 -640 0 3
rlabel polysilicon 2046 -634 2046 -634 0 1
rlabel polysilicon 2046 -640 2046 -640 0 3
rlabel polysilicon 2053 -634 2053 -634 0 1
rlabel polysilicon 2053 -640 2053 -640 0 3
rlabel polysilicon 2060 -634 2060 -634 0 1
rlabel polysilicon 2060 -640 2060 -640 0 3
rlabel polysilicon 2067 -634 2067 -634 0 1
rlabel polysilicon 2067 -640 2067 -640 0 3
rlabel polysilicon 2074 -634 2074 -634 0 1
rlabel polysilicon 2074 -640 2074 -640 0 3
rlabel polysilicon 2081 -634 2081 -634 0 1
rlabel polysilicon 2081 -640 2081 -640 0 3
rlabel polysilicon 2088 -634 2088 -634 0 1
rlabel polysilicon 2088 -640 2088 -640 0 3
rlabel polysilicon 2095 -634 2095 -634 0 1
rlabel polysilicon 2095 -640 2095 -640 0 3
rlabel polysilicon 2102 -634 2102 -634 0 1
rlabel polysilicon 2102 -640 2102 -640 0 3
rlabel polysilicon 2109 -634 2109 -634 0 1
rlabel polysilicon 2109 -640 2109 -640 0 3
rlabel polysilicon 2116 -634 2116 -634 0 1
rlabel polysilicon 2116 -640 2116 -640 0 3
rlabel polysilicon 2123 -634 2123 -634 0 1
rlabel polysilicon 2123 -640 2123 -640 0 3
rlabel polysilicon 2130 -634 2130 -634 0 1
rlabel polysilicon 2130 -640 2130 -640 0 3
rlabel polysilicon 2137 -634 2137 -634 0 1
rlabel polysilicon 2137 -640 2137 -640 0 3
rlabel polysilicon 2144 -634 2144 -634 0 1
rlabel polysilicon 2144 -640 2144 -640 0 3
rlabel polysilicon 2151 -634 2151 -634 0 1
rlabel polysilicon 2151 -640 2151 -640 0 3
rlabel polysilicon 2158 -634 2158 -634 0 1
rlabel polysilicon 2158 -640 2158 -640 0 3
rlabel polysilicon 2165 -634 2165 -634 0 1
rlabel polysilicon 2165 -640 2165 -640 0 3
rlabel polysilicon 2172 -634 2172 -634 0 1
rlabel polysilicon 2172 -640 2172 -640 0 3
rlabel polysilicon 2179 -634 2179 -634 0 1
rlabel polysilicon 2179 -640 2179 -640 0 3
rlabel polysilicon 2186 -634 2186 -634 0 1
rlabel polysilicon 2186 -640 2186 -640 0 3
rlabel polysilicon 2193 -634 2193 -634 0 1
rlabel polysilicon 2193 -640 2193 -640 0 3
rlabel polysilicon 2200 -634 2200 -634 0 1
rlabel polysilicon 2200 -640 2200 -640 0 3
rlabel polysilicon 2207 -634 2207 -634 0 1
rlabel polysilicon 2210 -634 2210 -634 0 2
rlabel polysilicon 2207 -640 2207 -640 0 3
rlabel polysilicon 2214 -634 2214 -634 0 1
rlabel polysilicon 2214 -640 2214 -640 0 3
rlabel polysilicon 2217 -640 2217 -640 0 4
rlabel polysilicon 2221 -634 2221 -634 0 1
rlabel polysilicon 2224 -634 2224 -634 0 2
rlabel polysilicon 2224 -640 2224 -640 0 4
rlabel polysilicon 2291 -634 2291 -634 0 1
rlabel polysilicon 2291 -640 2291 -640 0 3
rlabel polysilicon 2326 -634 2326 -634 0 1
rlabel polysilicon 2326 -640 2326 -640 0 3
rlabel polysilicon 2361 -634 2361 -634 0 1
rlabel polysilicon 2361 -640 2361 -640 0 3
rlabel polysilicon 2 -811 2 -811 0 1
rlabel polysilicon 2 -817 2 -817 0 3
rlabel polysilicon 12 -811 12 -811 0 2
rlabel polysilicon 9 -817 9 -817 0 3
rlabel polysilicon 19 -811 19 -811 0 2
rlabel polysilicon 16 -817 16 -817 0 3
rlabel polysilicon 19 -817 19 -817 0 4
rlabel polysilicon 23 -811 23 -811 0 1
rlabel polysilicon 23 -817 23 -817 0 3
rlabel polysilicon 30 -811 30 -811 0 1
rlabel polysilicon 30 -817 30 -817 0 3
rlabel polysilicon 37 -811 37 -811 0 1
rlabel polysilicon 37 -817 37 -817 0 3
rlabel polysilicon 44 -811 44 -811 0 1
rlabel polysilicon 47 -811 47 -811 0 2
rlabel polysilicon 44 -817 44 -817 0 3
rlabel polysilicon 47 -817 47 -817 0 4
rlabel polysilicon 51 -811 51 -811 0 1
rlabel polysilicon 51 -817 51 -817 0 3
rlabel polysilicon 58 -811 58 -811 0 1
rlabel polysilicon 58 -817 58 -817 0 3
rlabel polysilicon 65 -811 65 -811 0 1
rlabel polysilicon 68 -811 68 -811 0 2
rlabel polysilicon 65 -817 65 -817 0 3
rlabel polysilicon 72 -811 72 -811 0 1
rlabel polysilicon 72 -817 72 -817 0 3
rlabel polysilicon 79 -811 79 -811 0 1
rlabel polysilicon 82 -811 82 -811 0 2
rlabel polysilicon 79 -817 79 -817 0 3
rlabel polysilicon 86 -811 86 -811 0 1
rlabel polysilicon 86 -817 86 -817 0 3
rlabel polysilicon 93 -811 93 -811 0 1
rlabel polysilicon 93 -817 93 -817 0 3
rlabel polysilicon 100 -811 100 -811 0 1
rlabel polysilicon 100 -817 100 -817 0 3
rlabel polysilicon 107 -811 107 -811 0 1
rlabel polysilicon 107 -817 107 -817 0 3
rlabel polysilicon 114 -811 114 -811 0 1
rlabel polysilicon 114 -817 114 -817 0 3
rlabel polysilicon 121 -817 121 -817 0 3
rlabel polysilicon 124 -817 124 -817 0 4
rlabel polysilicon 128 -811 128 -811 0 1
rlabel polysilicon 131 -811 131 -811 0 2
rlabel polysilicon 128 -817 128 -817 0 3
rlabel polysilicon 135 -811 135 -811 0 1
rlabel polysilicon 135 -817 135 -817 0 3
rlabel polysilicon 142 -811 142 -811 0 1
rlabel polysilicon 145 -811 145 -811 0 2
rlabel polysilicon 145 -817 145 -817 0 4
rlabel polysilicon 149 -811 149 -811 0 1
rlabel polysilicon 149 -817 149 -817 0 3
rlabel polysilicon 156 -811 156 -811 0 1
rlabel polysilicon 156 -817 156 -817 0 3
rlabel polysilicon 163 -811 163 -811 0 1
rlabel polysilicon 163 -817 163 -817 0 3
rlabel polysilicon 170 -811 170 -811 0 1
rlabel polysilicon 170 -817 170 -817 0 3
rlabel polysilicon 177 -811 177 -811 0 1
rlabel polysilicon 177 -817 177 -817 0 3
rlabel polysilicon 184 -811 184 -811 0 1
rlabel polysilicon 187 -811 187 -811 0 2
rlabel polysilicon 184 -817 184 -817 0 3
rlabel polysilicon 187 -817 187 -817 0 4
rlabel polysilicon 191 -811 191 -811 0 1
rlabel polysilicon 191 -817 191 -817 0 3
rlabel polysilicon 198 -811 198 -811 0 1
rlabel polysilicon 198 -817 198 -817 0 3
rlabel polysilicon 205 -811 205 -811 0 1
rlabel polysilicon 208 -811 208 -811 0 2
rlabel polysilicon 205 -817 205 -817 0 3
rlabel polysilicon 212 -811 212 -811 0 1
rlabel polysilicon 212 -817 212 -817 0 3
rlabel polysilicon 219 -811 219 -811 0 1
rlabel polysilicon 222 -811 222 -811 0 2
rlabel polysilicon 222 -817 222 -817 0 4
rlabel polysilicon 226 -811 226 -811 0 1
rlabel polysilicon 226 -817 226 -817 0 3
rlabel polysilicon 233 -811 233 -811 0 1
rlabel polysilicon 236 -811 236 -811 0 2
rlabel polysilicon 233 -817 233 -817 0 3
rlabel polysilicon 240 -811 240 -811 0 1
rlabel polysilicon 240 -817 240 -817 0 3
rlabel polysilicon 247 -811 247 -811 0 1
rlabel polysilicon 247 -817 247 -817 0 3
rlabel polysilicon 254 -811 254 -811 0 1
rlabel polysilicon 254 -817 254 -817 0 3
rlabel polysilicon 261 -811 261 -811 0 1
rlabel polysilicon 261 -817 261 -817 0 3
rlabel polysilicon 268 -811 268 -811 0 1
rlabel polysilicon 268 -817 268 -817 0 3
rlabel polysilicon 275 -811 275 -811 0 1
rlabel polysilicon 275 -817 275 -817 0 3
rlabel polysilicon 282 -811 282 -811 0 1
rlabel polysilicon 282 -817 282 -817 0 3
rlabel polysilicon 289 -811 289 -811 0 1
rlabel polysilicon 289 -817 289 -817 0 3
rlabel polysilicon 296 -811 296 -811 0 1
rlabel polysilicon 296 -817 296 -817 0 3
rlabel polysilicon 303 -811 303 -811 0 1
rlabel polysilicon 303 -817 303 -817 0 3
rlabel polysilicon 310 -811 310 -811 0 1
rlabel polysilicon 310 -817 310 -817 0 3
rlabel polysilicon 317 -811 317 -811 0 1
rlabel polysilicon 317 -817 317 -817 0 3
rlabel polysilicon 324 -811 324 -811 0 1
rlabel polysilicon 324 -817 324 -817 0 3
rlabel polysilicon 331 -811 331 -811 0 1
rlabel polysilicon 331 -817 331 -817 0 3
rlabel polysilicon 338 -811 338 -811 0 1
rlabel polysilicon 338 -817 338 -817 0 3
rlabel polysilicon 345 -811 345 -811 0 1
rlabel polysilicon 345 -817 345 -817 0 3
rlabel polysilicon 352 -811 352 -811 0 1
rlabel polysilicon 352 -817 352 -817 0 3
rlabel polysilicon 359 -811 359 -811 0 1
rlabel polysilicon 362 -811 362 -811 0 2
rlabel polysilicon 359 -817 359 -817 0 3
rlabel polysilicon 362 -817 362 -817 0 4
rlabel polysilicon 366 -811 366 -811 0 1
rlabel polysilicon 366 -817 366 -817 0 3
rlabel polysilicon 373 -811 373 -811 0 1
rlabel polysilicon 373 -817 373 -817 0 3
rlabel polysilicon 380 -811 380 -811 0 1
rlabel polysilicon 380 -817 380 -817 0 3
rlabel polysilicon 387 -811 387 -811 0 1
rlabel polysilicon 387 -817 387 -817 0 3
rlabel polysilicon 394 -811 394 -811 0 1
rlabel polysilicon 394 -817 394 -817 0 3
rlabel polysilicon 401 -811 401 -811 0 1
rlabel polysilicon 401 -817 401 -817 0 3
rlabel polysilicon 408 -811 408 -811 0 1
rlabel polysilicon 408 -817 408 -817 0 3
rlabel polysilicon 415 -811 415 -811 0 1
rlabel polysilicon 415 -817 415 -817 0 3
rlabel polysilicon 422 -811 422 -811 0 1
rlabel polysilicon 422 -817 422 -817 0 3
rlabel polysilicon 429 -811 429 -811 0 1
rlabel polysilicon 429 -817 429 -817 0 3
rlabel polysilicon 436 -811 436 -811 0 1
rlabel polysilicon 436 -817 436 -817 0 3
rlabel polysilicon 443 -811 443 -811 0 1
rlabel polysilicon 443 -817 443 -817 0 3
rlabel polysilicon 450 -811 450 -811 0 1
rlabel polysilicon 450 -817 450 -817 0 3
rlabel polysilicon 457 -811 457 -811 0 1
rlabel polysilicon 457 -817 457 -817 0 3
rlabel polysilicon 464 -811 464 -811 0 1
rlabel polysilicon 464 -817 464 -817 0 3
rlabel polysilicon 471 -811 471 -811 0 1
rlabel polysilicon 471 -817 471 -817 0 3
rlabel polysilicon 478 -811 478 -811 0 1
rlabel polysilicon 478 -817 478 -817 0 3
rlabel polysilicon 485 -811 485 -811 0 1
rlabel polysilicon 485 -817 485 -817 0 3
rlabel polysilicon 492 -811 492 -811 0 1
rlabel polysilicon 492 -817 492 -817 0 3
rlabel polysilicon 499 -811 499 -811 0 1
rlabel polysilicon 499 -817 499 -817 0 3
rlabel polysilicon 506 -811 506 -811 0 1
rlabel polysilicon 506 -817 506 -817 0 3
rlabel polysilicon 513 -811 513 -811 0 1
rlabel polysilicon 513 -817 513 -817 0 3
rlabel polysilicon 520 -811 520 -811 0 1
rlabel polysilicon 523 -811 523 -811 0 2
rlabel polysilicon 520 -817 520 -817 0 3
rlabel polysilicon 527 -811 527 -811 0 1
rlabel polysilicon 527 -817 527 -817 0 3
rlabel polysilicon 534 -811 534 -811 0 1
rlabel polysilicon 534 -817 534 -817 0 3
rlabel polysilicon 541 -811 541 -811 0 1
rlabel polysilicon 541 -817 541 -817 0 3
rlabel polysilicon 548 -811 548 -811 0 1
rlabel polysilicon 548 -817 548 -817 0 3
rlabel polysilicon 555 -811 555 -811 0 1
rlabel polysilicon 555 -817 555 -817 0 3
rlabel polysilicon 562 -811 562 -811 0 1
rlabel polysilicon 562 -817 562 -817 0 3
rlabel polysilicon 569 -811 569 -811 0 1
rlabel polysilicon 569 -817 569 -817 0 3
rlabel polysilicon 576 -811 576 -811 0 1
rlabel polysilicon 576 -817 576 -817 0 3
rlabel polysilicon 583 -811 583 -811 0 1
rlabel polysilicon 586 -811 586 -811 0 2
rlabel polysilicon 583 -817 583 -817 0 3
rlabel polysilicon 586 -817 586 -817 0 4
rlabel polysilicon 590 -811 590 -811 0 1
rlabel polysilicon 590 -817 590 -817 0 3
rlabel polysilicon 593 -817 593 -817 0 4
rlabel polysilicon 597 -811 597 -811 0 1
rlabel polysilicon 597 -817 597 -817 0 3
rlabel polysilicon 604 -811 604 -811 0 1
rlabel polysilicon 604 -817 604 -817 0 3
rlabel polysilicon 611 -811 611 -811 0 1
rlabel polysilicon 611 -817 611 -817 0 3
rlabel polysilicon 618 -811 618 -811 0 1
rlabel polysilicon 618 -817 618 -817 0 3
rlabel polysilicon 625 -811 625 -811 0 1
rlabel polysilicon 625 -817 625 -817 0 3
rlabel polysilicon 632 -811 632 -811 0 1
rlabel polysilicon 632 -817 632 -817 0 3
rlabel polysilicon 639 -811 639 -811 0 1
rlabel polysilicon 639 -817 639 -817 0 3
rlabel polysilicon 646 -811 646 -811 0 1
rlabel polysilicon 646 -817 646 -817 0 3
rlabel polysilicon 653 -811 653 -811 0 1
rlabel polysilicon 653 -817 653 -817 0 3
rlabel polysilicon 660 -811 660 -811 0 1
rlabel polysilicon 660 -817 660 -817 0 3
rlabel polysilicon 667 -811 667 -811 0 1
rlabel polysilicon 667 -817 667 -817 0 3
rlabel polysilicon 674 -811 674 -811 0 1
rlabel polysilicon 674 -817 674 -817 0 3
rlabel polysilicon 681 -811 681 -811 0 1
rlabel polysilicon 684 -811 684 -811 0 2
rlabel polysilicon 684 -817 684 -817 0 4
rlabel polysilicon 688 -811 688 -811 0 1
rlabel polysilicon 688 -817 688 -817 0 3
rlabel polysilicon 698 -811 698 -811 0 2
rlabel polysilicon 695 -817 695 -817 0 3
rlabel polysilicon 698 -817 698 -817 0 4
rlabel polysilicon 702 -811 702 -811 0 1
rlabel polysilicon 702 -817 702 -817 0 3
rlabel polysilicon 709 -811 709 -811 0 1
rlabel polysilicon 709 -817 709 -817 0 3
rlabel polysilicon 716 -811 716 -811 0 1
rlabel polysilicon 716 -817 716 -817 0 3
rlabel polysilicon 726 -811 726 -811 0 2
rlabel polysilicon 723 -817 723 -817 0 3
rlabel polysilicon 726 -817 726 -817 0 4
rlabel polysilicon 730 -811 730 -811 0 1
rlabel polysilicon 730 -817 730 -817 0 3
rlabel polysilicon 737 -811 737 -811 0 1
rlabel polysilicon 737 -817 737 -817 0 3
rlabel polysilicon 744 -811 744 -811 0 1
rlabel polysilicon 747 -811 747 -811 0 2
rlabel polysilicon 744 -817 744 -817 0 3
rlabel polysilicon 747 -817 747 -817 0 4
rlabel polysilicon 751 -811 751 -811 0 1
rlabel polysilicon 754 -811 754 -811 0 2
rlabel polysilicon 751 -817 751 -817 0 3
rlabel polysilicon 754 -817 754 -817 0 4
rlabel polysilicon 758 -811 758 -811 0 1
rlabel polysilicon 758 -817 758 -817 0 3
rlabel polysilicon 765 -811 765 -811 0 1
rlabel polysilicon 765 -817 765 -817 0 3
rlabel polysilicon 772 -811 772 -811 0 1
rlabel polysilicon 772 -817 772 -817 0 3
rlabel polysilicon 779 -811 779 -811 0 1
rlabel polysilicon 779 -817 779 -817 0 3
rlabel polysilicon 786 -811 786 -811 0 1
rlabel polysilicon 786 -817 786 -817 0 3
rlabel polysilicon 793 -811 793 -811 0 1
rlabel polysilicon 793 -817 793 -817 0 3
rlabel polysilicon 800 -811 800 -811 0 1
rlabel polysilicon 800 -817 800 -817 0 3
rlabel polysilicon 807 -811 807 -811 0 1
rlabel polysilicon 807 -817 807 -817 0 3
rlabel polysilicon 814 -811 814 -811 0 1
rlabel polysilicon 814 -817 814 -817 0 3
rlabel polysilicon 821 -811 821 -811 0 1
rlabel polysilicon 821 -817 821 -817 0 3
rlabel polysilicon 828 -811 828 -811 0 1
rlabel polysilicon 828 -817 828 -817 0 3
rlabel polysilicon 831 -817 831 -817 0 4
rlabel polysilicon 835 -811 835 -811 0 1
rlabel polysilicon 835 -817 835 -817 0 3
rlabel polysilicon 842 -811 842 -811 0 1
rlabel polysilicon 842 -817 842 -817 0 3
rlabel polysilicon 849 -811 849 -811 0 1
rlabel polysilicon 849 -817 849 -817 0 3
rlabel polysilicon 856 -811 856 -811 0 1
rlabel polysilicon 856 -817 856 -817 0 3
rlabel polysilicon 863 -811 863 -811 0 1
rlabel polysilicon 863 -817 863 -817 0 3
rlabel polysilicon 870 -811 870 -811 0 1
rlabel polysilicon 870 -817 870 -817 0 3
rlabel polysilicon 880 -811 880 -811 0 2
rlabel polysilicon 877 -817 877 -817 0 3
rlabel polysilicon 884 -811 884 -811 0 1
rlabel polysilicon 884 -817 884 -817 0 3
rlabel polysilicon 891 -811 891 -811 0 1
rlabel polysilicon 891 -817 891 -817 0 3
rlabel polysilicon 898 -811 898 -811 0 1
rlabel polysilicon 898 -817 898 -817 0 3
rlabel polysilicon 905 -811 905 -811 0 1
rlabel polysilicon 905 -817 905 -817 0 3
rlabel polysilicon 912 -811 912 -811 0 1
rlabel polysilicon 912 -817 912 -817 0 3
rlabel polysilicon 919 -811 919 -811 0 1
rlabel polysilicon 919 -817 919 -817 0 3
rlabel polysilicon 926 -811 926 -811 0 1
rlabel polysilicon 926 -817 926 -817 0 3
rlabel polysilicon 933 -811 933 -811 0 1
rlabel polysilicon 933 -817 933 -817 0 3
rlabel polysilicon 940 -811 940 -811 0 1
rlabel polysilicon 940 -817 940 -817 0 3
rlabel polysilicon 947 -811 947 -811 0 1
rlabel polysilicon 947 -817 947 -817 0 3
rlabel polysilicon 954 -811 954 -811 0 1
rlabel polysilicon 957 -811 957 -811 0 2
rlabel polysilicon 954 -817 954 -817 0 3
rlabel polysilicon 957 -817 957 -817 0 4
rlabel polysilicon 961 -811 961 -811 0 1
rlabel polysilicon 961 -817 961 -817 0 3
rlabel polysilicon 968 -811 968 -811 0 1
rlabel polysilicon 968 -817 968 -817 0 3
rlabel polysilicon 975 -811 975 -811 0 1
rlabel polysilicon 975 -817 975 -817 0 3
rlabel polysilicon 982 -811 982 -811 0 1
rlabel polysilicon 982 -817 982 -817 0 3
rlabel polysilicon 989 -811 989 -811 0 1
rlabel polysilicon 989 -817 989 -817 0 3
rlabel polysilicon 996 -811 996 -811 0 1
rlabel polysilicon 996 -817 996 -817 0 3
rlabel polysilicon 1003 -811 1003 -811 0 1
rlabel polysilicon 1003 -817 1003 -817 0 3
rlabel polysilicon 1010 -811 1010 -811 0 1
rlabel polysilicon 1010 -817 1010 -817 0 3
rlabel polysilicon 1013 -817 1013 -817 0 4
rlabel polysilicon 1017 -811 1017 -811 0 1
rlabel polysilicon 1017 -817 1017 -817 0 3
rlabel polysilicon 1024 -811 1024 -811 0 1
rlabel polysilicon 1024 -817 1024 -817 0 3
rlabel polysilicon 1031 -811 1031 -811 0 1
rlabel polysilicon 1031 -817 1031 -817 0 3
rlabel polysilicon 1038 -811 1038 -811 0 1
rlabel polysilicon 1038 -817 1038 -817 0 3
rlabel polysilicon 1045 -811 1045 -811 0 1
rlabel polysilicon 1045 -817 1045 -817 0 3
rlabel polysilicon 1052 -811 1052 -811 0 1
rlabel polysilicon 1052 -817 1052 -817 0 3
rlabel polysilicon 1059 -811 1059 -811 0 1
rlabel polysilicon 1059 -817 1059 -817 0 3
rlabel polysilicon 1066 -811 1066 -811 0 1
rlabel polysilicon 1066 -817 1066 -817 0 3
rlabel polysilicon 1073 -811 1073 -811 0 1
rlabel polysilicon 1073 -817 1073 -817 0 3
rlabel polysilicon 1080 -811 1080 -811 0 1
rlabel polysilicon 1080 -817 1080 -817 0 3
rlabel polysilicon 1087 -811 1087 -811 0 1
rlabel polysilicon 1087 -817 1087 -817 0 3
rlabel polysilicon 1094 -811 1094 -811 0 1
rlabel polysilicon 1094 -817 1094 -817 0 3
rlabel polysilicon 1101 -811 1101 -811 0 1
rlabel polysilicon 1101 -817 1101 -817 0 3
rlabel polysilicon 1108 -811 1108 -811 0 1
rlabel polysilicon 1111 -811 1111 -811 0 2
rlabel polysilicon 1108 -817 1108 -817 0 3
rlabel polysilicon 1111 -817 1111 -817 0 4
rlabel polysilicon 1115 -811 1115 -811 0 1
rlabel polysilicon 1115 -817 1115 -817 0 3
rlabel polysilicon 1122 -811 1122 -811 0 1
rlabel polysilicon 1122 -817 1122 -817 0 3
rlabel polysilicon 1129 -811 1129 -811 0 1
rlabel polysilicon 1129 -817 1129 -817 0 3
rlabel polysilicon 1132 -817 1132 -817 0 4
rlabel polysilicon 1136 -811 1136 -811 0 1
rlabel polysilicon 1139 -811 1139 -811 0 2
rlabel polysilicon 1136 -817 1136 -817 0 3
rlabel polysilicon 1139 -817 1139 -817 0 4
rlabel polysilicon 1143 -811 1143 -811 0 1
rlabel polysilicon 1146 -811 1146 -811 0 2
rlabel polysilicon 1143 -817 1143 -817 0 3
rlabel polysilicon 1146 -817 1146 -817 0 4
rlabel polysilicon 1150 -811 1150 -811 0 1
rlabel polysilicon 1150 -817 1150 -817 0 3
rlabel polysilicon 1157 -811 1157 -811 0 1
rlabel polysilicon 1157 -817 1157 -817 0 3
rlabel polysilicon 1160 -817 1160 -817 0 4
rlabel polysilicon 1164 -811 1164 -811 0 1
rlabel polysilicon 1164 -817 1164 -817 0 3
rlabel polysilicon 1171 -811 1171 -811 0 1
rlabel polysilicon 1174 -811 1174 -811 0 2
rlabel polysilicon 1171 -817 1171 -817 0 3
rlabel polysilicon 1174 -817 1174 -817 0 4
rlabel polysilicon 1178 -811 1178 -811 0 1
rlabel polysilicon 1178 -817 1178 -817 0 3
rlabel polysilicon 1185 -811 1185 -811 0 1
rlabel polysilicon 1185 -817 1185 -817 0 3
rlabel polysilicon 1192 -811 1192 -811 0 1
rlabel polysilicon 1192 -817 1192 -817 0 3
rlabel polysilicon 1199 -811 1199 -811 0 1
rlabel polysilicon 1199 -817 1199 -817 0 3
rlabel polysilicon 1206 -811 1206 -811 0 1
rlabel polysilicon 1209 -811 1209 -811 0 2
rlabel polysilicon 1206 -817 1206 -817 0 3
rlabel polysilicon 1209 -817 1209 -817 0 4
rlabel polysilicon 1213 -811 1213 -811 0 1
rlabel polysilicon 1213 -817 1213 -817 0 3
rlabel polysilicon 1216 -817 1216 -817 0 4
rlabel polysilicon 1220 -811 1220 -811 0 1
rlabel polysilicon 1223 -811 1223 -811 0 2
rlabel polysilicon 1220 -817 1220 -817 0 3
rlabel polysilicon 1223 -817 1223 -817 0 4
rlabel polysilicon 1227 -811 1227 -811 0 1
rlabel polysilicon 1227 -817 1227 -817 0 3
rlabel polysilicon 1234 -811 1234 -811 0 1
rlabel polysilicon 1234 -817 1234 -817 0 3
rlabel polysilicon 1241 -811 1241 -811 0 1
rlabel polysilicon 1241 -817 1241 -817 0 3
rlabel polysilicon 1248 -811 1248 -811 0 1
rlabel polysilicon 1248 -817 1248 -817 0 3
rlabel polysilicon 1255 -811 1255 -811 0 1
rlabel polysilicon 1255 -817 1255 -817 0 3
rlabel polysilicon 1262 -811 1262 -811 0 1
rlabel polysilicon 1262 -817 1262 -817 0 3
rlabel polysilicon 1269 -811 1269 -811 0 1
rlabel polysilicon 1269 -817 1269 -817 0 3
rlabel polysilicon 1276 -811 1276 -811 0 1
rlabel polysilicon 1276 -817 1276 -817 0 3
rlabel polysilicon 1283 -811 1283 -811 0 1
rlabel polysilicon 1283 -817 1283 -817 0 3
rlabel polysilicon 1290 -811 1290 -811 0 1
rlabel polysilicon 1290 -817 1290 -817 0 3
rlabel polysilicon 1297 -811 1297 -811 0 1
rlabel polysilicon 1297 -817 1297 -817 0 3
rlabel polysilicon 1304 -811 1304 -811 0 1
rlabel polysilicon 1304 -817 1304 -817 0 3
rlabel polysilicon 1311 -811 1311 -811 0 1
rlabel polysilicon 1311 -817 1311 -817 0 3
rlabel polysilicon 1318 -811 1318 -811 0 1
rlabel polysilicon 1318 -817 1318 -817 0 3
rlabel polysilicon 1325 -811 1325 -811 0 1
rlabel polysilicon 1325 -817 1325 -817 0 3
rlabel polysilicon 1332 -811 1332 -811 0 1
rlabel polysilicon 1335 -817 1335 -817 0 4
rlabel polysilicon 1339 -811 1339 -811 0 1
rlabel polysilicon 1339 -817 1339 -817 0 3
rlabel polysilicon 1346 -811 1346 -811 0 1
rlabel polysilicon 1346 -817 1346 -817 0 3
rlabel polysilicon 1353 -811 1353 -811 0 1
rlabel polysilicon 1353 -817 1353 -817 0 3
rlabel polysilicon 1360 -811 1360 -811 0 1
rlabel polysilicon 1360 -817 1360 -817 0 3
rlabel polysilicon 1363 -817 1363 -817 0 4
rlabel polysilicon 1370 -811 1370 -811 0 2
rlabel polysilicon 1367 -817 1367 -817 0 3
rlabel polysilicon 1370 -817 1370 -817 0 4
rlabel polysilicon 1374 -811 1374 -811 0 1
rlabel polysilicon 1374 -817 1374 -817 0 3
rlabel polysilicon 1381 -811 1381 -811 0 1
rlabel polysilicon 1381 -817 1381 -817 0 3
rlabel polysilicon 1388 -811 1388 -811 0 1
rlabel polysilicon 1388 -817 1388 -817 0 3
rlabel polysilicon 1395 -811 1395 -811 0 1
rlabel polysilicon 1395 -817 1395 -817 0 3
rlabel polysilicon 1402 -811 1402 -811 0 1
rlabel polysilicon 1402 -817 1402 -817 0 3
rlabel polysilicon 1409 -811 1409 -811 0 1
rlabel polysilicon 1409 -817 1409 -817 0 3
rlabel polysilicon 1416 -811 1416 -811 0 1
rlabel polysilicon 1416 -817 1416 -817 0 3
rlabel polysilicon 1423 -811 1423 -811 0 1
rlabel polysilicon 1423 -817 1423 -817 0 3
rlabel polysilicon 1430 -811 1430 -811 0 1
rlabel polysilicon 1430 -817 1430 -817 0 3
rlabel polysilicon 1437 -811 1437 -811 0 1
rlabel polysilicon 1437 -817 1437 -817 0 3
rlabel polysilicon 1444 -811 1444 -811 0 1
rlabel polysilicon 1444 -817 1444 -817 0 3
rlabel polysilicon 1451 -811 1451 -811 0 1
rlabel polysilicon 1451 -817 1451 -817 0 3
rlabel polysilicon 1458 -811 1458 -811 0 1
rlabel polysilicon 1458 -817 1458 -817 0 3
rlabel polysilicon 1465 -811 1465 -811 0 1
rlabel polysilicon 1465 -817 1465 -817 0 3
rlabel polysilicon 1472 -811 1472 -811 0 1
rlabel polysilicon 1472 -817 1472 -817 0 3
rlabel polysilicon 1479 -811 1479 -811 0 1
rlabel polysilicon 1479 -817 1479 -817 0 3
rlabel polysilicon 1486 -811 1486 -811 0 1
rlabel polysilicon 1486 -817 1486 -817 0 3
rlabel polysilicon 1493 -811 1493 -811 0 1
rlabel polysilicon 1493 -817 1493 -817 0 3
rlabel polysilicon 1500 -811 1500 -811 0 1
rlabel polysilicon 1500 -817 1500 -817 0 3
rlabel polysilicon 1507 -811 1507 -811 0 1
rlabel polysilicon 1507 -817 1507 -817 0 3
rlabel polysilicon 1514 -811 1514 -811 0 1
rlabel polysilicon 1514 -817 1514 -817 0 3
rlabel polysilicon 1521 -811 1521 -811 0 1
rlabel polysilicon 1521 -817 1521 -817 0 3
rlabel polysilicon 1528 -811 1528 -811 0 1
rlabel polysilicon 1528 -817 1528 -817 0 3
rlabel polysilicon 1535 -811 1535 -811 0 1
rlabel polysilicon 1538 -811 1538 -811 0 2
rlabel polysilicon 1535 -817 1535 -817 0 3
rlabel polysilicon 1538 -817 1538 -817 0 4
rlabel polysilicon 1542 -811 1542 -811 0 1
rlabel polysilicon 1542 -817 1542 -817 0 3
rlabel polysilicon 1549 -811 1549 -811 0 1
rlabel polysilicon 1549 -817 1549 -817 0 3
rlabel polysilicon 1556 -811 1556 -811 0 1
rlabel polysilicon 1556 -817 1556 -817 0 3
rlabel polysilicon 1563 -811 1563 -811 0 1
rlabel polysilicon 1563 -817 1563 -817 0 3
rlabel polysilicon 1570 -811 1570 -811 0 1
rlabel polysilicon 1570 -817 1570 -817 0 3
rlabel polysilicon 1577 -811 1577 -811 0 1
rlabel polysilicon 1577 -817 1577 -817 0 3
rlabel polysilicon 1584 -811 1584 -811 0 1
rlabel polysilicon 1584 -817 1584 -817 0 3
rlabel polysilicon 1591 -811 1591 -811 0 1
rlabel polysilicon 1591 -817 1591 -817 0 3
rlabel polysilicon 1598 -811 1598 -811 0 1
rlabel polysilicon 1598 -817 1598 -817 0 3
rlabel polysilicon 1605 -811 1605 -811 0 1
rlabel polysilicon 1605 -817 1605 -817 0 3
rlabel polysilicon 1612 -811 1612 -811 0 1
rlabel polysilicon 1612 -817 1612 -817 0 3
rlabel polysilicon 1619 -811 1619 -811 0 1
rlabel polysilicon 1619 -817 1619 -817 0 3
rlabel polysilicon 1626 -811 1626 -811 0 1
rlabel polysilicon 1626 -817 1626 -817 0 3
rlabel polysilicon 1633 -811 1633 -811 0 1
rlabel polysilicon 1633 -817 1633 -817 0 3
rlabel polysilicon 1640 -811 1640 -811 0 1
rlabel polysilicon 1640 -817 1640 -817 0 3
rlabel polysilicon 1647 -811 1647 -811 0 1
rlabel polysilicon 1647 -817 1647 -817 0 3
rlabel polysilicon 1654 -811 1654 -811 0 1
rlabel polysilicon 1654 -817 1654 -817 0 3
rlabel polysilicon 1661 -811 1661 -811 0 1
rlabel polysilicon 1661 -817 1661 -817 0 3
rlabel polysilicon 1668 -811 1668 -811 0 1
rlabel polysilicon 1668 -817 1668 -817 0 3
rlabel polysilicon 1675 -811 1675 -811 0 1
rlabel polysilicon 1675 -817 1675 -817 0 3
rlabel polysilicon 1682 -811 1682 -811 0 1
rlabel polysilicon 1682 -817 1682 -817 0 3
rlabel polysilicon 1689 -811 1689 -811 0 1
rlabel polysilicon 1689 -817 1689 -817 0 3
rlabel polysilicon 1696 -811 1696 -811 0 1
rlabel polysilicon 1696 -817 1696 -817 0 3
rlabel polysilicon 1703 -811 1703 -811 0 1
rlabel polysilicon 1703 -817 1703 -817 0 3
rlabel polysilicon 1710 -811 1710 -811 0 1
rlabel polysilicon 1710 -817 1710 -817 0 3
rlabel polysilicon 1717 -811 1717 -811 0 1
rlabel polysilicon 1717 -817 1717 -817 0 3
rlabel polysilicon 1724 -811 1724 -811 0 1
rlabel polysilicon 1724 -817 1724 -817 0 3
rlabel polysilicon 1731 -811 1731 -811 0 1
rlabel polysilicon 1731 -817 1731 -817 0 3
rlabel polysilicon 1738 -811 1738 -811 0 1
rlabel polysilicon 1738 -817 1738 -817 0 3
rlabel polysilicon 1745 -811 1745 -811 0 1
rlabel polysilicon 1745 -817 1745 -817 0 3
rlabel polysilicon 1752 -811 1752 -811 0 1
rlabel polysilicon 1752 -817 1752 -817 0 3
rlabel polysilicon 1759 -811 1759 -811 0 1
rlabel polysilicon 1759 -817 1759 -817 0 3
rlabel polysilicon 1766 -811 1766 -811 0 1
rlabel polysilicon 1766 -817 1766 -817 0 3
rlabel polysilicon 1773 -811 1773 -811 0 1
rlabel polysilicon 1773 -817 1773 -817 0 3
rlabel polysilicon 1780 -811 1780 -811 0 1
rlabel polysilicon 1780 -817 1780 -817 0 3
rlabel polysilicon 1787 -811 1787 -811 0 1
rlabel polysilicon 1787 -817 1787 -817 0 3
rlabel polysilicon 1794 -811 1794 -811 0 1
rlabel polysilicon 1794 -817 1794 -817 0 3
rlabel polysilicon 1801 -811 1801 -811 0 1
rlabel polysilicon 1801 -817 1801 -817 0 3
rlabel polysilicon 1808 -811 1808 -811 0 1
rlabel polysilicon 1808 -817 1808 -817 0 3
rlabel polysilicon 1815 -811 1815 -811 0 1
rlabel polysilicon 1815 -817 1815 -817 0 3
rlabel polysilicon 1822 -811 1822 -811 0 1
rlabel polysilicon 1822 -817 1822 -817 0 3
rlabel polysilicon 1829 -811 1829 -811 0 1
rlabel polysilicon 1829 -817 1829 -817 0 3
rlabel polysilicon 1836 -811 1836 -811 0 1
rlabel polysilicon 1836 -817 1836 -817 0 3
rlabel polysilicon 1843 -811 1843 -811 0 1
rlabel polysilicon 1843 -817 1843 -817 0 3
rlabel polysilicon 1850 -811 1850 -811 0 1
rlabel polysilicon 1850 -817 1850 -817 0 3
rlabel polysilicon 1857 -811 1857 -811 0 1
rlabel polysilicon 1857 -817 1857 -817 0 3
rlabel polysilicon 1864 -811 1864 -811 0 1
rlabel polysilicon 1864 -817 1864 -817 0 3
rlabel polysilicon 1871 -811 1871 -811 0 1
rlabel polysilicon 1871 -817 1871 -817 0 3
rlabel polysilicon 1878 -811 1878 -811 0 1
rlabel polysilicon 1878 -817 1878 -817 0 3
rlabel polysilicon 1885 -811 1885 -811 0 1
rlabel polysilicon 1885 -817 1885 -817 0 3
rlabel polysilicon 1892 -811 1892 -811 0 1
rlabel polysilicon 1892 -817 1892 -817 0 3
rlabel polysilicon 1899 -811 1899 -811 0 1
rlabel polysilicon 1899 -817 1899 -817 0 3
rlabel polysilicon 1906 -811 1906 -811 0 1
rlabel polysilicon 1906 -817 1906 -817 0 3
rlabel polysilicon 1913 -811 1913 -811 0 1
rlabel polysilicon 1913 -817 1913 -817 0 3
rlabel polysilicon 1920 -811 1920 -811 0 1
rlabel polysilicon 1920 -817 1920 -817 0 3
rlabel polysilicon 1927 -811 1927 -811 0 1
rlabel polysilicon 1927 -817 1927 -817 0 3
rlabel polysilicon 1934 -811 1934 -811 0 1
rlabel polysilicon 1934 -817 1934 -817 0 3
rlabel polysilicon 1941 -811 1941 -811 0 1
rlabel polysilicon 1941 -817 1941 -817 0 3
rlabel polysilicon 1948 -811 1948 -811 0 1
rlabel polysilicon 1948 -817 1948 -817 0 3
rlabel polysilicon 1955 -811 1955 -811 0 1
rlabel polysilicon 1955 -817 1955 -817 0 3
rlabel polysilicon 1962 -811 1962 -811 0 1
rlabel polysilicon 1962 -817 1962 -817 0 3
rlabel polysilicon 1969 -811 1969 -811 0 1
rlabel polysilicon 1969 -817 1969 -817 0 3
rlabel polysilicon 1976 -811 1976 -811 0 1
rlabel polysilicon 1976 -817 1976 -817 0 3
rlabel polysilicon 1983 -811 1983 -811 0 1
rlabel polysilicon 1983 -817 1983 -817 0 3
rlabel polysilicon 1990 -811 1990 -811 0 1
rlabel polysilicon 1990 -817 1990 -817 0 3
rlabel polysilicon 1997 -811 1997 -811 0 1
rlabel polysilicon 1997 -817 1997 -817 0 3
rlabel polysilicon 2004 -811 2004 -811 0 1
rlabel polysilicon 2004 -817 2004 -817 0 3
rlabel polysilicon 2011 -811 2011 -811 0 1
rlabel polysilicon 2011 -817 2011 -817 0 3
rlabel polysilicon 2018 -811 2018 -811 0 1
rlabel polysilicon 2018 -817 2018 -817 0 3
rlabel polysilicon 2025 -811 2025 -811 0 1
rlabel polysilicon 2025 -817 2025 -817 0 3
rlabel polysilicon 2032 -811 2032 -811 0 1
rlabel polysilicon 2032 -817 2032 -817 0 3
rlabel polysilicon 2039 -811 2039 -811 0 1
rlabel polysilicon 2039 -817 2039 -817 0 3
rlabel polysilicon 2046 -811 2046 -811 0 1
rlabel polysilicon 2046 -817 2046 -817 0 3
rlabel polysilicon 2053 -811 2053 -811 0 1
rlabel polysilicon 2053 -817 2053 -817 0 3
rlabel polysilicon 2060 -811 2060 -811 0 1
rlabel polysilicon 2060 -817 2060 -817 0 3
rlabel polysilicon 2067 -811 2067 -811 0 1
rlabel polysilicon 2067 -817 2067 -817 0 3
rlabel polysilicon 2074 -811 2074 -811 0 1
rlabel polysilicon 2074 -817 2074 -817 0 3
rlabel polysilicon 2081 -811 2081 -811 0 1
rlabel polysilicon 2081 -817 2081 -817 0 3
rlabel polysilicon 2088 -811 2088 -811 0 1
rlabel polysilicon 2088 -817 2088 -817 0 3
rlabel polysilicon 2095 -811 2095 -811 0 1
rlabel polysilicon 2095 -817 2095 -817 0 3
rlabel polysilicon 2102 -811 2102 -811 0 1
rlabel polysilicon 2102 -817 2102 -817 0 3
rlabel polysilicon 2109 -811 2109 -811 0 1
rlabel polysilicon 2109 -817 2109 -817 0 3
rlabel polysilicon 2116 -811 2116 -811 0 1
rlabel polysilicon 2116 -817 2116 -817 0 3
rlabel polysilicon 2123 -811 2123 -811 0 1
rlabel polysilicon 2123 -817 2123 -817 0 3
rlabel polysilicon 2130 -811 2130 -811 0 1
rlabel polysilicon 2130 -817 2130 -817 0 3
rlabel polysilicon 2137 -811 2137 -811 0 1
rlabel polysilicon 2137 -817 2137 -817 0 3
rlabel polysilicon 2144 -811 2144 -811 0 1
rlabel polysilicon 2144 -817 2144 -817 0 3
rlabel polysilicon 2151 -811 2151 -811 0 1
rlabel polysilicon 2151 -817 2151 -817 0 3
rlabel polysilicon 2158 -811 2158 -811 0 1
rlabel polysilicon 2158 -817 2158 -817 0 3
rlabel polysilicon 2165 -811 2165 -811 0 1
rlabel polysilicon 2165 -817 2165 -817 0 3
rlabel polysilicon 2172 -811 2172 -811 0 1
rlabel polysilicon 2172 -817 2172 -817 0 3
rlabel polysilicon 2179 -811 2179 -811 0 1
rlabel polysilicon 2179 -817 2179 -817 0 3
rlabel polysilicon 2186 -811 2186 -811 0 1
rlabel polysilicon 2186 -817 2186 -817 0 3
rlabel polysilicon 2193 -811 2193 -811 0 1
rlabel polysilicon 2193 -817 2193 -817 0 3
rlabel polysilicon 2200 -811 2200 -811 0 1
rlabel polysilicon 2200 -817 2200 -817 0 3
rlabel polysilicon 2207 -811 2207 -811 0 1
rlabel polysilicon 2207 -817 2207 -817 0 3
rlabel polysilicon 2214 -811 2214 -811 0 1
rlabel polysilicon 2214 -817 2214 -817 0 3
rlabel polysilicon 2221 -811 2221 -811 0 1
rlabel polysilicon 2221 -817 2221 -817 0 3
rlabel polysilicon 2228 -811 2228 -811 0 1
rlabel polysilicon 2228 -817 2228 -817 0 3
rlabel polysilicon 2235 -811 2235 -811 0 1
rlabel polysilicon 2235 -817 2235 -817 0 3
rlabel polysilicon 2242 -811 2242 -811 0 1
rlabel polysilicon 2242 -817 2242 -817 0 3
rlabel polysilicon 2249 -811 2249 -811 0 1
rlabel polysilicon 2249 -817 2249 -817 0 3
rlabel polysilicon 2256 -811 2256 -811 0 1
rlabel polysilicon 2256 -817 2256 -817 0 3
rlabel polysilicon 2263 -811 2263 -811 0 1
rlabel polysilicon 2263 -817 2263 -817 0 3
rlabel polysilicon 2270 -811 2270 -811 0 1
rlabel polysilicon 2270 -817 2270 -817 0 3
rlabel polysilicon 2277 -811 2277 -811 0 1
rlabel polysilicon 2277 -817 2277 -817 0 3
rlabel polysilicon 2284 -811 2284 -811 0 1
rlabel polysilicon 2284 -817 2284 -817 0 3
rlabel polysilicon 2291 -811 2291 -811 0 1
rlabel polysilicon 2291 -817 2291 -817 0 3
rlabel polysilicon 2298 -811 2298 -811 0 1
rlabel polysilicon 2298 -817 2298 -817 0 3
rlabel polysilicon 2305 -811 2305 -811 0 1
rlabel polysilicon 2305 -817 2305 -817 0 3
rlabel polysilicon 2312 -811 2312 -811 0 1
rlabel polysilicon 2312 -817 2312 -817 0 3
rlabel polysilicon 2319 -811 2319 -811 0 1
rlabel polysilicon 2319 -817 2319 -817 0 3
rlabel polysilicon 2326 -811 2326 -811 0 1
rlabel polysilicon 2326 -817 2326 -817 0 3
rlabel polysilicon 2347 -811 2347 -811 0 1
rlabel polysilicon 2347 -817 2347 -817 0 3
rlabel polysilicon 2403 -811 2403 -811 0 1
rlabel polysilicon 2403 -817 2403 -817 0 3
rlabel polysilicon 2 -1000 2 -1000 0 1
rlabel polysilicon 2 -1006 2 -1006 0 3
rlabel polysilicon 9 -1000 9 -1000 0 1
rlabel polysilicon 9 -1006 9 -1006 0 3
rlabel polysilicon 16 -1000 16 -1000 0 1
rlabel polysilicon 16 -1006 16 -1006 0 3
rlabel polysilicon 23 -1000 23 -1000 0 1
rlabel polysilicon 23 -1006 23 -1006 0 3
rlabel polysilicon 30 -1000 30 -1000 0 1
rlabel polysilicon 30 -1006 30 -1006 0 3
rlabel polysilicon 37 -1000 37 -1000 0 1
rlabel polysilicon 37 -1006 37 -1006 0 3
rlabel polysilicon 44 -1000 44 -1000 0 1
rlabel polysilicon 44 -1006 44 -1006 0 3
rlabel polysilicon 51 -1000 51 -1000 0 1
rlabel polysilicon 51 -1006 51 -1006 0 3
rlabel polysilicon 58 -1000 58 -1000 0 1
rlabel polysilicon 58 -1006 58 -1006 0 3
rlabel polysilicon 65 -1000 65 -1000 0 1
rlabel polysilicon 65 -1006 65 -1006 0 3
rlabel polysilicon 72 -1000 72 -1000 0 1
rlabel polysilicon 72 -1006 72 -1006 0 3
rlabel polysilicon 79 -1000 79 -1000 0 1
rlabel polysilicon 79 -1006 79 -1006 0 3
rlabel polysilicon 86 -1000 86 -1000 0 1
rlabel polysilicon 86 -1006 86 -1006 0 3
rlabel polysilicon 93 -1006 93 -1006 0 3
rlabel polysilicon 96 -1006 96 -1006 0 4
rlabel polysilicon 100 -1000 100 -1000 0 1
rlabel polysilicon 103 -1000 103 -1000 0 2
rlabel polysilicon 100 -1006 100 -1006 0 3
rlabel polysilicon 103 -1006 103 -1006 0 4
rlabel polysilicon 107 -1000 107 -1000 0 1
rlabel polysilicon 107 -1006 107 -1006 0 3
rlabel polysilicon 114 -1000 114 -1000 0 1
rlabel polysilicon 114 -1006 114 -1006 0 3
rlabel polysilicon 121 -1000 121 -1000 0 1
rlabel polysilicon 121 -1006 121 -1006 0 3
rlabel polysilicon 128 -1000 128 -1000 0 1
rlabel polysilicon 128 -1006 128 -1006 0 3
rlabel polysilicon 135 -1000 135 -1000 0 1
rlabel polysilicon 135 -1006 135 -1006 0 3
rlabel polysilicon 138 -1006 138 -1006 0 4
rlabel polysilicon 142 -1000 142 -1000 0 1
rlabel polysilicon 142 -1006 142 -1006 0 3
rlabel polysilicon 149 -1000 149 -1000 0 1
rlabel polysilicon 149 -1006 149 -1006 0 3
rlabel polysilicon 156 -1000 156 -1000 0 1
rlabel polysilicon 156 -1006 156 -1006 0 3
rlabel polysilicon 163 -1000 163 -1000 0 1
rlabel polysilicon 163 -1006 163 -1006 0 3
rlabel polysilicon 170 -1000 170 -1000 0 1
rlabel polysilicon 170 -1006 170 -1006 0 3
rlabel polysilicon 177 -1000 177 -1000 0 1
rlabel polysilicon 180 -1000 180 -1000 0 2
rlabel polysilicon 177 -1006 177 -1006 0 3
rlabel polysilicon 180 -1006 180 -1006 0 4
rlabel polysilicon 184 -1000 184 -1000 0 1
rlabel polysilicon 187 -1000 187 -1000 0 2
rlabel polysilicon 187 -1006 187 -1006 0 4
rlabel polysilicon 191 -1000 191 -1000 0 1
rlabel polysilicon 191 -1006 191 -1006 0 3
rlabel polysilicon 198 -1000 198 -1000 0 1
rlabel polysilicon 198 -1006 198 -1006 0 3
rlabel polysilicon 205 -1000 205 -1000 0 1
rlabel polysilicon 205 -1006 205 -1006 0 3
rlabel polysilicon 212 -1000 212 -1000 0 1
rlabel polysilicon 212 -1006 212 -1006 0 3
rlabel polysilicon 219 -1000 219 -1000 0 1
rlabel polysilicon 222 -1000 222 -1000 0 2
rlabel polysilicon 222 -1006 222 -1006 0 4
rlabel polysilicon 226 -1000 226 -1000 0 1
rlabel polysilicon 226 -1006 226 -1006 0 3
rlabel polysilicon 233 -1000 233 -1000 0 1
rlabel polysilicon 233 -1006 233 -1006 0 3
rlabel polysilicon 240 -1000 240 -1000 0 1
rlabel polysilicon 240 -1006 240 -1006 0 3
rlabel polysilicon 247 -1000 247 -1000 0 1
rlabel polysilicon 247 -1006 247 -1006 0 3
rlabel polysilicon 254 -1000 254 -1000 0 1
rlabel polysilicon 254 -1006 254 -1006 0 3
rlabel polysilicon 261 -1000 261 -1000 0 1
rlabel polysilicon 261 -1006 261 -1006 0 3
rlabel polysilicon 268 -1000 268 -1000 0 1
rlabel polysilicon 271 -1000 271 -1000 0 2
rlabel polysilicon 271 -1006 271 -1006 0 4
rlabel polysilicon 275 -1000 275 -1000 0 1
rlabel polysilicon 275 -1006 275 -1006 0 3
rlabel polysilicon 282 -1000 282 -1000 0 1
rlabel polysilicon 282 -1006 282 -1006 0 3
rlabel polysilicon 289 -1000 289 -1000 0 1
rlabel polysilicon 289 -1006 289 -1006 0 3
rlabel polysilicon 296 -1000 296 -1000 0 1
rlabel polysilicon 296 -1006 296 -1006 0 3
rlabel polysilicon 303 -1000 303 -1000 0 1
rlabel polysilicon 303 -1006 303 -1006 0 3
rlabel polysilicon 310 -1000 310 -1000 0 1
rlabel polysilicon 310 -1006 310 -1006 0 3
rlabel polysilicon 317 -1000 317 -1000 0 1
rlabel polysilicon 317 -1006 317 -1006 0 3
rlabel polysilicon 324 -1000 324 -1000 0 1
rlabel polysilicon 324 -1006 324 -1006 0 3
rlabel polysilicon 331 -1000 331 -1000 0 1
rlabel polysilicon 331 -1006 331 -1006 0 3
rlabel polysilicon 338 -1000 338 -1000 0 1
rlabel polysilicon 338 -1006 338 -1006 0 3
rlabel polysilicon 345 -1000 345 -1000 0 1
rlabel polysilicon 345 -1006 345 -1006 0 3
rlabel polysilicon 352 -1000 352 -1000 0 1
rlabel polysilicon 352 -1006 352 -1006 0 3
rlabel polysilicon 359 -1000 359 -1000 0 1
rlabel polysilicon 359 -1006 359 -1006 0 3
rlabel polysilicon 366 -1000 366 -1000 0 1
rlabel polysilicon 366 -1006 366 -1006 0 3
rlabel polysilicon 373 -1000 373 -1000 0 1
rlabel polysilicon 376 -1000 376 -1000 0 2
rlabel polysilicon 373 -1006 373 -1006 0 3
rlabel polysilicon 376 -1006 376 -1006 0 4
rlabel polysilicon 380 -1000 380 -1000 0 1
rlabel polysilicon 380 -1006 380 -1006 0 3
rlabel polysilicon 387 -1000 387 -1000 0 1
rlabel polysilicon 390 -1000 390 -1000 0 2
rlabel polysilicon 390 -1006 390 -1006 0 4
rlabel polysilicon 394 -1000 394 -1000 0 1
rlabel polysilicon 394 -1006 394 -1006 0 3
rlabel polysilicon 401 -1000 401 -1000 0 1
rlabel polysilicon 401 -1006 401 -1006 0 3
rlabel polysilicon 408 -1000 408 -1000 0 1
rlabel polysilicon 408 -1006 408 -1006 0 3
rlabel polysilicon 415 -1000 415 -1000 0 1
rlabel polysilicon 415 -1006 415 -1006 0 3
rlabel polysilicon 422 -1000 422 -1000 0 1
rlabel polysilicon 422 -1006 422 -1006 0 3
rlabel polysilicon 429 -1000 429 -1000 0 1
rlabel polysilicon 429 -1006 429 -1006 0 3
rlabel polysilicon 436 -1000 436 -1000 0 1
rlabel polysilicon 436 -1006 436 -1006 0 3
rlabel polysilicon 443 -1000 443 -1000 0 1
rlabel polysilicon 443 -1006 443 -1006 0 3
rlabel polysilicon 450 -1000 450 -1000 0 1
rlabel polysilicon 450 -1006 450 -1006 0 3
rlabel polysilicon 457 -1000 457 -1000 0 1
rlabel polysilicon 457 -1006 457 -1006 0 3
rlabel polysilicon 464 -1000 464 -1000 0 1
rlabel polysilicon 464 -1006 464 -1006 0 3
rlabel polysilicon 471 -1000 471 -1000 0 1
rlabel polysilicon 471 -1006 471 -1006 0 3
rlabel polysilicon 478 -1000 478 -1000 0 1
rlabel polysilicon 478 -1006 478 -1006 0 3
rlabel polysilicon 485 -1000 485 -1000 0 1
rlabel polysilicon 485 -1006 485 -1006 0 3
rlabel polysilicon 492 -1000 492 -1000 0 1
rlabel polysilicon 492 -1006 492 -1006 0 3
rlabel polysilicon 499 -1000 499 -1000 0 1
rlabel polysilicon 499 -1006 499 -1006 0 3
rlabel polysilicon 506 -1000 506 -1000 0 1
rlabel polysilicon 506 -1006 506 -1006 0 3
rlabel polysilicon 513 -1000 513 -1000 0 1
rlabel polysilicon 513 -1006 513 -1006 0 3
rlabel polysilicon 520 -1000 520 -1000 0 1
rlabel polysilicon 520 -1006 520 -1006 0 3
rlabel polysilicon 527 -1000 527 -1000 0 1
rlabel polysilicon 530 -1000 530 -1000 0 2
rlabel polysilicon 534 -1000 534 -1000 0 1
rlabel polysilicon 534 -1006 534 -1006 0 3
rlabel polysilicon 541 -1000 541 -1000 0 1
rlabel polysilicon 541 -1006 541 -1006 0 3
rlabel polysilicon 548 -1000 548 -1000 0 1
rlabel polysilicon 548 -1006 548 -1006 0 3
rlabel polysilicon 555 -1000 555 -1000 0 1
rlabel polysilicon 555 -1006 555 -1006 0 3
rlabel polysilicon 562 -1000 562 -1000 0 1
rlabel polysilicon 562 -1006 562 -1006 0 3
rlabel polysilicon 569 -1000 569 -1000 0 1
rlabel polysilicon 569 -1006 569 -1006 0 3
rlabel polysilicon 576 -1000 576 -1000 0 1
rlabel polysilicon 576 -1006 576 -1006 0 3
rlabel polysilicon 583 -1000 583 -1000 0 1
rlabel polysilicon 583 -1006 583 -1006 0 3
rlabel polysilicon 590 -1000 590 -1000 0 1
rlabel polysilicon 590 -1006 590 -1006 0 3
rlabel polysilicon 597 -1000 597 -1000 0 1
rlabel polysilicon 597 -1006 597 -1006 0 3
rlabel polysilicon 604 -1000 604 -1000 0 1
rlabel polysilicon 604 -1006 604 -1006 0 3
rlabel polysilicon 611 -1000 611 -1000 0 1
rlabel polysilicon 614 -1000 614 -1000 0 2
rlabel polysilicon 611 -1006 611 -1006 0 3
rlabel polysilicon 618 -1000 618 -1000 0 1
rlabel polysilicon 618 -1006 618 -1006 0 3
rlabel polysilicon 625 -1000 625 -1000 0 1
rlabel polysilicon 628 -1000 628 -1000 0 2
rlabel polysilicon 625 -1006 625 -1006 0 3
rlabel polysilicon 628 -1006 628 -1006 0 4
rlabel polysilicon 632 -1000 632 -1000 0 1
rlabel polysilicon 635 -1000 635 -1000 0 2
rlabel polysilicon 632 -1006 632 -1006 0 3
rlabel polysilicon 635 -1006 635 -1006 0 4
rlabel polysilicon 639 -1000 639 -1000 0 1
rlabel polysilicon 639 -1006 639 -1006 0 3
rlabel polysilicon 646 -1000 646 -1000 0 1
rlabel polysilicon 646 -1006 646 -1006 0 3
rlabel polysilicon 653 -1000 653 -1000 0 1
rlabel polysilicon 653 -1006 653 -1006 0 3
rlabel polysilicon 660 -1000 660 -1000 0 1
rlabel polysilicon 660 -1006 660 -1006 0 3
rlabel polysilicon 667 -1000 667 -1000 0 1
rlabel polysilicon 667 -1006 667 -1006 0 3
rlabel polysilicon 674 -1000 674 -1000 0 1
rlabel polysilicon 674 -1006 674 -1006 0 3
rlabel polysilicon 681 -1000 681 -1000 0 1
rlabel polysilicon 681 -1006 681 -1006 0 3
rlabel polysilicon 688 -1000 688 -1000 0 1
rlabel polysilicon 688 -1006 688 -1006 0 3
rlabel polysilicon 695 -1000 695 -1000 0 1
rlabel polysilicon 695 -1006 695 -1006 0 3
rlabel polysilicon 702 -1000 702 -1000 0 1
rlabel polysilicon 702 -1006 702 -1006 0 3
rlabel polysilicon 709 -1000 709 -1000 0 1
rlabel polysilicon 709 -1006 709 -1006 0 3
rlabel polysilicon 716 -1000 716 -1000 0 1
rlabel polysilicon 719 -1000 719 -1000 0 2
rlabel polysilicon 719 -1006 719 -1006 0 4
rlabel polysilicon 723 -1000 723 -1000 0 1
rlabel polysilicon 723 -1006 723 -1006 0 3
rlabel polysilicon 730 -1000 730 -1000 0 1
rlabel polysilicon 730 -1006 730 -1006 0 3
rlabel polysilicon 737 -1000 737 -1000 0 1
rlabel polysilicon 737 -1006 737 -1006 0 3
rlabel polysilicon 744 -1000 744 -1000 0 1
rlabel polysilicon 744 -1006 744 -1006 0 3
rlabel polysilicon 751 -1000 751 -1000 0 1
rlabel polysilicon 751 -1006 751 -1006 0 3
rlabel polysilicon 758 -1000 758 -1000 0 1
rlabel polysilicon 758 -1006 758 -1006 0 3
rlabel polysilicon 765 -1000 765 -1000 0 1
rlabel polysilicon 765 -1006 765 -1006 0 3
rlabel polysilicon 772 -1000 772 -1000 0 1
rlabel polysilicon 775 -1000 775 -1000 0 2
rlabel polysilicon 772 -1006 772 -1006 0 3
rlabel polysilicon 775 -1006 775 -1006 0 4
rlabel polysilicon 782 -1000 782 -1000 0 2
rlabel polysilicon 779 -1006 779 -1006 0 3
rlabel polysilicon 782 -1006 782 -1006 0 4
rlabel polysilicon 786 -1000 786 -1000 0 1
rlabel polysilicon 786 -1006 786 -1006 0 3
rlabel polysilicon 793 -1000 793 -1000 0 1
rlabel polysilicon 796 -1000 796 -1000 0 2
rlabel polysilicon 793 -1006 793 -1006 0 3
rlabel polysilicon 796 -1006 796 -1006 0 4
rlabel polysilicon 800 -1000 800 -1000 0 1
rlabel polysilicon 800 -1006 800 -1006 0 3
rlabel polysilicon 807 -1000 807 -1000 0 1
rlabel polysilicon 807 -1006 807 -1006 0 3
rlabel polysilicon 814 -1000 814 -1000 0 1
rlabel polysilicon 817 -1000 817 -1000 0 2
rlabel polysilicon 814 -1006 814 -1006 0 3
rlabel polysilicon 817 -1006 817 -1006 0 4
rlabel polysilicon 821 -1000 821 -1000 0 1
rlabel polysilicon 821 -1006 821 -1006 0 3
rlabel polysilicon 828 -1000 828 -1000 0 1
rlabel polysilicon 828 -1006 828 -1006 0 3
rlabel polysilicon 831 -1006 831 -1006 0 4
rlabel polysilicon 835 -1000 835 -1000 0 1
rlabel polysilicon 835 -1006 835 -1006 0 3
rlabel polysilicon 842 -1000 842 -1000 0 1
rlabel polysilicon 842 -1006 842 -1006 0 3
rlabel polysilicon 849 -1000 849 -1000 0 1
rlabel polysilicon 849 -1006 849 -1006 0 3
rlabel polysilicon 856 -1000 856 -1000 0 1
rlabel polysilicon 856 -1006 856 -1006 0 3
rlabel polysilicon 863 -1000 863 -1000 0 1
rlabel polysilicon 863 -1006 863 -1006 0 3
rlabel polysilicon 870 -1000 870 -1000 0 1
rlabel polysilicon 870 -1006 870 -1006 0 3
rlabel polysilicon 877 -1000 877 -1000 0 1
rlabel polysilicon 877 -1006 877 -1006 0 3
rlabel polysilicon 884 -1000 884 -1000 0 1
rlabel polysilicon 884 -1006 884 -1006 0 3
rlabel polysilicon 891 -1000 891 -1000 0 1
rlabel polysilicon 891 -1006 891 -1006 0 3
rlabel polysilicon 898 -1000 898 -1000 0 1
rlabel polysilicon 898 -1006 898 -1006 0 3
rlabel polysilicon 905 -1000 905 -1000 0 1
rlabel polysilicon 905 -1006 905 -1006 0 3
rlabel polysilicon 912 -1000 912 -1000 0 1
rlabel polysilicon 912 -1006 912 -1006 0 3
rlabel polysilicon 919 -1000 919 -1000 0 1
rlabel polysilicon 919 -1006 919 -1006 0 3
rlabel polysilicon 926 -1000 926 -1000 0 1
rlabel polysilicon 926 -1006 926 -1006 0 3
rlabel polysilicon 933 -1000 933 -1000 0 1
rlabel polysilicon 936 -1000 936 -1000 0 2
rlabel polysilicon 936 -1006 936 -1006 0 4
rlabel polysilicon 940 -1000 940 -1000 0 1
rlabel polysilicon 940 -1006 940 -1006 0 3
rlabel polysilicon 947 -1000 947 -1000 0 1
rlabel polysilicon 947 -1006 947 -1006 0 3
rlabel polysilicon 954 -1000 954 -1000 0 1
rlabel polysilicon 954 -1006 954 -1006 0 3
rlabel polysilicon 957 -1006 957 -1006 0 4
rlabel polysilicon 961 -1000 961 -1000 0 1
rlabel polysilicon 961 -1006 961 -1006 0 3
rlabel polysilicon 968 -1000 968 -1000 0 1
rlabel polysilicon 968 -1006 968 -1006 0 3
rlabel polysilicon 975 -1000 975 -1000 0 1
rlabel polysilicon 975 -1006 975 -1006 0 3
rlabel polysilicon 982 -1000 982 -1000 0 1
rlabel polysilicon 982 -1006 982 -1006 0 3
rlabel polysilicon 989 -1000 989 -1000 0 1
rlabel polysilicon 989 -1006 989 -1006 0 3
rlabel polysilicon 996 -1000 996 -1000 0 1
rlabel polysilicon 996 -1006 996 -1006 0 3
rlabel polysilicon 1003 -1000 1003 -1000 0 1
rlabel polysilicon 1003 -1006 1003 -1006 0 3
rlabel polysilicon 1010 -1000 1010 -1000 0 1
rlabel polysilicon 1010 -1006 1010 -1006 0 3
rlabel polysilicon 1017 -1000 1017 -1000 0 1
rlabel polysilicon 1020 -1000 1020 -1000 0 2
rlabel polysilicon 1017 -1006 1017 -1006 0 3
rlabel polysilicon 1020 -1006 1020 -1006 0 4
rlabel polysilicon 1024 -1000 1024 -1000 0 1
rlabel polysilicon 1024 -1006 1024 -1006 0 3
rlabel polysilicon 1031 -1000 1031 -1000 0 1
rlabel polysilicon 1031 -1006 1031 -1006 0 3
rlabel polysilicon 1041 -1000 1041 -1000 0 2
rlabel polysilicon 1038 -1006 1038 -1006 0 3
rlabel polysilicon 1041 -1006 1041 -1006 0 4
rlabel polysilicon 1045 -1000 1045 -1000 0 1
rlabel polysilicon 1045 -1006 1045 -1006 0 3
rlabel polysilicon 1052 -1000 1052 -1000 0 1
rlabel polysilicon 1055 -1000 1055 -1000 0 2
rlabel polysilicon 1052 -1006 1052 -1006 0 3
rlabel polysilicon 1055 -1006 1055 -1006 0 4
rlabel polysilicon 1059 -1000 1059 -1000 0 1
rlabel polysilicon 1062 -1006 1062 -1006 0 4
rlabel polysilicon 1066 -1000 1066 -1000 0 1
rlabel polysilicon 1066 -1006 1066 -1006 0 3
rlabel polysilicon 1073 -1000 1073 -1000 0 1
rlabel polysilicon 1073 -1006 1073 -1006 0 3
rlabel polysilicon 1080 -1000 1080 -1000 0 1
rlabel polysilicon 1080 -1006 1080 -1006 0 3
rlabel polysilicon 1087 -1000 1087 -1000 0 1
rlabel polysilicon 1087 -1006 1087 -1006 0 3
rlabel polysilicon 1094 -1000 1094 -1000 0 1
rlabel polysilicon 1094 -1006 1094 -1006 0 3
rlabel polysilicon 1101 -1000 1101 -1000 0 1
rlabel polysilicon 1101 -1006 1101 -1006 0 3
rlabel polysilicon 1108 -1000 1108 -1000 0 1
rlabel polysilicon 1108 -1006 1108 -1006 0 3
rlabel polysilicon 1115 -1000 1115 -1000 0 1
rlabel polysilicon 1115 -1006 1115 -1006 0 3
rlabel polysilicon 1122 -1000 1122 -1000 0 1
rlabel polysilicon 1125 -1000 1125 -1000 0 2
rlabel polysilicon 1122 -1006 1122 -1006 0 3
rlabel polysilicon 1125 -1006 1125 -1006 0 4
rlabel polysilicon 1129 -1000 1129 -1000 0 1
rlabel polysilicon 1129 -1006 1129 -1006 0 3
rlabel polysilicon 1136 -1000 1136 -1000 0 1
rlabel polysilicon 1136 -1006 1136 -1006 0 3
rlabel polysilicon 1143 -1000 1143 -1000 0 1
rlabel polysilicon 1143 -1006 1143 -1006 0 3
rlabel polysilicon 1150 -1000 1150 -1000 0 1
rlabel polysilicon 1150 -1006 1150 -1006 0 3
rlabel polysilicon 1157 -1000 1157 -1000 0 1
rlabel polysilicon 1157 -1006 1157 -1006 0 3
rlabel polysilicon 1164 -1000 1164 -1000 0 1
rlabel polysilicon 1164 -1006 1164 -1006 0 3
rlabel polysilicon 1171 -1000 1171 -1000 0 1
rlabel polysilicon 1174 -1000 1174 -1000 0 2
rlabel polysilicon 1171 -1006 1171 -1006 0 3
rlabel polysilicon 1174 -1006 1174 -1006 0 4
rlabel polysilicon 1178 -1000 1178 -1000 0 1
rlabel polysilicon 1178 -1006 1178 -1006 0 3
rlabel polysilicon 1185 -1000 1185 -1000 0 1
rlabel polysilicon 1185 -1006 1185 -1006 0 3
rlabel polysilicon 1192 -1000 1192 -1000 0 1
rlabel polysilicon 1195 -1000 1195 -1000 0 2
rlabel polysilicon 1192 -1006 1192 -1006 0 3
rlabel polysilicon 1195 -1006 1195 -1006 0 4
rlabel polysilicon 1199 -1000 1199 -1000 0 1
rlabel polysilicon 1199 -1006 1199 -1006 0 3
rlabel polysilicon 1206 -1000 1206 -1000 0 1
rlabel polysilicon 1206 -1006 1206 -1006 0 3
rlabel polysilicon 1213 -1000 1213 -1000 0 1
rlabel polysilicon 1213 -1006 1213 -1006 0 3
rlabel polysilicon 1220 -1000 1220 -1000 0 1
rlabel polysilicon 1220 -1006 1220 -1006 0 3
rlabel polysilicon 1227 -1000 1227 -1000 0 1
rlabel polysilicon 1227 -1006 1227 -1006 0 3
rlabel polysilicon 1234 -1000 1234 -1000 0 1
rlabel polysilicon 1234 -1006 1234 -1006 0 3
rlabel polysilicon 1241 -1000 1241 -1000 0 1
rlabel polysilicon 1244 -1000 1244 -1000 0 2
rlabel polysilicon 1241 -1006 1241 -1006 0 3
rlabel polysilicon 1244 -1006 1244 -1006 0 4
rlabel polysilicon 1248 -1000 1248 -1000 0 1
rlabel polysilicon 1248 -1006 1248 -1006 0 3
rlabel polysilicon 1255 -1000 1255 -1000 0 1
rlabel polysilicon 1255 -1006 1255 -1006 0 3
rlabel polysilicon 1262 -1000 1262 -1000 0 1
rlabel polysilicon 1262 -1006 1262 -1006 0 3
rlabel polysilicon 1269 -1000 1269 -1000 0 1
rlabel polysilicon 1272 -1000 1272 -1000 0 2
rlabel polysilicon 1269 -1006 1269 -1006 0 3
rlabel polysilicon 1272 -1006 1272 -1006 0 4
rlabel polysilicon 1276 -1000 1276 -1000 0 1
rlabel polysilicon 1276 -1006 1276 -1006 0 3
rlabel polysilicon 1283 -1000 1283 -1000 0 1
rlabel polysilicon 1286 -1000 1286 -1000 0 2
rlabel polysilicon 1283 -1006 1283 -1006 0 3
rlabel polysilicon 1286 -1006 1286 -1006 0 4
rlabel polysilicon 1290 -1000 1290 -1000 0 1
rlabel polysilicon 1290 -1006 1290 -1006 0 3
rlabel polysilicon 1297 -1000 1297 -1000 0 1
rlabel polysilicon 1297 -1006 1297 -1006 0 3
rlabel polysilicon 1304 -1000 1304 -1000 0 1
rlabel polysilicon 1304 -1006 1304 -1006 0 3
rlabel polysilicon 1311 -1000 1311 -1000 0 1
rlabel polysilicon 1314 -1000 1314 -1000 0 2
rlabel polysilicon 1311 -1006 1311 -1006 0 3
rlabel polysilicon 1314 -1006 1314 -1006 0 4
rlabel polysilicon 1318 -1000 1318 -1000 0 1
rlabel polysilicon 1318 -1006 1318 -1006 0 3
rlabel polysilicon 1325 -1000 1325 -1000 0 1
rlabel polysilicon 1325 -1006 1325 -1006 0 3
rlabel polysilicon 1332 -1000 1332 -1000 0 1
rlabel polysilicon 1332 -1006 1332 -1006 0 3
rlabel polysilicon 1339 -1000 1339 -1000 0 1
rlabel polysilicon 1339 -1006 1339 -1006 0 3
rlabel polysilicon 1346 -1000 1346 -1000 0 1
rlabel polysilicon 1346 -1006 1346 -1006 0 3
rlabel polysilicon 1353 -1000 1353 -1000 0 1
rlabel polysilicon 1353 -1006 1353 -1006 0 3
rlabel polysilicon 1360 -1000 1360 -1000 0 1
rlabel polysilicon 1360 -1006 1360 -1006 0 3
rlabel polysilicon 1367 -1000 1367 -1000 0 1
rlabel polysilicon 1367 -1006 1367 -1006 0 3
rlabel polysilicon 1374 -1000 1374 -1000 0 1
rlabel polysilicon 1374 -1006 1374 -1006 0 3
rlabel polysilicon 1381 -1000 1381 -1000 0 1
rlabel polysilicon 1381 -1006 1381 -1006 0 3
rlabel polysilicon 1388 -1000 1388 -1000 0 1
rlabel polysilicon 1388 -1006 1388 -1006 0 3
rlabel polysilicon 1395 -1000 1395 -1000 0 1
rlabel polysilicon 1398 -1000 1398 -1000 0 2
rlabel polysilicon 1395 -1006 1395 -1006 0 3
rlabel polysilicon 1398 -1006 1398 -1006 0 4
rlabel polysilicon 1402 -1000 1402 -1000 0 1
rlabel polysilicon 1402 -1006 1402 -1006 0 3
rlabel polysilicon 1409 -1000 1409 -1000 0 1
rlabel polysilicon 1409 -1006 1409 -1006 0 3
rlabel polysilicon 1416 -1000 1416 -1000 0 1
rlabel polysilicon 1416 -1006 1416 -1006 0 3
rlabel polysilicon 1423 -1000 1423 -1000 0 1
rlabel polysilicon 1423 -1006 1423 -1006 0 3
rlabel polysilicon 1430 -1000 1430 -1000 0 1
rlabel polysilicon 1430 -1006 1430 -1006 0 3
rlabel polysilicon 1437 -1000 1437 -1000 0 1
rlabel polysilicon 1437 -1006 1437 -1006 0 3
rlabel polysilicon 1444 -1000 1444 -1000 0 1
rlabel polysilicon 1444 -1006 1444 -1006 0 3
rlabel polysilicon 1451 -1000 1451 -1000 0 1
rlabel polysilicon 1451 -1006 1451 -1006 0 3
rlabel polysilicon 1458 -1000 1458 -1000 0 1
rlabel polysilicon 1458 -1006 1458 -1006 0 3
rlabel polysilicon 1465 -1000 1465 -1000 0 1
rlabel polysilicon 1465 -1006 1465 -1006 0 3
rlabel polysilicon 1472 -1000 1472 -1000 0 1
rlabel polysilicon 1472 -1006 1472 -1006 0 3
rlabel polysilicon 1479 -1000 1479 -1000 0 1
rlabel polysilicon 1479 -1006 1479 -1006 0 3
rlabel polysilicon 1486 -1000 1486 -1000 0 1
rlabel polysilicon 1486 -1006 1486 -1006 0 3
rlabel polysilicon 1493 -1000 1493 -1000 0 1
rlabel polysilicon 1493 -1006 1493 -1006 0 3
rlabel polysilicon 1500 -1000 1500 -1000 0 1
rlabel polysilicon 1500 -1006 1500 -1006 0 3
rlabel polysilicon 1507 -1000 1507 -1000 0 1
rlabel polysilicon 1507 -1006 1507 -1006 0 3
rlabel polysilicon 1514 -1000 1514 -1000 0 1
rlabel polysilicon 1517 -1000 1517 -1000 0 2
rlabel polysilicon 1514 -1006 1514 -1006 0 3
rlabel polysilicon 1517 -1006 1517 -1006 0 4
rlabel polysilicon 1521 -1000 1521 -1000 0 1
rlabel polysilicon 1521 -1006 1521 -1006 0 3
rlabel polysilicon 1528 -1000 1528 -1000 0 1
rlabel polysilicon 1528 -1006 1528 -1006 0 3
rlabel polysilicon 1535 -1000 1535 -1000 0 1
rlabel polysilicon 1535 -1006 1535 -1006 0 3
rlabel polysilicon 1542 -1000 1542 -1000 0 1
rlabel polysilicon 1542 -1006 1542 -1006 0 3
rlabel polysilicon 1549 -1000 1549 -1000 0 1
rlabel polysilicon 1549 -1006 1549 -1006 0 3
rlabel polysilicon 1556 -1000 1556 -1000 0 1
rlabel polysilicon 1556 -1006 1556 -1006 0 3
rlabel polysilicon 1563 -1000 1563 -1000 0 1
rlabel polysilicon 1563 -1006 1563 -1006 0 3
rlabel polysilicon 1570 -1000 1570 -1000 0 1
rlabel polysilicon 1573 -1000 1573 -1000 0 2
rlabel polysilicon 1570 -1006 1570 -1006 0 3
rlabel polysilicon 1577 -1000 1577 -1000 0 1
rlabel polysilicon 1580 -1006 1580 -1006 0 4
rlabel polysilicon 1584 -1000 1584 -1000 0 1
rlabel polysilicon 1584 -1006 1584 -1006 0 3
rlabel polysilicon 1591 -1000 1591 -1000 0 1
rlabel polysilicon 1591 -1006 1591 -1006 0 3
rlabel polysilicon 1598 -1000 1598 -1000 0 1
rlabel polysilicon 1598 -1006 1598 -1006 0 3
rlabel polysilicon 1605 -1000 1605 -1000 0 1
rlabel polysilicon 1605 -1006 1605 -1006 0 3
rlabel polysilicon 1612 -1000 1612 -1000 0 1
rlabel polysilicon 1612 -1006 1612 -1006 0 3
rlabel polysilicon 1619 -1000 1619 -1000 0 1
rlabel polysilicon 1619 -1006 1619 -1006 0 3
rlabel polysilicon 1626 -1000 1626 -1000 0 1
rlabel polysilicon 1626 -1006 1626 -1006 0 3
rlabel polysilicon 1633 -1000 1633 -1000 0 1
rlabel polysilicon 1633 -1006 1633 -1006 0 3
rlabel polysilicon 1640 -1000 1640 -1000 0 1
rlabel polysilicon 1640 -1006 1640 -1006 0 3
rlabel polysilicon 1647 -1000 1647 -1000 0 1
rlabel polysilicon 1647 -1006 1647 -1006 0 3
rlabel polysilicon 1654 -1000 1654 -1000 0 1
rlabel polysilicon 1654 -1006 1654 -1006 0 3
rlabel polysilicon 1661 -1000 1661 -1000 0 1
rlabel polysilicon 1661 -1006 1661 -1006 0 3
rlabel polysilicon 1668 -1000 1668 -1000 0 1
rlabel polysilicon 1668 -1006 1668 -1006 0 3
rlabel polysilicon 1675 -1000 1675 -1000 0 1
rlabel polysilicon 1675 -1006 1675 -1006 0 3
rlabel polysilicon 1682 -1000 1682 -1000 0 1
rlabel polysilicon 1682 -1006 1682 -1006 0 3
rlabel polysilicon 1689 -1000 1689 -1000 0 1
rlabel polysilicon 1689 -1006 1689 -1006 0 3
rlabel polysilicon 1696 -1000 1696 -1000 0 1
rlabel polysilicon 1696 -1006 1696 -1006 0 3
rlabel polysilicon 1703 -1000 1703 -1000 0 1
rlabel polysilicon 1703 -1006 1703 -1006 0 3
rlabel polysilicon 1710 -1000 1710 -1000 0 1
rlabel polysilicon 1710 -1006 1710 -1006 0 3
rlabel polysilicon 1717 -1000 1717 -1000 0 1
rlabel polysilicon 1717 -1006 1717 -1006 0 3
rlabel polysilicon 1724 -1000 1724 -1000 0 1
rlabel polysilicon 1724 -1006 1724 -1006 0 3
rlabel polysilicon 1731 -1000 1731 -1000 0 1
rlabel polysilicon 1731 -1006 1731 -1006 0 3
rlabel polysilicon 1738 -1000 1738 -1000 0 1
rlabel polysilicon 1738 -1006 1738 -1006 0 3
rlabel polysilicon 1745 -1000 1745 -1000 0 1
rlabel polysilicon 1745 -1006 1745 -1006 0 3
rlabel polysilicon 1752 -1000 1752 -1000 0 1
rlabel polysilicon 1752 -1006 1752 -1006 0 3
rlabel polysilicon 1759 -1000 1759 -1000 0 1
rlabel polysilicon 1759 -1006 1759 -1006 0 3
rlabel polysilicon 1766 -1000 1766 -1000 0 1
rlabel polysilicon 1766 -1006 1766 -1006 0 3
rlabel polysilicon 1773 -1000 1773 -1000 0 1
rlabel polysilicon 1773 -1006 1773 -1006 0 3
rlabel polysilicon 1780 -1000 1780 -1000 0 1
rlabel polysilicon 1780 -1006 1780 -1006 0 3
rlabel polysilicon 1787 -1000 1787 -1000 0 1
rlabel polysilicon 1787 -1006 1787 -1006 0 3
rlabel polysilicon 1794 -1000 1794 -1000 0 1
rlabel polysilicon 1794 -1006 1794 -1006 0 3
rlabel polysilicon 1801 -1000 1801 -1000 0 1
rlabel polysilicon 1801 -1006 1801 -1006 0 3
rlabel polysilicon 1808 -1000 1808 -1000 0 1
rlabel polysilicon 1808 -1006 1808 -1006 0 3
rlabel polysilicon 1815 -1000 1815 -1000 0 1
rlabel polysilicon 1815 -1006 1815 -1006 0 3
rlabel polysilicon 1822 -1000 1822 -1000 0 1
rlabel polysilicon 1822 -1006 1822 -1006 0 3
rlabel polysilicon 1829 -1000 1829 -1000 0 1
rlabel polysilicon 1829 -1006 1829 -1006 0 3
rlabel polysilicon 1836 -1000 1836 -1000 0 1
rlabel polysilicon 1836 -1006 1836 -1006 0 3
rlabel polysilicon 1843 -1000 1843 -1000 0 1
rlabel polysilicon 1843 -1006 1843 -1006 0 3
rlabel polysilicon 1850 -1000 1850 -1000 0 1
rlabel polysilicon 1850 -1006 1850 -1006 0 3
rlabel polysilicon 1857 -1000 1857 -1000 0 1
rlabel polysilicon 1857 -1006 1857 -1006 0 3
rlabel polysilicon 1864 -1000 1864 -1000 0 1
rlabel polysilicon 1864 -1006 1864 -1006 0 3
rlabel polysilicon 1871 -1000 1871 -1000 0 1
rlabel polysilicon 1871 -1006 1871 -1006 0 3
rlabel polysilicon 1878 -1000 1878 -1000 0 1
rlabel polysilicon 1878 -1006 1878 -1006 0 3
rlabel polysilicon 1885 -1000 1885 -1000 0 1
rlabel polysilicon 1885 -1006 1885 -1006 0 3
rlabel polysilicon 1892 -1000 1892 -1000 0 1
rlabel polysilicon 1892 -1006 1892 -1006 0 3
rlabel polysilicon 1899 -1000 1899 -1000 0 1
rlabel polysilicon 1899 -1006 1899 -1006 0 3
rlabel polysilicon 1906 -1000 1906 -1000 0 1
rlabel polysilicon 1906 -1006 1906 -1006 0 3
rlabel polysilicon 1913 -1000 1913 -1000 0 1
rlabel polysilicon 1913 -1006 1913 -1006 0 3
rlabel polysilicon 1920 -1000 1920 -1000 0 1
rlabel polysilicon 1920 -1006 1920 -1006 0 3
rlabel polysilicon 1927 -1000 1927 -1000 0 1
rlabel polysilicon 1927 -1006 1927 -1006 0 3
rlabel polysilicon 1934 -1000 1934 -1000 0 1
rlabel polysilicon 1934 -1006 1934 -1006 0 3
rlabel polysilicon 1941 -1000 1941 -1000 0 1
rlabel polysilicon 1941 -1006 1941 -1006 0 3
rlabel polysilicon 1948 -1000 1948 -1000 0 1
rlabel polysilicon 1948 -1006 1948 -1006 0 3
rlabel polysilicon 1955 -1000 1955 -1000 0 1
rlabel polysilicon 1955 -1006 1955 -1006 0 3
rlabel polysilicon 1962 -1000 1962 -1000 0 1
rlabel polysilicon 1962 -1006 1962 -1006 0 3
rlabel polysilicon 1969 -1000 1969 -1000 0 1
rlabel polysilicon 1969 -1006 1969 -1006 0 3
rlabel polysilicon 1976 -1000 1976 -1000 0 1
rlabel polysilicon 1976 -1006 1976 -1006 0 3
rlabel polysilicon 1983 -1000 1983 -1000 0 1
rlabel polysilicon 1983 -1006 1983 -1006 0 3
rlabel polysilicon 1990 -1000 1990 -1000 0 1
rlabel polysilicon 1990 -1006 1990 -1006 0 3
rlabel polysilicon 1997 -1000 1997 -1000 0 1
rlabel polysilicon 1997 -1006 1997 -1006 0 3
rlabel polysilicon 2004 -1000 2004 -1000 0 1
rlabel polysilicon 2004 -1006 2004 -1006 0 3
rlabel polysilicon 2011 -1000 2011 -1000 0 1
rlabel polysilicon 2011 -1006 2011 -1006 0 3
rlabel polysilicon 2018 -1000 2018 -1000 0 1
rlabel polysilicon 2018 -1006 2018 -1006 0 3
rlabel polysilicon 2025 -1000 2025 -1000 0 1
rlabel polysilicon 2025 -1006 2025 -1006 0 3
rlabel polysilicon 2032 -1000 2032 -1000 0 1
rlabel polysilicon 2032 -1006 2032 -1006 0 3
rlabel polysilicon 2039 -1000 2039 -1000 0 1
rlabel polysilicon 2039 -1006 2039 -1006 0 3
rlabel polysilicon 2046 -1000 2046 -1000 0 1
rlabel polysilicon 2046 -1006 2046 -1006 0 3
rlabel polysilicon 2053 -1000 2053 -1000 0 1
rlabel polysilicon 2053 -1006 2053 -1006 0 3
rlabel polysilicon 2060 -1000 2060 -1000 0 1
rlabel polysilicon 2060 -1006 2060 -1006 0 3
rlabel polysilicon 2067 -1000 2067 -1000 0 1
rlabel polysilicon 2067 -1006 2067 -1006 0 3
rlabel polysilicon 2074 -1000 2074 -1000 0 1
rlabel polysilicon 2074 -1006 2074 -1006 0 3
rlabel polysilicon 2081 -1000 2081 -1000 0 1
rlabel polysilicon 2081 -1006 2081 -1006 0 3
rlabel polysilicon 2088 -1000 2088 -1000 0 1
rlabel polysilicon 2088 -1006 2088 -1006 0 3
rlabel polysilicon 2095 -1000 2095 -1000 0 1
rlabel polysilicon 2095 -1006 2095 -1006 0 3
rlabel polysilicon 2102 -1000 2102 -1000 0 1
rlabel polysilicon 2102 -1006 2102 -1006 0 3
rlabel polysilicon 2109 -1000 2109 -1000 0 1
rlabel polysilicon 2109 -1006 2109 -1006 0 3
rlabel polysilicon 2116 -1000 2116 -1000 0 1
rlabel polysilicon 2116 -1006 2116 -1006 0 3
rlabel polysilicon 2123 -1000 2123 -1000 0 1
rlabel polysilicon 2123 -1006 2123 -1006 0 3
rlabel polysilicon 2130 -1000 2130 -1000 0 1
rlabel polysilicon 2130 -1006 2130 -1006 0 3
rlabel polysilicon 2137 -1000 2137 -1000 0 1
rlabel polysilicon 2137 -1006 2137 -1006 0 3
rlabel polysilicon 2144 -1000 2144 -1000 0 1
rlabel polysilicon 2144 -1006 2144 -1006 0 3
rlabel polysilicon 2151 -1000 2151 -1000 0 1
rlabel polysilicon 2151 -1006 2151 -1006 0 3
rlabel polysilicon 2158 -1000 2158 -1000 0 1
rlabel polysilicon 2158 -1006 2158 -1006 0 3
rlabel polysilicon 2165 -1000 2165 -1000 0 1
rlabel polysilicon 2165 -1006 2165 -1006 0 3
rlabel polysilicon 2172 -1000 2172 -1000 0 1
rlabel polysilicon 2172 -1006 2172 -1006 0 3
rlabel polysilicon 2179 -1000 2179 -1000 0 1
rlabel polysilicon 2179 -1006 2179 -1006 0 3
rlabel polysilicon 2186 -1000 2186 -1000 0 1
rlabel polysilicon 2186 -1006 2186 -1006 0 3
rlabel polysilicon 2193 -1000 2193 -1000 0 1
rlabel polysilicon 2193 -1006 2193 -1006 0 3
rlabel polysilicon 2200 -1000 2200 -1000 0 1
rlabel polysilicon 2200 -1006 2200 -1006 0 3
rlabel polysilicon 2207 -1000 2207 -1000 0 1
rlabel polysilicon 2207 -1006 2207 -1006 0 3
rlabel polysilicon 2214 -1000 2214 -1000 0 1
rlabel polysilicon 2214 -1006 2214 -1006 0 3
rlabel polysilicon 2221 -1000 2221 -1000 0 1
rlabel polysilicon 2221 -1006 2221 -1006 0 3
rlabel polysilicon 2228 -1000 2228 -1000 0 1
rlabel polysilicon 2228 -1006 2228 -1006 0 3
rlabel polysilicon 2235 -1000 2235 -1000 0 1
rlabel polysilicon 2235 -1006 2235 -1006 0 3
rlabel polysilicon 2242 -1000 2242 -1000 0 1
rlabel polysilicon 2242 -1006 2242 -1006 0 3
rlabel polysilicon 2249 -1000 2249 -1000 0 1
rlabel polysilicon 2249 -1006 2249 -1006 0 3
rlabel polysilicon 2256 -1000 2256 -1000 0 1
rlabel polysilicon 2256 -1006 2256 -1006 0 3
rlabel polysilicon 2263 -1000 2263 -1000 0 1
rlabel polysilicon 2263 -1006 2263 -1006 0 3
rlabel polysilicon 2270 -1000 2270 -1000 0 1
rlabel polysilicon 2270 -1006 2270 -1006 0 3
rlabel polysilicon 2277 -1000 2277 -1000 0 1
rlabel polysilicon 2277 -1006 2277 -1006 0 3
rlabel polysilicon 2284 -1000 2284 -1000 0 1
rlabel polysilicon 2284 -1006 2284 -1006 0 3
rlabel polysilicon 2291 -1000 2291 -1000 0 1
rlabel polysilicon 2291 -1006 2291 -1006 0 3
rlabel polysilicon 2298 -1000 2298 -1000 0 1
rlabel polysilicon 2298 -1006 2298 -1006 0 3
rlabel polysilicon 2305 -1000 2305 -1000 0 1
rlabel polysilicon 2305 -1006 2305 -1006 0 3
rlabel polysilicon 2312 -1000 2312 -1000 0 1
rlabel polysilicon 2312 -1006 2312 -1006 0 3
rlabel polysilicon 2319 -1000 2319 -1000 0 1
rlabel polysilicon 2319 -1006 2319 -1006 0 3
rlabel polysilicon 2326 -1000 2326 -1000 0 1
rlabel polysilicon 2326 -1006 2326 -1006 0 3
rlabel polysilicon 2336 -1000 2336 -1000 0 2
rlabel polysilicon 2333 -1006 2333 -1006 0 3
rlabel polysilicon 2336 -1006 2336 -1006 0 4
rlabel polysilicon 2340 -1000 2340 -1000 0 1
rlabel polysilicon 2343 -1000 2343 -1000 0 2
rlabel polysilicon 2343 -1006 2343 -1006 0 4
rlabel polysilicon 2347 -1000 2347 -1000 0 1
rlabel polysilicon 2350 -1000 2350 -1000 0 2
rlabel polysilicon 2347 -1006 2347 -1006 0 3
rlabel polysilicon 2354 -1000 2354 -1000 0 1
rlabel polysilicon 2354 -1006 2354 -1006 0 3
rlabel polysilicon 2361 -1000 2361 -1000 0 1
rlabel polysilicon 2361 -1006 2361 -1006 0 3
rlabel polysilicon 2368 -1000 2368 -1000 0 1
rlabel polysilicon 2368 -1006 2368 -1006 0 3
rlabel polysilicon 2375 -1000 2375 -1000 0 1
rlabel polysilicon 2375 -1006 2375 -1006 0 3
rlabel polysilicon 2403 -1000 2403 -1000 0 1
rlabel polysilicon 2403 -1006 2403 -1006 0 3
rlabel polysilicon 2417 -1000 2417 -1000 0 1
rlabel polysilicon 2417 -1006 2417 -1006 0 3
rlabel polysilicon 9 -1167 9 -1167 0 1
rlabel polysilicon 9 -1173 9 -1173 0 3
rlabel polysilicon 16 -1167 16 -1167 0 1
rlabel polysilicon 16 -1173 16 -1173 0 3
rlabel polysilicon 23 -1167 23 -1167 0 1
rlabel polysilicon 23 -1173 23 -1173 0 3
rlabel polysilicon 30 -1167 30 -1167 0 1
rlabel polysilicon 30 -1173 30 -1173 0 3
rlabel polysilicon 37 -1167 37 -1167 0 1
rlabel polysilicon 37 -1173 37 -1173 0 3
rlabel polysilicon 44 -1167 44 -1167 0 1
rlabel polysilicon 44 -1173 44 -1173 0 3
rlabel polysilicon 51 -1167 51 -1167 0 1
rlabel polysilicon 51 -1173 51 -1173 0 3
rlabel polysilicon 58 -1167 58 -1167 0 1
rlabel polysilicon 58 -1173 58 -1173 0 3
rlabel polysilicon 65 -1167 65 -1167 0 1
rlabel polysilicon 65 -1173 65 -1173 0 3
rlabel polysilicon 72 -1167 72 -1167 0 1
rlabel polysilicon 72 -1173 72 -1173 0 3
rlabel polysilicon 79 -1167 79 -1167 0 1
rlabel polysilicon 79 -1173 79 -1173 0 3
rlabel polysilicon 86 -1167 86 -1167 0 1
rlabel polysilicon 89 -1167 89 -1167 0 2
rlabel polysilicon 86 -1173 86 -1173 0 3
rlabel polysilicon 89 -1173 89 -1173 0 4
rlabel polysilicon 93 -1167 93 -1167 0 1
rlabel polysilicon 93 -1173 93 -1173 0 3
rlabel polysilicon 100 -1167 100 -1167 0 1
rlabel polysilicon 100 -1173 100 -1173 0 3
rlabel polysilicon 107 -1167 107 -1167 0 1
rlabel polysilicon 110 -1167 110 -1167 0 2
rlabel polysilicon 110 -1173 110 -1173 0 4
rlabel polysilicon 114 -1167 114 -1167 0 1
rlabel polysilicon 117 -1167 117 -1167 0 2
rlabel polysilicon 114 -1173 114 -1173 0 3
rlabel polysilicon 121 -1167 121 -1167 0 1
rlabel polysilicon 121 -1173 121 -1173 0 3
rlabel polysilicon 128 -1167 128 -1167 0 1
rlabel polysilicon 128 -1173 128 -1173 0 3
rlabel polysilicon 135 -1167 135 -1167 0 1
rlabel polysilicon 138 -1167 138 -1167 0 2
rlabel polysilicon 135 -1173 135 -1173 0 3
rlabel polysilicon 138 -1173 138 -1173 0 4
rlabel polysilicon 142 -1167 142 -1167 0 1
rlabel polysilicon 145 -1167 145 -1167 0 2
rlabel polysilicon 142 -1173 142 -1173 0 3
rlabel polysilicon 145 -1173 145 -1173 0 4
rlabel polysilicon 149 -1167 149 -1167 0 1
rlabel polysilicon 149 -1173 149 -1173 0 3
rlabel polysilicon 156 -1167 156 -1167 0 1
rlabel polysilicon 156 -1173 156 -1173 0 3
rlabel polysilicon 163 -1167 163 -1167 0 1
rlabel polysilicon 163 -1173 163 -1173 0 3
rlabel polysilicon 170 -1167 170 -1167 0 1
rlabel polysilicon 170 -1173 170 -1173 0 3
rlabel polysilicon 177 -1167 177 -1167 0 1
rlabel polysilicon 177 -1173 177 -1173 0 3
rlabel polysilicon 184 -1167 184 -1167 0 1
rlabel polysilicon 184 -1173 184 -1173 0 3
rlabel polysilicon 191 -1167 191 -1167 0 1
rlabel polysilicon 191 -1173 191 -1173 0 3
rlabel polysilicon 198 -1167 198 -1167 0 1
rlabel polysilicon 198 -1173 198 -1173 0 3
rlabel polysilicon 205 -1167 205 -1167 0 1
rlabel polysilicon 205 -1173 205 -1173 0 3
rlabel polysilicon 212 -1167 212 -1167 0 1
rlabel polysilicon 212 -1173 212 -1173 0 3
rlabel polysilicon 219 -1167 219 -1167 0 1
rlabel polysilicon 219 -1173 219 -1173 0 3
rlabel polysilicon 226 -1167 226 -1167 0 1
rlabel polysilicon 226 -1173 226 -1173 0 3
rlabel polysilicon 233 -1167 233 -1167 0 1
rlabel polysilicon 233 -1173 233 -1173 0 3
rlabel polysilicon 240 -1167 240 -1167 0 1
rlabel polysilicon 240 -1173 240 -1173 0 3
rlabel polysilicon 243 -1173 243 -1173 0 4
rlabel polysilicon 247 -1167 247 -1167 0 1
rlabel polysilicon 247 -1173 247 -1173 0 3
rlabel polysilicon 254 -1167 254 -1167 0 1
rlabel polysilicon 254 -1173 254 -1173 0 3
rlabel polysilicon 261 -1167 261 -1167 0 1
rlabel polysilicon 261 -1173 261 -1173 0 3
rlabel polysilicon 268 -1167 268 -1167 0 1
rlabel polysilicon 268 -1173 268 -1173 0 3
rlabel polysilicon 275 -1167 275 -1167 0 1
rlabel polysilicon 275 -1173 275 -1173 0 3
rlabel polysilicon 282 -1167 282 -1167 0 1
rlabel polysilicon 282 -1173 282 -1173 0 3
rlabel polysilicon 289 -1167 289 -1167 0 1
rlabel polysilicon 289 -1173 289 -1173 0 3
rlabel polysilicon 296 -1167 296 -1167 0 1
rlabel polysilicon 296 -1173 296 -1173 0 3
rlabel polysilicon 303 -1167 303 -1167 0 1
rlabel polysilicon 303 -1173 303 -1173 0 3
rlabel polysilicon 310 -1167 310 -1167 0 1
rlabel polysilicon 310 -1173 310 -1173 0 3
rlabel polysilicon 317 -1167 317 -1167 0 1
rlabel polysilicon 317 -1173 317 -1173 0 3
rlabel polysilicon 324 -1167 324 -1167 0 1
rlabel polysilicon 324 -1173 324 -1173 0 3
rlabel polysilicon 331 -1167 331 -1167 0 1
rlabel polysilicon 331 -1173 331 -1173 0 3
rlabel polysilicon 338 -1167 338 -1167 0 1
rlabel polysilicon 338 -1173 338 -1173 0 3
rlabel polysilicon 345 -1167 345 -1167 0 1
rlabel polysilicon 345 -1173 345 -1173 0 3
rlabel polysilicon 352 -1167 352 -1167 0 1
rlabel polysilicon 352 -1173 352 -1173 0 3
rlabel polysilicon 359 -1167 359 -1167 0 1
rlabel polysilicon 359 -1173 359 -1173 0 3
rlabel polysilicon 366 -1167 366 -1167 0 1
rlabel polysilicon 366 -1173 366 -1173 0 3
rlabel polysilicon 373 -1167 373 -1167 0 1
rlabel polysilicon 373 -1173 373 -1173 0 3
rlabel polysilicon 380 -1167 380 -1167 0 1
rlabel polysilicon 380 -1173 380 -1173 0 3
rlabel polysilicon 387 -1167 387 -1167 0 1
rlabel polysilicon 387 -1173 387 -1173 0 3
rlabel polysilicon 394 -1167 394 -1167 0 1
rlabel polysilicon 394 -1173 394 -1173 0 3
rlabel polysilicon 401 -1167 401 -1167 0 1
rlabel polysilicon 401 -1173 401 -1173 0 3
rlabel polysilicon 408 -1167 408 -1167 0 1
rlabel polysilicon 408 -1173 408 -1173 0 3
rlabel polysilicon 415 -1167 415 -1167 0 1
rlabel polysilicon 415 -1173 415 -1173 0 3
rlabel polysilicon 422 -1167 422 -1167 0 1
rlabel polysilicon 425 -1167 425 -1167 0 2
rlabel polysilicon 422 -1173 422 -1173 0 3
rlabel polysilicon 429 -1167 429 -1167 0 1
rlabel polysilicon 432 -1167 432 -1167 0 2
rlabel polysilicon 432 -1173 432 -1173 0 4
rlabel polysilicon 436 -1167 436 -1167 0 1
rlabel polysilicon 436 -1173 436 -1173 0 3
rlabel polysilicon 443 -1167 443 -1167 0 1
rlabel polysilicon 443 -1173 443 -1173 0 3
rlabel polysilicon 450 -1167 450 -1167 0 1
rlabel polysilicon 450 -1173 450 -1173 0 3
rlabel polysilicon 457 -1167 457 -1167 0 1
rlabel polysilicon 457 -1173 457 -1173 0 3
rlabel polysilicon 464 -1167 464 -1167 0 1
rlabel polysilicon 464 -1173 464 -1173 0 3
rlabel polysilicon 471 -1167 471 -1167 0 1
rlabel polysilicon 471 -1173 471 -1173 0 3
rlabel polysilicon 478 -1167 478 -1167 0 1
rlabel polysilicon 478 -1173 478 -1173 0 3
rlabel polysilicon 485 -1167 485 -1167 0 1
rlabel polysilicon 485 -1173 485 -1173 0 3
rlabel polysilicon 492 -1167 492 -1167 0 1
rlabel polysilicon 492 -1173 492 -1173 0 3
rlabel polysilicon 499 -1167 499 -1167 0 1
rlabel polysilicon 499 -1173 499 -1173 0 3
rlabel polysilicon 506 -1167 506 -1167 0 1
rlabel polysilicon 506 -1173 506 -1173 0 3
rlabel polysilicon 509 -1173 509 -1173 0 4
rlabel polysilicon 513 -1167 513 -1167 0 1
rlabel polysilicon 513 -1173 513 -1173 0 3
rlabel polysilicon 520 -1167 520 -1167 0 1
rlabel polysilicon 520 -1173 520 -1173 0 3
rlabel polysilicon 527 -1167 527 -1167 0 1
rlabel polysilicon 527 -1173 527 -1173 0 3
rlabel polysilicon 534 -1167 534 -1167 0 1
rlabel polysilicon 534 -1173 534 -1173 0 3
rlabel polysilicon 541 -1167 541 -1167 0 1
rlabel polysilicon 541 -1173 541 -1173 0 3
rlabel polysilicon 548 -1167 548 -1167 0 1
rlabel polysilicon 548 -1173 548 -1173 0 3
rlabel polysilicon 555 -1167 555 -1167 0 1
rlabel polysilicon 555 -1173 555 -1173 0 3
rlabel polysilicon 562 -1167 562 -1167 0 1
rlabel polysilicon 562 -1173 562 -1173 0 3
rlabel polysilicon 569 -1167 569 -1167 0 1
rlabel polysilicon 569 -1173 569 -1173 0 3
rlabel polysilicon 576 -1167 576 -1167 0 1
rlabel polysilicon 576 -1173 576 -1173 0 3
rlabel polysilicon 583 -1167 583 -1167 0 1
rlabel polysilicon 583 -1173 583 -1173 0 3
rlabel polysilicon 590 -1167 590 -1167 0 1
rlabel polysilicon 593 -1167 593 -1167 0 2
rlabel polysilicon 590 -1173 590 -1173 0 3
rlabel polysilicon 597 -1167 597 -1167 0 1
rlabel polysilicon 597 -1173 597 -1173 0 3
rlabel polysilicon 604 -1167 604 -1167 0 1
rlabel polysilicon 607 -1167 607 -1167 0 2
rlabel polysilicon 607 -1173 607 -1173 0 4
rlabel polysilicon 611 -1167 611 -1167 0 1
rlabel polysilicon 611 -1173 611 -1173 0 3
rlabel polysilicon 618 -1167 618 -1167 0 1
rlabel polysilicon 618 -1173 618 -1173 0 3
rlabel polysilicon 625 -1167 625 -1167 0 1
rlabel polysilicon 625 -1173 625 -1173 0 3
rlabel polysilicon 632 -1167 632 -1167 0 1
rlabel polysilicon 632 -1173 632 -1173 0 3
rlabel polysilicon 639 -1167 639 -1167 0 1
rlabel polysilicon 639 -1173 639 -1173 0 3
rlabel polysilicon 646 -1167 646 -1167 0 1
rlabel polysilicon 646 -1173 646 -1173 0 3
rlabel polysilicon 656 -1167 656 -1167 0 2
rlabel polysilicon 653 -1173 653 -1173 0 3
rlabel polysilicon 656 -1173 656 -1173 0 4
rlabel polysilicon 660 -1167 660 -1167 0 1
rlabel polysilicon 660 -1173 660 -1173 0 3
rlabel polysilicon 667 -1167 667 -1167 0 1
rlabel polysilicon 667 -1173 667 -1173 0 3
rlabel polysilicon 674 -1167 674 -1167 0 1
rlabel polysilicon 674 -1173 674 -1173 0 3
rlabel polysilicon 681 -1167 681 -1167 0 1
rlabel polysilicon 681 -1173 681 -1173 0 3
rlabel polysilicon 688 -1167 688 -1167 0 1
rlabel polysilicon 688 -1173 688 -1173 0 3
rlabel polysilicon 695 -1167 695 -1167 0 1
rlabel polysilicon 695 -1173 695 -1173 0 3
rlabel polysilicon 702 -1167 702 -1167 0 1
rlabel polysilicon 702 -1173 702 -1173 0 3
rlabel polysilicon 709 -1167 709 -1167 0 1
rlabel polysilicon 709 -1173 709 -1173 0 3
rlabel polysilicon 716 -1167 716 -1167 0 1
rlabel polysilicon 716 -1173 716 -1173 0 3
rlabel polysilicon 723 -1167 723 -1167 0 1
rlabel polysilicon 723 -1173 723 -1173 0 3
rlabel polysilicon 730 -1167 730 -1167 0 1
rlabel polysilicon 733 -1167 733 -1167 0 2
rlabel polysilicon 730 -1173 730 -1173 0 3
rlabel polysilicon 737 -1167 737 -1167 0 1
rlabel polysilicon 737 -1173 737 -1173 0 3
rlabel polysilicon 744 -1167 744 -1167 0 1
rlabel polysilicon 744 -1173 744 -1173 0 3
rlabel polysilicon 751 -1167 751 -1167 0 1
rlabel polysilicon 751 -1173 751 -1173 0 3
rlabel polysilicon 761 -1167 761 -1167 0 2
rlabel polysilicon 758 -1173 758 -1173 0 3
rlabel polysilicon 761 -1173 761 -1173 0 4
rlabel polysilicon 765 -1167 765 -1167 0 1
rlabel polysilicon 765 -1173 765 -1173 0 3
rlabel polysilicon 772 -1167 772 -1167 0 1
rlabel polysilicon 775 -1167 775 -1167 0 2
rlabel polysilicon 772 -1173 772 -1173 0 3
rlabel polysilicon 779 -1167 779 -1167 0 1
rlabel polysilicon 779 -1173 779 -1173 0 3
rlabel polysilicon 786 -1167 786 -1167 0 1
rlabel polysilicon 786 -1173 786 -1173 0 3
rlabel polysilicon 793 -1167 793 -1167 0 1
rlabel polysilicon 793 -1173 793 -1173 0 3
rlabel polysilicon 800 -1167 800 -1167 0 1
rlabel polysilicon 800 -1173 800 -1173 0 3
rlabel polysilicon 807 -1167 807 -1167 0 1
rlabel polysilicon 807 -1173 807 -1173 0 3
rlabel polysilicon 814 -1167 814 -1167 0 1
rlabel polysilicon 814 -1173 814 -1173 0 3
rlabel polysilicon 821 -1167 821 -1167 0 1
rlabel polysilicon 824 -1167 824 -1167 0 2
rlabel polysilicon 821 -1173 821 -1173 0 3
rlabel polysilicon 824 -1173 824 -1173 0 4
rlabel polysilicon 828 -1167 828 -1167 0 1
rlabel polysilicon 828 -1173 828 -1173 0 3
rlabel polysilicon 835 -1167 835 -1167 0 1
rlabel polysilicon 835 -1173 835 -1173 0 3
rlabel polysilicon 842 -1167 842 -1167 0 1
rlabel polysilicon 842 -1173 842 -1173 0 3
rlabel polysilicon 849 -1167 849 -1167 0 1
rlabel polysilicon 852 -1173 852 -1173 0 4
rlabel polysilicon 856 -1167 856 -1167 0 1
rlabel polysilicon 856 -1173 856 -1173 0 3
rlabel polysilicon 863 -1167 863 -1167 0 1
rlabel polysilicon 866 -1167 866 -1167 0 2
rlabel polysilicon 866 -1173 866 -1173 0 4
rlabel polysilicon 870 -1167 870 -1167 0 1
rlabel polysilicon 877 -1167 877 -1167 0 1
rlabel polysilicon 880 -1167 880 -1167 0 2
rlabel polysilicon 877 -1173 877 -1173 0 3
rlabel polysilicon 880 -1173 880 -1173 0 4
rlabel polysilicon 884 -1167 884 -1167 0 1
rlabel polysilicon 884 -1173 884 -1173 0 3
rlabel polysilicon 891 -1167 891 -1167 0 1
rlabel polysilicon 891 -1173 891 -1173 0 3
rlabel polysilicon 898 -1167 898 -1167 0 1
rlabel polysilicon 898 -1173 898 -1173 0 3
rlabel polysilicon 905 -1167 905 -1167 0 1
rlabel polysilicon 908 -1173 908 -1173 0 4
rlabel polysilicon 912 -1167 912 -1167 0 1
rlabel polysilicon 912 -1173 912 -1173 0 3
rlabel polysilicon 919 -1167 919 -1167 0 1
rlabel polysilicon 919 -1173 919 -1173 0 3
rlabel polysilicon 926 -1167 926 -1167 0 1
rlabel polysilicon 926 -1173 926 -1173 0 3
rlabel polysilicon 933 -1167 933 -1167 0 1
rlabel polysilicon 933 -1173 933 -1173 0 3
rlabel polysilicon 940 -1167 940 -1167 0 1
rlabel polysilicon 940 -1173 940 -1173 0 3
rlabel polysilicon 947 -1167 947 -1167 0 1
rlabel polysilicon 950 -1167 950 -1167 0 2
rlabel polysilicon 947 -1173 947 -1173 0 3
rlabel polysilicon 950 -1173 950 -1173 0 4
rlabel polysilicon 957 -1167 957 -1167 0 2
rlabel polysilicon 954 -1173 954 -1173 0 3
rlabel polysilicon 961 -1167 961 -1167 0 1
rlabel polysilicon 964 -1167 964 -1167 0 2
rlabel polysilicon 961 -1173 961 -1173 0 3
rlabel polysilicon 964 -1173 964 -1173 0 4
rlabel polysilicon 968 -1167 968 -1167 0 1
rlabel polysilicon 968 -1173 968 -1173 0 3
rlabel polysilicon 975 -1167 975 -1167 0 1
rlabel polysilicon 975 -1173 975 -1173 0 3
rlabel polysilicon 982 -1167 982 -1167 0 1
rlabel polysilicon 982 -1173 982 -1173 0 3
rlabel polysilicon 989 -1167 989 -1167 0 1
rlabel polysilicon 989 -1173 989 -1173 0 3
rlabel polysilicon 996 -1167 996 -1167 0 1
rlabel polysilicon 996 -1173 996 -1173 0 3
rlabel polysilicon 1003 -1167 1003 -1167 0 1
rlabel polysilicon 1006 -1167 1006 -1167 0 2
rlabel polysilicon 1003 -1173 1003 -1173 0 3
rlabel polysilicon 1006 -1173 1006 -1173 0 4
rlabel polysilicon 1010 -1167 1010 -1167 0 1
rlabel polysilicon 1010 -1173 1010 -1173 0 3
rlabel polysilicon 1017 -1167 1017 -1167 0 1
rlabel polysilicon 1017 -1173 1017 -1173 0 3
rlabel polysilicon 1024 -1167 1024 -1167 0 1
rlabel polysilicon 1024 -1173 1024 -1173 0 3
rlabel polysilicon 1031 -1167 1031 -1167 0 1
rlabel polysilicon 1031 -1173 1031 -1173 0 3
rlabel polysilicon 1038 -1167 1038 -1167 0 1
rlabel polysilicon 1038 -1173 1038 -1173 0 3
rlabel polysilicon 1045 -1167 1045 -1167 0 1
rlabel polysilicon 1045 -1173 1045 -1173 0 3
rlabel polysilicon 1048 -1173 1048 -1173 0 4
rlabel polysilicon 1052 -1167 1052 -1167 0 1
rlabel polysilicon 1052 -1173 1052 -1173 0 3
rlabel polysilicon 1059 -1167 1059 -1167 0 1
rlabel polysilicon 1059 -1173 1059 -1173 0 3
rlabel polysilicon 1066 -1167 1066 -1167 0 1
rlabel polysilicon 1066 -1173 1066 -1173 0 3
rlabel polysilicon 1073 -1167 1073 -1167 0 1
rlabel polysilicon 1073 -1173 1073 -1173 0 3
rlabel polysilicon 1080 -1167 1080 -1167 0 1
rlabel polysilicon 1080 -1173 1080 -1173 0 3
rlabel polysilicon 1087 -1167 1087 -1167 0 1
rlabel polysilicon 1087 -1173 1087 -1173 0 3
rlabel polysilicon 1094 -1167 1094 -1167 0 1
rlabel polysilicon 1094 -1173 1094 -1173 0 3
rlabel polysilicon 1101 -1167 1101 -1167 0 1
rlabel polysilicon 1101 -1173 1101 -1173 0 3
rlabel polysilicon 1108 -1167 1108 -1167 0 1
rlabel polysilicon 1108 -1173 1108 -1173 0 3
rlabel polysilicon 1115 -1167 1115 -1167 0 1
rlabel polysilicon 1115 -1173 1115 -1173 0 3
rlabel polysilicon 1122 -1167 1122 -1167 0 1
rlabel polysilicon 1122 -1173 1122 -1173 0 3
rlabel polysilicon 1129 -1167 1129 -1167 0 1
rlabel polysilicon 1129 -1173 1129 -1173 0 3
rlabel polysilicon 1136 -1167 1136 -1167 0 1
rlabel polysilicon 1136 -1173 1136 -1173 0 3
rlabel polysilicon 1143 -1167 1143 -1167 0 1
rlabel polysilicon 1143 -1173 1143 -1173 0 3
rlabel polysilicon 1150 -1167 1150 -1167 0 1
rlabel polysilicon 1150 -1173 1150 -1173 0 3
rlabel polysilicon 1157 -1167 1157 -1167 0 1
rlabel polysilicon 1160 -1167 1160 -1167 0 2
rlabel polysilicon 1157 -1173 1157 -1173 0 3
rlabel polysilicon 1160 -1173 1160 -1173 0 4
rlabel polysilicon 1164 -1167 1164 -1167 0 1
rlabel polysilicon 1167 -1167 1167 -1167 0 2
rlabel polysilicon 1164 -1173 1164 -1173 0 3
rlabel polysilicon 1167 -1173 1167 -1173 0 4
rlabel polysilicon 1171 -1167 1171 -1167 0 1
rlabel polysilicon 1171 -1173 1171 -1173 0 3
rlabel polysilicon 1178 -1167 1178 -1167 0 1
rlabel polysilicon 1181 -1167 1181 -1167 0 2
rlabel polysilicon 1178 -1173 1178 -1173 0 3
rlabel polysilicon 1181 -1173 1181 -1173 0 4
rlabel polysilicon 1185 -1167 1185 -1167 0 1
rlabel polysilicon 1185 -1173 1185 -1173 0 3
rlabel polysilicon 1192 -1167 1192 -1167 0 1
rlabel polysilicon 1192 -1173 1192 -1173 0 3
rlabel polysilicon 1199 -1167 1199 -1167 0 1
rlabel polysilicon 1202 -1167 1202 -1167 0 2
rlabel polysilicon 1199 -1173 1199 -1173 0 3
rlabel polysilicon 1202 -1173 1202 -1173 0 4
rlabel polysilicon 1206 -1167 1206 -1167 0 1
rlabel polysilicon 1206 -1173 1206 -1173 0 3
rlabel polysilicon 1213 -1167 1213 -1167 0 1
rlabel polysilicon 1213 -1173 1213 -1173 0 3
rlabel polysilicon 1220 -1167 1220 -1167 0 1
rlabel polysilicon 1223 -1167 1223 -1167 0 2
rlabel polysilicon 1220 -1173 1220 -1173 0 3
rlabel polysilicon 1227 -1167 1227 -1167 0 1
rlabel polysilicon 1227 -1173 1227 -1173 0 3
rlabel polysilicon 1234 -1167 1234 -1167 0 1
rlabel polysilicon 1237 -1167 1237 -1167 0 2
rlabel polysilicon 1234 -1173 1234 -1173 0 3
rlabel polysilicon 1237 -1173 1237 -1173 0 4
rlabel polysilicon 1241 -1167 1241 -1167 0 1
rlabel polysilicon 1241 -1173 1241 -1173 0 3
rlabel polysilicon 1248 -1167 1248 -1167 0 1
rlabel polysilicon 1248 -1173 1248 -1173 0 3
rlabel polysilicon 1255 -1167 1255 -1167 0 1
rlabel polysilicon 1255 -1173 1255 -1173 0 3
rlabel polysilicon 1262 -1167 1262 -1167 0 1
rlabel polysilicon 1262 -1173 1262 -1173 0 3
rlabel polysilicon 1269 -1167 1269 -1167 0 1
rlabel polysilicon 1269 -1173 1269 -1173 0 3
rlabel polysilicon 1276 -1167 1276 -1167 0 1
rlabel polysilicon 1276 -1173 1276 -1173 0 3
rlabel polysilicon 1283 -1167 1283 -1167 0 1
rlabel polysilicon 1283 -1173 1283 -1173 0 3
rlabel polysilicon 1290 -1167 1290 -1167 0 1
rlabel polysilicon 1290 -1173 1290 -1173 0 3
rlabel polysilicon 1297 -1167 1297 -1167 0 1
rlabel polysilicon 1297 -1173 1297 -1173 0 3
rlabel polysilicon 1304 -1167 1304 -1167 0 1
rlabel polysilicon 1307 -1167 1307 -1167 0 2
rlabel polysilicon 1304 -1173 1304 -1173 0 3
rlabel polysilicon 1307 -1173 1307 -1173 0 4
rlabel polysilicon 1311 -1167 1311 -1167 0 1
rlabel polysilicon 1311 -1173 1311 -1173 0 3
rlabel polysilicon 1318 -1167 1318 -1167 0 1
rlabel polysilicon 1318 -1173 1318 -1173 0 3
rlabel polysilicon 1325 -1167 1325 -1167 0 1
rlabel polysilicon 1325 -1173 1325 -1173 0 3
rlabel polysilicon 1332 -1167 1332 -1167 0 1
rlabel polysilicon 1335 -1167 1335 -1167 0 2
rlabel polysilicon 1332 -1173 1332 -1173 0 3
rlabel polysilicon 1335 -1173 1335 -1173 0 4
rlabel polysilicon 1339 -1167 1339 -1167 0 1
rlabel polysilicon 1339 -1173 1339 -1173 0 3
rlabel polysilicon 1346 -1167 1346 -1167 0 1
rlabel polysilicon 1346 -1173 1346 -1173 0 3
rlabel polysilicon 1353 -1167 1353 -1167 0 1
rlabel polysilicon 1353 -1173 1353 -1173 0 3
rlabel polysilicon 1360 -1167 1360 -1167 0 1
rlabel polysilicon 1360 -1173 1360 -1173 0 3
rlabel polysilicon 1367 -1167 1367 -1167 0 1
rlabel polysilicon 1367 -1173 1367 -1173 0 3
rlabel polysilicon 1374 -1167 1374 -1167 0 1
rlabel polysilicon 1374 -1173 1374 -1173 0 3
rlabel polysilicon 1381 -1167 1381 -1167 0 1
rlabel polysilicon 1381 -1173 1381 -1173 0 3
rlabel polysilicon 1388 -1167 1388 -1167 0 1
rlabel polysilicon 1388 -1173 1388 -1173 0 3
rlabel polysilicon 1391 -1173 1391 -1173 0 4
rlabel polysilicon 1395 -1167 1395 -1167 0 1
rlabel polysilicon 1395 -1173 1395 -1173 0 3
rlabel polysilicon 1402 -1167 1402 -1167 0 1
rlabel polysilicon 1402 -1173 1402 -1173 0 3
rlabel polysilicon 1409 -1167 1409 -1167 0 1
rlabel polysilicon 1409 -1173 1409 -1173 0 3
rlabel polysilicon 1416 -1167 1416 -1167 0 1
rlabel polysilicon 1416 -1173 1416 -1173 0 3
rlabel polysilicon 1423 -1167 1423 -1167 0 1
rlabel polysilicon 1423 -1173 1423 -1173 0 3
rlabel polysilicon 1430 -1167 1430 -1167 0 1
rlabel polysilicon 1430 -1173 1430 -1173 0 3
rlabel polysilicon 1437 -1167 1437 -1167 0 1
rlabel polysilicon 1437 -1173 1437 -1173 0 3
rlabel polysilicon 1447 -1167 1447 -1167 0 2
rlabel polysilicon 1444 -1173 1444 -1173 0 3
rlabel polysilicon 1447 -1173 1447 -1173 0 4
rlabel polysilicon 1451 -1167 1451 -1167 0 1
rlabel polysilicon 1451 -1173 1451 -1173 0 3
rlabel polysilicon 1458 -1167 1458 -1167 0 1
rlabel polysilicon 1458 -1173 1458 -1173 0 3
rlabel polysilicon 1465 -1167 1465 -1167 0 1
rlabel polysilicon 1465 -1173 1465 -1173 0 3
rlabel polysilicon 1472 -1167 1472 -1167 0 1
rlabel polysilicon 1472 -1173 1472 -1173 0 3
rlabel polysilicon 1479 -1167 1479 -1167 0 1
rlabel polysilicon 1479 -1173 1479 -1173 0 3
rlabel polysilicon 1486 -1167 1486 -1167 0 1
rlabel polysilicon 1486 -1173 1486 -1173 0 3
rlabel polysilicon 1493 -1167 1493 -1167 0 1
rlabel polysilicon 1493 -1173 1493 -1173 0 3
rlabel polysilicon 1500 -1167 1500 -1167 0 1
rlabel polysilicon 1500 -1173 1500 -1173 0 3
rlabel polysilicon 1507 -1167 1507 -1167 0 1
rlabel polysilicon 1507 -1173 1507 -1173 0 3
rlabel polysilicon 1514 -1167 1514 -1167 0 1
rlabel polysilicon 1514 -1173 1514 -1173 0 3
rlabel polysilicon 1521 -1167 1521 -1167 0 1
rlabel polysilicon 1521 -1173 1521 -1173 0 3
rlabel polysilicon 1528 -1167 1528 -1167 0 1
rlabel polysilicon 1528 -1173 1528 -1173 0 3
rlabel polysilicon 1535 -1167 1535 -1167 0 1
rlabel polysilicon 1535 -1173 1535 -1173 0 3
rlabel polysilicon 1542 -1167 1542 -1167 0 1
rlabel polysilicon 1542 -1173 1542 -1173 0 3
rlabel polysilicon 1549 -1167 1549 -1167 0 1
rlabel polysilicon 1549 -1173 1549 -1173 0 3
rlabel polysilicon 1552 -1173 1552 -1173 0 4
rlabel polysilicon 1556 -1167 1556 -1167 0 1
rlabel polysilicon 1556 -1173 1556 -1173 0 3
rlabel polysilicon 1563 -1167 1563 -1167 0 1
rlabel polysilicon 1563 -1173 1563 -1173 0 3
rlabel polysilicon 1570 -1167 1570 -1167 0 1
rlabel polysilicon 1570 -1173 1570 -1173 0 3
rlabel polysilicon 1577 -1167 1577 -1167 0 1
rlabel polysilicon 1577 -1173 1577 -1173 0 3
rlabel polysilicon 1584 -1167 1584 -1167 0 1
rlabel polysilicon 1584 -1173 1584 -1173 0 3
rlabel polysilicon 1591 -1167 1591 -1167 0 1
rlabel polysilicon 1591 -1173 1591 -1173 0 3
rlabel polysilicon 1598 -1167 1598 -1167 0 1
rlabel polysilicon 1598 -1173 1598 -1173 0 3
rlabel polysilicon 1605 -1167 1605 -1167 0 1
rlabel polysilicon 1605 -1173 1605 -1173 0 3
rlabel polysilicon 1612 -1167 1612 -1167 0 1
rlabel polysilicon 1612 -1173 1612 -1173 0 3
rlabel polysilicon 1619 -1167 1619 -1167 0 1
rlabel polysilicon 1619 -1173 1619 -1173 0 3
rlabel polysilicon 1626 -1167 1626 -1167 0 1
rlabel polysilicon 1626 -1173 1626 -1173 0 3
rlabel polysilicon 1633 -1167 1633 -1167 0 1
rlabel polysilicon 1633 -1173 1633 -1173 0 3
rlabel polysilicon 1640 -1167 1640 -1167 0 1
rlabel polysilicon 1640 -1173 1640 -1173 0 3
rlabel polysilicon 1647 -1167 1647 -1167 0 1
rlabel polysilicon 1647 -1173 1647 -1173 0 3
rlabel polysilicon 1654 -1167 1654 -1167 0 1
rlabel polysilicon 1654 -1173 1654 -1173 0 3
rlabel polysilicon 1661 -1167 1661 -1167 0 1
rlabel polysilicon 1661 -1173 1661 -1173 0 3
rlabel polysilicon 1668 -1167 1668 -1167 0 1
rlabel polysilicon 1668 -1173 1668 -1173 0 3
rlabel polysilicon 1675 -1167 1675 -1167 0 1
rlabel polysilicon 1675 -1173 1675 -1173 0 3
rlabel polysilicon 1682 -1167 1682 -1167 0 1
rlabel polysilicon 1682 -1173 1682 -1173 0 3
rlabel polysilicon 1689 -1167 1689 -1167 0 1
rlabel polysilicon 1689 -1173 1689 -1173 0 3
rlabel polysilicon 1696 -1167 1696 -1167 0 1
rlabel polysilicon 1696 -1173 1696 -1173 0 3
rlabel polysilicon 1703 -1167 1703 -1167 0 1
rlabel polysilicon 1703 -1173 1703 -1173 0 3
rlabel polysilicon 1710 -1167 1710 -1167 0 1
rlabel polysilicon 1710 -1173 1710 -1173 0 3
rlabel polysilicon 1717 -1167 1717 -1167 0 1
rlabel polysilicon 1717 -1173 1717 -1173 0 3
rlabel polysilicon 1724 -1167 1724 -1167 0 1
rlabel polysilicon 1724 -1173 1724 -1173 0 3
rlabel polysilicon 1731 -1167 1731 -1167 0 1
rlabel polysilicon 1731 -1173 1731 -1173 0 3
rlabel polysilicon 1741 -1167 1741 -1167 0 2
rlabel polysilicon 1738 -1173 1738 -1173 0 3
rlabel polysilicon 1741 -1173 1741 -1173 0 4
rlabel polysilicon 1745 -1167 1745 -1167 0 1
rlabel polysilicon 1745 -1173 1745 -1173 0 3
rlabel polysilicon 1752 -1167 1752 -1167 0 1
rlabel polysilicon 1752 -1173 1752 -1173 0 3
rlabel polysilicon 1759 -1167 1759 -1167 0 1
rlabel polysilicon 1759 -1173 1759 -1173 0 3
rlabel polysilicon 1766 -1167 1766 -1167 0 1
rlabel polysilicon 1766 -1173 1766 -1173 0 3
rlabel polysilicon 1773 -1167 1773 -1167 0 1
rlabel polysilicon 1773 -1173 1773 -1173 0 3
rlabel polysilicon 1780 -1167 1780 -1167 0 1
rlabel polysilicon 1780 -1173 1780 -1173 0 3
rlabel polysilicon 1787 -1167 1787 -1167 0 1
rlabel polysilicon 1787 -1173 1787 -1173 0 3
rlabel polysilicon 1794 -1167 1794 -1167 0 1
rlabel polysilicon 1794 -1173 1794 -1173 0 3
rlabel polysilicon 1801 -1167 1801 -1167 0 1
rlabel polysilicon 1801 -1173 1801 -1173 0 3
rlabel polysilicon 1808 -1167 1808 -1167 0 1
rlabel polysilicon 1808 -1173 1808 -1173 0 3
rlabel polysilicon 1815 -1167 1815 -1167 0 1
rlabel polysilicon 1815 -1173 1815 -1173 0 3
rlabel polysilicon 1822 -1167 1822 -1167 0 1
rlabel polysilicon 1822 -1173 1822 -1173 0 3
rlabel polysilicon 1829 -1167 1829 -1167 0 1
rlabel polysilicon 1829 -1173 1829 -1173 0 3
rlabel polysilicon 1836 -1167 1836 -1167 0 1
rlabel polysilicon 1836 -1173 1836 -1173 0 3
rlabel polysilicon 1843 -1167 1843 -1167 0 1
rlabel polysilicon 1843 -1173 1843 -1173 0 3
rlabel polysilicon 1850 -1167 1850 -1167 0 1
rlabel polysilicon 1850 -1173 1850 -1173 0 3
rlabel polysilicon 1857 -1167 1857 -1167 0 1
rlabel polysilicon 1857 -1173 1857 -1173 0 3
rlabel polysilicon 1864 -1167 1864 -1167 0 1
rlabel polysilicon 1864 -1173 1864 -1173 0 3
rlabel polysilicon 1871 -1167 1871 -1167 0 1
rlabel polysilicon 1871 -1173 1871 -1173 0 3
rlabel polysilicon 1878 -1167 1878 -1167 0 1
rlabel polysilicon 1878 -1173 1878 -1173 0 3
rlabel polysilicon 1885 -1167 1885 -1167 0 1
rlabel polysilicon 1885 -1173 1885 -1173 0 3
rlabel polysilicon 1892 -1167 1892 -1167 0 1
rlabel polysilicon 1892 -1173 1892 -1173 0 3
rlabel polysilicon 1899 -1167 1899 -1167 0 1
rlabel polysilicon 1899 -1173 1899 -1173 0 3
rlabel polysilicon 1906 -1167 1906 -1167 0 1
rlabel polysilicon 1906 -1173 1906 -1173 0 3
rlabel polysilicon 1913 -1167 1913 -1167 0 1
rlabel polysilicon 1913 -1173 1913 -1173 0 3
rlabel polysilicon 1920 -1167 1920 -1167 0 1
rlabel polysilicon 1920 -1173 1920 -1173 0 3
rlabel polysilicon 1927 -1167 1927 -1167 0 1
rlabel polysilicon 1927 -1173 1927 -1173 0 3
rlabel polysilicon 1934 -1167 1934 -1167 0 1
rlabel polysilicon 1934 -1173 1934 -1173 0 3
rlabel polysilicon 1941 -1167 1941 -1167 0 1
rlabel polysilicon 1941 -1173 1941 -1173 0 3
rlabel polysilicon 1948 -1167 1948 -1167 0 1
rlabel polysilicon 1948 -1173 1948 -1173 0 3
rlabel polysilicon 1955 -1167 1955 -1167 0 1
rlabel polysilicon 1955 -1173 1955 -1173 0 3
rlabel polysilicon 1962 -1167 1962 -1167 0 1
rlabel polysilicon 1962 -1173 1962 -1173 0 3
rlabel polysilicon 1969 -1167 1969 -1167 0 1
rlabel polysilicon 1969 -1173 1969 -1173 0 3
rlabel polysilicon 1976 -1167 1976 -1167 0 1
rlabel polysilicon 1976 -1173 1976 -1173 0 3
rlabel polysilicon 1983 -1167 1983 -1167 0 1
rlabel polysilicon 1983 -1173 1983 -1173 0 3
rlabel polysilicon 1990 -1167 1990 -1167 0 1
rlabel polysilicon 1990 -1173 1990 -1173 0 3
rlabel polysilicon 1997 -1167 1997 -1167 0 1
rlabel polysilicon 1997 -1173 1997 -1173 0 3
rlabel polysilicon 2004 -1167 2004 -1167 0 1
rlabel polysilicon 2004 -1173 2004 -1173 0 3
rlabel polysilicon 2011 -1167 2011 -1167 0 1
rlabel polysilicon 2011 -1173 2011 -1173 0 3
rlabel polysilicon 2018 -1167 2018 -1167 0 1
rlabel polysilicon 2018 -1173 2018 -1173 0 3
rlabel polysilicon 2025 -1167 2025 -1167 0 1
rlabel polysilicon 2025 -1173 2025 -1173 0 3
rlabel polysilicon 2032 -1167 2032 -1167 0 1
rlabel polysilicon 2032 -1173 2032 -1173 0 3
rlabel polysilicon 2039 -1167 2039 -1167 0 1
rlabel polysilicon 2039 -1173 2039 -1173 0 3
rlabel polysilicon 2046 -1167 2046 -1167 0 1
rlabel polysilicon 2046 -1173 2046 -1173 0 3
rlabel polysilicon 2053 -1167 2053 -1167 0 1
rlabel polysilicon 2053 -1173 2053 -1173 0 3
rlabel polysilicon 2060 -1167 2060 -1167 0 1
rlabel polysilicon 2060 -1173 2060 -1173 0 3
rlabel polysilicon 2067 -1167 2067 -1167 0 1
rlabel polysilicon 2067 -1173 2067 -1173 0 3
rlabel polysilicon 2074 -1167 2074 -1167 0 1
rlabel polysilicon 2074 -1173 2074 -1173 0 3
rlabel polysilicon 2081 -1167 2081 -1167 0 1
rlabel polysilicon 2081 -1173 2081 -1173 0 3
rlabel polysilicon 2088 -1167 2088 -1167 0 1
rlabel polysilicon 2088 -1173 2088 -1173 0 3
rlabel polysilicon 2095 -1167 2095 -1167 0 1
rlabel polysilicon 2095 -1173 2095 -1173 0 3
rlabel polysilicon 2102 -1167 2102 -1167 0 1
rlabel polysilicon 2102 -1173 2102 -1173 0 3
rlabel polysilicon 2109 -1167 2109 -1167 0 1
rlabel polysilicon 2109 -1173 2109 -1173 0 3
rlabel polysilicon 2116 -1167 2116 -1167 0 1
rlabel polysilicon 2116 -1173 2116 -1173 0 3
rlabel polysilicon 2123 -1167 2123 -1167 0 1
rlabel polysilicon 2123 -1173 2123 -1173 0 3
rlabel polysilicon 2130 -1167 2130 -1167 0 1
rlabel polysilicon 2130 -1173 2130 -1173 0 3
rlabel polysilicon 2137 -1167 2137 -1167 0 1
rlabel polysilicon 2137 -1173 2137 -1173 0 3
rlabel polysilicon 2144 -1167 2144 -1167 0 1
rlabel polysilicon 2144 -1173 2144 -1173 0 3
rlabel polysilicon 2151 -1167 2151 -1167 0 1
rlabel polysilicon 2151 -1173 2151 -1173 0 3
rlabel polysilicon 2158 -1167 2158 -1167 0 1
rlabel polysilicon 2158 -1173 2158 -1173 0 3
rlabel polysilicon 2165 -1167 2165 -1167 0 1
rlabel polysilicon 2165 -1173 2165 -1173 0 3
rlabel polysilicon 2172 -1167 2172 -1167 0 1
rlabel polysilicon 2172 -1173 2172 -1173 0 3
rlabel polysilicon 2179 -1167 2179 -1167 0 1
rlabel polysilicon 2179 -1173 2179 -1173 0 3
rlabel polysilicon 2186 -1167 2186 -1167 0 1
rlabel polysilicon 2186 -1173 2186 -1173 0 3
rlabel polysilicon 2193 -1167 2193 -1167 0 1
rlabel polysilicon 2193 -1173 2193 -1173 0 3
rlabel polysilicon 2200 -1167 2200 -1167 0 1
rlabel polysilicon 2200 -1173 2200 -1173 0 3
rlabel polysilicon 2207 -1167 2207 -1167 0 1
rlabel polysilicon 2207 -1173 2207 -1173 0 3
rlabel polysilicon 2214 -1167 2214 -1167 0 1
rlabel polysilicon 2214 -1173 2214 -1173 0 3
rlabel polysilicon 2221 -1167 2221 -1167 0 1
rlabel polysilicon 2221 -1173 2221 -1173 0 3
rlabel polysilicon 2228 -1167 2228 -1167 0 1
rlabel polysilicon 2228 -1173 2228 -1173 0 3
rlabel polysilicon 2235 -1167 2235 -1167 0 1
rlabel polysilicon 2235 -1173 2235 -1173 0 3
rlabel polysilicon 2242 -1167 2242 -1167 0 1
rlabel polysilicon 2242 -1173 2242 -1173 0 3
rlabel polysilicon 2249 -1167 2249 -1167 0 1
rlabel polysilicon 2249 -1173 2249 -1173 0 3
rlabel polysilicon 2256 -1167 2256 -1167 0 1
rlabel polysilicon 2256 -1173 2256 -1173 0 3
rlabel polysilicon 2263 -1167 2263 -1167 0 1
rlabel polysilicon 2263 -1173 2263 -1173 0 3
rlabel polysilicon 2270 -1167 2270 -1167 0 1
rlabel polysilicon 2270 -1173 2270 -1173 0 3
rlabel polysilicon 2277 -1167 2277 -1167 0 1
rlabel polysilicon 2277 -1173 2277 -1173 0 3
rlabel polysilicon 2284 -1167 2284 -1167 0 1
rlabel polysilicon 2284 -1173 2284 -1173 0 3
rlabel polysilicon 2291 -1167 2291 -1167 0 1
rlabel polysilicon 2291 -1173 2291 -1173 0 3
rlabel polysilicon 2298 -1167 2298 -1167 0 1
rlabel polysilicon 2298 -1173 2298 -1173 0 3
rlabel polysilicon 2305 -1167 2305 -1167 0 1
rlabel polysilicon 2305 -1173 2305 -1173 0 3
rlabel polysilicon 2312 -1167 2312 -1167 0 1
rlabel polysilicon 2312 -1173 2312 -1173 0 3
rlabel polysilicon 2319 -1167 2319 -1167 0 1
rlabel polysilicon 2319 -1173 2319 -1173 0 3
rlabel polysilicon 2326 -1167 2326 -1167 0 1
rlabel polysilicon 2326 -1173 2326 -1173 0 3
rlabel polysilicon 2333 -1167 2333 -1167 0 1
rlabel polysilicon 2333 -1173 2333 -1173 0 3
rlabel polysilicon 2340 -1167 2340 -1167 0 1
rlabel polysilicon 2340 -1173 2340 -1173 0 3
rlabel polysilicon 2347 -1167 2347 -1167 0 1
rlabel polysilicon 2347 -1173 2347 -1173 0 3
rlabel polysilicon 2354 -1167 2354 -1167 0 1
rlabel polysilicon 2354 -1173 2354 -1173 0 3
rlabel polysilicon 2361 -1167 2361 -1167 0 1
rlabel polysilicon 2361 -1173 2361 -1173 0 3
rlabel polysilicon 2368 -1167 2368 -1167 0 1
rlabel polysilicon 2368 -1173 2368 -1173 0 3
rlabel polysilicon 2375 -1167 2375 -1167 0 1
rlabel polysilicon 2375 -1173 2375 -1173 0 3
rlabel polysilicon 2382 -1167 2382 -1167 0 1
rlabel polysilicon 2382 -1173 2382 -1173 0 3
rlabel polysilicon 2389 -1167 2389 -1167 0 1
rlabel polysilicon 2392 -1167 2392 -1167 0 2
rlabel polysilicon 2389 -1173 2389 -1173 0 3
rlabel polysilicon 2392 -1173 2392 -1173 0 4
rlabel polysilicon 2396 -1167 2396 -1167 0 1
rlabel polysilicon 2399 -1167 2399 -1167 0 2
rlabel polysilicon 2396 -1173 2396 -1173 0 3
rlabel polysilicon 2403 -1167 2403 -1167 0 1
rlabel polysilicon 2403 -1173 2403 -1173 0 3
rlabel polysilicon 2424 -1167 2424 -1167 0 1
rlabel polysilicon 2424 -1173 2424 -1173 0 3
rlabel polysilicon 2431 -1167 2431 -1167 0 1
rlabel polysilicon 2431 -1173 2431 -1173 0 3
rlabel polysilicon 2438 -1167 2438 -1167 0 1
rlabel polysilicon 2438 -1173 2438 -1173 0 3
rlabel polysilicon 5 -1350 5 -1350 0 2
rlabel polysilicon 2 -1356 2 -1356 0 3
rlabel polysilicon 9 -1350 9 -1350 0 1
rlabel polysilicon 9 -1356 9 -1356 0 3
rlabel polysilicon 19 -1350 19 -1350 0 2
rlabel polysilicon 16 -1356 16 -1356 0 3
rlabel polysilicon 23 -1350 23 -1350 0 1
rlabel polysilicon 23 -1356 23 -1356 0 3
rlabel polysilicon 30 -1350 30 -1350 0 1
rlabel polysilicon 30 -1356 30 -1356 0 3
rlabel polysilicon 37 -1350 37 -1350 0 1
rlabel polysilicon 37 -1356 37 -1356 0 3
rlabel polysilicon 44 -1350 44 -1350 0 1
rlabel polysilicon 44 -1356 44 -1356 0 3
rlabel polysilicon 51 -1350 51 -1350 0 1
rlabel polysilicon 51 -1356 51 -1356 0 3
rlabel polysilicon 58 -1350 58 -1350 0 1
rlabel polysilicon 58 -1356 58 -1356 0 3
rlabel polysilicon 65 -1350 65 -1350 0 1
rlabel polysilicon 72 -1350 72 -1350 0 1
rlabel polysilicon 72 -1356 72 -1356 0 3
rlabel polysilicon 79 -1350 79 -1350 0 1
rlabel polysilicon 82 -1356 82 -1356 0 4
rlabel polysilicon 86 -1350 86 -1350 0 1
rlabel polysilicon 86 -1356 86 -1356 0 3
rlabel polysilicon 93 -1350 93 -1350 0 1
rlabel polysilicon 93 -1356 93 -1356 0 3
rlabel polysilicon 100 -1350 100 -1350 0 1
rlabel polysilicon 100 -1356 100 -1356 0 3
rlabel polysilicon 107 -1350 107 -1350 0 1
rlabel polysilicon 107 -1356 107 -1356 0 3
rlabel polysilicon 114 -1350 114 -1350 0 1
rlabel polysilicon 114 -1356 114 -1356 0 3
rlabel polysilicon 121 -1350 121 -1350 0 1
rlabel polysilicon 124 -1350 124 -1350 0 2
rlabel polysilicon 121 -1356 121 -1356 0 3
rlabel polysilicon 124 -1356 124 -1356 0 4
rlabel polysilicon 128 -1350 128 -1350 0 1
rlabel polysilicon 128 -1356 128 -1356 0 3
rlabel polysilicon 135 -1350 135 -1350 0 1
rlabel polysilicon 135 -1356 135 -1356 0 3
rlabel polysilicon 142 -1350 142 -1350 0 1
rlabel polysilicon 142 -1356 142 -1356 0 3
rlabel polysilicon 149 -1350 149 -1350 0 1
rlabel polysilicon 149 -1356 149 -1356 0 3
rlabel polysilicon 156 -1350 156 -1350 0 1
rlabel polysilicon 156 -1356 156 -1356 0 3
rlabel polysilicon 163 -1350 163 -1350 0 1
rlabel polysilicon 163 -1356 163 -1356 0 3
rlabel polysilicon 170 -1350 170 -1350 0 1
rlabel polysilicon 170 -1356 170 -1356 0 3
rlabel polysilicon 177 -1350 177 -1350 0 1
rlabel polysilicon 177 -1356 177 -1356 0 3
rlabel polysilicon 184 -1350 184 -1350 0 1
rlabel polysilicon 184 -1356 184 -1356 0 3
rlabel polysilicon 191 -1350 191 -1350 0 1
rlabel polysilicon 191 -1356 191 -1356 0 3
rlabel polysilicon 198 -1350 198 -1350 0 1
rlabel polysilicon 198 -1356 198 -1356 0 3
rlabel polysilicon 205 -1350 205 -1350 0 1
rlabel polysilicon 208 -1350 208 -1350 0 2
rlabel polysilicon 205 -1356 205 -1356 0 3
rlabel polysilicon 208 -1356 208 -1356 0 4
rlabel polysilicon 212 -1350 212 -1350 0 1
rlabel polysilicon 212 -1356 212 -1356 0 3
rlabel polysilicon 219 -1350 219 -1350 0 1
rlabel polysilicon 219 -1356 219 -1356 0 3
rlabel polysilicon 229 -1350 229 -1350 0 2
rlabel polysilicon 226 -1356 226 -1356 0 3
rlabel polysilicon 229 -1356 229 -1356 0 4
rlabel polysilicon 233 -1350 233 -1350 0 1
rlabel polysilicon 233 -1356 233 -1356 0 3
rlabel polysilicon 240 -1350 240 -1350 0 1
rlabel polysilicon 240 -1356 240 -1356 0 3
rlabel polysilicon 247 -1350 247 -1350 0 1
rlabel polysilicon 247 -1356 247 -1356 0 3
rlabel polysilicon 250 -1356 250 -1356 0 4
rlabel polysilicon 254 -1356 254 -1356 0 3
rlabel polysilicon 257 -1356 257 -1356 0 4
rlabel polysilicon 261 -1350 261 -1350 0 1
rlabel polysilicon 261 -1356 261 -1356 0 3
rlabel polysilicon 268 -1350 268 -1350 0 1
rlabel polysilicon 271 -1356 271 -1356 0 4
rlabel polysilicon 275 -1350 275 -1350 0 1
rlabel polysilicon 275 -1356 275 -1356 0 3
rlabel polysilicon 282 -1350 282 -1350 0 1
rlabel polysilicon 282 -1356 282 -1356 0 3
rlabel polysilicon 289 -1350 289 -1350 0 1
rlabel polysilicon 289 -1356 289 -1356 0 3
rlabel polysilicon 296 -1350 296 -1350 0 1
rlabel polysilicon 296 -1356 296 -1356 0 3
rlabel polysilicon 303 -1350 303 -1350 0 1
rlabel polysilicon 303 -1356 303 -1356 0 3
rlabel polysilicon 310 -1350 310 -1350 0 1
rlabel polysilicon 310 -1356 310 -1356 0 3
rlabel polysilicon 317 -1350 317 -1350 0 1
rlabel polysilicon 317 -1356 317 -1356 0 3
rlabel polysilicon 324 -1350 324 -1350 0 1
rlabel polysilicon 324 -1356 324 -1356 0 3
rlabel polysilicon 331 -1350 331 -1350 0 1
rlabel polysilicon 331 -1356 331 -1356 0 3
rlabel polysilicon 338 -1350 338 -1350 0 1
rlabel polysilicon 338 -1356 338 -1356 0 3
rlabel polysilicon 345 -1350 345 -1350 0 1
rlabel polysilicon 345 -1356 345 -1356 0 3
rlabel polysilicon 352 -1350 352 -1350 0 1
rlabel polysilicon 352 -1356 352 -1356 0 3
rlabel polysilicon 359 -1350 359 -1350 0 1
rlabel polysilicon 359 -1356 359 -1356 0 3
rlabel polysilicon 366 -1350 366 -1350 0 1
rlabel polysilicon 366 -1356 366 -1356 0 3
rlabel polysilicon 373 -1350 373 -1350 0 1
rlabel polysilicon 373 -1356 373 -1356 0 3
rlabel polysilicon 380 -1350 380 -1350 0 1
rlabel polysilicon 380 -1356 380 -1356 0 3
rlabel polysilicon 387 -1350 387 -1350 0 1
rlabel polysilicon 387 -1356 387 -1356 0 3
rlabel polysilicon 394 -1350 394 -1350 0 1
rlabel polysilicon 394 -1356 394 -1356 0 3
rlabel polysilicon 401 -1350 401 -1350 0 1
rlabel polysilicon 401 -1356 401 -1356 0 3
rlabel polysilicon 408 -1350 408 -1350 0 1
rlabel polysilicon 408 -1356 408 -1356 0 3
rlabel polysilicon 415 -1350 415 -1350 0 1
rlabel polysilicon 415 -1356 415 -1356 0 3
rlabel polysilicon 422 -1350 422 -1350 0 1
rlabel polysilicon 422 -1356 422 -1356 0 3
rlabel polysilicon 429 -1350 429 -1350 0 1
rlabel polysilicon 429 -1356 429 -1356 0 3
rlabel polysilicon 436 -1350 436 -1350 0 1
rlabel polysilicon 436 -1356 436 -1356 0 3
rlabel polysilicon 443 -1350 443 -1350 0 1
rlabel polysilicon 443 -1356 443 -1356 0 3
rlabel polysilicon 450 -1350 450 -1350 0 1
rlabel polysilicon 450 -1356 450 -1356 0 3
rlabel polysilicon 457 -1350 457 -1350 0 1
rlabel polysilicon 457 -1356 457 -1356 0 3
rlabel polysilicon 464 -1350 464 -1350 0 1
rlabel polysilicon 464 -1356 464 -1356 0 3
rlabel polysilicon 471 -1350 471 -1350 0 1
rlabel polysilicon 471 -1356 471 -1356 0 3
rlabel polysilicon 478 -1350 478 -1350 0 1
rlabel polysilicon 478 -1356 478 -1356 0 3
rlabel polysilicon 485 -1350 485 -1350 0 1
rlabel polysilicon 485 -1356 485 -1356 0 3
rlabel polysilicon 492 -1350 492 -1350 0 1
rlabel polysilicon 492 -1356 492 -1356 0 3
rlabel polysilicon 499 -1350 499 -1350 0 1
rlabel polysilicon 499 -1356 499 -1356 0 3
rlabel polysilicon 506 -1350 506 -1350 0 1
rlabel polysilicon 506 -1356 506 -1356 0 3
rlabel polysilicon 513 -1350 513 -1350 0 1
rlabel polysilicon 513 -1356 513 -1356 0 3
rlabel polysilicon 520 -1350 520 -1350 0 1
rlabel polysilicon 520 -1356 520 -1356 0 3
rlabel polysilicon 527 -1350 527 -1350 0 1
rlabel polysilicon 527 -1356 527 -1356 0 3
rlabel polysilicon 534 -1350 534 -1350 0 1
rlabel polysilicon 534 -1356 534 -1356 0 3
rlabel polysilicon 541 -1350 541 -1350 0 1
rlabel polysilicon 541 -1356 541 -1356 0 3
rlabel polysilicon 548 -1350 548 -1350 0 1
rlabel polysilicon 548 -1356 548 -1356 0 3
rlabel polysilicon 555 -1350 555 -1350 0 1
rlabel polysilicon 555 -1356 555 -1356 0 3
rlabel polysilicon 562 -1350 562 -1350 0 1
rlabel polysilicon 562 -1356 562 -1356 0 3
rlabel polysilicon 569 -1350 569 -1350 0 1
rlabel polysilicon 569 -1356 569 -1356 0 3
rlabel polysilicon 576 -1350 576 -1350 0 1
rlabel polysilicon 576 -1356 576 -1356 0 3
rlabel polysilicon 583 -1350 583 -1350 0 1
rlabel polysilicon 583 -1356 583 -1356 0 3
rlabel polysilicon 590 -1350 590 -1350 0 1
rlabel polysilicon 590 -1356 590 -1356 0 3
rlabel polysilicon 597 -1350 597 -1350 0 1
rlabel polysilicon 597 -1356 597 -1356 0 3
rlabel polysilicon 604 -1350 604 -1350 0 1
rlabel polysilicon 607 -1350 607 -1350 0 2
rlabel polysilicon 604 -1356 604 -1356 0 3
rlabel polysilicon 607 -1356 607 -1356 0 4
rlabel polysilicon 611 -1350 611 -1350 0 1
rlabel polysilicon 611 -1356 611 -1356 0 3
rlabel polysilicon 618 -1350 618 -1350 0 1
rlabel polysilicon 618 -1356 618 -1356 0 3
rlabel polysilicon 625 -1350 625 -1350 0 1
rlabel polysilicon 625 -1356 625 -1356 0 3
rlabel polysilicon 632 -1350 632 -1350 0 1
rlabel polysilicon 632 -1356 632 -1356 0 3
rlabel polysilicon 639 -1350 639 -1350 0 1
rlabel polysilicon 642 -1350 642 -1350 0 2
rlabel polysilicon 639 -1356 639 -1356 0 3
rlabel polysilicon 642 -1356 642 -1356 0 4
rlabel polysilicon 646 -1350 646 -1350 0 1
rlabel polysilicon 646 -1356 646 -1356 0 3
rlabel polysilicon 653 -1350 653 -1350 0 1
rlabel polysilicon 653 -1356 653 -1356 0 3
rlabel polysilicon 660 -1350 660 -1350 0 1
rlabel polysilicon 660 -1356 660 -1356 0 3
rlabel polysilicon 667 -1350 667 -1350 0 1
rlabel polysilicon 667 -1356 667 -1356 0 3
rlabel polysilicon 674 -1350 674 -1350 0 1
rlabel polysilicon 677 -1350 677 -1350 0 2
rlabel polysilicon 674 -1356 674 -1356 0 3
rlabel polysilicon 677 -1356 677 -1356 0 4
rlabel polysilicon 681 -1350 681 -1350 0 1
rlabel polysilicon 681 -1356 681 -1356 0 3
rlabel polysilicon 688 -1350 688 -1350 0 1
rlabel polysilicon 688 -1356 688 -1356 0 3
rlabel polysilicon 695 -1350 695 -1350 0 1
rlabel polysilicon 695 -1356 695 -1356 0 3
rlabel polysilicon 702 -1350 702 -1350 0 1
rlabel polysilicon 702 -1356 702 -1356 0 3
rlabel polysilicon 709 -1350 709 -1350 0 1
rlabel polysilicon 709 -1356 709 -1356 0 3
rlabel polysilicon 716 -1350 716 -1350 0 1
rlabel polysilicon 716 -1356 716 -1356 0 3
rlabel polysilicon 723 -1350 723 -1350 0 1
rlabel polysilicon 726 -1350 726 -1350 0 2
rlabel polysilicon 726 -1356 726 -1356 0 4
rlabel polysilicon 730 -1350 730 -1350 0 1
rlabel polysilicon 730 -1356 730 -1356 0 3
rlabel polysilicon 737 -1350 737 -1350 0 1
rlabel polysilicon 737 -1356 737 -1356 0 3
rlabel polysilicon 744 -1350 744 -1350 0 1
rlabel polysilicon 744 -1356 744 -1356 0 3
rlabel polysilicon 751 -1350 751 -1350 0 1
rlabel polysilicon 751 -1356 751 -1356 0 3
rlabel polysilicon 758 -1350 758 -1350 0 1
rlabel polysilicon 758 -1356 758 -1356 0 3
rlabel polysilicon 765 -1350 765 -1350 0 1
rlabel polysilicon 765 -1356 765 -1356 0 3
rlabel polysilicon 772 -1350 772 -1350 0 1
rlabel polysilicon 772 -1356 772 -1356 0 3
rlabel polysilicon 779 -1350 779 -1350 0 1
rlabel polysilicon 782 -1350 782 -1350 0 2
rlabel polysilicon 779 -1356 779 -1356 0 3
rlabel polysilicon 782 -1356 782 -1356 0 4
rlabel polysilicon 786 -1350 786 -1350 0 1
rlabel polysilicon 789 -1350 789 -1350 0 2
rlabel polysilicon 786 -1356 786 -1356 0 3
rlabel polysilicon 789 -1356 789 -1356 0 4
rlabel polysilicon 793 -1350 793 -1350 0 1
rlabel polysilicon 796 -1350 796 -1350 0 2
rlabel polysilicon 796 -1356 796 -1356 0 4
rlabel polysilicon 800 -1350 800 -1350 0 1
rlabel polysilicon 800 -1356 800 -1356 0 3
rlabel polysilicon 807 -1350 807 -1350 0 1
rlabel polysilicon 807 -1356 807 -1356 0 3
rlabel polysilicon 814 -1350 814 -1350 0 1
rlabel polysilicon 814 -1356 814 -1356 0 3
rlabel polysilicon 821 -1350 821 -1350 0 1
rlabel polysilicon 821 -1356 821 -1356 0 3
rlabel polysilicon 828 -1350 828 -1350 0 1
rlabel polysilicon 831 -1350 831 -1350 0 2
rlabel polysilicon 828 -1356 828 -1356 0 3
rlabel polysilicon 831 -1356 831 -1356 0 4
rlabel polysilicon 835 -1350 835 -1350 0 1
rlabel polysilicon 835 -1356 835 -1356 0 3
rlabel polysilicon 838 -1356 838 -1356 0 4
rlabel polysilicon 842 -1350 842 -1350 0 1
rlabel polysilicon 842 -1356 842 -1356 0 3
rlabel polysilicon 849 -1350 849 -1350 0 1
rlabel polysilicon 849 -1356 849 -1356 0 3
rlabel polysilicon 856 -1350 856 -1350 0 1
rlabel polysilicon 856 -1356 856 -1356 0 3
rlabel polysilicon 863 -1350 863 -1350 0 1
rlabel polysilicon 866 -1350 866 -1350 0 2
rlabel polysilicon 866 -1356 866 -1356 0 4
rlabel polysilicon 870 -1356 870 -1356 0 3
rlabel polysilicon 880 -1350 880 -1350 0 2
rlabel polysilicon 877 -1356 877 -1356 0 3
rlabel polysilicon 880 -1356 880 -1356 0 4
rlabel polysilicon 884 -1350 884 -1350 0 1
rlabel polysilicon 884 -1356 884 -1356 0 3
rlabel polysilicon 891 -1350 891 -1350 0 1
rlabel polysilicon 894 -1350 894 -1350 0 2
rlabel polysilicon 891 -1356 891 -1356 0 3
rlabel polysilicon 894 -1356 894 -1356 0 4
rlabel polysilicon 898 -1350 898 -1350 0 1
rlabel polysilicon 898 -1356 898 -1356 0 3
rlabel polysilicon 905 -1350 905 -1350 0 1
rlabel polysilicon 905 -1356 905 -1356 0 3
rlabel polysilicon 912 -1350 912 -1350 0 1
rlabel polysilicon 912 -1356 912 -1356 0 3
rlabel polysilicon 919 -1350 919 -1350 0 1
rlabel polysilicon 919 -1356 919 -1356 0 3
rlabel polysilicon 926 -1350 926 -1350 0 1
rlabel polysilicon 926 -1356 926 -1356 0 3
rlabel polysilicon 933 -1350 933 -1350 0 1
rlabel polysilicon 933 -1356 933 -1356 0 3
rlabel polysilicon 940 -1350 940 -1350 0 1
rlabel polysilicon 940 -1356 940 -1356 0 3
rlabel polysilicon 947 -1350 947 -1350 0 1
rlabel polysilicon 947 -1356 947 -1356 0 3
rlabel polysilicon 954 -1350 954 -1350 0 1
rlabel polysilicon 957 -1350 957 -1350 0 2
rlabel polysilicon 954 -1356 954 -1356 0 3
rlabel polysilicon 957 -1356 957 -1356 0 4
rlabel polysilicon 961 -1350 961 -1350 0 1
rlabel polysilicon 961 -1356 961 -1356 0 3
rlabel polysilicon 968 -1350 968 -1350 0 1
rlabel polysilicon 968 -1356 968 -1356 0 3
rlabel polysilicon 975 -1350 975 -1350 0 1
rlabel polysilicon 975 -1356 975 -1356 0 3
rlabel polysilicon 985 -1350 985 -1350 0 2
rlabel polysilicon 982 -1356 982 -1356 0 3
rlabel polysilicon 985 -1356 985 -1356 0 4
rlabel polysilicon 989 -1350 989 -1350 0 1
rlabel polysilicon 992 -1350 992 -1350 0 2
rlabel polysilicon 989 -1356 989 -1356 0 3
rlabel polysilicon 992 -1356 992 -1356 0 4
rlabel polysilicon 996 -1350 996 -1350 0 1
rlabel polysilicon 999 -1350 999 -1350 0 2
rlabel polysilicon 996 -1356 996 -1356 0 3
rlabel polysilicon 999 -1356 999 -1356 0 4
rlabel polysilicon 1003 -1350 1003 -1350 0 1
rlabel polysilicon 1006 -1350 1006 -1350 0 2
rlabel polysilicon 1003 -1356 1003 -1356 0 3
rlabel polysilicon 1006 -1356 1006 -1356 0 4
rlabel polysilicon 1010 -1350 1010 -1350 0 1
rlabel polysilicon 1013 -1350 1013 -1350 0 2
rlabel polysilicon 1010 -1356 1010 -1356 0 3
rlabel polysilicon 1013 -1356 1013 -1356 0 4
rlabel polysilicon 1017 -1350 1017 -1350 0 1
rlabel polysilicon 1017 -1356 1017 -1356 0 3
rlabel polysilicon 1024 -1350 1024 -1350 0 1
rlabel polysilicon 1024 -1356 1024 -1356 0 3
rlabel polysilicon 1031 -1350 1031 -1350 0 1
rlabel polysilicon 1031 -1356 1031 -1356 0 3
rlabel polysilicon 1038 -1350 1038 -1350 0 1
rlabel polysilicon 1041 -1350 1041 -1350 0 2
rlabel polysilicon 1038 -1356 1038 -1356 0 3
rlabel polysilicon 1041 -1356 1041 -1356 0 4
rlabel polysilicon 1045 -1350 1045 -1350 0 1
rlabel polysilicon 1045 -1356 1045 -1356 0 3
rlabel polysilicon 1052 -1350 1052 -1350 0 1
rlabel polysilicon 1052 -1356 1052 -1356 0 3
rlabel polysilicon 1059 -1350 1059 -1350 0 1
rlabel polysilicon 1059 -1356 1059 -1356 0 3
rlabel polysilicon 1066 -1350 1066 -1350 0 1
rlabel polysilicon 1066 -1356 1066 -1356 0 3
rlabel polysilicon 1073 -1350 1073 -1350 0 1
rlabel polysilicon 1073 -1356 1073 -1356 0 3
rlabel polysilicon 1080 -1350 1080 -1350 0 1
rlabel polysilicon 1080 -1356 1080 -1356 0 3
rlabel polysilicon 1087 -1350 1087 -1350 0 1
rlabel polysilicon 1087 -1356 1087 -1356 0 3
rlabel polysilicon 1094 -1350 1094 -1350 0 1
rlabel polysilicon 1094 -1356 1094 -1356 0 3
rlabel polysilicon 1101 -1350 1101 -1350 0 1
rlabel polysilicon 1104 -1350 1104 -1350 0 2
rlabel polysilicon 1101 -1356 1101 -1356 0 3
rlabel polysilicon 1104 -1356 1104 -1356 0 4
rlabel polysilicon 1108 -1350 1108 -1350 0 1
rlabel polysilicon 1108 -1356 1108 -1356 0 3
rlabel polysilicon 1115 -1350 1115 -1350 0 1
rlabel polysilicon 1115 -1356 1115 -1356 0 3
rlabel polysilicon 1122 -1350 1122 -1350 0 1
rlabel polysilicon 1122 -1356 1122 -1356 0 3
rlabel polysilicon 1129 -1350 1129 -1350 0 1
rlabel polysilicon 1129 -1356 1129 -1356 0 3
rlabel polysilicon 1136 -1350 1136 -1350 0 1
rlabel polysilicon 1136 -1356 1136 -1356 0 3
rlabel polysilicon 1143 -1350 1143 -1350 0 1
rlabel polysilicon 1143 -1356 1143 -1356 0 3
rlabel polysilicon 1150 -1350 1150 -1350 0 1
rlabel polysilicon 1153 -1350 1153 -1350 0 2
rlabel polysilicon 1150 -1356 1150 -1356 0 3
rlabel polysilicon 1153 -1356 1153 -1356 0 4
rlabel polysilicon 1157 -1350 1157 -1350 0 1
rlabel polysilicon 1157 -1356 1157 -1356 0 3
rlabel polysilicon 1164 -1350 1164 -1350 0 1
rlabel polysilicon 1164 -1356 1164 -1356 0 3
rlabel polysilicon 1171 -1350 1171 -1350 0 1
rlabel polysilicon 1171 -1356 1171 -1356 0 3
rlabel polysilicon 1178 -1350 1178 -1350 0 1
rlabel polysilicon 1178 -1356 1178 -1356 0 3
rlabel polysilicon 1185 -1350 1185 -1350 0 1
rlabel polysilicon 1185 -1356 1185 -1356 0 3
rlabel polysilicon 1192 -1350 1192 -1350 0 1
rlabel polysilicon 1192 -1356 1192 -1356 0 3
rlabel polysilicon 1199 -1350 1199 -1350 0 1
rlabel polysilicon 1199 -1356 1199 -1356 0 3
rlabel polysilicon 1206 -1350 1206 -1350 0 1
rlabel polysilicon 1206 -1356 1206 -1356 0 3
rlabel polysilicon 1213 -1350 1213 -1350 0 1
rlabel polysilicon 1216 -1350 1216 -1350 0 2
rlabel polysilicon 1213 -1356 1213 -1356 0 3
rlabel polysilicon 1220 -1350 1220 -1350 0 1
rlabel polysilicon 1220 -1356 1220 -1356 0 3
rlabel polysilicon 1227 -1350 1227 -1350 0 1
rlabel polysilicon 1227 -1356 1227 -1356 0 3
rlabel polysilicon 1234 -1350 1234 -1350 0 1
rlabel polysilicon 1234 -1356 1234 -1356 0 3
rlabel polysilicon 1241 -1350 1241 -1350 0 1
rlabel polysilicon 1241 -1356 1241 -1356 0 3
rlabel polysilicon 1248 -1350 1248 -1350 0 1
rlabel polysilicon 1248 -1356 1248 -1356 0 3
rlabel polysilicon 1255 -1350 1255 -1350 0 1
rlabel polysilicon 1255 -1356 1255 -1356 0 3
rlabel polysilicon 1262 -1350 1262 -1350 0 1
rlabel polysilicon 1262 -1356 1262 -1356 0 3
rlabel polysilicon 1269 -1350 1269 -1350 0 1
rlabel polysilicon 1269 -1356 1269 -1356 0 3
rlabel polysilicon 1276 -1350 1276 -1350 0 1
rlabel polysilicon 1276 -1356 1276 -1356 0 3
rlabel polysilicon 1283 -1350 1283 -1350 0 1
rlabel polysilicon 1283 -1356 1283 -1356 0 3
rlabel polysilicon 1290 -1350 1290 -1350 0 1
rlabel polysilicon 1290 -1356 1290 -1356 0 3
rlabel polysilicon 1297 -1350 1297 -1350 0 1
rlabel polysilicon 1297 -1356 1297 -1356 0 3
rlabel polysilicon 1304 -1350 1304 -1350 0 1
rlabel polysilicon 1304 -1356 1304 -1356 0 3
rlabel polysilicon 1311 -1350 1311 -1350 0 1
rlabel polysilicon 1311 -1356 1311 -1356 0 3
rlabel polysilicon 1318 -1350 1318 -1350 0 1
rlabel polysilicon 1318 -1356 1318 -1356 0 3
rlabel polysilicon 1325 -1350 1325 -1350 0 1
rlabel polysilicon 1325 -1356 1325 -1356 0 3
rlabel polysilicon 1332 -1350 1332 -1350 0 1
rlabel polysilicon 1332 -1356 1332 -1356 0 3
rlabel polysilicon 1339 -1350 1339 -1350 0 1
rlabel polysilicon 1339 -1356 1339 -1356 0 3
rlabel polysilicon 1346 -1350 1346 -1350 0 1
rlabel polysilicon 1346 -1356 1346 -1356 0 3
rlabel polysilicon 1353 -1350 1353 -1350 0 1
rlabel polysilicon 1353 -1356 1353 -1356 0 3
rlabel polysilicon 1360 -1350 1360 -1350 0 1
rlabel polysilicon 1360 -1356 1360 -1356 0 3
rlabel polysilicon 1367 -1350 1367 -1350 0 1
rlabel polysilicon 1370 -1350 1370 -1350 0 2
rlabel polysilicon 1367 -1356 1367 -1356 0 3
rlabel polysilicon 1370 -1356 1370 -1356 0 4
rlabel polysilicon 1374 -1350 1374 -1350 0 1
rlabel polysilicon 1374 -1356 1374 -1356 0 3
rlabel polysilicon 1381 -1350 1381 -1350 0 1
rlabel polysilicon 1384 -1350 1384 -1350 0 2
rlabel polysilicon 1381 -1356 1381 -1356 0 3
rlabel polysilicon 1384 -1356 1384 -1356 0 4
rlabel polysilicon 1388 -1350 1388 -1350 0 1
rlabel polysilicon 1391 -1350 1391 -1350 0 2
rlabel polysilicon 1388 -1356 1388 -1356 0 3
rlabel polysilicon 1395 -1350 1395 -1350 0 1
rlabel polysilicon 1395 -1356 1395 -1356 0 3
rlabel polysilicon 1402 -1350 1402 -1350 0 1
rlabel polysilicon 1402 -1356 1402 -1356 0 3
rlabel polysilicon 1409 -1350 1409 -1350 0 1
rlabel polysilicon 1409 -1356 1409 -1356 0 3
rlabel polysilicon 1416 -1350 1416 -1350 0 1
rlabel polysilicon 1416 -1356 1416 -1356 0 3
rlabel polysilicon 1419 -1356 1419 -1356 0 4
rlabel polysilicon 1423 -1350 1423 -1350 0 1
rlabel polysilicon 1423 -1356 1423 -1356 0 3
rlabel polysilicon 1430 -1350 1430 -1350 0 1
rlabel polysilicon 1433 -1350 1433 -1350 0 2
rlabel polysilicon 1430 -1356 1430 -1356 0 3
rlabel polysilicon 1433 -1356 1433 -1356 0 4
rlabel polysilicon 1437 -1350 1437 -1350 0 1
rlabel polysilicon 1437 -1356 1437 -1356 0 3
rlabel polysilicon 1447 -1350 1447 -1350 0 2
rlabel polysilicon 1444 -1356 1444 -1356 0 3
rlabel polysilicon 1451 -1350 1451 -1350 0 1
rlabel polysilicon 1451 -1356 1451 -1356 0 3
rlabel polysilicon 1458 -1350 1458 -1350 0 1
rlabel polysilicon 1458 -1356 1458 -1356 0 3
rlabel polysilicon 1465 -1350 1465 -1350 0 1
rlabel polysilicon 1465 -1356 1465 -1356 0 3
rlabel polysilicon 1472 -1350 1472 -1350 0 1
rlabel polysilicon 1472 -1356 1472 -1356 0 3
rlabel polysilicon 1479 -1350 1479 -1350 0 1
rlabel polysilicon 1479 -1356 1479 -1356 0 3
rlabel polysilicon 1486 -1350 1486 -1350 0 1
rlabel polysilicon 1486 -1356 1486 -1356 0 3
rlabel polysilicon 1493 -1350 1493 -1350 0 1
rlabel polysilicon 1493 -1356 1493 -1356 0 3
rlabel polysilicon 1500 -1350 1500 -1350 0 1
rlabel polysilicon 1500 -1356 1500 -1356 0 3
rlabel polysilicon 1507 -1350 1507 -1350 0 1
rlabel polysilicon 1510 -1350 1510 -1350 0 2
rlabel polysilicon 1510 -1356 1510 -1356 0 4
rlabel polysilicon 1514 -1350 1514 -1350 0 1
rlabel polysilicon 1514 -1356 1514 -1356 0 3
rlabel polysilicon 1521 -1350 1521 -1350 0 1
rlabel polysilicon 1521 -1356 1521 -1356 0 3
rlabel polysilicon 1528 -1350 1528 -1350 0 1
rlabel polysilicon 1528 -1356 1528 -1356 0 3
rlabel polysilicon 1535 -1350 1535 -1350 0 1
rlabel polysilicon 1535 -1356 1535 -1356 0 3
rlabel polysilicon 1542 -1350 1542 -1350 0 1
rlabel polysilicon 1542 -1356 1542 -1356 0 3
rlabel polysilicon 1549 -1350 1549 -1350 0 1
rlabel polysilicon 1549 -1356 1549 -1356 0 3
rlabel polysilicon 1556 -1350 1556 -1350 0 1
rlabel polysilicon 1556 -1356 1556 -1356 0 3
rlabel polysilicon 1563 -1350 1563 -1350 0 1
rlabel polysilicon 1563 -1356 1563 -1356 0 3
rlabel polysilicon 1570 -1350 1570 -1350 0 1
rlabel polysilicon 1570 -1356 1570 -1356 0 3
rlabel polysilicon 1577 -1350 1577 -1350 0 1
rlabel polysilicon 1577 -1356 1577 -1356 0 3
rlabel polysilicon 1584 -1350 1584 -1350 0 1
rlabel polysilicon 1584 -1356 1584 -1356 0 3
rlabel polysilicon 1591 -1350 1591 -1350 0 1
rlabel polysilicon 1591 -1356 1591 -1356 0 3
rlabel polysilicon 1598 -1350 1598 -1350 0 1
rlabel polysilicon 1598 -1356 1598 -1356 0 3
rlabel polysilicon 1605 -1350 1605 -1350 0 1
rlabel polysilicon 1605 -1356 1605 -1356 0 3
rlabel polysilicon 1612 -1350 1612 -1350 0 1
rlabel polysilicon 1612 -1356 1612 -1356 0 3
rlabel polysilicon 1619 -1350 1619 -1350 0 1
rlabel polysilicon 1619 -1356 1619 -1356 0 3
rlabel polysilicon 1626 -1350 1626 -1350 0 1
rlabel polysilicon 1626 -1356 1626 -1356 0 3
rlabel polysilicon 1633 -1350 1633 -1350 0 1
rlabel polysilicon 1633 -1356 1633 -1356 0 3
rlabel polysilicon 1640 -1350 1640 -1350 0 1
rlabel polysilicon 1640 -1356 1640 -1356 0 3
rlabel polysilicon 1647 -1350 1647 -1350 0 1
rlabel polysilicon 1647 -1356 1647 -1356 0 3
rlabel polysilicon 1654 -1350 1654 -1350 0 1
rlabel polysilicon 1654 -1356 1654 -1356 0 3
rlabel polysilicon 1661 -1350 1661 -1350 0 1
rlabel polysilicon 1661 -1356 1661 -1356 0 3
rlabel polysilicon 1668 -1350 1668 -1350 0 1
rlabel polysilicon 1668 -1356 1668 -1356 0 3
rlabel polysilicon 1675 -1350 1675 -1350 0 1
rlabel polysilicon 1675 -1356 1675 -1356 0 3
rlabel polysilicon 1678 -1356 1678 -1356 0 4
rlabel polysilicon 1682 -1350 1682 -1350 0 1
rlabel polysilicon 1682 -1356 1682 -1356 0 3
rlabel polysilicon 1689 -1350 1689 -1350 0 1
rlabel polysilicon 1689 -1356 1689 -1356 0 3
rlabel polysilicon 1696 -1350 1696 -1350 0 1
rlabel polysilicon 1696 -1356 1696 -1356 0 3
rlabel polysilicon 1703 -1350 1703 -1350 0 1
rlabel polysilicon 1703 -1356 1703 -1356 0 3
rlabel polysilicon 1710 -1350 1710 -1350 0 1
rlabel polysilicon 1710 -1356 1710 -1356 0 3
rlabel polysilicon 1717 -1350 1717 -1350 0 1
rlabel polysilicon 1717 -1356 1717 -1356 0 3
rlabel polysilicon 1724 -1350 1724 -1350 0 1
rlabel polysilicon 1724 -1356 1724 -1356 0 3
rlabel polysilicon 1731 -1350 1731 -1350 0 1
rlabel polysilicon 1731 -1356 1731 -1356 0 3
rlabel polysilicon 1738 -1350 1738 -1350 0 1
rlabel polysilicon 1738 -1356 1738 -1356 0 3
rlabel polysilicon 1745 -1350 1745 -1350 0 1
rlabel polysilicon 1745 -1356 1745 -1356 0 3
rlabel polysilicon 1752 -1350 1752 -1350 0 1
rlabel polysilicon 1752 -1356 1752 -1356 0 3
rlabel polysilicon 1759 -1350 1759 -1350 0 1
rlabel polysilicon 1759 -1356 1759 -1356 0 3
rlabel polysilicon 1766 -1350 1766 -1350 0 1
rlabel polysilicon 1766 -1356 1766 -1356 0 3
rlabel polysilicon 1773 -1350 1773 -1350 0 1
rlabel polysilicon 1773 -1356 1773 -1356 0 3
rlabel polysilicon 1780 -1350 1780 -1350 0 1
rlabel polysilicon 1780 -1356 1780 -1356 0 3
rlabel polysilicon 1787 -1350 1787 -1350 0 1
rlabel polysilicon 1787 -1356 1787 -1356 0 3
rlabel polysilicon 1794 -1350 1794 -1350 0 1
rlabel polysilicon 1794 -1356 1794 -1356 0 3
rlabel polysilicon 1797 -1356 1797 -1356 0 4
rlabel polysilicon 1801 -1350 1801 -1350 0 1
rlabel polysilicon 1801 -1356 1801 -1356 0 3
rlabel polysilicon 1808 -1350 1808 -1350 0 1
rlabel polysilicon 1808 -1356 1808 -1356 0 3
rlabel polysilicon 1815 -1350 1815 -1350 0 1
rlabel polysilicon 1815 -1356 1815 -1356 0 3
rlabel polysilicon 1822 -1350 1822 -1350 0 1
rlabel polysilicon 1822 -1356 1822 -1356 0 3
rlabel polysilicon 1829 -1350 1829 -1350 0 1
rlabel polysilicon 1829 -1356 1829 -1356 0 3
rlabel polysilicon 1836 -1350 1836 -1350 0 1
rlabel polysilicon 1836 -1356 1836 -1356 0 3
rlabel polysilicon 1843 -1350 1843 -1350 0 1
rlabel polysilicon 1843 -1356 1843 -1356 0 3
rlabel polysilicon 1850 -1350 1850 -1350 0 1
rlabel polysilicon 1850 -1356 1850 -1356 0 3
rlabel polysilicon 1857 -1350 1857 -1350 0 1
rlabel polysilicon 1857 -1356 1857 -1356 0 3
rlabel polysilicon 1864 -1350 1864 -1350 0 1
rlabel polysilicon 1864 -1356 1864 -1356 0 3
rlabel polysilicon 1871 -1350 1871 -1350 0 1
rlabel polysilicon 1871 -1356 1871 -1356 0 3
rlabel polysilicon 1878 -1350 1878 -1350 0 1
rlabel polysilicon 1878 -1356 1878 -1356 0 3
rlabel polysilicon 1885 -1350 1885 -1350 0 1
rlabel polysilicon 1885 -1356 1885 -1356 0 3
rlabel polysilicon 1892 -1350 1892 -1350 0 1
rlabel polysilicon 1892 -1356 1892 -1356 0 3
rlabel polysilicon 1899 -1350 1899 -1350 0 1
rlabel polysilicon 1899 -1356 1899 -1356 0 3
rlabel polysilicon 1906 -1350 1906 -1350 0 1
rlabel polysilicon 1906 -1356 1906 -1356 0 3
rlabel polysilicon 1913 -1350 1913 -1350 0 1
rlabel polysilicon 1913 -1356 1913 -1356 0 3
rlabel polysilicon 1920 -1350 1920 -1350 0 1
rlabel polysilicon 1920 -1356 1920 -1356 0 3
rlabel polysilicon 1927 -1350 1927 -1350 0 1
rlabel polysilicon 1927 -1356 1927 -1356 0 3
rlabel polysilicon 1934 -1350 1934 -1350 0 1
rlabel polysilicon 1934 -1356 1934 -1356 0 3
rlabel polysilicon 1941 -1350 1941 -1350 0 1
rlabel polysilicon 1941 -1356 1941 -1356 0 3
rlabel polysilicon 1948 -1350 1948 -1350 0 1
rlabel polysilicon 1948 -1356 1948 -1356 0 3
rlabel polysilicon 1955 -1350 1955 -1350 0 1
rlabel polysilicon 1955 -1356 1955 -1356 0 3
rlabel polysilicon 1962 -1350 1962 -1350 0 1
rlabel polysilicon 1962 -1356 1962 -1356 0 3
rlabel polysilicon 1969 -1350 1969 -1350 0 1
rlabel polysilicon 1969 -1356 1969 -1356 0 3
rlabel polysilicon 1976 -1350 1976 -1350 0 1
rlabel polysilicon 1976 -1356 1976 -1356 0 3
rlabel polysilicon 1983 -1350 1983 -1350 0 1
rlabel polysilicon 1983 -1356 1983 -1356 0 3
rlabel polysilicon 1990 -1350 1990 -1350 0 1
rlabel polysilicon 1990 -1356 1990 -1356 0 3
rlabel polysilicon 1997 -1350 1997 -1350 0 1
rlabel polysilicon 1997 -1356 1997 -1356 0 3
rlabel polysilicon 2004 -1350 2004 -1350 0 1
rlabel polysilicon 2004 -1356 2004 -1356 0 3
rlabel polysilicon 2011 -1350 2011 -1350 0 1
rlabel polysilicon 2011 -1356 2011 -1356 0 3
rlabel polysilicon 2018 -1350 2018 -1350 0 1
rlabel polysilicon 2018 -1356 2018 -1356 0 3
rlabel polysilicon 2025 -1350 2025 -1350 0 1
rlabel polysilicon 2025 -1356 2025 -1356 0 3
rlabel polysilicon 2032 -1350 2032 -1350 0 1
rlabel polysilicon 2032 -1356 2032 -1356 0 3
rlabel polysilicon 2039 -1350 2039 -1350 0 1
rlabel polysilicon 2039 -1356 2039 -1356 0 3
rlabel polysilicon 2046 -1350 2046 -1350 0 1
rlabel polysilicon 2046 -1356 2046 -1356 0 3
rlabel polysilicon 2053 -1350 2053 -1350 0 1
rlabel polysilicon 2053 -1356 2053 -1356 0 3
rlabel polysilicon 2060 -1350 2060 -1350 0 1
rlabel polysilicon 2060 -1356 2060 -1356 0 3
rlabel polysilicon 2067 -1350 2067 -1350 0 1
rlabel polysilicon 2067 -1356 2067 -1356 0 3
rlabel polysilicon 2074 -1350 2074 -1350 0 1
rlabel polysilicon 2074 -1356 2074 -1356 0 3
rlabel polysilicon 2081 -1350 2081 -1350 0 1
rlabel polysilicon 2081 -1356 2081 -1356 0 3
rlabel polysilicon 2088 -1350 2088 -1350 0 1
rlabel polysilicon 2088 -1356 2088 -1356 0 3
rlabel polysilicon 2095 -1350 2095 -1350 0 1
rlabel polysilicon 2095 -1356 2095 -1356 0 3
rlabel polysilicon 2102 -1350 2102 -1350 0 1
rlabel polysilicon 2102 -1356 2102 -1356 0 3
rlabel polysilicon 2109 -1350 2109 -1350 0 1
rlabel polysilicon 2109 -1356 2109 -1356 0 3
rlabel polysilicon 2116 -1350 2116 -1350 0 1
rlabel polysilicon 2116 -1356 2116 -1356 0 3
rlabel polysilicon 2123 -1350 2123 -1350 0 1
rlabel polysilicon 2123 -1356 2123 -1356 0 3
rlabel polysilicon 2130 -1350 2130 -1350 0 1
rlabel polysilicon 2130 -1356 2130 -1356 0 3
rlabel polysilicon 2137 -1350 2137 -1350 0 1
rlabel polysilicon 2137 -1356 2137 -1356 0 3
rlabel polysilicon 2144 -1350 2144 -1350 0 1
rlabel polysilicon 2144 -1356 2144 -1356 0 3
rlabel polysilicon 2151 -1350 2151 -1350 0 1
rlabel polysilicon 2151 -1356 2151 -1356 0 3
rlabel polysilicon 2158 -1350 2158 -1350 0 1
rlabel polysilicon 2158 -1356 2158 -1356 0 3
rlabel polysilicon 2165 -1350 2165 -1350 0 1
rlabel polysilicon 2165 -1356 2165 -1356 0 3
rlabel polysilicon 2172 -1350 2172 -1350 0 1
rlabel polysilicon 2172 -1356 2172 -1356 0 3
rlabel polysilicon 2179 -1350 2179 -1350 0 1
rlabel polysilicon 2179 -1356 2179 -1356 0 3
rlabel polysilicon 2186 -1350 2186 -1350 0 1
rlabel polysilicon 2186 -1356 2186 -1356 0 3
rlabel polysilicon 2193 -1350 2193 -1350 0 1
rlabel polysilicon 2193 -1356 2193 -1356 0 3
rlabel polysilicon 2200 -1350 2200 -1350 0 1
rlabel polysilicon 2200 -1356 2200 -1356 0 3
rlabel polysilicon 2207 -1350 2207 -1350 0 1
rlabel polysilicon 2207 -1356 2207 -1356 0 3
rlabel polysilicon 2214 -1350 2214 -1350 0 1
rlabel polysilicon 2214 -1356 2214 -1356 0 3
rlabel polysilicon 2221 -1350 2221 -1350 0 1
rlabel polysilicon 2221 -1356 2221 -1356 0 3
rlabel polysilicon 2228 -1350 2228 -1350 0 1
rlabel polysilicon 2228 -1356 2228 -1356 0 3
rlabel polysilicon 2235 -1350 2235 -1350 0 1
rlabel polysilicon 2235 -1356 2235 -1356 0 3
rlabel polysilicon 2242 -1350 2242 -1350 0 1
rlabel polysilicon 2242 -1356 2242 -1356 0 3
rlabel polysilicon 2249 -1350 2249 -1350 0 1
rlabel polysilicon 2249 -1356 2249 -1356 0 3
rlabel polysilicon 2256 -1350 2256 -1350 0 1
rlabel polysilicon 2256 -1356 2256 -1356 0 3
rlabel polysilicon 2263 -1350 2263 -1350 0 1
rlabel polysilicon 2263 -1356 2263 -1356 0 3
rlabel polysilicon 2270 -1350 2270 -1350 0 1
rlabel polysilicon 2270 -1356 2270 -1356 0 3
rlabel polysilicon 2277 -1350 2277 -1350 0 1
rlabel polysilicon 2277 -1356 2277 -1356 0 3
rlabel polysilicon 2284 -1350 2284 -1350 0 1
rlabel polysilicon 2284 -1356 2284 -1356 0 3
rlabel polysilicon 2291 -1350 2291 -1350 0 1
rlabel polysilicon 2291 -1356 2291 -1356 0 3
rlabel polysilicon 2298 -1350 2298 -1350 0 1
rlabel polysilicon 2298 -1356 2298 -1356 0 3
rlabel polysilicon 2305 -1350 2305 -1350 0 1
rlabel polysilicon 2305 -1356 2305 -1356 0 3
rlabel polysilicon 2312 -1350 2312 -1350 0 1
rlabel polysilicon 2312 -1356 2312 -1356 0 3
rlabel polysilicon 2319 -1350 2319 -1350 0 1
rlabel polysilicon 2319 -1356 2319 -1356 0 3
rlabel polysilicon 2326 -1350 2326 -1350 0 1
rlabel polysilicon 2326 -1356 2326 -1356 0 3
rlabel polysilicon 2333 -1350 2333 -1350 0 1
rlabel polysilicon 2333 -1356 2333 -1356 0 3
rlabel polysilicon 2340 -1350 2340 -1350 0 1
rlabel polysilicon 2343 -1350 2343 -1350 0 2
rlabel polysilicon 2340 -1356 2340 -1356 0 3
rlabel polysilicon 2343 -1356 2343 -1356 0 4
rlabel polysilicon 2347 -1350 2347 -1350 0 1
rlabel polysilicon 2347 -1356 2347 -1356 0 3
rlabel polysilicon 2354 -1350 2354 -1350 0 1
rlabel polysilicon 2354 -1356 2354 -1356 0 3
rlabel polysilicon 2361 -1350 2361 -1350 0 1
rlabel polysilicon 2361 -1356 2361 -1356 0 3
rlabel polysilicon 2368 -1350 2368 -1350 0 1
rlabel polysilicon 2368 -1356 2368 -1356 0 3
rlabel polysilicon 2375 -1350 2375 -1350 0 1
rlabel polysilicon 2375 -1356 2375 -1356 0 3
rlabel polysilicon 2382 -1350 2382 -1350 0 1
rlabel polysilicon 2382 -1356 2382 -1356 0 3
rlabel polysilicon 2389 -1350 2389 -1350 0 1
rlabel polysilicon 2389 -1356 2389 -1356 0 3
rlabel polysilicon 2396 -1350 2396 -1350 0 1
rlabel polysilicon 2396 -1356 2396 -1356 0 3
rlabel polysilicon 2403 -1350 2403 -1350 0 1
rlabel polysilicon 2403 -1356 2403 -1356 0 3
rlabel polysilicon 2410 -1350 2410 -1350 0 1
rlabel polysilicon 2410 -1356 2410 -1356 0 3
rlabel polysilicon 2417 -1350 2417 -1350 0 1
rlabel polysilicon 2417 -1356 2417 -1356 0 3
rlabel polysilicon 2424 -1350 2424 -1350 0 1
rlabel polysilicon 2424 -1356 2424 -1356 0 3
rlabel polysilicon 2431 -1350 2431 -1350 0 1
rlabel polysilicon 2431 -1356 2431 -1356 0 3
rlabel polysilicon 2438 -1350 2438 -1350 0 1
rlabel polysilicon 2438 -1356 2438 -1356 0 3
rlabel polysilicon 2445 -1350 2445 -1350 0 1
rlabel polysilicon 2445 -1356 2445 -1356 0 3
rlabel polysilicon 2452 -1350 2452 -1350 0 1
rlabel polysilicon 2452 -1356 2452 -1356 0 3
rlabel polysilicon 2459 -1350 2459 -1350 0 1
rlabel polysilicon 2459 -1356 2459 -1356 0 3
rlabel polysilicon 2466 -1350 2466 -1350 0 1
rlabel polysilicon 2466 -1356 2466 -1356 0 3
rlabel polysilicon 2473 -1350 2473 -1350 0 1
rlabel polysilicon 2473 -1356 2473 -1356 0 3
rlabel polysilicon 2480 -1350 2480 -1350 0 1
rlabel polysilicon 2480 -1356 2480 -1356 0 3
rlabel polysilicon 2487 -1350 2487 -1350 0 1
rlabel polysilicon 2487 -1356 2487 -1356 0 3
rlabel polysilicon 2494 -1350 2494 -1350 0 1
rlabel polysilicon 2494 -1356 2494 -1356 0 3
rlabel polysilicon 2501 -1350 2501 -1350 0 1
rlabel polysilicon 2501 -1356 2501 -1356 0 3
rlabel polysilicon 2508 -1350 2508 -1350 0 1
rlabel polysilicon 2508 -1356 2508 -1356 0 3
rlabel polysilicon 2515 -1350 2515 -1350 0 1
rlabel polysilicon 2515 -1356 2515 -1356 0 3
rlabel polysilicon 2522 -1350 2522 -1350 0 1
rlabel polysilicon 2522 -1356 2522 -1356 0 3
rlabel polysilicon 2529 -1350 2529 -1350 0 1
rlabel polysilicon 2529 -1356 2529 -1356 0 3
rlabel polysilicon 2536 -1350 2536 -1350 0 1
rlabel polysilicon 2536 -1356 2536 -1356 0 3
rlabel polysilicon 2543 -1350 2543 -1350 0 1
rlabel polysilicon 2543 -1356 2543 -1356 0 3
rlabel polysilicon 2550 -1350 2550 -1350 0 1
rlabel polysilicon 2550 -1356 2550 -1356 0 3
rlabel polysilicon 2557 -1350 2557 -1350 0 1
rlabel polysilicon 2557 -1356 2557 -1356 0 3
rlabel polysilicon 2564 -1350 2564 -1350 0 1
rlabel polysilicon 2564 -1356 2564 -1356 0 3
rlabel polysilicon 2571 -1350 2571 -1350 0 1
rlabel polysilicon 2571 -1356 2571 -1356 0 3
rlabel polysilicon 2578 -1350 2578 -1350 0 1
rlabel polysilicon 2578 -1356 2578 -1356 0 3
rlabel polysilicon 2 -1527 2 -1527 0 1
rlabel polysilicon 2 -1533 2 -1533 0 3
rlabel polysilicon 9 -1527 9 -1527 0 1
rlabel polysilicon 9 -1533 9 -1533 0 3
rlabel polysilicon 16 -1527 16 -1527 0 1
rlabel polysilicon 19 -1527 19 -1527 0 2
rlabel polysilicon 23 -1527 23 -1527 0 1
rlabel polysilicon 26 -1527 26 -1527 0 2
rlabel polysilicon 23 -1533 23 -1533 0 3
rlabel polysilicon 30 -1527 30 -1527 0 1
rlabel polysilicon 30 -1533 30 -1533 0 3
rlabel polysilicon 37 -1527 37 -1527 0 1
rlabel polysilicon 40 -1527 40 -1527 0 2
rlabel polysilicon 37 -1533 37 -1533 0 3
rlabel polysilicon 40 -1533 40 -1533 0 4
rlabel polysilicon 44 -1527 44 -1527 0 1
rlabel polysilicon 47 -1527 47 -1527 0 2
rlabel polysilicon 44 -1533 44 -1533 0 3
rlabel polysilicon 47 -1533 47 -1533 0 4
rlabel polysilicon 51 -1527 51 -1527 0 1
rlabel polysilicon 54 -1527 54 -1527 0 2
rlabel polysilicon 51 -1533 51 -1533 0 3
rlabel polysilicon 58 -1527 58 -1527 0 1
rlabel polysilicon 58 -1533 58 -1533 0 3
rlabel polysilicon 65 -1533 65 -1533 0 3
rlabel polysilicon 72 -1527 72 -1527 0 1
rlabel polysilicon 72 -1533 72 -1533 0 3
rlabel polysilicon 79 -1527 79 -1527 0 1
rlabel polysilicon 79 -1533 79 -1533 0 3
rlabel polysilicon 86 -1527 86 -1527 0 1
rlabel polysilicon 89 -1527 89 -1527 0 2
rlabel polysilicon 86 -1533 86 -1533 0 3
rlabel polysilicon 89 -1533 89 -1533 0 4
rlabel polysilicon 93 -1527 93 -1527 0 1
rlabel polysilicon 93 -1533 93 -1533 0 3
rlabel polysilicon 100 -1527 100 -1527 0 1
rlabel polysilicon 100 -1533 100 -1533 0 3
rlabel polysilicon 107 -1527 107 -1527 0 1
rlabel polysilicon 110 -1527 110 -1527 0 2
rlabel polysilicon 110 -1533 110 -1533 0 4
rlabel polysilicon 114 -1527 114 -1527 0 1
rlabel polysilicon 117 -1527 117 -1527 0 2
rlabel polysilicon 114 -1533 114 -1533 0 3
rlabel polysilicon 117 -1533 117 -1533 0 4
rlabel polysilicon 121 -1527 121 -1527 0 1
rlabel polysilicon 121 -1533 121 -1533 0 3
rlabel polysilicon 128 -1527 128 -1527 0 1
rlabel polysilicon 128 -1533 128 -1533 0 3
rlabel polysilicon 135 -1527 135 -1527 0 1
rlabel polysilicon 135 -1533 135 -1533 0 3
rlabel polysilicon 142 -1527 142 -1527 0 1
rlabel polysilicon 142 -1533 142 -1533 0 3
rlabel polysilicon 149 -1527 149 -1527 0 1
rlabel polysilicon 149 -1533 149 -1533 0 3
rlabel polysilicon 156 -1527 156 -1527 0 1
rlabel polysilicon 156 -1533 156 -1533 0 3
rlabel polysilicon 163 -1527 163 -1527 0 1
rlabel polysilicon 163 -1533 163 -1533 0 3
rlabel polysilicon 170 -1527 170 -1527 0 1
rlabel polysilicon 170 -1533 170 -1533 0 3
rlabel polysilicon 177 -1527 177 -1527 0 1
rlabel polysilicon 177 -1533 177 -1533 0 3
rlabel polysilicon 184 -1527 184 -1527 0 1
rlabel polysilicon 184 -1533 184 -1533 0 3
rlabel polysilicon 191 -1527 191 -1527 0 1
rlabel polysilicon 191 -1533 191 -1533 0 3
rlabel polysilicon 198 -1527 198 -1527 0 1
rlabel polysilicon 201 -1527 201 -1527 0 2
rlabel polysilicon 198 -1533 198 -1533 0 3
rlabel polysilicon 201 -1533 201 -1533 0 4
rlabel polysilicon 208 -1527 208 -1527 0 2
rlabel polysilicon 205 -1533 205 -1533 0 3
rlabel polysilicon 208 -1533 208 -1533 0 4
rlabel polysilicon 212 -1527 212 -1527 0 1
rlabel polysilicon 212 -1533 212 -1533 0 3
rlabel polysilicon 219 -1527 219 -1527 0 1
rlabel polysilicon 219 -1533 219 -1533 0 3
rlabel polysilicon 226 -1527 226 -1527 0 1
rlabel polysilicon 226 -1533 226 -1533 0 3
rlabel polysilicon 233 -1527 233 -1527 0 1
rlabel polysilicon 236 -1527 236 -1527 0 2
rlabel polysilicon 233 -1533 233 -1533 0 3
rlabel polysilicon 236 -1533 236 -1533 0 4
rlabel polysilicon 240 -1527 240 -1527 0 1
rlabel polysilicon 240 -1533 240 -1533 0 3
rlabel polysilicon 247 -1527 247 -1527 0 1
rlabel polysilicon 247 -1533 247 -1533 0 3
rlabel polysilicon 254 -1527 254 -1527 0 1
rlabel polysilicon 254 -1533 254 -1533 0 3
rlabel polysilicon 261 -1527 261 -1527 0 1
rlabel polysilicon 261 -1533 261 -1533 0 3
rlabel polysilicon 268 -1527 268 -1527 0 1
rlabel polysilicon 268 -1533 268 -1533 0 3
rlabel polysilicon 275 -1527 275 -1527 0 1
rlabel polysilicon 275 -1533 275 -1533 0 3
rlabel polysilicon 282 -1527 282 -1527 0 1
rlabel polysilicon 282 -1533 282 -1533 0 3
rlabel polysilicon 289 -1527 289 -1527 0 1
rlabel polysilicon 289 -1533 289 -1533 0 3
rlabel polysilicon 296 -1527 296 -1527 0 1
rlabel polysilicon 296 -1533 296 -1533 0 3
rlabel polysilicon 303 -1527 303 -1527 0 1
rlabel polysilicon 303 -1533 303 -1533 0 3
rlabel polysilicon 310 -1527 310 -1527 0 1
rlabel polysilicon 310 -1533 310 -1533 0 3
rlabel polysilicon 317 -1527 317 -1527 0 1
rlabel polysilicon 317 -1533 317 -1533 0 3
rlabel polysilicon 324 -1527 324 -1527 0 1
rlabel polysilicon 324 -1533 324 -1533 0 3
rlabel polysilicon 331 -1527 331 -1527 0 1
rlabel polysilicon 331 -1533 331 -1533 0 3
rlabel polysilicon 338 -1527 338 -1527 0 1
rlabel polysilicon 338 -1533 338 -1533 0 3
rlabel polysilicon 345 -1527 345 -1527 0 1
rlabel polysilicon 345 -1533 345 -1533 0 3
rlabel polysilicon 352 -1527 352 -1527 0 1
rlabel polysilicon 352 -1533 352 -1533 0 3
rlabel polysilicon 359 -1527 359 -1527 0 1
rlabel polysilicon 359 -1533 359 -1533 0 3
rlabel polysilicon 366 -1527 366 -1527 0 1
rlabel polysilicon 366 -1533 366 -1533 0 3
rlabel polysilicon 373 -1527 373 -1527 0 1
rlabel polysilicon 373 -1533 373 -1533 0 3
rlabel polysilicon 380 -1527 380 -1527 0 1
rlabel polysilicon 380 -1533 380 -1533 0 3
rlabel polysilicon 387 -1527 387 -1527 0 1
rlabel polysilicon 387 -1533 387 -1533 0 3
rlabel polysilicon 394 -1527 394 -1527 0 1
rlabel polysilicon 394 -1533 394 -1533 0 3
rlabel polysilicon 401 -1527 401 -1527 0 1
rlabel polysilicon 401 -1533 401 -1533 0 3
rlabel polysilicon 408 -1527 408 -1527 0 1
rlabel polysilicon 408 -1533 408 -1533 0 3
rlabel polysilicon 415 -1527 415 -1527 0 1
rlabel polysilicon 415 -1533 415 -1533 0 3
rlabel polysilicon 422 -1527 422 -1527 0 1
rlabel polysilicon 422 -1533 422 -1533 0 3
rlabel polysilicon 429 -1527 429 -1527 0 1
rlabel polysilicon 429 -1533 429 -1533 0 3
rlabel polysilicon 436 -1527 436 -1527 0 1
rlabel polysilicon 436 -1533 436 -1533 0 3
rlabel polysilicon 443 -1527 443 -1527 0 1
rlabel polysilicon 443 -1533 443 -1533 0 3
rlabel polysilicon 450 -1527 450 -1527 0 1
rlabel polysilicon 450 -1533 450 -1533 0 3
rlabel polysilicon 457 -1527 457 -1527 0 1
rlabel polysilicon 457 -1533 457 -1533 0 3
rlabel polysilicon 464 -1527 464 -1527 0 1
rlabel polysilicon 464 -1533 464 -1533 0 3
rlabel polysilicon 471 -1527 471 -1527 0 1
rlabel polysilicon 471 -1533 471 -1533 0 3
rlabel polysilicon 478 -1527 478 -1527 0 1
rlabel polysilicon 478 -1533 478 -1533 0 3
rlabel polysilicon 485 -1527 485 -1527 0 1
rlabel polysilicon 485 -1533 485 -1533 0 3
rlabel polysilicon 492 -1527 492 -1527 0 1
rlabel polysilicon 492 -1533 492 -1533 0 3
rlabel polysilicon 499 -1527 499 -1527 0 1
rlabel polysilicon 499 -1533 499 -1533 0 3
rlabel polysilicon 506 -1527 506 -1527 0 1
rlabel polysilicon 506 -1533 506 -1533 0 3
rlabel polysilicon 513 -1527 513 -1527 0 1
rlabel polysilicon 516 -1527 516 -1527 0 2
rlabel polysilicon 513 -1533 513 -1533 0 3
rlabel polysilicon 516 -1533 516 -1533 0 4
rlabel polysilicon 520 -1527 520 -1527 0 1
rlabel polysilicon 520 -1533 520 -1533 0 3
rlabel polysilicon 527 -1527 527 -1527 0 1
rlabel polysilicon 527 -1533 527 -1533 0 3
rlabel polysilicon 534 -1527 534 -1527 0 1
rlabel polysilicon 534 -1533 534 -1533 0 3
rlabel polysilicon 541 -1527 541 -1527 0 1
rlabel polysilicon 541 -1533 541 -1533 0 3
rlabel polysilicon 548 -1527 548 -1527 0 1
rlabel polysilicon 548 -1533 548 -1533 0 3
rlabel polysilicon 555 -1527 555 -1527 0 1
rlabel polysilicon 555 -1533 555 -1533 0 3
rlabel polysilicon 562 -1527 562 -1527 0 1
rlabel polysilicon 562 -1533 562 -1533 0 3
rlabel polysilicon 569 -1527 569 -1527 0 1
rlabel polysilicon 569 -1533 569 -1533 0 3
rlabel polysilicon 576 -1527 576 -1527 0 1
rlabel polysilicon 576 -1533 576 -1533 0 3
rlabel polysilicon 583 -1527 583 -1527 0 1
rlabel polysilicon 583 -1533 583 -1533 0 3
rlabel polysilicon 593 -1527 593 -1527 0 2
rlabel polysilicon 590 -1533 590 -1533 0 3
rlabel polysilicon 593 -1533 593 -1533 0 4
rlabel polysilicon 597 -1527 597 -1527 0 1
rlabel polysilicon 597 -1533 597 -1533 0 3
rlabel polysilicon 604 -1527 604 -1527 0 1
rlabel polysilicon 604 -1533 604 -1533 0 3
rlabel polysilicon 611 -1527 611 -1527 0 1
rlabel polysilicon 611 -1533 611 -1533 0 3
rlabel polysilicon 618 -1527 618 -1527 0 1
rlabel polysilicon 618 -1533 618 -1533 0 3
rlabel polysilicon 625 -1527 625 -1527 0 1
rlabel polysilicon 628 -1527 628 -1527 0 2
rlabel polysilicon 625 -1533 625 -1533 0 3
rlabel polysilicon 628 -1533 628 -1533 0 4
rlabel polysilicon 632 -1527 632 -1527 0 1
rlabel polysilicon 632 -1533 632 -1533 0 3
rlabel polysilicon 639 -1527 639 -1527 0 1
rlabel polysilicon 642 -1527 642 -1527 0 2
rlabel polysilicon 639 -1533 639 -1533 0 3
rlabel polysilicon 642 -1533 642 -1533 0 4
rlabel polysilicon 646 -1527 646 -1527 0 1
rlabel polysilicon 646 -1533 646 -1533 0 3
rlabel polysilicon 653 -1527 653 -1527 0 1
rlabel polysilicon 653 -1533 653 -1533 0 3
rlabel polysilicon 660 -1527 660 -1527 0 1
rlabel polysilicon 660 -1533 660 -1533 0 3
rlabel polysilicon 667 -1527 667 -1527 0 1
rlabel polysilicon 667 -1533 667 -1533 0 3
rlabel polysilicon 674 -1527 674 -1527 0 1
rlabel polysilicon 674 -1533 674 -1533 0 3
rlabel polysilicon 681 -1527 681 -1527 0 1
rlabel polysilicon 681 -1533 681 -1533 0 3
rlabel polysilicon 688 -1527 688 -1527 0 1
rlabel polysilicon 691 -1527 691 -1527 0 2
rlabel polysilicon 688 -1533 688 -1533 0 3
rlabel polysilicon 691 -1533 691 -1533 0 4
rlabel polysilicon 695 -1527 695 -1527 0 1
rlabel polysilicon 695 -1533 695 -1533 0 3
rlabel polysilicon 702 -1527 702 -1527 0 1
rlabel polysilicon 702 -1533 702 -1533 0 3
rlabel polysilicon 709 -1527 709 -1527 0 1
rlabel polysilicon 709 -1533 709 -1533 0 3
rlabel polysilicon 716 -1527 716 -1527 0 1
rlabel polysilicon 716 -1533 716 -1533 0 3
rlabel polysilicon 723 -1527 723 -1527 0 1
rlabel polysilicon 723 -1533 723 -1533 0 3
rlabel polysilicon 730 -1527 730 -1527 0 1
rlabel polysilicon 730 -1533 730 -1533 0 3
rlabel polysilicon 737 -1527 737 -1527 0 1
rlabel polysilicon 740 -1527 740 -1527 0 2
rlabel polysilicon 737 -1533 737 -1533 0 3
rlabel polysilicon 744 -1527 744 -1527 0 1
rlabel polysilicon 744 -1533 744 -1533 0 3
rlabel polysilicon 751 -1527 751 -1527 0 1
rlabel polysilicon 751 -1533 751 -1533 0 3
rlabel polysilicon 758 -1527 758 -1527 0 1
rlabel polysilicon 758 -1533 758 -1533 0 3
rlabel polysilicon 765 -1527 765 -1527 0 1
rlabel polysilicon 765 -1533 765 -1533 0 3
rlabel polysilicon 772 -1527 772 -1527 0 1
rlabel polysilicon 772 -1533 772 -1533 0 3
rlabel polysilicon 779 -1527 779 -1527 0 1
rlabel polysilicon 779 -1533 779 -1533 0 3
rlabel polysilicon 786 -1527 786 -1527 0 1
rlabel polysilicon 786 -1533 786 -1533 0 3
rlabel polysilicon 793 -1527 793 -1527 0 1
rlabel polysilicon 796 -1527 796 -1527 0 2
rlabel polysilicon 793 -1533 793 -1533 0 3
rlabel polysilicon 796 -1533 796 -1533 0 4
rlabel polysilicon 800 -1527 800 -1527 0 1
rlabel polysilicon 800 -1533 800 -1533 0 3
rlabel polysilicon 807 -1527 807 -1527 0 1
rlabel polysilicon 807 -1533 807 -1533 0 3
rlabel polysilicon 810 -1533 810 -1533 0 4
rlabel polysilicon 814 -1527 814 -1527 0 1
rlabel polysilicon 814 -1533 814 -1533 0 3
rlabel polysilicon 824 -1527 824 -1527 0 2
rlabel polysilicon 821 -1533 821 -1533 0 3
rlabel polysilicon 824 -1533 824 -1533 0 4
rlabel polysilicon 828 -1527 828 -1527 0 1
rlabel polysilicon 828 -1533 828 -1533 0 3
rlabel polysilicon 835 -1527 835 -1527 0 1
rlabel polysilicon 835 -1533 835 -1533 0 3
rlabel polysilicon 842 -1527 842 -1527 0 1
rlabel polysilicon 842 -1533 842 -1533 0 3
rlabel polysilicon 849 -1527 849 -1527 0 1
rlabel polysilicon 849 -1533 849 -1533 0 3
rlabel polysilicon 856 -1527 856 -1527 0 1
rlabel polysilicon 856 -1533 856 -1533 0 3
rlabel polysilicon 863 -1527 863 -1527 0 1
rlabel polysilicon 866 -1527 866 -1527 0 2
rlabel polysilicon 863 -1533 863 -1533 0 3
rlabel polysilicon 866 -1533 866 -1533 0 4
rlabel polysilicon 870 -1527 870 -1527 0 1
rlabel polysilicon 870 -1533 870 -1533 0 3
rlabel polysilicon 877 -1527 877 -1527 0 1
rlabel polysilicon 880 -1527 880 -1527 0 2
rlabel polysilicon 880 -1533 880 -1533 0 4
rlabel polysilicon 884 -1527 884 -1527 0 1
rlabel polysilicon 887 -1527 887 -1527 0 2
rlabel polysilicon 887 -1533 887 -1533 0 4
rlabel polysilicon 891 -1527 891 -1527 0 1
rlabel polysilicon 891 -1533 891 -1533 0 3
rlabel polysilicon 898 -1527 898 -1527 0 1
rlabel polysilicon 898 -1533 898 -1533 0 3
rlabel polysilicon 905 -1527 905 -1527 0 1
rlabel polysilicon 908 -1527 908 -1527 0 2
rlabel polysilicon 905 -1533 905 -1533 0 3
rlabel polysilicon 912 -1527 912 -1527 0 1
rlabel polysilicon 912 -1533 912 -1533 0 3
rlabel polysilicon 919 -1527 919 -1527 0 1
rlabel polysilicon 919 -1533 919 -1533 0 3
rlabel polysilicon 926 -1527 926 -1527 0 1
rlabel polysilicon 926 -1533 926 -1533 0 3
rlabel polysilicon 933 -1527 933 -1527 0 1
rlabel polysilicon 933 -1533 933 -1533 0 3
rlabel polysilicon 940 -1527 940 -1527 0 1
rlabel polysilicon 943 -1527 943 -1527 0 2
rlabel polysilicon 940 -1533 940 -1533 0 3
rlabel polysilicon 943 -1533 943 -1533 0 4
rlabel polysilicon 947 -1527 947 -1527 0 1
rlabel polysilicon 947 -1533 947 -1533 0 3
rlabel polysilicon 954 -1527 954 -1527 0 1
rlabel polysilicon 954 -1533 954 -1533 0 3
rlabel polysilicon 961 -1527 961 -1527 0 1
rlabel polysilicon 961 -1533 961 -1533 0 3
rlabel polysilicon 964 -1533 964 -1533 0 4
rlabel polysilicon 968 -1527 968 -1527 0 1
rlabel polysilicon 968 -1533 968 -1533 0 3
rlabel polysilicon 975 -1527 975 -1527 0 1
rlabel polysilicon 975 -1533 975 -1533 0 3
rlabel polysilicon 982 -1527 982 -1527 0 1
rlabel polysilicon 982 -1533 982 -1533 0 3
rlabel polysilicon 989 -1527 989 -1527 0 1
rlabel polysilicon 989 -1533 989 -1533 0 3
rlabel polysilicon 996 -1527 996 -1527 0 1
rlabel polysilicon 996 -1533 996 -1533 0 3
rlabel polysilicon 1003 -1527 1003 -1527 0 1
rlabel polysilicon 1003 -1533 1003 -1533 0 3
rlabel polysilicon 1010 -1527 1010 -1527 0 1
rlabel polysilicon 1010 -1533 1010 -1533 0 3
rlabel polysilicon 1017 -1527 1017 -1527 0 1
rlabel polysilicon 1017 -1533 1017 -1533 0 3
rlabel polysilicon 1024 -1527 1024 -1527 0 1
rlabel polysilicon 1024 -1533 1024 -1533 0 3
rlabel polysilicon 1031 -1527 1031 -1527 0 1
rlabel polysilicon 1031 -1533 1031 -1533 0 3
rlabel polysilicon 1038 -1527 1038 -1527 0 1
rlabel polysilicon 1038 -1533 1038 -1533 0 3
rlabel polysilicon 1045 -1527 1045 -1527 0 1
rlabel polysilicon 1045 -1533 1045 -1533 0 3
rlabel polysilicon 1052 -1527 1052 -1527 0 1
rlabel polysilicon 1052 -1533 1052 -1533 0 3
rlabel polysilicon 1059 -1527 1059 -1527 0 1
rlabel polysilicon 1059 -1533 1059 -1533 0 3
rlabel polysilicon 1066 -1527 1066 -1527 0 1
rlabel polysilicon 1066 -1533 1066 -1533 0 3
rlabel polysilicon 1073 -1527 1073 -1527 0 1
rlabel polysilicon 1073 -1533 1073 -1533 0 3
rlabel polysilicon 1080 -1527 1080 -1527 0 1
rlabel polysilicon 1080 -1533 1080 -1533 0 3
rlabel polysilicon 1087 -1527 1087 -1527 0 1
rlabel polysilicon 1090 -1527 1090 -1527 0 2
rlabel polysilicon 1087 -1533 1087 -1533 0 3
rlabel polysilicon 1090 -1533 1090 -1533 0 4
rlabel polysilicon 1094 -1527 1094 -1527 0 1
rlabel polysilicon 1094 -1533 1094 -1533 0 3
rlabel polysilicon 1101 -1527 1101 -1527 0 1
rlabel polysilicon 1101 -1533 1101 -1533 0 3
rlabel polysilicon 1108 -1527 1108 -1527 0 1
rlabel polysilicon 1108 -1533 1108 -1533 0 3
rlabel polysilicon 1115 -1527 1115 -1527 0 1
rlabel polysilicon 1115 -1533 1115 -1533 0 3
rlabel polysilicon 1122 -1527 1122 -1527 0 1
rlabel polysilicon 1122 -1533 1122 -1533 0 3
rlabel polysilicon 1129 -1527 1129 -1527 0 1
rlabel polysilicon 1129 -1533 1129 -1533 0 3
rlabel polysilicon 1136 -1527 1136 -1527 0 1
rlabel polysilicon 1136 -1533 1136 -1533 0 3
rlabel polysilicon 1143 -1527 1143 -1527 0 1
rlabel polysilicon 1143 -1533 1143 -1533 0 3
rlabel polysilicon 1150 -1527 1150 -1527 0 1
rlabel polysilicon 1153 -1527 1153 -1527 0 2
rlabel polysilicon 1150 -1533 1150 -1533 0 3
rlabel polysilicon 1153 -1533 1153 -1533 0 4
rlabel polysilicon 1157 -1527 1157 -1527 0 1
rlabel polysilicon 1160 -1527 1160 -1527 0 2
rlabel polysilicon 1157 -1533 1157 -1533 0 3
rlabel polysilicon 1160 -1533 1160 -1533 0 4
rlabel polysilicon 1164 -1527 1164 -1527 0 1
rlabel polysilicon 1164 -1533 1164 -1533 0 3
rlabel polysilicon 1171 -1527 1171 -1527 0 1
rlabel polysilicon 1171 -1533 1171 -1533 0 3
rlabel polysilicon 1178 -1527 1178 -1527 0 1
rlabel polysilicon 1178 -1533 1178 -1533 0 3
rlabel polysilicon 1185 -1527 1185 -1527 0 1
rlabel polysilicon 1185 -1533 1185 -1533 0 3
rlabel polysilicon 1192 -1527 1192 -1527 0 1
rlabel polysilicon 1192 -1533 1192 -1533 0 3
rlabel polysilicon 1199 -1527 1199 -1527 0 1
rlabel polysilicon 1199 -1533 1199 -1533 0 3
rlabel polysilicon 1206 -1527 1206 -1527 0 1
rlabel polysilicon 1206 -1533 1206 -1533 0 3
rlabel polysilicon 1213 -1527 1213 -1527 0 1
rlabel polysilicon 1213 -1533 1213 -1533 0 3
rlabel polysilicon 1220 -1527 1220 -1527 0 1
rlabel polysilicon 1220 -1533 1220 -1533 0 3
rlabel polysilicon 1227 -1527 1227 -1527 0 1
rlabel polysilicon 1227 -1533 1227 -1533 0 3
rlabel polysilicon 1234 -1527 1234 -1527 0 1
rlabel polysilicon 1234 -1533 1234 -1533 0 3
rlabel polysilicon 1241 -1527 1241 -1527 0 1
rlabel polysilicon 1241 -1533 1241 -1533 0 3
rlabel polysilicon 1248 -1527 1248 -1527 0 1
rlabel polysilicon 1251 -1527 1251 -1527 0 2
rlabel polysilicon 1248 -1533 1248 -1533 0 3
rlabel polysilicon 1251 -1533 1251 -1533 0 4
rlabel polysilicon 1255 -1527 1255 -1527 0 1
rlabel polysilicon 1258 -1527 1258 -1527 0 2
rlabel polysilicon 1258 -1533 1258 -1533 0 4
rlabel polysilicon 1262 -1527 1262 -1527 0 1
rlabel polysilicon 1265 -1527 1265 -1527 0 2
rlabel polysilicon 1262 -1533 1262 -1533 0 3
rlabel polysilicon 1269 -1527 1269 -1527 0 1
rlabel polysilicon 1269 -1533 1269 -1533 0 3
rlabel polysilicon 1276 -1527 1276 -1527 0 1
rlabel polysilicon 1276 -1533 1276 -1533 0 3
rlabel polysilicon 1283 -1527 1283 -1527 0 1
rlabel polysilicon 1286 -1527 1286 -1527 0 2
rlabel polysilicon 1286 -1533 1286 -1533 0 4
rlabel polysilicon 1290 -1527 1290 -1527 0 1
rlabel polysilicon 1290 -1533 1290 -1533 0 3
rlabel polysilicon 1297 -1527 1297 -1527 0 1
rlabel polysilicon 1297 -1533 1297 -1533 0 3
rlabel polysilicon 1304 -1527 1304 -1527 0 1
rlabel polysilicon 1304 -1533 1304 -1533 0 3
rlabel polysilicon 1311 -1527 1311 -1527 0 1
rlabel polysilicon 1311 -1533 1311 -1533 0 3
rlabel polysilicon 1318 -1527 1318 -1527 0 1
rlabel polysilicon 1318 -1533 1318 -1533 0 3
rlabel polysilicon 1325 -1527 1325 -1527 0 1
rlabel polysilicon 1325 -1533 1325 -1533 0 3
rlabel polysilicon 1332 -1527 1332 -1527 0 1
rlabel polysilicon 1332 -1533 1332 -1533 0 3
rlabel polysilicon 1339 -1527 1339 -1527 0 1
rlabel polysilicon 1339 -1533 1339 -1533 0 3
rlabel polysilicon 1346 -1527 1346 -1527 0 1
rlabel polysilicon 1349 -1527 1349 -1527 0 2
rlabel polysilicon 1346 -1533 1346 -1533 0 3
rlabel polysilicon 1349 -1533 1349 -1533 0 4
rlabel polysilicon 1353 -1527 1353 -1527 0 1
rlabel polysilicon 1353 -1533 1353 -1533 0 3
rlabel polysilicon 1360 -1527 1360 -1527 0 1
rlabel polysilicon 1360 -1533 1360 -1533 0 3
rlabel polysilicon 1367 -1527 1367 -1527 0 1
rlabel polysilicon 1367 -1533 1367 -1533 0 3
rlabel polysilicon 1374 -1527 1374 -1527 0 1
rlabel polysilicon 1374 -1533 1374 -1533 0 3
rlabel polysilicon 1381 -1527 1381 -1527 0 1
rlabel polysilicon 1381 -1533 1381 -1533 0 3
rlabel polysilicon 1388 -1527 1388 -1527 0 1
rlabel polysilicon 1388 -1533 1388 -1533 0 3
rlabel polysilicon 1395 -1527 1395 -1527 0 1
rlabel polysilicon 1395 -1533 1395 -1533 0 3
rlabel polysilicon 1402 -1527 1402 -1527 0 1
rlabel polysilicon 1402 -1533 1402 -1533 0 3
rlabel polysilicon 1409 -1527 1409 -1527 0 1
rlabel polysilicon 1409 -1533 1409 -1533 0 3
rlabel polysilicon 1416 -1527 1416 -1527 0 1
rlabel polysilicon 1416 -1533 1416 -1533 0 3
rlabel polysilicon 1426 -1527 1426 -1527 0 2
rlabel polysilicon 1423 -1533 1423 -1533 0 3
rlabel polysilicon 1430 -1527 1430 -1527 0 1
rlabel polysilicon 1430 -1533 1430 -1533 0 3
rlabel polysilicon 1437 -1527 1437 -1527 0 1
rlabel polysilicon 1437 -1533 1437 -1533 0 3
rlabel polysilicon 1444 -1527 1444 -1527 0 1
rlabel polysilicon 1444 -1533 1444 -1533 0 3
rlabel polysilicon 1451 -1527 1451 -1527 0 1
rlabel polysilicon 1451 -1533 1451 -1533 0 3
rlabel polysilicon 1458 -1527 1458 -1527 0 1
rlabel polysilicon 1458 -1533 1458 -1533 0 3
rlabel polysilicon 1465 -1527 1465 -1527 0 1
rlabel polysilicon 1465 -1533 1465 -1533 0 3
rlabel polysilicon 1472 -1527 1472 -1527 0 1
rlabel polysilicon 1472 -1533 1472 -1533 0 3
rlabel polysilicon 1479 -1527 1479 -1527 0 1
rlabel polysilicon 1482 -1527 1482 -1527 0 2
rlabel polysilicon 1479 -1533 1479 -1533 0 3
rlabel polysilicon 1486 -1527 1486 -1527 0 1
rlabel polysilicon 1489 -1527 1489 -1527 0 2
rlabel polysilicon 1489 -1533 1489 -1533 0 4
rlabel polysilicon 1493 -1527 1493 -1527 0 1
rlabel polysilicon 1493 -1533 1493 -1533 0 3
rlabel polysilicon 1500 -1527 1500 -1527 0 1
rlabel polysilicon 1503 -1527 1503 -1527 0 2
rlabel polysilicon 1500 -1533 1500 -1533 0 3
rlabel polysilicon 1503 -1533 1503 -1533 0 4
rlabel polysilicon 1507 -1527 1507 -1527 0 1
rlabel polysilicon 1507 -1533 1507 -1533 0 3
rlabel polysilicon 1514 -1527 1514 -1527 0 1
rlabel polysilicon 1514 -1533 1514 -1533 0 3
rlabel polysilicon 1521 -1527 1521 -1527 0 1
rlabel polysilicon 1521 -1533 1521 -1533 0 3
rlabel polysilicon 1528 -1527 1528 -1527 0 1
rlabel polysilicon 1528 -1533 1528 -1533 0 3
rlabel polysilicon 1535 -1527 1535 -1527 0 1
rlabel polysilicon 1535 -1533 1535 -1533 0 3
rlabel polysilicon 1542 -1527 1542 -1527 0 1
rlabel polysilicon 1542 -1533 1542 -1533 0 3
rlabel polysilicon 1549 -1527 1549 -1527 0 1
rlabel polysilicon 1549 -1533 1549 -1533 0 3
rlabel polysilicon 1556 -1527 1556 -1527 0 1
rlabel polysilicon 1556 -1533 1556 -1533 0 3
rlabel polysilicon 1563 -1527 1563 -1527 0 1
rlabel polysilicon 1563 -1533 1563 -1533 0 3
rlabel polysilicon 1570 -1527 1570 -1527 0 1
rlabel polysilicon 1570 -1533 1570 -1533 0 3
rlabel polysilicon 1577 -1527 1577 -1527 0 1
rlabel polysilicon 1577 -1533 1577 -1533 0 3
rlabel polysilicon 1584 -1527 1584 -1527 0 1
rlabel polysilicon 1584 -1533 1584 -1533 0 3
rlabel polysilicon 1591 -1527 1591 -1527 0 1
rlabel polysilicon 1591 -1533 1591 -1533 0 3
rlabel polysilicon 1598 -1527 1598 -1527 0 1
rlabel polysilicon 1598 -1533 1598 -1533 0 3
rlabel polysilicon 1605 -1527 1605 -1527 0 1
rlabel polysilicon 1605 -1533 1605 -1533 0 3
rlabel polysilicon 1612 -1527 1612 -1527 0 1
rlabel polysilicon 1612 -1533 1612 -1533 0 3
rlabel polysilicon 1619 -1527 1619 -1527 0 1
rlabel polysilicon 1619 -1533 1619 -1533 0 3
rlabel polysilicon 1626 -1527 1626 -1527 0 1
rlabel polysilicon 1626 -1533 1626 -1533 0 3
rlabel polysilicon 1633 -1527 1633 -1527 0 1
rlabel polysilicon 1633 -1533 1633 -1533 0 3
rlabel polysilicon 1640 -1527 1640 -1527 0 1
rlabel polysilicon 1640 -1533 1640 -1533 0 3
rlabel polysilicon 1647 -1527 1647 -1527 0 1
rlabel polysilicon 1647 -1533 1647 -1533 0 3
rlabel polysilicon 1654 -1527 1654 -1527 0 1
rlabel polysilicon 1654 -1533 1654 -1533 0 3
rlabel polysilicon 1661 -1527 1661 -1527 0 1
rlabel polysilicon 1661 -1533 1661 -1533 0 3
rlabel polysilicon 1668 -1527 1668 -1527 0 1
rlabel polysilicon 1668 -1533 1668 -1533 0 3
rlabel polysilicon 1675 -1527 1675 -1527 0 1
rlabel polysilicon 1675 -1533 1675 -1533 0 3
rlabel polysilicon 1682 -1527 1682 -1527 0 1
rlabel polysilicon 1682 -1533 1682 -1533 0 3
rlabel polysilicon 1689 -1527 1689 -1527 0 1
rlabel polysilicon 1689 -1533 1689 -1533 0 3
rlabel polysilicon 1696 -1527 1696 -1527 0 1
rlabel polysilicon 1696 -1533 1696 -1533 0 3
rlabel polysilicon 1703 -1527 1703 -1527 0 1
rlabel polysilicon 1703 -1533 1703 -1533 0 3
rlabel polysilicon 1710 -1527 1710 -1527 0 1
rlabel polysilicon 1710 -1533 1710 -1533 0 3
rlabel polysilicon 1717 -1527 1717 -1527 0 1
rlabel polysilicon 1717 -1533 1717 -1533 0 3
rlabel polysilicon 1724 -1527 1724 -1527 0 1
rlabel polysilicon 1724 -1533 1724 -1533 0 3
rlabel polysilicon 1731 -1527 1731 -1527 0 1
rlabel polysilicon 1731 -1533 1731 -1533 0 3
rlabel polysilicon 1738 -1527 1738 -1527 0 1
rlabel polysilicon 1738 -1533 1738 -1533 0 3
rlabel polysilicon 1745 -1527 1745 -1527 0 1
rlabel polysilicon 1745 -1533 1745 -1533 0 3
rlabel polysilicon 1752 -1527 1752 -1527 0 1
rlabel polysilicon 1752 -1533 1752 -1533 0 3
rlabel polysilicon 1759 -1527 1759 -1527 0 1
rlabel polysilicon 1759 -1533 1759 -1533 0 3
rlabel polysilicon 1766 -1527 1766 -1527 0 1
rlabel polysilicon 1766 -1533 1766 -1533 0 3
rlabel polysilicon 1773 -1527 1773 -1527 0 1
rlabel polysilicon 1773 -1533 1773 -1533 0 3
rlabel polysilicon 1780 -1527 1780 -1527 0 1
rlabel polysilicon 1780 -1533 1780 -1533 0 3
rlabel polysilicon 1787 -1527 1787 -1527 0 1
rlabel polysilicon 1787 -1533 1787 -1533 0 3
rlabel polysilicon 1794 -1527 1794 -1527 0 1
rlabel polysilicon 1797 -1527 1797 -1527 0 2
rlabel polysilicon 1794 -1533 1794 -1533 0 3
rlabel polysilicon 1801 -1527 1801 -1527 0 1
rlabel polysilicon 1801 -1533 1801 -1533 0 3
rlabel polysilicon 1808 -1527 1808 -1527 0 1
rlabel polysilicon 1808 -1533 1808 -1533 0 3
rlabel polysilicon 1815 -1527 1815 -1527 0 1
rlabel polysilicon 1815 -1533 1815 -1533 0 3
rlabel polysilicon 1822 -1527 1822 -1527 0 1
rlabel polysilicon 1822 -1533 1822 -1533 0 3
rlabel polysilicon 1829 -1527 1829 -1527 0 1
rlabel polysilicon 1829 -1533 1829 -1533 0 3
rlabel polysilicon 1836 -1527 1836 -1527 0 1
rlabel polysilicon 1836 -1533 1836 -1533 0 3
rlabel polysilicon 1843 -1527 1843 -1527 0 1
rlabel polysilicon 1843 -1533 1843 -1533 0 3
rlabel polysilicon 1850 -1527 1850 -1527 0 1
rlabel polysilicon 1850 -1533 1850 -1533 0 3
rlabel polysilicon 1857 -1527 1857 -1527 0 1
rlabel polysilicon 1857 -1533 1857 -1533 0 3
rlabel polysilicon 1864 -1527 1864 -1527 0 1
rlabel polysilicon 1864 -1533 1864 -1533 0 3
rlabel polysilicon 1871 -1527 1871 -1527 0 1
rlabel polysilicon 1871 -1533 1871 -1533 0 3
rlabel polysilicon 1878 -1527 1878 -1527 0 1
rlabel polysilicon 1878 -1533 1878 -1533 0 3
rlabel polysilicon 1885 -1527 1885 -1527 0 1
rlabel polysilicon 1885 -1533 1885 -1533 0 3
rlabel polysilicon 1892 -1527 1892 -1527 0 1
rlabel polysilicon 1892 -1533 1892 -1533 0 3
rlabel polysilicon 1899 -1527 1899 -1527 0 1
rlabel polysilicon 1899 -1533 1899 -1533 0 3
rlabel polysilicon 1906 -1527 1906 -1527 0 1
rlabel polysilicon 1906 -1533 1906 -1533 0 3
rlabel polysilicon 1913 -1527 1913 -1527 0 1
rlabel polysilicon 1913 -1533 1913 -1533 0 3
rlabel polysilicon 1920 -1527 1920 -1527 0 1
rlabel polysilicon 1920 -1533 1920 -1533 0 3
rlabel polysilicon 1927 -1527 1927 -1527 0 1
rlabel polysilicon 1927 -1533 1927 -1533 0 3
rlabel polysilicon 1934 -1527 1934 -1527 0 1
rlabel polysilicon 1934 -1533 1934 -1533 0 3
rlabel polysilicon 1941 -1527 1941 -1527 0 1
rlabel polysilicon 1941 -1533 1941 -1533 0 3
rlabel polysilicon 1948 -1527 1948 -1527 0 1
rlabel polysilicon 1948 -1533 1948 -1533 0 3
rlabel polysilicon 1955 -1527 1955 -1527 0 1
rlabel polysilicon 1955 -1533 1955 -1533 0 3
rlabel polysilicon 1962 -1527 1962 -1527 0 1
rlabel polysilicon 1962 -1533 1962 -1533 0 3
rlabel polysilicon 1969 -1527 1969 -1527 0 1
rlabel polysilicon 1969 -1533 1969 -1533 0 3
rlabel polysilicon 1976 -1527 1976 -1527 0 1
rlabel polysilicon 1976 -1533 1976 -1533 0 3
rlabel polysilicon 1983 -1527 1983 -1527 0 1
rlabel polysilicon 1983 -1533 1983 -1533 0 3
rlabel polysilicon 1990 -1527 1990 -1527 0 1
rlabel polysilicon 1990 -1533 1990 -1533 0 3
rlabel polysilicon 1997 -1527 1997 -1527 0 1
rlabel polysilicon 1997 -1533 1997 -1533 0 3
rlabel polysilicon 2004 -1527 2004 -1527 0 1
rlabel polysilicon 2004 -1533 2004 -1533 0 3
rlabel polysilicon 2011 -1527 2011 -1527 0 1
rlabel polysilicon 2011 -1533 2011 -1533 0 3
rlabel polysilicon 2018 -1527 2018 -1527 0 1
rlabel polysilicon 2018 -1533 2018 -1533 0 3
rlabel polysilicon 2025 -1527 2025 -1527 0 1
rlabel polysilicon 2025 -1533 2025 -1533 0 3
rlabel polysilicon 2032 -1527 2032 -1527 0 1
rlabel polysilicon 2032 -1533 2032 -1533 0 3
rlabel polysilicon 2039 -1527 2039 -1527 0 1
rlabel polysilicon 2039 -1533 2039 -1533 0 3
rlabel polysilicon 2046 -1527 2046 -1527 0 1
rlabel polysilicon 2046 -1533 2046 -1533 0 3
rlabel polysilicon 2053 -1527 2053 -1527 0 1
rlabel polysilicon 2053 -1533 2053 -1533 0 3
rlabel polysilicon 2060 -1527 2060 -1527 0 1
rlabel polysilicon 2060 -1533 2060 -1533 0 3
rlabel polysilicon 2067 -1527 2067 -1527 0 1
rlabel polysilicon 2067 -1533 2067 -1533 0 3
rlabel polysilicon 2074 -1527 2074 -1527 0 1
rlabel polysilicon 2074 -1533 2074 -1533 0 3
rlabel polysilicon 2081 -1527 2081 -1527 0 1
rlabel polysilicon 2081 -1533 2081 -1533 0 3
rlabel polysilicon 2088 -1527 2088 -1527 0 1
rlabel polysilicon 2088 -1533 2088 -1533 0 3
rlabel polysilicon 2095 -1527 2095 -1527 0 1
rlabel polysilicon 2095 -1533 2095 -1533 0 3
rlabel polysilicon 2102 -1527 2102 -1527 0 1
rlabel polysilicon 2102 -1533 2102 -1533 0 3
rlabel polysilicon 2109 -1527 2109 -1527 0 1
rlabel polysilicon 2109 -1533 2109 -1533 0 3
rlabel polysilicon 2116 -1527 2116 -1527 0 1
rlabel polysilicon 2116 -1533 2116 -1533 0 3
rlabel polysilicon 2123 -1527 2123 -1527 0 1
rlabel polysilicon 2123 -1533 2123 -1533 0 3
rlabel polysilicon 2130 -1527 2130 -1527 0 1
rlabel polysilicon 2130 -1533 2130 -1533 0 3
rlabel polysilicon 2137 -1527 2137 -1527 0 1
rlabel polysilicon 2137 -1533 2137 -1533 0 3
rlabel polysilicon 2144 -1527 2144 -1527 0 1
rlabel polysilicon 2144 -1533 2144 -1533 0 3
rlabel polysilicon 2151 -1527 2151 -1527 0 1
rlabel polysilicon 2151 -1533 2151 -1533 0 3
rlabel polysilicon 2158 -1527 2158 -1527 0 1
rlabel polysilicon 2158 -1533 2158 -1533 0 3
rlabel polysilicon 2165 -1527 2165 -1527 0 1
rlabel polysilicon 2165 -1533 2165 -1533 0 3
rlabel polysilicon 2172 -1527 2172 -1527 0 1
rlabel polysilicon 2172 -1533 2172 -1533 0 3
rlabel polysilicon 2179 -1527 2179 -1527 0 1
rlabel polysilicon 2179 -1533 2179 -1533 0 3
rlabel polysilicon 2186 -1527 2186 -1527 0 1
rlabel polysilicon 2186 -1533 2186 -1533 0 3
rlabel polysilicon 2193 -1527 2193 -1527 0 1
rlabel polysilicon 2193 -1533 2193 -1533 0 3
rlabel polysilicon 2200 -1527 2200 -1527 0 1
rlabel polysilicon 2200 -1533 2200 -1533 0 3
rlabel polysilicon 2207 -1527 2207 -1527 0 1
rlabel polysilicon 2207 -1533 2207 -1533 0 3
rlabel polysilicon 2214 -1527 2214 -1527 0 1
rlabel polysilicon 2214 -1533 2214 -1533 0 3
rlabel polysilicon 2221 -1527 2221 -1527 0 1
rlabel polysilicon 2221 -1533 2221 -1533 0 3
rlabel polysilicon 2228 -1527 2228 -1527 0 1
rlabel polysilicon 2228 -1533 2228 -1533 0 3
rlabel polysilicon 2235 -1527 2235 -1527 0 1
rlabel polysilicon 2235 -1533 2235 -1533 0 3
rlabel polysilicon 2242 -1527 2242 -1527 0 1
rlabel polysilicon 2242 -1533 2242 -1533 0 3
rlabel polysilicon 2249 -1527 2249 -1527 0 1
rlabel polysilicon 2249 -1533 2249 -1533 0 3
rlabel polysilicon 2256 -1527 2256 -1527 0 1
rlabel polysilicon 2256 -1533 2256 -1533 0 3
rlabel polysilicon 2263 -1527 2263 -1527 0 1
rlabel polysilicon 2263 -1533 2263 -1533 0 3
rlabel polysilicon 2270 -1527 2270 -1527 0 1
rlabel polysilicon 2270 -1533 2270 -1533 0 3
rlabel polysilicon 2277 -1527 2277 -1527 0 1
rlabel polysilicon 2277 -1533 2277 -1533 0 3
rlabel polysilicon 2284 -1527 2284 -1527 0 1
rlabel polysilicon 2284 -1533 2284 -1533 0 3
rlabel polysilicon 2291 -1527 2291 -1527 0 1
rlabel polysilicon 2291 -1533 2291 -1533 0 3
rlabel polysilicon 2298 -1527 2298 -1527 0 1
rlabel polysilicon 2298 -1533 2298 -1533 0 3
rlabel polysilicon 2305 -1527 2305 -1527 0 1
rlabel polysilicon 2305 -1533 2305 -1533 0 3
rlabel polysilicon 2312 -1527 2312 -1527 0 1
rlabel polysilicon 2312 -1533 2312 -1533 0 3
rlabel polysilicon 2319 -1527 2319 -1527 0 1
rlabel polysilicon 2319 -1533 2319 -1533 0 3
rlabel polysilicon 2326 -1527 2326 -1527 0 1
rlabel polysilicon 2326 -1533 2326 -1533 0 3
rlabel polysilicon 2333 -1527 2333 -1527 0 1
rlabel polysilicon 2333 -1533 2333 -1533 0 3
rlabel polysilicon 2340 -1527 2340 -1527 0 1
rlabel polysilicon 2340 -1533 2340 -1533 0 3
rlabel polysilicon 2347 -1527 2347 -1527 0 1
rlabel polysilicon 2347 -1533 2347 -1533 0 3
rlabel polysilicon 2354 -1527 2354 -1527 0 1
rlabel polysilicon 2354 -1533 2354 -1533 0 3
rlabel polysilicon 2361 -1527 2361 -1527 0 1
rlabel polysilicon 2361 -1533 2361 -1533 0 3
rlabel polysilicon 2368 -1527 2368 -1527 0 1
rlabel polysilicon 2368 -1533 2368 -1533 0 3
rlabel polysilicon 2375 -1527 2375 -1527 0 1
rlabel polysilicon 2375 -1533 2375 -1533 0 3
rlabel polysilicon 2382 -1527 2382 -1527 0 1
rlabel polysilicon 2382 -1533 2382 -1533 0 3
rlabel polysilicon 2389 -1527 2389 -1527 0 1
rlabel polysilicon 2389 -1533 2389 -1533 0 3
rlabel polysilicon 2396 -1527 2396 -1527 0 1
rlabel polysilicon 2396 -1533 2396 -1533 0 3
rlabel polysilicon 2403 -1527 2403 -1527 0 1
rlabel polysilicon 2403 -1533 2403 -1533 0 3
rlabel polysilicon 2410 -1527 2410 -1527 0 1
rlabel polysilicon 2410 -1533 2410 -1533 0 3
rlabel polysilicon 2417 -1527 2417 -1527 0 1
rlabel polysilicon 2417 -1533 2417 -1533 0 3
rlabel polysilicon 2424 -1527 2424 -1527 0 1
rlabel polysilicon 2424 -1533 2424 -1533 0 3
rlabel polysilicon 2431 -1527 2431 -1527 0 1
rlabel polysilicon 2431 -1533 2431 -1533 0 3
rlabel polysilicon 2438 -1527 2438 -1527 0 1
rlabel polysilicon 2438 -1533 2438 -1533 0 3
rlabel polysilicon 2445 -1527 2445 -1527 0 1
rlabel polysilicon 2445 -1533 2445 -1533 0 3
rlabel polysilicon 2452 -1527 2452 -1527 0 1
rlabel polysilicon 2452 -1533 2452 -1533 0 3
rlabel polysilicon 2459 -1527 2459 -1527 0 1
rlabel polysilicon 2459 -1533 2459 -1533 0 3
rlabel polysilicon 2466 -1527 2466 -1527 0 1
rlabel polysilicon 2466 -1533 2466 -1533 0 3
rlabel polysilicon 2473 -1527 2473 -1527 0 1
rlabel polysilicon 2473 -1533 2473 -1533 0 3
rlabel polysilicon 2480 -1527 2480 -1527 0 1
rlabel polysilicon 2480 -1533 2480 -1533 0 3
rlabel polysilicon 2487 -1527 2487 -1527 0 1
rlabel polysilicon 2487 -1533 2487 -1533 0 3
rlabel polysilicon 2494 -1527 2494 -1527 0 1
rlabel polysilicon 2494 -1533 2494 -1533 0 3
rlabel polysilicon 2501 -1527 2501 -1527 0 1
rlabel polysilicon 2501 -1533 2501 -1533 0 3
rlabel polysilicon 2508 -1527 2508 -1527 0 1
rlabel polysilicon 2508 -1533 2508 -1533 0 3
rlabel polysilicon 2515 -1527 2515 -1527 0 1
rlabel polysilicon 2515 -1533 2515 -1533 0 3
rlabel polysilicon 2522 -1527 2522 -1527 0 1
rlabel polysilicon 2522 -1533 2522 -1533 0 3
rlabel polysilicon 2529 -1527 2529 -1527 0 1
rlabel polysilicon 2529 -1533 2529 -1533 0 3
rlabel polysilicon 2536 -1527 2536 -1527 0 1
rlabel polysilicon 2536 -1533 2536 -1533 0 3
rlabel polysilicon 2543 -1527 2543 -1527 0 1
rlabel polysilicon 2543 -1533 2543 -1533 0 3
rlabel polysilicon 2550 -1527 2550 -1527 0 1
rlabel polysilicon 2550 -1533 2550 -1533 0 3
rlabel polysilicon 2557 -1527 2557 -1527 0 1
rlabel polysilicon 2557 -1533 2557 -1533 0 3
rlabel polysilicon 16 -1700 16 -1700 0 1
rlabel polysilicon 16 -1706 16 -1706 0 3
rlabel polysilicon 23 -1700 23 -1700 0 1
rlabel polysilicon 23 -1706 23 -1706 0 3
rlabel polysilicon 30 -1700 30 -1700 0 1
rlabel polysilicon 30 -1706 30 -1706 0 3
rlabel polysilicon 37 -1700 37 -1700 0 1
rlabel polysilicon 37 -1706 37 -1706 0 3
rlabel polysilicon 44 -1700 44 -1700 0 1
rlabel polysilicon 44 -1706 44 -1706 0 3
rlabel polysilicon 51 -1700 51 -1700 0 1
rlabel polysilicon 51 -1706 51 -1706 0 3
rlabel polysilicon 58 -1700 58 -1700 0 1
rlabel polysilicon 58 -1706 58 -1706 0 3
rlabel polysilicon 65 -1700 65 -1700 0 1
rlabel polysilicon 65 -1706 65 -1706 0 3
rlabel polysilicon 72 -1700 72 -1700 0 1
rlabel polysilicon 72 -1706 72 -1706 0 3
rlabel polysilicon 79 -1700 79 -1700 0 1
rlabel polysilicon 79 -1706 79 -1706 0 3
rlabel polysilicon 86 -1700 86 -1700 0 1
rlabel polysilicon 86 -1706 86 -1706 0 3
rlabel polysilicon 93 -1700 93 -1700 0 1
rlabel polysilicon 96 -1700 96 -1700 0 2
rlabel polysilicon 93 -1706 93 -1706 0 3
rlabel polysilicon 96 -1706 96 -1706 0 4
rlabel polysilicon 100 -1700 100 -1700 0 1
rlabel polysilicon 100 -1706 100 -1706 0 3
rlabel polysilicon 107 -1700 107 -1700 0 1
rlabel polysilicon 107 -1706 107 -1706 0 3
rlabel polysilicon 114 -1700 114 -1700 0 1
rlabel polysilicon 114 -1706 114 -1706 0 3
rlabel polysilicon 121 -1700 121 -1700 0 1
rlabel polysilicon 121 -1706 121 -1706 0 3
rlabel polysilicon 128 -1700 128 -1700 0 1
rlabel polysilicon 128 -1706 128 -1706 0 3
rlabel polysilicon 135 -1700 135 -1700 0 1
rlabel polysilicon 135 -1706 135 -1706 0 3
rlabel polysilicon 142 -1700 142 -1700 0 1
rlabel polysilicon 142 -1706 142 -1706 0 3
rlabel polysilicon 149 -1700 149 -1700 0 1
rlabel polysilicon 149 -1706 149 -1706 0 3
rlabel polysilicon 156 -1700 156 -1700 0 1
rlabel polysilicon 156 -1706 156 -1706 0 3
rlabel polysilicon 163 -1700 163 -1700 0 1
rlabel polysilicon 163 -1706 163 -1706 0 3
rlabel polysilicon 170 -1700 170 -1700 0 1
rlabel polysilicon 170 -1706 170 -1706 0 3
rlabel polysilicon 180 -1700 180 -1700 0 2
rlabel polysilicon 177 -1706 177 -1706 0 3
rlabel polysilicon 180 -1706 180 -1706 0 4
rlabel polysilicon 184 -1700 184 -1700 0 1
rlabel polysilicon 184 -1706 184 -1706 0 3
rlabel polysilicon 191 -1700 191 -1700 0 1
rlabel polysilicon 194 -1700 194 -1700 0 2
rlabel polysilicon 191 -1706 191 -1706 0 3
rlabel polysilicon 194 -1706 194 -1706 0 4
rlabel polysilicon 198 -1700 198 -1700 0 1
rlabel polysilicon 198 -1706 198 -1706 0 3
rlabel polysilicon 205 -1700 205 -1700 0 1
rlabel polysilicon 205 -1706 205 -1706 0 3
rlabel polysilicon 212 -1700 212 -1700 0 1
rlabel polysilicon 212 -1706 212 -1706 0 3
rlabel polysilicon 215 -1706 215 -1706 0 4
rlabel polysilicon 219 -1700 219 -1700 0 1
rlabel polysilicon 219 -1706 219 -1706 0 3
rlabel polysilicon 226 -1700 226 -1700 0 1
rlabel polysilicon 229 -1700 229 -1700 0 2
rlabel polysilicon 229 -1706 229 -1706 0 4
rlabel polysilicon 233 -1700 233 -1700 0 1
rlabel polysilicon 233 -1706 233 -1706 0 3
rlabel polysilicon 240 -1700 240 -1700 0 1
rlabel polysilicon 240 -1706 240 -1706 0 3
rlabel polysilicon 250 -1700 250 -1700 0 2
rlabel polysilicon 247 -1706 247 -1706 0 3
rlabel polysilicon 254 -1700 254 -1700 0 1
rlabel polysilicon 254 -1706 254 -1706 0 3
rlabel polysilicon 261 -1700 261 -1700 0 1
rlabel polysilicon 261 -1706 261 -1706 0 3
rlabel polysilicon 268 -1700 268 -1700 0 1
rlabel polysilicon 268 -1706 268 -1706 0 3
rlabel polysilicon 275 -1700 275 -1700 0 1
rlabel polysilicon 275 -1706 275 -1706 0 3
rlabel polysilicon 282 -1700 282 -1700 0 1
rlabel polysilicon 282 -1706 282 -1706 0 3
rlabel polysilicon 289 -1700 289 -1700 0 1
rlabel polysilicon 289 -1706 289 -1706 0 3
rlabel polysilicon 296 -1700 296 -1700 0 1
rlabel polysilicon 296 -1706 296 -1706 0 3
rlabel polysilicon 303 -1700 303 -1700 0 1
rlabel polysilicon 303 -1706 303 -1706 0 3
rlabel polysilicon 310 -1700 310 -1700 0 1
rlabel polysilicon 310 -1706 310 -1706 0 3
rlabel polysilicon 317 -1700 317 -1700 0 1
rlabel polysilicon 317 -1706 317 -1706 0 3
rlabel polysilicon 324 -1700 324 -1700 0 1
rlabel polysilicon 324 -1706 324 -1706 0 3
rlabel polysilicon 331 -1700 331 -1700 0 1
rlabel polysilicon 331 -1706 331 -1706 0 3
rlabel polysilicon 338 -1700 338 -1700 0 1
rlabel polysilicon 338 -1706 338 -1706 0 3
rlabel polysilicon 345 -1700 345 -1700 0 1
rlabel polysilicon 345 -1706 345 -1706 0 3
rlabel polysilicon 352 -1700 352 -1700 0 1
rlabel polysilicon 352 -1706 352 -1706 0 3
rlabel polysilicon 359 -1700 359 -1700 0 1
rlabel polysilicon 359 -1706 359 -1706 0 3
rlabel polysilicon 366 -1700 366 -1700 0 1
rlabel polysilicon 366 -1706 366 -1706 0 3
rlabel polysilicon 373 -1700 373 -1700 0 1
rlabel polysilicon 373 -1706 373 -1706 0 3
rlabel polysilicon 380 -1700 380 -1700 0 1
rlabel polysilicon 380 -1706 380 -1706 0 3
rlabel polysilicon 387 -1700 387 -1700 0 1
rlabel polysilicon 387 -1706 387 -1706 0 3
rlabel polysilicon 394 -1700 394 -1700 0 1
rlabel polysilicon 394 -1706 394 -1706 0 3
rlabel polysilicon 401 -1700 401 -1700 0 1
rlabel polysilicon 401 -1706 401 -1706 0 3
rlabel polysilicon 408 -1700 408 -1700 0 1
rlabel polysilicon 408 -1706 408 -1706 0 3
rlabel polysilicon 415 -1700 415 -1700 0 1
rlabel polysilicon 415 -1706 415 -1706 0 3
rlabel polysilicon 422 -1700 422 -1700 0 1
rlabel polysilicon 422 -1706 422 -1706 0 3
rlabel polysilicon 429 -1700 429 -1700 0 1
rlabel polysilicon 429 -1706 429 -1706 0 3
rlabel polysilicon 436 -1700 436 -1700 0 1
rlabel polysilicon 436 -1706 436 -1706 0 3
rlabel polysilicon 443 -1700 443 -1700 0 1
rlabel polysilicon 443 -1706 443 -1706 0 3
rlabel polysilicon 450 -1700 450 -1700 0 1
rlabel polysilicon 453 -1700 453 -1700 0 2
rlabel polysilicon 453 -1706 453 -1706 0 4
rlabel polysilicon 457 -1700 457 -1700 0 1
rlabel polysilicon 460 -1700 460 -1700 0 2
rlabel polysilicon 460 -1706 460 -1706 0 4
rlabel polysilicon 464 -1700 464 -1700 0 1
rlabel polysilicon 464 -1706 464 -1706 0 3
rlabel polysilicon 471 -1700 471 -1700 0 1
rlabel polysilicon 471 -1706 471 -1706 0 3
rlabel polysilicon 478 -1700 478 -1700 0 1
rlabel polysilicon 481 -1700 481 -1700 0 2
rlabel polysilicon 478 -1706 478 -1706 0 3
rlabel polysilicon 481 -1706 481 -1706 0 4
rlabel polysilicon 485 -1700 485 -1700 0 1
rlabel polysilicon 485 -1706 485 -1706 0 3
rlabel polysilicon 492 -1700 492 -1700 0 1
rlabel polysilicon 492 -1706 492 -1706 0 3
rlabel polysilicon 499 -1700 499 -1700 0 1
rlabel polysilicon 499 -1706 499 -1706 0 3
rlabel polysilicon 506 -1700 506 -1700 0 1
rlabel polysilicon 506 -1706 506 -1706 0 3
rlabel polysilicon 513 -1700 513 -1700 0 1
rlabel polysilicon 513 -1706 513 -1706 0 3
rlabel polysilicon 520 -1700 520 -1700 0 1
rlabel polysilicon 520 -1706 520 -1706 0 3
rlabel polysilicon 527 -1700 527 -1700 0 1
rlabel polysilicon 527 -1706 527 -1706 0 3
rlabel polysilicon 534 -1700 534 -1700 0 1
rlabel polysilicon 534 -1706 534 -1706 0 3
rlabel polysilicon 541 -1700 541 -1700 0 1
rlabel polysilicon 541 -1706 541 -1706 0 3
rlabel polysilicon 548 -1700 548 -1700 0 1
rlabel polysilicon 548 -1706 548 -1706 0 3
rlabel polysilicon 555 -1700 555 -1700 0 1
rlabel polysilicon 555 -1706 555 -1706 0 3
rlabel polysilicon 562 -1700 562 -1700 0 1
rlabel polysilicon 562 -1706 562 -1706 0 3
rlabel polysilicon 569 -1700 569 -1700 0 1
rlabel polysilicon 569 -1706 569 -1706 0 3
rlabel polysilicon 576 -1706 576 -1706 0 3
rlabel polysilicon 579 -1706 579 -1706 0 4
rlabel polysilicon 583 -1700 583 -1700 0 1
rlabel polysilicon 583 -1706 583 -1706 0 3
rlabel polysilicon 590 -1700 590 -1700 0 1
rlabel polysilicon 590 -1706 590 -1706 0 3
rlabel polysilicon 597 -1700 597 -1700 0 1
rlabel polysilicon 597 -1706 597 -1706 0 3
rlabel polysilicon 604 -1700 604 -1700 0 1
rlabel polysilicon 604 -1706 604 -1706 0 3
rlabel polysilicon 611 -1700 611 -1700 0 1
rlabel polysilicon 611 -1706 611 -1706 0 3
rlabel polysilicon 618 -1700 618 -1700 0 1
rlabel polysilicon 618 -1706 618 -1706 0 3
rlabel polysilicon 625 -1700 625 -1700 0 1
rlabel polysilicon 625 -1706 625 -1706 0 3
rlabel polysilicon 632 -1700 632 -1700 0 1
rlabel polysilicon 632 -1706 632 -1706 0 3
rlabel polysilicon 639 -1700 639 -1700 0 1
rlabel polysilicon 642 -1700 642 -1700 0 2
rlabel polysilicon 642 -1706 642 -1706 0 4
rlabel polysilicon 646 -1700 646 -1700 0 1
rlabel polysilicon 646 -1706 646 -1706 0 3
rlabel polysilicon 653 -1700 653 -1700 0 1
rlabel polysilicon 653 -1706 653 -1706 0 3
rlabel polysilicon 660 -1700 660 -1700 0 1
rlabel polysilicon 660 -1706 660 -1706 0 3
rlabel polysilicon 667 -1700 667 -1700 0 1
rlabel polysilicon 667 -1706 667 -1706 0 3
rlabel polysilicon 674 -1700 674 -1700 0 1
rlabel polysilicon 674 -1706 674 -1706 0 3
rlabel polysilicon 681 -1700 681 -1700 0 1
rlabel polysilicon 681 -1706 681 -1706 0 3
rlabel polysilicon 688 -1700 688 -1700 0 1
rlabel polysilicon 688 -1706 688 -1706 0 3
rlabel polysilicon 695 -1700 695 -1700 0 1
rlabel polysilicon 698 -1700 698 -1700 0 2
rlabel polysilicon 695 -1706 695 -1706 0 3
rlabel polysilicon 698 -1706 698 -1706 0 4
rlabel polysilicon 702 -1700 702 -1700 0 1
rlabel polysilicon 702 -1706 702 -1706 0 3
rlabel polysilicon 709 -1700 709 -1700 0 1
rlabel polysilicon 709 -1706 709 -1706 0 3
rlabel polysilicon 716 -1700 716 -1700 0 1
rlabel polysilicon 719 -1700 719 -1700 0 2
rlabel polysilicon 716 -1706 716 -1706 0 3
rlabel polysilicon 719 -1706 719 -1706 0 4
rlabel polysilicon 723 -1700 723 -1700 0 1
rlabel polysilicon 723 -1706 723 -1706 0 3
rlabel polysilicon 730 -1700 730 -1700 0 1
rlabel polysilicon 730 -1706 730 -1706 0 3
rlabel polysilicon 737 -1700 737 -1700 0 1
rlabel polysilicon 737 -1706 737 -1706 0 3
rlabel polysilicon 744 -1700 744 -1700 0 1
rlabel polysilicon 744 -1706 744 -1706 0 3
rlabel polysilicon 751 -1700 751 -1700 0 1
rlabel polysilicon 751 -1706 751 -1706 0 3
rlabel polysilicon 758 -1700 758 -1700 0 1
rlabel polysilicon 758 -1706 758 -1706 0 3
rlabel polysilicon 765 -1700 765 -1700 0 1
rlabel polysilicon 765 -1706 765 -1706 0 3
rlabel polysilicon 772 -1700 772 -1700 0 1
rlabel polysilicon 772 -1706 772 -1706 0 3
rlabel polysilicon 779 -1700 779 -1700 0 1
rlabel polysilicon 779 -1706 779 -1706 0 3
rlabel polysilicon 786 -1700 786 -1700 0 1
rlabel polysilicon 786 -1706 786 -1706 0 3
rlabel polysilicon 793 -1700 793 -1700 0 1
rlabel polysilicon 793 -1706 793 -1706 0 3
rlabel polysilicon 800 -1700 800 -1700 0 1
rlabel polysilicon 800 -1706 800 -1706 0 3
rlabel polysilicon 807 -1700 807 -1700 0 1
rlabel polysilicon 807 -1706 807 -1706 0 3
rlabel polysilicon 814 -1700 814 -1700 0 1
rlabel polysilicon 814 -1706 814 -1706 0 3
rlabel polysilicon 821 -1700 821 -1700 0 1
rlabel polysilicon 821 -1706 821 -1706 0 3
rlabel polysilicon 828 -1700 828 -1700 0 1
rlabel polysilicon 828 -1706 828 -1706 0 3
rlabel polysilicon 835 -1700 835 -1700 0 1
rlabel polysilicon 835 -1706 835 -1706 0 3
rlabel polysilicon 842 -1700 842 -1700 0 1
rlabel polysilicon 842 -1706 842 -1706 0 3
rlabel polysilicon 849 -1700 849 -1700 0 1
rlabel polysilicon 849 -1706 849 -1706 0 3
rlabel polysilicon 856 -1700 856 -1700 0 1
rlabel polysilicon 859 -1700 859 -1700 0 2
rlabel polysilicon 856 -1706 856 -1706 0 3
rlabel polysilicon 859 -1706 859 -1706 0 4
rlabel polysilicon 863 -1700 863 -1700 0 1
rlabel polysilicon 863 -1706 863 -1706 0 3
rlabel polysilicon 870 -1700 870 -1700 0 1
rlabel polysilicon 870 -1706 870 -1706 0 3
rlabel polysilicon 877 -1700 877 -1700 0 1
rlabel polysilicon 877 -1706 877 -1706 0 3
rlabel polysilicon 884 -1700 884 -1700 0 1
rlabel polysilicon 884 -1706 884 -1706 0 3
rlabel polysilicon 891 -1700 891 -1700 0 1
rlabel polysilicon 891 -1706 891 -1706 0 3
rlabel polysilicon 898 -1700 898 -1700 0 1
rlabel polysilicon 898 -1706 898 -1706 0 3
rlabel polysilicon 905 -1700 905 -1700 0 1
rlabel polysilicon 905 -1706 905 -1706 0 3
rlabel polysilicon 912 -1700 912 -1700 0 1
rlabel polysilicon 912 -1706 912 -1706 0 3
rlabel polysilicon 919 -1700 919 -1700 0 1
rlabel polysilicon 919 -1706 919 -1706 0 3
rlabel polysilicon 926 -1700 926 -1700 0 1
rlabel polysilicon 926 -1706 926 -1706 0 3
rlabel polysilicon 933 -1700 933 -1700 0 1
rlabel polysilicon 936 -1700 936 -1700 0 2
rlabel polysilicon 933 -1706 933 -1706 0 3
rlabel polysilicon 936 -1706 936 -1706 0 4
rlabel polysilicon 940 -1700 940 -1700 0 1
rlabel polysilicon 940 -1706 940 -1706 0 3
rlabel polysilicon 947 -1700 947 -1700 0 1
rlabel polysilicon 947 -1706 947 -1706 0 3
rlabel polysilicon 954 -1700 954 -1700 0 1
rlabel polysilicon 954 -1706 954 -1706 0 3
rlabel polysilicon 961 -1700 961 -1700 0 1
rlabel polysilicon 961 -1706 961 -1706 0 3
rlabel polysilicon 968 -1700 968 -1700 0 1
rlabel polysilicon 968 -1706 968 -1706 0 3
rlabel polysilicon 971 -1706 971 -1706 0 4
rlabel polysilicon 975 -1700 975 -1700 0 1
rlabel polysilicon 975 -1706 975 -1706 0 3
rlabel polysilicon 982 -1700 982 -1700 0 1
rlabel polysilicon 982 -1706 982 -1706 0 3
rlabel polysilicon 989 -1700 989 -1700 0 1
rlabel polysilicon 989 -1706 989 -1706 0 3
rlabel polysilicon 996 -1700 996 -1700 0 1
rlabel polysilicon 996 -1706 996 -1706 0 3
rlabel polysilicon 1003 -1700 1003 -1700 0 1
rlabel polysilicon 1003 -1706 1003 -1706 0 3
rlabel polysilicon 1010 -1700 1010 -1700 0 1
rlabel polysilicon 1010 -1706 1010 -1706 0 3
rlabel polysilicon 1017 -1700 1017 -1700 0 1
rlabel polysilicon 1020 -1700 1020 -1700 0 2
rlabel polysilicon 1017 -1706 1017 -1706 0 3
rlabel polysilicon 1020 -1706 1020 -1706 0 4
rlabel polysilicon 1024 -1700 1024 -1700 0 1
rlabel polysilicon 1024 -1706 1024 -1706 0 3
rlabel polysilicon 1034 -1700 1034 -1700 0 2
rlabel polysilicon 1031 -1706 1031 -1706 0 3
rlabel polysilicon 1038 -1700 1038 -1700 0 1
rlabel polysilicon 1038 -1706 1038 -1706 0 3
rlabel polysilicon 1045 -1700 1045 -1700 0 1
rlabel polysilicon 1045 -1706 1045 -1706 0 3
rlabel polysilicon 1052 -1700 1052 -1700 0 1
rlabel polysilicon 1052 -1706 1052 -1706 0 3
rlabel polysilicon 1059 -1700 1059 -1700 0 1
rlabel polysilicon 1059 -1706 1059 -1706 0 3
rlabel polysilicon 1066 -1700 1066 -1700 0 1
rlabel polysilicon 1066 -1706 1066 -1706 0 3
rlabel polysilicon 1073 -1700 1073 -1700 0 1
rlabel polysilicon 1076 -1700 1076 -1700 0 2
rlabel polysilicon 1073 -1706 1073 -1706 0 3
rlabel polysilicon 1076 -1706 1076 -1706 0 4
rlabel polysilicon 1080 -1700 1080 -1700 0 1
rlabel polysilicon 1080 -1706 1080 -1706 0 3
rlabel polysilicon 1087 -1700 1087 -1700 0 1
rlabel polysilicon 1087 -1706 1087 -1706 0 3
rlabel polysilicon 1094 -1700 1094 -1700 0 1
rlabel polysilicon 1094 -1706 1094 -1706 0 3
rlabel polysilicon 1101 -1700 1101 -1700 0 1
rlabel polysilicon 1101 -1706 1101 -1706 0 3
rlabel polysilicon 1108 -1700 1108 -1700 0 1
rlabel polysilicon 1111 -1700 1111 -1700 0 2
rlabel polysilicon 1108 -1706 1108 -1706 0 3
rlabel polysilicon 1111 -1706 1111 -1706 0 4
rlabel polysilicon 1115 -1700 1115 -1700 0 1
rlabel polysilicon 1115 -1706 1115 -1706 0 3
rlabel polysilicon 1122 -1700 1122 -1700 0 1
rlabel polysilicon 1122 -1706 1122 -1706 0 3
rlabel polysilicon 1129 -1700 1129 -1700 0 1
rlabel polysilicon 1129 -1706 1129 -1706 0 3
rlabel polysilicon 1136 -1700 1136 -1700 0 1
rlabel polysilicon 1136 -1706 1136 -1706 0 3
rlabel polysilicon 1143 -1700 1143 -1700 0 1
rlabel polysilicon 1143 -1706 1143 -1706 0 3
rlabel polysilicon 1153 -1700 1153 -1700 0 2
rlabel polysilicon 1150 -1706 1150 -1706 0 3
rlabel polysilicon 1153 -1706 1153 -1706 0 4
rlabel polysilicon 1157 -1700 1157 -1700 0 1
rlabel polysilicon 1157 -1706 1157 -1706 0 3
rlabel polysilicon 1164 -1700 1164 -1700 0 1
rlabel polysilicon 1164 -1706 1164 -1706 0 3
rlabel polysilicon 1171 -1700 1171 -1700 0 1
rlabel polysilicon 1171 -1706 1171 -1706 0 3
rlabel polysilicon 1178 -1700 1178 -1700 0 1
rlabel polysilicon 1178 -1706 1178 -1706 0 3
rlabel polysilicon 1185 -1700 1185 -1700 0 1
rlabel polysilicon 1185 -1706 1185 -1706 0 3
rlabel polysilicon 1192 -1700 1192 -1700 0 1
rlabel polysilicon 1192 -1706 1192 -1706 0 3
rlabel polysilicon 1199 -1700 1199 -1700 0 1
rlabel polysilicon 1199 -1706 1199 -1706 0 3
rlabel polysilicon 1206 -1700 1206 -1700 0 1
rlabel polysilicon 1206 -1706 1206 -1706 0 3
rlabel polysilicon 1213 -1700 1213 -1700 0 1
rlabel polysilicon 1213 -1706 1213 -1706 0 3
rlabel polysilicon 1220 -1700 1220 -1700 0 1
rlabel polysilicon 1220 -1706 1220 -1706 0 3
rlabel polysilicon 1227 -1700 1227 -1700 0 1
rlabel polysilicon 1227 -1706 1227 -1706 0 3
rlabel polysilicon 1234 -1700 1234 -1700 0 1
rlabel polysilicon 1234 -1706 1234 -1706 0 3
rlabel polysilicon 1241 -1700 1241 -1700 0 1
rlabel polysilicon 1241 -1706 1241 -1706 0 3
rlabel polysilicon 1248 -1700 1248 -1700 0 1
rlabel polysilicon 1248 -1706 1248 -1706 0 3
rlabel polysilicon 1255 -1700 1255 -1700 0 1
rlabel polysilicon 1255 -1706 1255 -1706 0 3
rlabel polysilicon 1262 -1700 1262 -1700 0 1
rlabel polysilicon 1265 -1700 1265 -1700 0 2
rlabel polysilicon 1262 -1706 1262 -1706 0 3
rlabel polysilicon 1265 -1706 1265 -1706 0 4
rlabel polysilicon 1269 -1700 1269 -1700 0 1
rlabel polysilicon 1269 -1706 1269 -1706 0 3
rlabel polysilicon 1276 -1700 1276 -1700 0 1
rlabel polysilicon 1276 -1706 1276 -1706 0 3
rlabel polysilicon 1279 -1706 1279 -1706 0 4
rlabel polysilicon 1283 -1700 1283 -1700 0 1
rlabel polysilicon 1283 -1706 1283 -1706 0 3
rlabel polysilicon 1290 -1700 1290 -1700 0 1
rlabel polysilicon 1293 -1700 1293 -1700 0 2
rlabel polysilicon 1290 -1706 1290 -1706 0 3
rlabel polysilicon 1293 -1706 1293 -1706 0 4
rlabel polysilicon 1297 -1700 1297 -1700 0 1
rlabel polysilicon 1297 -1706 1297 -1706 0 3
rlabel polysilicon 1304 -1700 1304 -1700 0 1
rlabel polysilicon 1304 -1706 1304 -1706 0 3
rlabel polysilicon 1311 -1700 1311 -1700 0 1
rlabel polysilicon 1311 -1706 1311 -1706 0 3
rlabel polysilicon 1318 -1700 1318 -1700 0 1
rlabel polysilicon 1318 -1706 1318 -1706 0 3
rlabel polysilicon 1325 -1700 1325 -1700 0 1
rlabel polysilicon 1325 -1706 1325 -1706 0 3
rlabel polysilicon 1332 -1700 1332 -1700 0 1
rlabel polysilicon 1332 -1706 1332 -1706 0 3
rlabel polysilicon 1339 -1700 1339 -1700 0 1
rlabel polysilicon 1339 -1706 1339 -1706 0 3
rlabel polysilicon 1346 -1700 1346 -1700 0 1
rlabel polysilicon 1346 -1706 1346 -1706 0 3
rlabel polysilicon 1353 -1700 1353 -1700 0 1
rlabel polysilicon 1353 -1706 1353 -1706 0 3
rlabel polysilicon 1360 -1700 1360 -1700 0 1
rlabel polysilicon 1363 -1700 1363 -1700 0 2
rlabel polysilicon 1360 -1706 1360 -1706 0 3
rlabel polysilicon 1363 -1706 1363 -1706 0 4
rlabel polysilicon 1367 -1700 1367 -1700 0 1
rlabel polysilicon 1367 -1706 1367 -1706 0 3
rlabel polysilicon 1374 -1700 1374 -1700 0 1
rlabel polysilicon 1374 -1706 1374 -1706 0 3
rlabel polysilicon 1381 -1700 1381 -1700 0 1
rlabel polysilicon 1381 -1706 1381 -1706 0 3
rlabel polysilicon 1388 -1700 1388 -1700 0 1
rlabel polysilicon 1388 -1706 1388 -1706 0 3
rlabel polysilicon 1395 -1700 1395 -1700 0 1
rlabel polysilicon 1395 -1706 1395 -1706 0 3
rlabel polysilicon 1402 -1700 1402 -1700 0 1
rlabel polysilicon 1402 -1706 1402 -1706 0 3
rlabel polysilicon 1409 -1700 1409 -1700 0 1
rlabel polysilicon 1409 -1706 1409 -1706 0 3
rlabel polysilicon 1416 -1700 1416 -1700 0 1
rlabel polysilicon 1416 -1706 1416 -1706 0 3
rlabel polysilicon 1423 -1700 1423 -1700 0 1
rlabel polysilicon 1423 -1706 1423 -1706 0 3
rlabel polysilicon 1430 -1700 1430 -1700 0 1
rlabel polysilicon 1430 -1706 1430 -1706 0 3
rlabel polysilicon 1437 -1700 1437 -1700 0 1
rlabel polysilicon 1440 -1700 1440 -1700 0 2
rlabel polysilicon 1437 -1706 1437 -1706 0 3
rlabel polysilicon 1440 -1706 1440 -1706 0 4
rlabel polysilicon 1444 -1700 1444 -1700 0 1
rlabel polysilicon 1444 -1706 1444 -1706 0 3
rlabel polysilicon 1451 -1700 1451 -1700 0 1
rlabel polysilicon 1451 -1706 1451 -1706 0 3
rlabel polysilicon 1458 -1700 1458 -1700 0 1
rlabel polysilicon 1458 -1706 1458 -1706 0 3
rlabel polysilicon 1465 -1700 1465 -1700 0 1
rlabel polysilicon 1468 -1700 1468 -1700 0 2
rlabel polysilicon 1465 -1706 1465 -1706 0 3
rlabel polysilicon 1468 -1706 1468 -1706 0 4
rlabel polysilicon 1472 -1700 1472 -1700 0 1
rlabel polysilicon 1472 -1706 1472 -1706 0 3
rlabel polysilicon 1479 -1700 1479 -1700 0 1
rlabel polysilicon 1479 -1706 1479 -1706 0 3
rlabel polysilicon 1486 -1700 1486 -1700 0 1
rlabel polysilicon 1486 -1706 1486 -1706 0 3
rlabel polysilicon 1493 -1700 1493 -1700 0 1
rlabel polysilicon 1496 -1700 1496 -1700 0 2
rlabel polysilicon 1493 -1706 1493 -1706 0 3
rlabel polysilicon 1496 -1706 1496 -1706 0 4
rlabel polysilicon 1500 -1700 1500 -1700 0 1
rlabel polysilicon 1500 -1706 1500 -1706 0 3
rlabel polysilicon 1507 -1700 1507 -1700 0 1
rlabel polysilicon 1510 -1700 1510 -1700 0 2
rlabel polysilicon 1507 -1706 1507 -1706 0 3
rlabel polysilicon 1510 -1706 1510 -1706 0 4
rlabel polysilicon 1514 -1700 1514 -1700 0 1
rlabel polysilicon 1514 -1706 1514 -1706 0 3
rlabel polysilicon 1521 -1700 1521 -1700 0 1
rlabel polysilicon 1521 -1706 1521 -1706 0 3
rlabel polysilicon 1528 -1700 1528 -1700 0 1
rlabel polysilicon 1531 -1700 1531 -1700 0 2
rlabel polysilicon 1528 -1706 1528 -1706 0 3
rlabel polysilicon 1531 -1706 1531 -1706 0 4
rlabel polysilicon 1535 -1700 1535 -1700 0 1
rlabel polysilicon 1538 -1700 1538 -1700 0 2
rlabel polysilicon 1535 -1706 1535 -1706 0 3
rlabel polysilicon 1538 -1706 1538 -1706 0 4
rlabel polysilicon 1542 -1700 1542 -1700 0 1
rlabel polysilicon 1542 -1706 1542 -1706 0 3
rlabel polysilicon 1549 -1700 1549 -1700 0 1
rlabel polysilicon 1549 -1706 1549 -1706 0 3
rlabel polysilicon 1556 -1700 1556 -1700 0 1
rlabel polysilicon 1556 -1706 1556 -1706 0 3
rlabel polysilicon 1563 -1700 1563 -1700 0 1
rlabel polysilicon 1563 -1706 1563 -1706 0 3
rlabel polysilicon 1570 -1700 1570 -1700 0 1
rlabel polysilicon 1570 -1706 1570 -1706 0 3
rlabel polysilicon 1577 -1700 1577 -1700 0 1
rlabel polysilicon 1577 -1706 1577 -1706 0 3
rlabel polysilicon 1584 -1700 1584 -1700 0 1
rlabel polysilicon 1584 -1706 1584 -1706 0 3
rlabel polysilicon 1591 -1700 1591 -1700 0 1
rlabel polysilicon 1591 -1706 1591 -1706 0 3
rlabel polysilicon 1598 -1700 1598 -1700 0 1
rlabel polysilicon 1598 -1706 1598 -1706 0 3
rlabel polysilicon 1605 -1700 1605 -1700 0 1
rlabel polysilicon 1605 -1706 1605 -1706 0 3
rlabel polysilicon 1612 -1700 1612 -1700 0 1
rlabel polysilicon 1612 -1706 1612 -1706 0 3
rlabel polysilicon 1619 -1700 1619 -1700 0 1
rlabel polysilicon 1619 -1706 1619 -1706 0 3
rlabel polysilicon 1626 -1700 1626 -1700 0 1
rlabel polysilicon 1626 -1706 1626 -1706 0 3
rlabel polysilicon 1633 -1700 1633 -1700 0 1
rlabel polysilicon 1633 -1706 1633 -1706 0 3
rlabel polysilicon 1640 -1700 1640 -1700 0 1
rlabel polysilicon 1640 -1706 1640 -1706 0 3
rlabel polysilicon 1647 -1700 1647 -1700 0 1
rlabel polysilicon 1647 -1706 1647 -1706 0 3
rlabel polysilicon 1654 -1700 1654 -1700 0 1
rlabel polysilicon 1654 -1706 1654 -1706 0 3
rlabel polysilicon 1661 -1700 1661 -1700 0 1
rlabel polysilicon 1661 -1706 1661 -1706 0 3
rlabel polysilicon 1668 -1700 1668 -1700 0 1
rlabel polysilicon 1668 -1706 1668 -1706 0 3
rlabel polysilicon 1675 -1700 1675 -1700 0 1
rlabel polysilicon 1675 -1706 1675 -1706 0 3
rlabel polysilicon 1682 -1700 1682 -1700 0 1
rlabel polysilicon 1682 -1706 1682 -1706 0 3
rlabel polysilicon 1689 -1700 1689 -1700 0 1
rlabel polysilicon 1689 -1706 1689 -1706 0 3
rlabel polysilicon 1696 -1700 1696 -1700 0 1
rlabel polysilicon 1696 -1706 1696 -1706 0 3
rlabel polysilicon 1703 -1700 1703 -1700 0 1
rlabel polysilicon 1706 -1706 1706 -1706 0 4
rlabel polysilicon 1710 -1700 1710 -1700 0 1
rlabel polysilicon 1710 -1706 1710 -1706 0 3
rlabel polysilicon 1717 -1700 1717 -1700 0 1
rlabel polysilicon 1717 -1706 1717 -1706 0 3
rlabel polysilicon 1724 -1700 1724 -1700 0 1
rlabel polysilicon 1724 -1706 1724 -1706 0 3
rlabel polysilicon 1731 -1700 1731 -1700 0 1
rlabel polysilicon 1731 -1706 1731 -1706 0 3
rlabel polysilicon 1738 -1700 1738 -1700 0 1
rlabel polysilicon 1738 -1706 1738 -1706 0 3
rlabel polysilicon 1745 -1700 1745 -1700 0 1
rlabel polysilicon 1745 -1706 1745 -1706 0 3
rlabel polysilicon 1752 -1700 1752 -1700 0 1
rlabel polysilicon 1752 -1706 1752 -1706 0 3
rlabel polysilicon 1759 -1700 1759 -1700 0 1
rlabel polysilicon 1759 -1706 1759 -1706 0 3
rlabel polysilicon 1766 -1700 1766 -1700 0 1
rlabel polysilicon 1766 -1706 1766 -1706 0 3
rlabel polysilicon 1773 -1700 1773 -1700 0 1
rlabel polysilicon 1773 -1706 1773 -1706 0 3
rlabel polysilicon 1780 -1700 1780 -1700 0 1
rlabel polysilicon 1780 -1706 1780 -1706 0 3
rlabel polysilicon 1787 -1700 1787 -1700 0 1
rlabel polysilicon 1787 -1706 1787 -1706 0 3
rlabel polysilicon 1794 -1700 1794 -1700 0 1
rlabel polysilicon 1794 -1706 1794 -1706 0 3
rlabel polysilicon 1801 -1700 1801 -1700 0 1
rlabel polysilicon 1801 -1706 1801 -1706 0 3
rlabel polysilicon 1808 -1700 1808 -1700 0 1
rlabel polysilicon 1811 -1700 1811 -1700 0 2
rlabel polysilicon 1808 -1706 1808 -1706 0 3
rlabel polysilicon 1811 -1706 1811 -1706 0 4
rlabel polysilicon 1815 -1700 1815 -1700 0 1
rlabel polysilicon 1815 -1706 1815 -1706 0 3
rlabel polysilicon 1822 -1700 1822 -1700 0 1
rlabel polysilicon 1822 -1706 1822 -1706 0 3
rlabel polysilicon 1829 -1700 1829 -1700 0 1
rlabel polysilicon 1829 -1706 1829 -1706 0 3
rlabel polysilicon 1836 -1700 1836 -1700 0 1
rlabel polysilicon 1836 -1706 1836 -1706 0 3
rlabel polysilicon 1843 -1700 1843 -1700 0 1
rlabel polysilicon 1843 -1706 1843 -1706 0 3
rlabel polysilicon 1850 -1700 1850 -1700 0 1
rlabel polysilicon 1850 -1706 1850 -1706 0 3
rlabel polysilicon 1857 -1700 1857 -1700 0 1
rlabel polysilicon 1857 -1706 1857 -1706 0 3
rlabel polysilicon 1864 -1700 1864 -1700 0 1
rlabel polysilicon 1864 -1706 1864 -1706 0 3
rlabel polysilicon 1871 -1700 1871 -1700 0 1
rlabel polysilicon 1871 -1706 1871 -1706 0 3
rlabel polysilicon 1878 -1700 1878 -1700 0 1
rlabel polysilicon 1878 -1706 1878 -1706 0 3
rlabel polysilicon 1885 -1700 1885 -1700 0 1
rlabel polysilicon 1885 -1706 1885 -1706 0 3
rlabel polysilicon 1892 -1700 1892 -1700 0 1
rlabel polysilicon 1892 -1706 1892 -1706 0 3
rlabel polysilicon 1899 -1700 1899 -1700 0 1
rlabel polysilicon 1899 -1706 1899 -1706 0 3
rlabel polysilicon 1906 -1700 1906 -1700 0 1
rlabel polysilicon 1906 -1706 1906 -1706 0 3
rlabel polysilicon 1913 -1700 1913 -1700 0 1
rlabel polysilicon 1913 -1706 1913 -1706 0 3
rlabel polysilicon 1920 -1700 1920 -1700 0 1
rlabel polysilicon 1920 -1706 1920 -1706 0 3
rlabel polysilicon 1927 -1700 1927 -1700 0 1
rlabel polysilicon 1927 -1706 1927 -1706 0 3
rlabel polysilicon 1934 -1700 1934 -1700 0 1
rlabel polysilicon 1934 -1706 1934 -1706 0 3
rlabel polysilicon 1941 -1700 1941 -1700 0 1
rlabel polysilicon 1941 -1706 1941 -1706 0 3
rlabel polysilicon 1948 -1700 1948 -1700 0 1
rlabel polysilicon 1948 -1706 1948 -1706 0 3
rlabel polysilicon 1955 -1700 1955 -1700 0 1
rlabel polysilicon 1955 -1706 1955 -1706 0 3
rlabel polysilicon 1962 -1700 1962 -1700 0 1
rlabel polysilicon 1962 -1706 1962 -1706 0 3
rlabel polysilicon 1969 -1700 1969 -1700 0 1
rlabel polysilicon 1969 -1706 1969 -1706 0 3
rlabel polysilicon 1976 -1700 1976 -1700 0 1
rlabel polysilicon 1976 -1706 1976 -1706 0 3
rlabel polysilicon 1983 -1700 1983 -1700 0 1
rlabel polysilicon 1983 -1706 1983 -1706 0 3
rlabel polysilicon 1990 -1700 1990 -1700 0 1
rlabel polysilicon 1990 -1706 1990 -1706 0 3
rlabel polysilicon 1997 -1700 1997 -1700 0 1
rlabel polysilicon 1997 -1706 1997 -1706 0 3
rlabel polysilicon 2004 -1700 2004 -1700 0 1
rlabel polysilicon 2004 -1706 2004 -1706 0 3
rlabel polysilicon 2011 -1700 2011 -1700 0 1
rlabel polysilicon 2011 -1706 2011 -1706 0 3
rlabel polysilicon 2018 -1700 2018 -1700 0 1
rlabel polysilicon 2018 -1706 2018 -1706 0 3
rlabel polysilicon 2025 -1700 2025 -1700 0 1
rlabel polysilicon 2025 -1706 2025 -1706 0 3
rlabel polysilicon 2032 -1700 2032 -1700 0 1
rlabel polysilicon 2032 -1706 2032 -1706 0 3
rlabel polysilicon 2039 -1700 2039 -1700 0 1
rlabel polysilicon 2039 -1706 2039 -1706 0 3
rlabel polysilicon 2042 -1706 2042 -1706 0 4
rlabel polysilicon 2046 -1700 2046 -1700 0 1
rlabel polysilicon 2046 -1706 2046 -1706 0 3
rlabel polysilicon 2053 -1700 2053 -1700 0 1
rlabel polysilicon 2053 -1706 2053 -1706 0 3
rlabel polysilicon 2060 -1700 2060 -1700 0 1
rlabel polysilicon 2060 -1706 2060 -1706 0 3
rlabel polysilicon 2067 -1700 2067 -1700 0 1
rlabel polysilicon 2067 -1706 2067 -1706 0 3
rlabel polysilicon 2074 -1700 2074 -1700 0 1
rlabel polysilicon 2074 -1706 2074 -1706 0 3
rlabel polysilicon 2081 -1700 2081 -1700 0 1
rlabel polysilicon 2081 -1706 2081 -1706 0 3
rlabel polysilicon 2088 -1700 2088 -1700 0 1
rlabel polysilicon 2088 -1706 2088 -1706 0 3
rlabel polysilicon 2095 -1700 2095 -1700 0 1
rlabel polysilicon 2095 -1706 2095 -1706 0 3
rlabel polysilicon 2102 -1700 2102 -1700 0 1
rlabel polysilicon 2102 -1706 2102 -1706 0 3
rlabel polysilicon 2109 -1700 2109 -1700 0 1
rlabel polysilicon 2109 -1706 2109 -1706 0 3
rlabel polysilicon 2116 -1700 2116 -1700 0 1
rlabel polysilicon 2116 -1706 2116 -1706 0 3
rlabel polysilicon 2123 -1700 2123 -1700 0 1
rlabel polysilicon 2123 -1706 2123 -1706 0 3
rlabel polysilicon 2130 -1700 2130 -1700 0 1
rlabel polysilicon 2130 -1706 2130 -1706 0 3
rlabel polysilicon 2137 -1700 2137 -1700 0 1
rlabel polysilicon 2137 -1706 2137 -1706 0 3
rlabel polysilicon 2144 -1700 2144 -1700 0 1
rlabel polysilicon 2144 -1706 2144 -1706 0 3
rlabel polysilicon 2151 -1700 2151 -1700 0 1
rlabel polysilicon 2151 -1706 2151 -1706 0 3
rlabel polysilicon 2158 -1700 2158 -1700 0 1
rlabel polysilicon 2158 -1706 2158 -1706 0 3
rlabel polysilicon 2165 -1700 2165 -1700 0 1
rlabel polysilicon 2165 -1706 2165 -1706 0 3
rlabel polysilicon 2172 -1700 2172 -1700 0 1
rlabel polysilicon 2172 -1706 2172 -1706 0 3
rlabel polysilicon 2179 -1700 2179 -1700 0 1
rlabel polysilicon 2179 -1706 2179 -1706 0 3
rlabel polysilicon 2186 -1700 2186 -1700 0 1
rlabel polysilicon 2186 -1706 2186 -1706 0 3
rlabel polysilicon 2193 -1700 2193 -1700 0 1
rlabel polysilicon 2193 -1706 2193 -1706 0 3
rlabel polysilicon 2200 -1700 2200 -1700 0 1
rlabel polysilicon 2200 -1706 2200 -1706 0 3
rlabel polysilicon 2207 -1700 2207 -1700 0 1
rlabel polysilicon 2207 -1706 2207 -1706 0 3
rlabel polysilicon 2214 -1700 2214 -1700 0 1
rlabel polysilicon 2214 -1706 2214 -1706 0 3
rlabel polysilicon 2221 -1700 2221 -1700 0 1
rlabel polysilicon 2221 -1706 2221 -1706 0 3
rlabel polysilicon 2228 -1700 2228 -1700 0 1
rlabel polysilicon 2228 -1706 2228 -1706 0 3
rlabel polysilicon 2235 -1700 2235 -1700 0 1
rlabel polysilicon 2235 -1706 2235 -1706 0 3
rlabel polysilicon 2242 -1700 2242 -1700 0 1
rlabel polysilicon 2242 -1706 2242 -1706 0 3
rlabel polysilicon 2249 -1700 2249 -1700 0 1
rlabel polysilicon 2249 -1706 2249 -1706 0 3
rlabel polysilicon 2256 -1700 2256 -1700 0 1
rlabel polysilicon 2256 -1706 2256 -1706 0 3
rlabel polysilicon 2263 -1700 2263 -1700 0 1
rlabel polysilicon 2263 -1706 2263 -1706 0 3
rlabel polysilicon 2270 -1700 2270 -1700 0 1
rlabel polysilicon 2270 -1706 2270 -1706 0 3
rlabel polysilicon 2277 -1700 2277 -1700 0 1
rlabel polysilicon 2277 -1706 2277 -1706 0 3
rlabel polysilicon 2284 -1700 2284 -1700 0 1
rlabel polysilicon 2284 -1706 2284 -1706 0 3
rlabel polysilicon 2291 -1700 2291 -1700 0 1
rlabel polysilicon 2291 -1706 2291 -1706 0 3
rlabel polysilicon 2298 -1700 2298 -1700 0 1
rlabel polysilicon 2298 -1706 2298 -1706 0 3
rlabel polysilicon 2305 -1700 2305 -1700 0 1
rlabel polysilicon 2305 -1706 2305 -1706 0 3
rlabel polysilicon 2312 -1700 2312 -1700 0 1
rlabel polysilicon 2312 -1706 2312 -1706 0 3
rlabel polysilicon 2319 -1700 2319 -1700 0 1
rlabel polysilicon 2319 -1706 2319 -1706 0 3
rlabel polysilicon 2326 -1700 2326 -1700 0 1
rlabel polysilicon 2326 -1706 2326 -1706 0 3
rlabel polysilicon 2333 -1700 2333 -1700 0 1
rlabel polysilicon 2333 -1706 2333 -1706 0 3
rlabel polysilicon 2340 -1700 2340 -1700 0 1
rlabel polysilicon 2340 -1706 2340 -1706 0 3
rlabel polysilicon 2347 -1700 2347 -1700 0 1
rlabel polysilicon 2347 -1706 2347 -1706 0 3
rlabel polysilicon 2354 -1700 2354 -1700 0 1
rlabel polysilicon 2354 -1706 2354 -1706 0 3
rlabel polysilicon 2361 -1700 2361 -1700 0 1
rlabel polysilicon 2361 -1706 2361 -1706 0 3
rlabel polysilicon 2368 -1700 2368 -1700 0 1
rlabel polysilicon 2368 -1706 2368 -1706 0 3
rlabel polysilicon 2375 -1700 2375 -1700 0 1
rlabel polysilicon 2375 -1706 2375 -1706 0 3
rlabel polysilicon 2382 -1700 2382 -1700 0 1
rlabel polysilicon 2382 -1706 2382 -1706 0 3
rlabel polysilicon 2389 -1700 2389 -1700 0 1
rlabel polysilicon 2389 -1706 2389 -1706 0 3
rlabel polysilicon 2396 -1700 2396 -1700 0 1
rlabel polysilicon 2396 -1706 2396 -1706 0 3
rlabel polysilicon 2403 -1700 2403 -1700 0 1
rlabel polysilicon 2403 -1706 2403 -1706 0 3
rlabel polysilicon 2410 -1700 2410 -1700 0 1
rlabel polysilicon 2410 -1706 2410 -1706 0 3
rlabel polysilicon 2417 -1700 2417 -1700 0 1
rlabel polysilicon 2417 -1706 2417 -1706 0 3
rlabel polysilicon 2424 -1700 2424 -1700 0 1
rlabel polysilicon 2427 -1700 2427 -1700 0 2
rlabel polysilicon 2424 -1706 2424 -1706 0 3
rlabel polysilicon 2427 -1706 2427 -1706 0 4
rlabel polysilicon 2434 -1700 2434 -1700 0 2
rlabel polysilicon 2431 -1706 2431 -1706 0 3
rlabel polysilicon 2434 -1706 2434 -1706 0 4
rlabel polysilicon 2438 -1700 2438 -1700 0 1
rlabel polysilicon 2441 -1700 2441 -1700 0 2
rlabel polysilicon 2441 -1706 2441 -1706 0 4
rlabel polysilicon 2445 -1700 2445 -1700 0 1
rlabel polysilicon 2445 -1706 2445 -1706 0 3
rlabel polysilicon 2452 -1700 2452 -1700 0 1
rlabel polysilicon 2452 -1706 2452 -1706 0 3
rlabel polysilicon 2494 -1700 2494 -1700 0 1
rlabel polysilicon 2494 -1706 2494 -1706 0 3
rlabel polysilicon 2 -1851 2 -1851 0 1
rlabel polysilicon 2 -1857 2 -1857 0 3
rlabel polysilicon 9 -1851 9 -1851 0 1
rlabel polysilicon 9 -1857 9 -1857 0 3
rlabel polysilicon 16 -1851 16 -1851 0 1
rlabel polysilicon 16 -1857 16 -1857 0 3
rlabel polysilicon 23 -1851 23 -1851 0 1
rlabel polysilicon 23 -1857 23 -1857 0 3
rlabel polysilicon 30 -1851 30 -1851 0 1
rlabel polysilicon 30 -1857 30 -1857 0 3
rlabel polysilicon 37 -1851 37 -1851 0 1
rlabel polysilicon 37 -1857 37 -1857 0 3
rlabel polysilicon 47 -1851 47 -1851 0 2
rlabel polysilicon 44 -1857 44 -1857 0 3
rlabel polysilicon 47 -1857 47 -1857 0 4
rlabel polysilicon 51 -1851 51 -1851 0 1
rlabel polysilicon 51 -1857 51 -1857 0 3
rlabel polysilicon 58 -1851 58 -1851 0 1
rlabel polysilicon 58 -1857 58 -1857 0 3
rlabel polysilicon 65 -1851 65 -1851 0 1
rlabel polysilicon 65 -1857 65 -1857 0 3
rlabel polysilicon 72 -1851 72 -1851 0 1
rlabel polysilicon 72 -1857 72 -1857 0 3
rlabel polysilicon 79 -1851 79 -1851 0 1
rlabel polysilicon 79 -1857 79 -1857 0 3
rlabel polysilicon 86 -1851 86 -1851 0 1
rlabel polysilicon 86 -1857 86 -1857 0 3
rlabel polysilicon 93 -1851 93 -1851 0 1
rlabel polysilicon 93 -1857 93 -1857 0 3
rlabel polysilicon 100 -1851 100 -1851 0 1
rlabel polysilicon 100 -1857 100 -1857 0 3
rlabel polysilicon 107 -1851 107 -1851 0 1
rlabel polysilicon 107 -1857 107 -1857 0 3
rlabel polysilicon 114 -1851 114 -1851 0 1
rlabel polysilicon 114 -1857 114 -1857 0 3
rlabel polysilicon 121 -1851 121 -1851 0 1
rlabel polysilicon 124 -1851 124 -1851 0 2
rlabel polysilicon 121 -1857 121 -1857 0 3
rlabel polysilicon 124 -1857 124 -1857 0 4
rlabel polysilicon 128 -1851 128 -1851 0 1
rlabel polysilicon 128 -1857 128 -1857 0 3
rlabel polysilicon 135 -1851 135 -1851 0 1
rlabel polysilicon 135 -1857 135 -1857 0 3
rlabel polysilicon 142 -1851 142 -1851 0 1
rlabel polysilicon 142 -1857 142 -1857 0 3
rlabel polysilicon 149 -1851 149 -1851 0 1
rlabel polysilicon 149 -1857 149 -1857 0 3
rlabel polysilicon 159 -1851 159 -1851 0 2
rlabel polysilicon 159 -1857 159 -1857 0 4
rlabel polysilicon 163 -1851 163 -1851 0 1
rlabel polysilicon 163 -1857 163 -1857 0 3
rlabel polysilicon 170 -1851 170 -1851 0 1
rlabel polysilicon 170 -1857 170 -1857 0 3
rlabel polysilicon 177 -1851 177 -1851 0 1
rlabel polysilicon 177 -1857 177 -1857 0 3
rlabel polysilicon 184 -1851 184 -1851 0 1
rlabel polysilicon 187 -1851 187 -1851 0 2
rlabel polysilicon 184 -1857 184 -1857 0 3
rlabel polysilicon 187 -1857 187 -1857 0 4
rlabel polysilicon 191 -1851 191 -1851 0 1
rlabel polysilicon 191 -1857 191 -1857 0 3
rlabel polysilicon 198 -1851 198 -1851 0 1
rlabel polysilicon 201 -1851 201 -1851 0 2
rlabel polysilicon 198 -1857 198 -1857 0 3
rlabel polysilicon 205 -1851 205 -1851 0 1
rlabel polysilicon 205 -1857 205 -1857 0 3
rlabel polysilicon 212 -1851 212 -1851 0 1
rlabel polysilicon 212 -1857 212 -1857 0 3
rlabel polysilicon 219 -1851 219 -1851 0 1
rlabel polysilicon 219 -1857 219 -1857 0 3
rlabel polysilicon 226 -1851 226 -1851 0 1
rlabel polysilicon 226 -1857 226 -1857 0 3
rlabel polysilicon 229 -1857 229 -1857 0 4
rlabel polysilicon 233 -1851 233 -1851 0 1
rlabel polysilicon 236 -1851 236 -1851 0 2
rlabel polysilicon 233 -1857 233 -1857 0 3
rlabel polysilicon 240 -1851 240 -1851 0 1
rlabel polysilicon 240 -1857 240 -1857 0 3
rlabel polysilicon 250 -1851 250 -1851 0 2
rlabel polysilicon 247 -1857 247 -1857 0 3
rlabel polysilicon 250 -1857 250 -1857 0 4
rlabel polysilicon 254 -1851 254 -1851 0 1
rlabel polysilicon 254 -1857 254 -1857 0 3
rlabel polysilicon 261 -1851 261 -1851 0 1
rlabel polysilicon 261 -1857 261 -1857 0 3
rlabel polysilicon 268 -1851 268 -1851 0 1
rlabel polysilicon 268 -1857 268 -1857 0 3
rlabel polysilicon 275 -1851 275 -1851 0 1
rlabel polysilicon 275 -1857 275 -1857 0 3
rlabel polysilicon 282 -1851 282 -1851 0 1
rlabel polysilicon 282 -1857 282 -1857 0 3
rlabel polysilicon 289 -1851 289 -1851 0 1
rlabel polysilicon 289 -1857 289 -1857 0 3
rlabel polysilicon 296 -1851 296 -1851 0 1
rlabel polysilicon 296 -1857 296 -1857 0 3
rlabel polysilicon 303 -1851 303 -1851 0 1
rlabel polysilicon 303 -1857 303 -1857 0 3
rlabel polysilicon 310 -1851 310 -1851 0 1
rlabel polysilicon 310 -1857 310 -1857 0 3
rlabel polysilicon 317 -1851 317 -1851 0 1
rlabel polysilicon 317 -1857 317 -1857 0 3
rlabel polysilicon 324 -1851 324 -1851 0 1
rlabel polysilicon 324 -1857 324 -1857 0 3
rlabel polysilicon 331 -1851 331 -1851 0 1
rlabel polysilicon 331 -1857 331 -1857 0 3
rlabel polysilicon 338 -1851 338 -1851 0 1
rlabel polysilicon 338 -1857 338 -1857 0 3
rlabel polysilicon 345 -1851 345 -1851 0 1
rlabel polysilicon 345 -1857 345 -1857 0 3
rlabel polysilicon 352 -1851 352 -1851 0 1
rlabel polysilicon 352 -1857 352 -1857 0 3
rlabel polysilicon 359 -1851 359 -1851 0 1
rlabel polysilicon 359 -1857 359 -1857 0 3
rlabel polysilicon 366 -1851 366 -1851 0 1
rlabel polysilicon 366 -1857 366 -1857 0 3
rlabel polysilicon 373 -1851 373 -1851 0 1
rlabel polysilicon 373 -1857 373 -1857 0 3
rlabel polysilicon 380 -1851 380 -1851 0 1
rlabel polysilicon 380 -1857 380 -1857 0 3
rlabel polysilicon 387 -1851 387 -1851 0 1
rlabel polysilicon 387 -1857 387 -1857 0 3
rlabel polysilicon 394 -1851 394 -1851 0 1
rlabel polysilicon 394 -1857 394 -1857 0 3
rlabel polysilicon 401 -1851 401 -1851 0 1
rlabel polysilicon 401 -1857 401 -1857 0 3
rlabel polysilicon 408 -1851 408 -1851 0 1
rlabel polysilicon 408 -1857 408 -1857 0 3
rlabel polysilicon 415 -1851 415 -1851 0 1
rlabel polysilicon 415 -1857 415 -1857 0 3
rlabel polysilicon 422 -1851 422 -1851 0 1
rlabel polysilicon 422 -1857 422 -1857 0 3
rlabel polysilicon 429 -1851 429 -1851 0 1
rlabel polysilicon 429 -1857 429 -1857 0 3
rlabel polysilicon 432 -1857 432 -1857 0 4
rlabel polysilicon 436 -1851 436 -1851 0 1
rlabel polysilicon 436 -1857 436 -1857 0 3
rlabel polysilicon 443 -1851 443 -1851 0 1
rlabel polysilicon 446 -1851 446 -1851 0 2
rlabel polysilicon 443 -1857 443 -1857 0 3
rlabel polysilicon 446 -1857 446 -1857 0 4
rlabel polysilicon 450 -1857 450 -1857 0 3
rlabel polysilicon 457 -1851 457 -1851 0 1
rlabel polysilicon 457 -1857 457 -1857 0 3
rlabel polysilicon 464 -1851 464 -1851 0 1
rlabel polysilicon 464 -1857 464 -1857 0 3
rlabel polysilicon 471 -1851 471 -1851 0 1
rlabel polysilicon 471 -1857 471 -1857 0 3
rlabel polysilicon 478 -1851 478 -1851 0 1
rlabel polysilicon 478 -1857 478 -1857 0 3
rlabel polysilicon 485 -1851 485 -1851 0 1
rlabel polysilicon 485 -1857 485 -1857 0 3
rlabel polysilicon 492 -1851 492 -1851 0 1
rlabel polysilicon 492 -1857 492 -1857 0 3
rlabel polysilicon 499 -1851 499 -1851 0 1
rlabel polysilicon 499 -1857 499 -1857 0 3
rlabel polysilicon 506 -1851 506 -1851 0 1
rlabel polysilicon 506 -1857 506 -1857 0 3
rlabel polysilicon 513 -1851 513 -1851 0 1
rlabel polysilicon 516 -1851 516 -1851 0 2
rlabel polysilicon 513 -1857 513 -1857 0 3
rlabel polysilicon 516 -1857 516 -1857 0 4
rlabel polysilicon 520 -1851 520 -1851 0 1
rlabel polysilicon 520 -1857 520 -1857 0 3
rlabel polysilicon 527 -1851 527 -1851 0 1
rlabel polysilicon 527 -1857 527 -1857 0 3
rlabel polysilicon 534 -1851 534 -1851 0 1
rlabel polysilicon 534 -1857 534 -1857 0 3
rlabel polysilicon 541 -1851 541 -1851 0 1
rlabel polysilicon 541 -1857 541 -1857 0 3
rlabel polysilicon 548 -1851 548 -1851 0 1
rlabel polysilicon 548 -1857 548 -1857 0 3
rlabel polysilicon 555 -1851 555 -1851 0 1
rlabel polysilicon 555 -1857 555 -1857 0 3
rlabel polysilicon 562 -1851 562 -1851 0 1
rlabel polysilicon 565 -1851 565 -1851 0 2
rlabel polysilicon 562 -1857 562 -1857 0 3
rlabel polysilicon 565 -1857 565 -1857 0 4
rlabel polysilicon 569 -1851 569 -1851 0 1
rlabel polysilicon 569 -1857 569 -1857 0 3
rlabel polysilicon 576 -1851 576 -1851 0 1
rlabel polysilicon 576 -1857 576 -1857 0 3
rlabel polysilicon 583 -1851 583 -1851 0 1
rlabel polysilicon 583 -1857 583 -1857 0 3
rlabel polysilicon 590 -1851 590 -1851 0 1
rlabel polysilicon 590 -1857 590 -1857 0 3
rlabel polysilicon 597 -1851 597 -1851 0 1
rlabel polysilicon 597 -1857 597 -1857 0 3
rlabel polysilicon 604 -1851 604 -1851 0 1
rlabel polysilicon 604 -1857 604 -1857 0 3
rlabel polysilicon 611 -1851 611 -1851 0 1
rlabel polysilicon 614 -1851 614 -1851 0 2
rlabel polysilicon 611 -1857 611 -1857 0 3
rlabel polysilicon 614 -1857 614 -1857 0 4
rlabel polysilicon 618 -1851 618 -1851 0 1
rlabel polysilicon 618 -1857 618 -1857 0 3
rlabel polysilicon 625 -1851 625 -1851 0 1
rlabel polysilicon 625 -1857 625 -1857 0 3
rlabel polysilicon 632 -1857 632 -1857 0 3
rlabel polysilicon 635 -1857 635 -1857 0 4
rlabel polysilicon 639 -1851 639 -1851 0 1
rlabel polysilicon 639 -1857 639 -1857 0 3
rlabel polysilicon 646 -1851 646 -1851 0 1
rlabel polysilicon 649 -1851 649 -1851 0 2
rlabel polysilicon 646 -1857 646 -1857 0 3
rlabel polysilicon 649 -1857 649 -1857 0 4
rlabel polysilicon 653 -1851 653 -1851 0 1
rlabel polysilicon 653 -1857 653 -1857 0 3
rlabel polysilicon 660 -1851 660 -1851 0 1
rlabel polysilicon 660 -1857 660 -1857 0 3
rlabel polysilicon 667 -1851 667 -1851 0 1
rlabel polysilicon 667 -1857 667 -1857 0 3
rlabel polysilicon 674 -1851 674 -1851 0 1
rlabel polysilicon 674 -1857 674 -1857 0 3
rlabel polysilicon 681 -1851 681 -1851 0 1
rlabel polysilicon 681 -1857 681 -1857 0 3
rlabel polysilicon 688 -1851 688 -1851 0 1
rlabel polysilicon 688 -1857 688 -1857 0 3
rlabel polysilicon 695 -1851 695 -1851 0 1
rlabel polysilicon 695 -1857 695 -1857 0 3
rlabel polysilicon 702 -1851 702 -1851 0 1
rlabel polysilicon 702 -1857 702 -1857 0 3
rlabel polysilicon 709 -1851 709 -1851 0 1
rlabel polysilicon 709 -1857 709 -1857 0 3
rlabel polysilicon 716 -1851 716 -1851 0 1
rlabel polysilicon 716 -1857 716 -1857 0 3
rlabel polysilicon 723 -1851 723 -1851 0 1
rlabel polysilicon 723 -1857 723 -1857 0 3
rlabel polysilicon 726 -1857 726 -1857 0 4
rlabel polysilicon 730 -1851 730 -1851 0 1
rlabel polysilicon 733 -1851 733 -1851 0 2
rlabel polysilicon 730 -1857 730 -1857 0 3
rlabel polysilicon 737 -1851 737 -1851 0 1
rlabel polysilicon 740 -1851 740 -1851 0 2
rlabel polysilicon 737 -1857 737 -1857 0 3
rlabel polysilicon 740 -1857 740 -1857 0 4
rlabel polysilicon 744 -1851 744 -1851 0 1
rlabel polysilicon 744 -1857 744 -1857 0 3
rlabel polysilicon 751 -1851 751 -1851 0 1
rlabel polysilicon 751 -1857 751 -1857 0 3
rlabel polysilicon 758 -1851 758 -1851 0 1
rlabel polysilicon 758 -1857 758 -1857 0 3
rlabel polysilicon 765 -1851 765 -1851 0 1
rlabel polysilicon 765 -1857 765 -1857 0 3
rlabel polysilicon 772 -1851 772 -1851 0 1
rlabel polysilicon 772 -1857 772 -1857 0 3
rlabel polysilicon 779 -1851 779 -1851 0 1
rlabel polysilicon 779 -1857 779 -1857 0 3
rlabel polysilicon 786 -1851 786 -1851 0 1
rlabel polysilicon 786 -1857 786 -1857 0 3
rlabel polysilicon 793 -1851 793 -1851 0 1
rlabel polysilicon 793 -1857 793 -1857 0 3
rlabel polysilicon 800 -1851 800 -1851 0 1
rlabel polysilicon 803 -1851 803 -1851 0 2
rlabel polysilicon 800 -1857 800 -1857 0 3
rlabel polysilicon 803 -1857 803 -1857 0 4
rlabel polysilicon 807 -1851 807 -1851 0 1
rlabel polysilicon 807 -1857 807 -1857 0 3
rlabel polysilicon 814 -1851 814 -1851 0 1
rlabel polysilicon 814 -1857 814 -1857 0 3
rlabel polysilicon 821 -1851 821 -1851 0 1
rlabel polysilicon 821 -1857 821 -1857 0 3
rlabel polysilicon 828 -1851 828 -1851 0 1
rlabel polysilicon 828 -1857 828 -1857 0 3
rlabel polysilicon 835 -1851 835 -1851 0 1
rlabel polysilicon 835 -1857 835 -1857 0 3
rlabel polysilicon 842 -1851 842 -1851 0 1
rlabel polysilicon 842 -1857 842 -1857 0 3
rlabel polysilicon 849 -1857 849 -1857 0 3
rlabel polysilicon 852 -1857 852 -1857 0 4
rlabel polysilicon 856 -1851 856 -1851 0 1
rlabel polysilicon 856 -1857 856 -1857 0 3
rlabel polysilicon 863 -1851 863 -1851 0 1
rlabel polysilicon 863 -1857 863 -1857 0 3
rlabel polysilicon 870 -1851 870 -1851 0 1
rlabel polysilicon 870 -1857 870 -1857 0 3
rlabel polysilicon 877 -1851 877 -1851 0 1
rlabel polysilicon 877 -1857 877 -1857 0 3
rlabel polysilicon 884 -1851 884 -1851 0 1
rlabel polysilicon 884 -1857 884 -1857 0 3
rlabel polysilicon 891 -1851 891 -1851 0 1
rlabel polysilicon 894 -1851 894 -1851 0 2
rlabel polysilicon 891 -1857 891 -1857 0 3
rlabel polysilicon 894 -1857 894 -1857 0 4
rlabel polysilicon 898 -1851 898 -1851 0 1
rlabel polysilicon 898 -1857 898 -1857 0 3
rlabel polysilicon 905 -1851 905 -1851 0 1
rlabel polysilicon 908 -1851 908 -1851 0 2
rlabel polysilicon 908 -1857 908 -1857 0 4
rlabel polysilicon 912 -1851 912 -1851 0 1
rlabel polysilicon 912 -1857 912 -1857 0 3
rlabel polysilicon 919 -1851 919 -1851 0 1
rlabel polysilicon 919 -1857 919 -1857 0 3
rlabel polysilicon 926 -1851 926 -1851 0 1
rlabel polysilicon 926 -1857 926 -1857 0 3
rlabel polysilicon 933 -1851 933 -1851 0 1
rlabel polysilicon 933 -1857 933 -1857 0 3
rlabel polysilicon 940 -1851 940 -1851 0 1
rlabel polysilicon 943 -1851 943 -1851 0 2
rlabel polysilicon 940 -1857 940 -1857 0 3
rlabel polysilicon 943 -1857 943 -1857 0 4
rlabel polysilicon 947 -1851 947 -1851 0 1
rlabel polysilicon 947 -1857 947 -1857 0 3
rlabel polysilicon 954 -1851 954 -1851 0 1
rlabel polysilicon 957 -1851 957 -1851 0 2
rlabel polysilicon 954 -1857 954 -1857 0 3
rlabel polysilicon 957 -1857 957 -1857 0 4
rlabel polysilicon 961 -1851 961 -1851 0 1
rlabel polysilicon 961 -1857 961 -1857 0 3
rlabel polysilicon 968 -1851 968 -1851 0 1
rlabel polysilicon 968 -1857 968 -1857 0 3
rlabel polysilicon 975 -1851 975 -1851 0 1
rlabel polysilicon 975 -1857 975 -1857 0 3
rlabel polysilicon 982 -1851 982 -1851 0 1
rlabel polysilicon 982 -1857 982 -1857 0 3
rlabel polysilicon 989 -1851 989 -1851 0 1
rlabel polysilicon 989 -1857 989 -1857 0 3
rlabel polysilicon 996 -1851 996 -1851 0 1
rlabel polysilicon 996 -1857 996 -1857 0 3
rlabel polysilicon 1003 -1851 1003 -1851 0 1
rlabel polysilicon 1003 -1857 1003 -1857 0 3
rlabel polysilicon 1010 -1851 1010 -1851 0 1
rlabel polysilicon 1010 -1857 1010 -1857 0 3
rlabel polysilicon 1017 -1851 1017 -1851 0 1
rlabel polysilicon 1017 -1857 1017 -1857 0 3
rlabel polysilicon 1024 -1851 1024 -1851 0 1
rlabel polysilicon 1024 -1857 1024 -1857 0 3
rlabel polysilicon 1031 -1851 1031 -1851 0 1
rlabel polysilicon 1031 -1857 1031 -1857 0 3
rlabel polysilicon 1038 -1851 1038 -1851 0 1
rlabel polysilicon 1038 -1857 1038 -1857 0 3
rlabel polysilicon 1045 -1851 1045 -1851 0 1
rlabel polysilicon 1045 -1857 1045 -1857 0 3
rlabel polysilicon 1052 -1851 1052 -1851 0 1
rlabel polysilicon 1052 -1857 1052 -1857 0 3
rlabel polysilicon 1059 -1851 1059 -1851 0 1
rlabel polysilicon 1059 -1857 1059 -1857 0 3
rlabel polysilicon 1066 -1851 1066 -1851 0 1
rlabel polysilicon 1066 -1857 1066 -1857 0 3
rlabel polysilicon 1073 -1851 1073 -1851 0 1
rlabel polysilicon 1073 -1857 1073 -1857 0 3
rlabel polysilicon 1080 -1851 1080 -1851 0 1
rlabel polysilicon 1080 -1857 1080 -1857 0 3
rlabel polysilicon 1087 -1851 1087 -1851 0 1
rlabel polysilicon 1087 -1857 1087 -1857 0 3
rlabel polysilicon 1094 -1851 1094 -1851 0 1
rlabel polysilicon 1094 -1857 1094 -1857 0 3
rlabel polysilicon 1101 -1851 1101 -1851 0 1
rlabel polysilicon 1101 -1857 1101 -1857 0 3
rlabel polysilicon 1108 -1851 1108 -1851 0 1
rlabel polysilicon 1108 -1857 1108 -1857 0 3
rlabel polysilicon 1115 -1851 1115 -1851 0 1
rlabel polysilicon 1115 -1857 1115 -1857 0 3
rlabel polysilicon 1122 -1851 1122 -1851 0 1
rlabel polysilicon 1122 -1857 1122 -1857 0 3
rlabel polysilicon 1129 -1851 1129 -1851 0 1
rlabel polysilicon 1129 -1857 1129 -1857 0 3
rlabel polysilicon 1136 -1851 1136 -1851 0 1
rlabel polysilicon 1136 -1857 1136 -1857 0 3
rlabel polysilicon 1139 -1857 1139 -1857 0 4
rlabel polysilicon 1143 -1851 1143 -1851 0 1
rlabel polysilicon 1143 -1857 1143 -1857 0 3
rlabel polysilicon 1150 -1851 1150 -1851 0 1
rlabel polysilicon 1150 -1857 1150 -1857 0 3
rlabel polysilicon 1157 -1851 1157 -1851 0 1
rlabel polysilicon 1157 -1857 1157 -1857 0 3
rlabel polysilicon 1164 -1851 1164 -1851 0 1
rlabel polysilicon 1164 -1857 1164 -1857 0 3
rlabel polysilicon 1171 -1851 1171 -1851 0 1
rlabel polysilicon 1171 -1857 1171 -1857 0 3
rlabel polysilicon 1178 -1851 1178 -1851 0 1
rlabel polysilicon 1181 -1851 1181 -1851 0 2
rlabel polysilicon 1178 -1857 1178 -1857 0 3
rlabel polysilicon 1181 -1857 1181 -1857 0 4
rlabel polysilicon 1185 -1851 1185 -1851 0 1
rlabel polysilicon 1185 -1857 1185 -1857 0 3
rlabel polysilicon 1192 -1851 1192 -1851 0 1
rlabel polysilicon 1192 -1857 1192 -1857 0 3
rlabel polysilicon 1199 -1851 1199 -1851 0 1
rlabel polysilicon 1199 -1857 1199 -1857 0 3
rlabel polysilicon 1209 -1851 1209 -1851 0 2
rlabel polysilicon 1206 -1857 1206 -1857 0 3
rlabel polysilicon 1209 -1857 1209 -1857 0 4
rlabel polysilicon 1213 -1851 1213 -1851 0 1
rlabel polysilicon 1213 -1857 1213 -1857 0 3
rlabel polysilicon 1220 -1851 1220 -1851 0 1
rlabel polysilicon 1220 -1857 1220 -1857 0 3
rlabel polysilicon 1227 -1851 1227 -1851 0 1
rlabel polysilicon 1227 -1857 1227 -1857 0 3
rlabel polysilicon 1234 -1851 1234 -1851 0 1
rlabel polysilicon 1234 -1857 1234 -1857 0 3
rlabel polysilicon 1241 -1851 1241 -1851 0 1
rlabel polysilicon 1241 -1857 1241 -1857 0 3
rlabel polysilicon 1248 -1851 1248 -1851 0 1
rlabel polysilicon 1248 -1857 1248 -1857 0 3
rlabel polysilicon 1255 -1851 1255 -1851 0 1
rlabel polysilicon 1255 -1857 1255 -1857 0 3
rlabel polysilicon 1262 -1851 1262 -1851 0 1
rlabel polysilicon 1262 -1857 1262 -1857 0 3
rlabel polysilicon 1269 -1851 1269 -1851 0 1
rlabel polysilicon 1269 -1857 1269 -1857 0 3
rlabel polysilicon 1276 -1851 1276 -1851 0 1
rlabel polysilicon 1279 -1851 1279 -1851 0 2
rlabel polysilicon 1276 -1857 1276 -1857 0 3
rlabel polysilicon 1279 -1857 1279 -1857 0 4
rlabel polysilicon 1283 -1851 1283 -1851 0 1
rlabel polysilicon 1283 -1857 1283 -1857 0 3
rlabel polysilicon 1290 -1851 1290 -1851 0 1
rlabel polysilicon 1293 -1851 1293 -1851 0 2
rlabel polysilicon 1290 -1857 1290 -1857 0 3
rlabel polysilicon 1297 -1851 1297 -1851 0 1
rlabel polysilicon 1297 -1857 1297 -1857 0 3
rlabel polysilicon 1304 -1851 1304 -1851 0 1
rlabel polysilicon 1307 -1851 1307 -1851 0 2
rlabel polysilicon 1304 -1857 1304 -1857 0 3
rlabel polysilicon 1307 -1857 1307 -1857 0 4
rlabel polysilicon 1311 -1851 1311 -1851 0 1
rlabel polysilicon 1311 -1857 1311 -1857 0 3
rlabel polysilicon 1318 -1851 1318 -1851 0 1
rlabel polysilicon 1318 -1857 1318 -1857 0 3
rlabel polysilicon 1325 -1851 1325 -1851 0 1
rlabel polysilicon 1332 -1851 1332 -1851 0 1
rlabel polysilicon 1332 -1857 1332 -1857 0 3
rlabel polysilicon 1335 -1857 1335 -1857 0 4
rlabel polysilicon 1339 -1851 1339 -1851 0 1
rlabel polysilicon 1339 -1857 1339 -1857 0 3
rlabel polysilicon 1346 -1851 1346 -1851 0 1
rlabel polysilicon 1346 -1857 1346 -1857 0 3
rlabel polysilicon 1353 -1851 1353 -1851 0 1
rlabel polysilicon 1353 -1857 1353 -1857 0 3
rlabel polysilicon 1360 -1851 1360 -1851 0 1
rlabel polysilicon 1360 -1857 1360 -1857 0 3
rlabel polysilicon 1367 -1851 1367 -1851 0 1
rlabel polysilicon 1367 -1857 1367 -1857 0 3
rlabel polysilicon 1374 -1851 1374 -1851 0 1
rlabel polysilicon 1374 -1857 1374 -1857 0 3
rlabel polysilicon 1381 -1851 1381 -1851 0 1
rlabel polysilicon 1381 -1857 1381 -1857 0 3
rlabel polysilicon 1388 -1851 1388 -1851 0 1
rlabel polysilicon 1388 -1857 1388 -1857 0 3
rlabel polysilicon 1395 -1851 1395 -1851 0 1
rlabel polysilicon 1395 -1857 1395 -1857 0 3
rlabel polysilicon 1402 -1851 1402 -1851 0 1
rlabel polysilicon 1402 -1857 1402 -1857 0 3
rlabel polysilicon 1409 -1851 1409 -1851 0 1
rlabel polysilicon 1409 -1857 1409 -1857 0 3
rlabel polysilicon 1416 -1851 1416 -1851 0 1
rlabel polysilicon 1416 -1857 1416 -1857 0 3
rlabel polysilicon 1423 -1851 1423 -1851 0 1
rlabel polysilicon 1423 -1857 1423 -1857 0 3
rlabel polysilicon 1430 -1851 1430 -1851 0 1
rlabel polysilicon 1430 -1857 1430 -1857 0 3
rlabel polysilicon 1437 -1851 1437 -1851 0 1
rlabel polysilicon 1440 -1851 1440 -1851 0 2
rlabel polysilicon 1437 -1857 1437 -1857 0 3
rlabel polysilicon 1440 -1857 1440 -1857 0 4
rlabel polysilicon 1444 -1851 1444 -1851 0 1
rlabel polysilicon 1444 -1857 1444 -1857 0 3
rlabel polysilicon 1451 -1851 1451 -1851 0 1
rlabel polysilicon 1451 -1857 1451 -1857 0 3
rlabel polysilicon 1458 -1851 1458 -1851 0 1
rlabel polysilicon 1458 -1857 1458 -1857 0 3
rlabel polysilicon 1465 -1851 1465 -1851 0 1
rlabel polysilicon 1468 -1851 1468 -1851 0 2
rlabel polysilicon 1465 -1857 1465 -1857 0 3
rlabel polysilicon 1468 -1857 1468 -1857 0 4
rlabel polysilicon 1472 -1851 1472 -1851 0 1
rlabel polysilicon 1472 -1857 1472 -1857 0 3
rlabel polysilicon 1479 -1851 1479 -1851 0 1
rlabel polysilicon 1479 -1857 1479 -1857 0 3
rlabel polysilicon 1486 -1851 1486 -1851 0 1
rlabel polysilicon 1486 -1857 1486 -1857 0 3
rlabel polysilicon 1493 -1851 1493 -1851 0 1
rlabel polysilicon 1493 -1857 1493 -1857 0 3
rlabel polysilicon 1500 -1851 1500 -1851 0 1
rlabel polysilicon 1500 -1857 1500 -1857 0 3
rlabel polysilicon 1507 -1851 1507 -1851 0 1
rlabel polysilicon 1507 -1857 1507 -1857 0 3
rlabel polysilicon 1510 -1857 1510 -1857 0 4
rlabel polysilicon 1514 -1851 1514 -1851 0 1
rlabel polysilicon 1514 -1857 1514 -1857 0 3
rlabel polysilicon 1521 -1851 1521 -1851 0 1
rlabel polysilicon 1521 -1857 1521 -1857 0 3
rlabel polysilicon 1528 -1851 1528 -1851 0 1
rlabel polysilicon 1528 -1857 1528 -1857 0 3
rlabel polysilicon 1535 -1851 1535 -1851 0 1
rlabel polysilicon 1535 -1857 1535 -1857 0 3
rlabel polysilicon 1542 -1851 1542 -1851 0 1
rlabel polysilicon 1542 -1857 1542 -1857 0 3
rlabel polysilicon 1549 -1851 1549 -1851 0 1
rlabel polysilicon 1549 -1857 1549 -1857 0 3
rlabel polysilicon 1556 -1851 1556 -1851 0 1
rlabel polysilicon 1556 -1857 1556 -1857 0 3
rlabel polysilicon 1563 -1851 1563 -1851 0 1
rlabel polysilicon 1563 -1857 1563 -1857 0 3
rlabel polysilicon 1570 -1851 1570 -1851 0 1
rlabel polysilicon 1570 -1857 1570 -1857 0 3
rlabel polysilicon 1577 -1851 1577 -1851 0 1
rlabel polysilicon 1577 -1857 1577 -1857 0 3
rlabel polysilicon 1584 -1851 1584 -1851 0 1
rlabel polysilicon 1584 -1857 1584 -1857 0 3
rlabel polysilicon 1591 -1851 1591 -1851 0 1
rlabel polysilicon 1591 -1857 1591 -1857 0 3
rlabel polysilicon 1598 -1851 1598 -1851 0 1
rlabel polysilicon 1598 -1857 1598 -1857 0 3
rlabel polysilicon 1605 -1851 1605 -1851 0 1
rlabel polysilicon 1605 -1857 1605 -1857 0 3
rlabel polysilicon 1612 -1851 1612 -1851 0 1
rlabel polysilicon 1612 -1857 1612 -1857 0 3
rlabel polysilicon 1619 -1851 1619 -1851 0 1
rlabel polysilicon 1619 -1857 1619 -1857 0 3
rlabel polysilicon 1626 -1851 1626 -1851 0 1
rlabel polysilicon 1629 -1851 1629 -1851 0 2
rlabel polysilicon 1629 -1857 1629 -1857 0 4
rlabel polysilicon 1633 -1851 1633 -1851 0 1
rlabel polysilicon 1633 -1857 1633 -1857 0 3
rlabel polysilicon 1640 -1851 1640 -1851 0 1
rlabel polysilicon 1640 -1857 1640 -1857 0 3
rlabel polysilicon 1647 -1851 1647 -1851 0 1
rlabel polysilicon 1647 -1857 1647 -1857 0 3
rlabel polysilicon 1654 -1851 1654 -1851 0 1
rlabel polysilicon 1654 -1857 1654 -1857 0 3
rlabel polysilicon 1664 -1851 1664 -1851 0 2
rlabel polysilicon 1661 -1857 1661 -1857 0 3
rlabel polysilicon 1664 -1857 1664 -1857 0 4
rlabel polysilicon 1668 -1851 1668 -1851 0 1
rlabel polysilicon 1668 -1857 1668 -1857 0 3
rlabel polysilicon 1675 -1851 1675 -1851 0 1
rlabel polysilicon 1675 -1857 1675 -1857 0 3
rlabel polysilicon 1682 -1851 1682 -1851 0 1
rlabel polysilicon 1682 -1857 1682 -1857 0 3
rlabel polysilicon 1689 -1851 1689 -1851 0 1
rlabel polysilicon 1689 -1857 1689 -1857 0 3
rlabel polysilicon 1696 -1851 1696 -1851 0 1
rlabel polysilicon 1696 -1857 1696 -1857 0 3
rlabel polysilicon 1703 -1851 1703 -1851 0 1
rlabel polysilicon 1703 -1857 1703 -1857 0 3
rlabel polysilicon 1710 -1851 1710 -1851 0 1
rlabel polysilicon 1710 -1857 1710 -1857 0 3
rlabel polysilicon 1717 -1851 1717 -1851 0 1
rlabel polysilicon 1717 -1857 1717 -1857 0 3
rlabel polysilicon 1724 -1851 1724 -1851 0 1
rlabel polysilicon 1724 -1857 1724 -1857 0 3
rlabel polysilicon 1731 -1851 1731 -1851 0 1
rlabel polysilicon 1731 -1857 1731 -1857 0 3
rlabel polysilicon 1738 -1851 1738 -1851 0 1
rlabel polysilicon 1738 -1857 1738 -1857 0 3
rlabel polysilicon 1745 -1851 1745 -1851 0 1
rlabel polysilicon 1745 -1857 1745 -1857 0 3
rlabel polysilicon 1752 -1851 1752 -1851 0 1
rlabel polysilicon 1752 -1857 1752 -1857 0 3
rlabel polysilicon 1759 -1851 1759 -1851 0 1
rlabel polysilicon 1759 -1857 1759 -1857 0 3
rlabel polysilicon 1766 -1851 1766 -1851 0 1
rlabel polysilicon 1766 -1857 1766 -1857 0 3
rlabel polysilicon 1773 -1851 1773 -1851 0 1
rlabel polysilicon 1773 -1857 1773 -1857 0 3
rlabel polysilicon 1780 -1851 1780 -1851 0 1
rlabel polysilicon 1780 -1857 1780 -1857 0 3
rlabel polysilicon 1787 -1851 1787 -1851 0 1
rlabel polysilicon 1787 -1857 1787 -1857 0 3
rlabel polysilicon 1794 -1851 1794 -1851 0 1
rlabel polysilicon 1794 -1857 1794 -1857 0 3
rlabel polysilicon 1801 -1851 1801 -1851 0 1
rlabel polysilicon 1801 -1857 1801 -1857 0 3
rlabel polysilicon 1808 -1851 1808 -1851 0 1
rlabel polysilicon 1808 -1857 1808 -1857 0 3
rlabel polysilicon 1815 -1851 1815 -1851 0 1
rlabel polysilicon 1815 -1857 1815 -1857 0 3
rlabel polysilicon 1822 -1851 1822 -1851 0 1
rlabel polysilicon 1822 -1857 1822 -1857 0 3
rlabel polysilicon 1829 -1851 1829 -1851 0 1
rlabel polysilicon 1829 -1857 1829 -1857 0 3
rlabel polysilicon 1836 -1851 1836 -1851 0 1
rlabel polysilicon 1836 -1857 1836 -1857 0 3
rlabel polysilicon 1843 -1851 1843 -1851 0 1
rlabel polysilicon 1843 -1857 1843 -1857 0 3
rlabel polysilicon 1850 -1851 1850 -1851 0 1
rlabel polysilicon 1853 -1851 1853 -1851 0 2
rlabel polysilicon 1850 -1857 1850 -1857 0 3
rlabel polysilicon 1853 -1857 1853 -1857 0 4
rlabel polysilicon 1857 -1851 1857 -1851 0 1
rlabel polysilicon 1857 -1857 1857 -1857 0 3
rlabel polysilicon 1864 -1857 1864 -1857 0 3
rlabel polysilicon 1867 -1857 1867 -1857 0 4
rlabel polysilicon 1871 -1851 1871 -1851 0 1
rlabel polysilicon 1871 -1857 1871 -1857 0 3
rlabel polysilicon 1878 -1851 1878 -1851 0 1
rlabel polysilicon 1878 -1857 1878 -1857 0 3
rlabel polysilicon 1885 -1851 1885 -1851 0 1
rlabel polysilicon 1885 -1857 1885 -1857 0 3
rlabel polysilicon 1892 -1851 1892 -1851 0 1
rlabel polysilicon 1892 -1857 1892 -1857 0 3
rlabel polysilicon 1899 -1851 1899 -1851 0 1
rlabel polysilicon 1899 -1857 1899 -1857 0 3
rlabel polysilicon 1906 -1851 1906 -1851 0 1
rlabel polysilicon 1906 -1857 1906 -1857 0 3
rlabel polysilicon 1913 -1851 1913 -1851 0 1
rlabel polysilicon 1913 -1857 1913 -1857 0 3
rlabel polysilicon 1920 -1851 1920 -1851 0 1
rlabel polysilicon 1920 -1857 1920 -1857 0 3
rlabel polysilicon 1927 -1851 1927 -1851 0 1
rlabel polysilicon 1927 -1857 1927 -1857 0 3
rlabel polysilicon 1934 -1851 1934 -1851 0 1
rlabel polysilicon 1934 -1857 1934 -1857 0 3
rlabel polysilicon 1941 -1851 1941 -1851 0 1
rlabel polysilicon 1941 -1857 1941 -1857 0 3
rlabel polysilicon 1948 -1851 1948 -1851 0 1
rlabel polysilicon 1948 -1857 1948 -1857 0 3
rlabel polysilicon 1955 -1851 1955 -1851 0 1
rlabel polysilicon 1955 -1857 1955 -1857 0 3
rlabel polysilicon 1962 -1851 1962 -1851 0 1
rlabel polysilicon 1962 -1857 1962 -1857 0 3
rlabel polysilicon 1969 -1851 1969 -1851 0 1
rlabel polysilicon 1969 -1857 1969 -1857 0 3
rlabel polysilicon 1976 -1851 1976 -1851 0 1
rlabel polysilicon 1976 -1857 1976 -1857 0 3
rlabel polysilicon 1983 -1851 1983 -1851 0 1
rlabel polysilicon 1983 -1857 1983 -1857 0 3
rlabel polysilicon 1990 -1851 1990 -1851 0 1
rlabel polysilicon 1990 -1857 1990 -1857 0 3
rlabel polysilicon 1997 -1851 1997 -1851 0 1
rlabel polysilicon 1997 -1857 1997 -1857 0 3
rlabel polysilicon 2004 -1851 2004 -1851 0 1
rlabel polysilicon 2004 -1857 2004 -1857 0 3
rlabel polysilicon 2011 -1851 2011 -1851 0 1
rlabel polysilicon 2011 -1857 2011 -1857 0 3
rlabel polysilicon 2018 -1851 2018 -1851 0 1
rlabel polysilicon 2018 -1857 2018 -1857 0 3
rlabel polysilicon 2025 -1851 2025 -1851 0 1
rlabel polysilicon 2025 -1857 2025 -1857 0 3
rlabel polysilicon 2032 -1851 2032 -1851 0 1
rlabel polysilicon 2032 -1857 2032 -1857 0 3
rlabel polysilicon 2039 -1851 2039 -1851 0 1
rlabel polysilicon 2042 -1851 2042 -1851 0 2
rlabel polysilicon 2039 -1857 2039 -1857 0 3
rlabel polysilicon 2046 -1851 2046 -1851 0 1
rlabel polysilicon 2046 -1857 2046 -1857 0 3
rlabel polysilicon 2053 -1851 2053 -1851 0 1
rlabel polysilicon 2053 -1857 2053 -1857 0 3
rlabel polysilicon 2060 -1851 2060 -1851 0 1
rlabel polysilicon 2060 -1857 2060 -1857 0 3
rlabel polysilicon 2067 -1851 2067 -1851 0 1
rlabel polysilicon 2067 -1857 2067 -1857 0 3
rlabel polysilicon 2074 -1851 2074 -1851 0 1
rlabel polysilicon 2074 -1857 2074 -1857 0 3
rlabel polysilicon 2081 -1851 2081 -1851 0 1
rlabel polysilicon 2081 -1857 2081 -1857 0 3
rlabel polysilicon 2088 -1851 2088 -1851 0 1
rlabel polysilicon 2088 -1857 2088 -1857 0 3
rlabel polysilicon 2095 -1851 2095 -1851 0 1
rlabel polysilicon 2095 -1857 2095 -1857 0 3
rlabel polysilicon 2102 -1851 2102 -1851 0 1
rlabel polysilicon 2102 -1857 2102 -1857 0 3
rlabel polysilicon 2109 -1851 2109 -1851 0 1
rlabel polysilicon 2109 -1857 2109 -1857 0 3
rlabel polysilicon 2116 -1851 2116 -1851 0 1
rlabel polysilicon 2116 -1857 2116 -1857 0 3
rlabel polysilicon 2123 -1851 2123 -1851 0 1
rlabel polysilicon 2123 -1857 2123 -1857 0 3
rlabel polysilicon 2130 -1851 2130 -1851 0 1
rlabel polysilicon 2130 -1857 2130 -1857 0 3
rlabel polysilicon 2137 -1851 2137 -1851 0 1
rlabel polysilicon 2137 -1857 2137 -1857 0 3
rlabel polysilicon 2144 -1851 2144 -1851 0 1
rlabel polysilicon 2144 -1857 2144 -1857 0 3
rlabel polysilicon 2151 -1851 2151 -1851 0 1
rlabel polysilicon 2151 -1857 2151 -1857 0 3
rlabel polysilicon 2158 -1851 2158 -1851 0 1
rlabel polysilicon 2158 -1857 2158 -1857 0 3
rlabel polysilicon 2165 -1851 2165 -1851 0 1
rlabel polysilicon 2165 -1857 2165 -1857 0 3
rlabel polysilicon 2172 -1851 2172 -1851 0 1
rlabel polysilicon 2172 -1857 2172 -1857 0 3
rlabel polysilicon 2179 -1851 2179 -1851 0 1
rlabel polysilicon 2179 -1857 2179 -1857 0 3
rlabel polysilicon 2186 -1851 2186 -1851 0 1
rlabel polysilicon 2186 -1857 2186 -1857 0 3
rlabel polysilicon 2193 -1851 2193 -1851 0 1
rlabel polysilicon 2193 -1857 2193 -1857 0 3
rlabel polysilicon 2200 -1851 2200 -1851 0 1
rlabel polysilicon 2200 -1857 2200 -1857 0 3
rlabel polysilicon 2207 -1851 2207 -1851 0 1
rlabel polysilicon 2207 -1857 2207 -1857 0 3
rlabel polysilicon 2214 -1851 2214 -1851 0 1
rlabel polysilicon 2214 -1857 2214 -1857 0 3
rlabel polysilicon 2221 -1851 2221 -1851 0 1
rlabel polysilicon 2221 -1857 2221 -1857 0 3
rlabel polysilicon 2228 -1851 2228 -1851 0 1
rlabel polysilicon 2228 -1857 2228 -1857 0 3
rlabel polysilicon 2235 -1851 2235 -1851 0 1
rlabel polysilicon 2235 -1857 2235 -1857 0 3
rlabel polysilicon 2242 -1851 2242 -1851 0 1
rlabel polysilicon 2242 -1857 2242 -1857 0 3
rlabel polysilicon 2249 -1851 2249 -1851 0 1
rlabel polysilicon 2249 -1857 2249 -1857 0 3
rlabel polysilicon 2256 -1851 2256 -1851 0 1
rlabel polysilicon 2256 -1857 2256 -1857 0 3
rlabel polysilicon 2263 -1851 2263 -1851 0 1
rlabel polysilicon 2263 -1857 2263 -1857 0 3
rlabel polysilicon 2270 -1851 2270 -1851 0 1
rlabel polysilicon 2270 -1857 2270 -1857 0 3
rlabel polysilicon 2277 -1851 2277 -1851 0 1
rlabel polysilicon 2277 -1857 2277 -1857 0 3
rlabel polysilicon 2284 -1851 2284 -1851 0 1
rlabel polysilicon 2284 -1857 2284 -1857 0 3
rlabel polysilicon 2291 -1851 2291 -1851 0 1
rlabel polysilicon 2291 -1857 2291 -1857 0 3
rlabel polysilicon 2298 -1851 2298 -1851 0 1
rlabel polysilicon 2298 -1857 2298 -1857 0 3
rlabel polysilicon 2305 -1851 2305 -1851 0 1
rlabel polysilicon 2305 -1857 2305 -1857 0 3
rlabel polysilicon 2312 -1851 2312 -1851 0 1
rlabel polysilicon 2312 -1857 2312 -1857 0 3
rlabel polysilicon 2319 -1851 2319 -1851 0 1
rlabel polysilicon 2319 -1857 2319 -1857 0 3
rlabel polysilicon 2326 -1851 2326 -1851 0 1
rlabel polysilicon 2326 -1857 2326 -1857 0 3
rlabel polysilicon 2333 -1851 2333 -1851 0 1
rlabel polysilicon 2333 -1857 2333 -1857 0 3
rlabel polysilicon 2340 -1851 2340 -1851 0 1
rlabel polysilicon 2340 -1857 2340 -1857 0 3
rlabel polysilicon 2347 -1851 2347 -1851 0 1
rlabel polysilicon 2347 -1857 2347 -1857 0 3
rlabel polysilicon 2354 -1851 2354 -1851 0 1
rlabel polysilicon 2354 -1857 2354 -1857 0 3
rlabel polysilicon 2361 -1851 2361 -1851 0 1
rlabel polysilicon 2361 -1857 2361 -1857 0 3
rlabel polysilicon 2368 -1851 2368 -1851 0 1
rlabel polysilicon 2368 -1857 2368 -1857 0 3
rlabel polysilicon 2375 -1851 2375 -1851 0 1
rlabel polysilicon 2375 -1857 2375 -1857 0 3
rlabel polysilicon 2382 -1851 2382 -1851 0 1
rlabel polysilicon 2382 -1857 2382 -1857 0 3
rlabel polysilicon 2389 -1851 2389 -1851 0 1
rlabel polysilicon 2389 -1857 2389 -1857 0 3
rlabel polysilicon 2396 -1851 2396 -1851 0 1
rlabel polysilicon 2396 -1857 2396 -1857 0 3
rlabel polysilicon 2403 -1851 2403 -1851 0 1
rlabel polysilicon 2403 -1857 2403 -1857 0 3
rlabel polysilicon 2410 -1851 2410 -1851 0 1
rlabel polysilicon 2410 -1857 2410 -1857 0 3
rlabel polysilicon 2417 -1851 2417 -1851 0 1
rlabel polysilicon 2417 -1857 2417 -1857 0 3
rlabel polysilicon 2424 -1851 2424 -1851 0 1
rlabel polysilicon 2424 -1857 2424 -1857 0 3
rlabel polysilicon 2431 -1851 2431 -1851 0 1
rlabel polysilicon 2431 -1857 2431 -1857 0 3
rlabel polysilicon 2438 -1851 2438 -1851 0 1
rlabel polysilicon 2438 -1857 2438 -1857 0 3
rlabel polysilicon 2445 -1851 2445 -1851 0 1
rlabel polysilicon 2445 -1857 2445 -1857 0 3
rlabel polysilicon 2452 -1851 2452 -1851 0 1
rlabel polysilicon 2452 -1857 2452 -1857 0 3
rlabel polysilicon 2459 -1851 2459 -1851 0 1
rlabel polysilicon 2459 -1857 2459 -1857 0 3
rlabel polysilicon 2466 -1851 2466 -1851 0 1
rlabel polysilicon 2469 -1851 2469 -1851 0 2
rlabel polysilicon 2466 -1857 2466 -1857 0 3
rlabel polysilicon 2469 -1857 2469 -1857 0 4
rlabel polysilicon 2473 -1851 2473 -1851 0 1
rlabel polysilicon 2476 -1851 2476 -1851 0 2
rlabel polysilicon 2473 -1857 2473 -1857 0 3
rlabel polysilicon 2 -2026 2 -2026 0 1
rlabel polysilicon 2 -2032 2 -2032 0 3
rlabel polysilicon 9 -2026 9 -2026 0 1
rlabel polysilicon 9 -2032 9 -2032 0 3
rlabel polysilicon 16 -2026 16 -2026 0 1
rlabel polysilicon 16 -2032 16 -2032 0 3
rlabel polysilicon 23 -2026 23 -2026 0 1
rlabel polysilicon 23 -2032 23 -2032 0 3
rlabel polysilicon 30 -2026 30 -2026 0 1
rlabel polysilicon 30 -2032 30 -2032 0 3
rlabel polysilicon 37 -2026 37 -2026 0 1
rlabel polysilicon 37 -2032 37 -2032 0 3
rlabel polysilicon 44 -2026 44 -2026 0 1
rlabel polysilicon 44 -2032 44 -2032 0 3
rlabel polysilicon 51 -2026 51 -2026 0 1
rlabel polysilicon 51 -2032 51 -2032 0 3
rlabel polysilicon 54 -2032 54 -2032 0 4
rlabel polysilicon 58 -2026 58 -2026 0 1
rlabel polysilicon 58 -2032 58 -2032 0 3
rlabel polysilicon 65 -2026 65 -2026 0 1
rlabel polysilicon 65 -2032 65 -2032 0 3
rlabel polysilicon 72 -2026 72 -2026 0 1
rlabel polysilicon 72 -2032 72 -2032 0 3
rlabel polysilicon 79 -2026 79 -2026 0 1
rlabel polysilicon 79 -2032 79 -2032 0 3
rlabel polysilicon 86 -2026 86 -2026 0 1
rlabel polysilicon 89 -2026 89 -2026 0 2
rlabel polysilicon 89 -2032 89 -2032 0 4
rlabel polysilicon 93 -2026 93 -2026 0 1
rlabel polysilicon 93 -2032 93 -2032 0 3
rlabel polysilicon 100 -2026 100 -2026 0 1
rlabel polysilicon 103 -2026 103 -2026 0 2
rlabel polysilicon 100 -2032 100 -2032 0 3
rlabel polysilicon 103 -2032 103 -2032 0 4
rlabel polysilicon 107 -2026 107 -2026 0 1
rlabel polysilicon 107 -2032 107 -2032 0 3
rlabel polysilicon 114 -2026 114 -2026 0 1
rlabel polysilicon 114 -2032 114 -2032 0 3
rlabel polysilicon 121 -2026 121 -2026 0 1
rlabel polysilicon 121 -2032 121 -2032 0 3
rlabel polysilicon 128 -2026 128 -2026 0 1
rlabel polysilicon 131 -2026 131 -2026 0 2
rlabel polysilicon 131 -2032 131 -2032 0 4
rlabel polysilicon 135 -2026 135 -2026 0 1
rlabel polysilicon 135 -2032 135 -2032 0 3
rlabel polysilicon 142 -2026 142 -2026 0 1
rlabel polysilicon 142 -2032 142 -2032 0 3
rlabel polysilicon 149 -2026 149 -2026 0 1
rlabel polysilicon 149 -2032 149 -2032 0 3
rlabel polysilicon 156 -2026 156 -2026 0 1
rlabel polysilicon 159 -2026 159 -2026 0 2
rlabel polysilicon 156 -2032 156 -2032 0 3
rlabel polysilicon 159 -2032 159 -2032 0 4
rlabel polysilicon 163 -2026 163 -2026 0 1
rlabel polysilicon 163 -2032 163 -2032 0 3
rlabel polysilicon 170 -2026 170 -2026 0 1
rlabel polysilicon 173 -2026 173 -2026 0 2
rlabel polysilicon 170 -2032 170 -2032 0 3
rlabel polysilicon 173 -2032 173 -2032 0 4
rlabel polysilicon 177 -2026 177 -2026 0 1
rlabel polysilicon 177 -2032 177 -2032 0 3
rlabel polysilicon 184 -2026 184 -2026 0 1
rlabel polysilicon 184 -2032 184 -2032 0 3
rlabel polysilicon 191 -2026 191 -2026 0 1
rlabel polysilicon 194 -2026 194 -2026 0 2
rlabel polysilicon 191 -2032 191 -2032 0 3
rlabel polysilicon 194 -2032 194 -2032 0 4
rlabel polysilicon 198 -2026 198 -2026 0 1
rlabel polysilicon 198 -2032 198 -2032 0 3
rlabel polysilicon 205 -2026 205 -2026 0 1
rlabel polysilicon 205 -2032 205 -2032 0 3
rlabel polysilicon 212 -2026 212 -2026 0 1
rlabel polysilicon 215 -2026 215 -2026 0 2
rlabel polysilicon 212 -2032 212 -2032 0 3
rlabel polysilicon 215 -2032 215 -2032 0 4
rlabel polysilicon 219 -2026 219 -2026 0 1
rlabel polysilicon 219 -2032 219 -2032 0 3
rlabel polysilicon 226 -2026 226 -2026 0 1
rlabel polysilicon 226 -2032 226 -2032 0 3
rlabel polysilicon 233 -2026 233 -2026 0 1
rlabel polysilicon 233 -2032 233 -2032 0 3
rlabel polysilicon 240 -2026 240 -2026 0 1
rlabel polysilicon 240 -2032 240 -2032 0 3
rlabel polysilicon 247 -2026 247 -2026 0 1
rlabel polysilicon 247 -2032 247 -2032 0 3
rlabel polysilicon 254 -2026 254 -2026 0 1
rlabel polysilicon 254 -2032 254 -2032 0 3
rlabel polysilicon 261 -2026 261 -2026 0 1
rlabel polysilicon 261 -2032 261 -2032 0 3
rlabel polysilicon 268 -2026 268 -2026 0 1
rlabel polysilicon 268 -2032 268 -2032 0 3
rlabel polysilicon 275 -2026 275 -2026 0 1
rlabel polysilicon 275 -2032 275 -2032 0 3
rlabel polysilicon 282 -2026 282 -2026 0 1
rlabel polysilicon 282 -2032 282 -2032 0 3
rlabel polysilicon 289 -2026 289 -2026 0 1
rlabel polysilicon 289 -2032 289 -2032 0 3
rlabel polysilicon 296 -2026 296 -2026 0 1
rlabel polysilicon 296 -2032 296 -2032 0 3
rlabel polysilicon 303 -2026 303 -2026 0 1
rlabel polysilicon 303 -2032 303 -2032 0 3
rlabel polysilicon 310 -2026 310 -2026 0 1
rlabel polysilicon 310 -2032 310 -2032 0 3
rlabel polysilicon 317 -2026 317 -2026 0 1
rlabel polysilicon 317 -2032 317 -2032 0 3
rlabel polysilicon 324 -2026 324 -2026 0 1
rlabel polysilicon 324 -2032 324 -2032 0 3
rlabel polysilicon 331 -2026 331 -2026 0 1
rlabel polysilicon 331 -2032 331 -2032 0 3
rlabel polysilicon 338 -2026 338 -2026 0 1
rlabel polysilicon 338 -2032 338 -2032 0 3
rlabel polysilicon 345 -2026 345 -2026 0 1
rlabel polysilicon 345 -2032 345 -2032 0 3
rlabel polysilicon 352 -2026 352 -2026 0 1
rlabel polysilicon 352 -2032 352 -2032 0 3
rlabel polysilicon 359 -2026 359 -2026 0 1
rlabel polysilicon 359 -2032 359 -2032 0 3
rlabel polysilicon 366 -2026 366 -2026 0 1
rlabel polysilicon 366 -2032 366 -2032 0 3
rlabel polysilicon 373 -2026 373 -2026 0 1
rlabel polysilicon 373 -2032 373 -2032 0 3
rlabel polysilicon 380 -2026 380 -2026 0 1
rlabel polysilicon 380 -2032 380 -2032 0 3
rlabel polysilicon 387 -2026 387 -2026 0 1
rlabel polysilicon 387 -2032 387 -2032 0 3
rlabel polysilicon 394 -2026 394 -2026 0 1
rlabel polysilicon 394 -2032 394 -2032 0 3
rlabel polysilicon 401 -2026 401 -2026 0 1
rlabel polysilicon 401 -2032 401 -2032 0 3
rlabel polysilicon 408 -2026 408 -2026 0 1
rlabel polysilicon 408 -2032 408 -2032 0 3
rlabel polysilicon 415 -2026 415 -2026 0 1
rlabel polysilicon 415 -2032 415 -2032 0 3
rlabel polysilicon 422 -2026 422 -2026 0 1
rlabel polysilicon 422 -2032 422 -2032 0 3
rlabel polysilicon 429 -2026 429 -2026 0 1
rlabel polysilicon 429 -2032 429 -2032 0 3
rlabel polysilicon 436 -2026 436 -2026 0 1
rlabel polysilicon 436 -2032 436 -2032 0 3
rlabel polysilicon 443 -2026 443 -2026 0 1
rlabel polysilicon 443 -2032 443 -2032 0 3
rlabel polysilicon 450 -2026 450 -2026 0 1
rlabel polysilicon 450 -2032 450 -2032 0 3
rlabel polysilicon 457 -2026 457 -2026 0 1
rlabel polysilicon 457 -2032 457 -2032 0 3
rlabel polysilicon 464 -2026 464 -2026 0 1
rlabel polysilicon 464 -2032 464 -2032 0 3
rlabel polysilicon 471 -2026 471 -2026 0 1
rlabel polysilicon 471 -2032 471 -2032 0 3
rlabel polysilicon 478 -2026 478 -2026 0 1
rlabel polysilicon 478 -2032 478 -2032 0 3
rlabel polysilicon 485 -2026 485 -2026 0 1
rlabel polysilicon 485 -2032 485 -2032 0 3
rlabel polysilicon 492 -2026 492 -2026 0 1
rlabel polysilicon 492 -2032 492 -2032 0 3
rlabel polysilicon 499 -2026 499 -2026 0 1
rlabel polysilicon 499 -2032 499 -2032 0 3
rlabel polysilicon 506 -2026 506 -2026 0 1
rlabel polysilicon 506 -2032 506 -2032 0 3
rlabel polysilicon 513 -2026 513 -2026 0 1
rlabel polysilicon 513 -2032 513 -2032 0 3
rlabel polysilicon 520 -2026 520 -2026 0 1
rlabel polysilicon 520 -2032 520 -2032 0 3
rlabel polysilicon 527 -2026 527 -2026 0 1
rlabel polysilicon 527 -2032 527 -2032 0 3
rlabel polysilicon 534 -2026 534 -2026 0 1
rlabel polysilicon 534 -2032 534 -2032 0 3
rlabel polysilicon 541 -2026 541 -2026 0 1
rlabel polysilicon 544 -2026 544 -2026 0 2
rlabel polysilicon 548 -2026 548 -2026 0 1
rlabel polysilicon 548 -2032 548 -2032 0 3
rlabel polysilicon 555 -2026 555 -2026 0 1
rlabel polysilicon 555 -2032 555 -2032 0 3
rlabel polysilicon 562 -2026 562 -2026 0 1
rlabel polysilicon 562 -2032 562 -2032 0 3
rlabel polysilicon 569 -2026 569 -2026 0 1
rlabel polysilicon 569 -2032 569 -2032 0 3
rlabel polysilicon 576 -2026 576 -2026 0 1
rlabel polysilicon 576 -2032 576 -2032 0 3
rlabel polysilicon 583 -2026 583 -2026 0 1
rlabel polysilicon 586 -2026 586 -2026 0 2
rlabel polysilicon 586 -2032 586 -2032 0 4
rlabel polysilicon 590 -2026 590 -2026 0 1
rlabel polysilicon 590 -2032 590 -2032 0 3
rlabel polysilicon 597 -2026 597 -2026 0 1
rlabel polysilicon 597 -2032 597 -2032 0 3
rlabel polysilicon 604 -2026 604 -2026 0 1
rlabel polysilicon 604 -2032 604 -2032 0 3
rlabel polysilicon 611 -2026 611 -2026 0 1
rlabel polysilicon 611 -2032 611 -2032 0 3
rlabel polysilicon 618 -2026 618 -2026 0 1
rlabel polysilicon 618 -2032 618 -2032 0 3
rlabel polysilicon 625 -2026 625 -2026 0 1
rlabel polysilicon 625 -2032 625 -2032 0 3
rlabel polysilicon 632 -2026 632 -2026 0 1
rlabel polysilicon 635 -2026 635 -2026 0 2
rlabel polysilicon 632 -2032 632 -2032 0 3
rlabel polysilicon 639 -2026 639 -2026 0 1
rlabel polysilicon 639 -2032 639 -2032 0 3
rlabel polysilicon 646 -2026 646 -2026 0 1
rlabel polysilicon 646 -2032 646 -2032 0 3
rlabel polysilicon 653 -2026 653 -2026 0 1
rlabel polysilicon 653 -2032 653 -2032 0 3
rlabel polysilicon 660 -2026 660 -2026 0 1
rlabel polysilicon 660 -2032 660 -2032 0 3
rlabel polysilicon 667 -2026 667 -2026 0 1
rlabel polysilicon 667 -2032 667 -2032 0 3
rlabel polysilicon 674 -2026 674 -2026 0 1
rlabel polysilicon 674 -2032 674 -2032 0 3
rlabel polysilicon 681 -2026 681 -2026 0 1
rlabel polysilicon 681 -2032 681 -2032 0 3
rlabel polysilicon 688 -2026 688 -2026 0 1
rlabel polysilicon 688 -2032 688 -2032 0 3
rlabel polysilicon 695 -2026 695 -2026 0 1
rlabel polysilicon 695 -2032 695 -2032 0 3
rlabel polysilicon 702 -2026 702 -2026 0 1
rlabel polysilicon 702 -2032 702 -2032 0 3
rlabel polysilicon 709 -2026 709 -2026 0 1
rlabel polysilicon 709 -2032 709 -2032 0 3
rlabel polysilicon 716 -2026 716 -2026 0 1
rlabel polysilicon 716 -2032 716 -2032 0 3
rlabel polysilicon 723 -2026 723 -2026 0 1
rlabel polysilicon 723 -2032 723 -2032 0 3
rlabel polysilicon 730 -2026 730 -2026 0 1
rlabel polysilicon 730 -2032 730 -2032 0 3
rlabel polysilicon 737 -2026 737 -2026 0 1
rlabel polysilicon 740 -2026 740 -2026 0 2
rlabel polysilicon 737 -2032 737 -2032 0 3
rlabel polysilicon 740 -2032 740 -2032 0 4
rlabel polysilicon 744 -2026 744 -2026 0 1
rlabel polysilicon 744 -2032 744 -2032 0 3
rlabel polysilicon 751 -2026 751 -2026 0 1
rlabel polysilicon 751 -2032 751 -2032 0 3
rlabel polysilicon 758 -2026 758 -2026 0 1
rlabel polysilicon 758 -2032 758 -2032 0 3
rlabel polysilicon 765 -2026 765 -2026 0 1
rlabel polysilicon 765 -2032 765 -2032 0 3
rlabel polysilicon 772 -2026 772 -2026 0 1
rlabel polysilicon 772 -2032 772 -2032 0 3
rlabel polysilicon 779 -2026 779 -2026 0 1
rlabel polysilicon 782 -2026 782 -2026 0 2
rlabel polysilicon 779 -2032 779 -2032 0 3
rlabel polysilicon 786 -2026 786 -2026 0 1
rlabel polysilicon 786 -2032 786 -2032 0 3
rlabel polysilicon 793 -2026 793 -2026 0 1
rlabel polysilicon 793 -2032 793 -2032 0 3
rlabel polysilicon 800 -2032 800 -2032 0 3
rlabel polysilicon 803 -2032 803 -2032 0 4
rlabel polysilicon 807 -2026 807 -2026 0 1
rlabel polysilicon 807 -2032 807 -2032 0 3
rlabel polysilicon 814 -2026 814 -2026 0 1
rlabel polysilicon 814 -2032 814 -2032 0 3
rlabel polysilicon 821 -2026 821 -2026 0 1
rlabel polysilicon 821 -2032 821 -2032 0 3
rlabel polysilicon 828 -2026 828 -2026 0 1
rlabel polysilicon 831 -2026 831 -2026 0 2
rlabel polysilicon 828 -2032 828 -2032 0 3
rlabel polysilicon 831 -2032 831 -2032 0 4
rlabel polysilicon 835 -2026 835 -2026 0 1
rlabel polysilicon 835 -2032 835 -2032 0 3
rlabel polysilicon 842 -2026 842 -2026 0 1
rlabel polysilicon 842 -2032 842 -2032 0 3
rlabel polysilicon 849 -2026 849 -2026 0 1
rlabel polysilicon 849 -2032 849 -2032 0 3
rlabel polysilicon 856 -2026 856 -2026 0 1
rlabel polysilicon 856 -2032 856 -2032 0 3
rlabel polysilicon 863 -2026 863 -2026 0 1
rlabel polysilicon 863 -2032 863 -2032 0 3
rlabel polysilicon 870 -2026 870 -2026 0 1
rlabel polysilicon 870 -2032 870 -2032 0 3
rlabel polysilicon 877 -2026 877 -2026 0 1
rlabel polysilicon 877 -2032 877 -2032 0 3
rlabel polysilicon 884 -2026 884 -2026 0 1
rlabel polysilicon 884 -2032 884 -2032 0 3
rlabel polysilicon 891 -2026 891 -2026 0 1
rlabel polysilicon 891 -2032 891 -2032 0 3
rlabel polysilicon 898 -2026 898 -2026 0 1
rlabel polysilicon 898 -2032 898 -2032 0 3
rlabel polysilicon 905 -2026 905 -2026 0 1
rlabel polysilicon 905 -2032 905 -2032 0 3
rlabel polysilicon 912 -2026 912 -2026 0 1
rlabel polysilicon 912 -2032 912 -2032 0 3
rlabel polysilicon 919 -2026 919 -2026 0 1
rlabel polysilicon 922 -2026 922 -2026 0 2
rlabel polysilicon 919 -2032 919 -2032 0 3
rlabel polysilicon 922 -2032 922 -2032 0 4
rlabel polysilicon 926 -2026 926 -2026 0 1
rlabel polysilicon 926 -2032 926 -2032 0 3
rlabel polysilicon 933 -2026 933 -2026 0 1
rlabel polysilicon 933 -2032 933 -2032 0 3
rlabel polysilicon 940 -2026 940 -2026 0 1
rlabel polysilicon 940 -2032 940 -2032 0 3
rlabel polysilicon 947 -2026 947 -2026 0 1
rlabel polysilicon 947 -2032 947 -2032 0 3
rlabel polysilicon 954 -2026 954 -2026 0 1
rlabel polysilicon 957 -2026 957 -2026 0 2
rlabel polysilicon 954 -2032 954 -2032 0 3
rlabel polysilicon 957 -2032 957 -2032 0 4
rlabel polysilicon 961 -2026 961 -2026 0 1
rlabel polysilicon 961 -2032 961 -2032 0 3
rlabel polysilicon 968 -2026 968 -2026 0 1
rlabel polysilicon 968 -2032 968 -2032 0 3
rlabel polysilicon 975 -2026 975 -2026 0 1
rlabel polysilicon 978 -2026 978 -2026 0 2
rlabel polysilicon 978 -2032 978 -2032 0 4
rlabel polysilicon 982 -2026 982 -2026 0 1
rlabel polysilicon 982 -2032 982 -2032 0 3
rlabel polysilicon 989 -2026 989 -2026 0 1
rlabel polysilicon 989 -2032 989 -2032 0 3
rlabel polysilicon 996 -2026 996 -2026 0 1
rlabel polysilicon 996 -2032 996 -2032 0 3
rlabel polysilicon 1003 -2026 1003 -2026 0 1
rlabel polysilicon 1003 -2032 1003 -2032 0 3
rlabel polysilicon 1010 -2026 1010 -2026 0 1
rlabel polysilicon 1010 -2032 1010 -2032 0 3
rlabel polysilicon 1017 -2026 1017 -2026 0 1
rlabel polysilicon 1017 -2032 1017 -2032 0 3
rlabel polysilicon 1024 -2026 1024 -2026 0 1
rlabel polysilicon 1024 -2032 1024 -2032 0 3
rlabel polysilicon 1031 -2026 1031 -2026 0 1
rlabel polysilicon 1031 -2032 1031 -2032 0 3
rlabel polysilicon 1038 -2026 1038 -2026 0 1
rlabel polysilicon 1038 -2032 1038 -2032 0 3
rlabel polysilicon 1045 -2026 1045 -2026 0 1
rlabel polysilicon 1045 -2032 1045 -2032 0 3
rlabel polysilicon 1052 -2026 1052 -2026 0 1
rlabel polysilicon 1052 -2032 1052 -2032 0 3
rlabel polysilicon 1059 -2026 1059 -2026 0 1
rlabel polysilicon 1062 -2026 1062 -2026 0 2
rlabel polysilicon 1059 -2032 1059 -2032 0 3
rlabel polysilicon 1062 -2032 1062 -2032 0 4
rlabel polysilicon 1066 -2026 1066 -2026 0 1
rlabel polysilicon 1066 -2032 1066 -2032 0 3
rlabel polysilicon 1073 -2026 1073 -2026 0 1
rlabel polysilicon 1073 -2032 1073 -2032 0 3
rlabel polysilicon 1080 -2026 1080 -2026 0 1
rlabel polysilicon 1080 -2032 1080 -2032 0 3
rlabel polysilicon 1087 -2026 1087 -2026 0 1
rlabel polysilicon 1087 -2032 1087 -2032 0 3
rlabel polysilicon 1094 -2026 1094 -2026 0 1
rlabel polysilicon 1094 -2032 1094 -2032 0 3
rlabel polysilicon 1101 -2026 1101 -2026 0 1
rlabel polysilicon 1101 -2032 1101 -2032 0 3
rlabel polysilicon 1108 -2026 1108 -2026 0 1
rlabel polysilicon 1111 -2026 1111 -2026 0 2
rlabel polysilicon 1108 -2032 1108 -2032 0 3
rlabel polysilicon 1111 -2032 1111 -2032 0 4
rlabel polysilicon 1115 -2026 1115 -2026 0 1
rlabel polysilicon 1115 -2032 1115 -2032 0 3
rlabel polysilicon 1125 -2026 1125 -2026 0 2
rlabel polysilicon 1122 -2032 1122 -2032 0 3
rlabel polysilicon 1125 -2032 1125 -2032 0 4
rlabel polysilicon 1129 -2026 1129 -2026 0 1
rlabel polysilicon 1129 -2032 1129 -2032 0 3
rlabel polysilicon 1136 -2026 1136 -2026 0 1
rlabel polysilicon 1136 -2032 1136 -2032 0 3
rlabel polysilicon 1143 -2026 1143 -2026 0 1
rlabel polysilicon 1143 -2032 1143 -2032 0 3
rlabel polysilicon 1153 -2026 1153 -2026 0 2
rlabel polysilicon 1153 -2032 1153 -2032 0 4
rlabel polysilicon 1157 -2026 1157 -2026 0 1
rlabel polysilicon 1157 -2032 1157 -2032 0 3
rlabel polysilicon 1164 -2026 1164 -2026 0 1
rlabel polysilicon 1167 -2026 1167 -2026 0 2
rlabel polysilicon 1164 -2032 1164 -2032 0 3
rlabel polysilicon 1167 -2032 1167 -2032 0 4
rlabel polysilicon 1171 -2026 1171 -2026 0 1
rlabel polysilicon 1171 -2032 1171 -2032 0 3
rlabel polysilicon 1178 -2026 1178 -2026 0 1
rlabel polysilicon 1178 -2032 1178 -2032 0 3
rlabel polysilicon 1185 -2026 1185 -2026 0 1
rlabel polysilicon 1185 -2032 1185 -2032 0 3
rlabel polysilicon 1188 -2032 1188 -2032 0 4
rlabel polysilicon 1192 -2026 1192 -2026 0 1
rlabel polysilicon 1192 -2032 1192 -2032 0 3
rlabel polysilicon 1199 -2026 1199 -2026 0 1
rlabel polysilicon 1199 -2032 1199 -2032 0 3
rlabel polysilicon 1206 -2026 1206 -2026 0 1
rlabel polysilicon 1206 -2032 1206 -2032 0 3
rlabel polysilicon 1213 -2026 1213 -2026 0 1
rlabel polysilicon 1213 -2032 1213 -2032 0 3
rlabel polysilicon 1220 -2026 1220 -2026 0 1
rlabel polysilicon 1220 -2032 1220 -2032 0 3
rlabel polysilicon 1227 -2026 1227 -2026 0 1
rlabel polysilicon 1230 -2032 1230 -2032 0 4
rlabel polysilicon 1234 -2026 1234 -2026 0 1
rlabel polysilicon 1234 -2032 1234 -2032 0 3
rlabel polysilicon 1241 -2026 1241 -2026 0 1
rlabel polysilicon 1241 -2032 1241 -2032 0 3
rlabel polysilicon 1248 -2026 1248 -2026 0 1
rlabel polysilicon 1248 -2032 1248 -2032 0 3
rlabel polysilicon 1255 -2026 1255 -2026 0 1
rlabel polysilicon 1255 -2032 1255 -2032 0 3
rlabel polysilicon 1262 -2026 1262 -2026 0 1
rlabel polysilicon 1262 -2032 1262 -2032 0 3
rlabel polysilicon 1269 -2026 1269 -2026 0 1
rlabel polysilicon 1269 -2032 1269 -2032 0 3
rlabel polysilicon 1276 -2026 1276 -2026 0 1
rlabel polysilicon 1276 -2032 1276 -2032 0 3
rlabel polysilicon 1283 -2026 1283 -2026 0 1
rlabel polysilicon 1283 -2032 1283 -2032 0 3
rlabel polysilicon 1290 -2026 1290 -2026 0 1
rlabel polysilicon 1290 -2032 1290 -2032 0 3
rlabel polysilicon 1297 -2026 1297 -2026 0 1
rlabel polysilicon 1300 -2026 1300 -2026 0 2
rlabel polysilicon 1297 -2032 1297 -2032 0 3
rlabel polysilicon 1300 -2032 1300 -2032 0 4
rlabel polysilicon 1304 -2026 1304 -2026 0 1
rlabel polysilicon 1304 -2032 1304 -2032 0 3
rlabel polysilicon 1311 -2026 1311 -2026 0 1
rlabel polysilicon 1311 -2032 1311 -2032 0 3
rlabel polysilicon 1318 -2026 1318 -2026 0 1
rlabel polysilicon 1318 -2032 1318 -2032 0 3
rlabel polysilicon 1325 -2032 1325 -2032 0 3
rlabel polysilicon 1332 -2026 1332 -2026 0 1
rlabel polysilicon 1335 -2026 1335 -2026 0 2
rlabel polysilicon 1332 -2032 1332 -2032 0 3
rlabel polysilicon 1339 -2026 1339 -2026 0 1
rlabel polysilicon 1339 -2032 1339 -2032 0 3
rlabel polysilicon 1346 -2026 1346 -2026 0 1
rlabel polysilicon 1346 -2032 1346 -2032 0 3
rlabel polysilicon 1353 -2026 1353 -2026 0 1
rlabel polysilicon 1353 -2032 1353 -2032 0 3
rlabel polysilicon 1360 -2026 1360 -2026 0 1
rlabel polysilicon 1363 -2026 1363 -2026 0 2
rlabel polysilicon 1360 -2032 1360 -2032 0 3
rlabel polysilicon 1363 -2032 1363 -2032 0 4
rlabel polysilicon 1367 -2026 1367 -2026 0 1
rlabel polysilicon 1367 -2032 1367 -2032 0 3
rlabel polysilicon 1374 -2026 1374 -2026 0 1
rlabel polysilicon 1374 -2032 1374 -2032 0 3
rlabel polysilicon 1381 -2026 1381 -2026 0 1
rlabel polysilicon 1381 -2032 1381 -2032 0 3
rlabel polysilicon 1388 -2026 1388 -2026 0 1
rlabel polysilicon 1388 -2032 1388 -2032 0 3
rlabel polysilicon 1395 -2026 1395 -2026 0 1
rlabel polysilicon 1395 -2032 1395 -2032 0 3
rlabel polysilicon 1402 -2026 1402 -2026 0 1
rlabel polysilicon 1402 -2032 1402 -2032 0 3
rlabel polysilicon 1409 -2026 1409 -2026 0 1
rlabel polysilicon 1409 -2032 1409 -2032 0 3
rlabel polysilicon 1416 -2026 1416 -2026 0 1
rlabel polysilicon 1416 -2032 1416 -2032 0 3
rlabel polysilicon 1423 -2026 1423 -2026 0 1
rlabel polysilicon 1423 -2032 1423 -2032 0 3
rlabel polysilicon 1430 -2026 1430 -2026 0 1
rlabel polysilicon 1430 -2032 1430 -2032 0 3
rlabel polysilicon 1437 -2026 1437 -2026 0 1
rlabel polysilicon 1440 -2026 1440 -2026 0 2
rlabel polysilicon 1437 -2032 1437 -2032 0 3
rlabel polysilicon 1440 -2032 1440 -2032 0 4
rlabel polysilicon 1444 -2026 1444 -2026 0 1
rlabel polysilicon 1444 -2032 1444 -2032 0 3
rlabel polysilicon 1451 -2026 1451 -2026 0 1
rlabel polysilicon 1451 -2032 1451 -2032 0 3
rlabel polysilicon 1458 -2026 1458 -2026 0 1
rlabel polysilicon 1458 -2032 1458 -2032 0 3
rlabel polysilicon 1465 -2026 1465 -2026 0 1
rlabel polysilicon 1465 -2032 1465 -2032 0 3
rlabel polysilicon 1472 -2026 1472 -2026 0 1
rlabel polysilicon 1475 -2026 1475 -2026 0 2
rlabel polysilicon 1475 -2032 1475 -2032 0 4
rlabel polysilicon 1479 -2026 1479 -2026 0 1
rlabel polysilicon 1479 -2032 1479 -2032 0 3
rlabel polysilicon 1486 -2026 1486 -2026 0 1
rlabel polysilicon 1489 -2026 1489 -2026 0 2
rlabel polysilicon 1486 -2032 1486 -2032 0 3
rlabel polysilicon 1489 -2032 1489 -2032 0 4
rlabel polysilicon 1493 -2026 1493 -2026 0 1
rlabel polysilicon 1496 -2026 1496 -2026 0 2
rlabel polysilicon 1493 -2032 1493 -2032 0 3
rlabel polysilicon 1496 -2032 1496 -2032 0 4
rlabel polysilicon 1500 -2026 1500 -2026 0 1
rlabel polysilicon 1500 -2032 1500 -2032 0 3
rlabel polysilicon 1507 -2026 1507 -2026 0 1
rlabel polysilicon 1507 -2032 1507 -2032 0 3
rlabel polysilicon 1514 -2026 1514 -2026 0 1
rlabel polysilicon 1514 -2032 1514 -2032 0 3
rlabel polysilicon 1524 -2026 1524 -2026 0 2
rlabel polysilicon 1521 -2032 1521 -2032 0 3
rlabel polysilicon 1528 -2026 1528 -2026 0 1
rlabel polysilicon 1528 -2032 1528 -2032 0 3
rlabel polysilicon 1535 -2026 1535 -2026 0 1
rlabel polysilicon 1535 -2032 1535 -2032 0 3
rlabel polysilicon 1538 -2032 1538 -2032 0 4
rlabel polysilicon 1542 -2026 1542 -2026 0 1
rlabel polysilicon 1542 -2032 1542 -2032 0 3
rlabel polysilicon 1549 -2026 1549 -2026 0 1
rlabel polysilicon 1549 -2032 1549 -2032 0 3
rlabel polysilicon 1552 -2032 1552 -2032 0 4
rlabel polysilicon 1556 -2026 1556 -2026 0 1
rlabel polysilicon 1556 -2032 1556 -2032 0 3
rlabel polysilicon 1563 -2026 1563 -2026 0 1
rlabel polysilicon 1563 -2032 1563 -2032 0 3
rlabel polysilicon 1570 -2026 1570 -2026 0 1
rlabel polysilicon 1570 -2032 1570 -2032 0 3
rlabel polysilicon 1577 -2026 1577 -2026 0 1
rlabel polysilicon 1577 -2032 1577 -2032 0 3
rlabel polysilicon 1584 -2026 1584 -2026 0 1
rlabel polysilicon 1584 -2032 1584 -2032 0 3
rlabel polysilicon 1591 -2026 1591 -2026 0 1
rlabel polysilicon 1591 -2032 1591 -2032 0 3
rlabel polysilicon 1598 -2026 1598 -2026 0 1
rlabel polysilicon 1598 -2032 1598 -2032 0 3
rlabel polysilicon 1605 -2026 1605 -2026 0 1
rlabel polysilicon 1605 -2032 1605 -2032 0 3
rlabel polysilicon 1612 -2026 1612 -2026 0 1
rlabel polysilicon 1612 -2032 1612 -2032 0 3
rlabel polysilicon 1619 -2026 1619 -2026 0 1
rlabel polysilicon 1622 -2026 1622 -2026 0 2
rlabel polysilicon 1619 -2032 1619 -2032 0 3
rlabel polysilicon 1622 -2032 1622 -2032 0 4
rlabel polysilicon 1626 -2026 1626 -2026 0 1
rlabel polysilicon 1626 -2032 1626 -2032 0 3
rlabel polysilicon 1633 -2026 1633 -2026 0 1
rlabel polysilicon 1636 -2026 1636 -2026 0 2
rlabel polysilicon 1633 -2032 1633 -2032 0 3
rlabel polysilicon 1636 -2032 1636 -2032 0 4
rlabel polysilicon 1640 -2026 1640 -2026 0 1
rlabel polysilicon 1640 -2032 1640 -2032 0 3
rlabel polysilicon 1647 -2026 1647 -2026 0 1
rlabel polysilicon 1647 -2032 1647 -2032 0 3
rlabel polysilicon 1654 -2026 1654 -2026 0 1
rlabel polysilicon 1654 -2032 1654 -2032 0 3
rlabel polysilicon 1661 -2026 1661 -2026 0 1
rlabel polysilicon 1664 -2026 1664 -2026 0 2
rlabel polysilicon 1661 -2032 1661 -2032 0 3
rlabel polysilicon 1664 -2032 1664 -2032 0 4
rlabel polysilicon 1668 -2026 1668 -2026 0 1
rlabel polysilicon 1668 -2032 1668 -2032 0 3
rlabel polysilicon 1675 -2026 1675 -2026 0 1
rlabel polysilicon 1675 -2032 1675 -2032 0 3
rlabel polysilicon 1682 -2026 1682 -2026 0 1
rlabel polysilicon 1682 -2032 1682 -2032 0 3
rlabel polysilicon 1689 -2026 1689 -2026 0 1
rlabel polysilicon 1689 -2032 1689 -2032 0 3
rlabel polysilicon 1696 -2026 1696 -2026 0 1
rlabel polysilicon 1696 -2032 1696 -2032 0 3
rlabel polysilicon 1703 -2026 1703 -2026 0 1
rlabel polysilicon 1703 -2032 1703 -2032 0 3
rlabel polysilicon 1710 -2026 1710 -2026 0 1
rlabel polysilicon 1710 -2032 1710 -2032 0 3
rlabel polysilicon 1717 -2026 1717 -2026 0 1
rlabel polysilicon 1717 -2032 1717 -2032 0 3
rlabel polysilicon 1724 -2026 1724 -2026 0 1
rlabel polysilicon 1724 -2032 1724 -2032 0 3
rlabel polysilicon 1731 -2026 1731 -2026 0 1
rlabel polysilicon 1734 -2026 1734 -2026 0 2
rlabel polysilicon 1738 -2026 1738 -2026 0 1
rlabel polysilicon 1738 -2032 1738 -2032 0 3
rlabel polysilicon 1745 -2026 1745 -2026 0 1
rlabel polysilicon 1745 -2032 1745 -2032 0 3
rlabel polysilicon 1752 -2026 1752 -2026 0 1
rlabel polysilicon 1752 -2032 1752 -2032 0 3
rlabel polysilicon 1759 -2026 1759 -2026 0 1
rlabel polysilicon 1759 -2032 1759 -2032 0 3
rlabel polysilicon 1766 -2026 1766 -2026 0 1
rlabel polysilicon 1766 -2032 1766 -2032 0 3
rlabel polysilicon 1773 -2026 1773 -2026 0 1
rlabel polysilicon 1773 -2032 1773 -2032 0 3
rlabel polysilicon 1780 -2026 1780 -2026 0 1
rlabel polysilicon 1780 -2032 1780 -2032 0 3
rlabel polysilicon 1787 -2026 1787 -2026 0 1
rlabel polysilicon 1787 -2032 1787 -2032 0 3
rlabel polysilicon 1794 -2026 1794 -2026 0 1
rlabel polysilicon 1794 -2032 1794 -2032 0 3
rlabel polysilicon 1801 -2026 1801 -2026 0 1
rlabel polysilicon 1801 -2032 1801 -2032 0 3
rlabel polysilicon 1808 -2026 1808 -2026 0 1
rlabel polysilicon 1808 -2032 1808 -2032 0 3
rlabel polysilicon 1815 -2026 1815 -2026 0 1
rlabel polysilicon 1815 -2032 1815 -2032 0 3
rlabel polysilicon 1822 -2026 1822 -2026 0 1
rlabel polysilicon 1822 -2032 1822 -2032 0 3
rlabel polysilicon 1829 -2026 1829 -2026 0 1
rlabel polysilicon 1829 -2032 1829 -2032 0 3
rlabel polysilicon 1836 -2026 1836 -2026 0 1
rlabel polysilicon 1836 -2032 1836 -2032 0 3
rlabel polysilicon 1843 -2026 1843 -2026 0 1
rlabel polysilicon 1843 -2032 1843 -2032 0 3
rlabel polysilicon 1850 -2026 1850 -2026 0 1
rlabel polysilicon 1850 -2032 1850 -2032 0 3
rlabel polysilicon 1857 -2026 1857 -2026 0 1
rlabel polysilicon 1857 -2032 1857 -2032 0 3
rlabel polysilicon 1864 -2026 1864 -2026 0 1
rlabel polysilicon 1864 -2032 1864 -2032 0 3
rlabel polysilicon 1871 -2026 1871 -2026 0 1
rlabel polysilicon 1871 -2032 1871 -2032 0 3
rlabel polysilicon 1878 -2026 1878 -2026 0 1
rlabel polysilicon 1878 -2032 1878 -2032 0 3
rlabel polysilicon 1885 -2026 1885 -2026 0 1
rlabel polysilicon 1885 -2032 1885 -2032 0 3
rlabel polysilicon 1892 -2026 1892 -2026 0 1
rlabel polysilicon 1892 -2032 1892 -2032 0 3
rlabel polysilicon 1899 -2026 1899 -2026 0 1
rlabel polysilicon 1899 -2032 1899 -2032 0 3
rlabel polysilicon 1906 -2026 1906 -2026 0 1
rlabel polysilicon 1906 -2032 1906 -2032 0 3
rlabel polysilicon 1913 -2026 1913 -2026 0 1
rlabel polysilicon 1913 -2032 1913 -2032 0 3
rlabel polysilicon 1920 -2026 1920 -2026 0 1
rlabel polysilicon 1920 -2032 1920 -2032 0 3
rlabel polysilicon 1927 -2026 1927 -2026 0 1
rlabel polysilicon 1927 -2032 1927 -2032 0 3
rlabel polysilicon 1934 -2026 1934 -2026 0 1
rlabel polysilicon 1934 -2032 1934 -2032 0 3
rlabel polysilicon 1941 -2026 1941 -2026 0 1
rlabel polysilicon 1941 -2032 1941 -2032 0 3
rlabel polysilicon 1948 -2026 1948 -2026 0 1
rlabel polysilicon 1948 -2032 1948 -2032 0 3
rlabel polysilicon 1955 -2026 1955 -2026 0 1
rlabel polysilicon 1955 -2032 1955 -2032 0 3
rlabel polysilicon 1962 -2026 1962 -2026 0 1
rlabel polysilicon 1962 -2032 1962 -2032 0 3
rlabel polysilicon 1969 -2026 1969 -2026 0 1
rlabel polysilicon 1969 -2032 1969 -2032 0 3
rlabel polysilicon 1976 -2026 1976 -2026 0 1
rlabel polysilicon 1976 -2032 1976 -2032 0 3
rlabel polysilicon 1983 -2026 1983 -2026 0 1
rlabel polysilicon 1983 -2032 1983 -2032 0 3
rlabel polysilicon 1990 -2026 1990 -2026 0 1
rlabel polysilicon 1990 -2032 1990 -2032 0 3
rlabel polysilicon 1997 -2026 1997 -2026 0 1
rlabel polysilicon 1997 -2032 1997 -2032 0 3
rlabel polysilicon 2004 -2026 2004 -2026 0 1
rlabel polysilicon 2004 -2032 2004 -2032 0 3
rlabel polysilicon 2011 -2026 2011 -2026 0 1
rlabel polysilicon 2011 -2032 2011 -2032 0 3
rlabel polysilicon 2018 -2026 2018 -2026 0 1
rlabel polysilicon 2018 -2032 2018 -2032 0 3
rlabel polysilicon 2025 -2026 2025 -2026 0 1
rlabel polysilicon 2025 -2032 2025 -2032 0 3
rlabel polysilicon 2032 -2026 2032 -2026 0 1
rlabel polysilicon 2032 -2032 2032 -2032 0 3
rlabel polysilicon 2039 -2026 2039 -2026 0 1
rlabel polysilicon 2039 -2032 2039 -2032 0 3
rlabel polysilicon 2046 -2026 2046 -2026 0 1
rlabel polysilicon 2046 -2032 2046 -2032 0 3
rlabel polysilicon 2053 -2026 2053 -2026 0 1
rlabel polysilicon 2053 -2032 2053 -2032 0 3
rlabel polysilicon 2060 -2026 2060 -2026 0 1
rlabel polysilicon 2060 -2032 2060 -2032 0 3
rlabel polysilicon 2067 -2026 2067 -2026 0 1
rlabel polysilicon 2067 -2032 2067 -2032 0 3
rlabel polysilicon 2074 -2026 2074 -2026 0 1
rlabel polysilicon 2074 -2032 2074 -2032 0 3
rlabel polysilicon 2081 -2026 2081 -2026 0 1
rlabel polysilicon 2081 -2032 2081 -2032 0 3
rlabel polysilicon 2088 -2026 2088 -2026 0 1
rlabel polysilicon 2088 -2032 2088 -2032 0 3
rlabel polysilicon 2095 -2026 2095 -2026 0 1
rlabel polysilicon 2095 -2032 2095 -2032 0 3
rlabel polysilicon 2102 -2026 2102 -2026 0 1
rlabel polysilicon 2102 -2032 2102 -2032 0 3
rlabel polysilicon 2109 -2026 2109 -2026 0 1
rlabel polysilicon 2109 -2032 2109 -2032 0 3
rlabel polysilicon 2116 -2026 2116 -2026 0 1
rlabel polysilicon 2116 -2032 2116 -2032 0 3
rlabel polysilicon 2123 -2026 2123 -2026 0 1
rlabel polysilicon 2123 -2032 2123 -2032 0 3
rlabel polysilicon 2130 -2026 2130 -2026 0 1
rlabel polysilicon 2130 -2032 2130 -2032 0 3
rlabel polysilicon 2137 -2026 2137 -2026 0 1
rlabel polysilicon 2137 -2032 2137 -2032 0 3
rlabel polysilicon 2144 -2026 2144 -2026 0 1
rlabel polysilicon 2144 -2032 2144 -2032 0 3
rlabel polysilicon 2151 -2026 2151 -2026 0 1
rlabel polysilicon 2151 -2032 2151 -2032 0 3
rlabel polysilicon 2158 -2026 2158 -2026 0 1
rlabel polysilicon 2158 -2032 2158 -2032 0 3
rlabel polysilicon 2165 -2026 2165 -2026 0 1
rlabel polysilicon 2165 -2032 2165 -2032 0 3
rlabel polysilicon 2172 -2026 2172 -2026 0 1
rlabel polysilicon 2172 -2032 2172 -2032 0 3
rlabel polysilicon 2179 -2026 2179 -2026 0 1
rlabel polysilicon 2179 -2032 2179 -2032 0 3
rlabel polysilicon 2186 -2026 2186 -2026 0 1
rlabel polysilicon 2186 -2032 2186 -2032 0 3
rlabel polysilicon 2193 -2026 2193 -2026 0 1
rlabel polysilicon 2193 -2032 2193 -2032 0 3
rlabel polysilicon 2200 -2026 2200 -2026 0 1
rlabel polysilicon 2200 -2032 2200 -2032 0 3
rlabel polysilicon 2207 -2026 2207 -2026 0 1
rlabel polysilicon 2207 -2032 2207 -2032 0 3
rlabel polysilicon 2214 -2026 2214 -2026 0 1
rlabel polysilicon 2214 -2032 2214 -2032 0 3
rlabel polysilicon 2221 -2026 2221 -2026 0 1
rlabel polysilicon 2221 -2032 2221 -2032 0 3
rlabel polysilicon 2228 -2026 2228 -2026 0 1
rlabel polysilicon 2228 -2032 2228 -2032 0 3
rlabel polysilicon 2235 -2026 2235 -2026 0 1
rlabel polysilicon 2235 -2032 2235 -2032 0 3
rlabel polysilicon 2242 -2026 2242 -2026 0 1
rlabel polysilicon 2242 -2032 2242 -2032 0 3
rlabel polysilicon 2249 -2026 2249 -2026 0 1
rlabel polysilicon 2249 -2032 2249 -2032 0 3
rlabel polysilicon 2256 -2026 2256 -2026 0 1
rlabel polysilicon 2256 -2032 2256 -2032 0 3
rlabel polysilicon 2263 -2026 2263 -2026 0 1
rlabel polysilicon 2263 -2032 2263 -2032 0 3
rlabel polysilicon 2270 -2026 2270 -2026 0 1
rlabel polysilicon 2270 -2032 2270 -2032 0 3
rlabel polysilicon 2277 -2026 2277 -2026 0 1
rlabel polysilicon 2277 -2032 2277 -2032 0 3
rlabel polysilicon 2284 -2026 2284 -2026 0 1
rlabel polysilicon 2284 -2032 2284 -2032 0 3
rlabel polysilicon 2291 -2026 2291 -2026 0 1
rlabel polysilicon 2291 -2032 2291 -2032 0 3
rlabel polysilicon 2298 -2026 2298 -2026 0 1
rlabel polysilicon 2298 -2032 2298 -2032 0 3
rlabel polysilicon 2305 -2026 2305 -2026 0 1
rlabel polysilicon 2305 -2032 2305 -2032 0 3
rlabel polysilicon 2312 -2026 2312 -2026 0 1
rlabel polysilicon 2312 -2032 2312 -2032 0 3
rlabel polysilicon 2319 -2026 2319 -2026 0 1
rlabel polysilicon 2319 -2032 2319 -2032 0 3
rlabel polysilicon 2326 -2026 2326 -2026 0 1
rlabel polysilicon 2326 -2032 2326 -2032 0 3
rlabel polysilicon 2333 -2026 2333 -2026 0 1
rlabel polysilicon 2333 -2032 2333 -2032 0 3
rlabel polysilicon 2340 -2026 2340 -2026 0 1
rlabel polysilicon 2340 -2032 2340 -2032 0 3
rlabel polysilicon 2347 -2026 2347 -2026 0 1
rlabel polysilicon 2347 -2032 2347 -2032 0 3
rlabel polysilicon 2354 -2026 2354 -2026 0 1
rlabel polysilicon 2354 -2032 2354 -2032 0 3
rlabel polysilicon 2361 -2026 2361 -2026 0 1
rlabel polysilicon 2361 -2032 2361 -2032 0 3
rlabel polysilicon 2368 -2026 2368 -2026 0 1
rlabel polysilicon 2368 -2032 2368 -2032 0 3
rlabel polysilicon 2375 -2026 2375 -2026 0 1
rlabel polysilicon 2375 -2032 2375 -2032 0 3
rlabel polysilicon 2382 -2026 2382 -2026 0 1
rlabel polysilicon 2382 -2032 2382 -2032 0 3
rlabel polysilicon 2389 -2026 2389 -2026 0 1
rlabel polysilicon 2389 -2032 2389 -2032 0 3
rlabel polysilicon 2396 -2026 2396 -2026 0 1
rlabel polysilicon 2396 -2032 2396 -2032 0 3
rlabel polysilicon 2403 -2026 2403 -2026 0 1
rlabel polysilicon 2403 -2032 2403 -2032 0 3
rlabel polysilicon 2410 -2026 2410 -2026 0 1
rlabel polysilicon 2410 -2032 2410 -2032 0 3
rlabel polysilicon 2420 -2026 2420 -2026 0 2
rlabel polysilicon 2424 -2026 2424 -2026 0 1
rlabel polysilicon 2424 -2032 2424 -2032 0 3
rlabel polysilicon 9 -2177 9 -2177 0 1
rlabel polysilicon 9 -2183 9 -2183 0 3
rlabel polysilicon 16 -2177 16 -2177 0 1
rlabel polysilicon 16 -2183 16 -2183 0 3
rlabel polysilicon 23 -2177 23 -2177 0 1
rlabel polysilicon 23 -2183 23 -2183 0 3
rlabel polysilicon 30 -2177 30 -2177 0 1
rlabel polysilicon 30 -2183 30 -2183 0 3
rlabel polysilicon 37 -2177 37 -2177 0 1
rlabel polysilicon 40 -2183 40 -2183 0 4
rlabel polysilicon 44 -2177 44 -2177 0 1
rlabel polysilicon 44 -2183 44 -2183 0 3
rlabel polysilicon 51 -2177 51 -2177 0 1
rlabel polysilicon 51 -2183 51 -2183 0 3
rlabel polysilicon 54 -2183 54 -2183 0 4
rlabel polysilicon 58 -2177 58 -2177 0 1
rlabel polysilicon 58 -2183 58 -2183 0 3
rlabel polysilicon 65 -2177 65 -2177 0 1
rlabel polysilicon 65 -2183 65 -2183 0 3
rlabel polysilicon 72 -2177 72 -2177 0 1
rlabel polysilicon 72 -2183 72 -2183 0 3
rlabel polysilicon 79 -2177 79 -2177 0 1
rlabel polysilicon 79 -2183 79 -2183 0 3
rlabel polysilicon 86 -2177 86 -2177 0 1
rlabel polysilicon 86 -2183 86 -2183 0 3
rlabel polysilicon 93 -2177 93 -2177 0 1
rlabel polysilicon 96 -2177 96 -2177 0 2
rlabel polysilicon 93 -2183 93 -2183 0 3
rlabel polysilicon 96 -2183 96 -2183 0 4
rlabel polysilicon 100 -2177 100 -2177 0 1
rlabel polysilicon 100 -2183 100 -2183 0 3
rlabel polysilicon 107 -2177 107 -2177 0 1
rlabel polysilicon 107 -2183 107 -2183 0 3
rlabel polysilicon 114 -2177 114 -2177 0 1
rlabel polysilicon 114 -2183 114 -2183 0 3
rlabel polysilicon 121 -2177 121 -2177 0 1
rlabel polysilicon 124 -2177 124 -2177 0 2
rlabel polysilicon 121 -2183 121 -2183 0 3
rlabel polysilicon 124 -2183 124 -2183 0 4
rlabel polysilicon 131 -2177 131 -2177 0 2
rlabel polysilicon 128 -2183 128 -2183 0 3
rlabel polysilicon 131 -2183 131 -2183 0 4
rlabel polysilicon 135 -2177 135 -2177 0 1
rlabel polysilicon 138 -2177 138 -2177 0 2
rlabel polysilicon 135 -2183 135 -2183 0 3
rlabel polysilicon 138 -2183 138 -2183 0 4
rlabel polysilicon 142 -2177 142 -2177 0 1
rlabel polysilicon 142 -2183 142 -2183 0 3
rlabel polysilicon 149 -2177 149 -2177 0 1
rlabel polysilicon 149 -2183 149 -2183 0 3
rlabel polysilicon 156 -2177 156 -2177 0 1
rlabel polysilicon 156 -2183 156 -2183 0 3
rlabel polysilicon 163 -2177 163 -2177 0 1
rlabel polysilicon 163 -2183 163 -2183 0 3
rlabel polysilicon 170 -2177 170 -2177 0 1
rlabel polysilicon 170 -2183 170 -2183 0 3
rlabel polysilicon 177 -2177 177 -2177 0 1
rlabel polysilicon 177 -2183 177 -2183 0 3
rlabel polysilicon 184 -2177 184 -2177 0 1
rlabel polysilicon 184 -2183 184 -2183 0 3
rlabel polysilicon 191 -2177 191 -2177 0 1
rlabel polysilicon 191 -2183 191 -2183 0 3
rlabel polysilicon 198 -2177 198 -2177 0 1
rlabel polysilicon 198 -2183 198 -2183 0 3
rlabel polysilicon 205 -2177 205 -2177 0 1
rlabel polysilicon 205 -2183 205 -2183 0 3
rlabel polysilicon 212 -2177 212 -2177 0 1
rlabel polysilicon 212 -2183 212 -2183 0 3
rlabel polysilicon 219 -2177 219 -2177 0 1
rlabel polysilicon 219 -2183 219 -2183 0 3
rlabel polysilicon 226 -2177 226 -2177 0 1
rlabel polysilicon 226 -2183 226 -2183 0 3
rlabel polysilicon 233 -2177 233 -2177 0 1
rlabel polysilicon 236 -2177 236 -2177 0 2
rlabel polysilicon 233 -2183 233 -2183 0 3
rlabel polysilicon 236 -2183 236 -2183 0 4
rlabel polysilicon 240 -2177 240 -2177 0 1
rlabel polysilicon 243 -2177 243 -2177 0 2
rlabel polysilicon 247 -2177 247 -2177 0 1
rlabel polysilicon 247 -2183 247 -2183 0 3
rlabel polysilicon 257 -2177 257 -2177 0 2
rlabel polysilicon 257 -2183 257 -2183 0 4
rlabel polysilicon 261 -2177 261 -2177 0 1
rlabel polysilicon 261 -2183 261 -2183 0 3
rlabel polysilicon 268 -2177 268 -2177 0 1
rlabel polysilicon 268 -2183 268 -2183 0 3
rlabel polysilicon 275 -2177 275 -2177 0 1
rlabel polysilicon 275 -2183 275 -2183 0 3
rlabel polysilicon 282 -2177 282 -2177 0 1
rlabel polysilicon 282 -2183 282 -2183 0 3
rlabel polysilicon 289 -2177 289 -2177 0 1
rlabel polysilicon 289 -2183 289 -2183 0 3
rlabel polysilicon 296 -2177 296 -2177 0 1
rlabel polysilicon 296 -2183 296 -2183 0 3
rlabel polysilicon 303 -2177 303 -2177 0 1
rlabel polysilicon 303 -2183 303 -2183 0 3
rlabel polysilicon 310 -2177 310 -2177 0 1
rlabel polysilicon 310 -2183 310 -2183 0 3
rlabel polysilicon 317 -2177 317 -2177 0 1
rlabel polysilicon 317 -2183 317 -2183 0 3
rlabel polysilicon 324 -2177 324 -2177 0 1
rlabel polysilicon 324 -2183 324 -2183 0 3
rlabel polysilicon 331 -2177 331 -2177 0 1
rlabel polysilicon 331 -2183 331 -2183 0 3
rlabel polysilicon 338 -2177 338 -2177 0 1
rlabel polysilicon 338 -2183 338 -2183 0 3
rlabel polysilicon 345 -2177 345 -2177 0 1
rlabel polysilicon 345 -2183 345 -2183 0 3
rlabel polysilicon 352 -2177 352 -2177 0 1
rlabel polysilicon 352 -2183 352 -2183 0 3
rlabel polysilicon 359 -2177 359 -2177 0 1
rlabel polysilicon 359 -2183 359 -2183 0 3
rlabel polysilicon 366 -2177 366 -2177 0 1
rlabel polysilicon 366 -2183 366 -2183 0 3
rlabel polysilicon 373 -2177 373 -2177 0 1
rlabel polysilicon 373 -2183 373 -2183 0 3
rlabel polysilicon 380 -2177 380 -2177 0 1
rlabel polysilicon 380 -2183 380 -2183 0 3
rlabel polysilicon 387 -2177 387 -2177 0 1
rlabel polysilicon 387 -2183 387 -2183 0 3
rlabel polysilicon 394 -2177 394 -2177 0 1
rlabel polysilicon 394 -2183 394 -2183 0 3
rlabel polysilicon 401 -2177 401 -2177 0 1
rlabel polysilicon 404 -2177 404 -2177 0 2
rlabel polysilicon 401 -2183 401 -2183 0 3
rlabel polysilicon 408 -2177 408 -2177 0 1
rlabel polysilicon 408 -2183 408 -2183 0 3
rlabel polysilicon 415 -2177 415 -2177 0 1
rlabel polysilicon 415 -2183 415 -2183 0 3
rlabel polysilicon 422 -2177 422 -2177 0 1
rlabel polysilicon 422 -2183 422 -2183 0 3
rlabel polysilicon 429 -2177 429 -2177 0 1
rlabel polysilicon 429 -2183 429 -2183 0 3
rlabel polysilicon 436 -2177 436 -2177 0 1
rlabel polysilicon 436 -2183 436 -2183 0 3
rlabel polysilicon 443 -2177 443 -2177 0 1
rlabel polysilicon 443 -2183 443 -2183 0 3
rlabel polysilicon 450 -2177 450 -2177 0 1
rlabel polysilicon 450 -2183 450 -2183 0 3
rlabel polysilicon 457 -2177 457 -2177 0 1
rlabel polysilicon 457 -2183 457 -2183 0 3
rlabel polysilicon 464 -2177 464 -2177 0 1
rlabel polysilicon 464 -2183 464 -2183 0 3
rlabel polysilicon 471 -2177 471 -2177 0 1
rlabel polysilicon 471 -2183 471 -2183 0 3
rlabel polysilicon 478 -2177 478 -2177 0 1
rlabel polysilicon 478 -2183 478 -2183 0 3
rlabel polysilicon 485 -2177 485 -2177 0 1
rlabel polysilicon 485 -2183 485 -2183 0 3
rlabel polysilicon 492 -2177 492 -2177 0 1
rlabel polysilicon 492 -2183 492 -2183 0 3
rlabel polysilicon 495 -2183 495 -2183 0 4
rlabel polysilicon 499 -2177 499 -2177 0 1
rlabel polysilicon 499 -2183 499 -2183 0 3
rlabel polysilicon 506 -2177 506 -2177 0 1
rlabel polysilicon 506 -2183 506 -2183 0 3
rlabel polysilicon 513 -2177 513 -2177 0 1
rlabel polysilicon 516 -2177 516 -2177 0 2
rlabel polysilicon 513 -2183 513 -2183 0 3
rlabel polysilicon 516 -2183 516 -2183 0 4
rlabel polysilicon 520 -2177 520 -2177 0 1
rlabel polysilicon 520 -2183 520 -2183 0 3
rlabel polysilicon 527 -2177 527 -2177 0 1
rlabel polysilicon 527 -2183 527 -2183 0 3
rlabel polysilicon 534 -2177 534 -2177 0 1
rlabel polysilicon 534 -2183 534 -2183 0 3
rlabel polysilicon 541 -2177 541 -2177 0 1
rlabel polysilicon 541 -2183 541 -2183 0 3
rlabel polysilicon 548 -2177 548 -2177 0 1
rlabel polysilicon 548 -2183 548 -2183 0 3
rlabel polysilicon 555 -2177 555 -2177 0 1
rlabel polysilicon 555 -2183 555 -2183 0 3
rlabel polysilicon 562 -2177 562 -2177 0 1
rlabel polysilicon 562 -2183 562 -2183 0 3
rlabel polysilicon 569 -2177 569 -2177 0 1
rlabel polysilicon 569 -2183 569 -2183 0 3
rlabel polysilicon 576 -2177 576 -2177 0 1
rlabel polysilicon 576 -2183 576 -2183 0 3
rlabel polysilicon 583 -2177 583 -2177 0 1
rlabel polysilicon 583 -2183 583 -2183 0 3
rlabel polysilicon 590 -2177 590 -2177 0 1
rlabel polysilicon 590 -2183 590 -2183 0 3
rlabel polysilicon 597 -2177 597 -2177 0 1
rlabel polysilicon 597 -2183 597 -2183 0 3
rlabel polysilicon 604 -2177 604 -2177 0 1
rlabel polysilicon 604 -2183 604 -2183 0 3
rlabel polysilicon 611 -2177 611 -2177 0 1
rlabel polysilicon 611 -2183 611 -2183 0 3
rlabel polysilicon 618 -2177 618 -2177 0 1
rlabel polysilicon 618 -2183 618 -2183 0 3
rlabel polysilicon 625 -2177 625 -2177 0 1
rlabel polysilicon 625 -2183 625 -2183 0 3
rlabel polysilicon 632 -2177 632 -2177 0 1
rlabel polysilicon 632 -2183 632 -2183 0 3
rlabel polysilicon 639 -2177 639 -2177 0 1
rlabel polysilicon 639 -2183 639 -2183 0 3
rlabel polysilicon 646 -2177 646 -2177 0 1
rlabel polysilicon 646 -2183 646 -2183 0 3
rlabel polysilicon 653 -2177 653 -2177 0 1
rlabel polysilicon 656 -2177 656 -2177 0 2
rlabel polysilicon 656 -2183 656 -2183 0 4
rlabel polysilicon 660 -2177 660 -2177 0 1
rlabel polysilicon 660 -2183 660 -2183 0 3
rlabel polysilicon 667 -2177 667 -2177 0 1
rlabel polysilicon 670 -2177 670 -2177 0 2
rlabel polysilicon 670 -2183 670 -2183 0 4
rlabel polysilicon 674 -2177 674 -2177 0 1
rlabel polysilicon 674 -2183 674 -2183 0 3
rlabel polysilicon 681 -2177 681 -2177 0 1
rlabel polysilicon 681 -2183 681 -2183 0 3
rlabel polysilicon 688 -2177 688 -2177 0 1
rlabel polysilicon 688 -2183 688 -2183 0 3
rlabel polysilicon 695 -2177 695 -2177 0 1
rlabel polysilicon 695 -2183 695 -2183 0 3
rlabel polysilicon 702 -2177 702 -2177 0 1
rlabel polysilicon 702 -2183 702 -2183 0 3
rlabel polysilicon 709 -2177 709 -2177 0 1
rlabel polysilicon 709 -2183 709 -2183 0 3
rlabel polysilicon 716 -2177 716 -2177 0 1
rlabel polysilicon 716 -2183 716 -2183 0 3
rlabel polysilicon 723 -2177 723 -2177 0 1
rlabel polysilicon 723 -2183 723 -2183 0 3
rlabel polysilicon 730 -2177 730 -2177 0 1
rlabel polysilicon 730 -2183 730 -2183 0 3
rlabel polysilicon 737 -2177 737 -2177 0 1
rlabel polysilicon 737 -2183 737 -2183 0 3
rlabel polysilicon 744 -2177 744 -2177 0 1
rlabel polysilicon 747 -2177 747 -2177 0 2
rlabel polysilicon 744 -2183 744 -2183 0 3
rlabel polysilicon 747 -2183 747 -2183 0 4
rlabel polysilicon 751 -2177 751 -2177 0 1
rlabel polysilicon 751 -2183 751 -2183 0 3
rlabel polysilicon 758 -2177 758 -2177 0 1
rlabel polysilicon 761 -2177 761 -2177 0 2
rlabel polysilicon 758 -2183 758 -2183 0 3
rlabel polysilicon 765 -2177 765 -2177 0 1
rlabel polysilicon 765 -2183 765 -2183 0 3
rlabel polysilicon 772 -2177 772 -2177 0 1
rlabel polysilicon 772 -2183 772 -2183 0 3
rlabel polysilicon 779 -2177 779 -2177 0 1
rlabel polysilicon 779 -2183 779 -2183 0 3
rlabel polysilicon 786 -2177 786 -2177 0 1
rlabel polysilicon 786 -2183 786 -2183 0 3
rlabel polysilicon 789 -2183 789 -2183 0 4
rlabel polysilicon 793 -2177 793 -2177 0 1
rlabel polysilicon 793 -2183 793 -2183 0 3
rlabel polysilicon 800 -2177 800 -2177 0 1
rlabel polysilicon 800 -2183 800 -2183 0 3
rlabel polysilicon 807 -2177 807 -2177 0 1
rlabel polysilicon 807 -2183 807 -2183 0 3
rlabel polysilicon 814 -2177 814 -2177 0 1
rlabel polysilicon 814 -2183 814 -2183 0 3
rlabel polysilicon 821 -2177 821 -2177 0 1
rlabel polysilicon 821 -2183 821 -2183 0 3
rlabel polysilicon 828 -2177 828 -2177 0 1
rlabel polysilicon 828 -2183 828 -2183 0 3
rlabel polysilicon 835 -2177 835 -2177 0 1
rlabel polysilicon 835 -2183 835 -2183 0 3
rlabel polysilicon 842 -2177 842 -2177 0 1
rlabel polysilicon 842 -2183 842 -2183 0 3
rlabel polysilicon 849 -2177 849 -2177 0 1
rlabel polysilicon 849 -2183 849 -2183 0 3
rlabel polysilicon 856 -2177 856 -2177 0 1
rlabel polysilicon 856 -2183 856 -2183 0 3
rlabel polysilicon 863 -2177 863 -2177 0 1
rlabel polysilicon 863 -2183 863 -2183 0 3
rlabel polysilicon 870 -2177 870 -2177 0 1
rlabel polysilicon 870 -2183 870 -2183 0 3
rlabel polysilicon 877 -2177 877 -2177 0 1
rlabel polysilicon 877 -2183 877 -2183 0 3
rlabel polysilicon 884 -2177 884 -2177 0 1
rlabel polysilicon 884 -2183 884 -2183 0 3
rlabel polysilicon 891 -2177 891 -2177 0 1
rlabel polysilicon 891 -2183 891 -2183 0 3
rlabel polysilicon 898 -2177 898 -2177 0 1
rlabel polysilicon 898 -2183 898 -2183 0 3
rlabel polysilicon 905 -2177 905 -2177 0 1
rlabel polysilicon 905 -2183 905 -2183 0 3
rlabel polysilicon 912 -2177 912 -2177 0 1
rlabel polysilicon 912 -2183 912 -2183 0 3
rlabel polysilicon 919 -2177 919 -2177 0 1
rlabel polysilicon 919 -2183 919 -2183 0 3
rlabel polysilicon 926 -2177 926 -2177 0 1
rlabel polysilicon 926 -2183 926 -2183 0 3
rlabel polysilicon 933 -2177 933 -2177 0 1
rlabel polysilicon 933 -2183 933 -2183 0 3
rlabel polysilicon 940 -2177 940 -2177 0 1
rlabel polysilicon 940 -2183 940 -2183 0 3
rlabel polysilicon 947 -2177 947 -2177 0 1
rlabel polysilicon 947 -2183 947 -2183 0 3
rlabel polysilicon 954 -2177 954 -2177 0 1
rlabel polysilicon 954 -2183 954 -2183 0 3
rlabel polysilicon 961 -2177 961 -2177 0 1
rlabel polysilicon 961 -2183 961 -2183 0 3
rlabel polysilicon 968 -2177 968 -2177 0 1
rlabel polysilicon 968 -2183 968 -2183 0 3
rlabel polysilicon 975 -2177 975 -2177 0 1
rlabel polysilicon 978 -2177 978 -2177 0 2
rlabel polysilicon 975 -2183 975 -2183 0 3
rlabel polysilicon 978 -2183 978 -2183 0 4
rlabel polysilicon 982 -2177 982 -2177 0 1
rlabel polysilicon 982 -2183 982 -2183 0 3
rlabel polysilicon 989 -2177 989 -2177 0 1
rlabel polysilicon 989 -2183 989 -2183 0 3
rlabel polysilicon 996 -2177 996 -2177 0 1
rlabel polysilicon 996 -2183 996 -2183 0 3
rlabel polysilicon 1003 -2177 1003 -2177 0 1
rlabel polysilicon 1003 -2183 1003 -2183 0 3
rlabel polysilicon 1010 -2177 1010 -2177 0 1
rlabel polysilicon 1010 -2183 1010 -2183 0 3
rlabel polysilicon 1017 -2177 1017 -2177 0 1
rlabel polysilicon 1017 -2183 1017 -2183 0 3
rlabel polysilicon 1024 -2177 1024 -2177 0 1
rlabel polysilicon 1024 -2183 1024 -2183 0 3
rlabel polysilicon 1031 -2177 1031 -2177 0 1
rlabel polysilicon 1031 -2183 1031 -2183 0 3
rlabel polysilicon 1038 -2177 1038 -2177 0 1
rlabel polysilicon 1038 -2183 1038 -2183 0 3
rlabel polysilicon 1045 -2177 1045 -2177 0 1
rlabel polysilicon 1045 -2183 1045 -2183 0 3
rlabel polysilicon 1052 -2177 1052 -2177 0 1
rlabel polysilicon 1055 -2177 1055 -2177 0 2
rlabel polysilicon 1052 -2183 1052 -2183 0 3
rlabel polysilicon 1055 -2183 1055 -2183 0 4
rlabel polysilicon 1059 -2177 1059 -2177 0 1
rlabel polysilicon 1059 -2183 1059 -2183 0 3
rlabel polysilicon 1066 -2177 1066 -2177 0 1
rlabel polysilicon 1066 -2183 1066 -2183 0 3
rlabel polysilicon 1073 -2177 1073 -2177 0 1
rlabel polysilicon 1073 -2183 1073 -2183 0 3
rlabel polysilicon 1080 -2177 1080 -2177 0 1
rlabel polysilicon 1080 -2183 1080 -2183 0 3
rlabel polysilicon 1087 -2177 1087 -2177 0 1
rlabel polysilicon 1087 -2183 1087 -2183 0 3
rlabel polysilicon 1094 -2177 1094 -2177 0 1
rlabel polysilicon 1094 -2183 1094 -2183 0 3
rlabel polysilicon 1101 -2177 1101 -2177 0 1
rlabel polysilicon 1101 -2183 1101 -2183 0 3
rlabel polysilicon 1108 -2177 1108 -2177 0 1
rlabel polysilicon 1108 -2183 1108 -2183 0 3
rlabel polysilicon 1115 -2177 1115 -2177 0 1
rlabel polysilicon 1115 -2183 1115 -2183 0 3
rlabel polysilicon 1122 -2177 1122 -2177 0 1
rlabel polysilicon 1122 -2183 1122 -2183 0 3
rlabel polysilicon 1129 -2177 1129 -2177 0 1
rlabel polysilicon 1129 -2183 1129 -2183 0 3
rlabel polysilicon 1136 -2177 1136 -2177 0 1
rlabel polysilicon 1136 -2183 1136 -2183 0 3
rlabel polysilicon 1143 -2177 1143 -2177 0 1
rlabel polysilicon 1143 -2183 1143 -2183 0 3
rlabel polysilicon 1150 -2177 1150 -2177 0 1
rlabel polysilicon 1153 -2177 1153 -2177 0 2
rlabel polysilicon 1157 -2177 1157 -2177 0 1
rlabel polysilicon 1157 -2183 1157 -2183 0 3
rlabel polysilicon 1164 -2177 1164 -2177 0 1
rlabel polysilicon 1164 -2183 1164 -2183 0 3
rlabel polysilicon 1171 -2177 1171 -2177 0 1
rlabel polysilicon 1171 -2183 1171 -2183 0 3
rlabel polysilicon 1178 -2177 1178 -2177 0 1
rlabel polysilicon 1178 -2183 1178 -2183 0 3
rlabel polysilicon 1185 -2177 1185 -2177 0 1
rlabel polysilicon 1188 -2177 1188 -2177 0 2
rlabel polysilicon 1185 -2183 1185 -2183 0 3
rlabel polysilicon 1188 -2183 1188 -2183 0 4
rlabel polysilicon 1192 -2177 1192 -2177 0 1
rlabel polysilicon 1192 -2183 1192 -2183 0 3
rlabel polysilicon 1199 -2177 1199 -2177 0 1
rlabel polysilicon 1202 -2177 1202 -2177 0 2
rlabel polysilicon 1199 -2183 1199 -2183 0 3
rlabel polysilicon 1202 -2183 1202 -2183 0 4
rlabel polysilicon 1206 -2177 1206 -2177 0 1
rlabel polysilicon 1206 -2183 1206 -2183 0 3
rlabel polysilicon 1213 -2177 1213 -2177 0 1
rlabel polysilicon 1213 -2183 1213 -2183 0 3
rlabel polysilicon 1220 -2177 1220 -2177 0 1
rlabel polysilicon 1223 -2177 1223 -2177 0 2
rlabel polysilicon 1220 -2183 1220 -2183 0 3
rlabel polysilicon 1223 -2183 1223 -2183 0 4
rlabel polysilicon 1230 -2177 1230 -2177 0 2
rlabel polysilicon 1227 -2183 1227 -2183 0 3
rlabel polysilicon 1230 -2183 1230 -2183 0 4
rlabel polysilicon 1234 -2177 1234 -2177 0 1
rlabel polysilicon 1234 -2183 1234 -2183 0 3
rlabel polysilicon 1241 -2177 1241 -2177 0 1
rlabel polysilicon 1241 -2183 1241 -2183 0 3
rlabel polysilicon 1248 -2177 1248 -2177 0 1
rlabel polysilicon 1248 -2183 1248 -2183 0 3
rlabel polysilicon 1255 -2177 1255 -2177 0 1
rlabel polysilicon 1258 -2177 1258 -2177 0 2
rlabel polysilicon 1255 -2183 1255 -2183 0 3
rlabel polysilicon 1258 -2183 1258 -2183 0 4
rlabel polysilicon 1262 -2177 1262 -2177 0 1
rlabel polysilicon 1262 -2183 1262 -2183 0 3
rlabel polysilicon 1269 -2177 1269 -2177 0 1
rlabel polysilicon 1269 -2183 1269 -2183 0 3
rlabel polysilicon 1276 -2177 1276 -2177 0 1
rlabel polysilicon 1276 -2183 1276 -2183 0 3
rlabel polysilicon 1283 -2177 1283 -2177 0 1
rlabel polysilicon 1283 -2183 1283 -2183 0 3
rlabel polysilicon 1290 -2177 1290 -2177 0 1
rlabel polysilicon 1290 -2183 1290 -2183 0 3
rlabel polysilicon 1297 -2177 1297 -2177 0 1
rlabel polysilicon 1297 -2183 1297 -2183 0 3
rlabel polysilicon 1304 -2177 1304 -2177 0 1
rlabel polysilicon 1307 -2177 1307 -2177 0 2
rlabel polysilicon 1304 -2183 1304 -2183 0 3
rlabel polysilicon 1307 -2183 1307 -2183 0 4
rlabel polysilicon 1311 -2177 1311 -2177 0 1
rlabel polysilicon 1311 -2183 1311 -2183 0 3
rlabel polysilicon 1318 -2177 1318 -2177 0 1
rlabel polysilicon 1318 -2183 1318 -2183 0 3
rlabel polysilicon 1325 -2177 1325 -2177 0 1
rlabel polysilicon 1325 -2183 1325 -2183 0 3
rlabel polysilicon 1332 -2177 1332 -2177 0 1
rlabel polysilicon 1335 -2177 1335 -2177 0 2
rlabel polysilicon 1332 -2183 1332 -2183 0 3
rlabel polysilicon 1335 -2183 1335 -2183 0 4
rlabel polysilicon 1339 -2177 1339 -2177 0 1
rlabel polysilicon 1342 -2177 1342 -2177 0 2
rlabel polysilicon 1339 -2183 1339 -2183 0 3
rlabel polysilicon 1342 -2183 1342 -2183 0 4
rlabel polysilicon 1346 -2177 1346 -2177 0 1
rlabel polysilicon 1346 -2183 1346 -2183 0 3
rlabel polysilicon 1353 -2177 1353 -2177 0 1
rlabel polysilicon 1353 -2183 1353 -2183 0 3
rlabel polysilicon 1360 -2177 1360 -2177 0 1
rlabel polysilicon 1360 -2183 1360 -2183 0 3
rlabel polysilicon 1367 -2177 1367 -2177 0 1
rlabel polysilicon 1367 -2183 1367 -2183 0 3
rlabel polysilicon 1370 -2183 1370 -2183 0 4
rlabel polysilicon 1374 -2177 1374 -2177 0 1
rlabel polysilicon 1374 -2183 1374 -2183 0 3
rlabel polysilicon 1381 -2177 1381 -2177 0 1
rlabel polysilicon 1384 -2177 1384 -2177 0 2
rlabel polysilicon 1381 -2183 1381 -2183 0 3
rlabel polysilicon 1384 -2183 1384 -2183 0 4
rlabel polysilicon 1388 -2177 1388 -2177 0 1
rlabel polysilicon 1388 -2183 1388 -2183 0 3
rlabel polysilicon 1395 -2177 1395 -2177 0 1
rlabel polysilicon 1395 -2183 1395 -2183 0 3
rlabel polysilicon 1402 -2177 1402 -2177 0 1
rlabel polysilicon 1405 -2177 1405 -2177 0 2
rlabel polysilicon 1402 -2183 1402 -2183 0 3
rlabel polysilicon 1405 -2183 1405 -2183 0 4
rlabel polysilicon 1409 -2177 1409 -2177 0 1
rlabel polysilicon 1409 -2183 1409 -2183 0 3
rlabel polysilicon 1416 -2177 1416 -2177 0 1
rlabel polysilicon 1416 -2183 1416 -2183 0 3
rlabel polysilicon 1423 -2177 1423 -2177 0 1
rlabel polysilicon 1423 -2183 1423 -2183 0 3
rlabel polysilicon 1430 -2177 1430 -2177 0 1
rlabel polysilicon 1430 -2183 1430 -2183 0 3
rlabel polysilicon 1437 -2177 1437 -2177 0 1
rlabel polysilicon 1437 -2183 1437 -2183 0 3
rlabel polysilicon 1444 -2177 1444 -2177 0 1
rlabel polysilicon 1444 -2183 1444 -2183 0 3
rlabel polysilicon 1451 -2177 1451 -2177 0 1
rlabel polysilicon 1451 -2183 1451 -2183 0 3
rlabel polysilicon 1458 -2177 1458 -2177 0 1
rlabel polysilicon 1458 -2183 1458 -2183 0 3
rlabel polysilicon 1465 -2177 1465 -2177 0 1
rlabel polysilicon 1465 -2183 1465 -2183 0 3
rlabel polysilicon 1472 -2177 1472 -2177 0 1
rlabel polysilicon 1472 -2183 1472 -2183 0 3
rlabel polysilicon 1479 -2177 1479 -2177 0 1
rlabel polysilicon 1479 -2183 1479 -2183 0 3
rlabel polysilicon 1486 -2177 1486 -2177 0 1
rlabel polysilicon 1489 -2177 1489 -2177 0 2
rlabel polysilicon 1486 -2183 1486 -2183 0 3
rlabel polysilicon 1489 -2183 1489 -2183 0 4
rlabel polysilicon 1493 -2177 1493 -2177 0 1
rlabel polysilicon 1493 -2183 1493 -2183 0 3
rlabel polysilicon 1500 -2177 1500 -2177 0 1
rlabel polysilicon 1500 -2183 1500 -2183 0 3
rlabel polysilicon 1507 -2177 1507 -2177 0 1
rlabel polysilicon 1507 -2183 1507 -2183 0 3
rlabel polysilicon 1514 -2177 1514 -2177 0 1
rlabel polysilicon 1514 -2183 1514 -2183 0 3
rlabel polysilicon 1521 -2177 1521 -2177 0 1
rlabel polysilicon 1521 -2183 1521 -2183 0 3
rlabel polysilicon 1528 -2177 1528 -2177 0 1
rlabel polysilicon 1528 -2183 1528 -2183 0 3
rlabel polysilicon 1535 -2177 1535 -2177 0 1
rlabel polysilicon 1535 -2183 1535 -2183 0 3
rlabel polysilicon 1542 -2177 1542 -2177 0 1
rlabel polysilicon 1542 -2183 1542 -2183 0 3
rlabel polysilicon 1549 -2177 1549 -2177 0 1
rlabel polysilicon 1549 -2183 1549 -2183 0 3
rlabel polysilicon 1556 -2177 1556 -2177 0 1
rlabel polysilicon 1556 -2183 1556 -2183 0 3
rlabel polysilicon 1563 -2177 1563 -2177 0 1
rlabel polysilicon 1563 -2183 1563 -2183 0 3
rlabel polysilicon 1570 -2177 1570 -2177 0 1
rlabel polysilicon 1570 -2183 1570 -2183 0 3
rlabel polysilicon 1577 -2177 1577 -2177 0 1
rlabel polysilicon 1580 -2177 1580 -2177 0 2
rlabel polysilicon 1580 -2183 1580 -2183 0 4
rlabel polysilicon 1584 -2177 1584 -2177 0 1
rlabel polysilicon 1584 -2183 1584 -2183 0 3
rlabel polysilicon 1591 -2177 1591 -2177 0 1
rlabel polysilicon 1591 -2183 1591 -2183 0 3
rlabel polysilicon 1598 -2177 1598 -2177 0 1
rlabel polysilicon 1598 -2183 1598 -2183 0 3
rlabel polysilicon 1605 -2177 1605 -2177 0 1
rlabel polysilicon 1605 -2183 1605 -2183 0 3
rlabel polysilicon 1612 -2177 1612 -2177 0 1
rlabel polysilicon 1612 -2183 1612 -2183 0 3
rlabel polysilicon 1619 -2177 1619 -2177 0 1
rlabel polysilicon 1619 -2183 1619 -2183 0 3
rlabel polysilicon 1626 -2177 1626 -2177 0 1
rlabel polysilicon 1626 -2183 1626 -2183 0 3
rlabel polysilicon 1633 -2177 1633 -2177 0 1
rlabel polysilicon 1633 -2183 1633 -2183 0 3
rlabel polysilicon 1640 -2177 1640 -2177 0 1
rlabel polysilicon 1640 -2183 1640 -2183 0 3
rlabel polysilicon 1647 -2177 1647 -2177 0 1
rlabel polysilicon 1650 -2177 1650 -2177 0 2
rlabel polysilicon 1647 -2183 1647 -2183 0 3
rlabel polysilicon 1650 -2183 1650 -2183 0 4
rlabel polysilicon 1654 -2177 1654 -2177 0 1
rlabel polysilicon 1654 -2183 1654 -2183 0 3
rlabel polysilicon 1661 -2177 1661 -2177 0 1
rlabel polysilicon 1661 -2183 1661 -2183 0 3
rlabel polysilicon 1668 -2177 1668 -2177 0 1
rlabel polysilicon 1668 -2183 1668 -2183 0 3
rlabel polysilicon 1675 -2177 1675 -2177 0 1
rlabel polysilicon 1675 -2183 1675 -2183 0 3
rlabel polysilicon 1682 -2177 1682 -2177 0 1
rlabel polysilicon 1682 -2183 1682 -2183 0 3
rlabel polysilicon 1689 -2177 1689 -2177 0 1
rlabel polysilicon 1689 -2183 1689 -2183 0 3
rlabel polysilicon 1696 -2177 1696 -2177 0 1
rlabel polysilicon 1696 -2183 1696 -2183 0 3
rlabel polysilicon 1703 -2177 1703 -2177 0 1
rlabel polysilicon 1703 -2183 1703 -2183 0 3
rlabel polysilicon 1713 -2177 1713 -2177 0 2
rlabel polysilicon 1717 -2177 1717 -2177 0 1
rlabel polysilicon 1717 -2183 1717 -2183 0 3
rlabel polysilicon 1724 -2177 1724 -2177 0 1
rlabel polysilicon 1724 -2183 1724 -2183 0 3
rlabel polysilicon 1731 -2177 1731 -2177 0 1
rlabel polysilicon 1731 -2183 1731 -2183 0 3
rlabel polysilicon 1738 -2177 1738 -2177 0 1
rlabel polysilicon 1738 -2183 1738 -2183 0 3
rlabel polysilicon 1745 -2177 1745 -2177 0 1
rlabel polysilicon 1745 -2183 1745 -2183 0 3
rlabel polysilicon 1752 -2177 1752 -2177 0 1
rlabel polysilicon 1752 -2183 1752 -2183 0 3
rlabel polysilicon 1759 -2177 1759 -2177 0 1
rlabel polysilicon 1759 -2183 1759 -2183 0 3
rlabel polysilicon 1766 -2177 1766 -2177 0 1
rlabel polysilicon 1766 -2183 1766 -2183 0 3
rlabel polysilicon 1773 -2177 1773 -2177 0 1
rlabel polysilicon 1773 -2183 1773 -2183 0 3
rlabel polysilicon 1780 -2177 1780 -2177 0 1
rlabel polysilicon 1780 -2183 1780 -2183 0 3
rlabel polysilicon 1787 -2177 1787 -2177 0 1
rlabel polysilicon 1787 -2183 1787 -2183 0 3
rlabel polysilicon 1794 -2177 1794 -2177 0 1
rlabel polysilicon 1794 -2183 1794 -2183 0 3
rlabel polysilicon 1801 -2177 1801 -2177 0 1
rlabel polysilicon 1801 -2183 1801 -2183 0 3
rlabel polysilicon 1808 -2177 1808 -2177 0 1
rlabel polysilicon 1808 -2183 1808 -2183 0 3
rlabel polysilicon 1815 -2177 1815 -2177 0 1
rlabel polysilicon 1815 -2183 1815 -2183 0 3
rlabel polysilicon 1822 -2177 1822 -2177 0 1
rlabel polysilicon 1822 -2183 1822 -2183 0 3
rlabel polysilicon 1829 -2177 1829 -2177 0 1
rlabel polysilicon 1829 -2183 1829 -2183 0 3
rlabel polysilicon 1836 -2177 1836 -2177 0 1
rlabel polysilicon 1843 -2177 1843 -2177 0 1
rlabel polysilicon 1843 -2183 1843 -2183 0 3
rlabel polysilicon 1850 -2177 1850 -2177 0 1
rlabel polysilicon 1850 -2183 1850 -2183 0 3
rlabel polysilicon 1857 -2177 1857 -2177 0 1
rlabel polysilicon 1857 -2183 1857 -2183 0 3
rlabel polysilicon 1860 -2183 1860 -2183 0 4
rlabel polysilicon 1864 -2177 1864 -2177 0 1
rlabel polysilicon 1864 -2183 1864 -2183 0 3
rlabel polysilicon 1871 -2177 1871 -2177 0 1
rlabel polysilicon 1871 -2183 1871 -2183 0 3
rlabel polysilicon 1878 -2177 1878 -2177 0 1
rlabel polysilicon 1878 -2183 1878 -2183 0 3
rlabel polysilicon 1885 -2177 1885 -2177 0 1
rlabel polysilicon 1885 -2183 1885 -2183 0 3
rlabel polysilicon 1892 -2177 1892 -2177 0 1
rlabel polysilicon 1892 -2183 1892 -2183 0 3
rlabel polysilicon 1899 -2177 1899 -2177 0 1
rlabel polysilicon 1899 -2183 1899 -2183 0 3
rlabel polysilicon 1906 -2177 1906 -2177 0 1
rlabel polysilicon 1906 -2183 1906 -2183 0 3
rlabel polysilicon 1913 -2177 1913 -2177 0 1
rlabel polysilicon 1913 -2183 1913 -2183 0 3
rlabel polysilicon 1920 -2177 1920 -2177 0 1
rlabel polysilicon 1920 -2183 1920 -2183 0 3
rlabel polysilicon 1927 -2177 1927 -2177 0 1
rlabel polysilicon 1927 -2183 1927 -2183 0 3
rlabel polysilicon 1934 -2177 1934 -2177 0 1
rlabel polysilicon 1934 -2183 1934 -2183 0 3
rlabel polysilicon 1941 -2177 1941 -2177 0 1
rlabel polysilicon 1941 -2183 1941 -2183 0 3
rlabel polysilicon 1948 -2177 1948 -2177 0 1
rlabel polysilicon 1948 -2183 1948 -2183 0 3
rlabel polysilicon 1955 -2177 1955 -2177 0 1
rlabel polysilicon 1955 -2183 1955 -2183 0 3
rlabel polysilicon 1962 -2177 1962 -2177 0 1
rlabel polysilicon 1962 -2183 1962 -2183 0 3
rlabel polysilicon 1969 -2177 1969 -2177 0 1
rlabel polysilicon 1969 -2183 1969 -2183 0 3
rlabel polysilicon 1976 -2177 1976 -2177 0 1
rlabel polysilicon 1976 -2183 1976 -2183 0 3
rlabel polysilicon 1983 -2177 1983 -2177 0 1
rlabel polysilicon 1983 -2183 1983 -2183 0 3
rlabel polysilicon 1990 -2177 1990 -2177 0 1
rlabel polysilicon 1990 -2183 1990 -2183 0 3
rlabel polysilicon 1997 -2177 1997 -2177 0 1
rlabel polysilicon 1997 -2183 1997 -2183 0 3
rlabel polysilicon 2004 -2177 2004 -2177 0 1
rlabel polysilicon 2004 -2183 2004 -2183 0 3
rlabel polysilicon 2011 -2177 2011 -2177 0 1
rlabel polysilicon 2011 -2183 2011 -2183 0 3
rlabel polysilicon 2018 -2177 2018 -2177 0 1
rlabel polysilicon 2018 -2183 2018 -2183 0 3
rlabel polysilicon 2025 -2177 2025 -2177 0 1
rlabel polysilicon 2025 -2183 2025 -2183 0 3
rlabel polysilicon 2032 -2177 2032 -2177 0 1
rlabel polysilicon 2032 -2183 2032 -2183 0 3
rlabel polysilicon 2039 -2177 2039 -2177 0 1
rlabel polysilicon 2039 -2183 2039 -2183 0 3
rlabel polysilicon 2046 -2177 2046 -2177 0 1
rlabel polysilicon 2046 -2183 2046 -2183 0 3
rlabel polysilicon 2053 -2177 2053 -2177 0 1
rlabel polysilicon 2053 -2183 2053 -2183 0 3
rlabel polysilicon 2060 -2177 2060 -2177 0 1
rlabel polysilicon 2060 -2183 2060 -2183 0 3
rlabel polysilicon 2067 -2177 2067 -2177 0 1
rlabel polysilicon 2067 -2183 2067 -2183 0 3
rlabel polysilicon 2074 -2177 2074 -2177 0 1
rlabel polysilicon 2074 -2183 2074 -2183 0 3
rlabel polysilicon 2081 -2177 2081 -2177 0 1
rlabel polysilicon 2081 -2183 2081 -2183 0 3
rlabel polysilicon 2088 -2177 2088 -2177 0 1
rlabel polysilicon 2088 -2183 2088 -2183 0 3
rlabel polysilicon 2095 -2177 2095 -2177 0 1
rlabel polysilicon 2095 -2183 2095 -2183 0 3
rlabel polysilicon 2102 -2177 2102 -2177 0 1
rlabel polysilicon 2102 -2183 2102 -2183 0 3
rlabel polysilicon 2109 -2177 2109 -2177 0 1
rlabel polysilicon 2109 -2183 2109 -2183 0 3
rlabel polysilicon 2116 -2177 2116 -2177 0 1
rlabel polysilicon 2116 -2183 2116 -2183 0 3
rlabel polysilicon 2123 -2177 2123 -2177 0 1
rlabel polysilicon 2123 -2183 2123 -2183 0 3
rlabel polysilicon 2130 -2177 2130 -2177 0 1
rlabel polysilicon 2130 -2183 2130 -2183 0 3
rlabel polysilicon 2137 -2177 2137 -2177 0 1
rlabel polysilicon 2137 -2183 2137 -2183 0 3
rlabel polysilicon 2144 -2177 2144 -2177 0 1
rlabel polysilicon 2144 -2183 2144 -2183 0 3
rlabel polysilicon 2151 -2177 2151 -2177 0 1
rlabel polysilicon 2151 -2183 2151 -2183 0 3
rlabel polysilicon 2158 -2177 2158 -2177 0 1
rlabel polysilicon 2158 -2183 2158 -2183 0 3
rlabel polysilicon 2165 -2177 2165 -2177 0 1
rlabel polysilicon 2165 -2183 2165 -2183 0 3
rlabel polysilicon 2172 -2177 2172 -2177 0 1
rlabel polysilicon 2172 -2183 2172 -2183 0 3
rlabel polysilicon 2179 -2177 2179 -2177 0 1
rlabel polysilicon 2179 -2183 2179 -2183 0 3
rlabel polysilicon 2186 -2177 2186 -2177 0 1
rlabel polysilicon 2186 -2183 2186 -2183 0 3
rlabel polysilicon 2193 -2177 2193 -2177 0 1
rlabel polysilicon 2193 -2183 2193 -2183 0 3
rlabel polysilicon 2200 -2177 2200 -2177 0 1
rlabel polysilicon 2200 -2183 2200 -2183 0 3
rlabel polysilicon 2207 -2177 2207 -2177 0 1
rlabel polysilicon 2207 -2183 2207 -2183 0 3
rlabel polysilicon 2214 -2177 2214 -2177 0 1
rlabel polysilicon 2214 -2183 2214 -2183 0 3
rlabel polysilicon 2221 -2177 2221 -2177 0 1
rlabel polysilicon 2221 -2183 2221 -2183 0 3
rlabel polysilicon 2228 -2177 2228 -2177 0 1
rlabel polysilicon 2228 -2183 2228 -2183 0 3
rlabel polysilicon 2235 -2177 2235 -2177 0 1
rlabel polysilicon 2235 -2183 2235 -2183 0 3
rlabel polysilicon 2242 -2177 2242 -2177 0 1
rlabel polysilicon 2242 -2183 2242 -2183 0 3
rlabel polysilicon 2249 -2177 2249 -2177 0 1
rlabel polysilicon 2249 -2183 2249 -2183 0 3
rlabel polysilicon 2256 -2177 2256 -2177 0 1
rlabel polysilicon 2256 -2183 2256 -2183 0 3
rlabel polysilicon 2263 -2177 2263 -2177 0 1
rlabel polysilicon 2263 -2183 2263 -2183 0 3
rlabel polysilicon 2270 -2177 2270 -2177 0 1
rlabel polysilicon 2270 -2183 2270 -2183 0 3
rlabel polysilicon 2277 -2177 2277 -2177 0 1
rlabel polysilicon 2277 -2183 2277 -2183 0 3
rlabel polysilicon 2284 -2177 2284 -2177 0 1
rlabel polysilicon 2284 -2183 2284 -2183 0 3
rlabel polysilicon 2291 -2177 2291 -2177 0 1
rlabel polysilicon 2291 -2183 2291 -2183 0 3
rlabel polysilicon 2298 -2177 2298 -2177 0 1
rlabel polysilicon 2298 -2183 2298 -2183 0 3
rlabel polysilicon 2305 -2177 2305 -2177 0 1
rlabel polysilicon 2305 -2183 2305 -2183 0 3
rlabel polysilicon 2312 -2177 2312 -2177 0 1
rlabel polysilicon 2312 -2183 2312 -2183 0 3
rlabel polysilicon 2319 -2177 2319 -2177 0 1
rlabel polysilicon 2319 -2183 2319 -2183 0 3
rlabel polysilicon 2326 -2177 2326 -2177 0 1
rlabel polysilicon 2326 -2183 2326 -2183 0 3
rlabel polysilicon 2333 -2177 2333 -2177 0 1
rlabel polysilicon 2333 -2183 2333 -2183 0 3
rlabel polysilicon 2340 -2177 2340 -2177 0 1
rlabel polysilicon 2340 -2183 2340 -2183 0 3
rlabel polysilicon 2347 -2177 2347 -2177 0 1
rlabel polysilicon 2347 -2183 2347 -2183 0 3
rlabel polysilicon 2354 -2177 2354 -2177 0 1
rlabel polysilicon 2354 -2183 2354 -2183 0 3
rlabel polysilicon 2361 -2177 2361 -2177 0 1
rlabel polysilicon 2361 -2183 2361 -2183 0 3
rlabel polysilicon 2368 -2177 2368 -2177 0 1
rlabel polysilicon 2368 -2183 2368 -2183 0 3
rlabel polysilicon 2375 -2177 2375 -2177 0 1
rlabel polysilicon 2375 -2183 2375 -2183 0 3
rlabel polysilicon 2382 -2177 2382 -2177 0 1
rlabel polysilicon 2382 -2183 2382 -2183 0 3
rlabel polysilicon 2389 -2177 2389 -2177 0 1
rlabel polysilicon 2389 -2183 2389 -2183 0 3
rlabel polysilicon 2396 -2177 2396 -2177 0 1
rlabel polysilicon 2396 -2183 2396 -2183 0 3
rlabel polysilicon 2403 -2177 2403 -2177 0 1
rlabel polysilicon 2403 -2183 2403 -2183 0 3
rlabel polysilicon 2410 -2177 2410 -2177 0 1
rlabel polysilicon 2410 -2183 2410 -2183 0 3
rlabel polysilicon 2417 -2177 2417 -2177 0 1
rlabel polysilicon 2417 -2183 2417 -2183 0 3
rlabel polysilicon 2424 -2177 2424 -2177 0 1
rlabel polysilicon 2424 -2183 2424 -2183 0 3
rlabel polysilicon 2 -2326 2 -2326 0 1
rlabel polysilicon 2 -2332 2 -2332 0 3
rlabel polysilicon 16 -2326 16 -2326 0 1
rlabel polysilicon 16 -2332 16 -2332 0 3
rlabel polysilicon 23 -2326 23 -2326 0 1
rlabel polysilicon 23 -2332 23 -2332 0 3
rlabel polysilicon 33 -2326 33 -2326 0 2
rlabel polysilicon 30 -2332 30 -2332 0 3
rlabel polysilicon 33 -2332 33 -2332 0 4
rlabel polysilicon 37 -2326 37 -2326 0 1
rlabel polysilicon 37 -2332 37 -2332 0 3
rlabel polysilicon 44 -2326 44 -2326 0 1
rlabel polysilicon 44 -2332 44 -2332 0 3
rlabel polysilicon 51 -2326 51 -2326 0 1
rlabel polysilicon 51 -2332 51 -2332 0 3
rlabel polysilicon 58 -2326 58 -2326 0 1
rlabel polysilicon 58 -2332 58 -2332 0 3
rlabel polysilicon 65 -2326 65 -2326 0 1
rlabel polysilicon 65 -2332 65 -2332 0 3
rlabel polysilicon 72 -2326 72 -2326 0 1
rlabel polysilicon 72 -2332 72 -2332 0 3
rlabel polysilicon 79 -2326 79 -2326 0 1
rlabel polysilicon 79 -2332 79 -2332 0 3
rlabel polysilicon 86 -2326 86 -2326 0 1
rlabel polysilicon 86 -2332 86 -2332 0 3
rlabel polysilicon 93 -2326 93 -2326 0 1
rlabel polysilicon 93 -2332 93 -2332 0 3
rlabel polysilicon 96 -2332 96 -2332 0 4
rlabel polysilicon 100 -2326 100 -2326 0 1
rlabel polysilicon 100 -2332 100 -2332 0 3
rlabel polysilicon 107 -2326 107 -2326 0 1
rlabel polysilicon 107 -2332 107 -2332 0 3
rlabel polysilicon 114 -2326 114 -2326 0 1
rlabel polysilicon 114 -2332 114 -2332 0 3
rlabel polysilicon 121 -2326 121 -2326 0 1
rlabel polysilicon 121 -2332 121 -2332 0 3
rlabel polysilicon 128 -2326 128 -2326 0 1
rlabel polysilicon 128 -2332 128 -2332 0 3
rlabel polysilicon 135 -2326 135 -2326 0 1
rlabel polysilicon 135 -2332 135 -2332 0 3
rlabel polysilicon 142 -2326 142 -2326 0 1
rlabel polysilicon 145 -2326 145 -2326 0 2
rlabel polysilicon 142 -2332 142 -2332 0 3
rlabel polysilicon 145 -2332 145 -2332 0 4
rlabel polysilicon 149 -2326 149 -2326 0 1
rlabel polysilicon 149 -2332 149 -2332 0 3
rlabel polysilicon 156 -2326 156 -2326 0 1
rlabel polysilicon 156 -2332 156 -2332 0 3
rlabel polysilicon 163 -2326 163 -2326 0 1
rlabel polysilicon 166 -2326 166 -2326 0 2
rlabel polysilicon 163 -2332 163 -2332 0 3
rlabel polysilicon 166 -2332 166 -2332 0 4
rlabel polysilicon 170 -2326 170 -2326 0 1
rlabel polysilicon 170 -2332 170 -2332 0 3
rlabel polysilicon 177 -2326 177 -2326 0 1
rlabel polysilicon 184 -2326 184 -2326 0 1
rlabel polysilicon 184 -2332 184 -2332 0 3
rlabel polysilicon 191 -2326 191 -2326 0 1
rlabel polysilicon 191 -2332 191 -2332 0 3
rlabel polysilicon 198 -2326 198 -2326 0 1
rlabel polysilicon 198 -2332 198 -2332 0 3
rlabel polysilicon 205 -2326 205 -2326 0 1
rlabel polysilicon 205 -2332 205 -2332 0 3
rlabel polysilicon 212 -2326 212 -2326 0 1
rlabel polysilicon 212 -2332 212 -2332 0 3
rlabel polysilicon 219 -2326 219 -2326 0 1
rlabel polysilicon 219 -2332 219 -2332 0 3
rlabel polysilicon 226 -2326 226 -2326 0 1
rlabel polysilicon 226 -2332 226 -2332 0 3
rlabel polysilicon 233 -2326 233 -2326 0 1
rlabel polysilicon 233 -2332 233 -2332 0 3
rlabel polysilicon 243 -2326 243 -2326 0 2
rlabel polysilicon 243 -2332 243 -2332 0 4
rlabel polysilicon 247 -2326 247 -2326 0 1
rlabel polysilicon 250 -2326 250 -2326 0 2
rlabel polysilicon 247 -2332 247 -2332 0 3
rlabel polysilicon 254 -2326 254 -2326 0 1
rlabel polysilicon 254 -2332 254 -2332 0 3
rlabel polysilicon 261 -2326 261 -2326 0 1
rlabel polysilicon 261 -2332 261 -2332 0 3
rlabel polysilicon 268 -2326 268 -2326 0 1
rlabel polysilicon 268 -2332 268 -2332 0 3
rlabel polysilicon 275 -2326 275 -2326 0 1
rlabel polysilicon 275 -2332 275 -2332 0 3
rlabel polysilicon 282 -2326 282 -2326 0 1
rlabel polysilicon 282 -2332 282 -2332 0 3
rlabel polysilicon 289 -2326 289 -2326 0 1
rlabel polysilicon 289 -2332 289 -2332 0 3
rlabel polysilicon 296 -2326 296 -2326 0 1
rlabel polysilicon 296 -2332 296 -2332 0 3
rlabel polysilicon 303 -2326 303 -2326 0 1
rlabel polysilicon 303 -2332 303 -2332 0 3
rlabel polysilicon 310 -2326 310 -2326 0 1
rlabel polysilicon 310 -2332 310 -2332 0 3
rlabel polysilicon 317 -2326 317 -2326 0 1
rlabel polysilicon 317 -2332 317 -2332 0 3
rlabel polysilicon 324 -2326 324 -2326 0 1
rlabel polysilicon 324 -2332 324 -2332 0 3
rlabel polysilicon 331 -2326 331 -2326 0 1
rlabel polysilicon 331 -2332 331 -2332 0 3
rlabel polysilicon 338 -2326 338 -2326 0 1
rlabel polysilicon 338 -2332 338 -2332 0 3
rlabel polysilicon 345 -2326 345 -2326 0 1
rlabel polysilicon 345 -2332 345 -2332 0 3
rlabel polysilicon 352 -2326 352 -2326 0 1
rlabel polysilicon 352 -2332 352 -2332 0 3
rlabel polysilicon 359 -2326 359 -2326 0 1
rlabel polysilicon 359 -2332 359 -2332 0 3
rlabel polysilicon 366 -2326 366 -2326 0 1
rlabel polysilicon 366 -2332 366 -2332 0 3
rlabel polysilicon 373 -2326 373 -2326 0 1
rlabel polysilicon 373 -2332 373 -2332 0 3
rlabel polysilicon 380 -2326 380 -2326 0 1
rlabel polysilicon 380 -2332 380 -2332 0 3
rlabel polysilicon 387 -2326 387 -2326 0 1
rlabel polysilicon 387 -2332 387 -2332 0 3
rlabel polysilicon 394 -2326 394 -2326 0 1
rlabel polysilicon 394 -2332 394 -2332 0 3
rlabel polysilicon 401 -2326 401 -2326 0 1
rlabel polysilicon 401 -2332 401 -2332 0 3
rlabel polysilicon 408 -2326 408 -2326 0 1
rlabel polysilicon 408 -2332 408 -2332 0 3
rlabel polysilicon 415 -2326 415 -2326 0 1
rlabel polysilicon 415 -2332 415 -2332 0 3
rlabel polysilicon 422 -2326 422 -2326 0 1
rlabel polysilicon 422 -2332 422 -2332 0 3
rlabel polysilicon 429 -2326 429 -2326 0 1
rlabel polysilicon 436 -2326 436 -2326 0 1
rlabel polysilicon 436 -2332 436 -2332 0 3
rlabel polysilicon 443 -2326 443 -2326 0 1
rlabel polysilicon 443 -2332 443 -2332 0 3
rlabel polysilicon 450 -2326 450 -2326 0 1
rlabel polysilicon 450 -2332 450 -2332 0 3
rlabel polysilicon 457 -2326 457 -2326 0 1
rlabel polysilicon 457 -2332 457 -2332 0 3
rlabel polysilicon 464 -2326 464 -2326 0 1
rlabel polysilicon 464 -2332 464 -2332 0 3
rlabel polysilicon 471 -2326 471 -2326 0 1
rlabel polysilicon 471 -2332 471 -2332 0 3
rlabel polysilicon 478 -2326 478 -2326 0 1
rlabel polysilicon 478 -2332 478 -2332 0 3
rlabel polysilicon 485 -2326 485 -2326 0 1
rlabel polysilicon 485 -2332 485 -2332 0 3
rlabel polysilicon 492 -2326 492 -2326 0 1
rlabel polysilicon 492 -2332 492 -2332 0 3
rlabel polysilicon 499 -2326 499 -2326 0 1
rlabel polysilicon 499 -2332 499 -2332 0 3
rlabel polysilicon 506 -2326 506 -2326 0 1
rlabel polysilicon 506 -2332 506 -2332 0 3
rlabel polysilicon 513 -2326 513 -2326 0 1
rlabel polysilicon 513 -2332 513 -2332 0 3
rlabel polysilicon 520 -2326 520 -2326 0 1
rlabel polysilicon 520 -2332 520 -2332 0 3
rlabel polysilicon 527 -2326 527 -2326 0 1
rlabel polysilicon 527 -2332 527 -2332 0 3
rlabel polysilicon 534 -2326 534 -2326 0 1
rlabel polysilicon 534 -2332 534 -2332 0 3
rlabel polysilicon 541 -2326 541 -2326 0 1
rlabel polysilicon 541 -2332 541 -2332 0 3
rlabel polysilicon 548 -2326 548 -2326 0 1
rlabel polysilicon 548 -2332 548 -2332 0 3
rlabel polysilicon 555 -2326 555 -2326 0 1
rlabel polysilicon 555 -2332 555 -2332 0 3
rlabel polysilicon 562 -2326 562 -2326 0 1
rlabel polysilicon 562 -2332 562 -2332 0 3
rlabel polysilicon 569 -2326 569 -2326 0 1
rlabel polysilicon 569 -2332 569 -2332 0 3
rlabel polysilicon 576 -2326 576 -2326 0 1
rlabel polysilicon 576 -2332 576 -2332 0 3
rlabel polysilicon 583 -2326 583 -2326 0 1
rlabel polysilicon 583 -2332 583 -2332 0 3
rlabel polysilicon 590 -2326 590 -2326 0 1
rlabel polysilicon 593 -2326 593 -2326 0 2
rlabel polysilicon 593 -2332 593 -2332 0 4
rlabel polysilicon 597 -2326 597 -2326 0 1
rlabel polysilicon 597 -2332 597 -2332 0 3
rlabel polysilicon 604 -2326 604 -2326 0 1
rlabel polysilicon 604 -2332 604 -2332 0 3
rlabel polysilicon 611 -2326 611 -2326 0 1
rlabel polysilicon 611 -2332 611 -2332 0 3
rlabel polysilicon 618 -2326 618 -2326 0 1
rlabel polysilicon 621 -2326 621 -2326 0 2
rlabel polysilicon 618 -2332 618 -2332 0 3
rlabel polysilicon 621 -2332 621 -2332 0 4
rlabel polysilicon 625 -2326 625 -2326 0 1
rlabel polysilicon 628 -2332 628 -2332 0 4
rlabel polysilicon 632 -2326 632 -2326 0 1
rlabel polysilicon 632 -2332 632 -2332 0 3
rlabel polysilicon 639 -2326 639 -2326 0 1
rlabel polysilicon 639 -2332 639 -2332 0 3
rlabel polysilicon 646 -2326 646 -2326 0 1
rlabel polysilicon 646 -2332 646 -2332 0 3
rlabel polysilicon 653 -2326 653 -2326 0 1
rlabel polysilicon 653 -2332 653 -2332 0 3
rlabel polysilicon 660 -2326 660 -2326 0 1
rlabel polysilicon 663 -2326 663 -2326 0 2
rlabel polysilicon 660 -2332 660 -2332 0 3
rlabel polysilicon 667 -2326 667 -2326 0 1
rlabel polysilicon 670 -2326 670 -2326 0 2
rlabel polysilicon 667 -2332 667 -2332 0 3
rlabel polysilicon 670 -2332 670 -2332 0 4
rlabel polysilicon 674 -2326 674 -2326 0 1
rlabel polysilicon 674 -2332 674 -2332 0 3
rlabel polysilicon 681 -2326 681 -2326 0 1
rlabel polysilicon 681 -2332 681 -2332 0 3
rlabel polysilicon 688 -2326 688 -2326 0 1
rlabel polysilicon 688 -2332 688 -2332 0 3
rlabel polysilicon 695 -2326 695 -2326 0 1
rlabel polysilicon 695 -2332 695 -2332 0 3
rlabel polysilicon 702 -2326 702 -2326 0 1
rlabel polysilicon 705 -2326 705 -2326 0 2
rlabel polysilicon 702 -2332 702 -2332 0 3
rlabel polysilicon 709 -2326 709 -2326 0 1
rlabel polysilicon 709 -2332 709 -2332 0 3
rlabel polysilicon 716 -2326 716 -2326 0 1
rlabel polysilicon 716 -2332 716 -2332 0 3
rlabel polysilicon 723 -2326 723 -2326 0 1
rlabel polysilicon 726 -2326 726 -2326 0 2
rlabel polysilicon 723 -2332 723 -2332 0 3
rlabel polysilicon 726 -2332 726 -2332 0 4
rlabel polysilicon 730 -2326 730 -2326 0 1
rlabel polysilicon 730 -2332 730 -2332 0 3
rlabel polysilicon 737 -2326 737 -2326 0 1
rlabel polysilicon 737 -2332 737 -2332 0 3
rlabel polysilicon 744 -2326 744 -2326 0 1
rlabel polysilicon 744 -2332 744 -2332 0 3
rlabel polysilicon 751 -2326 751 -2326 0 1
rlabel polysilicon 751 -2332 751 -2332 0 3
rlabel polysilicon 758 -2326 758 -2326 0 1
rlabel polysilicon 758 -2332 758 -2332 0 3
rlabel polysilicon 765 -2326 765 -2326 0 1
rlabel polysilicon 768 -2332 768 -2332 0 4
rlabel polysilicon 772 -2326 772 -2326 0 1
rlabel polysilicon 772 -2332 772 -2332 0 3
rlabel polysilicon 779 -2326 779 -2326 0 1
rlabel polysilicon 782 -2326 782 -2326 0 2
rlabel polysilicon 782 -2332 782 -2332 0 4
rlabel polysilicon 786 -2326 786 -2326 0 1
rlabel polysilicon 786 -2332 786 -2332 0 3
rlabel polysilicon 793 -2326 793 -2326 0 1
rlabel polysilicon 793 -2332 793 -2332 0 3
rlabel polysilicon 800 -2326 800 -2326 0 1
rlabel polysilicon 800 -2332 800 -2332 0 3
rlabel polysilicon 807 -2326 807 -2326 0 1
rlabel polysilicon 807 -2332 807 -2332 0 3
rlabel polysilicon 814 -2326 814 -2326 0 1
rlabel polysilicon 814 -2332 814 -2332 0 3
rlabel polysilicon 821 -2326 821 -2326 0 1
rlabel polysilicon 821 -2332 821 -2332 0 3
rlabel polysilicon 828 -2326 828 -2326 0 1
rlabel polysilicon 828 -2332 828 -2332 0 3
rlabel polysilicon 835 -2326 835 -2326 0 1
rlabel polysilicon 835 -2332 835 -2332 0 3
rlabel polysilicon 842 -2326 842 -2326 0 1
rlabel polysilicon 842 -2332 842 -2332 0 3
rlabel polysilicon 849 -2326 849 -2326 0 1
rlabel polysilicon 849 -2332 849 -2332 0 3
rlabel polysilicon 856 -2326 856 -2326 0 1
rlabel polysilicon 859 -2326 859 -2326 0 2
rlabel polysilicon 856 -2332 856 -2332 0 3
rlabel polysilicon 859 -2332 859 -2332 0 4
rlabel polysilicon 863 -2326 863 -2326 0 1
rlabel polysilicon 863 -2332 863 -2332 0 3
rlabel polysilicon 870 -2326 870 -2326 0 1
rlabel polysilicon 870 -2332 870 -2332 0 3
rlabel polysilicon 877 -2326 877 -2326 0 1
rlabel polysilicon 877 -2332 877 -2332 0 3
rlabel polysilicon 884 -2326 884 -2326 0 1
rlabel polysilicon 884 -2332 884 -2332 0 3
rlabel polysilicon 891 -2326 891 -2326 0 1
rlabel polysilicon 891 -2332 891 -2332 0 3
rlabel polysilicon 898 -2326 898 -2326 0 1
rlabel polysilicon 898 -2332 898 -2332 0 3
rlabel polysilicon 905 -2326 905 -2326 0 1
rlabel polysilicon 905 -2332 905 -2332 0 3
rlabel polysilicon 912 -2326 912 -2326 0 1
rlabel polysilicon 912 -2332 912 -2332 0 3
rlabel polysilicon 919 -2326 919 -2326 0 1
rlabel polysilicon 919 -2332 919 -2332 0 3
rlabel polysilicon 922 -2332 922 -2332 0 4
rlabel polysilicon 926 -2326 926 -2326 0 1
rlabel polysilicon 926 -2332 926 -2332 0 3
rlabel polysilicon 936 -2326 936 -2326 0 2
rlabel polysilicon 933 -2332 933 -2332 0 3
rlabel polysilicon 936 -2332 936 -2332 0 4
rlabel polysilicon 940 -2326 940 -2326 0 1
rlabel polysilicon 940 -2332 940 -2332 0 3
rlabel polysilicon 947 -2326 947 -2326 0 1
rlabel polysilicon 947 -2332 947 -2332 0 3
rlabel polysilicon 954 -2326 954 -2326 0 1
rlabel polysilicon 954 -2332 954 -2332 0 3
rlabel polysilicon 961 -2326 961 -2326 0 1
rlabel polysilicon 961 -2332 961 -2332 0 3
rlabel polysilicon 968 -2326 968 -2326 0 1
rlabel polysilicon 968 -2332 968 -2332 0 3
rlabel polysilicon 975 -2326 975 -2326 0 1
rlabel polysilicon 978 -2326 978 -2326 0 2
rlabel polysilicon 975 -2332 975 -2332 0 3
rlabel polysilicon 978 -2332 978 -2332 0 4
rlabel polysilicon 982 -2326 982 -2326 0 1
rlabel polysilicon 982 -2332 982 -2332 0 3
rlabel polysilicon 989 -2326 989 -2326 0 1
rlabel polysilicon 992 -2326 992 -2326 0 2
rlabel polysilicon 989 -2332 989 -2332 0 3
rlabel polysilicon 992 -2332 992 -2332 0 4
rlabel polysilicon 996 -2326 996 -2326 0 1
rlabel polysilicon 996 -2332 996 -2332 0 3
rlabel polysilicon 1003 -2326 1003 -2326 0 1
rlabel polysilicon 1003 -2332 1003 -2332 0 3
rlabel polysilicon 1010 -2326 1010 -2326 0 1
rlabel polysilicon 1010 -2332 1010 -2332 0 3
rlabel polysilicon 1017 -2326 1017 -2326 0 1
rlabel polysilicon 1017 -2332 1017 -2332 0 3
rlabel polysilicon 1024 -2326 1024 -2326 0 1
rlabel polysilicon 1024 -2332 1024 -2332 0 3
rlabel polysilicon 1031 -2326 1031 -2326 0 1
rlabel polysilicon 1031 -2332 1031 -2332 0 3
rlabel polysilicon 1041 -2326 1041 -2326 0 2
rlabel polysilicon 1038 -2332 1038 -2332 0 3
rlabel polysilicon 1041 -2332 1041 -2332 0 4
rlabel polysilicon 1045 -2326 1045 -2326 0 1
rlabel polysilicon 1045 -2332 1045 -2332 0 3
rlabel polysilicon 1052 -2326 1052 -2326 0 1
rlabel polysilicon 1052 -2332 1052 -2332 0 3
rlabel polysilicon 1059 -2326 1059 -2326 0 1
rlabel polysilicon 1059 -2332 1059 -2332 0 3
rlabel polysilicon 1066 -2326 1066 -2326 0 1
rlabel polysilicon 1066 -2332 1066 -2332 0 3
rlabel polysilicon 1073 -2326 1073 -2326 0 1
rlabel polysilicon 1073 -2332 1073 -2332 0 3
rlabel polysilicon 1080 -2326 1080 -2326 0 1
rlabel polysilicon 1080 -2332 1080 -2332 0 3
rlabel polysilicon 1087 -2326 1087 -2326 0 1
rlabel polysilicon 1087 -2332 1087 -2332 0 3
rlabel polysilicon 1094 -2326 1094 -2326 0 1
rlabel polysilicon 1094 -2332 1094 -2332 0 3
rlabel polysilicon 1101 -2326 1101 -2326 0 1
rlabel polysilicon 1101 -2332 1101 -2332 0 3
rlabel polysilicon 1108 -2326 1108 -2326 0 1
rlabel polysilicon 1108 -2332 1108 -2332 0 3
rlabel polysilicon 1115 -2326 1115 -2326 0 1
rlabel polysilicon 1115 -2332 1115 -2332 0 3
rlabel polysilicon 1122 -2326 1122 -2326 0 1
rlabel polysilicon 1122 -2332 1122 -2332 0 3
rlabel polysilicon 1129 -2326 1129 -2326 0 1
rlabel polysilicon 1129 -2332 1129 -2332 0 3
rlabel polysilicon 1136 -2326 1136 -2326 0 1
rlabel polysilicon 1139 -2326 1139 -2326 0 2
rlabel polysilicon 1136 -2332 1136 -2332 0 3
rlabel polysilicon 1139 -2332 1139 -2332 0 4
rlabel polysilicon 1143 -2326 1143 -2326 0 1
rlabel polysilicon 1143 -2332 1143 -2332 0 3
rlabel polysilicon 1150 -2326 1150 -2326 0 1
rlabel polysilicon 1150 -2332 1150 -2332 0 3
rlabel polysilicon 1157 -2326 1157 -2326 0 1
rlabel polysilicon 1157 -2332 1157 -2332 0 3
rlabel polysilicon 1164 -2326 1164 -2326 0 1
rlabel polysilicon 1164 -2332 1164 -2332 0 3
rlabel polysilicon 1171 -2326 1171 -2326 0 1
rlabel polysilicon 1171 -2332 1171 -2332 0 3
rlabel polysilicon 1178 -2326 1178 -2326 0 1
rlabel polysilicon 1178 -2332 1178 -2332 0 3
rlabel polysilicon 1185 -2326 1185 -2326 0 1
rlabel polysilicon 1185 -2332 1185 -2332 0 3
rlabel polysilicon 1192 -2326 1192 -2326 0 1
rlabel polysilicon 1192 -2332 1192 -2332 0 3
rlabel polysilicon 1199 -2326 1199 -2326 0 1
rlabel polysilicon 1199 -2332 1199 -2332 0 3
rlabel polysilicon 1206 -2326 1206 -2326 0 1
rlabel polysilicon 1206 -2332 1206 -2332 0 3
rlabel polysilicon 1213 -2326 1213 -2326 0 1
rlabel polysilicon 1213 -2332 1213 -2332 0 3
rlabel polysilicon 1220 -2326 1220 -2326 0 1
rlabel polysilicon 1220 -2332 1220 -2332 0 3
rlabel polysilicon 1227 -2326 1227 -2326 0 1
rlabel polysilicon 1227 -2332 1227 -2332 0 3
rlabel polysilicon 1234 -2326 1234 -2326 0 1
rlabel polysilicon 1234 -2332 1234 -2332 0 3
rlabel polysilicon 1241 -2326 1241 -2326 0 1
rlabel polysilicon 1241 -2332 1241 -2332 0 3
rlabel polysilicon 1248 -2326 1248 -2326 0 1
rlabel polysilicon 1248 -2332 1248 -2332 0 3
rlabel polysilicon 1251 -2332 1251 -2332 0 4
rlabel polysilicon 1255 -2326 1255 -2326 0 1
rlabel polysilicon 1255 -2332 1255 -2332 0 3
rlabel polysilicon 1262 -2326 1262 -2326 0 1
rlabel polysilicon 1262 -2332 1262 -2332 0 3
rlabel polysilicon 1269 -2326 1269 -2326 0 1
rlabel polysilicon 1269 -2332 1269 -2332 0 3
rlabel polysilicon 1276 -2326 1276 -2326 0 1
rlabel polysilicon 1276 -2332 1276 -2332 0 3
rlabel polysilicon 1283 -2326 1283 -2326 0 1
rlabel polysilicon 1283 -2332 1283 -2332 0 3
rlabel polysilicon 1290 -2326 1290 -2326 0 1
rlabel polysilicon 1293 -2326 1293 -2326 0 2
rlabel polysilicon 1290 -2332 1290 -2332 0 3
rlabel polysilicon 1293 -2332 1293 -2332 0 4
rlabel polysilicon 1297 -2326 1297 -2326 0 1
rlabel polysilicon 1297 -2332 1297 -2332 0 3
rlabel polysilicon 1304 -2326 1304 -2326 0 1
rlabel polysilicon 1304 -2332 1304 -2332 0 3
rlabel polysilicon 1311 -2326 1311 -2326 0 1
rlabel polysilicon 1311 -2332 1311 -2332 0 3
rlabel polysilicon 1318 -2326 1318 -2326 0 1
rlabel polysilicon 1321 -2326 1321 -2326 0 2
rlabel polysilicon 1318 -2332 1318 -2332 0 3
rlabel polysilicon 1321 -2332 1321 -2332 0 4
rlabel polysilicon 1325 -2326 1325 -2326 0 1
rlabel polysilicon 1325 -2332 1325 -2332 0 3
rlabel polysilicon 1332 -2326 1332 -2326 0 1
rlabel polysilicon 1332 -2332 1332 -2332 0 3
rlabel polysilicon 1339 -2326 1339 -2326 0 1
rlabel polysilicon 1339 -2332 1339 -2332 0 3
rlabel polysilicon 1346 -2326 1346 -2326 0 1
rlabel polysilicon 1346 -2332 1346 -2332 0 3
rlabel polysilicon 1353 -2326 1353 -2326 0 1
rlabel polysilicon 1353 -2332 1353 -2332 0 3
rlabel polysilicon 1360 -2326 1360 -2326 0 1
rlabel polysilicon 1360 -2332 1360 -2332 0 3
rlabel polysilicon 1367 -2326 1367 -2326 0 1
rlabel polysilicon 1367 -2332 1367 -2332 0 3
rlabel polysilicon 1374 -2326 1374 -2326 0 1
rlabel polysilicon 1374 -2332 1374 -2332 0 3
rlabel polysilicon 1381 -2326 1381 -2326 0 1
rlabel polysilicon 1381 -2332 1381 -2332 0 3
rlabel polysilicon 1388 -2326 1388 -2326 0 1
rlabel polysilicon 1388 -2332 1388 -2332 0 3
rlabel polysilicon 1395 -2326 1395 -2326 0 1
rlabel polysilicon 1398 -2326 1398 -2326 0 2
rlabel polysilicon 1398 -2332 1398 -2332 0 4
rlabel polysilicon 1402 -2326 1402 -2326 0 1
rlabel polysilicon 1402 -2332 1402 -2332 0 3
rlabel polysilicon 1409 -2326 1409 -2326 0 1
rlabel polysilicon 1409 -2332 1409 -2332 0 3
rlabel polysilicon 1416 -2326 1416 -2326 0 1
rlabel polysilicon 1416 -2332 1416 -2332 0 3
rlabel polysilicon 1423 -2326 1423 -2326 0 1
rlabel polysilicon 1423 -2332 1423 -2332 0 3
rlabel polysilicon 1430 -2326 1430 -2326 0 1
rlabel polysilicon 1430 -2332 1430 -2332 0 3
rlabel polysilicon 1437 -2326 1437 -2326 0 1
rlabel polysilicon 1437 -2332 1437 -2332 0 3
rlabel polysilicon 1444 -2326 1444 -2326 0 1
rlabel polysilicon 1444 -2332 1444 -2332 0 3
rlabel polysilicon 1451 -2326 1451 -2326 0 1
rlabel polysilicon 1451 -2332 1451 -2332 0 3
rlabel polysilicon 1458 -2326 1458 -2326 0 1
rlabel polysilicon 1458 -2332 1458 -2332 0 3
rlabel polysilicon 1465 -2326 1465 -2326 0 1
rlabel polysilicon 1465 -2332 1465 -2332 0 3
rlabel polysilicon 1472 -2326 1472 -2326 0 1
rlabel polysilicon 1472 -2332 1472 -2332 0 3
rlabel polysilicon 1479 -2326 1479 -2326 0 1
rlabel polysilicon 1479 -2332 1479 -2332 0 3
rlabel polysilicon 1486 -2326 1486 -2326 0 1
rlabel polysilicon 1486 -2332 1486 -2332 0 3
rlabel polysilicon 1493 -2326 1493 -2326 0 1
rlabel polysilicon 1496 -2326 1496 -2326 0 2
rlabel polysilicon 1493 -2332 1493 -2332 0 3
rlabel polysilicon 1496 -2332 1496 -2332 0 4
rlabel polysilicon 1500 -2326 1500 -2326 0 1
rlabel polysilicon 1503 -2326 1503 -2326 0 2
rlabel polysilicon 1500 -2332 1500 -2332 0 3
rlabel polysilicon 1507 -2326 1507 -2326 0 1
rlabel polysilicon 1507 -2332 1507 -2332 0 3
rlabel polysilicon 1514 -2326 1514 -2326 0 1
rlabel polysilicon 1517 -2326 1517 -2326 0 2
rlabel polysilicon 1517 -2332 1517 -2332 0 4
rlabel polysilicon 1521 -2326 1521 -2326 0 1
rlabel polysilicon 1521 -2332 1521 -2332 0 3
rlabel polysilicon 1528 -2326 1528 -2326 0 1
rlabel polysilicon 1528 -2332 1528 -2332 0 3
rlabel polysilicon 1535 -2326 1535 -2326 0 1
rlabel polysilicon 1535 -2332 1535 -2332 0 3
rlabel polysilicon 1542 -2326 1542 -2326 0 1
rlabel polysilicon 1545 -2326 1545 -2326 0 2
rlabel polysilicon 1542 -2332 1542 -2332 0 3
rlabel polysilicon 1545 -2332 1545 -2332 0 4
rlabel polysilicon 1549 -2326 1549 -2326 0 1
rlabel polysilicon 1549 -2332 1549 -2332 0 3
rlabel polysilicon 1556 -2326 1556 -2326 0 1
rlabel polysilicon 1556 -2332 1556 -2332 0 3
rlabel polysilicon 1563 -2326 1563 -2326 0 1
rlabel polysilicon 1563 -2332 1563 -2332 0 3
rlabel polysilicon 1570 -2326 1570 -2326 0 1
rlabel polysilicon 1570 -2332 1570 -2332 0 3
rlabel polysilicon 1577 -2326 1577 -2326 0 1
rlabel polysilicon 1577 -2332 1577 -2332 0 3
rlabel polysilicon 1584 -2326 1584 -2326 0 1
rlabel polysilicon 1584 -2332 1584 -2332 0 3
rlabel polysilicon 1591 -2326 1591 -2326 0 1
rlabel polysilicon 1591 -2332 1591 -2332 0 3
rlabel polysilicon 1598 -2326 1598 -2326 0 1
rlabel polysilicon 1598 -2332 1598 -2332 0 3
rlabel polysilicon 1605 -2326 1605 -2326 0 1
rlabel polysilicon 1605 -2332 1605 -2332 0 3
rlabel polysilicon 1612 -2326 1612 -2326 0 1
rlabel polysilicon 1612 -2332 1612 -2332 0 3
rlabel polysilicon 1619 -2326 1619 -2326 0 1
rlabel polysilicon 1619 -2332 1619 -2332 0 3
rlabel polysilicon 1626 -2326 1626 -2326 0 1
rlabel polysilicon 1629 -2326 1629 -2326 0 2
rlabel polysilicon 1626 -2332 1626 -2332 0 3
rlabel polysilicon 1629 -2332 1629 -2332 0 4
rlabel polysilicon 1633 -2326 1633 -2326 0 1
rlabel polysilicon 1633 -2332 1633 -2332 0 3
rlabel polysilicon 1640 -2326 1640 -2326 0 1
rlabel polysilicon 1640 -2332 1640 -2332 0 3
rlabel polysilicon 1647 -2326 1647 -2326 0 1
rlabel polysilicon 1647 -2332 1647 -2332 0 3
rlabel polysilicon 1654 -2326 1654 -2326 0 1
rlabel polysilicon 1654 -2332 1654 -2332 0 3
rlabel polysilicon 1661 -2326 1661 -2326 0 1
rlabel polysilicon 1661 -2332 1661 -2332 0 3
rlabel polysilicon 1668 -2326 1668 -2326 0 1
rlabel polysilicon 1668 -2332 1668 -2332 0 3
rlabel polysilicon 1675 -2326 1675 -2326 0 1
rlabel polysilicon 1675 -2332 1675 -2332 0 3
rlabel polysilicon 1685 -2326 1685 -2326 0 2
rlabel polysilicon 1682 -2332 1682 -2332 0 3
rlabel polysilicon 1685 -2332 1685 -2332 0 4
rlabel polysilicon 1689 -2326 1689 -2326 0 1
rlabel polysilicon 1689 -2332 1689 -2332 0 3
rlabel polysilicon 1696 -2326 1696 -2326 0 1
rlabel polysilicon 1696 -2332 1696 -2332 0 3
rlabel polysilicon 1703 -2326 1703 -2326 0 1
rlabel polysilicon 1703 -2332 1703 -2332 0 3
rlabel polysilicon 1710 -2326 1710 -2326 0 1
rlabel polysilicon 1710 -2332 1710 -2332 0 3
rlabel polysilicon 1717 -2326 1717 -2326 0 1
rlabel polysilicon 1717 -2332 1717 -2332 0 3
rlabel polysilicon 1724 -2326 1724 -2326 0 1
rlabel polysilicon 1724 -2332 1724 -2332 0 3
rlabel polysilicon 1731 -2326 1731 -2326 0 1
rlabel polysilicon 1731 -2332 1731 -2332 0 3
rlabel polysilicon 1738 -2326 1738 -2326 0 1
rlabel polysilicon 1738 -2332 1738 -2332 0 3
rlabel polysilicon 1745 -2326 1745 -2326 0 1
rlabel polysilicon 1745 -2332 1745 -2332 0 3
rlabel polysilicon 1752 -2326 1752 -2326 0 1
rlabel polysilicon 1752 -2332 1752 -2332 0 3
rlabel polysilicon 1759 -2326 1759 -2326 0 1
rlabel polysilicon 1759 -2332 1759 -2332 0 3
rlabel polysilicon 1766 -2326 1766 -2326 0 1
rlabel polysilicon 1766 -2332 1766 -2332 0 3
rlabel polysilicon 1773 -2326 1773 -2326 0 1
rlabel polysilicon 1773 -2332 1773 -2332 0 3
rlabel polysilicon 1780 -2326 1780 -2326 0 1
rlabel polysilicon 1780 -2332 1780 -2332 0 3
rlabel polysilicon 1787 -2326 1787 -2326 0 1
rlabel polysilicon 1787 -2332 1787 -2332 0 3
rlabel polysilicon 1794 -2326 1794 -2326 0 1
rlabel polysilicon 1794 -2332 1794 -2332 0 3
rlabel polysilicon 1801 -2326 1801 -2326 0 1
rlabel polysilicon 1801 -2332 1801 -2332 0 3
rlabel polysilicon 1808 -2326 1808 -2326 0 1
rlabel polysilicon 1808 -2332 1808 -2332 0 3
rlabel polysilicon 1815 -2326 1815 -2326 0 1
rlabel polysilicon 1815 -2332 1815 -2332 0 3
rlabel polysilicon 1822 -2326 1822 -2326 0 1
rlabel polysilicon 1822 -2332 1822 -2332 0 3
rlabel polysilicon 1829 -2326 1829 -2326 0 1
rlabel polysilicon 1829 -2332 1829 -2332 0 3
rlabel polysilicon 1836 -2326 1836 -2326 0 1
rlabel polysilicon 1836 -2332 1836 -2332 0 3
rlabel polysilicon 1843 -2326 1843 -2326 0 1
rlabel polysilicon 1843 -2332 1843 -2332 0 3
rlabel polysilicon 1850 -2326 1850 -2326 0 1
rlabel polysilicon 1850 -2332 1850 -2332 0 3
rlabel polysilicon 1853 -2332 1853 -2332 0 4
rlabel polysilicon 1857 -2326 1857 -2326 0 1
rlabel polysilicon 1857 -2332 1857 -2332 0 3
rlabel polysilicon 1864 -2326 1864 -2326 0 1
rlabel polysilicon 1864 -2332 1864 -2332 0 3
rlabel polysilicon 1871 -2326 1871 -2326 0 1
rlabel polysilicon 1871 -2332 1871 -2332 0 3
rlabel polysilicon 1878 -2326 1878 -2326 0 1
rlabel polysilicon 1878 -2332 1878 -2332 0 3
rlabel polysilicon 1885 -2326 1885 -2326 0 1
rlabel polysilicon 1885 -2332 1885 -2332 0 3
rlabel polysilicon 1895 -2326 1895 -2326 0 2
rlabel polysilicon 1895 -2332 1895 -2332 0 4
rlabel polysilicon 1899 -2326 1899 -2326 0 1
rlabel polysilicon 1899 -2332 1899 -2332 0 3
rlabel polysilicon 1906 -2326 1906 -2326 0 1
rlabel polysilicon 1906 -2332 1906 -2332 0 3
rlabel polysilicon 1913 -2326 1913 -2326 0 1
rlabel polysilicon 1913 -2332 1913 -2332 0 3
rlabel polysilicon 1920 -2326 1920 -2326 0 1
rlabel polysilicon 1920 -2332 1920 -2332 0 3
rlabel polysilicon 1927 -2326 1927 -2326 0 1
rlabel polysilicon 1927 -2332 1927 -2332 0 3
rlabel polysilicon 1934 -2326 1934 -2326 0 1
rlabel polysilicon 1937 -2326 1937 -2326 0 2
rlabel polysilicon 1934 -2332 1934 -2332 0 3
rlabel polysilicon 1937 -2332 1937 -2332 0 4
rlabel polysilicon 1941 -2326 1941 -2326 0 1
rlabel polysilicon 1941 -2332 1941 -2332 0 3
rlabel polysilicon 1948 -2326 1948 -2326 0 1
rlabel polysilicon 1948 -2332 1948 -2332 0 3
rlabel polysilicon 1955 -2326 1955 -2326 0 1
rlabel polysilicon 1955 -2332 1955 -2332 0 3
rlabel polysilicon 1962 -2326 1962 -2326 0 1
rlabel polysilicon 1962 -2332 1962 -2332 0 3
rlabel polysilicon 1969 -2326 1969 -2326 0 1
rlabel polysilicon 1969 -2332 1969 -2332 0 3
rlabel polysilicon 1976 -2326 1976 -2326 0 1
rlabel polysilicon 1979 -2326 1979 -2326 0 2
rlabel polysilicon 1979 -2332 1979 -2332 0 4
rlabel polysilicon 1983 -2326 1983 -2326 0 1
rlabel polysilicon 1983 -2332 1983 -2332 0 3
rlabel polysilicon 1990 -2326 1990 -2326 0 1
rlabel polysilicon 1990 -2332 1990 -2332 0 3
rlabel polysilicon 1997 -2326 1997 -2326 0 1
rlabel polysilicon 1997 -2332 1997 -2332 0 3
rlabel polysilicon 2004 -2326 2004 -2326 0 1
rlabel polysilicon 2004 -2332 2004 -2332 0 3
rlabel polysilicon 2011 -2326 2011 -2326 0 1
rlabel polysilicon 2011 -2332 2011 -2332 0 3
rlabel polysilicon 2018 -2326 2018 -2326 0 1
rlabel polysilicon 2018 -2332 2018 -2332 0 3
rlabel polysilicon 2025 -2326 2025 -2326 0 1
rlabel polysilicon 2025 -2332 2025 -2332 0 3
rlabel polysilicon 2032 -2326 2032 -2326 0 1
rlabel polysilicon 2032 -2332 2032 -2332 0 3
rlabel polysilicon 2039 -2326 2039 -2326 0 1
rlabel polysilicon 2039 -2332 2039 -2332 0 3
rlabel polysilicon 2046 -2326 2046 -2326 0 1
rlabel polysilicon 2046 -2332 2046 -2332 0 3
rlabel polysilicon 2053 -2326 2053 -2326 0 1
rlabel polysilicon 2053 -2332 2053 -2332 0 3
rlabel polysilicon 2060 -2326 2060 -2326 0 1
rlabel polysilicon 2060 -2332 2060 -2332 0 3
rlabel polysilicon 2067 -2326 2067 -2326 0 1
rlabel polysilicon 2067 -2332 2067 -2332 0 3
rlabel polysilicon 2074 -2326 2074 -2326 0 1
rlabel polysilicon 2074 -2332 2074 -2332 0 3
rlabel polysilicon 2081 -2326 2081 -2326 0 1
rlabel polysilicon 2081 -2332 2081 -2332 0 3
rlabel polysilicon 2088 -2326 2088 -2326 0 1
rlabel polysilicon 2088 -2332 2088 -2332 0 3
rlabel polysilicon 2095 -2326 2095 -2326 0 1
rlabel polysilicon 2095 -2332 2095 -2332 0 3
rlabel polysilicon 2102 -2326 2102 -2326 0 1
rlabel polysilicon 2102 -2332 2102 -2332 0 3
rlabel polysilicon 2109 -2326 2109 -2326 0 1
rlabel polysilicon 2109 -2332 2109 -2332 0 3
rlabel polysilicon 2116 -2326 2116 -2326 0 1
rlabel polysilicon 2116 -2332 2116 -2332 0 3
rlabel polysilicon 2123 -2326 2123 -2326 0 1
rlabel polysilicon 2123 -2332 2123 -2332 0 3
rlabel polysilicon 2130 -2326 2130 -2326 0 1
rlabel polysilicon 2130 -2332 2130 -2332 0 3
rlabel polysilicon 2137 -2326 2137 -2326 0 1
rlabel polysilicon 2137 -2332 2137 -2332 0 3
rlabel polysilicon 2144 -2326 2144 -2326 0 1
rlabel polysilicon 2144 -2332 2144 -2332 0 3
rlabel polysilicon 2151 -2326 2151 -2326 0 1
rlabel polysilicon 2151 -2332 2151 -2332 0 3
rlabel polysilicon 2158 -2326 2158 -2326 0 1
rlabel polysilicon 2158 -2332 2158 -2332 0 3
rlabel polysilicon 2165 -2326 2165 -2326 0 1
rlabel polysilicon 2165 -2332 2165 -2332 0 3
rlabel polysilicon 2172 -2326 2172 -2326 0 1
rlabel polysilicon 2172 -2332 2172 -2332 0 3
rlabel polysilicon 2179 -2326 2179 -2326 0 1
rlabel polysilicon 2179 -2332 2179 -2332 0 3
rlabel polysilicon 2186 -2326 2186 -2326 0 1
rlabel polysilicon 2186 -2332 2186 -2332 0 3
rlabel polysilicon 2193 -2326 2193 -2326 0 1
rlabel polysilicon 2193 -2332 2193 -2332 0 3
rlabel polysilicon 2200 -2326 2200 -2326 0 1
rlabel polysilicon 2200 -2332 2200 -2332 0 3
rlabel polysilicon 2207 -2326 2207 -2326 0 1
rlabel polysilicon 2207 -2332 2207 -2332 0 3
rlabel polysilicon 2214 -2326 2214 -2326 0 1
rlabel polysilicon 2214 -2332 2214 -2332 0 3
rlabel polysilicon 2221 -2326 2221 -2326 0 1
rlabel polysilicon 2221 -2332 2221 -2332 0 3
rlabel polysilicon 2228 -2326 2228 -2326 0 1
rlabel polysilicon 2228 -2332 2228 -2332 0 3
rlabel polysilicon 2235 -2326 2235 -2326 0 1
rlabel polysilicon 2235 -2332 2235 -2332 0 3
rlabel polysilicon 2242 -2326 2242 -2326 0 1
rlabel polysilicon 2242 -2332 2242 -2332 0 3
rlabel polysilicon 2249 -2326 2249 -2326 0 1
rlabel polysilicon 2249 -2332 2249 -2332 0 3
rlabel polysilicon 2256 -2326 2256 -2326 0 1
rlabel polysilicon 2256 -2332 2256 -2332 0 3
rlabel polysilicon 2263 -2326 2263 -2326 0 1
rlabel polysilicon 2263 -2332 2263 -2332 0 3
rlabel polysilicon 2270 -2326 2270 -2326 0 1
rlabel polysilicon 2270 -2332 2270 -2332 0 3
rlabel polysilicon 2277 -2326 2277 -2326 0 1
rlabel polysilicon 2277 -2332 2277 -2332 0 3
rlabel polysilicon 2284 -2326 2284 -2326 0 1
rlabel polysilicon 2284 -2332 2284 -2332 0 3
rlabel polysilicon 2291 -2326 2291 -2326 0 1
rlabel polysilicon 2291 -2332 2291 -2332 0 3
rlabel polysilicon 2298 -2326 2298 -2326 0 1
rlabel polysilicon 2298 -2332 2298 -2332 0 3
rlabel polysilicon 2305 -2326 2305 -2326 0 1
rlabel polysilicon 2305 -2332 2305 -2332 0 3
rlabel polysilicon 2312 -2326 2312 -2326 0 1
rlabel polysilicon 2312 -2332 2312 -2332 0 3
rlabel polysilicon 2319 -2326 2319 -2326 0 1
rlabel polysilicon 2319 -2332 2319 -2332 0 3
rlabel polysilicon 2326 -2326 2326 -2326 0 1
rlabel polysilicon 2326 -2332 2326 -2332 0 3
rlabel polysilicon 2333 -2326 2333 -2326 0 1
rlabel polysilicon 2336 -2326 2336 -2326 0 2
rlabel polysilicon 2333 -2332 2333 -2332 0 3
rlabel polysilicon 2336 -2332 2336 -2332 0 4
rlabel polysilicon 2343 -2326 2343 -2326 0 2
rlabel polysilicon 2343 -2332 2343 -2332 0 4
rlabel polysilicon 2347 -2326 2347 -2326 0 1
rlabel polysilicon 2347 -2332 2347 -2332 0 3
rlabel polysilicon 2 -2499 2 -2499 0 1
rlabel polysilicon 5 -2499 5 -2499 0 2
rlabel polysilicon 5 -2505 5 -2505 0 4
rlabel polysilicon 9 -2499 9 -2499 0 1
rlabel polysilicon 9 -2505 9 -2505 0 3
rlabel polysilicon 16 -2499 16 -2499 0 1
rlabel polysilicon 19 -2505 19 -2505 0 4
rlabel polysilicon 23 -2499 23 -2499 0 1
rlabel polysilicon 23 -2505 23 -2505 0 3
rlabel polysilicon 30 -2505 30 -2505 0 3
rlabel polysilicon 33 -2505 33 -2505 0 4
rlabel polysilicon 37 -2499 37 -2499 0 1
rlabel polysilicon 37 -2505 37 -2505 0 3
rlabel polysilicon 40 -2505 40 -2505 0 4
rlabel polysilicon 44 -2499 44 -2499 0 1
rlabel polysilicon 44 -2505 44 -2505 0 3
rlabel polysilicon 51 -2499 51 -2499 0 1
rlabel polysilicon 51 -2505 51 -2505 0 3
rlabel polysilicon 58 -2499 58 -2499 0 1
rlabel polysilicon 58 -2505 58 -2505 0 3
rlabel polysilicon 61 -2505 61 -2505 0 4
rlabel polysilicon 65 -2499 65 -2499 0 1
rlabel polysilicon 65 -2505 65 -2505 0 3
rlabel polysilicon 72 -2499 72 -2499 0 1
rlabel polysilicon 72 -2505 72 -2505 0 3
rlabel polysilicon 79 -2499 79 -2499 0 1
rlabel polysilicon 79 -2505 79 -2505 0 3
rlabel polysilicon 86 -2499 86 -2499 0 1
rlabel polysilicon 86 -2505 86 -2505 0 3
rlabel polysilicon 93 -2499 93 -2499 0 1
rlabel polysilicon 96 -2499 96 -2499 0 2
rlabel polysilicon 93 -2505 93 -2505 0 3
rlabel polysilicon 96 -2505 96 -2505 0 4
rlabel polysilicon 100 -2499 100 -2499 0 1
rlabel polysilicon 100 -2505 100 -2505 0 3
rlabel polysilicon 107 -2499 107 -2499 0 1
rlabel polysilicon 110 -2499 110 -2499 0 2
rlabel polysilicon 110 -2505 110 -2505 0 4
rlabel polysilicon 114 -2499 114 -2499 0 1
rlabel polysilicon 114 -2505 114 -2505 0 3
rlabel polysilicon 121 -2499 121 -2499 0 1
rlabel polysilicon 121 -2505 121 -2505 0 3
rlabel polysilicon 128 -2499 128 -2499 0 1
rlabel polysilicon 128 -2505 128 -2505 0 3
rlabel polysilicon 135 -2499 135 -2499 0 1
rlabel polysilicon 135 -2505 135 -2505 0 3
rlabel polysilicon 142 -2499 142 -2499 0 1
rlabel polysilicon 142 -2505 142 -2505 0 3
rlabel polysilicon 149 -2499 149 -2499 0 1
rlabel polysilicon 149 -2505 149 -2505 0 3
rlabel polysilicon 156 -2499 156 -2499 0 1
rlabel polysilicon 156 -2505 156 -2505 0 3
rlabel polysilicon 163 -2499 163 -2499 0 1
rlabel polysilicon 163 -2505 163 -2505 0 3
rlabel polysilicon 166 -2505 166 -2505 0 4
rlabel polysilicon 170 -2499 170 -2499 0 1
rlabel polysilicon 170 -2505 170 -2505 0 3
rlabel polysilicon 177 -2505 177 -2505 0 3
rlabel polysilicon 184 -2499 184 -2499 0 1
rlabel polysilicon 184 -2505 184 -2505 0 3
rlabel polysilicon 191 -2499 191 -2499 0 1
rlabel polysilicon 191 -2505 191 -2505 0 3
rlabel polysilicon 198 -2499 198 -2499 0 1
rlabel polysilicon 198 -2505 198 -2505 0 3
rlabel polysilicon 205 -2499 205 -2499 0 1
rlabel polysilicon 205 -2505 205 -2505 0 3
rlabel polysilicon 212 -2499 212 -2499 0 1
rlabel polysilicon 212 -2505 212 -2505 0 3
rlabel polysilicon 219 -2499 219 -2499 0 1
rlabel polysilicon 219 -2505 219 -2505 0 3
rlabel polysilicon 226 -2499 226 -2499 0 1
rlabel polysilicon 226 -2505 226 -2505 0 3
rlabel polysilicon 233 -2499 233 -2499 0 1
rlabel polysilicon 233 -2505 233 -2505 0 3
rlabel polysilicon 240 -2499 240 -2499 0 1
rlabel polysilicon 240 -2505 240 -2505 0 3
rlabel polysilicon 247 -2499 247 -2499 0 1
rlabel polysilicon 247 -2505 247 -2505 0 3
rlabel polysilicon 254 -2499 254 -2499 0 1
rlabel polysilicon 254 -2505 254 -2505 0 3
rlabel polysilicon 261 -2499 261 -2499 0 1
rlabel polysilicon 261 -2505 261 -2505 0 3
rlabel polysilicon 268 -2499 268 -2499 0 1
rlabel polysilicon 268 -2505 268 -2505 0 3
rlabel polysilicon 275 -2499 275 -2499 0 1
rlabel polysilicon 275 -2505 275 -2505 0 3
rlabel polysilicon 282 -2499 282 -2499 0 1
rlabel polysilicon 282 -2505 282 -2505 0 3
rlabel polysilicon 289 -2499 289 -2499 0 1
rlabel polysilicon 289 -2505 289 -2505 0 3
rlabel polysilicon 296 -2499 296 -2499 0 1
rlabel polysilicon 296 -2505 296 -2505 0 3
rlabel polysilicon 303 -2499 303 -2499 0 1
rlabel polysilicon 303 -2505 303 -2505 0 3
rlabel polysilicon 310 -2499 310 -2499 0 1
rlabel polysilicon 310 -2505 310 -2505 0 3
rlabel polysilicon 317 -2499 317 -2499 0 1
rlabel polysilicon 317 -2505 317 -2505 0 3
rlabel polysilicon 324 -2499 324 -2499 0 1
rlabel polysilicon 324 -2505 324 -2505 0 3
rlabel polysilicon 331 -2499 331 -2499 0 1
rlabel polysilicon 331 -2505 331 -2505 0 3
rlabel polysilicon 338 -2499 338 -2499 0 1
rlabel polysilicon 338 -2505 338 -2505 0 3
rlabel polysilicon 345 -2499 345 -2499 0 1
rlabel polysilicon 345 -2505 345 -2505 0 3
rlabel polysilicon 352 -2499 352 -2499 0 1
rlabel polysilicon 352 -2505 352 -2505 0 3
rlabel polysilicon 359 -2499 359 -2499 0 1
rlabel polysilicon 359 -2505 359 -2505 0 3
rlabel polysilicon 366 -2499 366 -2499 0 1
rlabel polysilicon 366 -2505 366 -2505 0 3
rlabel polysilicon 373 -2499 373 -2499 0 1
rlabel polysilicon 373 -2505 373 -2505 0 3
rlabel polysilicon 380 -2499 380 -2499 0 1
rlabel polysilicon 380 -2505 380 -2505 0 3
rlabel polysilicon 387 -2499 387 -2499 0 1
rlabel polysilicon 387 -2505 387 -2505 0 3
rlabel polysilicon 394 -2499 394 -2499 0 1
rlabel polysilicon 394 -2505 394 -2505 0 3
rlabel polysilicon 401 -2499 401 -2499 0 1
rlabel polysilicon 401 -2505 401 -2505 0 3
rlabel polysilicon 408 -2499 408 -2499 0 1
rlabel polysilicon 408 -2505 408 -2505 0 3
rlabel polysilicon 415 -2499 415 -2499 0 1
rlabel polysilicon 415 -2505 415 -2505 0 3
rlabel polysilicon 422 -2499 422 -2499 0 1
rlabel polysilicon 422 -2505 422 -2505 0 3
rlabel polysilicon 429 -2499 429 -2499 0 1
rlabel polysilicon 429 -2505 429 -2505 0 3
rlabel polysilicon 436 -2499 436 -2499 0 1
rlabel polysilicon 436 -2505 436 -2505 0 3
rlabel polysilicon 443 -2499 443 -2499 0 1
rlabel polysilicon 443 -2505 443 -2505 0 3
rlabel polysilicon 450 -2499 450 -2499 0 1
rlabel polysilicon 450 -2505 450 -2505 0 3
rlabel polysilicon 457 -2499 457 -2499 0 1
rlabel polysilicon 457 -2505 457 -2505 0 3
rlabel polysilicon 464 -2499 464 -2499 0 1
rlabel polysilicon 464 -2505 464 -2505 0 3
rlabel polysilicon 471 -2499 471 -2499 0 1
rlabel polysilicon 471 -2505 471 -2505 0 3
rlabel polysilicon 478 -2499 478 -2499 0 1
rlabel polysilicon 481 -2499 481 -2499 0 2
rlabel polysilicon 478 -2505 478 -2505 0 3
rlabel polysilicon 481 -2505 481 -2505 0 4
rlabel polysilicon 485 -2499 485 -2499 0 1
rlabel polysilicon 485 -2505 485 -2505 0 3
rlabel polysilicon 492 -2499 492 -2499 0 1
rlabel polysilicon 492 -2505 492 -2505 0 3
rlabel polysilicon 499 -2499 499 -2499 0 1
rlabel polysilicon 499 -2505 499 -2505 0 3
rlabel polysilicon 506 -2499 506 -2499 0 1
rlabel polysilicon 506 -2505 506 -2505 0 3
rlabel polysilicon 513 -2499 513 -2499 0 1
rlabel polysilicon 513 -2505 513 -2505 0 3
rlabel polysilicon 520 -2499 520 -2499 0 1
rlabel polysilicon 520 -2505 520 -2505 0 3
rlabel polysilicon 527 -2499 527 -2499 0 1
rlabel polysilicon 527 -2505 527 -2505 0 3
rlabel polysilicon 534 -2499 534 -2499 0 1
rlabel polysilicon 534 -2505 534 -2505 0 3
rlabel polysilicon 541 -2499 541 -2499 0 1
rlabel polysilicon 541 -2505 541 -2505 0 3
rlabel polysilicon 548 -2499 548 -2499 0 1
rlabel polysilicon 548 -2505 548 -2505 0 3
rlabel polysilicon 555 -2499 555 -2499 0 1
rlabel polysilicon 555 -2505 555 -2505 0 3
rlabel polysilicon 562 -2499 562 -2499 0 1
rlabel polysilicon 562 -2505 562 -2505 0 3
rlabel polysilicon 569 -2499 569 -2499 0 1
rlabel polysilicon 569 -2505 569 -2505 0 3
rlabel polysilicon 576 -2499 576 -2499 0 1
rlabel polysilicon 576 -2505 576 -2505 0 3
rlabel polysilicon 583 -2499 583 -2499 0 1
rlabel polysilicon 583 -2505 583 -2505 0 3
rlabel polysilicon 590 -2499 590 -2499 0 1
rlabel polysilicon 590 -2505 590 -2505 0 3
rlabel polysilicon 597 -2499 597 -2499 0 1
rlabel polysilicon 597 -2505 597 -2505 0 3
rlabel polysilicon 604 -2499 604 -2499 0 1
rlabel polysilicon 607 -2499 607 -2499 0 2
rlabel polysilicon 607 -2505 607 -2505 0 4
rlabel polysilicon 611 -2499 611 -2499 0 1
rlabel polysilicon 611 -2505 611 -2505 0 3
rlabel polysilicon 618 -2499 618 -2499 0 1
rlabel polysilicon 618 -2505 618 -2505 0 3
rlabel polysilicon 625 -2499 625 -2499 0 1
rlabel polysilicon 625 -2505 625 -2505 0 3
rlabel polysilicon 632 -2499 632 -2499 0 1
rlabel polysilicon 632 -2505 632 -2505 0 3
rlabel polysilicon 639 -2499 639 -2499 0 1
rlabel polysilicon 639 -2505 639 -2505 0 3
rlabel polysilicon 646 -2499 646 -2499 0 1
rlabel polysilicon 646 -2505 646 -2505 0 3
rlabel polysilicon 653 -2499 653 -2499 0 1
rlabel polysilicon 653 -2505 653 -2505 0 3
rlabel polysilicon 660 -2499 660 -2499 0 1
rlabel polysilicon 660 -2505 660 -2505 0 3
rlabel polysilicon 667 -2499 667 -2499 0 1
rlabel polysilicon 670 -2499 670 -2499 0 2
rlabel polysilicon 667 -2505 667 -2505 0 3
rlabel polysilicon 670 -2505 670 -2505 0 4
rlabel polysilicon 674 -2499 674 -2499 0 1
rlabel polysilicon 674 -2505 674 -2505 0 3
rlabel polysilicon 681 -2499 681 -2499 0 1
rlabel polysilicon 681 -2505 681 -2505 0 3
rlabel polysilicon 688 -2499 688 -2499 0 1
rlabel polysilicon 688 -2505 688 -2505 0 3
rlabel polysilicon 695 -2499 695 -2499 0 1
rlabel polysilicon 695 -2505 695 -2505 0 3
rlabel polysilicon 702 -2499 702 -2499 0 1
rlabel polysilicon 702 -2505 702 -2505 0 3
rlabel polysilicon 709 -2499 709 -2499 0 1
rlabel polysilicon 709 -2505 709 -2505 0 3
rlabel polysilicon 716 -2499 716 -2499 0 1
rlabel polysilicon 716 -2505 716 -2505 0 3
rlabel polysilicon 723 -2499 723 -2499 0 1
rlabel polysilicon 723 -2505 723 -2505 0 3
rlabel polysilicon 730 -2499 730 -2499 0 1
rlabel polysilicon 730 -2505 730 -2505 0 3
rlabel polysilicon 737 -2499 737 -2499 0 1
rlabel polysilicon 740 -2499 740 -2499 0 2
rlabel polysilicon 737 -2505 737 -2505 0 3
rlabel polysilicon 740 -2505 740 -2505 0 4
rlabel polysilicon 744 -2499 744 -2499 0 1
rlabel polysilicon 744 -2505 744 -2505 0 3
rlabel polysilicon 751 -2499 751 -2499 0 1
rlabel polysilicon 751 -2505 751 -2505 0 3
rlabel polysilicon 758 -2499 758 -2499 0 1
rlabel polysilicon 758 -2505 758 -2505 0 3
rlabel polysilicon 765 -2499 765 -2499 0 1
rlabel polysilicon 765 -2505 765 -2505 0 3
rlabel polysilicon 772 -2499 772 -2499 0 1
rlabel polysilicon 775 -2499 775 -2499 0 2
rlabel polysilicon 775 -2505 775 -2505 0 4
rlabel polysilicon 779 -2499 779 -2499 0 1
rlabel polysilicon 779 -2505 779 -2505 0 3
rlabel polysilicon 786 -2499 786 -2499 0 1
rlabel polysilicon 786 -2505 786 -2505 0 3
rlabel polysilicon 793 -2499 793 -2499 0 1
rlabel polysilicon 796 -2499 796 -2499 0 2
rlabel polysilicon 793 -2505 793 -2505 0 3
rlabel polysilicon 796 -2505 796 -2505 0 4
rlabel polysilicon 800 -2499 800 -2499 0 1
rlabel polysilicon 800 -2505 800 -2505 0 3
rlabel polysilicon 807 -2499 807 -2499 0 1
rlabel polysilicon 807 -2505 807 -2505 0 3
rlabel polysilicon 814 -2499 814 -2499 0 1
rlabel polysilicon 814 -2505 814 -2505 0 3
rlabel polysilicon 821 -2499 821 -2499 0 1
rlabel polysilicon 821 -2505 821 -2505 0 3
rlabel polysilicon 828 -2499 828 -2499 0 1
rlabel polysilicon 828 -2505 828 -2505 0 3
rlabel polysilicon 835 -2499 835 -2499 0 1
rlabel polysilicon 835 -2505 835 -2505 0 3
rlabel polysilicon 842 -2499 842 -2499 0 1
rlabel polysilicon 842 -2505 842 -2505 0 3
rlabel polysilicon 849 -2499 849 -2499 0 1
rlabel polysilicon 849 -2505 849 -2505 0 3
rlabel polysilicon 856 -2499 856 -2499 0 1
rlabel polysilicon 859 -2499 859 -2499 0 2
rlabel polysilicon 856 -2505 856 -2505 0 3
rlabel polysilicon 859 -2505 859 -2505 0 4
rlabel polysilicon 863 -2499 863 -2499 0 1
rlabel polysilicon 863 -2505 863 -2505 0 3
rlabel polysilicon 870 -2499 870 -2499 0 1
rlabel polysilicon 873 -2499 873 -2499 0 2
rlabel polysilicon 873 -2505 873 -2505 0 4
rlabel polysilicon 877 -2499 877 -2499 0 1
rlabel polysilicon 877 -2505 877 -2505 0 3
rlabel polysilicon 884 -2499 884 -2499 0 1
rlabel polysilicon 884 -2505 884 -2505 0 3
rlabel polysilicon 891 -2499 891 -2499 0 1
rlabel polysilicon 891 -2505 891 -2505 0 3
rlabel polysilicon 898 -2499 898 -2499 0 1
rlabel polysilicon 898 -2505 898 -2505 0 3
rlabel polysilicon 905 -2499 905 -2499 0 1
rlabel polysilicon 905 -2505 905 -2505 0 3
rlabel polysilicon 912 -2499 912 -2499 0 1
rlabel polysilicon 912 -2505 912 -2505 0 3
rlabel polysilicon 919 -2499 919 -2499 0 1
rlabel polysilicon 922 -2499 922 -2499 0 2
rlabel polysilicon 919 -2505 919 -2505 0 3
rlabel polysilicon 922 -2505 922 -2505 0 4
rlabel polysilicon 926 -2499 926 -2499 0 1
rlabel polysilicon 926 -2505 926 -2505 0 3
rlabel polysilicon 933 -2499 933 -2499 0 1
rlabel polysilicon 933 -2505 933 -2505 0 3
rlabel polysilicon 940 -2499 940 -2499 0 1
rlabel polysilicon 940 -2505 940 -2505 0 3
rlabel polysilicon 947 -2499 947 -2499 0 1
rlabel polysilicon 947 -2505 947 -2505 0 3
rlabel polysilicon 954 -2499 954 -2499 0 1
rlabel polysilicon 957 -2499 957 -2499 0 2
rlabel polysilicon 954 -2505 954 -2505 0 3
rlabel polysilicon 957 -2505 957 -2505 0 4
rlabel polysilicon 961 -2499 961 -2499 0 1
rlabel polysilicon 961 -2505 961 -2505 0 3
rlabel polysilicon 968 -2499 968 -2499 0 1
rlabel polysilicon 968 -2505 968 -2505 0 3
rlabel polysilicon 975 -2499 975 -2499 0 1
rlabel polysilicon 978 -2499 978 -2499 0 2
rlabel polysilicon 975 -2505 975 -2505 0 3
rlabel polysilicon 978 -2505 978 -2505 0 4
rlabel polysilicon 982 -2499 982 -2499 0 1
rlabel polysilicon 982 -2505 982 -2505 0 3
rlabel polysilicon 992 -2499 992 -2499 0 2
rlabel polysilicon 989 -2505 989 -2505 0 3
rlabel polysilicon 992 -2505 992 -2505 0 4
rlabel polysilicon 996 -2499 996 -2499 0 1
rlabel polysilicon 996 -2505 996 -2505 0 3
rlabel polysilicon 1003 -2499 1003 -2499 0 1
rlabel polysilicon 1003 -2505 1003 -2505 0 3
rlabel polysilicon 1010 -2499 1010 -2499 0 1
rlabel polysilicon 1013 -2499 1013 -2499 0 2
rlabel polysilicon 1010 -2505 1010 -2505 0 3
rlabel polysilicon 1013 -2505 1013 -2505 0 4
rlabel polysilicon 1017 -2499 1017 -2499 0 1
rlabel polysilicon 1017 -2505 1017 -2505 0 3
rlabel polysilicon 1024 -2499 1024 -2499 0 1
rlabel polysilicon 1024 -2505 1024 -2505 0 3
rlabel polysilicon 1031 -2499 1031 -2499 0 1
rlabel polysilicon 1031 -2505 1031 -2505 0 3
rlabel polysilicon 1038 -2499 1038 -2499 0 1
rlabel polysilicon 1038 -2505 1038 -2505 0 3
rlabel polysilicon 1045 -2499 1045 -2499 0 1
rlabel polysilicon 1045 -2505 1045 -2505 0 3
rlabel polysilicon 1052 -2499 1052 -2499 0 1
rlabel polysilicon 1055 -2499 1055 -2499 0 2
rlabel polysilicon 1052 -2505 1052 -2505 0 3
rlabel polysilicon 1055 -2505 1055 -2505 0 4
rlabel polysilicon 1059 -2499 1059 -2499 0 1
rlabel polysilicon 1059 -2505 1059 -2505 0 3
rlabel polysilicon 1066 -2499 1066 -2499 0 1
rlabel polysilicon 1066 -2505 1066 -2505 0 3
rlabel polysilicon 1073 -2499 1073 -2499 0 1
rlabel polysilicon 1076 -2499 1076 -2499 0 2
rlabel polysilicon 1073 -2505 1073 -2505 0 3
rlabel polysilicon 1080 -2499 1080 -2499 0 1
rlabel polysilicon 1083 -2499 1083 -2499 0 2
rlabel polysilicon 1080 -2505 1080 -2505 0 3
rlabel polysilicon 1083 -2505 1083 -2505 0 4
rlabel polysilicon 1087 -2499 1087 -2499 0 1
rlabel polysilicon 1087 -2505 1087 -2505 0 3
rlabel polysilicon 1094 -2499 1094 -2499 0 1
rlabel polysilicon 1094 -2505 1094 -2505 0 3
rlabel polysilicon 1101 -2499 1101 -2499 0 1
rlabel polysilicon 1101 -2505 1101 -2505 0 3
rlabel polysilicon 1108 -2499 1108 -2499 0 1
rlabel polysilicon 1108 -2505 1108 -2505 0 3
rlabel polysilicon 1115 -2499 1115 -2499 0 1
rlabel polysilicon 1115 -2505 1115 -2505 0 3
rlabel polysilicon 1122 -2499 1122 -2499 0 1
rlabel polysilicon 1122 -2505 1122 -2505 0 3
rlabel polysilicon 1129 -2499 1129 -2499 0 1
rlabel polysilicon 1129 -2505 1129 -2505 0 3
rlabel polysilicon 1136 -2499 1136 -2499 0 1
rlabel polysilicon 1136 -2505 1136 -2505 0 3
rlabel polysilicon 1143 -2499 1143 -2499 0 1
rlabel polysilicon 1143 -2505 1143 -2505 0 3
rlabel polysilicon 1150 -2499 1150 -2499 0 1
rlabel polysilicon 1150 -2505 1150 -2505 0 3
rlabel polysilicon 1157 -2499 1157 -2499 0 1
rlabel polysilicon 1157 -2505 1157 -2505 0 3
rlabel polysilicon 1164 -2499 1164 -2499 0 1
rlabel polysilicon 1164 -2505 1164 -2505 0 3
rlabel polysilicon 1171 -2499 1171 -2499 0 1
rlabel polysilicon 1174 -2499 1174 -2499 0 2
rlabel polysilicon 1171 -2505 1171 -2505 0 3
rlabel polysilicon 1174 -2505 1174 -2505 0 4
rlabel polysilicon 1178 -2499 1178 -2499 0 1
rlabel polysilicon 1178 -2505 1178 -2505 0 3
rlabel polysilicon 1185 -2499 1185 -2499 0 1
rlabel polysilicon 1185 -2505 1185 -2505 0 3
rlabel polysilicon 1192 -2499 1192 -2499 0 1
rlabel polysilicon 1192 -2505 1192 -2505 0 3
rlabel polysilicon 1199 -2499 1199 -2499 0 1
rlabel polysilicon 1199 -2505 1199 -2505 0 3
rlabel polysilicon 1206 -2499 1206 -2499 0 1
rlabel polysilicon 1206 -2505 1206 -2505 0 3
rlabel polysilicon 1213 -2499 1213 -2499 0 1
rlabel polysilicon 1213 -2505 1213 -2505 0 3
rlabel polysilicon 1216 -2505 1216 -2505 0 4
rlabel polysilicon 1220 -2499 1220 -2499 0 1
rlabel polysilicon 1220 -2505 1220 -2505 0 3
rlabel polysilicon 1227 -2499 1227 -2499 0 1
rlabel polysilicon 1227 -2505 1227 -2505 0 3
rlabel polysilicon 1234 -2499 1234 -2499 0 1
rlabel polysilicon 1234 -2505 1234 -2505 0 3
rlabel polysilicon 1241 -2499 1241 -2499 0 1
rlabel polysilicon 1241 -2505 1241 -2505 0 3
rlabel polysilicon 1248 -2499 1248 -2499 0 1
rlabel polysilicon 1248 -2505 1248 -2505 0 3
rlabel polysilicon 1255 -2499 1255 -2499 0 1
rlabel polysilicon 1255 -2505 1255 -2505 0 3
rlabel polysilicon 1262 -2499 1262 -2499 0 1
rlabel polysilicon 1262 -2505 1262 -2505 0 3
rlabel polysilicon 1269 -2499 1269 -2499 0 1
rlabel polysilicon 1272 -2499 1272 -2499 0 2
rlabel polysilicon 1269 -2505 1269 -2505 0 3
rlabel polysilicon 1272 -2505 1272 -2505 0 4
rlabel polysilicon 1276 -2499 1276 -2499 0 1
rlabel polysilicon 1276 -2505 1276 -2505 0 3
rlabel polysilicon 1283 -2499 1283 -2499 0 1
rlabel polysilicon 1283 -2505 1283 -2505 0 3
rlabel polysilicon 1290 -2505 1290 -2505 0 3
rlabel polysilicon 1297 -2499 1297 -2499 0 1
rlabel polysilicon 1297 -2505 1297 -2505 0 3
rlabel polysilicon 1304 -2499 1304 -2499 0 1
rlabel polysilicon 1304 -2505 1304 -2505 0 3
rlabel polysilicon 1311 -2499 1311 -2499 0 1
rlabel polysilicon 1311 -2505 1311 -2505 0 3
rlabel polysilicon 1318 -2499 1318 -2499 0 1
rlabel polysilicon 1318 -2505 1318 -2505 0 3
rlabel polysilicon 1325 -2499 1325 -2499 0 1
rlabel polysilicon 1325 -2505 1325 -2505 0 3
rlabel polysilicon 1332 -2499 1332 -2499 0 1
rlabel polysilicon 1335 -2499 1335 -2499 0 2
rlabel polysilicon 1332 -2505 1332 -2505 0 3
rlabel polysilicon 1335 -2505 1335 -2505 0 4
rlabel polysilicon 1339 -2499 1339 -2499 0 1
rlabel polysilicon 1339 -2505 1339 -2505 0 3
rlabel polysilicon 1346 -2499 1346 -2499 0 1
rlabel polysilicon 1346 -2505 1346 -2505 0 3
rlabel polysilicon 1353 -2499 1353 -2499 0 1
rlabel polysilicon 1356 -2499 1356 -2499 0 2
rlabel polysilicon 1353 -2505 1353 -2505 0 3
rlabel polysilicon 1356 -2505 1356 -2505 0 4
rlabel polysilicon 1363 -2499 1363 -2499 0 2
rlabel polysilicon 1360 -2505 1360 -2505 0 3
rlabel polysilicon 1363 -2505 1363 -2505 0 4
rlabel polysilicon 1367 -2499 1367 -2499 0 1
rlabel polysilicon 1367 -2505 1367 -2505 0 3
rlabel polysilicon 1374 -2499 1374 -2499 0 1
rlabel polysilicon 1377 -2499 1377 -2499 0 2
rlabel polysilicon 1374 -2505 1374 -2505 0 3
rlabel polysilicon 1377 -2505 1377 -2505 0 4
rlabel polysilicon 1381 -2499 1381 -2499 0 1
rlabel polysilicon 1381 -2505 1381 -2505 0 3
rlabel polysilicon 1388 -2499 1388 -2499 0 1
rlabel polysilicon 1388 -2505 1388 -2505 0 3
rlabel polysilicon 1395 -2499 1395 -2499 0 1
rlabel polysilicon 1395 -2505 1395 -2505 0 3
rlabel polysilicon 1402 -2499 1402 -2499 0 1
rlabel polysilicon 1402 -2505 1402 -2505 0 3
rlabel polysilicon 1409 -2499 1409 -2499 0 1
rlabel polysilicon 1409 -2505 1409 -2505 0 3
rlabel polysilicon 1416 -2499 1416 -2499 0 1
rlabel polysilicon 1416 -2505 1416 -2505 0 3
rlabel polysilicon 1423 -2499 1423 -2499 0 1
rlabel polysilicon 1423 -2505 1423 -2505 0 3
rlabel polysilicon 1430 -2499 1430 -2499 0 1
rlabel polysilicon 1430 -2505 1430 -2505 0 3
rlabel polysilicon 1437 -2499 1437 -2499 0 1
rlabel polysilicon 1437 -2505 1437 -2505 0 3
rlabel polysilicon 1444 -2499 1444 -2499 0 1
rlabel polysilicon 1444 -2505 1444 -2505 0 3
rlabel polysilicon 1451 -2499 1451 -2499 0 1
rlabel polysilicon 1451 -2505 1451 -2505 0 3
rlabel polysilicon 1458 -2499 1458 -2499 0 1
rlabel polysilicon 1458 -2505 1458 -2505 0 3
rlabel polysilicon 1465 -2499 1465 -2499 0 1
rlabel polysilicon 1465 -2505 1465 -2505 0 3
rlabel polysilicon 1472 -2499 1472 -2499 0 1
rlabel polysilicon 1472 -2505 1472 -2505 0 3
rlabel polysilicon 1479 -2499 1479 -2499 0 1
rlabel polysilicon 1479 -2505 1479 -2505 0 3
rlabel polysilicon 1486 -2499 1486 -2499 0 1
rlabel polysilicon 1486 -2505 1486 -2505 0 3
rlabel polysilicon 1493 -2499 1493 -2499 0 1
rlabel polysilicon 1493 -2505 1493 -2505 0 3
rlabel polysilicon 1500 -2499 1500 -2499 0 1
rlabel polysilicon 1500 -2505 1500 -2505 0 3
rlabel polysilicon 1507 -2499 1507 -2499 0 1
rlabel polysilicon 1507 -2505 1507 -2505 0 3
rlabel polysilicon 1514 -2499 1514 -2499 0 1
rlabel polysilicon 1514 -2505 1514 -2505 0 3
rlabel polysilicon 1521 -2499 1521 -2499 0 1
rlabel polysilicon 1521 -2505 1521 -2505 0 3
rlabel polysilicon 1528 -2499 1528 -2499 0 1
rlabel polysilicon 1528 -2505 1528 -2505 0 3
rlabel polysilicon 1535 -2499 1535 -2499 0 1
rlabel polysilicon 1535 -2505 1535 -2505 0 3
rlabel polysilicon 1542 -2499 1542 -2499 0 1
rlabel polysilicon 1542 -2505 1542 -2505 0 3
rlabel polysilicon 1549 -2499 1549 -2499 0 1
rlabel polysilicon 1549 -2505 1549 -2505 0 3
rlabel polysilicon 1556 -2499 1556 -2499 0 1
rlabel polysilicon 1556 -2505 1556 -2505 0 3
rlabel polysilicon 1563 -2499 1563 -2499 0 1
rlabel polysilicon 1563 -2505 1563 -2505 0 3
rlabel polysilicon 1570 -2499 1570 -2499 0 1
rlabel polysilicon 1570 -2505 1570 -2505 0 3
rlabel polysilicon 1577 -2499 1577 -2499 0 1
rlabel polysilicon 1580 -2499 1580 -2499 0 2
rlabel polysilicon 1577 -2505 1577 -2505 0 3
rlabel polysilicon 1580 -2505 1580 -2505 0 4
rlabel polysilicon 1584 -2499 1584 -2499 0 1
rlabel polysilicon 1584 -2505 1584 -2505 0 3
rlabel polysilicon 1591 -2499 1591 -2499 0 1
rlabel polysilicon 1591 -2505 1591 -2505 0 3
rlabel polysilicon 1598 -2499 1598 -2499 0 1
rlabel polysilicon 1601 -2499 1601 -2499 0 2
rlabel polysilicon 1598 -2505 1598 -2505 0 3
rlabel polysilicon 1601 -2505 1601 -2505 0 4
rlabel polysilicon 1605 -2499 1605 -2499 0 1
rlabel polysilicon 1605 -2505 1605 -2505 0 3
rlabel polysilicon 1612 -2499 1612 -2499 0 1
rlabel polysilicon 1612 -2505 1612 -2505 0 3
rlabel polysilicon 1619 -2499 1619 -2499 0 1
rlabel polysilicon 1619 -2505 1619 -2505 0 3
rlabel polysilicon 1626 -2499 1626 -2499 0 1
rlabel polysilicon 1626 -2505 1626 -2505 0 3
rlabel polysilicon 1633 -2499 1633 -2499 0 1
rlabel polysilicon 1633 -2505 1633 -2505 0 3
rlabel polysilicon 1640 -2499 1640 -2499 0 1
rlabel polysilicon 1640 -2505 1640 -2505 0 3
rlabel polysilicon 1647 -2499 1647 -2499 0 1
rlabel polysilicon 1647 -2505 1647 -2505 0 3
rlabel polysilicon 1654 -2499 1654 -2499 0 1
rlabel polysilicon 1654 -2505 1654 -2505 0 3
rlabel polysilicon 1661 -2499 1661 -2499 0 1
rlabel polysilicon 1661 -2505 1661 -2505 0 3
rlabel polysilicon 1668 -2499 1668 -2499 0 1
rlabel polysilicon 1668 -2505 1668 -2505 0 3
rlabel polysilicon 1678 -2499 1678 -2499 0 2
rlabel polysilicon 1678 -2505 1678 -2505 0 4
rlabel polysilicon 1682 -2499 1682 -2499 0 1
rlabel polysilicon 1682 -2505 1682 -2505 0 3
rlabel polysilicon 1689 -2499 1689 -2499 0 1
rlabel polysilicon 1689 -2505 1689 -2505 0 3
rlabel polysilicon 1696 -2499 1696 -2499 0 1
rlabel polysilicon 1696 -2505 1696 -2505 0 3
rlabel polysilicon 1703 -2499 1703 -2499 0 1
rlabel polysilicon 1703 -2505 1703 -2505 0 3
rlabel polysilicon 1710 -2499 1710 -2499 0 1
rlabel polysilicon 1710 -2505 1710 -2505 0 3
rlabel polysilicon 1717 -2499 1717 -2499 0 1
rlabel polysilicon 1717 -2505 1717 -2505 0 3
rlabel polysilicon 1724 -2499 1724 -2499 0 1
rlabel polysilicon 1724 -2505 1724 -2505 0 3
rlabel polysilicon 1731 -2499 1731 -2499 0 1
rlabel polysilicon 1731 -2505 1731 -2505 0 3
rlabel polysilicon 1738 -2499 1738 -2499 0 1
rlabel polysilicon 1738 -2505 1738 -2505 0 3
rlabel polysilicon 1745 -2499 1745 -2499 0 1
rlabel polysilicon 1745 -2505 1745 -2505 0 3
rlabel polysilicon 1752 -2499 1752 -2499 0 1
rlabel polysilicon 1752 -2505 1752 -2505 0 3
rlabel polysilicon 1759 -2499 1759 -2499 0 1
rlabel polysilicon 1759 -2505 1759 -2505 0 3
rlabel polysilicon 1766 -2499 1766 -2499 0 1
rlabel polysilicon 1766 -2505 1766 -2505 0 3
rlabel polysilicon 1773 -2499 1773 -2499 0 1
rlabel polysilicon 1773 -2505 1773 -2505 0 3
rlabel polysilicon 1780 -2499 1780 -2499 0 1
rlabel polysilicon 1780 -2505 1780 -2505 0 3
rlabel polysilicon 1787 -2499 1787 -2499 0 1
rlabel polysilicon 1787 -2505 1787 -2505 0 3
rlabel polysilicon 1794 -2499 1794 -2499 0 1
rlabel polysilicon 1794 -2505 1794 -2505 0 3
rlabel polysilicon 1801 -2499 1801 -2499 0 1
rlabel polysilicon 1804 -2499 1804 -2499 0 2
rlabel polysilicon 1804 -2505 1804 -2505 0 4
rlabel polysilicon 1808 -2499 1808 -2499 0 1
rlabel polysilicon 1808 -2505 1808 -2505 0 3
rlabel polysilicon 1815 -2499 1815 -2499 0 1
rlabel polysilicon 1815 -2505 1815 -2505 0 3
rlabel polysilicon 1822 -2499 1822 -2499 0 1
rlabel polysilicon 1822 -2505 1822 -2505 0 3
rlabel polysilicon 1829 -2499 1829 -2499 0 1
rlabel polysilicon 1829 -2505 1829 -2505 0 3
rlabel polysilicon 1836 -2499 1836 -2499 0 1
rlabel polysilicon 1836 -2505 1836 -2505 0 3
rlabel polysilicon 1843 -2499 1843 -2499 0 1
rlabel polysilicon 1843 -2505 1843 -2505 0 3
rlabel polysilicon 1850 -2499 1850 -2499 0 1
rlabel polysilicon 1853 -2499 1853 -2499 0 2
rlabel polysilicon 1850 -2505 1850 -2505 0 3
rlabel polysilicon 1857 -2499 1857 -2499 0 1
rlabel polysilicon 1857 -2505 1857 -2505 0 3
rlabel polysilicon 1864 -2499 1864 -2499 0 1
rlabel polysilicon 1864 -2505 1864 -2505 0 3
rlabel polysilicon 1871 -2499 1871 -2499 0 1
rlabel polysilicon 1871 -2505 1871 -2505 0 3
rlabel polysilicon 1878 -2499 1878 -2499 0 1
rlabel polysilicon 1878 -2505 1878 -2505 0 3
rlabel polysilicon 1885 -2499 1885 -2499 0 1
rlabel polysilicon 1885 -2505 1885 -2505 0 3
rlabel polysilicon 1892 -2499 1892 -2499 0 1
rlabel polysilicon 1892 -2505 1892 -2505 0 3
rlabel polysilicon 1899 -2499 1899 -2499 0 1
rlabel polysilicon 1899 -2505 1899 -2505 0 3
rlabel polysilicon 1906 -2499 1906 -2499 0 1
rlabel polysilicon 1906 -2505 1906 -2505 0 3
rlabel polysilicon 1913 -2499 1913 -2499 0 1
rlabel polysilicon 1913 -2505 1913 -2505 0 3
rlabel polysilicon 1920 -2499 1920 -2499 0 1
rlabel polysilicon 1920 -2505 1920 -2505 0 3
rlabel polysilicon 1927 -2499 1927 -2499 0 1
rlabel polysilicon 1927 -2505 1927 -2505 0 3
rlabel polysilicon 1934 -2499 1934 -2499 0 1
rlabel polysilicon 1934 -2505 1934 -2505 0 3
rlabel polysilicon 1941 -2499 1941 -2499 0 1
rlabel polysilicon 1941 -2505 1941 -2505 0 3
rlabel polysilicon 1948 -2499 1948 -2499 0 1
rlabel polysilicon 1948 -2505 1948 -2505 0 3
rlabel polysilicon 1955 -2499 1955 -2499 0 1
rlabel polysilicon 1955 -2505 1955 -2505 0 3
rlabel polysilicon 1962 -2499 1962 -2499 0 1
rlabel polysilicon 1962 -2505 1962 -2505 0 3
rlabel polysilicon 1969 -2499 1969 -2499 0 1
rlabel polysilicon 1969 -2505 1969 -2505 0 3
rlabel polysilicon 1976 -2499 1976 -2499 0 1
rlabel polysilicon 1976 -2505 1976 -2505 0 3
rlabel polysilicon 1983 -2499 1983 -2499 0 1
rlabel polysilicon 1983 -2505 1983 -2505 0 3
rlabel polysilicon 1990 -2499 1990 -2499 0 1
rlabel polysilicon 1990 -2505 1990 -2505 0 3
rlabel polysilicon 1997 -2499 1997 -2499 0 1
rlabel polysilicon 1997 -2505 1997 -2505 0 3
rlabel polysilicon 2004 -2499 2004 -2499 0 1
rlabel polysilicon 2004 -2505 2004 -2505 0 3
rlabel polysilicon 2011 -2499 2011 -2499 0 1
rlabel polysilicon 2011 -2505 2011 -2505 0 3
rlabel polysilicon 2018 -2499 2018 -2499 0 1
rlabel polysilicon 2018 -2505 2018 -2505 0 3
rlabel polysilicon 2025 -2499 2025 -2499 0 1
rlabel polysilicon 2025 -2505 2025 -2505 0 3
rlabel polysilicon 2032 -2499 2032 -2499 0 1
rlabel polysilicon 2032 -2505 2032 -2505 0 3
rlabel polysilicon 2039 -2499 2039 -2499 0 1
rlabel polysilicon 2039 -2505 2039 -2505 0 3
rlabel polysilicon 2046 -2499 2046 -2499 0 1
rlabel polysilicon 2046 -2505 2046 -2505 0 3
rlabel polysilicon 2053 -2499 2053 -2499 0 1
rlabel polysilicon 2053 -2505 2053 -2505 0 3
rlabel polysilicon 2060 -2499 2060 -2499 0 1
rlabel polysilicon 2060 -2505 2060 -2505 0 3
rlabel polysilicon 2067 -2499 2067 -2499 0 1
rlabel polysilicon 2067 -2505 2067 -2505 0 3
rlabel polysilicon 2074 -2499 2074 -2499 0 1
rlabel polysilicon 2074 -2505 2074 -2505 0 3
rlabel polysilicon 2081 -2499 2081 -2499 0 1
rlabel polysilicon 2081 -2505 2081 -2505 0 3
rlabel polysilicon 2088 -2499 2088 -2499 0 1
rlabel polysilicon 2088 -2505 2088 -2505 0 3
rlabel polysilicon 2095 -2499 2095 -2499 0 1
rlabel polysilicon 2095 -2505 2095 -2505 0 3
rlabel polysilicon 2102 -2499 2102 -2499 0 1
rlabel polysilicon 2102 -2505 2102 -2505 0 3
rlabel polysilicon 2109 -2499 2109 -2499 0 1
rlabel polysilicon 2109 -2505 2109 -2505 0 3
rlabel polysilicon 2116 -2499 2116 -2499 0 1
rlabel polysilicon 2116 -2505 2116 -2505 0 3
rlabel polysilicon 2123 -2499 2123 -2499 0 1
rlabel polysilicon 2123 -2505 2123 -2505 0 3
rlabel polysilicon 2130 -2499 2130 -2499 0 1
rlabel polysilicon 2130 -2505 2130 -2505 0 3
rlabel polysilicon 2137 -2499 2137 -2499 0 1
rlabel polysilicon 2137 -2505 2137 -2505 0 3
rlabel polysilicon 2144 -2499 2144 -2499 0 1
rlabel polysilicon 2144 -2505 2144 -2505 0 3
rlabel polysilicon 2151 -2499 2151 -2499 0 1
rlabel polysilicon 2151 -2505 2151 -2505 0 3
rlabel polysilicon 2158 -2499 2158 -2499 0 1
rlabel polysilicon 2158 -2505 2158 -2505 0 3
rlabel polysilicon 2165 -2499 2165 -2499 0 1
rlabel polysilicon 2165 -2505 2165 -2505 0 3
rlabel polysilicon 2172 -2499 2172 -2499 0 1
rlabel polysilicon 2172 -2505 2172 -2505 0 3
rlabel polysilicon 2179 -2499 2179 -2499 0 1
rlabel polysilicon 2179 -2505 2179 -2505 0 3
rlabel polysilicon 2186 -2499 2186 -2499 0 1
rlabel polysilicon 2186 -2505 2186 -2505 0 3
rlabel polysilicon 2193 -2499 2193 -2499 0 1
rlabel polysilicon 2193 -2505 2193 -2505 0 3
rlabel polysilicon 2200 -2499 2200 -2499 0 1
rlabel polysilicon 2200 -2505 2200 -2505 0 3
rlabel polysilicon 2207 -2499 2207 -2499 0 1
rlabel polysilicon 2207 -2505 2207 -2505 0 3
rlabel polysilicon 2214 -2499 2214 -2499 0 1
rlabel polysilicon 2214 -2505 2214 -2505 0 3
rlabel polysilicon 2221 -2499 2221 -2499 0 1
rlabel polysilicon 2221 -2505 2221 -2505 0 3
rlabel polysilicon 2228 -2499 2228 -2499 0 1
rlabel polysilicon 2228 -2505 2228 -2505 0 3
rlabel polysilicon 2235 -2499 2235 -2499 0 1
rlabel polysilicon 2235 -2505 2235 -2505 0 3
rlabel polysilicon 2242 -2499 2242 -2499 0 1
rlabel polysilicon 2242 -2505 2242 -2505 0 3
rlabel polysilicon 2249 -2499 2249 -2499 0 1
rlabel polysilicon 2249 -2505 2249 -2505 0 3
rlabel polysilicon 2256 -2499 2256 -2499 0 1
rlabel polysilicon 2256 -2505 2256 -2505 0 3
rlabel polysilicon 2263 -2499 2263 -2499 0 1
rlabel polysilicon 2263 -2505 2263 -2505 0 3
rlabel polysilicon 2270 -2499 2270 -2499 0 1
rlabel polysilicon 2270 -2505 2270 -2505 0 3
rlabel polysilicon 2280 -2499 2280 -2499 0 2
rlabel polysilicon 2280 -2505 2280 -2505 0 4
rlabel polysilicon 2284 -2499 2284 -2499 0 1
rlabel polysilicon 2284 -2505 2284 -2505 0 3
rlabel polysilicon 2291 -2499 2291 -2499 0 1
rlabel polysilicon 2291 -2505 2291 -2505 0 3
rlabel polysilicon 2298 -2499 2298 -2499 0 1
rlabel polysilicon 2298 -2505 2298 -2505 0 3
rlabel polysilicon 2305 -2499 2305 -2499 0 1
rlabel polysilicon 2305 -2505 2305 -2505 0 3
rlabel polysilicon 2312 -2499 2312 -2499 0 1
rlabel polysilicon 2312 -2505 2312 -2505 0 3
rlabel polysilicon 9 -2672 9 -2672 0 1
rlabel polysilicon 9 -2678 9 -2678 0 3
rlabel polysilicon 16 -2672 16 -2672 0 1
rlabel polysilicon 16 -2678 16 -2678 0 3
rlabel polysilicon 26 -2672 26 -2672 0 2
rlabel polysilicon 23 -2678 23 -2678 0 3
rlabel polysilicon 26 -2678 26 -2678 0 4
rlabel polysilicon 30 -2672 30 -2672 0 1
rlabel polysilicon 30 -2678 30 -2678 0 3
rlabel polysilicon 37 -2672 37 -2672 0 1
rlabel polysilicon 37 -2678 37 -2678 0 3
rlabel polysilicon 44 -2672 44 -2672 0 1
rlabel polysilicon 44 -2678 44 -2678 0 3
rlabel polysilicon 51 -2672 51 -2672 0 1
rlabel polysilicon 54 -2672 54 -2672 0 2
rlabel polysilicon 51 -2678 51 -2678 0 3
rlabel polysilicon 54 -2678 54 -2678 0 4
rlabel polysilicon 58 -2672 58 -2672 0 1
rlabel polysilicon 58 -2678 58 -2678 0 3
rlabel polysilicon 65 -2672 65 -2672 0 1
rlabel polysilicon 68 -2672 68 -2672 0 2
rlabel polysilicon 65 -2678 65 -2678 0 3
rlabel polysilicon 68 -2678 68 -2678 0 4
rlabel polysilicon 72 -2672 72 -2672 0 1
rlabel polysilicon 75 -2672 75 -2672 0 2
rlabel polysilicon 72 -2678 72 -2678 0 3
rlabel polysilicon 75 -2678 75 -2678 0 4
rlabel polysilicon 79 -2672 79 -2672 0 1
rlabel polysilicon 79 -2678 79 -2678 0 3
rlabel polysilicon 86 -2672 86 -2672 0 1
rlabel polysilicon 86 -2678 86 -2678 0 3
rlabel polysilicon 93 -2672 93 -2672 0 1
rlabel polysilicon 93 -2678 93 -2678 0 3
rlabel polysilicon 100 -2672 100 -2672 0 1
rlabel polysilicon 103 -2672 103 -2672 0 2
rlabel polysilicon 100 -2678 100 -2678 0 3
rlabel polysilicon 103 -2678 103 -2678 0 4
rlabel polysilicon 107 -2672 107 -2672 0 1
rlabel polysilicon 107 -2678 107 -2678 0 3
rlabel polysilicon 114 -2672 114 -2672 0 1
rlabel polysilicon 114 -2678 114 -2678 0 3
rlabel polysilicon 121 -2672 121 -2672 0 1
rlabel polysilicon 121 -2678 121 -2678 0 3
rlabel polysilicon 128 -2672 128 -2672 0 1
rlabel polysilicon 131 -2672 131 -2672 0 2
rlabel polysilicon 128 -2678 128 -2678 0 3
rlabel polysilicon 131 -2678 131 -2678 0 4
rlabel polysilicon 135 -2672 135 -2672 0 1
rlabel polysilicon 135 -2678 135 -2678 0 3
rlabel polysilicon 142 -2672 142 -2672 0 1
rlabel polysilicon 142 -2678 142 -2678 0 3
rlabel polysilicon 149 -2672 149 -2672 0 1
rlabel polysilicon 149 -2678 149 -2678 0 3
rlabel polysilicon 156 -2672 156 -2672 0 1
rlabel polysilicon 156 -2678 156 -2678 0 3
rlabel polysilicon 163 -2672 163 -2672 0 1
rlabel polysilicon 163 -2678 163 -2678 0 3
rlabel polysilicon 170 -2672 170 -2672 0 1
rlabel polysilicon 170 -2678 170 -2678 0 3
rlabel polysilicon 177 -2672 177 -2672 0 1
rlabel polysilicon 177 -2678 177 -2678 0 3
rlabel polysilicon 184 -2672 184 -2672 0 1
rlabel polysilicon 184 -2678 184 -2678 0 3
rlabel polysilicon 191 -2672 191 -2672 0 1
rlabel polysilicon 191 -2678 191 -2678 0 3
rlabel polysilicon 198 -2672 198 -2672 0 1
rlabel polysilicon 201 -2672 201 -2672 0 2
rlabel polysilicon 198 -2678 198 -2678 0 3
rlabel polysilicon 205 -2672 205 -2672 0 1
rlabel polysilicon 205 -2678 205 -2678 0 3
rlabel polysilicon 212 -2672 212 -2672 0 1
rlabel polysilicon 212 -2678 212 -2678 0 3
rlabel polysilicon 219 -2672 219 -2672 0 1
rlabel polysilicon 219 -2678 219 -2678 0 3
rlabel polysilicon 226 -2672 226 -2672 0 1
rlabel polysilicon 226 -2678 226 -2678 0 3
rlabel polysilicon 233 -2672 233 -2672 0 1
rlabel polysilicon 233 -2678 233 -2678 0 3
rlabel polysilicon 240 -2672 240 -2672 0 1
rlabel polysilicon 240 -2678 240 -2678 0 3
rlabel polysilicon 243 -2678 243 -2678 0 4
rlabel polysilicon 247 -2672 247 -2672 0 1
rlabel polysilicon 247 -2678 247 -2678 0 3
rlabel polysilicon 254 -2672 254 -2672 0 1
rlabel polysilicon 254 -2678 254 -2678 0 3
rlabel polysilicon 261 -2672 261 -2672 0 1
rlabel polysilicon 261 -2678 261 -2678 0 3
rlabel polysilicon 268 -2672 268 -2672 0 1
rlabel polysilicon 268 -2678 268 -2678 0 3
rlabel polysilicon 275 -2672 275 -2672 0 1
rlabel polysilicon 275 -2678 275 -2678 0 3
rlabel polysilicon 282 -2672 282 -2672 0 1
rlabel polysilicon 282 -2678 282 -2678 0 3
rlabel polysilicon 289 -2672 289 -2672 0 1
rlabel polysilicon 289 -2678 289 -2678 0 3
rlabel polysilicon 296 -2672 296 -2672 0 1
rlabel polysilicon 296 -2678 296 -2678 0 3
rlabel polysilicon 303 -2672 303 -2672 0 1
rlabel polysilicon 303 -2678 303 -2678 0 3
rlabel polysilicon 310 -2672 310 -2672 0 1
rlabel polysilicon 310 -2678 310 -2678 0 3
rlabel polysilicon 317 -2672 317 -2672 0 1
rlabel polysilicon 317 -2678 317 -2678 0 3
rlabel polysilicon 324 -2672 324 -2672 0 1
rlabel polysilicon 324 -2678 324 -2678 0 3
rlabel polysilicon 331 -2672 331 -2672 0 1
rlabel polysilicon 331 -2678 331 -2678 0 3
rlabel polysilicon 338 -2672 338 -2672 0 1
rlabel polysilicon 338 -2678 338 -2678 0 3
rlabel polysilicon 345 -2672 345 -2672 0 1
rlabel polysilicon 345 -2678 345 -2678 0 3
rlabel polysilicon 352 -2672 352 -2672 0 1
rlabel polysilicon 352 -2678 352 -2678 0 3
rlabel polysilicon 359 -2672 359 -2672 0 1
rlabel polysilicon 359 -2678 359 -2678 0 3
rlabel polysilicon 366 -2672 366 -2672 0 1
rlabel polysilicon 366 -2678 366 -2678 0 3
rlabel polysilicon 373 -2672 373 -2672 0 1
rlabel polysilicon 373 -2678 373 -2678 0 3
rlabel polysilicon 380 -2672 380 -2672 0 1
rlabel polysilicon 380 -2678 380 -2678 0 3
rlabel polysilicon 387 -2672 387 -2672 0 1
rlabel polysilicon 387 -2678 387 -2678 0 3
rlabel polysilicon 394 -2672 394 -2672 0 1
rlabel polysilicon 394 -2678 394 -2678 0 3
rlabel polysilicon 401 -2672 401 -2672 0 1
rlabel polysilicon 401 -2678 401 -2678 0 3
rlabel polysilicon 408 -2672 408 -2672 0 1
rlabel polysilicon 411 -2672 411 -2672 0 2
rlabel polysilicon 408 -2678 408 -2678 0 3
rlabel polysilicon 411 -2678 411 -2678 0 4
rlabel polysilicon 415 -2672 415 -2672 0 1
rlabel polysilicon 415 -2678 415 -2678 0 3
rlabel polysilicon 422 -2672 422 -2672 0 1
rlabel polysilicon 422 -2678 422 -2678 0 3
rlabel polysilicon 429 -2672 429 -2672 0 1
rlabel polysilicon 429 -2678 429 -2678 0 3
rlabel polysilicon 436 -2672 436 -2672 0 1
rlabel polysilicon 436 -2678 436 -2678 0 3
rlabel polysilicon 443 -2672 443 -2672 0 1
rlabel polysilicon 443 -2678 443 -2678 0 3
rlabel polysilicon 450 -2672 450 -2672 0 1
rlabel polysilicon 450 -2678 450 -2678 0 3
rlabel polysilicon 457 -2672 457 -2672 0 1
rlabel polysilicon 457 -2678 457 -2678 0 3
rlabel polysilicon 464 -2672 464 -2672 0 1
rlabel polysilicon 464 -2678 464 -2678 0 3
rlabel polysilicon 471 -2672 471 -2672 0 1
rlabel polysilicon 471 -2678 471 -2678 0 3
rlabel polysilicon 478 -2672 478 -2672 0 1
rlabel polysilicon 478 -2678 478 -2678 0 3
rlabel polysilicon 485 -2672 485 -2672 0 1
rlabel polysilicon 485 -2678 485 -2678 0 3
rlabel polysilicon 492 -2672 492 -2672 0 1
rlabel polysilicon 492 -2678 492 -2678 0 3
rlabel polysilicon 499 -2672 499 -2672 0 1
rlabel polysilicon 499 -2678 499 -2678 0 3
rlabel polysilicon 506 -2672 506 -2672 0 1
rlabel polysilicon 506 -2678 506 -2678 0 3
rlabel polysilicon 513 -2672 513 -2672 0 1
rlabel polysilicon 513 -2678 513 -2678 0 3
rlabel polysilicon 520 -2672 520 -2672 0 1
rlabel polysilicon 520 -2678 520 -2678 0 3
rlabel polysilicon 527 -2672 527 -2672 0 1
rlabel polysilicon 527 -2678 527 -2678 0 3
rlabel polysilicon 534 -2672 534 -2672 0 1
rlabel polysilicon 534 -2678 534 -2678 0 3
rlabel polysilicon 541 -2672 541 -2672 0 1
rlabel polysilicon 541 -2678 541 -2678 0 3
rlabel polysilicon 548 -2672 548 -2672 0 1
rlabel polysilicon 548 -2678 548 -2678 0 3
rlabel polysilicon 555 -2672 555 -2672 0 1
rlabel polysilicon 558 -2672 558 -2672 0 2
rlabel polysilicon 555 -2678 555 -2678 0 3
rlabel polysilicon 558 -2678 558 -2678 0 4
rlabel polysilicon 562 -2672 562 -2672 0 1
rlabel polysilicon 562 -2678 562 -2678 0 3
rlabel polysilicon 569 -2672 569 -2672 0 1
rlabel polysilicon 569 -2678 569 -2678 0 3
rlabel polysilicon 576 -2672 576 -2672 0 1
rlabel polysilicon 576 -2678 576 -2678 0 3
rlabel polysilicon 583 -2672 583 -2672 0 1
rlabel polysilicon 583 -2678 583 -2678 0 3
rlabel polysilicon 590 -2672 590 -2672 0 1
rlabel polysilicon 590 -2678 590 -2678 0 3
rlabel polysilicon 597 -2672 597 -2672 0 1
rlabel polysilicon 597 -2678 597 -2678 0 3
rlabel polysilicon 604 -2672 604 -2672 0 1
rlabel polysilicon 604 -2678 604 -2678 0 3
rlabel polysilicon 611 -2672 611 -2672 0 1
rlabel polysilicon 611 -2678 611 -2678 0 3
rlabel polysilicon 618 -2672 618 -2672 0 1
rlabel polysilicon 618 -2678 618 -2678 0 3
rlabel polysilicon 625 -2672 625 -2672 0 1
rlabel polysilicon 625 -2678 625 -2678 0 3
rlabel polysilicon 632 -2672 632 -2672 0 1
rlabel polysilicon 632 -2678 632 -2678 0 3
rlabel polysilicon 639 -2672 639 -2672 0 1
rlabel polysilicon 639 -2678 639 -2678 0 3
rlabel polysilicon 646 -2672 646 -2672 0 1
rlabel polysilicon 646 -2678 646 -2678 0 3
rlabel polysilicon 653 -2672 653 -2672 0 1
rlabel polysilicon 653 -2678 653 -2678 0 3
rlabel polysilicon 660 -2672 660 -2672 0 1
rlabel polysilicon 660 -2678 660 -2678 0 3
rlabel polysilicon 667 -2672 667 -2672 0 1
rlabel polysilicon 667 -2678 667 -2678 0 3
rlabel polysilicon 674 -2672 674 -2672 0 1
rlabel polysilicon 674 -2678 674 -2678 0 3
rlabel polysilicon 681 -2672 681 -2672 0 1
rlabel polysilicon 681 -2678 681 -2678 0 3
rlabel polysilicon 688 -2672 688 -2672 0 1
rlabel polysilicon 688 -2678 688 -2678 0 3
rlabel polysilicon 695 -2672 695 -2672 0 1
rlabel polysilicon 695 -2678 695 -2678 0 3
rlabel polysilicon 702 -2672 702 -2672 0 1
rlabel polysilicon 702 -2678 702 -2678 0 3
rlabel polysilicon 709 -2672 709 -2672 0 1
rlabel polysilicon 709 -2678 709 -2678 0 3
rlabel polysilicon 716 -2672 716 -2672 0 1
rlabel polysilicon 716 -2678 716 -2678 0 3
rlabel polysilicon 726 -2672 726 -2672 0 2
rlabel polysilicon 726 -2678 726 -2678 0 4
rlabel polysilicon 730 -2672 730 -2672 0 1
rlabel polysilicon 730 -2678 730 -2678 0 3
rlabel polysilicon 737 -2672 737 -2672 0 1
rlabel polysilicon 737 -2678 737 -2678 0 3
rlabel polysilicon 744 -2672 744 -2672 0 1
rlabel polysilicon 744 -2678 744 -2678 0 3
rlabel polysilicon 751 -2672 751 -2672 0 1
rlabel polysilicon 751 -2678 751 -2678 0 3
rlabel polysilicon 758 -2672 758 -2672 0 1
rlabel polysilicon 758 -2678 758 -2678 0 3
rlabel polysilicon 765 -2672 765 -2672 0 1
rlabel polysilicon 765 -2678 765 -2678 0 3
rlabel polysilicon 772 -2672 772 -2672 0 1
rlabel polysilicon 772 -2678 772 -2678 0 3
rlabel polysilicon 779 -2672 779 -2672 0 1
rlabel polysilicon 779 -2678 779 -2678 0 3
rlabel polysilicon 786 -2672 786 -2672 0 1
rlabel polysilicon 789 -2672 789 -2672 0 2
rlabel polysilicon 786 -2678 786 -2678 0 3
rlabel polysilicon 789 -2678 789 -2678 0 4
rlabel polysilicon 793 -2672 793 -2672 0 1
rlabel polysilicon 793 -2678 793 -2678 0 3
rlabel polysilicon 800 -2672 800 -2672 0 1
rlabel polysilicon 800 -2678 800 -2678 0 3
rlabel polysilicon 810 -2672 810 -2672 0 2
rlabel polysilicon 807 -2678 807 -2678 0 3
rlabel polysilicon 810 -2678 810 -2678 0 4
rlabel polysilicon 814 -2672 814 -2672 0 1
rlabel polysilicon 817 -2672 817 -2672 0 2
rlabel polysilicon 814 -2678 814 -2678 0 3
rlabel polysilicon 817 -2678 817 -2678 0 4
rlabel polysilicon 821 -2672 821 -2672 0 1
rlabel polysilicon 824 -2672 824 -2672 0 2
rlabel polysilicon 821 -2678 821 -2678 0 3
rlabel polysilicon 824 -2678 824 -2678 0 4
rlabel polysilicon 828 -2672 828 -2672 0 1
rlabel polysilicon 828 -2678 828 -2678 0 3
rlabel polysilicon 835 -2672 835 -2672 0 1
rlabel polysilicon 835 -2678 835 -2678 0 3
rlabel polysilicon 842 -2672 842 -2672 0 1
rlabel polysilicon 842 -2678 842 -2678 0 3
rlabel polysilicon 849 -2672 849 -2672 0 1
rlabel polysilicon 849 -2678 849 -2678 0 3
rlabel polysilicon 856 -2672 856 -2672 0 1
rlabel polysilicon 856 -2678 856 -2678 0 3
rlabel polysilicon 863 -2672 863 -2672 0 1
rlabel polysilicon 863 -2678 863 -2678 0 3
rlabel polysilicon 870 -2672 870 -2672 0 1
rlabel polysilicon 870 -2678 870 -2678 0 3
rlabel polysilicon 877 -2672 877 -2672 0 1
rlabel polysilicon 877 -2678 877 -2678 0 3
rlabel polysilicon 884 -2672 884 -2672 0 1
rlabel polysilicon 884 -2678 884 -2678 0 3
rlabel polysilicon 891 -2672 891 -2672 0 1
rlabel polysilicon 894 -2672 894 -2672 0 2
rlabel polysilicon 894 -2678 894 -2678 0 4
rlabel polysilicon 898 -2672 898 -2672 0 1
rlabel polysilicon 898 -2678 898 -2678 0 3
rlabel polysilicon 905 -2672 905 -2672 0 1
rlabel polysilicon 905 -2678 905 -2678 0 3
rlabel polysilicon 912 -2672 912 -2672 0 1
rlabel polysilicon 912 -2678 912 -2678 0 3
rlabel polysilicon 919 -2678 919 -2678 0 3
rlabel polysilicon 922 -2678 922 -2678 0 4
rlabel polysilicon 926 -2672 926 -2672 0 1
rlabel polysilicon 926 -2678 926 -2678 0 3
rlabel polysilicon 933 -2672 933 -2672 0 1
rlabel polysilicon 933 -2678 933 -2678 0 3
rlabel polysilicon 940 -2672 940 -2672 0 1
rlabel polysilicon 940 -2678 940 -2678 0 3
rlabel polysilicon 947 -2672 947 -2672 0 1
rlabel polysilicon 950 -2672 950 -2672 0 2
rlabel polysilicon 947 -2678 947 -2678 0 3
rlabel polysilicon 950 -2678 950 -2678 0 4
rlabel polysilicon 954 -2672 954 -2672 0 1
rlabel polysilicon 954 -2678 954 -2678 0 3
rlabel polysilicon 957 -2678 957 -2678 0 4
rlabel polysilicon 961 -2672 961 -2672 0 1
rlabel polysilicon 961 -2678 961 -2678 0 3
rlabel polysilicon 968 -2672 968 -2672 0 1
rlabel polysilicon 968 -2678 968 -2678 0 3
rlabel polysilicon 975 -2672 975 -2672 0 1
rlabel polysilicon 975 -2678 975 -2678 0 3
rlabel polysilicon 982 -2672 982 -2672 0 1
rlabel polysilicon 982 -2678 982 -2678 0 3
rlabel polysilicon 989 -2672 989 -2672 0 1
rlabel polysilicon 989 -2678 989 -2678 0 3
rlabel polysilicon 996 -2672 996 -2672 0 1
rlabel polysilicon 996 -2678 996 -2678 0 3
rlabel polysilicon 1003 -2672 1003 -2672 0 1
rlabel polysilicon 1006 -2672 1006 -2672 0 2
rlabel polysilicon 1003 -2678 1003 -2678 0 3
rlabel polysilicon 1010 -2672 1010 -2672 0 1
rlabel polysilicon 1013 -2672 1013 -2672 0 2
rlabel polysilicon 1010 -2678 1010 -2678 0 3
rlabel polysilicon 1013 -2678 1013 -2678 0 4
rlabel polysilicon 1017 -2672 1017 -2672 0 1
rlabel polysilicon 1017 -2678 1017 -2678 0 3
rlabel polysilicon 1024 -2672 1024 -2672 0 1
rlabel polysilicon 1024 -2678 1024 -2678 0 3
rlabel polysilicon 1031 -2672 1031 -2672 0 1
rlabel polysilicon 1031 -2678 1031 -2678 0 3
rlabel polysilicon 1038 -2672 1038 -2672 0 1
rlabel polysilicon 1038 -2678 1038 -2678 0 3
rlabel polysilicon 1041 -2678 1041 -2678 0 4
rlabel polysilicon 1045 -2672 1045 -2672 0 1
rlabel polysilicon 1045 -2678 1045 -2678 0 3
rlabel polysilicon 1052 -2672 1052 -2672 0 1
rlabel polysilicon 1052 -2678 1052 -2678 0 3
rlabel polysilicon 1059 -2672 1059 -2672 0 1
rlabel polysilicon 1059 -2678 1059 -2678 0 3
rlabel polysilicon 1066 -2672 1066 -2672 0 1
rlabel polysilicon 1066 -2678 1066 -2678 0 3
rlabel polysilicon 1073 -2672 1073 -2672 0 1
rlabel polysilicon 1073 -2678 1073 -2678 0 3
rlabel polysilicon 1080 -2672 1080 -2672 0 1
rlabel polysilicon 1080 -2678 1080 -2678 0 3
rlabel polysilicon 1087 -2672 1087 -2672 0 1
rlabel polysilicon 1087 -2678 1087 -2678 0 3
rlabel polysilicon 1094 -2672 1094 -2672 0 1
rlabel polysilicon 1094 -2678 1094 -2678 0 3
rlabel polysilicon 1101 -2672 1101 -2672 0 1
rlabel polysilicon 1101 -2678 1101 -2678 0 3
rlabel polysilicon 1108 -2672 1108 -2672 0 1
rlabel polysilicon 1108 -2678 1108 -2678 0 3
rlabel polysilicon 1115 -2672 1115 -2672 0 1
rlabel polysilicon 1115 -2678 1115 -2678 0 3
rlabel polysilicon 1122 -2672 1122 -2672 0 1
rlabel polysilicon 1125 -2672 1125 -2672 0 2
rlabel polysilicon 1122 -2678 1122 -2678 0 3
rlabel polysilicon 1125 -2678 1125 -2678 0 4
rlabel polysilicon 1129 -2672 1129 -2672 0 1
rlabel polysilicon 1129 -2678 1129 -2678 0 3
rlabel polysilicon 1136 -2672 1136 -2672 0 1
rlabel polysilicon 1139 -2678 1139 -2678 0 4
rlabel polysilicon 1143 -2672 1143 -2672 0 1
rlabel polysilicon 1143 -2678 1143 -2678 0 3
rlabel polysilicon 1150 -2672 1150 -2672 0 1
rlabel polysilicon 1150 -2678 1150 -2678 0 3
rlabel polysilicon 1157 -2672 1157 -2672 0 1
rlabel polysilicon 1157 -2678 1157 -2678 0 3
rlabel polysilicon 1164 -2672 1164 -2672 0 1
rlabel polysilicon 1164 -2678 1164 -2678 0 3
rlabel polysilicon 1171 -2672 1171 -2672 0 1
rlabel polysilicon 1171 -2678 1171 -2678 0 3
rlabel polysilicon 1178 -2672 1178 -2672 0 1
rlabel polysilicon 1178 -2678 1178 -2678 0 3
rlabel polysilicon 1185 -2672 1185 -2672 0 1
rlabel polysilicon 1188 -2672 1188 -2672 0 2
rlabel polysilicon 1185 -2678 1185 -2678 0 3
rlabel polysilicon 1192 -2672 1192 -2672 0 1
rlabel polysilicon 1195 -2672 1195 -2672 0 2
rlabel polysilicon 1192 -2678 1192 -2678 0 3
rlabel polysilicon 1195 -2678 1195 -2678 0 4
rlabel polysilicon 1199 -2672 1199 -2672 0 1
rlabel polysilicon 1199 -2678 1199 -2678 0 3
rlabel polysilicon 1206 -2672 1206 -2672 0 1
rlabel polysilicon 1206 -2678 1206 -2678 0 3
rlabel polysilicon 1213 -2672 1213 -2672 0 1
rlabel polysilicon 1213 -2678 1213 -2678 0 3
rlabel polysilicon 1220 -2672 1220 -2672 0 1
rlabel polysilicon 1220 -2678 1220 -2678 0 3
rlabel polysilicon 1227 -2672 1227 -2672 0 1
rlabel polysilicon 1227 -2678 1227 -2678 0 3
rlabel polysilicon 1234 -2672 1234 -2672 0 1
rlabel polysilicon 1237 -2672 1237 -2672 0 2
rlabel polysilicon 1234 -2678 1234 -2678 0 3
rlabel polysilicon 1241 -2672 1241 -2672 0 1
rlabel polysilicon 1241 -2678 1241 -2678 0 3
rlabel polysilicon 1244 -2678 1244 -2678 0 4
rlabel polysilicon 1248 -2672 1248 -2672 0 1
rlabel polysilicon 1248 -2678 1248 -2678 0 3
rlabel polysilicon 1255 -2672 1255 -2672 0 1
rlabel polysilicon 1255 -2678 1255 -2678 0 3
rlabel polysilicon 1262 -2672 1262 -2672 0 1
rlabel polysilicon 1262 -2678 1262 -2678 0 3
rlabel polysilicon 1269 -2672 1269 -2672 0 1
rlabel polysilicon 1269 -2678 1269 -2678 0 3
rlabel polysilicon 1276 -2672 1276 -2672 0 1
rlabel polysilicon 1276 -2678 1276 -2678 0 3
rlabel polysilicon 1283 -2672 1283 -2672 0 1
rlabel polysilicon 1283 -2678 1283 -2678 0 3
rlabel polysilicon 1290 -2672 1290 -2672 0 1
rlabel polysilicon 1290 -2678 1290 -2678 0 3
rlabel polysilicon 1297 -2672 1297 -2672 0 1
rlabel polysilicon 1297 -2678 1297 -2678 0 3
rlabel polysilicon 1304 -2672 1304 -2672 0 1
rlabel polysilicon 1304 -2678 1304 -2678 0 3
rlabel polysilicon 1311 -2672 1311 -2672 0 1
rlabel polysilicon 1314 -2672 1314 -2672 0 2
rlabel polysilicon 1311 -2678 1311 -2678 0 3
rlabel polysilicon 1314 -2678 1314 -2678 0 4
rlabel polysilicon 1318 -2672 1318 -2672 0 1
rlabel polysilicon 1318 -2678 1318 -2678 0 3
rlabel polysilicon 1325 -2678 1325 -2678 0 3
rlabel polysilicon 1328 -2678 1328 -2678 0 4
rlabel polysilicon 1332 -2672 1332 -2672 0 1
rlabel polysilicon 1332 -2678 1332 -2678 0 3
rlabel polysilicon 1339 -2672 1339 -2672 0 1
rlabel polysilicon 1339 -2678 1339 -2678 0 3
rlabel polysilicon 1346 -2672 1346 -2672 0 1
rlabel polysilicon 1346 -2678 1346 -2678 0 3
rlabel polysilicon 1353 -2672 1353 -2672 0 1
rlabel polysilicon 1353 -2678 1353 -2678 0 3
rlabel polysilicon 1360 -2672 1360 -2672 0 1
rlabel polysilicon 1360 -2678 1360 -2678 0 3
rlabel polysilicon 1367 -2672 1367 -2672 0 1
rlabel polysilicon 1367 -2678 1367 -2678 0 3
rlabel polysilicon 1374 -2672 1374 -2672 0 1
rlabel polysilicon 1374 -2678 1374 -2678 0 3
rlabel polysilicon 1381 -2672 1381 -2672 0 1
rlabel polysilicon 1381 -2678 1381 -2678 0 3
rlabel polysilicon 1388 -2672 1388 -2672 0 1
rlabel polysilicon 1388 -2678 1388 -2678 0 3
rlabel polysilicon 1395 -2672 1395 -2672 0 1
rlabel polysilicon 1398 -2672 1398 -2672 0 2
rlabel polysilicon 1395 -2678 1395 -2678 0 3
rlabel polysilicon 1398 -2678 1398 -2678 0 4
rlabel polysilicon 1402 -2672 1402 -2672 0 1
rlabel polysilicon 1402 -2678 1402 -2678 0 3
rlabel polysilicon 1409 -2672 1409 -2672 0 1
rlabel polysilicon 1412 -2672 1412 -2672 0 2
rlabel polysilicon 1409 -2678 1409 -2678 0 3
rlabel polysilicon 1416 -2672 1416 -2672 0 1
rlabel polysilicon 1416 -2678 1416 -2678 0 3
rlabel polysilicon 1423 -2672 1423 -2672 0 1
rlabel polysilicon 1423 -2678 1423 -2678 0 3
rlabel polysilicon 1430 -2672 1430 -2672 0 1
rlabel polysilicon 1430 -2678 1430 -2678 0 3
rlabel polysilicon 1433 -2678 1433 -2678 0 4
rlabel polysilicon 1437 -2672 1437 -2672 0 1
rlabel polysilicon 1440 -2672 1440 -2672 0 2
rlabel polysilicon 1437 -2678 1437 -2678 0 3
rlabel polysilicon 1440 -2678 1440 -2678 0 4
rlabel polysilicon 1444 -2672 1444 -2672 0 1
rlabel polysilicon 1447 -2672 1447 -2672 0 2
rlabel polysilicon 1444 -2678 1444 -2678 0 3
rlabel polysilicon 1451 -2672 1451 -2672 0 1
rlabel polysilicon 1451 -2678 1451 -2678 0 3
rlabel polysilicon 1458 -2672 1458 -2672 0 1
rlabel polysilicon 1458 -2678 1458 -2678 0 3
rlabel polysilicon 1465 -2672 1465 -2672 0 1
rlabel polysilicon 1465 -2678 1465 -2678 0 3
rlabel polysilicon 1472 -2672 1472 -2672 0 1
rlabel polysilicon 1472 -2678 1472 -2678 0 3
rlabel polysilicon 1479 -2672 1479 -2672 0 1
rlabel polysilicon 1479 -2678 1479 -2678 0 3
rlabel polysilicon 1486 -2672 1486 -2672 0 1
rlabel polysilicon 1486 -2678 1486 -2678 0 3
rlabel polysilicon 1493 -2672 1493 -2672 0 1
rlabel polysilicon 1493 -2678 1493 -2678 0 3
rlabel polysilicon 1500 -2672 1500 -2672 0 1
rlabel polysilicon 1500 -2678 1500 -2678 0 3
rlabel polysilicon 1507 -2672 1507 -2672 0 1
rlabel polysilicon 1510 -2672 1510 -2672 0 2
rlabel polysilicon 1507 -2678 1507 -2678 0 3
rlabel polysilicon 1510 -2678 1510 -2678 0 4
rlabel polysilicon 1514 -2672 1514 -2672 0 1
rlabel polysilicon 1514 -2678 1514 -2678 0 3
rlabel polysilicon 1521 -2672 1521 -2672 0 1
rlabel polysilicon 1521 -2678 1521 -2678 0 3
rlabel polysilicon 1528 -2672 1528 -2672 0 1
rlabel polysilicon 1528 -2678 1528 -2678 0 3
rlabel polysilicon 1535 -2672 1535 -2672 0 1
rlabel polysilicon 1535 -2678 1535 -2678 0 3
rlabel polysilicon 1542 -2672 1542 -2672 0 1
rlabel polysilicon 1542 -2678 1542 -2678 0 3
rlabel polysilicon 1549 -2672 1549 -2672 0 1
rlabel polysilicon 1549 -2678 1549 -2678 0 3
rlabel polysilicon 1556 -2672 1556 -2672 0 1
rlabel polysilicon 1556 -2678 1556 -2678 0 3
rlabel polysilicon 1563 -2672 1563 -2672 0 1
rlabel polysilicon 1563 -2678 1563 -2678 0 3
rlabel polysilicon 1570 -2672 1570 -2672 0 1
rlabel polysilicon 1570 -2678 1570 -2678 0 3
rlabel polysilicon 1577 -2672 1577 -2672 0 1
rlabel polysilicon 1580 -2672 1580 -2672 0 2
rlabel polysilicon 1577 -2678 1577 -2678 0 3
rlabel polysilicon 1580 -2678 1580 -2678 0 4
rlabel polysilicon 1584 -2672 1584 -2672 0 1
rlabel polysilicon 1584 -2678 1584 -2678 0 3
rlabel polysilicon 1591 -2672 1591 -2672 0 1
rlabel polysilicon 1591 -2678 1591 -2678 0 3
rlabel polysilicon 1598 -2672 1598 -2672 0 1
rlabel polysilicon 1598 -2678 1598 -2678 0 3
rlabel polysilicon 1605 -2672 1605 -2672 0 1
rlabel polysilicon 1605 -2678 1605 -2678 0 3
rlabel polysilicon 1612 -2672 1612 -2672 0 1
rlabel polysilicon 1612 -2678 1612 -2678 0 3
rlabel polysilicon 1619 -2672 1619 -2672 0 1
rlabel polysilicon 1619 -2678 1619 -2678 0 3
rlabel polysilicon 1626 -2672 1626 -2672 0 1
rlabel polysilicon 1626 -2678 1626 -2678 0 3
rlabel polysilicon 1633 -2672 1633 -2672 0 1
rlabel polysilicon 1633 -2678 1633 -2678 0 3
rlabel polysilicon 1640 -2672 1640 -2672 0 1
rlabel polysilicon 1640 -2678 1640 -2678 0 3
rlabel polysilicon 1647 -2672 1647 -2672 0 1
rlabel polysilicon 1647 -2678 1647 -2678 0 3
rlabel polysilicon 1654 -2672 1654 -2672 0 1
rlabel polysilicon 1654 -2678 1654 -2678 0 3
rlabel polysilicon 1661 -2672 1661 -2672 0 1
rlabel polysilicon 1661 -2678 1661 -2678 0 3
rlabel polysilicon 1668 -2672 1668 -2672 0 1
rlabel polysilicon 1668 -2678 1668 -2678 0 3
rlabel polysilicon 1675 -2672 1675 -2672 0 1
rlabel polysilicon 1675 -2678 1675 -2678 0 3
rlabel polysilicon 1682 -2672 1682 -2672 0 1
rlabel polysilicon 1682 -2678 1682 -2678 0 3
rlabel polysilicon 1689 -2672 1689 -2672 0 1
rlabel polysilicon 1689 -2678 1689 -2678 0 3
rlabel polysilicon 1696 -2672 1696 -2672 0 1
rlabel polysilicon 1696 -2678 1696 -2678 0 3
rlabel polysilicon 1703 -2672 1703 -2672 0 1
rlabel polysilicon 1703 -2678 1703 -2678 0 3
rlabel polysilicon 1710 -2672 1710 -2672 0 1
rlabel polysilicon 1710 -2678 1710 -2678 0 3
rlabel polysilicon 1717 -2672 1717 -2672 0 1
rlabel polysilicon 1717 -2678 1717 -2678 0 3
rlabel polysilicon 1724 -2672 1724 -2672 0 1
rlabel polysilicon 1724 -2678 1724 -2678 0 3
rlabel polysilicon 1731 -2672 1731 -2672 0 1
rlabel polysilicon 1731 -2678 1731 -2678 0 3
rlabel polysilicon 1738 -2672 1738 -2672 0 1
rlabel polysilicon 1738 -2678 1738 -2678 0 3
rlabel polysilicon 1745 -2672 1745 -2672 0 1
rlabel polysilicon 1745 -2678 1745 -2678 0 3
rlabel polysilicon 1752 -2672 1752 -2672 0 1
rlabel polysilicon 1755 -2672 1755 -2672 0 2
rlabel polysilicon 1752 -2678 1752 -2678 0 3
rlabel polysilicon 1755 -2678 1755 -2678 0 4
rlabel polysilicon 1759 -2672 1759 -2672 0 1
rlabel polysilicon 1759 -2678 1759 -2678 0 3
rlabel polysilicon 1766 -2672 1766 -2672 0 1
rlabel polysilicon 1766 -2678 1766 -2678 0 3
rlabel polysilicon 1773 -2672 1773 -2672 0 1
rlabel polysilicon 1773 -2678 1773 -2678 0 3
rlabel polysilicon 1780 -2672 1780 -2672 0 1
rlabel polysilicon 1780 -2678 1780 -2678 0 3
rlabel polysilicon 1787 -2672 1787 -2672 0 1
rlabel polysilicon 1787 -2678 1787 -2678 0 3
rlabel polysilicon 1794 -2672 1794 -2672 0 1
rlabel polysilicon 1794 -2678 1794 -2678 0 3
rlabel polysilicon 1801 -2672 1801 -2672 0 1
rlabel polysilicon 1801 -2678 1801 -2678 0 3
rlabel polysilicon 1808 -2672 1808 -2672 0 1
rlabel polysilicon 1808 -2678 1808 -2678 0 3
rlabel polysilicon 1815 -2672 1815 -2672 0 1
rlabel polysilicon 1815 -2678 1815 -2678 0 3
rlabel polysilicon 1822 -2672 1822 -2672 0 1
rlabel polysilicon 1822 -2678 1822 -2678 0 3
rlabel polysilicon 1829 -2672 1829 -2672 0 1
rlabel polysilicon 1829 -2678 1829 -2678 0 3
rlabel polysilicon 1836 -2672 1836 -2672 0 1
rlabel polysilicon 1836 -2678 1836 -2678 0 3
rlabel polysilicon 1843 -2672 1843 -2672 0 1
rlabel polysilicon 1843 -2678 1843 -2678 0 3
rlabel polysilicon 1850 -2672 1850 -2672 0 1
rlabel polysilicon 1850 -2678 1850 -2678 0 3
rlabel polysilicon 1857 -2672 1857 -2672 0 1
rlabel polysilicon 1857 -2678 1857 -2678 0 3
rlabel polysilicon 1864 -2672 1864 -2672 0 1
rlabel polysilicon 1864 -2678 1864 -2678 0 3
rlabel polysilicon 1871 -2672 1871 -2672 0 1
rlabel polysilicon 1871 -2678 1871 -2678 0 3
rlabel polysilicon 1878 -2672 1878 -2672 0 1
rlabel polysilicon 1878 -2678 1878 -2678 0 3
rlabel polysilicon 1885 -2672 1885 -2672 0 1
rlabel polysilicon 1885 -2678 1885 -2678 0 3
rlabel polysilicon 1892 -2672 1892 -2672 0 1
rlabel polysilicon 1892 -2678 1892 -2678 0 3
rlabel polysilicon 1899 -2672 1899 -2672 0 1
rlabel polysilicon 1899 -2678 1899 -2678 0 3
rlabel polysilicon 1906 -2672 1906 -2672 0 1
rlabel polysilicon 1906 -2678 1906 -2678 0 3
rlabel polysilicon 1913 -2672 1913 -2672 0 1
rlabel polysilicon 1913 -2678 1913 -2678 0 3
rlabel polysilicon 1920 -2672 1920 -2672 0 1
rlabel polysilicon 1920 -2678 1920 -2678 0 3
rlabel polysilicon 1927 -2672 1927 -2672 0 1
rlabel polysilicon 1927 -2678 1927 -2678 0 3
rlabel polysilicon 1934 -2672 1934 -2672 0 1
rlabel polysilicon 1934 -2678 1934 -2678 0 3
rlabel polysilicon 1941 -2672 1941 -2672 0 1
rlabel polysilicon 1941 -2678 1941 -2678 0 3
rlabel polysilicon 1948 -2672 1948 -2672 0 1
rlabel polysilicon 1948 -2678 1948 -2678 0 3
rlabel polysilicon 1955 -2672 1955 -2672 0 1
rlabel polysilicon 1955 -2678 1955 -2678 0 3
rlabel polysilicon 1962 -2672 1962 -2672 0 1
rlabel polysilicon 1962 -2678 1962 -2678 0 3
rlabel polysilicon 1969 -2672 1969 -2672 0 1
rlabel polysilicon 1969 -2678 1969 -2678 0 3
rlabel polysilicon 1976 -2672 1976 -2672 0 1
rlabel polysilicon 1976 -2678 1976 -2678 0 3
rlabel polysilicon 1983 -2672 1983 -2672 0 1
rlabel polysilicon 1983 -2678 1983 -2678 0 3
rlabel polysilicon 1990 -2672 1990 -2672 0 1
rlabel polysilicon 1990 -2678 1990 -2678 0 3
rlabel polysilicon 1997 -2672 1997 -2672 0 1
rlabel polysilicon 1997 -2678 1997 -2678 0 3
rlabel polysilicon 2004 -2672 2004 -2672 0 1
rlabel polysilicon 2004 -2678 2004 -2678 0 3
rlabel polysilicon 2011 -2672 2011 -2672 0 1
rlabel polysilicon 2011 -2678 2011 -2678 0 3
rlabel polysilicon 2018 -2672 2018 -2672 0 1
rlabel polysilicon 2018 -2678 2018 -2678 0 3
rlabel polysilicon 2025 -2672 2025 -2672 0 1
rlabel polysilicon 2025 -2678 2025 -2678 0 3
rlabel polysilicon 2032 -2672 2032 -2672 0 1
rlabel polysilicon 2032 -2678 2032 -2678 0 3
rlabel polysilicon 2039 -2672 2039 -2672 0 1
rlabel polysilicon 2039 -2678 2039 -2678 0 3
rlabel polysilicon 2046 -2672 2046 -2672 0 1
rlabel polysilicon 2046 -2678 2046 -2678 0 3
rlabel polysilicon 2053 -2672 2053 -2672 0 1
rlabel polysilicon 2053 -2678 2053 -2678 0 3
rlabel polysilicon 2060 -2672 2060 -2672 0 1
rlabel polysilicon 2060 -2678 2060 -2678 0 3
rlabel polysilicon 2067 -2672 2067 -2672 0 1
rlabel polysilicon 2067 -2678 2067 -2678 0 3
rlabel polysilicon 2074 -2672 2074 -2672 0 1
rlabel polysilicon 2074 -2678 2074 -2678 0 3
rlabel polysilicon 2081 -2672 2081 -2672 0 1
rlabel polysilicon 2081 -2678 2081 -2678 0 3
rlabel polysilicon 2088 -2672 2088 -2672 0 1
rlabel polysilicon 2088 -2678 2088 -2678 0 3
rlabel polysilicon 2095 -2672 2095 -2672 0 1
rlabel polysilicon 2095 -2678 2095 -2678 0 3
rlabel polysilicon 2102 -2672 2102 -2672 0 1
rlabel polysilicon 2102 -2678 2102 -2678 0 3
rlabel polysilicon 2109 -2672 2109 -2672 0 1
rlabel polysilicon 2109 -2678 2109 -2678 0 3
rlabel polysilicon 2116 -2672 2116 -2672 0 1
rlabel polysilicon 2116 -2678 2116 -2678 0 3
rlabel polysilicon 2123 -2672 2123 -2672 0 1
rlabel polysilicon 2123 -2678 2123 -2678 0 3
rlabel polysilicon 2130 -2672 2130 -2672 0 1
rlabel polysilicon 2130 -2678 2130 -2678 0 3
rlabel polysilicon 2137 -2672 2137 -2672 0 1
rlabel polysilicon 2137 -2678 2137 -2678 0 3
rlabel polysilicon 2144 -2672 2144 -2672 0 1
rlabel polysilicon 2144 -2678 2144 -2678 0 3
rlabel polysilicon 2151 -2672 2151 -2672 0 1
rlabel polysilicon 2151 -2678 2151 -2678 0 3
rlabel polysilicon 2158 -2672 2158 -2672 0 1
rlabel polysilicon 2158 -2678 2158 -2678 0 3
rlabel polysilicon 2165 -2672 2165 -2672 0 1
rlabel polysilicon 2165 -2678 2165 -2678 0 3
rlabel polysilicon 2172 -2672 2172 -2672 0 1
rlabel polysilicon 2172 -2678 2172 -2678 0 3
rlabel polysilicon 2179 -2672 2179 -2672 0 1
rlabel polysilicon 2179 -2678 2179 -2678 0 3
rlabel polysilicon 2186 -2672 2186 -2672 0 1
rlabel polysilicon 2186 -2678 2186 -2678 0 3
rlabel polysilicon 2193 -2672 2193 -2672 0 1
rlabel polysilicon 2193 -2678 2193 -2678 0 3
rlabel polysilicon 2200 -2672 2200 -2672 0 1
rlabel polysilicon 2200 -2678 2200 -2678 0 3
rlabel polysilicon 2207 -2672 2207 -2672 0 1
rlabel polysilicon 2207 -2678 2207 -2678 0 3
rlabel polysilicon 2214 -2672 2214 -2672 0 1
rlabel polysilicon 2214 -2678 2214 -2678 0 3
rlabel polysilicon 2221 -2672 2221 -2672 0 1
rlabel polysilicon 2221 -2678 2221 -2678 0 3
rlabel polysilicon 2228 -2672 2228 -2672 0 1
rlabel polysilicon 2228 -2678 2228 -2678 0 3
rlabel polysilicon 2235 -2672 2235 -2672 0 1
rlabel polysilicon 2235 -2678 2235 -2678 0 3
rlabel polysilicon 2242 -2672 2242 -2672 0 1
rlabel polysilicon 2242 -2678 2242 -2678 0 3
rlabel polysilicon 2263 -2672 2263 -2672 0 1
rlabel polysilicon 2263 -2678 2263 -2678 0 3
rlabel polysilicon 2270 -2672 2270 -2672 0 1
rlabel polysilicon 2270 -2678 2270 -2678 0 3
rlabel polysilicon 2 -2835 2 -2835 0 1
rlabel polysilicon 2 -2841 2 -2841 0 3
rlabel polysilicon 9 -2835 9 -2835 0 1
rlabel polysilicon 9 -2841 9 -2841 0 3
rlabel polysilicon 16 -2835 16 -2835 0 1
rlabel polysilicon 16 -2841 16 -2841 0 3
rlabel polysilicon 23 -2835 23 -2835 0 1
rlabel polysilicon 23 -2841 23 -2841 0 3
rlabel polysilicon 30 -2835 30 -2835 0 1
rlabel polysilicon 30 -2841 30 -2841 0 3
rlabel polysilicon 37 -2835 37 -2835 0 1
rlabel polysilicon 37 -2841 37 -2841 0 3
rlabel polysilicon 44 -2835 44 -2835 0 1
rlabel polysilicon 44 -2841 44 -2841 0 3
rlabel polysilicon 51 -2835 51 -2835 0 1
rlabel polysilicon 54 -2835 54 -2835 0 2
rlabel polysilicon 51 -2841 51 -2841 0 3
rlabel polysilicon 58 -2835 58 -2835 0 1
rlabel polysilicon 58 -2841 58 -2841 0 3
rlabel polysilicon 65 -2835 65 -2835 0 1
rlabel polysilicon 65 -2841 65 -2841 0 3
rlabel polysilicon 72 -2835 72 -2835 0 1
rlabel polysilicon 72 -2841 72 -2841 0 3
rlabel polysilicon 79 -2835 79 -2835 0 1
rlabel polysilicon 82 -2835 82 -2835 0 2
rlabel polysilicon 79 -2841 79 -2841 0 3
rlabel polysilicon 82 -2841 82 -2841 0 4
rlabel polysilicon 86 -2835 86 -2835 0 1
rlabel polysilicon 86 -2841 86 -2841 0 3
rlabel polysilicon 93 -2835 93 -2835 0 1
rlabel polysilicon 93 -2841 93 -2841 0 3
rlabel polysilicon 100 -2835 100 -2835 0 1
rlabel polysilicon 100 -2841 100 -2841 0 3
rlabel polysilicon 110 -2835 110 -2835 0 2
rlabel polysilicon 107 -2841 107 -2841 0 3
rlabel polysilicon 114 -2835 114 -2835 0 1
rlabel polysilicon 114 -2841 114 -2841 0 3
rlabel polysilicon 121 -2835 121 -2835 0 1
rlabel polysilicon 121 -2841 121 -2841 0 3
rlabel polysilicon 128 -2835 128 -2835 0 1
rlabel polysilicon 128 -2841 128 -2841 0 3
rlabel polysilicon 135 -2835 135 -2835 0 1
rlabel polysilicon 135 -2841 135 -2841 0 3
rlabel polysilicon 142 -2835 142 -2835 0 1
rlabel polysilicon 142 -2841 142 -2841 0 3
rlabel polysilicon 149 -2835 149 -2835 0 1
rlabel polysilicon 149 -2841 149 -2841 0 3
rlabel polysilicon 156 -2835 156 -2835 0 1
rlabel polysilicon 156 -2841 156 -2841 0 3
rlabel polysilicon 163 -2835 163 -2835 0 1
rlabel polysilicon 163 -2841 163 -2841 0 3
rlabel polysilicon 170 -2835 170 -2835 0 1
rlabel polysilicon 170 -2841 170 -2841 0 3
rlabel polysilicon 177 -2835 177 -2835 0 1
rlabel polysilicon 177 -2841 177 -2841 0 3
rlabel polysilicon 184 -2835 184 -2835 0 1
rlabel polysilicon 184 -2841 184 -2841 0 3
rlabel polysilicon 191 -2835 191 -2835 0 1
rlabel polysilicon 191 -2841 191 -2841 0 3
rlabel polysilicon 198 -2835 198 -2835 0 1
rlabel polysilicon 198 -2841 198 -2841 0 3
rlabel polysilicon 205 -2835 205 -2835 0 1
rlabel polysilicon 205 -2841 205 -2841 0 3
rlabel polysilicon 212 -2835 212 -2835 0 1
rlabel polysilicon 212 -2841 212 -2841 0 3
rlabel polysilicon 219 -2835 219 -2835 0 1
rlabel polysilicon 222 -2835 222 -2835 0 2
rlabel polysilicon 219 -2841 219 -2841 0 3
rlabel polysilicon 222 -2841 222 -2841 0 4
rlabel polysilicon 226 -2835 226 -2835 0 1
rlabel polysilicon 226 -2841 226 -2841 0 3
rlabel polysilicon 236 -2835 236 -2835 0 2
rlabel polysilicon 233 -2841 233 -2841 0 3
rlabel polysilicon 236 -2841 236 -2841 0 4
rlabel polysilicon 240 -2835 240 -2835 0 1
rlabel polysilicon 240 -2841 240 -2841 0 3
rlabel polysilicon 247 -2835 247 -2835 0 1
rlabel polysilicon 250 -2835 250 -2835 0 2
rlabel polysilicon 247 -2841 247 -2841 0 3
rlabel polysilicon 250 -2841 250 -2841 0 4
rlabel polysilicon 254 -2835 254 -2835 0 1
rlabel polysilicon 254 -2841 254 -2841 0 3
rlabel polysilicon 261 -2835 261 -2835 0 1
rlabel polysilicon 261 -2841 261 -2841 0 3
rlabel polysilicon 268 -2835 268 -2835 0 1
rlabel polysilicon 268 -2841 268 -2841 0 3
rlabel polysilicon 275 -2835 275 -2835 0 1
rlabel polysilicon 275 -2841 275 -2841 0 3
rlabel polysilicon 282 -2835 282 -2835 0 1
rlabel polysilicon 282 -2841 282 -2841 0 3
rlabel polysilicon 289 -2835 289 -2835 0 1
rlabel polysilicon 289 -2841 289 -2841 0 3
rlabel polysilicon 296 -2835 296 -2835 0 1
rlabel polysilicon 296 -2841 296 -2841 0 3
rlabel polysilicon 303 -2835 303 -2835 0 1
rlabel polysilicon 303 -2841 303 -2841 0 3
rlabel polysilicon 310 -2835 310 -2835 0 1
rlabel polysilicon 310 -2841 310 -2841 0 3
rlabel polysilicon 317 -2835 317 -2835 0 1
rlabel polysilicon 317 -2841 317 -2841 0 3
rlabel polysilicon 324 -2835 324 -2835 0 1
rlabel polysilicon 324 -2841 324 -2841 0 3
rlabel polysilicon 331 -2835 331 -2835 0 1
rlabel polysilicon 331 -2841 331 -2841 0 3
rlabel polysilicon 338 -2835 338 -2835 0 1
rlabel polysilicon 338 -2841 338 -2841 0 3
rlabel polysilicon 345 -2835 345 -2835 0 1
rlabel polysilicon 345 -2841 345 -2841 0 3
rlabel polysilicon 352 -2835 352 -2835 0 1
rlabel polysilicon 352 -2841 352 -2841 0 3
rlabel polysilicon 359 -2835 359 -2835 0 1
rlabel polysilicon 359 -2841 359 -2841 0 3
rlabel polysilicon 366 -2835 366 -2835 0 1
rlabel polysilicon 366 -2841 366 -2841 0 3
rlabel polysilicon 373 -2835 373 -2835 0 1
rlabel polysilicon 373 -2841 373 -2841 0 3
rlabel polysilicon 380 -2835 380 -2835 0 1
rlabel polysilicon 380 -2841 380 -2841 0 3
rlabel polysilicon 387 -2835 387 -2835 0 1
rlabel polysilicon 387 -2841 387 -2841 0 3
rlabel polysilicon 394 -2835 394 -2835 0 1
rlabel polysilicon 394 -2841 394 -2841 0 3
rlabel polysilicon 401 -2835 401 -2835 0 1
rlabel polysilicon 401 -2841 401 -2841 0 3
rlabel polysilicon 408 -2835 408 -2835 0 1
rlabel polysilicon 408 -2841 408 -2841 0 3
rlabel polysilicon 415 -2835 415 -2835 0 1
rlabel polysilicon 415 -2841 415 -2841 0 3
rlabel polysilicon 422 -2835 422 -2835 0 1
rlabel polysilicon 422 -2841 422 -2841 0 3
rlabel polysilicon 432 -2835 432 -2835 0 2
rlabel polysilicon 429 -2841 429 -2841 0 3
rlabel polysilicon 436 -2835 436 -2835 0 1
rlabel polysilicon 436 -2841 436 -2841 0 3
rlabel polysilicon 443 -2835 443 -2835 0 1
rlabel polysilicon 443 -2841 443 -2841 0 3
rlabel polysilicon 450 -2835 450 -2835 0 1
rlabel polysilicon 450 -2841 450 -2841 0 3
rlabel polysilicon 457 -2835 457 -2835 0 1
rlabel polysilicon 460 -2835 460 -2835 0 2
rlabel polysilicon 460 -2841 460 -2841 0 4
rlabel polysilicon 464 -2835 464 -2835 0 1
rlabel polysilicon 464 -2841 464 -2841 0 3
rlabel polysilicon 471 -2835 471 -2835 0 1
rlabel polysilicon 471 -2841 471 -2841 0 3
rlabel polysilicon 478 -2835 478 -2835 0 1
rlabel polysilicon 478 -2841 478 -2841 0 3
rlabel polysilicon 485 -2835 485 -2835 0 1
rlabel polysilicon 485 -2841 485 -2841 0 3
rlabel polysilicon 492 -2835 492 -2835 0 1
rlabel polysilicon 492 -2841 492 -2841 0 3
rlabel polysilicon 499 -2835 499 -2835 0 1
rlabel polysilicon 499 -2841 499 -2841 0 3
rlabel polysilicon 506 -2835 506 -2835 0 1
rlabel polysilicon 506 -2841 506 -2841 0 3
rlabel polysilicon 513 -2835 513 -2835 0 1
rlabel polysilicon 513 -2841 513 -2841 0 3
rlabel polysilicon 520 -2835 520 -2835 0 1
rlabel polysilicon 520 -2841 520 -2841 0 3
rlabel polysilicon 527 -2835 527 -2835 0 1
rlabel polysilicon 527 -2841 527 -2841 0 3
rlabel polysilicon 534 -2835 534 -2835 0 1
rlabel polysilicon 534 -2841 534 -2841 0 3
rlabel polysilicon 541 -2835 541 -2835 0 1
rlabel polysilicon 544 -2835 544 -2835 0 2
rlabel polysilicon 544 -2841 544 -2841 0 4
rlabel polysilicon 548 -2835 548 -2835 0 1
rlabel polysilicon 548 -2841 548 -2841 0 3
rlabel polysilicon 555 -2835 555 -2835 0 1
rlabel polysilicon 555 -2841 555 -2841 0 3
rlabel polysilicon 562 -2835 562 -2835 0 1
rlabel polysilicon 562 -2841 562 -2841 0 3
rlabel polysilicon 569 -2835 569 -2835 0 1
rlabel polysilicon 569 -2841 569 -2841 0 3
rlabel polysilicon 576 -2835 576 -2835 0 1
rlabel polysilicon 576 -2841 576 -2841 0 3
rlabel polysilicon 583 -2835 583 -2835 0 1
rlabel polysilicon 583 -2841 583 -2841 0 3
rlabel polysilicon 590 -2835 590 -2835 0 1
rlabel polysilicon 590 -2841 590 -2841 0 3
rlabel polysilicon 597 -2835 597 -2835 0 1
rlabel polysilicon 597 -2841 597 -2841 0 3
rlabel polysilicon 604 -2835 604 -2835 0 1
rlabel polysilicon 604 -2841 604 -2841 0 3
rlabel polysilicon 611 -2835 611 -2835 0 1
rlabel polysilicon 611 -2841 611 -2841 0 3
rlabel polysilicon 618 -2835 618 -2835 0 1
rlabel polysilicon 621 -2835 621 -2835 0 2
rlabel polysilicon 618 -2841 618 -2841 0 3
rlabel polysilicon 621 -2841 621 -2841 0 4
rlabel polysilicon 625 -2835 625 -2835 0 1
rlabel polysilicon 625 -2841 625 -2841 0 3
rlabel polysilicon 632 -2835 632 -2835 0 1
rlabel polysilicon 632 -2841 632 -2841 0 3
rlabel polysilicon 639 -2835 639 -2835 0 1
rlabel polysilicon 639 -2841 639 -2841 0 3
rlabel polysilicon 646 -2835 646 -2835 0 1
rlabel polysilicon 646 -2841 646 -2841 0 3
rlabel polysilicon 653 -2835 653 -2835 0 1
rlabel polysilicon 653 -2841 653 -2841 0 3
rlabel polysilicon 660 -2835 660 -2835 0 1
rlabel polysilicon 663 -2835 663 -2835 0 2
rlabel polysilicon 660 -2841 660 -2841 0 3
rlabel polysilicon 663 -2841 663 -2841 0 4
rlabel polysilicon 667 -2835 667 -2835 0 1
rlabel polysilicon 667 -2841 667 -2841 0 3
rlabel polysilicon 674 -2835 674 -2835 0 1
rlabel polysilicon 674 -2841 674 -2841 0 3
rlabel polysilicon 681 -2835 681 -2835 0 1
rlabel polysilicon 681 -2841 681 -2841 0 3
rlabel polysilicon 688 -2835 688 -2835 0 1
rlabel polysilicon 688 -2841 688 -2841 0 3
rlabel polysilicon 695 -2835 695 -2835 0 1
rlabel polysilicon 695 -2841 695 -2841 0 3
rlabel polysilicon 702 -2835 702 -2835 0 1
rlabel polysilicon 705 -2835 705 -2835 0 2
rlabel polysilicon 702 -2841 702 -2841 0 3
rlabel polysilicon 705 -2841 705 -2841 0 4
rlabel polysilicon 709 -2835 709 -2835 0 1
rlabel polysilicon 709 -2841 709 -2841 0 3
rlabel polysilicon 716 -2835 716 -2835 0 1
rlabel polysilicon 716 -2841 716 -2841 0 3
rlabel polysilicon 723 -2835 723 -2835 0 1
rlabel polysilicon 723 -2841 723 -2841 0 3
rlabel polysilicon 730 -2835 730 -2835 0 1
rlabel polysilicon 733 -2835 733 -2835 0 2
rlabel polysilicon 730 -2841 730 -2841 0 3
rlabel polysilicon 733 -2841 733 -2841 0 4
rlabel polysilicon 737 -2835 737 -2835 0 1
rlabel polysilicon 737 -2841 737 -2841 0 3
rlabel polysilicon 744 -2835 744 -2835 0 1
rlabel polysilicon 744 -2841 744 -2841 0 3
rlabel polysilicon 747 -2841 747 -2841 0 4
rlabel polysilicon 751 -2835 751 -2835 0 1
rlabel polysilicon 751 -2841 751 -2841 0 3
rlabel polysilicon 758 -2835 758 -2835 0 1
rlabel polysilicon 758 -2841 758 -2841 0 3
rlabel polysilicon 765 -2835 765 -2835 0 1
rlabel polysilicon 765 -2841 765 -2841 0 3
rlabel polysilicon 772 -2835 772 -2835 0 1
rlabel polysilicon 772 -2841 772 -2841 0 3
rlabel polysilicon 779 -2835 779 -2835 0 1
rlabel polysilicon 779 -2841 779 -2841 0 3
rlabel polysilicon 786 -2835 786 -2835 0 1
rlabel polysilicon 789 -2835 789 -2835 0 2
rlabel polysilicon 789 -2841 789 -2841 0 4
rlabel polysilicon 793 -2835 793 -2835 0 1
rlabel polysilicon 793 -2841 793 -2841 0 3
rlabel polysilicon 800 -2835 800 -2835 0 1
rlabel polysilicon 800 -2841 800 -2841 0 3
rlabel polysilicon 807 -2835 807 -2835 0 1
rlabel polysilicon 807 -2841 807 -2841 0 3
rlabel polysilicon 814 -2835 814 -2835 0 1
rlabel polysilicon 814 -2841 814 -2841 0 3
rlabel polysilicon 821 -2835 821 -2835 0 1
rlabel polysilicon 821 -2841 821 -2841 0 3
rlabel polysilicon 828 -2835 828 -2835 0 1
rlabel polysilicon 828 -2841 828 -2841 0 3
rlabel polysilicon 835 -2835 835 -2835 0 1
rlabel polysilicon 838 -2835 838 -2835 0 2
rlabel polysilicon 842 -2835 842 -2835 0 1
rlabel polysilicon 842 -2841 842 -2841 0 3
rlabel polysilicon 849 -2835 849 -2835 0 1
rlabel polysilicon 849 -2841 849 -2841 0 3
rlabel polysilicon 856 -2835 856 -2835 0 1
rlabel polysilicon 856 -2841 856 -2841 0 3
rlabel polysilicon 863 -2835 863 -2835 0 1
rlabel polysilicon 866 -2835 866 -2835 0 2
rlabel polysilicon 863 -2841 863 -2841 0 3
rlabel polysilicon 866 -2841 866 -2841 0 4
rlabel polysilicon 870 -2835 870 -2835 0 1
rlabel polysilicon 870 -2841 870 -2841 0 3
rlabel polysilicon 877 -2835 877 -2835 0 1
rlabel polysilicon 877 -2841 877 -2841 0 3
rlabel polysilicon 884 -2835 884 -2835 0 1
rlabel polysilicon 884 -2841 884 -2841 0 3
rlabel polysilicon 891 -2835 891 -2835 0 1
rlabel polysilicon 891 -2841 891 -2841 0 3
rlabel polysilicon 898 -2835 898 -2835 0 1
rlabel polysilicon 898 -2841 898 -2841 0 3
rlabel polysilicon 905 -2835 905 -2835 0 1
rlabel polysilicon 905 -2841 905 -2841 0 3
rlabel polysilicon 912 -2835 912 -2835 0 1
rlabel polysilicon 915 -2835 915 -2835 0 2
rlabel polysilicon 912 -2841 912 -2841 0 3
rlabel polysilicon 919 -2835 919 -2835 0 1
rlabel polysilicon 919 -2841 919 -2841 0 3
rlabel polysilicon 926 -2835 926 -2835 0 1
rlabel polysilicon 926 -2841 926 -2841 0 3
rlabel polysilicon 933 -2835 933 -2835 0 1
rlabel polysilicon 933 -2841 933 -2841 0 3
rlabel polysilicon 940 -2835 940 -2835 0 1
rlabel polysilicon 943 -2835 943 -2835 0 2
rlabel polysilicon 940 -2841 940 -2841 0 3
rlabel polysilicon 943 -2841 943 -2841 0 4
rlabel polysilicon 947 -2835 947 -2835 0 1
rlabel polysilicon 947 -2841 947 -2841 0 3
rlabel polysilicon 954 -2835 954 -2835 0 1
rlabel polysilicon 954 -2841 954 -2841 0 3
rlabel polysilicon 961 -2835 961 -2835 0 1
rlabel polysilicon 964 -2835 964 -2835 0 2
rlabel polysilicon 961 -2841 961 -2841 0 3
rlabel polysilicon 968 -2835 968 -2835 0 1
rlabel polysilicon 968 -2841 968 -2841 0 3
rlabel polysilicon 975 -2835 975 -2835 0 1
rlabel polysilicon 978 -2835 978 -2835 0 2
rlabel polysilicon 978 -2841 978 -2841 0 4
rlabel polysilicon 982 -2835 982 -2835 0 1
rlabel polysilicon 982 -2841 982 -2841 0 3
rlabel polysilicon 989 -2835 989 -2835 0 1
rlabel polysilicon 989 -2841 989 -2841 0 3
rlabel polysilicon 996 -2835 996 -2835 0 1
rlabel polysilicon 996 -2841 996 -2841 0 3
rlabel polysilicon 1003 -2835 1003 -2835 0 1
rlabel polysilicon 1003 -2841 1003 -2841 0 3
rlabel polysilicon 1010 -2835 1010 -2835 0 1
rlabel polysilicon 1010 -2841 1010 -2841 0 3
rlabel polysilicon 1017 -2835 1017 -2835 0 1
rlabel polysilicon 1017 -2841 1017 -2841 0 3
rlabel polysilicon 1024 -2835 1024 -2835 0 1
rlabel polysilicon 1024 -2841 1024 -2841 0 3
rlabel polysilicon 1031 -2835 1031 -2835 0 1
rlabel polysilicon 1031 -2841 1031 -2841 0 3
rlabel polysilicon 1038 -2835 1038 -2835 0 1
rlabel polysilicon 1038 -2841 1038 -2841 0 3
rlabel polysilicon 1045 -2835 1045 -2835 0 1
rlabel polysilicon 1045 -2841 1045 -2841 0 3
rlabel polysilicon 1052 -2835 1052 -2835 0 1
rlabel polysilicon 1055 -2835 1055 -2835 0 2
rlabel polysilicon 1052 -2841 1052 -2841 0 3
rlabel polysilicon 1055 -2841 1055 -2841 0 4
rlabel polysilicon 1059 -2835 1059 -2835 0 1
rlabel polysilicon 1062 -2835 1062 -2835 0 2
rlabel polysilicon 1059 -2841 1059 -2841 0 3
rlabel polysilicon 1066 -2835 1066 -2835 0 1
rlabel polysilicon 1066 -2841 1066 -2841 0 3
rlabel polysilicon 1073 -2835 1073 -2835 0 1
rlabel polysilicon 1073 -2841 1073 -2841 0 3
rlabel polysilicon 1080 -2835 1080 -2835 0 1
rlabel polysilicon 1080 -2841 1080 -2841 0 3
rlabel polysilicon 1087 -2835 1087 -2835 0 1
rlabel polysilicon 1087 -2841 1087 -2841 0 3
rlabel polysilicon 1094 -2835 1094 -2835 0 1
rlabel polysilicon 1097 -2835 1097 -2835 0 2
rlabel polysilicon 1094 -2841 1094 -2841 0 3
rlabel polysilicon 1097 -2841 1097 -2841 0 4
rlabel polysilicon 1101 -2835 1101 -2835 0 1
rlabel polysilicon 1101 -2841 1101 -2841 0 3
rlabel polysilicon 1108 -2835 1108 -2835 0 1
rlabel polysilicon 1108 -2841 1108 -2841 0 3
rlabel polysilicon 1115 -2835 1115 -2835 0 1
rlabel polysilicon 1115 -2841 1115 -2841 0 3
rlabel polysilicon 1122 -2835 1122 -2835 0 1
rlabel polysilicon 1122 -2841 1122 -2841 0 3
rlabel polysilicon 1129 -2835 1129 -2835 0 1
rlabel polysilicon 1129 -2841 1129 -2841 0 3
rlabel polysilicon 1136 -2835 1136 -2835 0 1
rlabel polysilicon 1136 -2841 1136 -2841 0 3
rlabel polysilicon 1143 -2835 1143 -2835 0 1
rlabel polysilicon 1143 -2841 1143 -2841 0 3
rlabel polysilicon 1150 -2835 1150 -2835 0 1
rlabel polysilicon 1150 -2841 1150 -2841 0 3
rlabel polysilicon 1157 -2835 1157 -2835 0 1
rlabel polysilicon 1157 -2841 1157 -2841 0 3
rlabel polysilicon 1164 -2835 1164 -2835 0 1
rlabel polysilicon 1164 -2841 1164 -2841 0 3
rlabel polysilicon 1171 -2835 1171 -2835 0 1
rlabel polysilicon 1171 -2841 1171 -2841 0 3
rlabel polysilicon 1178 -2835 1178 -2835 0 1
rlabel polysilicon 1178 -2841 1178 -2841 0 3
rlabel polysilicon 1185 -2835 1185 -2835 0 1
rlabel polysilicon 1185 -2841 1185 -2841 0 3
rlabel polysilicon 1192 -2835 1192 -2835 0 1
rlabel polysilicon 1192 -2841 1192 -2841 0 3
rlabel polysilicon 1199 -2835 1199 -2835 0 1
rlabel polysilicon 1199 -2841 1199 -2841 0 3
rlabel polysilicon 1206 -2835 1206 -2835 0 1
rlabel polysilicon 1206 -2841 1206 -2841 0 3
rlabel polysilicon 1213 -2835 1213 -2835 0 1
rlabel polysilicon 1213 -2841 1213 -2841 0 3
rlabel polysilicon 1220 -2835 1220 -2835 0 1
rlabel polysilicon 1220 -2841 1220 -2841 0 3
rlabel polysilicon 1227 -2835 1227 -2835 0 1
rlabel polysilicon 1227 -2841 1227 -2841 0 3
rlabel polysilicon 1234 -2835 1234 -2835 0 1
rlabel polysilicon 1234 -2841 1234 -2841 0 3
rlabel polysilicon 1241 -2835 1241 -2835 0 1
rlabel polysilicon 1241 -2841 1241 -2841 0 3
rlabel polysilicon 1248 -2835 1248 -2835 0 1
rlabel polysilicon 1248 -2841 1248 -2841 0 3
rlabel polysilicon 1255 -2835 1255 -2835 0 1
rlabel polysilicon 1258 -2835 1258 -2835 0 2
rlabel polysilicon 1258 -2841 1258 -2841 0 4
rlabel polysilicon 1262 -2835 1262 -2835 0 1
rlabel polysilicon 1262 -2841 1262 -2841 0 3
rlabel polysilicon 1269 -2835 1269 -2835 0 1
rlabel polysilicon 1269 -2841 1269 -2841 0 3
rlabel polysilicon 1276 -2835 1276 -2835 0 1
rlabel polysilicon 1276 -2841 1276 -2841 0 3
rlabel polysilicon 1283 -2835 1283 -2835 0 1
rlabel polysilicon 1286 -2835 1286 -2835 0 2
rlabel polysilicon 1286 -2841 1286 -2841 0 4
rlabel polysilicon 1290 -2835 1290 -2835 0 1
rlabel polysilicon 1290 -2841 1290 -2841 0 3
rlabel polysilicon 1297 -2835 1297 -2835 0 1
rlabel polysilicon 1297 -2841 1297 -2841 0 3
rlabel polysilicon 1304 -2835 1304 -2835 0 1
rlabel polysilicon 1304 -2841 1304 -2841 0 3
rlabel polysilicon 1311 -2835 1311 -2835 0 1
rlabel polysilicon 1314 -2835 1314 -2835 0 2
rlabel polysilicon 1311 -2841 1311 -2841 0 3
rlabel polysilicon 1314 -2841 1314 -2841 0 4
rlabel polysilicon 1318 -2835 1318 -2835 0 1
rlabel polysilicon 1318 -2841 1318 -2841 0 3
rlabel polysilicon 1325 -2835 1325 -2835 0 1
rlabel polysilicon 1325 -2841 1325 -2841 0 3
rlabel polysilicon 1332 -2835 1332 -2835 0 1
rlabel polysilicon 1332 -2841 1332 -2841 0 3
rlabel polysilicon 1339 -2835 1339 -2835 0 1
rlabel polysilicon 1339 -2841 1339 -2841 0 3
rlabel polysilicon 1346 -2835 1346 -2835 0 1
rlabel polysilicon 1346 -2841 1346 -2841 0 3
rlabel polysilicon 1349 -2841 1349 -2841 0 4
rlabel polysilicon 1353 -2835 1353 -2835 0 1
rlabel polysilicon 1353 -2841 1353 -2841 0 3
rlabel polysilicon 1360 -2835 1360 -2835 0 1
rlabel polysilicon 1360 -2841 1360 -2841 0 3
rlabel polysilicon 1367 -2835 1367 -2835 0 1
rlabel polysilicon 1367 -2841 1367 -2841 0 3
rlabel polysilicon 1374 -2835 1374 -2835 0 1
rlabel polysilicon 1374 -2841 1374 -2841 0 3
rlabel polysilicon 1381 -2835 1381 -2835 0 1
rlabel polysilicon 1381 -2841 1381 -2841 0 3
rlabel polysilicon 1391 -2835 1391 -2835 0 2
rlabel polysilicon 1388 -2841 1388 -2841 0 3
rlabel polysilicon 1391 -2841 1391 -2841 0 4
rlabel polysilicon 1395 -2835 1395 -2835 0 1
rlabel polysilicon 1395 -2841 1395 -2841 0 3
rlabel polysilicon 1402 -2835 1402 -2835 0 1
rlabel polysilicon 1402 -2841 1402 -2841 0 3
rlabel polysilicon 1409 -2835 1409 -2835 0 1
rlabel polysilicon 1409 -2841 1409 -2841 0 3
rlabel polysilicon 1416 -2835 1416 -2835 0 1
rlabel polysilicon 1416 -2841 1416 -2841 0 3
rlabel polysilicon 1423 -2835 1423 -2835 0 1
rlabel polysilicon 1423 -2841 1423 -2841 0 3
rlabel polysilicon 1433 -2835 1433 -2835 0 2
rlabel polysilicon 1430 -2841 1430 -2841 0 3
rlabel polysilicon 1433 -2841 1433 -2841 0 4
rlabel polysilicon 1437 -2835 1437 -2835 0 1
rlabel polysilicon 1437 -2841 1437 -2841 0 3
rlabel polysilicon 1444 -2835 1444 -2835 0 1
rlabel polysilicon 1444 -2841 1444 -2841 0 3
rlabel polysilicon 1451 -2835 1451 -2835 0 1
rlabel polysilicon 1451 -2841 1451 -2841 0 3
rlabel polysilicon 1458 -2835 1458 -2835 0 1
rlabel polysilicon 1458 -2841 1458 -2841 0 3
rlabel polysilicon 1465 -2835 1465 -2835 0 1
rlabel polysilicon 1465 -2841 1465 -2841 0 3
rlabel polysilicon 1472 -2835 1472 -2835 0 1
rlabel polysilicon 1472 -2841 1472 -2841 0 3
rlabel polysilicon 1479 -2835 1479 -2835 0 1
rlabel polysilicon 1479 -2841 1479 -2841 0 3
rlabel polysilicon 1489 -2835 1489 -2835 0 2
rlabel polysilicon 1486 -2841 1486 -2841 0 3
rlabel polysilicon 1489 -2841 1489 -2841 0 4
rlabel polysilicon 1493 -2835 1493 -2835 0 1
rlabel polysilicon 1496 -2835 1496 -2835 0 2
rlabel polysilicon 1493 -2841 1493 -2841 0 3
rlabel polysilicon 1496 -2841 1496 -2841 0 4
rlabel polysilicon 1500 -2835 1500 -2835 0 1
rlabel polysilicon 1500 -2841 1500 -2841 0 3
rlabel polysilicon 1507 -2835 1507 -2835 0 1
rlabel polysilicon 1507 -2841 1507 -2841 0 3
rlabel polysilicon 1514 -2835 1514 -2835 0 1
rlabel polysilicon 1514 -2841 1514 -2841 0 3
rlabel polysilicon 1521 -2835 1521 -2835 0 1
rlabel polysilicon 1521 -2841 1521 -2841 0 3
rlabel polysilicon 1528 -2835 1528 -2835 0 1
rlabel polysilicon 1528 -2841 1528 -2841 0 3
rlabel polysilicon 1535 -2835 1535 -2835 0 1
rlabel polysilicon 1535 -2841 1535 -2841 0 3
rlabel polysilicon 1542 -2835 1542 -2835 0 1
rlabel polysilicon 1542 -2841 1542 -2841 0 3
rlabel polysilicon 1549 -2835 1549 -2835 0 1
rlabel polysilicon 1549 -2841 1549 -2841 0 3
rlabel polysilicon 1556 -2835 1556 -2835 0 1
rlabel polysilicon 1556 -2841 1556 -2841 0 3
rlabel polysilicon 1563 -2841 1563 -2841 0 3
rlabel polysilicon 1566 -2841 1566 -2841 0 4
rlabel polysilicon 1570 -2835 1570 -2835 0 1
rlabel polysilicon 1570 -2841 1570 -2841 0 3
rlabel polysilicon 1577 -2835 1577 -2835 0 1
rlabel polysilicon 1577 -2841 1577 -2841 0 3
rlabel polysilicon 1584 -2835 1584 -2835 0 1
rlabel polysilicon 1584 -2841 1584 -2841 0 3
rlabel polysilicon 1591 -2835 1591 -2835 0 1
rlabel polysilicon 1591 -2841 1591 -2841 0 3
rlabel polysilicon 1598 -2835 1598 -2835 0 1
rlabel polysilicon 1598 -2841 1598 -2841 0 3
rlabel polysilicon 1605 -2835 1605 -2835 0 1
rlabel polysilicon 1605 -2841 1605 -2841 0 3
rlabel polysilicon 1612 -2835 1612 -2835 0 1
rlabel polysilicon 1612 -2841 1612 -2841 0 3
rlabel polysilicon 1619 -2835 1619 -2835 0 1
rlabel polysilicon 1619 -2841 1619 -2841 0 3
rlabel polysilicon 1626 -2835 1626 -2835 0 1
rlabel polysilicon 1626 -2841 1626 -2841 0 3
rlabel polysilicon 1633 -2835 1633 -2835 0 1
rlabel polysilicon 1633 -2841 1633 -2841 0 3
rlabel polysilicon 1640 -2835 1640 -2835 0 1
rlabel polysilicon 1640 -2841 1640 -2841 0 3
rlabel polysilicon 1647 -2835 1647 -2835 0 1
rlabel polysilicon 1647 -2841 1647 -2841 0 3
rlabel polysilicon 1654 -2835 1654 -2835 0 1
rlabel polysilicon 1654 -2841 1654 -2841 0 3
rlabel polysilicon 1661 -2835 1661 -2835 0 1
rlabel polysilicon 1661 -2841 1661 -2841 0 3
rlabel polysilicon 1668 -2835 1668 -2835 0 1
rlabel polysilicon 1668 -2841 1668 -2841 0 3
rlabel polysilicon 1675 -2835 1675 -2835 0 1
rlabel polysilicon 1675 -2841 1675 -2841 0 3
rlabel polysilicon 1685 -2835 1685 -2835 0 2
rlabel polysilicon 1682 -2841 1682 -2841 0 3
rlabel polysilicon 1685 -2841 1685 -2841 0 4
rlabel polysilicon 1689 -2835 1689 -2835 0 1
rlabel polysilicon 1689 -2841 1689 -2841 0 3
rlabel polysilicon 1696 -2835 1696 -2835 0 1
rlabel polysilicon 1696 -2841 1696 -2841 0 3
rlabel polysilicon 1706 -2835 1706 -2835 0 2
rlabel polysilicon 1703 -2841 1703 -2841 0 3
rlabel polysilicon 1706 -2841 1706 -2841 0 4
rlabel polysilicon 1710 -2835 1710 -2835 0 1
rlabel polysilicon 1710 -2841 1710 -2841 0 3
rlabel polysilicon 1717 -2835 1717 -2835 0 1
rlabel polysilicon 1717 -2841 1717 -2841 0 3
rlabel polysilicon 1724 -2835 1724 -2835 0 1
rlabel polysilicon 1724 -2841 1724 -2841 0 3
rlabel polysilicon 1731 -2835 1731 -2835 0 1
rlabel polysilicon 1731 -2841 1731 -2841 0 3
rlabel polysilicon 1738 -2835 1738 -2835 0 1
rlabel polysilicon 1738 -2841 1738 -2841 0 3
rlabel polysilicon 1745 -2835 1745 -2835 0 1
rlabel polysilicon 1745 -2841 1745 -2841 0 3
rlabel polysilicon 1755 -2835 1755 -2835 0 2
rlabel polysilicon 1752 -2841 1752 -2841 0 3
rlabel polysilicon 1755 -2841 1755 -2841 0 4
rlabel polysilicon 1759 -2835 1759 -2835 0 1
rlabel polysilicon 1759 -2841 1759 -2841 0 3
rlabel polysilicon 1766 -2835 1766 -2835 0 1
rlabel polysilicon 1766 -2841 1766 -2841 0 3
rlabel polysilicon 1773 -2835 1773 -2835 0 1
rlabel polysilicon 1773 -2841 1773 -2841 0 3
rlabel polysilicon 1780 -2835 1780 -2835 0 1
rlabel polysilicon 1780 -2841 1780 -2841 0 3
rlabel polysilicon 1787 -2835 1787 -2835 0 1
rlabel polysilicon 1787 -2841 1787 -2841 0 3
rlabel polysilicon 1794 -2835 1794 -2835 0 1
rlabel polysilicon 1794 -2841 1794 -2841 0 3
rlabel polysilicon 1801 -2835 1801 -2835 0 1
rlabel polysilicon 1801 -2841 1801 -2841 0 3
rlabel polysilicon 1808 -2835 1808 -2835 0 1
rlabel polysilicon 1808 -2841 1808 -2841 0 3
rlabel polysilicon 1815 -2835 1815 -2835 0 1
rlabel polysilicon 1815 -2841 1815 -2841 0 3
rlabel polysilicon 1822 -2835 1822 -2835 0 1
rlabel polysilicon 1822 -2841 1822 -2841 0 3
rlabel polysilicon 1829 -2835 1829 -2835 0 1
rlabel polysilicon 1829 -2841 1829 -2841 0 3
rlabel polysilicon 1836 -2835 1836 -2835 0 1
rlabel polysilicon 1836 -2841 1836 -2841 0 3
rlabel polysilicon 1843 -2835 1843 -2835 0 1
rlabel polysilicon 1843 -2841 1843 -2841 0 3
rlabel polysilicon 1850 -2835 1850 -2835 0 1
rlabel polysilicon 1850 -2841 1850 -2841 0 3
rlabel polysilicon 1857 -2835 1857 -2835 0 1
rlabel polysilicon 1857 -2841 1857 -2841 0 3
rlabel polysilicon 1864 -2835 1864 -2835 0 1
rlabel polysilicon 1864 -2841 1864 -2841 0 3
rlabel polysilicon 1871 -2835 1871 -2835 0 1
rlabel polysilicon 1871 -2841 1871 -2841 0 3
rlabel polysilicon 1878 -2835 1878 -2835 0 1
rlabel polysilicon 1878 -2841 1878 -2841 0 3
rlabel polysilicon 1885 -2835 1885 -2835 0 1
rlabel polysilicon 1885 -2841 1885 -2841 0 3
rlabel polysilicon 1892 -2835 1892 -2835 0 1
rlabel polysilicon 1892 -2841 1892 -2841 0 3
rlabel polysilicon 1899 -2835 1899 -2835 0 1
rlabel polysilicon 1899 -2841 1899 -2841 0 3
rlabel polysilicon 1906 -2835 1906 -2835 0 1
rlabel polysilicon 1906 -2841 1906 -2841 0 3
rlabel polysilicon 1913 -2835 1913 -2835 0 1
rlabel polysilicon 1913 -2841 1913 -2841 0 3
rlabel polysilicon 1920 -2835 1920 -2835 0 1
rlabel polysilicon 1920 -2841 1920 -2841 0 3
rlabel polysilicon 1927 -2835 1927 -2835 0 1
rlabel polysilicon 1927 -2841 1927 -2841 0 3
rlabel polysilicon 1934 -2835 1934 -2835 0 1
rlabel polysilicon 1934 -2841 1934 -2841 0 3
rlabel polysilicon 1941 -2835 1941 -2835 0 1
rlabel polysilicon 1941 -2841 1941 -2841 0 3
rlabel polysilicon 1948 -2835 1948 -2835 0 1
rlabel polysilicon 1948 -2841 1948 -2841 0 3
rlabel polysilicon 1955 -2835 1955 -2835 0 1
rlabel polysilicon 1955 -2841 1955 -2841 0 3
rlabel polysilicon 1962 -2835 1962 -2835 0 1
rlabel polysilicon 1962 -2841 1962 -2841 0 3
rlabel polysilicon 1969 -2835 1969 -2835 0 1
rlabel polysilicon 1969 -2841 1969 -2841 0 3
rlabel polysilicon 1976 -2835 1976 -2835 0 1
rlabel polysilicon 1976 -2841 1976 -2841 0 3
rlabel polysilicon 1983 -2835 1983 -2835 0 1
rlabel polysilicon 1983 -2841 1983 -2841 0 3
rlabel polysilicon 1990 -2835 1990 -2835 0 1
rlabel polysilicon 1990 -2841 1990 -2841 0 3
rlabel polysilicon 1997 -2835 1997 -2835 0 1
rlabel polysilicon 1997 -2841 1997 -2841 0 3
rlabel polysilicon 2004 -2835 2004 -2835 0 1
rlabel polysilicon 2004 -2841 2004 -2841 0 3
rlabel polysilicon 2011 -2835 2011 -2835 0 1
rlabel polysilicon 2011 -2841 2011 -2841 0 3
rlabel polysilicon 2018 -2835 2018 -2835 0 1
rlabel polysilicon 2018 -2841 2018 -2841 0 3
rlabel polysilicon 2025 -2835 2025 -2835 0 1
rlabel polysilicon 2025 -2841 2025 -2841 0 3
rlabel polysilicon 2032 -2835 2032 -2835 0 1
rlabel polysilicon 2032 -2841 2032 -2841 0 3
rlabel polysilicon 2039 -2835 2039 -2835 0 1
rlabel polysilicon 2039 -2841 2039 -2841 0 3
rlabel polysilicon 2046 -2835 2046 -2835 0 1
rlabel polysilicon 2046 -2841 2046 -2841 0 3
rlabel polysilicon 2053 -2835 2053 -2835 0 1
rlabel polysilicon 2053 -2841 2053 -2841 0 3
rlabel polysilicon 2060 -2835 2060 -2835 0 1
rlabel polysilicon 2060 -2841 2060 -2841 0 3
rlabel polysilicon 2067 -2835 2067 -2835 0 1
rlabel polysilicon 2067 -2841 2067 -2841 0 3
rlabel polysilicon 2074 -2835 2074 -2835 0 1
rlabel polysilicon 2074 -2841 2074 -2841 0 3
rlabel polysilicon 2081 -2835 2081 -2835 0 1
rlabel polysilicon 2081 -2841 2081 -2841 0 3
rlabel polysilicon 2088 -2835 2088 -2835 0 1
rlabel polysilicon 2088 -2841 2088 -2841 0 3
rlabel polysilicon 2095 -2835 2095 -2835 0 1
rlabel polysilicon 2095 -2841 2095 -2841 0 3
rlabel polysilicon 2102 -2835 2102 -2835 0 1
rlabel polysilicon 2102 -2841 2102 -2841 0 3
rlabel polysilicon 2109 -2835 2109 -2835 0 1
rlabel polysilicon 2109 -2841 2109 -2841 0 3
rlabel polysilicon 2116 -2835 2116 -2835 0 1
rlabel polysilicon 2116 -2841 2116 -2841 0 3
rlabel polysilicon 2123 -2835 2123 -2835 0 1
rlabel polysilicon 2123 -2841 2123 -2841 0 3
rlabel polysilicon 2130 -2835 2130 -2835 0 1
rlabel polysilicon 2130 -2841 2130 -2841 0 3
rlabel polysilicon 2137 -2835 2137 -2835 0 1
rlabel polysilicon 2137 -2841 2137 -2841 0 3
rlabel polysilicon 2144 -2835 2144 -2835 0 1
rlabel polysilicon 2144 -2841 2144 -2841 0 3
rlabel polysilicon 2151 -2835 2151 -2835 0 1
rlabel polysilicon 2151 -2841 2151 -2841 0 3
rlabel polysilicon 2158 -2835 2158 -2835 0 1
rlabel polysilicon 2158 -2841 2158 -2841 0 3
rlabel polysilicon 2165 -2835 2165 -2835 0 1
rlabel polysilicon 2165 -2841 2165 -2841 0 3
rlabel polysilicon 2172 -2835 2172 -2835 0 1
rlabel polysilicon 2172 -2841 2172 -2841 0 3
rlabel polysilicon 2179 -2835 2179 -2835 0 1
rlabel polysilicon 2179 -2841 2179 -2841 0 3
rlabel polysilicon 2186 -2835 2186 -2835 0 1
rlabel polysilicon 2186 -2841 2186 -2841 0 3
rlabel polysilicon 2193 -2835 2193 -2835 0 1
rlabel polysilicon 2193 -2841 2193 -2841 0 3
rlabel polysilicon 2200 -2835 2200 -2835 0 1
rlabel polysilicon 2200 -2841 2200 -2841 0 3
rlabel polysilicon 2207 -2835 2207 -2835 0 1
rlabel polysilicon 2207 -2841 2207 -2841 0 3
rlabel polysilicon 2214 -2835 2214 -2835 0 1
rlabel polysilicon 2214 -2841 2214 -2841 0 3
rlabel polysilicon 2221 -2835 2221 -2835 0 1
rlabel polysilicon 2224 -2835 2224 -2835 0 2
rlabel polysilicon 2221 -2841 2221 -2841 0 3
rlabel polysilicon 2224 -2841 2224 -2841 0 4
rlabel polysilicon 2228 -2835 2228 -2835 0 1
rlabel polysilicon 2228 -2841 2228 -2841 0 3
rlabel polysilicon 2235 -2835 2235 -2835 0 1
rlabel polysilicon 2235 -2841 2235 -2841 0 3
rlabel polysilicon 2242 -2835 2242 -2835 0 1
rlabel polysilicon 2242 -2841 2242 -2841 0 3
rlabel polysilicon 2249 -2835 2249 -2835 0 1
rlabel polysilicon 2249 -2841 2249 -2841 0 3
rlabel polysilicon 2259 -2835 2259 -2835 0 2
rlabel polysilicon 2256 -2841 2256 -2841 0 3
rlabel polysilicon 2259 -2841 2259 -2841 0 4
rlabel polysilicon 2263 -2835 2263 -2835 0 1
rlabel polysilicon 2263 -2841 2263 -2841 0 3
rlabel polysilicon 2270 -2835 2270 -2835 0 1
rlabel polysilicon 2270 -2841 2270 -2841 0 3
rlabel polysilicon 16 -2980 16 -2980 0 1
rlabel polysilicon 16 -2986 16 -2986 0 3
rlabel polysilicon 23 -2980 23 -2980 0 1
rlabel polysilicon 23 -2986 23 -2986 0 3
rlabel polysilicon 30 -2980 30 -2980 0 1
rlabel polysilicon 30 -2986 30 -2986 0 3
rlabel polysilicon 37 -2980 37 -2980 0 1
rlabel polysilicon 37 -2986 37 -2986 0 3
rlabel polysilicon 44 -2980 44 -2980 0 1
rlabel polysilicon 44 -2986 44 -2986 0 3
rlabel polysilicon 54 -2980 54 -2980 0 2
rlabel polysilicon 51 -2986 51 -2986 0 3
rlabel polysilicon 58 -2980 58 -2980 0 1
rlabel polysilicon 58 -2986 58 -2986 0 3
rlabel polysilicon 65 -2980 65 -2980 0 1
rlabel polysilicon 65 -2986 65 -2986 0 3
rlabel polysilicon 72 -2980 72 -2980 0 1
rlabel polysilicon 72 -2986 72 -2986 0 3
rlabel polysilicon 79 -2980 79 -2980 0 1
rlabel polysilicon 79 -2986 79 -2986 0 3
rlabel polysilicon 86 -2980 86 -2980 0 1
rlabel polysilicon 86 -2986 86 -2986 0 3
rlabel polysilicon 93 -2980 93 -2980 0 1
rlabel polysilicon 93 -2986 93 -2986 0 3
rlabel polysilicon 100 -2980 100 -2980 0 1
rlabel polysilicon 103 -2980 103 -2980 0 2
rlabel polysilicon 100 -2986 100 -2986 0 3
rlabel polysilicon 103 -2986 103 -2986 0 4
rlabel polysilicon 110 -2980 110 -2980 0 2
rlabel polysilicon 110 -2986 110 -2986 0 4
rlabel polysilicon 114 -2980 114 -2980 0 1
rlabel polysilicon 117 -2980 117 -2980 0 2
rlabel polysilicon 117 -2986 117 -2986 0 4
rlabel polysilicon 121 -2980 121 -2980 0 1
rlabel polysilicon 124 -2980 124 -2980 0 2
rlabel polysilicon 121 -2986 121 -2986 0 3
rlabel polysilicon 124 -2986 124 -2986 0 4
rlabel polysilicon 128 -2980 128 -2980 0 1
rlabel polysilicon 128 -2986 128 -2986 0 3
rlabel polysilicon 135 -2980 135 -2980 0 1
rlabel polysilicon 135 -2986 135 -2986 0 3
rlabel polysilicon 142 -2980 142 -2980 0 1
rlabel polysilicon 142 -2986 142 -2986 0 3
rlabel polysilicon 149 -2980 149 -2980 0 1
rlabel polysilicon 149 -2986 149 -2986 0 3
rlabel polysilicon 159 -2980 159 -2980 0 2
rlabel polysilicon 156 -2986 156 -2986 0 3
rlabel polysilicon 159 -2986 159 -2986 0 4
rlabel polysilicon 163 -2980 163 -2980 0 1
rlabel polysilicon 163 -2986 163 -2986 0 3
rlabel polysilicon 170 -2980 170 -2980 0 1
rlabel polysilicon 170 -2986 170 -2986 0 3
rlabel polysilicon 177 -2980 177 -2980 0 1
rlabel polysilicon 177 -2986 177 -2986 0 3
rlabel polysilicon 184 -2980 184 -2980 0 1
rlabel polysilicon 184 -2986 184 -2986 0 3
rlabel polysilicon 191 -2980 191 -2980 0 1
rlabel polysilicon 191 -2986 191 -2986 0 3
rlabel polysilicon 198 -2980 198 -2980 0 1
rlabel polysilicon 198 -2986 198 -2986 0 3
rlabel polysilicon 205 -2980 205 -2980 0 1
rlabel polysilicon 205 -2986 205 -2986 0 3
rlabel polysilicon 212 -2980 212 -2980 0 1
rlabel polysilicon 215 -2980 215 -2980 0 2
rlabel polysilicon 212 -2986 212 -2986 0 3
rlabel polysilicon 215 -2986 215 -2986 0 4
rlabel polysilicon 219 -2980 219 -2980 0 1
rlabel polysilicon 219 -2986 219 -2986 0 3
rlabel polysilicon 226 -2980 226 -2980 0 1
rlabel polysilicon 226 -2986 226 -2986 0 3
rlabel polysilicon 233 -2980 233 -2980 0 1
rlabel polysilicon 233 -2986 233 -2986 0 3
rlabel polysilicon 240 -2980 240 -2980 0 1
rlabel polysilicon 240 -2986 240 -2986 0 3
rlabel polysilicon 247 -2980 247 -2980 0 1
rlabel polysilicon 247 -2986 247 -2986 0 3
rlabel polysilicon 254 -2980 254 -2980 0 1
rlabel polysilicon 257 -2980 257 -2980 0 2
rlabel polysilicon 254 -2986 254 -2986 0 3
rlabel polysilicon 261 -2980 261 -2980 0 1
rlabel polysilicon 261 -2986 261 -2986 0 3
rlabel polysilicon 268 -2980 268 -2980 0 1
rlabel polysilicon 268 -2986 268 -2986 0 3
rlabel polysilicon 275 -2980 275 -2980 0 1
rlabel polysilicon 275 -2986 275 -2986 0 3
rlabel polysilicon 282 -2980 282 -2980 0 1
rlabel polysilicon 282 -2986 282 -2986 0 3
rlabel polysilicon 289 -2980 289 -2980 0 1
rlabel polysilicon 289 -2986 289 -2986 0 3
rlabel polysilicon 296 -2980 296 -2980 0 1
rlabel polysilicon 296 -2986 296 -2986 0 3
rlabel polysilicon 303 -2980 303 -2980 0 1
rlabel polysilicon 303 -2986 303 -2986 0 3
rlabel polysilicon 310 -2980 310 -2980 0 1
rlabel polysilicon 310 -2986 310 -2986 0 3
rlabel polysilicon 317 -2980 317 -2980 0 1
rlabel polysilicon 317 -2986 317 -2986 0 3
rlabel polysilicon 324 -2980 324 -2980 0 1
rlabel polysilicon 324 -2986 324 -2986 0 3
rlabel polysilicon 331 -2980 331 -2980 0 1
rlabel polysilicon 331 -2986 331 -2986 0 3
rlabel polysilicon 338 -2980 338 -2980 0 1
rlabel polysilicon 338 -2986 338 -2986 0 3
rlabel polysilicon 345 -2980 345 -2980 0 1
rlabel polysilicon 345 -2986 345 -2986 0 3
rlabel polysilicon 352 -2980 352 -2980 0 1
rlabel polysilicon 352 -2986 352 -2986 0 3
rlabel polysilicon 359 -2980 359 -2980 0 1
rlabel polysilicon 359 -2986 359 -2986 0 3
rlabel polysilicon 366 -2980 366 -2980 0 1
rlabel polysilicon 366 -2986 366 -2986 0 3
rlabel polysilicon 373 -2980 373 -2980 0 1
rlabel polysilicon 373 -2986 373 -2986 0 3
rlabel polysilicon 380 -2980 380 -2980 0 1
rlabel polysilicon 380 -2986 380 -2986 0 3
rlabel polysilicon 387 -2980 387 -2980 0 1
rlabel polysilicon 387 -2986 387 -2986 0 3
rlabel polysilicon 394 -2980 394 -2980 0 1
rlabel polysilicon 394 -2986 394 -2986 0 3
rlabel polysilicon 401 -2980 401 -2980 0 1
rlabel polysilicon 401 -2986 401 -2986 0 3
rlabel polysilicon 408 -2980 408 -2980 0 1
rlabel polysilicon 408 -2986 408 -2986 0 3
rlabel polysilicon 415 -2980 415 -2980 0 1
rlabel polysilicon 415 -2986 415 -2986 0 3
rlabel polysilicon 422 -2980 422 -2980 0 1
rlabel polysilicon 422 -2986 422 -2986 0 3
rlabel polysilicon 429 -2980 429 -2980 0 1
rlabel polysilicon 429 -2986 429 -2986 0 3
rlabel polysilicon 436 -2980 436 -2980 0 1
rlabel polysilicon 436 -2986 436 -2986 0 3
rlabel polysilicon 443 -2980 443 -2980 0 1
rlabel polysilicon 443 -2986 443 -2986 0 3
rlabel polysilicon 450 -2980 450 -2980 0 1
rlabel polysilicon 450 -2986 450 -2986 0 3
rlabel polysilicon 457 -2980 457 -2980 0 1
rlabel polysilicon 457 -2986 457 -2986 0 3
rlabel polysilicon 464 -2980 464 -2980 0 1
rlabel polysilicon 467 -2980 467 -2980 0 2
rlabel polysilicon 471 -2980 471 -2980 0 1
rlabel polysilicon 471 -2986 471 -2986 0 3
rlabel polysilicon 478 -2980 478 -2980 0 1
rlabel polysilicon 478 -2986 478 -2986 0 3
rlabel polysilicon 485 -2980 485 -2980 0 1
rlabel polysilicon 485 -2986 485 -2986 0 3
rlabel polysilicon 492 -2980 492 -2980 0 1
rlabel polysilicon 492 -2986 492 -2986 0 3
rlabel polysilicon 499 -2980 499 -2980 0 1
rlabel polysilicon 499 -2986 499 -2986 0 3
rlabel polysilicon 506 -2980 506 -2980 0 1
rlabel polysilicon 506 -2986 506 -2986 0 3
rlabel polysilicon 513 -2980 513 -2980 0 1
rlabel polysilicon 513 -2986 513 -2986 0 3
rlabel polysilicon 520 -2980 520 -2980 0 1
rlabel polysilicon 520 -2986 520 -2986 0 3
rlabel polysilicon 527 -2980 527 -2980 0 1
rlabel polysilicon 527 -2986 527 -2986 0 3
rlabel polysilicon 534 -2980 534 -2980 0 1
rlabel polysilicon 534 -2986 534 -2986 0 3
rlabel polysilicon 541 -2980 541 -2980 0 1
rlabel polysilicon 544 -2980 544 -2980 0 2
rlabel polysilicon 541 -2986 541 -2986 0 3
rlabel polysilicon 544 -2986 544 -2986 0 4
rlabel polysilicon 548 -2980 548 -2980 0 1
rlabel polysilicon 548 -2986 548 -2986 0 3
rlabel polysilicon 555 -2980 555 -2980 0 1
rlabel polysilicon 555 -2986 555 -2986 0 3
rlabel polysilicon 562 -2980 562 -2980 0 1
rlabel polysilicon 565 -2980 565 -2980 0 2
rlabel polysilicon 565 -2986 565 -2986 0 4
rlabel polysilicon 569 -2980 569 -2980 0 1
rlabel polysilicon 569 -2986 569 -2986 0 3
rlabel polysilicon 572 -2986 572 -2986 0 4
rlabel polysilicon 576 -2980 576 -2980 0 1
rlabel polysilicon 576 -2986 576 -2986 0 3
rlabel polysilicon 583 -2980 583 -2980 0 1
rlabel polysilicon 583 -2986 583 -2986 0 3
rlabel polysilicon 590 -2980 590 -2980 0 1
rlabel polysilicon 590 -2986 590 -2986 0 3
rlabel polysilicon 597 -2980 597 -2980 0 1
rlabel polysilicon 597 -2986 597 -2986 0 3
rlabel polysilicon 604 -2980 604 -2980 0 1
rlabel polysilicon 604 -2986 604 -2986 0 3
rlabel polysilicon 611 -2980 611 -2980 0 1
rlabel polysilicon 611 -2986 611 -2986 0 3
rlabel polysilicon 618 -2980 618 -2980 0 1
rlabel polysilicon 618 -2986 618 -2986 0 3
rlabel polysilicon 625 -2980 625 -2980 0 1
rlabel polysilicon 625 -2986 625 -2986 0 3
rlabel polysilicon 632 -2980 632 -2980 0 1
rlabel polysilicon 632 -2986 632 -2986 0 3
rlabel polysilicon 639 -2980 639 -2980 0 1
rlabel polysilicon 642 -2980 642 -2980 0 2
rlabel polysilicon 642 -2986 642 -2986 0 4
rlabel polysilicon 646 -2980 646 -2980 0 1
rlabel polysilicon 646 -2986 646 -2986 0 3
rlabel polysilicon 653 -2980 653 -2980 0 1
rlabel polysilicon 653 -2986 653 -2986 0 3
rlabel polysilicon 660 -2980 660 -2980 0 1
rlabel polysilicon 663 -2980 663 -2980 0 2
rlabel polysilicon 660 -2986 660 -2986 0 3
rlabel polysilicon 663 -2986 663 -2986 0 4
rlabel polysilicon 667 -2980 667 -2980 0 1
rlabel polysilicon 667 -2986 667 -2986 0 3
rlabel polysilicon 674 -2980 674 -2980 0 1
rlabel polysilicon 674 -2986 674 -2986 0 3
rlabel polysilicon 681 -2980 681 -2980 0 1
rlabel polysilicon 681 -2986 681 -2986 0 3
rlabel polysilicon 688 -2980 688 -2980 0 1
rlabel polysilicon 688 -2986 688 -2986 0 3
rlabel polysilicon 695 -2980 695 -2980 0 1
rlabel polysilicon 695 -2986 695 -2986 0 3
rlabel polysilicon 702 -2980 702 -2980 0 1
rlabel polysilicon 702 -2986 702 -2986 0 3
rlabel polysilicon 709 -2980 709 -2980 0 1
rlabel polysilicon 709 -2986 709 -2986 0 3
rlabel polysilicon 716 -2980 716 -2980 0 1
rlabel polysilicon 716 -2986 716 -2986 0 3
rlabel polysilicon 723 -2980 723 -2980 0 1
rlabel polysilicon 723 -2986 723 -2986 0 3
rlabel polysilicon 730 -2980 730 -2980 0 1
rlabel polysilicon 730 -2986 730 -2986 0 3
rlabel polysilicon 737 -2980 737 -2980 0 1
rlabel polysilicon 740 -2980 740 -2980 0 2
rlabel polysilicon 737 -2986 737 -2986 0 3
rlabel polysilicon 740 -2986 740 -2986 0 4
rlabel polysilicon 744 -2980 744 -2980 0 1
rlabel polysilicon 744 -2986 744 -2986 0 3
rlabel polysilicon 751 -2980 751 -2980 0 1
rlabel polysilicon 751 -2986 751 -2986 0 3
rlabel polysilicon 758 -2980 758 -2980 0 1
rlabel polysilicon 758 -2986 758 -2986 0 3
rlabel polysilicon 765 -2980 765 -2980 0 1
rlabel polysilicon 765 -2986 765 -2986 0 3
rlabel polysilicon 772 -2980 772 -2980 0 1
rlabel polysilicon 772 -2986 772 -2986 0 3
rlabel polysilicon 779 -2980 779 -2980 0 1
rlabel polysilicon 779 -2986 779 -2986 0 3
rlabel polysilicon 786 -2980 786 -2980 0 1
rlabel polysilicon 786 -2986 786 -2986 0 3
rlabel polysilicon 793 -2980 793 -2980 0 1
rlabel polysilicon 793 -2986 793 -2986 0 3
rlabel polysilicon 800 -2980 800 -2980 0 1
rlabel polysilicon 807 -2980 807 -2980 0 1
rlabel polysilicon 807 -2986 807 -2986 0 3
rlabel polysilicon 814 -2980 814 -2980 0 1
rlabel polysilicon 814 -2986 814 -2986 0 3
rlabel polysilicon 821 -2980 821 -2980 0 1
rlabel polysilicon 821 -2986 821 -2986 0 3
rlabel polysilicon 828 -2980 828 -2980 0 1
rlabel polysilicon 828 -2986 828 -2986 0 3
rlabel polysilicon 835 -2980 835 -2980 0 1
rlabel polysilicon 835 -2986 835 -2986 0 3
rlabel polysilicon 842 -2980 842 -2980 0 1
rlabel polysilicon 842 -2986 842 -2986 0 3
rlabel polysilicon 849 -2980 849 -2980 0 1
rlabel polysilicon 849 -2986 849 -2986 0 3
rlabel polysilicon 856 -2980 856 -2980 0 1
rlabel polysilicon 856 -2986 856 -2986 0 3
rlabel polysilicon 863 -2980 863 -2980 0 1
rlabel polysilicon 863 -2986 863 -2986 0 3
rlabel polysilicon 870 -2980 870 -2980 0 1
rlabel polysilicon 870 -2986 870 -2986 0 3
rlabel polysilicon 880 -2980 880 -2980 0 2
rlabel polysilicon 880 -2986 880 -2986 0 4
rlabel polysilicon 884 -2980 884 -2980 0 1
rlabel polysilicon 884 -2986 884 -2986 0 3
rlabel polysilicon 891 -2980 891 -2980 0 1
rlabel polysilicon 891 -2986 891 -2986 0 3
rlabel polysilicon 898 -2980 898 -2980 0 1
rlabel polysilicon 898 -2986 898 -2986 0 3
rlabel polysilicon 905 -2980 905 -2980 0 1
rlabel polysilicon 905 -2986 905 -2986 0 3
rlabel polysilicon 912 -2980 912 -2980 0 1
rlabel polysilicon 912 -2986 912 -2986 0 3
rlabel polysilicon 922 -2980 922 -2980 0 2
rlabel polysilicon 919 -2986 919 -2986 0 3
rlabel polysilicon 922 -2986 922 -2986 0 4
rlabel polysilicon 926 -2980 926 -2980 0 1
rlabel polysilicon 926 -2986 926 -2986 0 3
rlabel polysilicon 933 -2980 933 -2980 0 1
rlabel polysilicon 933 -2986 933 -2986 0 3
rlabel polysilicon 940 -2980 940 -2980 0 1
rlabel polysilicon 940 -2986 940 -2986 0 3
rlabel polysilicon 947 -2980 947 -2980 0 1
rlabel polysilicon 947 -2986 947 -2986 0 3
rlabel polysilicon 954 -2980 954 -2980 0 1
rlabel polysilicon 954 -2986 954 -2986 0 3
rlabel polysilicon 961 -2980 961 -2980 0 1
rlabel polysilicon 964 -2980 964 -2980 0 2
rlabel polysilicon 961 -2986 961 -2986 0 3
rlabel polysilicon 964 -2986 964 -2986 0 4
rlabel polysilicon 968 -2980 968 -2980 0 1
rlabel polysilicon 968 -2986 968 -2986 0 3
rlabel polysilicon 975 -2980 975 -2980 0 1
rlabel polysilicon 975 -2986 975 -2986 0 3
rlabel polysilicon 982 -2980 982 -2980 0 1
rlabel polysilicon 985 -2980 985 -2980 0 2
rlabel polysilicon 982 -2986 982 -2986 0 3
rlabel polysilicon 985 -2986 985 -2986 0 4
rlabel polysilicon 989 -2980 989 -2980 0 1
rlabel polysilicon 989 -2986 989 -2986 0 3
rlabel polysilicon 996 -2980 996 -2980 0 1
rlabel polysilicon 996 -2986 996 -2986 0 3
rlabel polysilicon 1003 -2980 1003 -2980 0 1
rlabel polysilicon 1003 -2986 1003 -2986 0 3
rlabel polysilicon 1010 -2980 1010 -2980 0 1
rlabel polysilicon 1010 -2986 1010 -2986 0 3
rlabel polysilicon 1017 -2980 1017 -2980 0 1
rlabel polysilicon 1017 -2986 1017 -2986 0 3
rlabel polysilicon 1024 -2980 1024 -2980 0 1
rlabel polysilicon 1024 -2986 1024 -2986 0 3
rlabel polysilicon 1031 -2980 1031 -2980 0 1
rlabel polysilicon 1031 -2986 1031 -2986 0 3
rlabel polysilicon 1034 -2986 1034 -2986 0 4
rlabel polysilicon 1038 -2980 1038 -2980 0 1
rlabel polysilicon 1041 -2980 1041 -2980 0 2
rlabel polysilicon 1038 -2986 1038 -2986 0 3
rlabel polysilicon 1041 -2986 1041 -2986 0 4
rlabel polysilicon 1045 -2980 1045 -2980 0 1
rlabel polysilicon 1045 -2986 1045 -2986 0 3
rlabel polysilicon 1055 -2980 1055 -2980 0 2
rlabel polysilicon 1052 -2986 1052 -2986 0 3
rlabel polysilicon 1055 -2986 1055 -2986 0 4
rlabel polysilicon 1059 -2980 1059 -2980 0 1
rlabel polysilicon 1062 -2980 1062 -2980 0 2
rlabel polysilicon 1059 -2986 1059 -2986 0 3
rlabel polysilicon 1062 -2986 1062 -2986 0 4
rlabel polysilicon 1066 -2980 1066 -2980 0 1
rlabel polysilicon 1069 -2980 1069 -2980 0 2
rlabel polysilicon 1066 -2986 1066 -2986 0 3
rlabel polysilicon 1069 -2986 1069 -2986 0 4
rlabel polysilicon 1073 -2980 1073 -2980 0 1
rlabel polysilicon 1073 -2986 1073 -2986 0 3
rlabel polysilicon 1080 -2980 1080 -2980 0 1
rlabel polysilicon 1080 -2986 1080 -2986 0 3
rlabel polysilicon 1087 -2980 1087 -2980 0 1
rlabel polysilicon 1087 -2986 1087 -2986 0 3
rlabel polysilicon 1094 -2980 1094 -2980 0 1
rlabel polysilicon 1097 -2980 1097 -2980 0 2
rlabel polysilicon 1097 -2986 1097 -2986 0 4
rlabel polysilicon 1101 -2980 1101 -2980 0 1
rlabel polysilicon 1101 -2986 1101 -2986 0 3
rlabel polysilicon 1108 -2980 1108 -2980 0 1
rlabel polysilicon 1108 -2986 1108 -2986 0 3
rlabel polysilicon 1115 -2980 1115 -2980 0 1
rlabel polysilicon 1115 -2986 1115 -2986 0 3
rlabel polysilicon 1122 -2980 1122 -2980 0 1
rlabel polysilicon 1125 -2980 1125 -2980 0 2
rlabel polysilicon 1125 -2986 1125 -2986 0 4
rlabel polysilicon 1129 -2980 1129 -2980 0 1
rlabel polysilicon 1129 -2986 1129 -2986 0 3
rlabel polysilicon 1136 -2980 1136 -2980 0 1
rlabel polysilicon 1139 -2980 1139 -2980 0 2
rlabel polysilicon 1136 -2986 1136 -2986 0 3
rlabel polysilicon 1139 -2986 1139 -2986 0 4
rlabel polysilicon 1143 -2980 1143 -2980 0 1
rlabel polysilicon 1143 -2986 1143 -2986 0 3
rlabel polysilicon 1150 -2980 1150 -2980 0 1
rlabel polysilicon 1150 -2986 1150 -2986 0 3
rlabel polysilicon 1157 -2980 1157 -2980 0 1
rlabel polysilicon 1160 -2980 1160 -2980 0 2
rlabel polysilicon 1157 -2986 1157 -2986 0 3
rlabel polysilicon 1160 -2986 1160 -2986 0 4
rlabel polysilicon 1164 -2980 1164 -2980 0 1
rlabel polysilicon 1164 -2986 1164 -2986 0 3
rlabel polysilicon 1171 -2980 1171 -2980 0 1
rlabel polysilicon 1171 -2986 1171 -2986 0 3
rlabel polysilicon 1178 -2980 1178 -2980 0 1
rlabel polysilicon 1178 -2986 1178 -2986 0 3
rlabel polysilicon 1185 -2980 1185 -2980 0 1
rlabel polysilicon 1185 -2986 1185 -2986 0 3
rlabel polysilicon 1192 -2980 1192 -2980 0 1
rlabel polysilicon 1192 -2986 1192 -2986 0 3
rlabel polysilicon 1199 -2980 1199 -2980 0 1
rlabel polysilicon 1202 -2980 1202 -2980 0 2
rlabel polysilicon 1199 -2986 1199 -2986 0 3
rlabel polysilicon 1202 -2986 1202 -2986 0 4
rlabel polysilicon 1206 -2980 1206 -2980 0 1
rlabel polysilicon 1209 -2980 1209 -2980 0 2
rlabel polysilicon 1209 -2986 1209 -2986 0 4
rlabel polysilicon 1213 -2980 1213 -2980 0 1
rlabel polysilicon 1213 -2986 1213 -2986 0 3
rlabel polysilicon 1220 -2980 1220 -2980 0 1
rlabel polysilicon 1220 -2986 1220 -2986 0 3
rlabel polysilicon 1227 -2980 1227 -2980 0 1
rlabel polysilicon 1227 -2986 1227 -2986 0 3
rlabel polysilicon 1234 -2980 1234 -2980 0 1
rlabel polysilicon 1234 -2986 1234 -2986 0 3
rlabel polysilicon 1241 -2980 1241 -2980 0 1
rlabel polysilicon 1241 -2986 1241 -2986 0 3
rlabel polysilicon 1248 -2980 1248 -2980 0 1
rlabel polysilicon 1248 -2986 1248 -2986 0 3
rlabel polysilicon 1255 -2980 1255 -2980 0 1
rlabel polysilicon 1255 -2986 1255 -2986 0 3
rlabel polysilicon 1262 -2980 1262 -2980 0 1
rlabel polysilicon 1262 -2986 1262 -2986 0 3
rlabel polysilicon 1269 -2980 1269 -2980 0 1
rlabel polysilicon 1269 -2986 1269 -2986 0 3
rlabel polysilicon 1276 -2980 1276 -2980 0 1
rlabel polysilicon 1276 -2986 1276 -2986 0 3
rlabel polysilicon 1283 -2980 1283 -2980 0 1
rlabel polysilicon 1283 -2986 1283 -2986 0 3
rlabel polysilicon 1290 -2980 1290 -2980 0 1
rlabel polysilicon 1290 -2986 1290 -2986 0 3
rlabel polysilicon 1297 -2980 1297 -2980 0 1
rlabel polysilicon 1297 -2986 1297 -2986 0 3
rlabel polysilicon 1304 -2980 1304 -2980 0 1
rlabel polysilicon 1304 -2986 1304 -2986 0 3
rlabel polysilicon 1314 -2980 1314 -2980 0 2
rlabel polysilicon 1311 -2986 1311 -2986 0 3
rlabel polysilicon 1314 -2986 1314 -2986 0 4
rlabel polysilicon 1318 -2980 1318 -2980 0 1
rlabel polysilicon 1318 -2986 1318 -2986 0 3
rlabel polysilicon 1325 -2980 1325 -2980 0 1
rlabel polysilicon 1325 -2986 1325 -2986 0 3
rlabel polysilicon 1332 -2980 1332 -2980 0 1
rlabel polysilicon 1332 -2986 1332 -2986 0 3
rlabel polysilicon 1339 -2980 1339 -2980 0 1
rlabel polysilicon 1339 -2986 1339 -2986 0 3
rlabel polysilicon 1346 -2980 1346 -2980 0 1
rlabel polysilicon 1346 -2986 1346 -2986 0 3
rlabel polysilicon 1353 -2980 1353 -2980 0 1
rlabel polysilicon 1353 -2986 1353 -2986 0 3
rlabel polysilicon 1360 -2980 1360 -2980 0 1
rlabel polysilicon 1363 -2980 1363 -2980 0 2
rlabel polysilicon 1363 -2986 1363 -2986 0 4
rlabel polysilicon 1367 -2980 1367 -2980 0 1
rlabel polysilicon 1367 -2986 1367 -2986 0 3
rlabel polysilicon 1374 -2980 1374 -2980 0 1
rlabel polysilicon 1374 -2986 1374 -2986 0 3
rlabel polysilicon 1381 -2980 1381 -2980 0 1
rlabel polysilicon 1381 -2986 1381 -2986 0 3
rlabel polysilicon 1388 -2980 1388 -2980 0 1
rlabel polysilicon 1388 -2986 1388 -2986 0 3
rlabel polysilicon 1395 -2980 1395 -2980 0 1
rlabel polysilicon 1395 -2986 1395 -2986 0 3
rlabel polysilicon 1402 -2980 1402 -2980 0 1
rlabel polysilicon 1402 -2986 1402 -2986 0 3
rlabel polysilicon 1409 -2980 1409 -2980 0 1
rlabel polysilicon 1409 -2986 1409 -2986 0 3
rlabel polysilicon 1419 -2980 1419 -2980 0 2
rlabel polysilicon 1416 -2986 1416 -2986 0 3
rlabel polysilicon 1419 -2986 1419 -2986 0 4
rlabel polysilicon 1423 -2980 1423 -2980 0 1
rlabel polysilicon 1423 -2986 1423 -2986 0 3
rlabel polysilicon 1430 -2980 1430 -2980 0 1
rlabel polysilicon 1430 -2986 1430 -2986 0 3
rlabel polysilicon 1437 -2980 1437 -2980 0 1
rlabel polysilicon 1437 -2986 1437 -2986 0 3
rlabel polysilicon 1444 -2980 1444 -2980 0 1
rlabel polysilicon 1444 -2986 1444 -2986 0 3
rlabel polysilicon 1451 -2980 1451 -2980 0 1
rlabel polysilicon 1451 -2986 1451 -2986 0 3
rlabel polysilicon 1458 -2980 1458 -2980 0 1
rlabel polysilicon 1458 -2986 1458 -2986 0 3
rlabel polysilicon 1465 -2980 1465 -2980 0 1
rlabel polysilicon 1465 -2986 1465 -2986 0 3
rlabel polysilicon 1472 -2980 1472 -2980 0 1
rlabel polysilicon 1472 -2986 1472 -2986 0 3
rlabel polysilicon 1479 -2980 1479 -2980 0 1
rlabel polysilicon 1479 -2986 1479 -2986 0 3
rlabel polysilicon 1486 -2980 1486 -2980 0 1
rlabel polysilicon 1486 -2986 1486 -2986 0 3
rlabel polysilicon 1493 -2980 1493 -2980 0 1
rlabel polysilicon 1493 -2986 1493 -2986 0 3
rlabel polysilicon 1500 -2980 1500 -2980 0 1
rlabel polysilicon 1500 -2986 1500 -2986 0 3
rlabel polysilicon 1507 -2980 1507 -2980 0 1
rlabel polysilicon 1507 -2986 1507 -2986 0 3
rlabel polysilicon 1514 -2980 1514 -2980 0 1
rlabel polysilicon 1514 -2986 1514 -2986 0 3
rlabel polysilicon 1521 -2980 1521 -2980 0 1
rlabel polysilicon 1521 -2986 1521 -2986 0 3
rlabel polysilicon 1528 -2980 1528 -2980 0 1
rlabel polysilicon 1528 -2986 1528 -2986 0 3
rlabel polysilicon 1535 -2980 1535 -2980 0 1
rlabel polysilicon 1535 -2986 1535 -2986 0 3
rlabel polysilicon 1542 -2980 1542 -2980 0 1
rlabel polysilicon 1542 -2986 1542 -2986 0 3
rlabel polysilicon 1549 -2980 1549 -2980 0 1
rlabel polysilicon 1549 -2986 1549 -2986 0 3
rlabel polysilicon 1556 -2980 1556 -2980 0 1
rlabel polysilicon 1556 -2986 1556 -2986 0 3
rlabel polysilicon 1563 -2980 1563 -2980 0 1
rlabel polysilicon 1563 -2986 1563 -2986 0 3
rlabel polysilicon 1570 -2980 1570 -2980 0 1
rlabel polysilicon 1570 -2986 1570 -2986 0 3
rlabel polysilicon 1573 -2986 1573 -2986 0 4
rlabel polysilicon 1577 -2980 1577 -2980 0 1
rlabel polysilicon 1577 -2986 1577 -2986 0 3
rlabel polysilicon 1584 -2980 1584 -2980 0 1
rlabel polysilicon 1584 -2986 1584 -2986 0 3
rlabel polysilicon 1591 -2980 1591 -2980 0 1
rlabel polysilicon 1591 -2986 1591 -2986 0 3
rlabel polysilicon 1598 -2980 1598 -2980 0 1
rlabel polysilicon 1598 -2986 1598 -2986 0 3
rlabel polysilicon 1605 -2980 1605 -2980 0 1
rlabel polysilicon 1605 -2986 1605 -2986 0 3
rlabel polysilicon 1612 -2980 1612 -2980 0 1
rlabel polysilicon 1612 -2986 1612 -2986 0 3
rlabel polysilicon 1619 -2980 1619 -2980 0 1
rlabel polysilicon 1619 -2986 1619 -2986 0 3
rlabel polysilicon 1626 -2980 1626 -2980 0 1
rlabel polysilicon 1626 -2986 1626 -2986 0 3
rlabel polysilicon 1633 -2980 1633 -2980 0 1
rlabel polysilicon 1633 -2986 1633 -2986 0 3
rlabel polysilicon 1640 -2980 1640 -2980 0 1
rlabel polysilicon 1640 -2986 1640 -2986 0 3
rlabel polysilicon 1647 -2980 1647 -2980 0 1
rlabel polysilicon 1647 -2986 1647 -2986 0 3
rlabel polysilicon 1654 -2980 1654 -2980 0 1
rlabel polysilicon 1654 -2986 1654 -2986 0 3
rlabel polysilicon 1661 -2980 1661 -2980 0 1
rlabel polysilicon 1661 -2986 1661 -2986 0 3
rlabel polysilicon 1668 -2980 1668 -2980 0 1
rlabel polysilicon 1668 -2986 1668 -2986 0 3
rlabel polysilicon 1675 -2980 1675 -2980 0 1
rlabel polysilicon 1675 -2986 1675 -2986 0 3
rlabel polysilicon 1682 -2980 1682 -2980 0 1
rlabel polysilicon 1682 -2986 1682 -2986 0 3
rlabel polysilicon 1689 -2980 1689 -2980 0 1
rlabel polysilicon 1689 -2986 1689 -2986 0 3
rlabel polysilicon 1696 -2980 1696 -2980 0 1
rlabel polysilicon 1696 -2986 1696 -2986 0 3
rlabel polysilicon 1703 -2980 1703 -2980 0 1
rlabel polysilicon 1703 -2986 1703 -2986 0 3
rlabel polysilicon 1710 -2980 1710 -2980 0 1
rlabel polysilicon 1710 -2986 1710 -2986 0 3
rlabel polysilicon 1717 -2980 1717 -2980 0 1
rlabel polysilicon 1717 -2986 1717 -2986 0 3
rlabel polysilicon 1724 -2980 1724 -2980 0 1
rlabel polysilicon 1724 -2986 1724 -2986 0 3
rlabel polysilicon 1731 -2980 1731 -2980 0 1
rlabel polysilicon 1731 -2986 1731 -2986 0 3
rlabel polysilicon 1738 -2980 1738 -2980 0 1
rlabel polysilicon 1738 -2986 1738 -2986 0 3
rlabel polysilicon 1745 -2980 1745 -2980 0 1
rlabel polysilicon 1745 -2986 1745 -2986 0 3
rlabel polysilicon 1752 -2980 1752 -2980 0 1
rlabel polysilicon 1752 -2986 1752 -2986 0 3
rlabel polysilicon 1759 -2980 1759 -2980 0 1
rlabel polysilicon 1759 -2986 1759 -2986 0 3
rlabel polysilicon 1766 -2986 1766 -2986 0 3
rlabel polysilicon 1769 -2986 1769 -2986 0 4
rlabel polysilicon 1773 -2980 1773 -2980 0 1
rlabel polysilicon 1773 -2986 1773 -2986 0 3
rlabel polysilicon 1780 -2980 1780 -2980 0 1
rlabel polysilicon 1780 -2986 1780 -2986 0 3
rlabel polysilicon 1787 -2980 1787 -2980 0 1
rlabel polysilicon 1787 -2986 1787 -2986 0 3
rlabel polysilicon 1794 -2980 1794 -2980 0 1
rlabel polysilicon 1794 -2986 1794 -2986 0 3
rlabel polysilicon 1801 -2980 1801 -2980 0 1
rlabel polysilicon 1801 -2986 1801 -2986 0 3
rlabel polysilicon 1808 -2980 1808 -2980 0 1
rlabel polysilicon 1808 -2986 1808 -2986 0 3
rlabel polysilicon 1815 -2980 1815 -2980 0 1
rlabel polysilicon 1815 -2986 1815 -2986 0 3
rlabel polysilicon 1822 -2980 1822 -2980 0 1
rlabel polysilicon 1822 -2986 1822 -2986 0 3
rlabel polysilicon 1829 -2980 1829 -2980 0 1
rlabel polysilicon 1829 -2986 1829 -2986 0 3
rlabel polysilicon 1836 -2980 1836 -2980 0 1
rlabel polysilicon 1836 -2986 1836 -2986 0 3
rlabel polysilicon 1843 -2980 1843 -2980 0 1
rlabel polysilicon 1843 -2986 1843 -2986 0 3
rlabel polysilicon 1850 -2980 1850 -2980 0 1
rlabel polysilicon 1850 -2986 1850 -2986 0 3
rlabel polysilicon 1857 -2980 1857 -2980 0 1
rlabel polysilicon 1857 -2986 1857 -2986 0 3
rlabel polysilicon 1864 -2980 1864 -2980 0 1
rlabel polysilicon 1864 -2986 1864 -2986 0 3
rlabel polysilicon 1871 -2980 1871 -2980 0 1
rlabel polysilicon 1871 -2986 1871 -2986 0 3
rlabel polysilicon 1874 -2986 1874 -2986 0 4
rlabel polysilicon 1878 -2980 1878 -2980 0 1
rlabel polysilicon 1878 -2986 1878 -2986 0 3
rlabel polysilicon 1885 -2980 1885 -2980 0 1
rlabel polysilicon 1885 -2986 1885 -2986 0 3
rlabel polysilicon 1892 -2980 1892 -2980 0 1
rlabel polysilicon 1892 -2986 1892 -2986 0 3
rlabel polysilicon 1899 -2980 1899 -2980 0 1
rlabel polysilicon 1899 -2986 1899 -2986 0 3
rlabel polysilicon 1906 -2980 1906 -2980 0 1
rlabel polysilicon 1906 -2986 1906 -2986 0 3
rlabel polysilicon 1913 -2980 1913 -2980 0 1
rlabel polysilicon 1913 -2986 1913 -2986 0 3
rlabel polysilicon 1920 -2980 1920 -2980 0 1
rlabel polysilicon 1920 -2986 1920 -2986 0 3
rlabel polysilicon 1927 -2980 1927 -2980 0 1
rlabel polysilicon 1927 -2986 1927 -2986 0 3
rlabel polysilicon 1934 -2980 1934 -2980 0 1
rlabel polysilicon 1934 -2986 1934 -2986 0 3
rlabel polysilicon 1941 -2980 1941 -2980 0 1
rlabel polysilicon 1941 -2986 1941 -2986 0 3
rlabel polysilicon 1948 -2980 1948 -2980 0 1
rlabel polysilicon 1948 -2986 1948 -2986 0 3
rlabel polysilicon 1955 -2980 1955 -2980 0 1
rlabel polysilicon 1955 -2986 1955 -2986 0 3
rlabel polysilicon 1962 -2980 1962 -2980 0 1
rlabel polysilicon 1962 -2986 1962 -2986 0 3
rlabel polysilicon 1969 -2980 1969 -2980 0 1
rlabel polysilicon 1969 -2986 1969 -2986 0 3
rlabel polysilicon 1976 -2980 1976 -2980 0 1
rlabel polysilicon 1976 -2986 1976 -2986 0 3
rlabel polysilicon 1983 -2980 1983 -2980 0 1
rlabel polysilicon 1983 -2986 1983 -2986 0 3
rlabel polysilicon 1990 -2980 1990 -2980 0 1
rlabel polysilicon 1990 -2986 1990 -2986 0 3
rlabel polysilicon 1997 -2980 1997 -2980 0 1
rlabel polysilicon 1997 -2986 1997 -2986 0 3
rlabel polysilicon 2004 -2980 2004 -2980 0 1
rlabel polysilicon 2004 -2986 2004 -2986 0 3
rlabel polysilicon 2011 -2980 2011 -2980 0 1
rlabel polysilicon 2011 -2986 2011 -2986 0 3
rlabel polysilicon 2018 -2980 2018 -2980 0 1
rlabel polysilicon 2018 -2986 2018 -2986 0 3
rlabel polysilicon 2025 -2980 2025 -2980 0 1
rlabel polysilicon 2025 -2986 2025 -2986 0 3
rlabel polysilicon 2032 -2980 2032 -2980 0 1
rlabel polysilicon 2032 -2986 2032 -2986 0 3
rlabel polysilicon 2039 -2980 2039 -2980 0 1
rlabel polysilicon 2039 -2986 2039 -2986 0 3
rlabel polysilicon 2046 -2980 2046 -2980 0 1
rlabel polysilicon 2046 -2986 2046 -2986 0 3
rlabel polysilicon 2053 -2980 2053 -2980 0 1
rlabel polysilicon 2053 -2986 2053 -2986 0 3
rlabel polysilicon 2060 -2980 2060 -2980 0 1
rlabel polysilicon 2060 -2986 2060 -2986 0 3
rlabel polysilicon 2067 -2980 2067 -2980 0 1
rlabel polysilicon 2067 -2986 2067 -2986 0 3
rlabel polysilicon 2074 -2980 2074 -2980 0 1
rlabel polysilicon 2074 -2986 2074 -2986 0 3
rlabel polysilicon 2081 -2980 2081 -2980 0 1
rlabel polysilicon 2081 -2986 2081 -2986 0 3
rlabel polysilicon 2088 -2980 2088 -2980 0 1
rlabel polysilicon 2088 -2986 2088 -2986 0 3
rlabel polysilicon 2095 -2980 2095 -2980 0 1
rlabel polysilicon 2098 -2980 2098 -2980 0 2
rlabel polysilicon 2095 -2986 2095 -2986 0 3
rlabel polysilicon 2098 -2986 2098 -2986 0 4
rlabel polysilicon 2102 -2980 2102 -2980 0 1
rlabel polysilicon 2102 -2986 2102 -2986 0 3
rlabel polysilicon 2109 -2980 2109 -2980 0 1
rlabel polysilicon 2109 -2986 2109 -2986 0 3
rlabel polysilicon 2116 -2980 2116 -2980 0 1
rlabel polysilicon 2116 -2986 2116 -2986 0 3
rlabel polysilicon 2123 -2980 2123 -2980 0 1
rlabel polysilicon 2123 -2986 2123 -2986 0 3
rlabel polysilicon 2130 -2980 2130 -2980 0 1
rlabel polysilicon 2130 -2986 2130 -2986 0 3
rlabel polysilicon 2137 -2980 2137 -2980 0 1
rlabel polysilicon 2137 -2986 2137 -2986 0 3
rlabel polysilicon 2144 -2980 2144 -2980 0 1
rlabel polysilicon 2144 -2986 2144 -2986 0 3
rlabel polysilicon 2151 -2980 2151 -2980 0 1
rlabel polysilicon 2151 -2986 2151 -2986 0 3
rlabel polysilicon 23 -3095 23 -3095 0 1
rlabel polysilicon 23 -3101 23 -3101 0 3
rlabel polysilicon 30 -3095 30 -3095 0 1
rlabel polysilicon 30 -3101 30 -3101 0 3
rlabel polysilicon 37 -3095 37 -3095 0 1
rlabel polysilicon 37 -3101 37 -3101 0 3
rlabel polysilicon 58 -3095 58 -3095 0 1
rlabel polysilicon 58 -3101 58 -3101 0 3
rlabel polysilicon 65 -3095 65 -3095 0 1
rlabel polysilicon 65 -3101 65 -3101 0 3
rlabel polysilicon 72 -3095 72 -3095 0 1
rlabel polysilicon 72 -3101 72 -3101 0 3
rlabel polysilicon 79 -3101 79 -3101 0 3
rlabel polysilicon 82 -3101 82 -3101 0 4
rlabel polysilicon 86 -3095 86 -3095 0 1
rlabel polysilicon 86 -3101 86 -3101 0 3
rlabel polysilicon 93 -3095 93 -3095 0 1
rlabel polysilicon 100 -3095 100 -3095 0 1
rlabel polysilicon 100 -3101 100 -3101 0 3
rlabel polysilicon 107 -3095 107 -3095 0 1
rlabel polysilicon 107 -3101 107 -3101 0 3
rlabel polysilicon 114 -3095 114 -3095 0 1
rlabel polysilicon 114 -3101 114 -3101 0 3
rlabel polysilicon 121 -3095 121 -3095 0 1
rlabel polysilicon 121 -3101 121 -3101 0 3
rlabel polysilicon 131 -3095 131 -3095 0 2
rlabel polysilicon 128 -3101 128 -3101 0 3
rlabel polysilicon 131 -3101 131 -3101 0 4
rlabel polysilicon 138 -3095 138 -3095 0 2
rlabel polysilicon 135 -3101 135 -3101 0 3
rlabel polysilicon 138 -3101 138 -3101 0 4
rlabel polysilicon 142 -3095 142 -3095 0 1
rlabel polysilicon 142 -3101 142 -3101 0 3
rlabel polysilicon 149 -3095 149 -3095 0 1
rlabel polysilicon 149 -3101 149 -3101 0 3
rlabel polysilicon 156 -3095 156 -3095 0 1
rlabel polysilicon 156 -3101 156 -3101 0 3
rlabel polysilicon 166 -3095 166 -3095 0 2
rlabel polysilicon 163 -3101 163 -3101 0 3
rlabel polysilicon 166 -3101 166 -3101 0 4
rlabel polysilicon 173 -3095 173 -3095 0 2
rlabel polysilicon 170 -3101 170 -3101 0 3
rlabel polysilicon 173 -3101 173 -3101 0 4
rlabel polysilicon 177 -3095 177 -3095 0 1
rlabel polysilicon 177 -3101 177 -3101 0 3
rlabel polysilicon 184 -3095 184 -3095 0 1
rlabel polysilicon 184 -3101 184 -3101 0 3
rlabel polysilicon 191 -3095 191 -3095 0 1
rlabel polysilicon 191 -3101 191 -3101 0 3
rlabel polysilicon 198 -3095 198 -3095 0 1
rlabel polysilicon 198 -3101 198 -3101 0 3
rlabel polysilicon 205 -3095 205 -3095 0 1
rlabel polysilicon 208 -3095 208 -3095 0 2
rlabel polysilicon 205 -3101 205 -3101 0 3
rlabel polysilicon 208 -3101 208 -3101 0 4
rlabel polysilicon 212 -3095 212 -3095 0 1
rlabel polysilicon 212 -3101 212 -3101 0 3
rlabel polysilicon 219 -3095 219 -3095 0 1
rlabel polysilicon 219 -3101 219 -3101 0 3
rlabel polysilicon 226 -3095 226 -3095 0 1
rlabel polysilicon 226 -3101 226 -3101 0 3
rlabel polysilicon 236 -3095 236 -3095 0 2
rlabel polysilicon 236 -3101 236 -3101 0 4
rlabel polysilicon 240 -3095 240 -3095 0 1
rlabel polysilicon 240 -3101 240 -3101 0 3
rlabel polysilicon 247 -3095 247 -3095 0 1
rlabel polysilicon 247 -3101 247 -3101 0 3
rlabel polysilicon 254 -3095 254 -3095 0 1
rlabel polysilicon 254 -3101 254 -3101 0 3
rlabel polysilicon 261 -3095 261 -3095 0 1
rlabel polysilicon 261 -3101 261 -3101 0 3
rlabel polysilicon 268 -3095 268 -3095 0 1
rlabel polysilicon 268 -3101 268 -3101 0 3
rlabel polysilicon 275 -3095 275 -3095 0 1
rlabel polysilicon 275 -3101 275 -3101 0 3
rlabel polysilicon 282 -3095 282 -3095 0 1
rlabel polysilicon 282 -3101 282 -3101 0 3
rlabel polysilicon 289 -3095 289 -3095 0 1
rlabel polysilicon 289 -3101 289 -3101 0 3
rlabel polysilicon 296 -3095 296 -3095 0 1
rlabel polysilicon 296 -3101 296 -3101 0 3
rlabel polysilicon 303 -3095 303 -3095 0 1
rlabel polysilicon 303 -3101 303 -3101 0 3
rlabel polysilicon 310 -3095 310 -3095 0 1
rlabel polysilicon 310 -3101 310 -3101 0 3
rlabel polysilicon 317 -3095 317 -3095 0 1
rlabel polysilicon 317 -3101 317 -3101 0 3
rlabel polysilicon 324 -3095 324 -3095 0 1
rlabel polysilicon 324 -3101 324 -3101 0 3
rlabel polysilicon 331 -3095 331 -3095 0 1
rlabel polysilicon 331 -3101 331 -3101 0 3
rlabel polysilicon 338 -3095 338 -3095 0 1
rlabel polysilicon 338 -3101 338 -3101 0 3
rlabel polysilicon 345 -3095 345 -3095 0 1
rlabel polysilicon 345 -3101 345 -3101 0 3
rlabel polysilicon 352 -3095 352 -3095 0 1
rlabel polysilicon 352 -3101 352 -3101 0 3
rlabel polysilicon 359 -3095 359 -3095 0 1
rlabel polysilicon 359 -3101 359 -3101 0 3
rlabel polysilicon 366 -3095 366 -3095 0 1
rlabel polysilicon 366 -3101 366 -3101 0 3
rlabel polysilicon 373 -3095 373 -3095 0 1
rlabel polysilicon 373 -3101 373 -3101 0 3
rlabel polysilicon 380 -3095 380 -3095 0 1
rlabel polysilicon 380 -3101 380 -3101 0 3
rlabel polysilicon 387 -3095 387 -3095 0 1
rlabel polysilicon 387 -3101 387 -3101 0 3
rlabel polysilicon 394 -3095 394 -3095 0 1
rlabel polysilicon 394 -3101 394 -3101 0 3
rlabel polysilicon 401 -3095 401 -3095 0 1
rlabel polysilicon 401 -3101 401 -3101 0 3
rlabel polysilicon 408 -3095 408 -3095 0 1
rlabel polysilicon 408 -3101 408 -3101 0 3
rlabel polysilicon 415 -3095 415 -3095 0 1
rlabel polysilicon 415 -3101 415 -3101 0 3
rlabel polysilicon 422 -3095 422 -3095 0 1
rlabel polysilicon 422 -3101 422 -3101 0 3
rlabel polysilicon 429 -3095 429 -3095 0 1
rlabel polysilicon 429 -3101 429 -3101 0 3
rlabel polysilicon 436 -3095 436 -3095 0 1
rlabel polysilicon 436 -3101 436 -3101 0 3
rlabel polysilicon 443 -3095 443 -3095 0 1
rlabel polysilicon 443 -3101 443 -3101 0 3
rlabel polysilicon 450 -3095 450 -3095 0 1
rlabel polysilicon 450 -3101 450 -3101 0 3
rlabel polysilicon 457 -3095 457 -3095 0 1
rlabel polysilicon 460 -3095 460 -3095 0 2
rlabel polysilicon 457 -3101 457 -3101 0 3
rlabel polysilicon 460 -3101 460 -3101 0 4
rlabel polysilicon 464 -3095 464 -3095 0 1
rlabel polysilicon 464 -3101 464 -3101 0 3
rlabel polysilicon 471 -3095 471 -3095 0 1
rlabel polysilicon 471 -3101 471 -3101 0 3
rlabel polysilicon 478 -3095 478 -3095 0 1
rlabel polysilicon 478 -3101 478 -3101 0 3
rlabel polysilicon 485 -3095 485 -3095 0 1
rlabel polysilicon 485 -3101 485 -3101 0 3
rlabel polysilicon 492 -3095 492 -3095 0 1
rlabel polysilicon 492 -3101 492 -3101 0 3
rlabel polysilicon 499 -3095 499 -3095 0 1
rlabel polysilicon 499 -3101 499 -3101 0 3
rlabel polysilicon 506 -3095 506 -3095 0 1
rlabel polysilicon 506 -3101 506 -3101 0 3
rlabel polysilicon 513 -3095 513 -3095 0 1
rlabel polysilicon 513 -3101 513 -3101 0 3
rlabel polysilicon 520 -3095 520 -3095 0 1
rlabel polysilicon 520 -3101 520 -3101 0 3
rlabel polysilicon 527 -3101 527 -3101 0 3
rlabel polysilicon 530 -3101 530 -3101 0 4
rlabel polysilicon 534 -3095 534 -3095 0 1
rlabel polysilicon 534 -3101 534 -3101 0 3
rlabel polysilicon 541 -3095 541 -3095 0 1
rlabel polysilicon 541 -3101 541 -3101 0 3
rlabel polysilicon 548 -3095 548 -3095 0 1
rlabel polysilicon 548 -3101 548 -3101 0 3
rlabel polysilicon 555 -3095 555 -3095 0 1
rlabel polysilicon 555 -3101 555 -3101 0 3
rlabel polysilicon 562 -3095 562 -3095 0 1
rlabel polysilicon 562 -3101 562 -3101 0 3
rlabel polysilicon 569 -3095 569 -3095 0 1
rlabel polysilicon 569 -3101 569 -3101 0 3
rlabel polysilicon 576 -3095 576 -3095 0 1
rlabel polysilicon 576 -3101 576 -3101 0 3
rlabel polysilicon 583 -3095 583 -3095 0 1
rlabel polysilicon 583 -3101 583 -3101 0 3
rlabel polysilicon 590 -3095 590 -3095 0 1
rlabel polysilicon 590 -3101 590 -3101 0 3
rlabel polysilicon 597 -3095 597 -3095 0 1
rlabel polysilicon 597 -3101 597 -3101 0 3
rlabel polysilicon 604 -3095 604 -3095 0 1
rlabel polysilicon 604 -3101 604 -3101 0 3
rlabel polysilicon 611 -3095 611 -3095 0 1
rlabel polysilicon 614 -3095 614 -3095 0 2
rlabel polysilicon 611 -3101 611 -3101 0 3
rlabel polysilicon 614 -3101 614 -3101 0 4
rlabel polysilicon 618 -3095 618 -3095 0 1
rlabel polysilicon 618 -3101 618 -3101 0 3
rlabel polysilicon 625 -3095 625 -3095 0 1
rlabel polysilicon 625 -3101 625 -3101 0 3
rlabel polysilicon 632 -3095 632 -3095 0 1
rlabel polysilicon 632 -3101 632 -3101 0 3
rlabel polysilicon 639 -3095 639 -3095 0 1
rlabel polysilicon 639 -3101 639 -3101 0 3
rlabel polysilicon 646 -3095 646 -3095 0 1
rlabel polysilicon 646 -3101 646 -3101 0 3
rlabel polysilicon 653 -3095 653 -3095 0 1
rlabel polysilicon 653 -3101 653 -3101 0 3
rlabel polysilicon 660 -3095 660 -3095 0 1
rlabel polysilicon 660 -3101 660 -3101 0 3
rlabel polysilicon 667 -3095 667 -3095 0 1
rlabel polysilicon 667 -3101 667 -3101 0 3
rlabel polysilicon 674 -3095 674 -3095 0 1
rlabel polysilicon 674 -3101 674 -3101 0 3
rlabel polysilicon 681 -3095 681 -3095 0 1
rlabel polysilicon 681 -3101 681 -3101 0 3
rlabel polysilicon 688 -3095 688 -3095 0 1
rlabel polysilicon 688 -3101 688 -3101 0 3
rlabel polysilicon 695 -3095 695 -3095 0 1
rlabel polysilicon 695 -3101 695 -3101 0 3
rlabel polysilicon 702 -3095 702 -3095 0 1
rlabel polysilicon 702 -3101 702 -3101 0 3
rlabel polysilicon 709 -3095 709 -3095 0 1
rlabel polysilicon 709 -3101 709 -3101 0 3
rlabel polysilicon 716 -3095 716 -3095 0 1
rlabel polysilicon 716 -3101 716 -3101 0 3
rlabel polysilicon 723 -3095 723 -3095 0 1
rlabel polysilicon 723 -3101 723 -3101 0 3
rlabel polysilicon 730 -3095 730 -3095 0 1
rlabel polysilicon 730 -3101 730 -3101 0 3
rlabel polysilicon 737 -3095 737 -3095 0 1
rlabel polysilicon 737 -3101 737 -3101 0 3
rlabel polysilicon 744 -3095 744 -3095 0 1
rlabel polysilicon 744 -3101 744 -3101 0 3
rlabel polysilicon 751 -3095 751 -3095 0 1
rlabel polysilicon 751 -3101 751 -3101 0 3
rlabel polysilicon 758 -3095 758 -3095 0 1
rlabel polysilicon 758 -3101 758 -3101 0 3
rlabel polysilicon 765 -3095 765 -3095 0 1
rlabel polysilicon 765 -3101 765 -3101 0 3
rlabel polysilicon 772 -3095 772 -3095 0 1
rlabel polysilicon 772 -3101 772 -3101 0 3
rlabel polysilicon 779 -3095 779 -3095 0 1
rlabel polysilicon 779 -3101 779 -3101 0 3
rlabel polysilicon 786 -3095 786 -3095 0 1
rlabel polysilicon 786 -3101 786 -3101 0 3
rlabel polysilicon 793 -3095 793 -3095 0 1
rlabel polysilicon 793 -3101 793 -3101 0 3
rlabel polysilicon 800 -3101 800 -3101 0 3
rlabel polysilicon 807 -3095 807 -3095 0 1
rlabel polysilicon 807 -3101 807 -3101 0 3
rlabel polysilicon 817 -3095 817 -3095 0 2
rlabel polysilicon 814 -3101 814 -3101 0 3
rlabel polysilicon 817 -3101 817 -3101 0 4
rlabel polysilicon 821 -3095 821 -3095 0 1
rlabel polysilicon 821 -3101 821 -3101 0 3
rlabel polysilicon 828 -3095 828 -3095 0 1
rlabel polysilicon 828 -3101 828 -3101 0 3
rlabel polysilicon 835 -3095 835 -3095 0 1
rlabel polysilicon 835 -3101 835 -3101 0 3
rlabel polysilicon 842 -3095 842 -3095 0 1
rlabel polysilicon 842 -3101 842 -3101 0 3
rlabel polysilicon 849 -3095 849 -3095 0 1
rlabel polysilicon 849 -3101 849 -3101 0 3
rlabel polysilicon 856 -3095 856 -3095 0 1
rlabel polysilicon 856 -3101 856 -3101 0 3
rlabel polysilicon 863 -3095 863 -3095 0 1
rlabel polysilicon 866 -3101 866 -3101 0 4
rlabel polysilicon 870 -3095 870 -3095 0 1
rlabel polysilicon 870 -3101 870 -3101 0 3
rlabel polysilicon 877 -3095 877 -3095 0 1
rlabel polysilicon 880 -3095 880 -3095 0 2
rlabel polysilicon 877 -3101 877 -3101 0 3
rlabel polysilicon 880 -3101 880 -3101 0 4
rlabel polysilicon 884 -3095 884 -3095 0 1
rlabel polysilicon 884 -3101 884 -3101 0 3
rlabel polysilicon 894 -3095 894 -3095 0 2
rlabel polysilicon 891 -3101 891 -3101 0 3
rlabel polysilicon 898 -3095 898 -3095 0 1
rlabel polysilicon 898 -3101 898 -3101 0 3
rlabel polysilicon 905 -3095 905 -3095 0 1
rlabel polysilicon 905 -3101 905 -3101 0 3
rlabel polysilicon 912 -3095 912 -3095 0 1
rlabel polysilicon 915 -3095 915 -3095 0 2
rlabel polysilicon 912 -3101 912 -3101 0 3
rlabel polysilicon 919 -3095 919 -3095 0 1
rlabel polysilicon 919 -3101 919 -3101 0 3
rlabel polysilicon 926 -3095 926 -3095 0 1
rlabel polysilicon 926 -3101 926 -3101 0 3
rlabel polysilicon 933 -3095 933 -3095 0 1
rlabel polysilicon 933 -3101 933 -3101 0 3
rlabel polysilicon 940 -3095 940 -3095 0 1
rlabel polysilicon 940 -3101 940 -3101 0 3
rlabel polysilicon 947 -3095 947 -3095 0 1
rlabel polysilicon 947 -3101 947 -3101 0 3
rlabel polysilicon 954 -3095 954 -3095 0 1
rlabel polysilicon 954 -3101 954 -3101 0 3
rlabel polysilicon 961 -3095 961 -3095 0 1
rlabel polysilicon 961 -3101 961 -3101 0 3
rlabel polysilicon 968 -3095 968 -3095 0 1
rlabel polysilicon 968 -3101 968 -3101 0 3
rlabel polysilicon 975 -3095 975 -3095 0 1
rlabel polysilicon 975 -3101 975 -3101 0 3
rlabel polysilicon 982 -3095 982 -3095 0 1
rlabel polysilicon 982 -3101 982 -3101 0 3
rlabel polysilicon 989 -3095 989 -3095 0 1
rlabel polysilicon 989 -3101 989 -3101 0 3
rlabel polysilicon 996 -3095 996 -3095 0 1
rlabel polysilicon 996 -3101 996 -3101 0 3
rlabel polysilicon 1003 -3095 1003 -3095 0 1
rlabel polysilicon 1003 -3101 1003 -3101 0 3
rlabel polysilicon 1010 -3095 1010 -3095 0 1
rlabel polysilicon 1010 -3101 1010 -3101 0 3
rlabel polysilicon 1017 -3095 1017 -3095 0 1
rlabel polysilicon 1017 -3101 1017 -3101 0 3
rlabel polysilicon 1024 -3095 1024 -3095 0 1
rlabel polysilicon 1024 -3101 1024 -3101 0 3
rlabel polysilicon 1031 -3095 1031 -3095 0 1
rlabel polysilicon 1031 -3101 1031 -3101 0 3
rlabel polysilicon 1038 -3095 1038 -3095 0 1
rlabel polysilicon 1038 -3101 1038 -3101 0 3
rlabel polysilicon 1045 -3095 1045 -3095 0 1
rlabel polysilicon 1045 -3101 1045 -3101 0 3
rlabel polysilicon 1055 -3095 1055 -3095 0 2
rlabel polysilicon 1055 -3101 1055 -3101 0 4
rlabel polysilicon 1059 -3095 1059 -3095 0 1
rlabel polysilicon 1059 -3101 1059 -3101 0 3
rlabel polysilicon 1066 -3095 1066 -3095 0 1
rlabel polysilicon 1066 -3101 1066 -3101 0 3
rlabel polysilicon 1073 -3095 1073 -3095 0 1
rlabel polysilicon 1076 -3095 1076 -3095 0 2
rlabel polysilicon 1073 -3101 1073 -3101 0 3
rlabel polysilicon 1076 -3101 1076 -3101 0 4
rlabel polysilicon 1083 -3095 1083 -3095 0 2
rlabel polysilicon 1080 -3101 1080 -3101 0 3
rlabel polysilicon 1083 -3101 1083 -3101 0 4
rlabel polysilicon 1087 -3095 1087 -3095 0 1
rlabel polysilicon 1087 -3101 1087 -3101 0 3
rlabel polysilicon 1094 -3095 1094 -3095 0 1
rlabel polysilicon 1094 -3101 1094 -3101 0 3
rlabel polysilicon 1101 -3095 1101 -3095 0 1
rlabel polysilicon 1101 -3101 1101 -3101 0 3
rlabel polysilicon 1108 -3095 1108 -3095 0 1
rlabel polysilicon 1108 -3101 1108 -3101 0 3
rlabel polysilicon 1115 -3095 1115 -3095 0 1
rlabel polysilicon 1115 -3101 1115 -3101 0 3
rlabel polysilicon 1122 -3095 1122 -3095 0 1
rlabel polysilicon 1122 -3101 1122 -3101 0 3
rlabel polysilicon 1125 -3101 1125 -3101 0 4
rlabel polysilicon 1129 -3095 1129 -3095 0 1
rlabel polysilicon 1129 -3101 1129 -3101 0 3
rlabel polysilicon 1136 -3095 1136 -3095 0 1
rlabel polysilicon 1136 -3101 1136 -3101 0 3
rlabel polysilicon 1143 -3095 1143 -3095 0 1
rlabel polysilicon 1143 -3101 1143 -3101 0 3
rlabel polysilicon 1150 -3095 1150 -3095 0 1
rlabel polysilicon 1150 -3101 1150 -3101 0 3
rlabel polysilicon 1157 -3095 1157 -3095 0 1
rlabel polysilicon 1160 -3095 1160 -3095 0 2
rlabel polysilicon 1157 -3101 1157 -3101 0 3
rlabel polysilicon 1160 -3101 1160 -3101 0 4
rlabel polysilicon 1164 -3095 1164 -3095 0 1
rlabel polysilicon 1164 -3101 1164 -3101 0 3
rlabel polysilicon 1171 -3095 1171 -3095 0 1
rlabel polysilicon 1171 -3101 1171 -3101 0 3
rlabel polysilicon 1178 -3095 1178 -3095 0 1
rlabel polysilicon 1178 -3101 1178 -3101 0 3
rlabel polysilicon 1185 -3095 1185 -3095 0 1
rlabel polysilicon 1185 -3101 1185 -3101 0 3
rlabel polysilicon 1192 -3095 1192 -3095 0 1
rlabel polysilicon 1192 -3101 1192 -3101 0 3
rlabel polysilicon 1199 -3095 1199 -3095 0 1
rlabel polysilicon 1199 -3101 1199 -3101 0 3
rlabel polysilicon 1206 -3095 1206 -3095 0 1
rlabel polysilicon 1206 -3101 1206 -3101 0 3
rlabel polysilicon 1213 -3095 1213 -3095 0 1
rlabel polysilicon 1216 -3095 1216 -3095 0 2
rlabel polysilicon 1213 -3101 1213 -3101 0 3
rlabel polysilicon 1216 -3101 1216 -3101 0 4
rlabel polysilicon 1220 -3095 1220 -3095 0 1
rlabel polysilicon 1220 -3101 1220 -3101 0 3
rlabel polysilicon 1227 -3095 1227 -3095 0 1
rlabel polysilicon 1227 -3101 1227 -3101 0 3
rlabel polysilicon 1234 -3095 1234 -3095 0 1
rlabel polysilicon 1237 -3095 1237 -3095 0 2
rlabel polysilicon 1234 -3101 1234 -3101 0 3
rlabel polysilicon 1237 -3101 1237 -3101 0 4
rlabel polysilicon 1241 -3095 1241 -3095 0 1
rlabel polysilicon 1241 -3101 1241 -3101 0 3
rlabel polysilicon 1248 -3101 1248 -3101 0 3
rlabel polysilicon 1255 -3095 1255 -3095 0 1
rlabel polysilicon 1255 -3101 1255 -3101 0 3
rlabel polysilicon 1262 -3095 1262 -3095 0 1
rlabel polysilicon 1262 -3101 1262 -3101 0 3
rlabel polysilicon 1269 -3095 1269 -3095 0 1
rlabel polysilicon 1269 -3101 1269 -3101 0 3
rlabel polysilicon 1276 -3101 1276 -3101 0 3
rlabel polysilicon 1283 -3095 1283 -3095 0 1
rlabel polysilicon 1283 -3101 1283 -3101 0 3
rlabel polysilicon 1290 -3095 1290 -3095 0 1
rlabel polysilicon 1290 -3101 1290 -3101 0 3
rlabel polysilicon 1297 -3095 1297 -3095 0 1
rlabel polysilicon 1297 -3101 1297 -3101 0 3
rlabel polysilicon 1304 -3095 1304 -3095 0 1
rlabel polysilicon 1304 -3101 1304 -3101 0 3
rlabel polysilicon 1311 -3095 1311 -3095 0 1
rlabel polysilicon 1311 -3101 1311 -3101 0 3
rlabel polysilicon 1314 -3101 1314 -3101 0 4
rlabel polysilicon 1318 -3095 1318 -3095 0 1
rlabel polysilicon 1318 -3101 1318 -3101 0 3
rlabel polysilicon 1325 -3095 1325 -3095 0 1
rlabel polysilicon 1325 -3101 1325 -3101 0 3
rlabel polysilicon 1332 -3095 1332 -3095 0 1
rlabel polysilicon 1332 -3101 1332 -3101 0 3
rlabel polysilicon 1339 -3095 1339 -3095 0 1
rlabel polysilicon 1339 -3101 1339 -3101 0 3
rlabel polysilicon 1346 -3095 1346 -3095 0 1
rlabel polysilicon 1346 -3101 1346 -3101 0 3
rlabel polysilicon 1353 -3095 1353 -3095 0 1
rlabel polysilicon 1353 -3101 1353 -3101 0 3
rlabel polysilicon 1360 -3095 1360 -3095 0 1
rlabel polysilicon 1360 -3101 1360 -3101 0 3
rlabel polysilicon 1367 -3095 1367 -3095 0 1
rlabel polysilicon 1367 -3101 1367 -3101 0 3
rlabel polysilicon 1374 -3095 1374 -3095 0 1
rlabel polysilicon 1374 -3101 1374 -3101 0 3
rlabel polysilicon 1381 -3095 1381 -3095 0 1
rlabel polysilicon 1381 -3101 1381 -3101 0 3
rlabel polysilicon 1388 -3095 1388 -3095 0 1
rlabel polysilicon 1388 -3101 1388 -3101 0 3
rlabel polysilicon 1398 -3095 1398 -3095 0 2
rlabel polysilicon 1395 -3101 1395 -3101 0 3
rlabel polysilicon 1398 -3101 1398 -3101 0 4
rlabel polysilicon 1402 -3095 1402 -3095 0 1
rlabel polysilicon 1405 -3095 1405 -3095 0 2
rlabel polysilicon 1402 -3101 1402 -3101 0 3
rlabel polysilicon 1409 -3095 1409 -3095 0 1
rlabel polysilicon 1409 -3101 1409 -3101 0 3
rlabel polysilicon 1416 -3095 1416 -3095 0 1
rlabel polysilicon 1416 -3101 1416 -3101 0 3
rlabel polysilicon 1423 -3095 1423 -3095 0 1
rlabel polysilicon 1423 -3101 1423 -3101 0 3
rlabel polysilicon 1430 -3095 1430 -3095 0 1
rlabel polysilicon 1430 -3101 1430 -3101 0 3
rlabel polysilicon 1437 -3095 1437 -3095 0 1
rlabel polysilicon 1437 -3101 1437 -3101 0 3
rlabel polysilicon 1444 -3101 1444 -3101 0 3
rlabel polysilicon 1447 -3101 1447 -3101 0 4
rlabel polysilicon 1451 -3095 1451 -3095 0 1
rlabel polysilicon 1451 -3101 1451 -3101 0 3
rlabel polysilicon 1458 -3095 1458 -3095 0 1
rlabel polysilicon 1458 -3101 1458 -3101 0 3
rlabel polysilicon 1465 -3095 1465 -3095 0 1
rlabel polysilicon 1465 -3101 1465 -3101 0 3
rlabel polysilicon 1472 -3095 1472 -3095 0 1
rlabel polysilicon 1472 -3101 1472 -3101 0 3
rlabel polysilicon 1479 -3095 1479 -3095 0 1
rlabel polysilicon 1479 -3101 1479 -3101 0 3
rlabel polysilicon 1486 -3095 1486 -3095 0 1
rlabel polysilicon 1486 -3101 1486 -3101 0 3
rlabel polysilicon 1493 -3095 1493 -3095 0 1
rlabel polysilicon 1493 -3101 1493 -3101 0 3
rlabel polysilicon 1500 -3095 1500 -3095 0 1
rlabel polysilicon 1500 -3101 1500 -3101 0 3
rlabel polysilicon 1507 -3095 1507 -3095 0 1
rlabel polysilicon 1507 -3101 1507 -3101 0 3
rlabel polysilicon 1514 -3095 1514 -3095 0 1
rlabel polysilicon 1514 -3101 1514 -3101 0 3
rlabel polysilicon 1521 -3095 1521 -3095 0 1
rlabel polysilicon 1521 -3101 1521 -3101 0 3
rlabel polysilicon 1528 -3095 1528 -3095 0 1
rlabel polysilicon 1528 -3101 1528 -3101 0 3
rlabel polysilicon 1535 -3095 1535 -3095 0 1
rlabel polysilicon 1535 -3101 1535 -3101 0 3
rlabel polysilicon 1542 -3095 1542 -3095 0 1
rlabel polysilicon 1542 -3101 1542 -3101 0 3
rlabel polysilicon 1549 -3095 1549 -3095 0 1
rlabel polysilicon 1549 -3101 1549 -3101 0 3
rlabel polysilicon 1556 -3095 1556 -3095 0 1
rlabel polysilicon 1559 -3095 1559 -3095 0 2
rlabel polysilicon 1556 -3101 1556 -3101 0 3
rlabel polysilicon 1559 -3101 1559 -3101 0 4
rlabel polysilicon 1566 -3095 1566 -3095 0 2
rlabel polysilicon 1563 -3101 1563 -3101 0 3
rlabel polysilicon 1566 -3101 1566 -3101 0 4
rlabel polysilicon 1570 -3095 1570 -3095 0 1
rlabel polysilicon 1570 -3101 1570 -3101 0 3
rlabel polysilicon 1577 -3095 1577 -3095 0 1
rlabel polysilicon 1577 -3101 1577 -3101 0 3
rlabel polysilicon 1584 -3095 1584 -3095 0 1
rlabel polysilicon 1584 -3101 1584 -3101 0 3
rlabel polysilicon 1591 -3095 1591 -3095 0 1
rlabel polysilicon 1591 -3101 1591 -3101 0 3
rlabel polysilicon 1598 -3095 1598 -3095 0 1
rlabel polysilicon 1598 -3101 1598 -3101 0 3
rlabel polysilicon 1605 -3095 1605 -3095 0 1
rlabel polysilicon 1605 -3101 1605 -3101 0 3
rlabel polysilicon 1612 -3095 1612 -3095 0 1
rlabel polysilicon 1612 -3101 1612 -3101 0 3
rlabel polysilicon 1619 -3095 1619 -3095 0 1
rlabel polysilicon 1619 -3101 1619 -3101 0 3
rlabel polysilicon 1626 -3095 1626 -3095 0 1
rlabel polysilicon 1626 -3101 1626 -3101 0 3
rlabel polysilicon 1633 -3095 1633 -3095 0 1
rlabel polysilicon 1633 -3101 1633 -3101 0 3
rlabel polysilicon 1640 -3095 1640 -3095 0 1
rlabel polysilicon 1640 -3101 1640 -3101 0 3
rlabel polysilicon 1647 -3095 1647 -3095 0 1
rlabel polysilicon 1647 -3101 1647 -3101 0 3
rlabel polysilicon 1654 -3095 1654 -3095 0 1
rlabel polysilicon 1654 -3101 1654 -3101 0 3
rlabel polysilicon 1661 -3095 1661 -3095 0 1
rlabel polysilicon 1661 -3101 1661 -3101 0 3
rlabel polysilicon 1668 -3095 1668 -3095 0 1
rlabel polysilicon 1668 -3101 1668 -3101 0 3
rlabel polysilicon 1675 -3095 1675 -3095 0 1
rlabel polysilicon 1675 -3101 1675 -3101 0 3
rlabel polysilicon 1682 -3095 1682 -3095 0 1
rlabel polysilicon 1685 -3095 1685 -3095 0 2
rlabel polysilicon 1685 -3101 1685 -3101 0 4
rlabel polysilicon 1689 -3095 1689 -3095 0 1
rlabel polysilicon 1689 -3101 1689 -3101 0 3
rlabel polysilicon 1696 -3095 1696 -3095 0 1
rlabel polysilicon 1696 -3101 1696 -3101 0 3
rlabel polysilicon 1703 -3095 1703 -3095 0 1
rlabel polysilicon 1703 -3101 1703 -3101 0 3
rlabel polysilicon 1710 -3095 1710 -3095 0 1
rlabel polysilicon 1710 -3101 1710 -3101 0 3
rlabel polysilicon 1717 -3095 1717 -3095 0 1
rlabel polysilicon 1717 -3101 1717 -3101 0 3
rlabel polysilicon 1724 -3095 1724 -3095 0 1
rlabel polysilicon 1724 -3101 1724 -3101 0 3
rlabel polysilicon 1731 -3095 1731 -3095 0 1
rlabel polysilicon 1731 -3101 1731 -3101 0 3
rlabel polysilicon 1738 -3095 1738 -3095 0 1
rlabel polysilicon 1738 -3101 1738 -3101 0 3
rlabel polysilicon 1745 -3095 1745 -3095 0 1
rlabel polysilicon 1745 -3101 1745 -3101 0 3
rlabel polysilicon 1752 -3095 1752 -3095 0 1
rlabel polysilicon 1752 -3101 1752 -3101 0 3
rlabel polysilicon 1759 -3095 1759 -3095 0 1
rlabel polysilicon 1759 -3101 1759 -3101 0 3
rlabel polysilicon 1766 -3095 1766 -3095 0 1
rlabel polysilicon 1766 -3101 1766 -3101 0 3
rlabel polysilicon 1773 -3095 1773 -3095 0 1
rlabel polysilicon 1773 -3101 1773 -3101 0 3
rlabel polysilicon 1780 -3095 1780 -3095 0 1
rlabel polysilicon 1780 -3101 1780 -3101 0 3
rlabel polysilicon 1787 -3095 1787 -3095 0 1
rlabel polysilicon 1787 -3101 1787 -3101 0 3
rlabel polysilicon 1794 -3095 1794 -3095 0 1
rlabel polysilicon 1794 -3101 1794 -3101 0 3
rlabel polysilicon 1801 -3095 1801 -3095 0 1
rlabel polysilicon 1801 -3101 1801 -3101 0 3
rlabel polysilicon 1808 -3095 1808 -3095 0 1
rlabel polysilicon 1808 -3101 1808 -3101 0 3
rlabel polysilicon 1815 -3095 1815 -3095 0 1
rlabel polysilicon 1815 -3101 1815 -3101 0 3
rlabel polysilicon 1822 -3095 1822 -3095 0 1
rlabel polysilicon 1822 -3101 1822 -3101 0 3
rlabel polysilicon 1829 -3095 1829 -3095 0 1
rlabel polysilicon 1829 -3101 1829 -3101 0 3
rlabel polysilicon 1836 -3095 1836 -3095 0 1
rlabel polysilicon 1836 -3101 1836 -3101 0 3
rlabel polysilicon 1843 -3095 1843 -3095 0 1
rlabel polysilicon 1843 -3101 1843 -3101 0 3
rlabel polysilicon 1850 -3095 1850 -3095 0 1
rlabel polysilicon 1850 -3101 1850 -3101 0 3
rlabel polysilicon 1857 -3095 1857 -3095 0 1
rlabel polysilicon 1857 -3101 1857 -3101 0 3
rlabel polysilicon 1864 -3095 1864 -3095 0 1
rlabel polysilicon 1864 -3101 1864 -3101 0 3
rlabel polysilicon 1871 -3095 1871 -3095 0 1
rlabel polysilicon 1874 -3095 1874 -3095 0 2
rlabel polysilicon 1871 -3101 1871 -3101 0 3
rlabel polysilicon 1881 -3095 1881 -3095 0 2
rlabel polysilicon 1878 -3101 1878 -3101 0 3
rlabel polysilicon 1881 -3101 1881 -3101 0 4
rlabel polysilicon 1885 -3095 1885 -3095 0 1
rlabel polysilicon 1885 -3101 1885 -3101 0 3
rlabel polysilicon 1892 -3095 1892 -3095 0 1
rlabel polysilicon 1892 -3101 1892 -3101 0 3
rlabel polysilicon 1899 -3095 1899 -3095 0 1
rlabel polysilicon 1899 -3101 1899 -3101 0 3
rlabel polysilicon 1906 -3095 1906 -3095 0 1
rlabel polysilicon 1906 -3101 1906 -3101 0 3
rlabel polysilicon 1913 -3095 1913 -3095 0 1
rlabel polysilicon 1913 -3101 1913 -3101 0 3
rlabel polysilicon 1920 -3095 1920 -3095 0 1
rlabel polysilicon 1920 -3101 1920 -3101 0 3
rlabel polysilicon 1927 -3095 1927 -3095 0 1
rlabel polysilicon 1927 -3101 1927 -3101 0 3
rlabel polysilicon 1934 -3095 1934 -3095 0 1
rlabel polysilicon 1934 -3101 1934 -3101 0 3
rlabel polysilicon 1941 -3095 1941 -3095 0 1
rlabel polysilicon 1941 -3101 1941 -3101 0 3
rlabel polysilicon 1948 -3095 1948 -3095 0 1
rlabel polysilicon 1948 -3101 1948 -3101 0 3
rlabel polysilicon 1955 -3095 1955 -3095 0 1
rlabel polysilicon 1955 -3101 1955 -3101 0 3
rlabel polysilicon 1962 -3095 1962 -3095 0 1
rlabel polysilicon 1965 -3095 1965 -3095 0 2
rlabel polysilicon 1962 -3101 1962 -3101 0 3
rlabel polysilicon 1965 -3101 1965 -3101 0 4
rlabel polysilicon 1969 -3095 1969 -3095 0 1
rlabel polysilicon 1969 -3101 1969 -3101 0 3
rlabel polysilicon 1976 -3095 1976 -3095 0 1
rlabel polysilicon 1976 -3101 1976 -3101 0 3
rlabel polysilicon 1983 -3095 1983 -3095 0 1
rlabel polysilicon 1983 -3101 1983 -3101 0 3
rlabel polysilicon 1990 -3095 1990 -3095 0 1
rlabel polysilicon 1990 -3101 1990 -3101 0 3
rlabel polysilicon 1997 -3095 1997 -3095 0 1
rlabel polysilicon 1997 -3101 1997 -3101 0 3
rlabel polysilicon 2004 -3095 2004 -3095 0 1
rlabel polysilicon 2004 -3101 2004 -3101 0 3
rlabel polysilicon 2032 -3095 2032 -3095 0 1
rlabel polysilicon 2032 -3101 2032 -3101 0 3
rlabel polysilicon 2046 -3095 2046 -3095 0 1
rlabel polysilicon 2046 -3101 2046 -3101 0 3
rlabel polysilicon 2074 -3095 2074 -3095 0 1
rlabel polysilicon 2074 -3101 2074 -3101 0 3
rlabel polysilicon 93 -3226 93 -3226 0 1
rlabel polysilicon 93 -3232 93 -3232 0 3
rlabel polysilicon 100 -3226 100 -3226 0 1
rlabel polysilicon 100 -3232 100 -3232 0 3
rlabel polysilicon 107 -3226 107 -3226 0 1
rlabel polysilicon 107 -3232 107 -3232 0 3
rlabel polysilicon 114 -3226 114 -3226 0 1
rlabel polysilicon 117 -3232 117 -3232 0 4
rlabel polysilicon 121 -3226 121 -3226 0 1
rlabel polysilicon 121 -3232 121 -3232 0 3
rlabel polysilicon 128 -3226 128 -3226 0 1
rlabel polysilicon 128 -3232 128 -3232 0 3
rlabel polysilicon 135 -3226 135 -3226 0 1
rlabel polysilicon 135 -3232 135 -3232 0 3
rlabel polysilicon 142 -3226 142 -3226 0 1
rlabel polysilicon 142 -3232 142 -3232 0 3
rlabel polysilicon 149 -3226 149 -3226 0 1
rlabel polysilicon 149 -3232 149 -3232 0 3
rlabel polysilicon 156 -3226 156 -3226 0 1
rlabel polysilicon 156 -3232 156 -3232 0 3
rlabel polysilicon 163 -3226 163 -3226 0 1
rlabel polysilicon 163 -3232 163 -3232 0 3
rlabel polysilicon 170 -3226 170 -3226 0 1
rlabel polysilicon 173 -3232 173 -3232 0 4
rlabel polysilicon 177 -3226 177 -3226 0 1
rlabel polysilicon 177 -3232 177 -3232 0 3
rlabel polysilicon 187 -3226 187 -3226 0 2
rlabel polysilicon 187 -3232 187 -3232 0 4
rlabel polysilicon 191 -3226 191 -3226 0 1
rlabel polysilicon 194 -3226 194 -3226 0 2
rlabel polysilicon 191 -3232 191 -3232 0 3
rlabel polysilicon 198 -3226 198 -3226 0 1
rlabel polysilicon 198 -3232 198 -3232 0 3
rlabel polysilicon 205 -3226 205 -3226 0 1
rlabel polysilicon 208 -3226 208 -3226 0 2
rlabel polysilicon 205 -3232 205 -3232 0 3
rlabel polysilicon 208 -3232 208 -3232 0 4
rlabel polysilicon 212 -3226 212 -3226 0 1
rlabel polysilicon 212 -3232 212 -3232 0 3
rlabel polysilicon 219 -3226 219 -3226 0 1
rlabel polysilicon 219 -3232 219 -3232 0 3
rlabel polysilicon 226 -3226 226 -3226 0 1
rlabel polysilicon 226 -3232 226 -3232 0 3
rlabel polysilicon 233 -3226 233 -3226 0 1
rlabel polysilicon 233 -3232 233 -3232 0 3
rlabel polysilicon 240 -3226 240 -3226 0 1
rlabel polysilicon 240 -3232 240 -3232 0 3
rlabel polysilicon 247 -3226 247 -3226 0 1
rlabel polysilicon 247 -3232 247 -3232 0 3
rlabel polysilicon 254 -3226 254 -3226 0 1
rlabel polysilicon 254 -3232 254 -3232 0 3
rlabel polysilicon 261 -3226 261 -3226 0 1
rlabel polysilicon 261 -3232 261 -3232 0 3
rlabel polysilicon 268 -3226 268 -3226 0 1
rlabel polysilicon 268 -3232 268 -3232 0 3
rlabel polysilicon 275 -3226 275 -3226 0 1
rlabel polysilicon 275 -3232 275 -3232 0 3
rlabel polysilicon 282 -3226 282 -3226 0 1
rlabel polysilicon 282 -3232 282 -3232 0 3
rlabel polysilicon 289 -3226 289 -3226 0 1
rlabel polysilicon 289 -3232 289 -3232 0 3
rlabel polysilicon 296 -3226 296 -3226 0 1
rlabel polysilicon 296 -3232 296 -3232 0 3
rlabel polysilicon 303 -3226 303 -3226 0 1
rlabel polysilicon 303 -3232 303 -3232 0 3
rlabel polysilicon 310 -3226 310 -3226 0 1
rlabel polysilicon 310 -3232 310 -3232 0 3
rlabel polysilicon 317 -3226 317 -3226 0 1
rlabel polysilicon 317 -3232 317 -3232 0 3
rlabel polysilicon 324 -3226 324 -3226 0 1
rlabel polysilicon 324 -3232 324 -3232 0 3
rlabel polysilicon 331 -3226 331 -3226 0 1
rlabel polysilicon 331 -3232 331 -3232 0 3
rlabel polysilicon 338 -3226 338 -3226 0 1
rlabel polysilicon 338 -3232 338 -3232 0 3
rlabel polysilicon 345 -3226 345 -3226 0 1
rlabel polysilicon 345 -3232 345 -3232 0 3
rlabel polysilicon 352 -3226 352 -3226 0 1
rlabel polysilicon 352 -3232 352 -3232 0 3
rlabel polysilicon 359 -3226 359 -3226 0 1
rlabel polysilicon 359 -3232 359 -3232 0 3
rlabel polysilicon 366 -3226 366 -3226 0 1
rlabel polysilicon 366 -3232 366 -3232 0 3
rlabel polysilicon 373 -3226 373 -3226 0 1
rlabel polysilicon 373 -3232 373 -3232 0 3
rlabel polysilicon 380 -3226 380 -3226 0 1
rlabel polysilicon 380 -3232 380 -3232 0 3
rlabel polysilicon 387 -3226 387 -3226 0 1
rlabel polysilicon 387 -3232 387 -3232 0 3
rlabel polysilicon 394 -3226 394 -3226 0 1
rlabel polysilicon 394 -3232 394 -3232 0 3
rlabel polysilicon 401 -3226 401 -3226 0 1
rlabel polysilicon 404 -3226 404 -3226 0 2
rlabel polysilicon 401 -3232 401 -3232 0 3
rlabel polysilicon 404 -3232 404 -3232 0 4
rlabel polysilicon 408 -3226 408 -3226 0 1
rlabel polysilicon 408 -3232 408 -3232 0 3
rlabel polysilicon 415 -3226 415 -3226 0 1
rlabel polysilicon 418 -3226 418 -3226 0 2
rlabel polysilicon 415 -3232 415 -3232 0 3
rlabel polysilicon 418 -3232 418 -3232 0 4
rlabel polysilicon 425 -3226 425 -3226 0 2
rlabel polysilicon 422 -3232 422 -3232 0 3
rlabel polysilicon 429 -3226 429 -3226 0 1
rlabel polysilicon 429 -3232 429 -3232 0 3
rlabel polysilicon 436 -3226 436 -3226 0 1
rlabel polysilicon 436 -3232 436 -3232 0 3
rlabel polysilicon 443 -3226 443 -3226 0 1
rlabel polysilicon 443 -3232 443 -3232 0 3
rlabel polysilicon 450 -3226 450 -3226 0 1
rlabel polysilicon 450 -3232 450 -3232 0 3
rlabel polysilicon 457 -3226 457 -3226 0 1
rlabel polysilicon 457 -3232 457 -3232 0 3
rlabel polysilicon 464 -3226 464 -3226 0 1
rlabel polysilicon 464 -3232 464 -3232 0 3
rlabel polysilicon 471 -3226 471 -3226 0 1
rlabel polysilicon 471 -3232 471 -3232 0 3
rlabel polysilicon 478 -3226 478 -3226 0 1
rlabel polysilicon 478 -3232 478 -3232 0 3
rlabel polysilicon 485 -3226 485 -3226 0 1
rlabel polysilicon 485 -3232 485 -3232 0 3
rlabel polysilicon 492 -3226 492 -3226 0 1
rlabel polysilicon 495 -3232 495 -3232 0 4
rlabel polysilicon 499 -3226 499 -3226 0 1
rlabel polysilicon 499 -3232 499 -3232 0 3
rlabel polysilicon 506 -3226 506 -3226 0 1
rlabel polysilicon 506 -3232 506 -3232 0 3
rlabel polysilicon 513 -3226 513 -3226 0 1
rlabel polysilicon 513 -3232 513 -3232 0 3
rlabel polysilicon 520 -3226 520 -3226 0 1
rlabel polysilicon 520 -3232 520 -3232 0 3
rlabel polysilicon 527 -3226 527 -3226 0 1
rlabel polysilicon 527 -3232 527 -3232 0 3
rlabel polysilicon 534 -3226 534 -3226 0 1
rlabel polysilicon 534 -3232 534 -3232 0 3
rlabel polysilicon 541 -3226 541 -3226 0 1
rlabel polysilicon 541 -3232 541 -3232 0 3
rlabel polysilicon 548 -3226 548 -3226 0 1
rlabel polysilicon 548 -3232 548 -3232 0 3
rlabel polysilicon 555 -3226 555 -3226 0 1
rlabel polysilicon 555 -3232 555 -3232 0 3
rlabel polysilicon 562 -3226 562 -3226 0 1
rlabel polysilicon 562 -3232 562 -3232 0 3
rlabel polysilicon 569 -3226 569 -3226 0 1
rlabel polysilicon 569 -3232 569 -3232 0 3
rlabel polysilicon 576 -3226 576 -3226 0 1
rlabel polysilicon 579 -3226 579 -3226 0 2
rlabel polysilicon 576 -3232 576 -3232 0 3
rlabel polysilicon 579 -3232 579 -3232 0 4
rlabel polysilicon 583 -3226 583 -3226 0 1
rlabel polysilicon 583 -3232 583 -3232 0 3
rlabel polysilicon 590 -3226 590 -3226 0 1
rlabel polysilicon 590 -3232 590 -3232 0 3
rlabel polysilicon 597 -3226 597 -3226 0 1
rlabel polysilicon 597 -3232 597 -3232 0 3
rlabel polysilicon 604 -3226 604 -3226 0 1
rlabel polysilicon 604 -3232 604 -3232 0 3
rlabel polysilicon 611 -3226 611 -3226 0 1
rlabel polysilicon 614 -3226 614 -3226 0 2
rlabel polysilicon 611 -3232 611 -3232 0 3
rlabel polysilicon 614 -3232 614 -3232 0 4
rlabel polysilicon 618 -3226 618 -3226 0 1
rlabel polysilicon 618 -3232 618 -3232 0 3
rlabel polysilicon 625 -3226 625 -3226 0 1
rlabel polysilicon 625 -3232 625 -3232 0 3
rlabel polysilicon 632 -3226 632 -3226 0 1
rlabel polysilicon 632 -3232 632 -3232 0 3
rlabel polysilicon 639 -3226 639 -3226 0 1
rlabel polysilicon 639 -3232 639 -3232 0 3
rlabel polysilicon 646 -3226 646 -3226 0 1
rlabel polysilicon 646 -3232 646 -3232 0 3
rlabel polysilicon 653 -3226 653 -3226 0 1
rlabel polysilicon 653 -3232 653 -3232 0 3
rlabel polysilicon 660 -3226 660 -3226 0 1
rlabel polysilicon 660 -3232 660 -3232 0 3
rlabel polysilicon 667 -3226 667 -3226 0 1
rlabel polysilicon 667 -3232 667 -3232 0 3
rlabel polysilicon 674 -3226 674 -3226 0 1
rlabel polysilicon 677 -3232 677 -3232 0 4
rlabel polysilicon 681 -3226 681 -3226 0 1
rlabel polysilicon 681 -3232 681 -3232 0 3
rlabel polysilicon 688 -3226 688 -3226 0 1
rlabel polysilicon 688 -3232 688 -3232 0 3
rlabel polysilicon 695 -3226 695 -3226 0 1
rlabel polysilicon 695 -3232 695 -3232 0 3
rlabel polysilicon 702 -3226 702 -3226 0 1
rlabel polysilicon 702 -3232 702 -3232 0 3
rlabel polysilicon 709 -3226 709 -3226 0 1
rlabel polysilicon 709 -3232 709 -3232 0 3
rlabel polysilicon 716 -3226 716 -3226 0 1
rlabel polysilicon 716 -3232 716 -3232 0 3
rlabel polysilicon 719 -3232 719 -3232 0 4
rlabel polysilicon 723 -3226 723 -3226 0 1
rlabel polysilicon 723 -3232 723 -3232 0 3
rlabel polysilicon 730 -3226 730 -3226 0 1
rlabel polysilicon 730 -3232 730 -3232 0 3
rlabel polysilicon 737 -3226 737 -3226 0 1
rlabel polysilicon 737 -3232 737 -3232 0 3
rlabel polysilicon 744 -3226 744 -3226 0 1
rlabel polysilicon 747 -3226 747 -3226 0 2
rlabel polysilicon 751 -3226 751 -3226 0 1
rlabel polysilicon 751 -3232 751 -3232 0 3
rlabel polysilicon 758 -3226 758 -3226 0 1
rlabel polysilicon 758 -3232 758 -3232 0 3
rlabel polysilicon 765 -3226 765 -3226 0 1
rlabel polysilicon 768 -3226 768 -3226 0 2
rlabel polysilicon 765 -3232 765 -3232 0 3
rlabel polysilicon 768 -3232 768 -3232 0 4
rlabel polysilicon 772 -3226 772 -3226 0 1
rlabel polysilicon 772 -3232 772 -3232 0 3
rlabel polysilicon 779 -3226 779 -3226 0 1
rlabel polysilicon 779 -3232 779 -3232 0 3
rlabel polysilicon 786 -3226 786 -3226 0 1
rlabel polysilicon 786 -3232 786 -3232 0 3
rlabel polysilicon 793 -3226 793 -3226 0 1
rlabel polysilicon 793 -3232 793 -3232 0 3
rlabel polysilicon 800 -3226 800 -3226 0 1
rlabel polysilicon 800 -3232 800 -3232 0 3
rlabel polysilicon 803 -3232 803 -3232 0 4
rlabel polysilicon 807 -3226 807 -3226 0 1
rlabel polysilicon 807 -3232 807 -3232 0 3
rlabel polysilicon 814 -3226 814 -3226 0 1
rlabel polysilicon 817 -3226 817 -3226 0 2
rlabel polysilicon 817 -3232 817 -3232 0 4
rlabel polysilicon 821 -3226 821 -3226 0 1
rlabel polysilicon 821 -3232 821 -3232 0 3
rlabel polysilicon 828 -3226 828 -3226 0 1
rlabel polysilicon 828 -3232 828 -3232 0 3
rlabel polysilicon 835 -3226 835 -3226 0 1
rlabel polysilicon 835 -3232 835 -3232 0 3
rlabel polysilicon 842 -3226 842 -3226 0 1
rlabel polysilicon 842 -3232 842 -3232 0 3
rlabel polysilicon 849 -3226 849 -3226 0 1
rlabel polysilicon 849 -3232 849 -3232 0 3
rlabel polysilicon 856 -3226 856 -3226 0 1
rlabel polysilicon 856 -3232 856 -3232 0 3
rlabel polysilicon 863 -3226 863 -3226 0 1
rlabel polysilicon 863 -3232 863 -3232 0 3
rlabel polysilicon 873 -3226 873 -3226 0 2
rlabel polysilicon 870 -3232 870 -3232 0 3
rlabel polysilicon 873 -3232 873 -3232 0 4
rlabel polysilicon 877 -3226 877 -3226 0 1
rlabel polysilicon 877 -3232 877 -3232 0 3
rlabel polysilicon 884 -3226 884 -3226 0 1
rlabel polysilicon 884 -3232 884 -3232 0 3
rlabel polysilicon 891 -3226 891 -3226 0 1
rlabel polysilicon 891 -3232 891 -3232 0 3
rlabel polysilicon 898 -3226 898 -3226 0 1
rlabel polysilicon 898 -3232 898 -3232 0 3
rlabel polysilicon 905 -3226 905 -3226 0 1
rlabel polysilicon 905 -3232 905 -3232 0 3
rlabel polysilicon 912 -3226 912 -3226 0 1
rlabel polysilicon 912 -3232 912 -3232 0 3
rlabel polysilicon 919 -3226 919 -3226 0 1
rlabel polysilicon 919 -3232 919 -3232 0 3
rlabel polysilicon 926 -3226 926 -3226 0 1
rlabel polysilicon 926 -3232 926 -3232 0 3
rlabel polysilicon 933 -3226 933 -3226 0 1
rlabel polysilicon 933 -3232 933 -3232 0 3
rlabel polysilicon 940 -3226 940 -3226 0 1
rlabel polysilicon 943 -3226 943 -3226 0 2
rlabel polysilicon 940 -3232 940 -3232 0 3
rlabel polysilicon 943 -3232 943 -3232 0 4
rlabel polysilicon 947 -3226 947 -3226 0 1
rlabel polysilicon 947 -3232 947 -3232 0 3
rlabel polysilicon 954 -3226 954 -3226 0 1
rlabel polysilicon 954 -3232 954 -3232 0 3
rlabel polysilicon 957 -3232 957 -3232 0 4
rlabel polysilicon 961 -3226 961 -3226 0 1
rlabel polysilicon 961 -3232 961 -3232 0 3
rlabel polysilicon 968 -3226 968 -3226 0 1
rlabel polysilicon 968 -3232 968 -3232 0 3
rlabel polysilicon 975 -3226 975 -3226 0 1
rlabel polysilicon 975 -3232 975 -3232 0 3
rlabel polysilicon 985 -3226 985 -3226 0 2
rlabel polysilicon 985 -3232 985 -3232 0 4
rlabel polysilicon 989 -3226 989 -3226 0 1
rlabel polysilicon 989 -3232 989 -3232 0 3
rlabel polysilicon 996 -3226 996 -3226 0 1
rlabel polysilicon 996 -3232 996 -3232 0 3
rlabel polysilicon 1003 -3226 1003 -3226 0 1
rlabel polysilicon 1003 -3232 1003 -3232 0 3
rlabel polysilicon 1010 -3226 1010 -3226 0 1
rlabel polysilicon 1010 -3232 1010 -3232 0 3
rlabel polysilicon 1017 -3226 1017 -3226 0 1
rlabel polysilicon 1017 -3232 1017 -3232 0 3
rlabel polysilicon 1024 -3226 1024 -3226 0 1
rlabel polysilicon 1024 -3232 1024 -3232 0 3
rlabel polysilicon 1031 -3226 1031 -3226 0 1
rlabel polysilicon 1031 -3232 1031 -3232 0 3
rlabel polysilicon 1038 -3226 1038 -3226 0 1
rlabel polysilicon 1038 -3232 1038 -3232 0 3
rlabel polysilicon 1045 -3226 1045 -3226 0 1
rlabel polysilicon 1045 -3232 1045 -3232 0 3
rlabel polysilicon 1052 -3226 1052 -3226 0 1
rlabel polysilicon 1052 -3232 1052 -3232 0 3
rlabel polysilicon 1059 -3226 1059 -3226 0 1
rlabel polysilicon 1059 -3232 1059 -3232 0 3
rlabel polysilicon 1066 -3226 1066 -3226 0 1
rlabel polysilicon 1066 -3232 1066 -3232 0 3
rlabel polysilicon 1073 -3226 1073 -3226 0 1
rlabel polysilicon 1073 -3232 1073 -3232 0 3
rlabel polysilicon 1080 -3226 1080 -3226 0 1
rlabel polysilicon 1080 -3232 1080 -3232 0 3
rlabel polysilicon 1087 -3226 1087 -3226 0 1
rlabel polysilicon 1087 -3232 1087 -3232 0 3
rlabel polysilicon 1094 -3226 1094 -3226 0 1
rlabel polysilicon 1094 -3232 1094 -3232 0 3
rlabel polysilicon 1101 -3226 1101 -3226 0 1
rlabel polysilicon 1101 -3232 1101 -3232 0 3
rlabel polysilicon 1108 -3226 1108 -3226 0 1
rlabel polysilicon 1111 -3226 1111 -3226 0 2
rlabel polysilicon 1108 -3232 1108 -3232 0 3
rlabel polysilicon 1115 -3226 1115 -3226 0 1
rlabel polysilicon 1115 -3232 1115 -3232 0 3
rlabel polysilicon 1122 -3226 1122 -3226 0 1
rlabel polysilicon 1122 -3232 1122 -3232 0 3
rlabel polysilicon 1129 -3226 1129 -3226 0 1
rlabel polysilicon 1129 -3232 1129 -3232 0 3
rlabel polysilicon 1136 -3226 1136 -3226 0 1
rlabel polysilicon 1136 -3232 1136 -3232 0 3
rlabel polysilicon 1143 -3226 1143 -3226 0 1
rlabel polysilicon 1143 -3232 1143 -3232 0 3
rlabel polysilicon 1150 -3226 1150 -3226 0 1
rlabel polysilicon 1150 -3232 1150 -3232 0 3
rlabel polysilicon 1157 -3226 1157 -3226 0 1
rlabel polysilicon 1157 -3232 1157 -3232 0 3
rlabel polysilicon 1164 -3226 1164 -3226 0 1
rlabel polysilicon 1167 -3226 1167 -3226 0 2
rlabel polysilicon 1164 -3232 1164 -3232 0 3
rlabel polysilicon 1167 -3232 1167 -3232 0 4
rlabel polysilicon 1171 -3226 1171 -3226 0 1
rlabel polysilicon 1171 -3232 1171 -3232 0 3
rlabel polysilicon 1178 -3226 1178 -3226 0 1
rlabel polysilicon 1178 -3232 1178 -3232 0 3
rlabel polysilicon 1185 -3226 1185 -3226 0 1
rlabel polysilicon 1185 -3232 1185 -3232 0 3
rlabel polysilicon 1192 -3226 1192 -3226 0 1
rlabel polysilicon 1192 -3232 1192 -3232 0 3
rlabel polysilicon 1199 -3226 1199 -3226 0 1
rlabel polysilicon 1199 -3232 1199 -3232 0 3
rlabel polysilicon 1206 -3226 1206 -3226 0 1
rlabel polysilicon 1206 -3232 1206 -3232 0 3
rlabel polysilicon 1213 -3226 1213 -3226 0 1
rlabel polysilicon 1216 -3226 1216 -3226 0 2
rlabel polysilicon 1213 -3232 1213 -3232 0 3
rlabel polysilicon 1216 -3232 1216 -3232 0 4
rlabel polysilicon 1220 -3226 1220 -3226 0 1
rlabel polysilicon 1220 -3232 1220 -3232 0 3
rlabel polysilicon 1227 -3226 1227 -3226 0 1
rlabel polysilicon 1227 -3232 1227 -3232 0 3
rlabel polysilicon 1234 -3232 1234 -3232 0 3
rlabel polysilicon 1237 -3232 1237 -3232 0 4
rlabel polysilicon 1241 -3226 1241 -3226 0 1
rlabel polysilicon 1241 -3232 1241 -3232 0 3
rlabel polysilicon 1248 -3226 1248 -3226 0 1
rlabel polysilicon 1248 -3232 1248 -3232 0 3
rlabel polysilicon 1255 -3226 1255 -3226 0 1
rlabel polysilicon 1258 -3226 1258 -3226 0 2
rlabel polysilicon 1255 -3232 1255 -3232 0 3
rlabel polysilicon 1262 -3226 1262 -3226 0 1
rlabel polysilicon 1262 -3232 1262 -3232 0 3
rlabel polysilicon 1269 -3226 1269 -3226 0 1
rlabel polysilicon 1269 -3232 1269 -3232 0 3
rlabel polysilicon 1276 -3226 1276 -3226 0 1
rlabel polysilicon 1276 -3232 1276 -3232 0 3
rlabel polysilicon 1283 -3226 1283 -3226 0 1
rlabel polysilicon 1283 -3232 1283 -3232 0 3
rlabel polysilicon 1290 -3226 1290 -3226 0 1
rlabel polysilicon 1290 -3232 1290 -3232 0 3
rlabel polysilicon 1297 -3226 1297 -3226 0 1
rlabel polysilicon 1297 -3232 1297 -3232 0 3
rlabel polysilicon 1304 -3226 1304 -3226 0 1
rlabel polysilicon 1304 -3232 1304 -3232 0 3
rlabel polysilicon 1311 -3226 1311 -3226 0 1
rlabel polysilicon 1311 -3232 1311 -3232 0 3
rlabel polysilicon 1318 -3226 1318 -3226 0 1
rlabel polysilicon 1318 -3232 1318 -3232 0 3
rlabel polysilicon 1325 -3226 1325 -3226 0 1
rlabel polysilicon 1325 -3232 1325 -3232 0 3
rlabel polysilicon 1332 -3226 1332 -3226 0 1
rlabel polysilicon 1332 -3232 1332 -3232 0 3
rlabel polysilicon 1339 -3226 1339 -3226 0 1
rlabel polysilicon 1339 -3232 1339 -3232 0 3
rlabel polysilicon 1346 -3226 1346 -3226 0 1
rlabel polysilicon 1346 -3232 1346 -3232 0 3
rlabel polysilicon 1353 -3226 1353 -3226 0 1
rlabel polysilicon 1356 -3226 1356 -3226 0 2
rlabel polysilicon 1353 -3232 1353 -3232 0 3
rlabel polysilicon 1360 -3226 1360 -3226 0 1
rlabel polysilicon 1360 -3232 1360 -3232 0 3
rlabel polysilicon 1367 -3226 1367 -3226 0 1
rlabel polysilicon 1367 -3232 1367 -3232 0 3
rlabel polysilicon 1374 -3226 1374 -3226 0 1
rlabel polysilicon 1374 -3232 1374 -3232 0 3
rlabel polysilicon 1381 -3226 1381 -3226 0 1
rlabel polysilicon 1381 -3232 1381 -3232 0 3
rlabel polysilicon 1388 -3226 1388 -3226 0 1
rlabel polysilicon 1388 -3232 1388 -3232 0 3
rlabel polysilicon 1395 -3226 1395 -3226 0 1
rlabel polysilicon 1395 -3232 1395 -3232 0 3
rlabel polysilicon 1402 -3226 1402 -3226 0 1
rlabel polysilicon 1402 -3232 1402 -3232 0 3
rlabel polysilicon 1409 -3226 1409 -3226 0 1
rlabel polysilicon 1409 -3232 1409 -3232 0 3
rlabel polysilicon 1416 -3226 1416 -3226 0 1
rlabel polysilicon 1416 -3232 1416 -3232 0 3
rlabel polysilicon 1423 -3226 1423 -3226 0 1
rlabel polysilicon 1423 -3232 1423 -3232 0 3
rlabel polysilicon 1430 -3226 1430 -3226 0 1
rlabel polysilicon 1430 -3232 1430 -3232 0 3
rlabel polysilicon 1437 -3226 1437 -3226 0 1
rlabel polysilicon 1437 -3232 1437 -3232 0 3
rlabel polysilicon 1444 -3226 1444 -3226 0 1
rlabel polysilicon 1444 -3232 1444 -3232 0 3
rlabel polysilicon 1451 -3226 1451 -3226 0 1
rlabel polysilicon 1451 -3232 1451 -3232 0 3
rlabel polysilicon 1458 -3226 1458 -3226 0 1
rlabel polysilicon 1461 -3226 1461 -3226 0 2
rlabel polysilicon 1458 -3232 1458 -3232 0 3
rlabel polysilicon 1465 -3226 1465 -3226 0 1
rlabel polysilicon 1465 -3232 1465 -3232 0 3
rlabel polysilicon 1472 -3226 1472 -3226 0 1
rlabel polysilicon 1472 -3232 1472 -3232 0 3
rlabel polysilicon 1479 -3226 1479 -3226 0 1
rlabel polysilicon 1479 -3232 1479 -3232 0 3
rlabel polysilicon 1486 -3226 1486 -3226 0 1
rlabel polysilicon 1486 -3232 1486 -3232 0 3
rlabel polysilicon 1493 -3226 1493 -3226 0 1
rlabel polysilicon 1493 -3232 1493 -3232 0 3
rlabel polysilicon 1500 -3226 1500 -3226 0 1
rlabel polysilicon 1500 -3232 1500 -3232 0 3
rlabel polysilicon 1507 -3226 1507 -3226 0 1
rlabel polysilicon 1507 -3232 1507 -3232 0 3
rlabel polysilicon 1514 -3226 1514 -3226 0 1
rlabel polysilicon 1514 -3232 1514 -3232 0 3
rlabel polysilicon 1521 -3226 1521 -3226 0 1
rlabel polysilicon 1521 -3232 1521 -3232 0 3
rlabel polysilicon 1528 -3226 1528 -3226 0 1
rlabel polysilicon 1528 -3232 1528 -3232 0 3
rlabel polysilicon 1535 -3226 1535 -3226 0 1
rlabel polysilicon 1535 -3232 1535 -3232 0 3
rlabel polysilicon 1542 -3226 1542 -3226 0 1
rlabel polysilicon 1542 -3232 1542 -3232 0 3
rlabel polysilicon 1549 -3226 1549 -3226 0 1
rlabel polysilicon 1549 -3232 1549 -3232 0 3
rlabel polysilicon 1556 -3226 1556 -3226 0 1
rlabel polysilicon 1556 -3232 1556 -3232 0 3
rlabel polysilicon 1563 -3226 1563 -3226 0 1
rlabel polysilicon 1563 -3232 1563 -3232 0 3
rlabel polysilicon 1570 -3226 1570 -3226 0 1
rlabel polysilicon 1570 -3232 1570 -3232 0 3
rlabel polysilicon 1577 -3226 1577 -3226 0 1
rlabel polysilicon 1580 -3232 1580 -3232 0 4
rlabel polysilicon 1584 -3226 1584 -3226 0 1
rlabel polysilicon 1584 -3232 1584 -3232 0 3
rlabel polysilicon 1591 -3226 1591 -3226 0 1
rlabel polysilicon 1591 -3232 1591 -3232 0 3
rlabel polysilicon 1598 -3226 1598 -3226 0 1
rlabel polysilicon 1598 -3232 1598 -3232 0 3
rlabel polysilicon 1605 -3226 1605 -3226 0 1
rlabel polysilicon 1605 -3232 1605 -3232 0 3
rlabel polysilicon 1612 -3226 1612 -3226 0 1
rlabel polysilicon 1612 -3232 1612 -3232 0 3
rlabel polysilicon 1619 -3226 1619 -3226 0 1
rlabel polysilicon 1619 -3232 1619 -3232 0 3
rlabel polysilicon 1626 -3226 1626 -3226 0 1
rlabel polysilicon 1626 -3232 1626 -3232 0 3
rlabel polysilicon 1633 -3226 1633 -3226 0 1
rlabel polysilicon 1633 -3232 1633 -3232 0 3
rlabel polysilicon 1640 -3226 1640 -3226 0 1
rlabel polysilicon 1643 -3226 1643 -3226 0 2
rlabel polysilicon 1640 -3232 1640 -3232 0 3
rlabel polysilicon 1643 -3232 1643 -3232 0 4
rlabel polysilicon 1647 -3226 1647 -3226 0 1
rlabel polysilicon 1650 -3226 1650 -3226 0 2
rlabel polysilicon 1647 -3232 1647 -3232 0 3
rlabel polysilicon 1650 -3232 1650 -3232 0 4
rlabel polysilicon 1654 -3226 1654 -3226 0 1
rlabel polysilicon 1657 -3226 1657 -3226 0 2
rlabel polysilicon 1654 -3232 1654 -3232 0 3
rlabel polysilicon 1661 -3226 1661 -3226 0 1
rlabel polysilicon 1661 -3232 1661 -3232 0 3
rlabel polysilicon 1671 -3226 1671 -3226 0 2
rlabel polysilicon 1671 -3232 1671 -3232 0 4
rlabel polysilicon 1675 -3226 1675 -3226 0 1
rlabel polysilicon 1675 -3232 1675 -3232 0 3
rlabel polysilicon 1682 -3226 1682 -3226 0 1
rlabel polysilicon 1685 -3226 1685 -3226 0 2
rlabel polysilicon 1682 -3232 1682 -3232 0 3
rlabel polysilicon 1685 -3232 1685 -3232 0 4
rlabel polysilicon 1689 -3226 1689 -3226 0 1
rlabel polysilicon 1689 -3232 1689 -3232 0 3
rlabel polysilicon 1696 -3226 1696 -3226 0 1
rlabel polysilicon 1696 -3232 1696 -3232 0 3
rlabel polysilicon 1703 -3226 1703 -3226 0 1
rlabel polysilicon 1703 -3232 1703 -3232 0 3
rlabel polysilicon 1710 -3226 1710 -3226 0 1
rlabel polysilicon 1710 -3232 1710 -3232 0 3
rlabel polysilicon 1717 -3226 1717 -3226 0 1
rlabel polysilicon 1717 -3232 1717 -3232 0 3
rlabel polysilicon 1724 -3226 1724 -3226 0 1
rlabel polysilicon 1724 -3232 1724 -3232 0 3
rlabel polysilicon 1731 -3226 1731 -3226 0 1
rlabel polysilicon 1731 -3232 1731 -3232 0 3
rlabel polysilicon 1738 -3226 1738 -3226 0 1
rlabel polysilicon 1738 -3232 1738 -3232 0 3
rlabel polysilicon 1745 -3226 1745 -3226 0 1
rlabel polysilicon 1745 -3232 1745 -3232 0 3
rlabel polysilicon 1752 -3226 1752 -3226 0 1
rlabel polysilicon 1752 -3232 1752 -3232 0 3
rlabel polysilicon 1759 -3226 1759 -3226 0 1
rlabel polysilicon 1759 -3232 1759 -3232 0 3
rlabel polysilicon 1766 -3226 1766 -3226 0 1
rlabel polysilicon 1766 -3232 1766 -3232 0 3
rlabel polysilicon 1773 -3226 1773 -3226 0 1
rlabel polysilicon 1773 -3232 1773 -3232 0 3
rlabel polysilicon 1780 -3226 1780 -3226 0 1
rlabel polysilicon 1780 -3232 1780 -3232 0 3
rlabel polysilicon 1808 -3226 1808 -3226 0 1
rlabel polysilicon 1808 -3232 1808 -3232 0 3
rlabel polysilicon 1815 -3226 1815 -3226 0 1
rlabel polysilicon 1815 -3232 1815 -3232 0 3
rlabel polysilicon 1822 -3226 1822 -3226 0 1
rlabel polysilicon 1822 -3232 1822 -3232 0 3
rlabel polysilicon 1850 -3226 1850 -3226 0 1
rlabel polysilicon 1853 -3226 1853 -3226 0 2
rlabel polysilicon 1850 -3232 1850 -3232 0 3
rlabel polysilicon 1853 -3232 1853 -3232 0 4
rlabel polysilicon 1857 -3226 1857 -3226 0 1
rlabel polysilicon 1857 -3232 1857 -3232 0 3
rlabel polysilicon 1864 -3226 1864 -3226 0 1
rlabel polysilicon 1864 -3232 1864 -3232 0 3
rlabel polysilicon 1878 -3226 1878 -3226 0 1
rlabel polysilicon 1878 -3232 1878 -3232 0 3
rlabel polysilicon 1885 -3226 1885 -3226 0 1
rlabel polysilicon 1885 -3232 1885 -3232 0 3
rlabel polysilicon 1892 -3226 1892 -3226 0 1
rlabel polysilicon 1892 -3232 1892 -3232 0 3
rlabel polysilicon 1906 -3226 1906 -3226 0 1
rlabel polysilicon 1906 -3232 1906 -3232 0 3
rlabel polysilicon 1920 -3226 1920 -3226 0 1
rlabel polysilicon 1920 -3232 1920 -3232 0 3
rlabel polysilicon 1962 -3226 1962 -3226 0 1
rlabel polysilicon 1965 -3226 1965 -3226 0 2
rlabel polysilicon 1962 -3232 1962 -3232 0 3
rlabel polysilicon 1965 -3232 1965 -3232 0 4
rlabel polysilicon 1969 -3226 1969 -3226 0 1
rlabel polysilicon 1969 -3232 1969 -3232 0 3
rlabel polysilicon 1976 -3226 1976 -3226 0 1
rlabel polysilicon 1976 -3232 1976 -3232 0 3
rlabel polysilicon 1983 -3226 1983 -3226 0 1
rlabel polysilicon 1983 -3232 1983 -3232 0 3
rlabel polysilicon 2018 -3226 2018 -3226 0 1
rlabel polysilicon 2018 -3232 2018 -3232 0 3
rlabel polysilicon 2046 -3226 2046 -3226 0 1
rlabel polysilicon 2046 -3232 2046 -3232 0 3
rlabel polysilicon 142 -3329 142 -3329 0 1
rlabel polysilicon 142 -3335 142 -3335 0 3
rlabel polysilicon 163 -3329 163 -3329 0 1
rlabel polysilicon 163 -3335 163 -3335 0 3
rlabel polysilicon 170 -3329 170 -3329 0 1
rlabel polysilicon 170 -3335 170 -3335 0 3
rlabel polysilicon 177 -3329 177 -3329 0 1
rlabel polysilicon 177 -3335 177 -3335 0 3
rlabel polysilicon 184 -3329 184 -3329 0 1
rlabel polysilicon 184 -3335 184 -3335 0 3
rlabel polysilicon 191 -3329 191 -3329 0 1
rlabel polysilicon 191 -3335 191 -3335 0 3
rlabel polysilicon 198 -3329 198 -3329 0 1
rlabel polysilicon 198 -3335 198 -3335 0 3
rlabel polysilicon 205 -3329 205 -3329 0 1
rlabel polysilicon 205 -3335 205 -3335 0 3
rlabel polysilicon 215 -3329 215 -3329 0 2
rlabel polysilicon 212 -3335 212 -3335 0 3
rlabel polysilicon 215 -3335 215 -3335 0 4
rlabel polysilicon 219 -3329 219 -3329 0 1
rlabel polysilicon 219 -3335 219 -3335 0 3
rlabel polysilicon 226 -3329 226 -3329 0 1
rlabel polysilicon 229 -3329 229 -3329 0 2
rlabel polysilicon 236 -3335 236 -3335 0 4
rlabel polysilicon 240 -3329 240 -3329 0 1
rlabel polysilicon 240 -3335 240 -3335 0 3
rlabel polysilicon 247 -3329 247 -3329 0 1
rlabel polysilicon 247 -3335 247 -3335 0 3
rlabel polysilicon 254 -3329 254 -3329 0 1
rlabel polysilicon 257 -3329 257 -3329 0 2
rlabel polysilicon 257 -3335 257 -3335 0 4
rlabel polysilicon 261 -3329 261 -3329 0 1
rlabel polysilicon 261 -3335 261 -3335 0 3
rlabel polysilicon 268 -3329 268 -3329 0 1
rlabel polysilicon 268 -3335 268 -3335 0 3
rlabel polysilicon 275 -3329 275 -3329 0 1
rlabel polysilicon 275 -3335 275 -3335 0 3
rlabel polysilicon 282 -3329 282 -3329 0 1
rlabel polysilicon 282 -3335 282 -3335 0 3
rlabel polysilicon 289 -3329 289 -3329 0 1
rlabel polysilicon 289 -3335 289 -3335 0 3
rlabel polysilicon 296 -3329 296 -3329 0 1
rlabel polysilicon 296 -3335 296 -3335 0 3
rlabel polysilicon 303 -3329 303 -3329 0 1
rlabel polysilicon 303 -3335 303 -3335 0 3
rlabel polysilicon 310 -3329 310 -3329 0 1
rlabel polysilicon 310 -3335 310 -3335 0 3
rlabel polysilicon 317 -3329 317 -3329 0 1
rlabel polysilicon 317 -3335 317 -3335 0 3
rlabel polysilicon 324 -3329 324 -3329 0 1
rlabel polysilicon 324 -3335 324 -3335 0 3
rlabel polysilicon 331 -3329 331 -3329 0 1
rlabel polysilicon 331 -3335 331 -3335 0 3
rlabel polysilicon 338 -3329 338 -3329 0 1
rlabel polysilicon 338 -3335 338 -3335 0 3
rlabel polysilicon 345 -3329 345 -3329 0 1
rlabel polysilicon 345 -3335 345 -3335 0 3
rlabel polysilicon 352 -3329 352 -3329 0 1
rlabel polysilicon 352 -3335 352 -3335 0 3
rlabel polysilicon 359 -3329 359 -3329 0 1
rlabel polysilicon 359 -3335 359 -3335 0 3
rlabel polysilicon 366 -3329 366 -3329 0 1
rlabel polysilicon 366 -3335 366 -3335 0 3
rlabel polysilicon 373 -3329 373 -3329 0 1
rlabel polysilicon 373 -3335 373 -3335 0 3
rlabel polysilicon 380 -3329 380 -3329 0 1
rlabel polysilicon 383 -3329 383 -3329 0 2
rlabel polysilicon 380 -3335 380 -3335 0 3
rlabel polysilicon 383 -3335 383 -3335 0 4
rlabel polysilicon 387 -3329 387 -3329 0 1
rlabel polysilicon 387 -3335 387 -3335 0 3
rlabel polysilicon 394 -3329 394 -3329 0 1
rlabel polysilicon 394 -3335 394 -3335 0 3
rlabel polysilicon 401 -3329 401 -3329 0 1
rlabel polysilicon 401 -3335 401 -3335 0 3
rlabel polysilicon 408 -3329 408 -3329 0 1
rlabel polysilicon 408 -3335 408 -3335 0 3
rlabel polysilicon 415 -3329 415 -3329 0 1
rlabel polysilicon 415 -3335 415 -3335 0 3
rlabel polysilicon 418 -3335 418 -3335 0 4
rlabel polysilicon 422 -3329 422 -3329 0 1
rlabel polysilicon 422 -3335 422 -3335 0 3
rlabel polysilicon 429 -3329 429 -3329 0 1
rlabel polysilicon 429 -3335 429 -3335 0 3
rlabel polysilicon 436 -3329 436 -3329 0 1
rlabel polysilicon 436 -3335 436 -3335 0 3
rlabel polysilicon 443 -3329 443 -3329 0 1
rlabel polysilicon 443 -3335 443 -3335 0 3
rlabel polysilicon 450 -3329 450 -3329 0 1
rlabel polysilicon 450 -3335 450 -3335 0 3
rlabel polysilicon 457 -3329 457 -3329 0 1
rlabel polysilicon 457 -3335 457 -3335 0 3
rlabel polysilicon 464 -3329 464 -3329 0 1
rlabel polysilicon 464 -3335 464 -3335 0 3
rlabel polysilicon 471 -3329 471 -3329 0 1
rlabel polysilicon 471 -3335 471 -3335 0 3
rlabel polysilicon 478 -3329 478 -3329 0 1
rlabel polysilicon 478 -3335 478 -3335 0 3
rlabel polysilicon 485 -3329 485 -3329 0 1
rlabel polysilicon 485 -3335 485 -3335 0 3
rlabel polysilicon 492 -3329 492 -3329 0 1
rlabel polysilicon 492 -3335 492 -3335 0 3
rlabel polysilicon 499 -3329 499 -3329 0 1
rlabel polysilicon 499 -3335 499 -3335 0 3
rlabel polysilicon 506 -3329 506 -3329 0 1
rlabel polysilicon 506 -3335 506 -3335 0 3
rlabel polysilicon 513 -3329 513 -3329 0 1
rlabel polysilicon 513 -3335 513 -3335 0 3
rlabel polysilicon 520 -3329 520 -3329 0 1
rlabel polysilicon 520 -3335 520 -3335 0 3
rlabel polysilicon 527 -3329 527 -3329 0 1
rlabel polysilicon 527 -3335 527 -3335 0 3
rlabel polysilicon 534 -3329 534 -3329 0 1
rlabel polysilicon 537 -3329 537 -3329 0 2
rlabel polysilicon 534 -3335 534 -3335 0 3
rlabel polysilicon 537 -3335 537 -3335 0 4
rlabel polysilicon 541 -3329 541 -3329 0 1
rlabel polysilicon 541 -3335 541 -3335 0 3
rlabel polysilicon 548 -3329 548 -3329 0 1
rlabel polysilicon 548 -3335 548 -3335 0 3
rlabel polysilicon 555 -3329 555 -3329 0 1
rlabel polysilicon 555 -3335 555 -3335 0 3
rlabel polysilicon 562 -3329 562 -3329 0 1
rlabel polysilicon 562 -3335 562 -3335 0 3
rlabel polysilicon 569 -3329 569 -3329 0 1
rlabel polysilicon 569 -3335 569 -3335 0 3
rlabel polysilicon 576 -3329 576 -3329 0 1
rlabel polysilicon 583 -3329 583 -3329 0 1
rlabel polysilicon 583 -3335 583 -3335 0 3
rlabel polysilicon 590 -3329 590 -3329 0 1
rlabel polysilicon 590 -3335 590 -3335 0 3
rlabel polysilicon 597 -3329 597 -3329 0 1
rlabel polysilicon 600 -3329 600 -3329 0 2
rlabel polysilicon 597 -3335 597 -3335 0 3
rlabel polysilicon 600 -3335 600 -3335 0 4
rlabel polysilicon 604 -3329 604 -3329 0 1
rlabel polysilicon 604 -3335 604 -3335 0 3
rlabel polysilicon 611 -3329 611 -3329 0 1
rlabel polysilicon 611 -3335 611 -3335 0 3
rlabel polysilicon 618 -3329 618 -3329 0 1
rlabel polysilicon 618 -3335 618 -3335 0 3
rlabel polysilicon 625 -3329 625 -3329 0 1
rlabel polysilicon 625 -3335 625 -3335 0 3
rlabel polysilicon 632 -3329 632 -3329 0 1
rlabel polysilicon 632 -3335 632 -3335 0 3
rlabel polysilicon 639 -3329 639 -3329 0 1
rlabel polysilicon 642 -3329 642 -3329 0 2
rlabel polysilicon 646 -3329 646 -3329 0 1
rlabel polysilicon 646 -3335 646 -3335 0 3
rlabel polysilicon 653 -3329 653 -3329 0 1
rlabel polysilicon 653 -3335 653 -3335 0 3
rlabel polysilicon 660 -3329 660 -3329 0 1
rlabel polysilicon 660 -3335 660 -3335 0 3
rlabel polysilicon 667 -3329 667 -3329 0 1
rlabel polysilicon 667 -3335 667 -3335 0 3
rlabel polysilicon 674 -3329 674 -3329 0 1
rlabel polysilicon 674 -3335 674 -3335 0 3
rlabel polysilicon 681 -3329 681 -3329 0 1
rlabel polysilicon 681 -3335 681 -3335 0 3
rlabel polysilicon 688 -3329 688 -3329 0 1
rlabel polysilicon 688 -3335 688 -3335 0 3
rlabel polysilicon 695 -3329 695 -3329 0 1
rlabel polysilicon 695 -3335 695 -3335 0 3
rlabel polysilicon 702 -3329 702 -3329 0 1
rlabel polysilicon 702 -3335 702 -3335 0 3
rlabel polysilicon 709 -3329 709 -3329 0 1
rlabel polysilicon 709 -3335 709 -3335 0 3
rlabel polysilicon 716 -3329 716 -3329 0 1
rlabel polysilicon 716 -3335 716 -3335 0 3
rlabel polysilicon 726 -3329 726 -3329 0 2
rlabel polysilicon 723 -3335 723 -3335 0 3
rlabel polysilicon 733 -3329 733 -3329 0 2
rlabel polysilicon 730 -3335 730 -3335 0 3
rlabel polysilicon 737 -3329 737 -3329 0 1
rlabel polysilicon 737 -3335 737 -3335 0 3
rlabel polysilicon 744 -3329 744 -3329 0 1
rlabel polysilicon 744 -3335 744 -3335 0 3
rlabel polysilicon 751 -3329 751 -3329 0 1
rlabel polysilicon 751 -3335 751 -3335 0 3
rlabel polysilicon 758 -3329 758 -3329 0 1
rlabel polysilicon 758 -3335 758 -3335 0 3
rlabel polysilicon 765 -3329 765 -3329 0 1
rlabel polysilicon 765 -3335 765 -3335 0 3
rlabel polysilicon 772 -3329 772 -3329 0 1
rlabel polysilicon 772 -3335 772 -3335 0 3
rlabel polysilicon 779 -3329 779 -3329 0 1
rlabel polysilicon 782 -3329 782 -3329 0 2
rlabel polysilicon 779 -3335 779 -3335 0 3
rlabel polysilicon 786 -3329 786 -3329 0 1
rlabel polysilicon 786 -3335 786 -3335 0 3
rlabel polysilicon 793 -3329 793 -3329 0 1
rlabel polysilicon 793 -3335 793 -3335 0 3
rlabel polysilicon 800 -3329 800 -3329 0 1
rlabel polysilicon 800 -3335 800 -3335 0 3
rlabel polysilicon 807 -3329 807 -3329 0 1
rlabel polysilicon 807 -3335 807 -3335 0 3
rlabel polysilicon 814 -3329 814 -3329 0 1
rlabel polysilicon 814 -3335 814 -3335 0 3
rlabel polysilicon 821 -3329 821 -3329 0 1
rlabel polysilicon 821 -3335 821 -3335 0 3
rlabel polysilicon 828 -3329 828 -3329 0 1
rlabel polysilicon 828 -3335 828 -3335 0 3
rlabel polysilicon 835 -3329 835 -3329 0 1
rlabel polysilicon 835 -3335 835 -3335 0 3
rlabel polysilicon 842 -3329 842 -3329 0 1
rlabel polysilicon 842 -3335 842 -3335 0 3
rlabel polysilicon 849 -3329 849 -3329 0 1
rlabel polysilicon 849 -3335 849 -3335 0 3
rlabel polysilicon 852 -3335 852 -3335 0 4
rlabel polysilicon 856 -3329 856 -3329 0 1
rlabel polysilicon 856 -3335 856 -3335 0 3
rlabel polysilicon 863 -3329 863 -3329 0 1
rlabel polysilicon 863 -3335 863 -3335 0 3
rlabel polysilicon 870 -3329 870 -3329 0 1
rlabel polysilicon 870 -3335 870 -3335 0 3
rlabel polysilicon 877 -3329 877 -3329 0 1
rlabel polysilicon 877 -3335 877 -3335 0 3
rlabel polysilicon 884 -3329 884 -3329 0 1
rlabel polysilicon 884 -3335 884 -3335 0 3
rlabel polysilicon 891 -3329 891 -3329 0 1
rlabel polysilicon 891 -3335 891 -3335 0 3
rlabel polysilicon 898 -3329 898 -3329 0 1
rlabel polysilicon 898 -3335 898 -3335 0 3
rlabel polysilicon 905 -3329 905 -3329 0 1
rlabel polysilicon 905 -3335 905 -3335 0 3
rlabel polysilicon 912 -3329 912 -3329 0 1
rlabel polysilicon 912 -3335 912 -3335 0 3
rlabel polysilicon 919 -3329 919 -3329 0 1
rlabel polysilicon 919 -3335 919 -3335 0 3
rlabel polysilicon 926 -3329 926 -3329 0 1
rlabel polysilicon 929 -3329 929 -3329 0 2
rlabel polysilicon 926 -3335 926 -3335 0 3
rlabel polysilicon 933 -3329 933 -3329 0 1
rlabel polysilicon 933 -3335 933 -3335 0 3
rlabel polysilicon 940 -3329 940 -3329 0 1
rlabel polysilicon 940 -3335 940 -3335 0 3
rlabel polysilicon 947 -3329 947 -3329 0 1
rlabel polysilicon 947 -3335 947 -3335 0 3
rlabel polysilicon 957 -3329 957 -3329 0 2
rlabel polysilicon 954 -3335 954 -3335 0 3
rlabel polysilicon 957 -3335 957 -3335 0 4
rlabel polysilicon 961 -3329 961 -3329 0 1
rlabel polysilicon 961 -3335 961 -3335 0 3
rlabel polysilicon 968 -3329 968 -3329 0 1
rlabel polysilicon 968 -3335 968 -3335 0 3
rlabel polysilicon 971 -3335 971 -3335 0 4
rlabel polysilicon 978 -3329 978 -3329 0 2
rlabel polysilicon 975 -3335 975 -3335 0 3
rlabel polysilicon 978 -3335 978 -3335 0 4
rlabel polysilicon 982 -3329 982 -3329 0 1
rlabel polysilicon 982 -3335 982 -3335 0 3
rlabel polysilicon 989 -3329 989 -3329 0 1
rlabel polysilicon 992 -3329 992 -3329 0 2
rlabel polysilicon 989 -3335 989 -3335 0 3
rlabel polysilicon 996 -3329 996 -3329 0 1
rlabel polysilicon 996 -3335 996 -3335 0 3
rlabel polysilicon 1003 -3329 1003 -3329 0 1
rlabel polysilicon 1003 -3335 1003 -3335 0 3
rlabel polysilicon 1010 -3329 1010 -3329 0 1
rlabel polysilicon 1010 -3335 1010 -3335 0 3
rlabel polysilicon 1017 -3329 1017 -3329 0 1
rlabel polysilicon 1017 -3335 1017 -3335 0 3
rlabel polysilicon 1024 -3329 1024 -3329 0 1
rlabel polysilicon 1024 -3335 1024 -3335 0 3
rlabel polysilicon 1031 -3329 1031 -3329 0 1
rlabel polysilicon 1031 -3335 1031 -3335 0 3
rlabel polysilicon 1038 -3329 1038 -3329 0 1
rlabel polysilicon 1038 -3335 1038 -3335 0 3
rlabel polysilicon 1045 -3329 1045 -3329 0 1
rlabel polysilicon 1045 -3335 1045 -3335 0 3
rlabel polysilicon 1052 -3329 1052 -3329 0 1
rlabel polysilicon 1052 -3335 1052 -3335 0 3
rlabel polysilicon 1059 -3329 1059 -3329 0 1
rlabel polysilicon 1059 -3335 1059 -3335 0 3
rlabel polysilicon 1066 -3329 1066 -3329 0 1
rlabel polysilicon 1069 -3329 1069 -3329 0 2
rlabel polysilicon 1066 -3335 1066 -3335 0 3
rlabel polysilicon 1073 -3329 1073 -3329 0 1
rlabel polysilicon 1073 -3335 1073 -3335 0 3
rlabel polysilicon 1080 -3329 1080 -3329 0 1
rlabel polysilicon 1080 -3335 1080 -3335 0 3
rlabel polysilicon 1083 -3335 1083 -3335 0 4
rlabel polysilicon 1087 -3329 1087 -3329 0 1
rlabel polysilicon 1087 -3335 1087 -3335 0 3
rlabel polysilicon 1094 -3329 1094 -3329 0 1
rlabel polysilicon 1094 -3335 1094 -3335 0 3
rlabel polysilicon 1097 -3335 1097 -3335 0 4
rlabel polysilicon 1104 -3329 1104 -3329 0 2
rlabel polysilicon 1104 -3335 1104 -3335 0 4
rlabel polysilicon 1108 -3329 1108 -3329 0 1
rlabel polysilicon 1108 -3335 1108 -3335 0 3
rlabel polysilicon 1115 -3329 1115 -3329 0 1
rlabel polysilicon 1115 -3335 1115 -3335 0 3
rlabel polysilicon 1122 -3329 1122 -3329 0 1
rlabel polysilicon 1122 -3335 1122 -3335 0 3
rlabel polysilicon 1129 -3329 1129 -3329 0 1
rlabel polysilicon 1129 -3335 1129 -3335 0 3
rlabel polysilicon 1136 -3329 1136 -3329 0 1
rlabel polysilicon 1136 -3335 1136 -3335 0 3
rlabel polysilicon 1143 -3329 1143 -3329 0 1
rlabel polysilicon 1143 -3335 1143 -3335 0 3
rlabel polysilicon 1150 -3329 1150 -3329 0 1
rlabel polysilicon 1150 -3335 1150 -3335 0 3
rlabel polysilicon 1157 -3329 1157 -3329 0 1
rlabel polysilicon 1157 -3335 1157 -3335 0 3
rlabel polysilicon 1164 -3329 1164 -3329 0 1
rlabel polysilicon 1164 -3335 1164 -3335 0 3
rlabel polysilicon 1171 -3329 1171 -3329 0 1
rlabel polysilicon 1171 -3335 1171 -3335 0 3
rlabel polysilicon 1178 -3329 1178 -3329 0 1
rlabel polysilicon 1178 -3335 1178 -3335 0 3
rlabel polysilicon 1185 -3329 1185 -3329 0 1
rlabel polysilicon 1185 -3335 1185 -3335 0 3
rlabel polysilicon 1192 -3329 1192 -3329 0 1
rlabel polysilicon 1192 -3335 1192 -3335 0 3
rlabel polysilicon 1199 -3329 1199 -3329 0 1
rlabel polysilicon 1199 -3335 1199 -3335 0 3
rlabel polysilicon 1206 -3329 1206 -3329 0 1
rlabel polysilicon 1206 -3335 1206 -3335 0 3
rlabel polysilicon 1216 -3329 1216 -3329 0 2
rlabel polysilicon 1213 -3335 1213 -3335 0 3
rlabel polysilicon 1216 -3335 1216 -3335 0 4
rlabel polysilicon 1220 -3329 1220 -3329 0 1
rlabel polysilicon 1220 -3335 1220 -3335 0 3
rlabel polysilicon 1227 -3329 1227 -3329 0 1
rlabel polysilicon 1227 -3335 1227 -3335 0 3
rlabel polysilicon 1234 -3329 1234 -3329 0 1
rlabel polysilicon 1237 -3329 1237 -3329 0 2
rlabel polysilicon 1234 -3335 1234 -3335 0 3
rlabel polysilicon 1237 -3335 1237 -3335 0 4
rlabel polysilicon 1241 -3329 1241 -3329 0 1
rlabel polysilicon 1241 -3335 1241 -3335 0 3
rlabel polysilicon 1248 -3329 1248 -3329 0 1
rlabel polysilicon 1248 -3335 1248 -3335 0 3
rlabel polysilicon 1255 -3329 1255 -3329 0 1
rlabel polysilicon 1255 -3335 1255 -3335 0 3
rlabel polysilicon 1262 -3329 1262 -3329 0 1
rlabel polysilicon 1262 -3335 1262 -3335 0 3
rlabel polysilicon 1269 -3329 1269 -3329 0 1
rlabel polysilicon 1269 -3335 1269 -3335 0 3
rlabel polysilicon 1272 -3335 1272 -3335 0 4
rlabel polysilicon 1276 -3329 1276 -3329 0 1
rlabel polysilicon 1276 -3335 1276 -3335 0 3
rlabel polysilicon 1283 -3329 1283 -3329 0 1
rlabel polysilicon 1283 -3335 1283 -3335 0 3
rlabel polysilicon 1290 -3329 1290 -3329 0 1
rlabel polysilicon 1290 -3335 1290 -3335 0 3
rlabel polysilicon 1297 -3329 1297 -3329 0 1
rlabel polysilicon 1297 -3335 1297 -3335 0 3
rlabel polysilicon 1304 -3329 1304 -3329 0 1
rlabel polysilicon 1304 -3335 1304 -3335 0 3
rlabel polysilicon 1311 -3329 1311 -3329 0 1
rlabel polysilicon 1311 -3335 1311 -3335 0 3
rlabel polysilicon 1318 -3329 1318 -3329 0 1
rlabel polysilicon 1318 -3335 1318 -3335 0 3
rlabel polysilicon 1325 -3329 1325 -3329 0 1
rlabel polysilicon 1325 -3335 1325 -3335 0 3
rlabel polysilicon 1332 -3329 1332 -3329 0 1
rlabel polysilicon 1332 -3335 1332 -3335 0 3
rlabel polysilicon 1339 -3329 1339 -3329 0 1
rlabel polysilicon 1339 -3335 1339 -3335 0 3
rlabel polysilicon 1346 -3329 1346 -3329 0 1
rlabel polysilicon 1346 -3335 1346 -3335 0 3
rlabel polysilicon 1353 -3329 1353 -3329 0 1
rlabel polysilicon 1353 -3335 1353 -3335 0 3
rlabel polysilicon 1360 -3329 1360 -3329 0 1
rlabel polysilicon 1360 -3335 1360 -3335 0 3
rlabel polysilicon 1367 -3329 1367 -3329 0 1
rlabel polysilicon 1370 -3335 1370 -3335 0 4
rlabel polysilicon 1374 -3329 1374 -3329 0 1
rlabel polysilicon 1374 -3335 1374 -3335 0 3
rlabel polysilicon 1381 -3335 1381 -3335 0 3
rlabel polysilicon 1384 -3335 1384 -3335 0 4
rlabel polysilicon 1388 -3329 1388 -3329 0 1
rlabel polysilicon 1388 -3335 1388 -3335 0 3
rlabel polysilicon 1395 -3329 1395 -3329 0 1
rlabel polysilicon 1395 -3335 1395 -3335 0 3
rlabel polysilicon 1402 -3329 1402 -3329 0 1
rlabel polysilicon 1402 -3335 1402 -3335 0 3
rlabel polysilicon 1409 -3329 1409 -3329 0 1
rlabel polysilicon 1409 -3335 1409 -3335 0 3
rlabel polysilicon 1416 -3335 1416 -3335 0 3
rlabel polysilicon 1419 -3335 1419 -3335 0 4
rlabel polysilicon 1423 -3329 1423 -3329 0 1
rlabel polysilicon 1423 -3335 1423 -3335 0 3
rlabel polysilicon 1430 -3329 1430 -3329 0 1
rlabel polysilicon 1430 -3335 1430 -3335 0 3
rlabel polysilicon 1437 -3329 1437 -3329 0 1
rlabel polysilicon 1437 -3335 1437 -3335 0 3
rlabel polysilicon 1444 -3329 1444 -3329 0 1
rlabel polysilicon 1444 -3335 1444 -3335 0 3
rlabel polysilicon 1451 -3329 1451 -3329 0 1
rlabel polysilicon 1451 -3335 1451 -3335 0 3
rlabel polysilicon 1458 -3329 1458 -3329 0 1
rlabel polysilicon 1458 -3335 1458 -3335 0 3
rlabel polysilicon 1465 -3329 1465 -3329 0 1
rlabel polysilicon 1465 -3335 1465 -3335 0 3
rlabel polysilicon 1472 -3329 1472 -3329 0 1
rlabel polysilicon 1472 -3335 1472 -3335 0 3
rlabel polysilicon 1479 -3329 1479 -3329 0 1
rlabel polysilicon 1479 -3335 1479 -3335 0 3
rlabel polysilicon 1486 -3329 1486 -3329 0 1
rlabel polysilicon 1486 -3335 1486 -3335 0 3
rlabel polysilicon 1493 -3329 1493 -3329 0 1
rlabel polysilicon 1493 -3335 1493 -3335 0 3
rlabel polysilicon 1500 -3329 1500 -3329 0 1
rlabel polysilicon 1500 -3335 1500 -3335 0 3
rlabel polysilicon 1507 -3329 1507 -3329 0 1
rlabel polysilicon 1507 -3335 1507 -3335 0 3
rlabel polysilicon 1514 -3329 1514 -3329 0 1
rlabel polysilicon 1514 -3335 1514 -3335 0 3
rlabel polysilicon 1521 -3329 1521 -3329 0 1
rlabel polysilicon 1521 -3335 1521 -3335 0 3
rlabel polysilicon 1528 -3329 1528 -3329 0 1
rlabel polysilicon 1528 -3335 1528 -3335 0 3
rlabel polysilicon 1556 -3329 1556 -3329 0 1
rlabel polysilicon 1556 -3335 1556 -3335 0 3
rlabel polysilicon 1563 -3329 1563 -3329 0 1
rlabel polysilicon 1563 -3335 1563 -3335 0 3
rlabel polysilicon 1591 -3329 1591 -3329 0 1
rlabel polysilicon 1591 -3335 1591 -3335 0 3
rlabel polysilicon 1598 -3329 1598 -3329 0 1
rlabel polysilicon 1598 -3335 1598 -3335 0 3
rlabel polysilicon 1605 -3329 1605 -3329 0 1
rlabel polysilicon 1605 -3335 1605 -3335 0 3
rlabel polysilicon 1608 -3335 1608 -3335 0 4
rlabel polysilicon 1626 -3329 1626 -3329 0 1
rlabel polysilicon 1626 -3335 1626 -3335 0 3
rlabel polysilicon 1654 -3329 1654 -3329 0 1
rlabel polysilicon 1654 -3335 1654 -3335 0 3
rlabel polysilicon 1661 -3329 1661 -3329 0 1
rlabel polysilicon 1661 -3335 1661 -3335 0 3
rlabel polysilicon 1668 -3329 1668 -3329 0 1
rlabel polysilicon 1668 -3335 1668 -3335 0 3
rlabel polysilicon 1717 -3329 1717 -3329 0 1
rlabel polysilicon 1717 -3335 1717 -3335 0 3
rlabel polysilicon 1724 -3329 1724 -3329 0 1
rlabel polysilicon 1727 -3329 1727 -3329 0 2
rlabel polysilicon 1727 -3335 1727 -3335 0 4
rlabel polysilicon 1731 -3329 1731 -3329 0 1
rlabel polysilicon 1731 -3335 1731 -3335 0 3
rlabel polysilicon 1738 -3329 1738 -3329 0 1
rlabel polysilicon 1738 -3335 1738 -3335 0 3
rlabel polysilicon 1745 -3329 1745 -3329 0 1
rlabel polysilicon 1745 -3335 1745 -3335 0 3
rlabel polysilicon 1752 -3329 1752 -3329 0 1
rlabel polysilicon 1752 -3335 1752 -3335 0 3
rlabel polysilicon 1766 -3329 1766 -3329 0 1
rlabel polysilicon 1766 -3335 1766 -3335 0 3
rlabel polysilicon 1780 -3329 1780 -3329 0 1
rlabel polysilicon 1780 -3335 1780 -3335 0 3
rlabel polysilicon 1787 -3329 1787 -3329 0 1
rlabel polysilicon 1787 -3335 1787 -3335 0 3
rlabel polysilicon 1794 -3329 1794 -3329 0 1
rlabel polysilicon 1794 -3335 1794 -3335 0 3
rlabel polysilicon 1801 -3329 1801 -3329 0 1
rlabel polysilicon 1801 -3335 1801 -3335 0 3
rlabel polysilicon 1815 -3329 1815 -3329 0 1
rlabel polysilicon 1815 -3335 1815 -3335 0 3
rlabel polysilicon 1836 -3329 1836 -3329 0 1
rlabel polysilicon 1836 -3335 1836 -3335 0 3
rlabel polysilicon 1843 -3329 1843 -3329 0 1
rlabel polysilicon 1843 -3335 1843 -3335 0 3
rlabel polysilicon 1850 -3329 1850 -3329 0 1
rlabel polysilicon 1853 -3329 1853 -3329 0 2
rlabel polysilicon 1850 -3335 1850 -3335 0 3
rlabel polysilicon 1853 -3335 1853 -3335 0 4
rlabel polysilicon 1857 -3329 1857 -3329 0 1
rlabel polysilicon 1857 -3335 1857 -3335 0 3
rlabel polysilicon 1864 -3329 1864 -3329 0 1
rlabel polysilicon 1864 -3335 1864 -3335 0 3
rlabel polysilicon 1871 -3329 1871 -3329 0 1
rlabel polysilicon 1871 -3335 1871 -3335 0 3
rlabel polysilicon 1878 -3329 1878 -3329 0 1
rlabel polysilicon 1878 -3335 1878 -3335 0 3
rlabel polysilicon 1885 -3335 1885 -3335 0 3
rlabel polysilicon 1888 -3335 1888 -3335 0 4
rlabel polysilicon 1892 -3329 1892 -3329 0 1
rlabel polysilicon 1892 -3335 1892 -3335 0 3
rlabel polysilicon 1906 -3329 1906 -3329 0 1
rlabel polysilicon 1906 -3335 1906 -3335 0 3
rlabel polysilicon 1962 -3329 1962 -3329 0 1
rlabel polysilicon 1962 -3335 1962 -3335 0 3
rlabel polysilicon 1969 -3329 1969 -3329 0 1
rlabel polysilicon 1969 -3335 1969 -3335 0 3
rlabel polysilicon 2025 -3329 2025 -3329 0 1
rlabel polysilicon 2025 -3335 2025 -3335 0 3
rlabel polysilicon 2028 -3335 2028 -3335 0 4
rlabel polysilicon 2032 -3329 2032 -3329 0 1
rlabel polysilicon 2032 -3335 2032 -3335 0 3
rlabel polysilicon 173 -3416 173 -3416 0 2
rlabel polysilicon 170 -3422 170 -3422 0 3
rlabel polysilicon 173 -3422 173 -3422 0 4
rlabel polysilicon 180 -3416 180 -3416 0 2
rlabel polysilicon 296 -3416 296 -3416 0 1
rlabel polysilicon 296 -3422 296 -3422 0 3
rlabel polysilicon 310 -3416 310 -3416 0 1
rlabel polysilicon 310 -3422 310 -3422 0 3
rlabel polysilicon 317 -3422 317 -3422 0 3
rlabel polysilicon 331 -3416 331 -3416 0 1
rlabel polysilicon 331 -3422 331 -3422 0 3
rlabel polysilicon 338 -3416 338 -3416 0 1
rlabel polysilicon 338 -3422 338 -3422 0 3
rlabel polysilicon 345 -3416 345 -3416 0 1
rlabel polysilicon 345 -3422 345 -3422 0 3
rlabel polysilicon 359 -3416 359 -3416 0 1
rlabel polysilicon 359 -3422 359 -3422 0 3
rlabel polysilicon 373 -3416 373 -3416 0 1
rlabel polysilicon 373 -3422 373 -3422 0 3
rlabel polysilicon 380 -3416 380 -3416 0 1
rlabel polysilicon 380 -3422 380 -3422 0 3
rlabel polysilicon 387 -3416 387 -3416 0 1
rlabel polysilicon 390 -3416 390 -3416 0 2
rlabel polysilicon 390 -3422 390 -3422 0 4
rlabel polysilicon 394 -3416 394 -3416 0 1
rlabel polysilicon 394 -3422 394 -3422 0 3
rlabel polysilicon 401 -3416 401 -3416 0 1
rlabel polysilicon 401 -3422 401 -3422 0 3
rlabel polysilicon 404 -3422 404 -3422 0 4
rlabel polysilicon 408 -3416 408 -3416 0 1
rlabel polysilicon 408 -3422 408 -3422 0 3
rlabel polysilicon 422 -3416 422 -3416 0 1
rlabel polysilicon 422 -3422 422 -3422 0 3
rlabel polysilicon 429 -3416 429 -3416 0 1
rlabel polysilicon 429 -3422 429 -3422 0 3
rlabel polysilicon 436 -3416 436 -3416 0 1
rlabel polysilicon 436 -3422 436 -3422 0 3
rlabel polysilicon 439 -3422 439 -3422 0 4
rlabel polysilicon 443 -3416 443 -3416 0 1
rlabel polysilicon 443 -3422 443 -3422 0 3
rlabel polysilicon 450 -3416 450 -3416 0 1
rlabel polysilicon 450 -3422 450 -3422 0 3
rlabel polysilicon 457 -3416 457 -3416 0 1
rlabel polysilicon 457 -3422 457 -3422 0 3
rlabel polysilicon 464 -3416 464 -3416 0 1
rlabel polysilicon 464 -3422 464 -3422 0 3
rlabel polysilicon 474 -3416 474 -3416 0 2
rlabel polysilicon 471 -3422 471 -3422 0 3
rlabel polysilicon 474 -3422 474 -3422 0 4
rlabel polysilicon 478 -3416 478 -3416 0 1
rlabel polysilicon 478 -3422 478 -3422 0 3
rlabel polysilicon 488 -3416 488 -3416 0 2
rlabel polysilicon 488 -3422 488 -3422 0 4
rlabel polysilicon 492 -3416 492 -3416 0 1
rlabel polysilicon 492 -3422 492 -3422 0 3
rlabel polysilicon 499 -3416 499 -3416 0 1
rlabel polysilicon 499 -3422 499 -3422 0 3
rlabel polysilicon 506 -3416 506 -3416 0 1
rlabel polysilicon 506 -3422 506 -3422 0 3
rlabel polysilicon 513 -3416 513 -3416 0 1
rlabel polysilicon 513 -3422 513 -3422 0 3
rlabel polysilicon 520 -3416 520 -3416 0 1
rlabel polysilicon 520 -3422 520 -3422 0 3
rlabel polysilicon 527 -3416 527 -3416 0 1
rlabel polysilicon 527 -3422 527 -3422 0 3
rlabel polysilicon 534 -3416 534 -3416 0 1
rlabel polysilicon 534 -3422 534 -3422 0 3
rlabel polysilicon 541 -3416 541 -3416 0 1
rlabel polysilicon 541 -3422 541 -3422 0 3
rlabel polysilicon 548 -3416 548 -3416 0 1
rlabel polysilicon 548 -3422 548 -3422 0 3
rlabel polysilicon 555 -3416 555 -3416 0 1
rlabel polysilicon 555 -3422 555 -3422 0 3
rlabel polysilicon 558 -3422 558 -3422 0 4
rlabel polysilicon 562 -3416 562 -3416 0 1
rlabel polysilicon 562 -3422 562 -3422 0 3
rlabel polysilicon 569 -3416 569 -3416 0 1
rlabel polysilicon 569 -3422 569 -3422 0 3
rlabel polysilicon 576 -3422 576 -3422 0 3
rlabel polysilicon 583 -3416 583 -3416 0 1
rlabel polysilicon 583 -3422 583 -3422 0 3
rlabel polysilicon 590 -3416 590 -3416 0 1
rlabel polysilicon 590 -3422 590 -3422 0 3
rlabel polysilicon 597 -3416 597 -3416 0 1
rlabel polysilicon 597 -3422 597 -3422 0 3
rlabel polysilicon 604 -3416 604 -3416 0 1
rlabel polysilicon 604 -3422 604 -3422 0 3
rlabel polysilicon 611 -3416 611 -3416 0 1
rlabel polysilicon 611 -3422 611 -3422 0 3
rlabel polysilicon 618 -3416 618 -3416 0 1
rlabel polysilicon 618 -3422 618 -3422 0 3
rlabel polysilicon 625 -3416 625 -3416 0 1
rlabel polysilicon 625 -3422 625 -3422 0 3
rlabel polysilicon 632 -3416 632 -3416 0 1
rlabel polysilicon 632 -3422 632 -3422 0 3
rlabel polysilicon 639 -3416 639 -3416 0 1
rlabel polysilicon 639 -3422 639 -3422 0 3
rlabel polysilicon 646 -3416 646 -3416 0 1
rlabel polysilicon 646 -3422 646 -3422 0 3
rlabel polysilicon 653 -3416 653 -3416 0 1
rlabel polysilicon 653 -3422 653 -3422 0 3
rlabel polysilicon 660 -3416 660 -3416 0 1
rlabel polysilicon 660 -3422 660 -3422 0 3
rlabel polysilicon 667 -3416 667 -3416 0 1
rlabel polysilicon 674 -3416 674 -3416 0 1
rlabel polysilicon 674 -3422 674 -3422 0 3
rlabel polysilicon 681 -3416 681 -3416 0 1
rlabel polysilicon 681 -3422 681 -3422 0 3
rlabel polysilicon 688 -3416 688 -3416 0 1
rlabel polysilicon 695 -3416 695 -3416 0 1
rlabel polysilicon 695 -3422 695 -3422 0 3
rlabel polysilicon 702 -3416 702 -3416 0 1
rlabel polysilicon 702 -3422 702 -3422 0 3
rlabel polysilicon 709 -3416 709 -3416 0 1
rlabel polysilicon 709 -3422 709 -3422 0 3
rlabel polysilicon 716 -3416 716 -3416 0 1
rlabel polysilicon 716 -3422 716 -3422 0 3
rlabel polysilicon 723 -3416 723 -3416 0 1
rlabel polysilicon 726 -3416 726 -3416 0 2
rlabel polysilicon 723 -3422 723 -3422 0 3
rlabel polysilicon 726 -3422 726 -3422 0 4
rlabel polysilicon 730 -3416 730 -3416 0 1
rlabel polysilicon 730 -3422 730 -3422 0 3
rlabel polysilicon 737 -3416 737 -3416 0 1
rlabel polysilicon 737 -3422 737 -3422 0 3
rlabel polysilicon 744 -3416 744 -3416 0 1
rlabel polysilicon 744 -3422 744 -3422 0 3
rlabel polysilicon 751 -3416 751 -3416 0 1
rlabel polysilicon 751 -3422 751 -3422 0 3
rlabel polysilicon 758 -3416 758 -3416 0 1
rlabel polysilicon 758 -3422 758 -3422 0 3
rlabel polysilicon 765 -3416 765 -3416 0 1
rlabel polysilicon 765 -3422 765 -3422 0 3
rlabel polysilicon 772 -3416 772 -3416 0 1
rlabel polysilicon 772 -3422 772 -3422 0 3
rlabel polysilicon 779 -3416 779 -3416 0 1
rlabel polysilicon 779 -3422 779 -3422 0 3
rlabel polysilicon 786 -3416 786 -3416 0 1
rlabel polysilicon 786 -3422 786 -3422 0 3
rlabel polysilicon 793 -3416 793 -3416 0 1
rlabel polysilicon 793 -3422 793 -3422 0 3
rlabel polysilicon 800 -3416 800 -3416 0 1
rlabel polysilicon 803 -3416 803 -3416 0 2
rlabel polysilicon 807 -3416 807 -3416 0 1
rlabel polysilicon 807 -3422 807 -3422 0 3
rlabel polysilicon 814 -3416 814 -3416 0 1
rlabel polysilicon 814 -3422 814 -3422 0 3
rlabel polysilicon 821 -3416 821 -3416 0 1
rlabel polysilicon 821 -3422 821 -3422 0 3
rlabel polysilicon 828 -3416 828 -3416 0 1
rlabel polysilicon 828 -3422 828 -3422 0 3
rlabel polysilicon 835 -3416 835 -3416 0 1
rlabel polysilicon 835 -3422 835 -3422 0 3
rlabel polysilicon 842 -3416 842 -3416 0 1
rlabel polysilicon 842 -3422 842 -3422 0 3
rlabel polysilicon 845 -3422 845 -3422 0 4
rlabel polysilicon 849 -3416 849 -3416 0 1
rlabel polysilicon 849 -3422 849 -3422 0 3
rlabel polysilicon 859 -3416 859 -3416 0 2
rlabel polysilicon 859 -3422 859 -3422 0 4
rlabel polysilicon 863 -3416 863 -3416 0 1
rlabel polysilicon 863 -3422 863 -3422 0 3
rlabel polysilicon 870 -3416 870 -3416 0 1
rlabel polysilicon 870 -3422 870 -3422 0 3
rlabel polysilicon 877 -3416 877 -3416 0 1
rlabel polysilicon 877 -3422 877 -3422 0 3
rlabel polysilicon 884 -3416 884 -3416 0 1
rlabel polysilicon 884 -3422 884 -3422 0 3
rlabel polysilicon 891 -3416 891 -3416 0 1
rlabel polysilicon 891 -3422 891 -3422 0 3
rlabel polysilicon 901 -3416 901 -3416 0 2
rlabel polysilicon 898 -3422 898 -3422 0 3
rlabel polysilicon 901 -3422 901 -3422 0 4
rlabel polysilicon 905 -3416 905 -3416 0 1
rlabel polysilicon 905 -3422 905 -3422 0 3
rlabel polysilicon 912 -3416 912 -3416 0 1
rlabel polysilicon 912 -3422 912 -3422 0 3
rlabel polysilicon 919 -3416 919 -3416 0 1
rlabel polysilicon 919 -3422 919 -3422 0 3
rlabel polysilicon 922 -3422 922 -3422 0 4
rlabel polysilicon 926 -3416 926 -3416 0 1
rlabel polysilicon 926 -3422 926 -3422 0 3
rlabel polysilicon 933 -3416 933 -3416 0 1
rlabel polysilicon 936 -3416 936 -3416 0 2
rlabel polysilicon 940 -3416 940 -3416 0 1
rlabel polysilicon 940 -3422 940 -3422 0 3
rlabel polysilicon 947 -3416 947 -3416 0 1
rlabel polysilicon 947 -3422 947 -3422 0 3
rlabel polysilicon 954 -3416 954 -3416 0 1
rlabel polysilicon 954 -3422 954 -3422 0 3
rlabel polysilicon 961 -3416 961 -3416 0 1
rlabel polysilicon 961 -3422 961 -3422 0 3
rlabel polysilicon 968 -3416 968 -3416 0 1
rlabel polysilicon 968 -3422 968 -3422 0 3
rlabel polysilicon 975 -3416 975 -3416 0 1
rlabel polysilicon 975 -3422 975 -3422 0 3
rlabel polysilicon 982 -3416 982 -3416 0 1
rlabel polysilicon 982 -3422 982 -3422 0 3
rlabel polysilicon 989 -3416 989 -3416 0 1
rlabel polysilicon 992 -3416 992 -3416 0 2
rlabel polysilicon 989 -3422 989 -3422 0 3
rlabel polysilicon 992 -3422 992 -3422 0 4
rlabel polysilicon 996 -3416 996 -3416 0 1
rlabel polysilicon 996 -3422 996 -3422 0 3
rlabel polysilicon 1003 -3416 1003 -3416 0 1
rlabel polysilicon 1003 -3422 1003 -3422 0 3
rlabel polysilicon 1010 -3416 1010 -3416 0 1
rlabel polysilicon 1010 -3422 1010 -3422 0 3
rlabel polysilicon 1017 -3416 1017 -3416 0 1
rlabel polysilicon 1017 -3422 1017 -3422 0 3
rlabel polysilicon 1024 -3416 1024 -3416 0 1
rlabel polysilicon 1027 -3416 1027 -3416 0 2
rlabel polysilicon 1031 -3416 1031 -3416 0 1
rlabel polysilicon 1034 -3416 1034 -3416 0 2
rlabel polysilicon 1031 -3422 1031 -3422 0 3
rlabel polysilicon 1034 -3422 1034 -3422 0 4
rlabel polysilicon 1038 -3416 1038 -3416 0 1
rlabel polysilicon 1038 -3422 1038 -3422 0 3
rlabel polysilicon 1045 -3416 1045 -3416 0 1
rlabel polysilicon 1045 -3422 1045 -3422 0 3
rlabel polysilicon 1052 -3416 1052 -3416 0 1
rlabel polysilicon 1052 -3422 1052 -3422 0 3
rlabel polysilicon 1059 -3416 1059 -3416 0 1
rlabel polysilicon 1059 -3422 1059 -3422 0 3
rlabel polysilicon 1066 -3416 1066 -3416 0 1
rlabel polysilicon 1066 -3422 1066 -3422 0 3
rlabel polysilicon 1069 -3422 1069 -3422 0 4
rlabel polysilicon 1073 -3416 1073 -3416 0 1
rlabel polysilicon 1073 -3422 1073 -3422 0 3
rlabel polysilicon 1080 -3416 1080 -3416 0 1
rlabel polysilicon 1080 -3422 1080 -3422 0 3
rlabel polysilicon 1087 -3416 1087 -3416 0 1
rlabel polysilicon 1087 -3422 1087 -3422 0 3
rlabel polysilicon 1094 -3416 1094 -3416 0 1
rlabel polysilicon 1094 -3422 1094 -3422 0 3
rlabel polysilicon 1101 -3416 1101 -3416 0 1
rlabel polysilicon 1101 -3422 1101 -3422 0 3
rlabel polysilicon 1108 -3416 1108 -3416 0 1
rlabel polysilicon 1108 -3422 1108 -3422 0 3
rlabel polysilicon 1115 -3416 1115 -3416 0 1
rlabel polysilicon 1115 -3422 1115 -3422 0 3
rlabel polysilicon 1122 -3416 1122 -3416 0 1
rlabel polysilicon 1125 -3416 1125 -3416 0 2
rlabel polysilicon 1122 -3422 1122 -3422 0 3
rlabel polysilicon 1125 -3422 1125 -3422 0 4
rlabel polysilicon 1136 -3416 1136 -3416 0 1
rlabel polysilicon 1136 -3422 1136 -3422 0 3
rlabel polysilicon 1143 -3416 1143 -3416 0 1
rlabel polysilicon 1143 -3422 1143 -3422 0 3
rlabel polysilicon 1160 -3416 1160 -3416 0 2
rlabel polysilicon 1157 -3422 1157 -3422 0 3
rlabel polysilicon 1171 -3416 1171 -3416 0 1
rlabel polysilicon 1171 -3422 1171 -3422 0 3
rlabel polysilicon 1178 -3416 1178 -3416 0 1
rlabel polysilicon 1178 -3422 1178 -3422 0 3
rlabel polysilicon 1185 -3416 1185 -3416 0 1
rlabel polysilicon 1185 -3422 1185 -3422 0 3
rlabel polysilicon 1192 -3416 1192 -3416 0 1
rlabel polysilicon 1192 -3422 1192 -3422 0 3
rlabel polysilicon 1199 -3416 1199 -3416 0 1
rlabel polysilicon 1199 -3422 1199 -3422 0 3
rlabel polysilicon 1206 -3416 1206 -3416 0 1
rlabel polysilicon 1209 -3416 1209 -3416 0 2
rlabel polysilicon 1206 -3422 1206 -3422 0 3
rlabel polysilicon 1213 -3416 1213 -3416 0 1
rlabel polysilicon 1213 -3422 1213 -3422 0 3
rlabel polysilicon 1220 -3416 1220 -3416 0 1
rlabel polysilicon 1220 -3422 1220 -3422 0 3
rlabel polysilicon 1227 -3416 1227 -3416 0 1
rlabel polysilicon 1227 -3422 1227 -3422 0 3
rlabel polysilicon 1234 -3416 1234 -3416 0 1
rlabel polysilicon 1234 -3422 1234 -3422 0 3
rlabel polysilicon 1241 -3416 1241 -3416 0 1
rlabel polysilicon 1241 -3422 1241 -3422 0 3
rlabel polysilicon 1248 -3416 1248 -3416 0 1
rlabel polysilicon 1248 -3422 1248 -3422 0 3
rlabel polysilicon 1255 -3416 1255 -3416 0 1
rlabel polysilicon 1255 -3422 1255 -3422 0 3
rlabel polysilicon 1262 -3416 1262 -3416 0 1
rlabel polysilicon 1262 -3422 1262 -3422 0 3
rlabel polysilicon 1269 -3416 1269 -3416 0 1
rlabel polysilicon 1269 -3422 1269 -3422 0 3
rlabel polysilicon 1276 -3422 1276 -3422 0 3
rlabel polysilicon 1283 -3416 1283 -3416 0 1
rlabel polysilicon 1283 -3422 1283 -3422 0 3
rlabel polysilicon 1290 -3416 1290 -3416 0 1
rlabel polysilicon 1290 -3422 1290 -3422 0 3
rlabel polysilicon 1297 -3416 1297 -3416 0 1
rlabel polysilicon 1297 -3422 1297 -3422 0 3
rlabel polysilicon 1304 -3416 1304 -3416 0 1
rlabel polysilicon 1307 -3422 1307 -3422 0 4
rlabel polysilicon 1332 -3416 1332 -3416 0 1
rlabel polysilicon 1332 -3422 1332 -3422 0 3
rlabel polysilicon 1346 -3416 1346 -3416 0 1
rlabel polysilicon 1346 -3422 1346 -3422 0 3
rlabel polysilicon 1360 -3416 1360 -3416 0 1
rlabel polysilicon 1360 -3422 1360 -3422 0 3
rlabel polysilicon 1367 -3416 1367 -3416 0 1
rlabel polysilicon 1367 -3422 1367 -3422 0 3
rlabel polysilicon 1374 -3416 1374 -3416 0 1
rlabel polysilicon 1377 -3416 1377 -3416 0 2
rlabel polysilicon 1374 -3422 1374 -3422 0 3
rlabel polysilicon 1381 -3416 1381 -3416 0 1
rlabel polysilicon 1381 -3422 1381 -3422 0 3
rlabel polysilicon 1451 -3416 1451 -3416 0 1
rlabel polysilicon 1451 -3422 1451 -3422 0 3
rlabel polysilicon 1458 -3416 1458 -3416 0 1
rlabel polysilicon 1458 -3422 1458 -3422 0 3
rlabel polysilicon 1465 -3416 1465 -3416 0 1
rlabel polysilicon 1465 -3422 1465 -3422 0 3
rlabel polysilicon 1472 -3416 1472 -3416 0 1
rlabel polysilicon 1472 -3422 1472 -3422 0 3
rlabel polysilicon 1500 -3416 1500 -3416 0 1
rlabel polysilicon 1500 -3422 1500 -3422 0 3
rlabel polysilicon 1521 -3416 1521 -3416 0 1
rlabel polysilicon 1521 -3422 1521 -3422 0 3
rlabel polysilicon 1528 -3416 1528 -3416 0 1
rlabel polysilicon 1528 -3422 1528 -3422 0 3
rlabel polysilicon 1549 -3416 1549 -3416 0 1
rlabel polysilicon 1552 -3416 1552 -3416 0 2
rlabel polysilicon 1584 -3416 1584 -3416 0 1
rlabel polysilicon 1587 -3416 1587 -3416 0 2
rlabel polysilicon 1584 -3422 1584 -3422 0 3
rlabel polysilicon 1612 -3416 1612 -3416 0 1
rlabel polysilicon 1612 -3422 1612 -3422 0 3
rlabel polysilicon 1647 -3416 1647 -3416 0 1
rlabel polysilicon 1647 -3422 1647 -3422 0 3
rlabel polysilicon 1654 -3416 1654 -3416 0 1
rlabel polysilicon 1654 -3422 1654 -3422 0 3
rlabel polysilicon 1724 -3416 1724 -3416 0 1
rlabel polysilicon 1724 -3422 1724 -3422 0 3
rlabel polysilicon 1731 -3416 1731 -3416 0 1
rlabel polysilicon 1731 -3422 1731 -3422 0 3
rlabel polysilicon 1738 -3416 1738 -3416 0 1
rlabel polysilicon 1738 -3422 1738 -3422 0 3
rlabel polysilicon 1759 -3416 1759 -3416 0 1
rlabel polysilicon 1759 -3422 1759 -3422 0 3
rlabel polysilicon 1769 -3416 1769 -3416 0 2
rlabel polysilicon 1766 -3422 1766 -3422 0 3
rlabel polysilicon 1780 -3416 1780 -3416 0 1
rlabel polysilicon 1780 -3422 1780 -3422 0 3
rlabel polysilicon 1787 -3416 1787 -3416 0 1
rlabel polysilicon 1787 -3422 1787 -3422 0 3
rlabel polysilicon 1801 -3416 1801 -3416 0 1
rlabel polysilicon 1801 -3422 1801 -3422 0 3
rlabel polysilicon 1808 -3416 1808 -3416 0 1
rlabel polysilicon 1811 -3416 1811 -3416 0 2
rlabel polysilicon 1808 -3422 1808 -3422 0 3
rlabel polysilicon 1822 -3416 1822 -3416 0 1
rlabel polysilicon 1822 -3422 1822 -3422 0 3
rlabel polysilicon 1829 -3416 1829 -3416 0 1
rlabel polysilicon 1829 -3422 1829 -3422 0 3
rlabel polysilicon 1836 -3416 1836 -3416 0 1
rlabel polysilicon 1836 -3422 1836 -3422 0 3
rlabel polysilicon 1843 -3416 1843 -3416 0 1
rlabel polysilicon 1843 -3422 1843 -3422 0 3
rlabel polysilicon 1850 -3416 1850 -3416 0 1
rlabel polysilicon 1850 -3422 1850 -3422 0 3
rlabel polysilicon 1857 -3416 1857 -3416 0 1
rlabel polysilicon 1857 -3422 1857 -3422 0 3
rlabel polysilicon 1864 -3416 1864 -3416 0 1
rlabel polysilicon 1864 -3422 1864 -3422 0 3
rlabel polysilicon 1867 -3422 1867 -3422 0 4
rlabel polysilicon 1871 -3416 1871 -3416 0 1
rlabel polysilicon 1871 -3422 1871 -3422 0 3
rlabel polysilicon 1955 -3416 1955 -3416 0 1
rlabel polysilicon 1955 -3422 1955 -3422 0 3
rlabel polysilicon 1962 -3416 1962 -3416 0 1
rlabel polysilicon 1962 -3422 1962 -3422 0 3
rlabel polysilicon 2025 -3416 2025 -3416 0 1
rlabel polysilicon 2028 -3416 2028 -3416 0 2
rlabel polysilicon 2025 -3422 2025 -3422 0 3
rlabel polysilicon 2032 -3416 2032 -3416 0 1
rlabel polysilicon 2032 -3422 2032 -3422 0 3
rlabel polysilicon 173 -3461 173 -3461 0 2
rlabel polysilicon 268 -3461 268 -3461 0 1
rlabel polysilicon 271 -3467 271 -3467 0 4
rlabel polysilicon 324 -3461 324 -3461 0 1
rlabel polysilicon 324 -3467 324 -3467 0 3
rlabel polysilicon 380 -3461 380 -3461 0 1
rlabel polysilicon 380 -3467 380 -3467 0 3
rlabel polysilicon 415 -3461 415 -3461 0 1
rlabel polysilicon 415 -3467 415 -3467 0 3
rlabel polysilicon 422 -3461 422 -3461 0 1
rlabel polysilicon 422 -3467 422 -3467 0 3
rlabel polysilicon 439 -3467 439 -3467 0 4
rlabel polysilicon 443 -3461 443 -3461 0 1
rlabel polysilicon 443 -3467 443 -3467 0 3
rlabel polysilicon 457 -3461 457 -3461 0 1
rlabel polysilicon 457 -3467 457 -3467 0 3
rlabel polysilicon 464 -3461 464 -3461 0 1
rlabel polysilicon 467 -3461 467 -3461 0 2
rlabel polysilicon 467 -3467 467 -3467 0 4
rlabel polysilicon 485 -3461 485 -3461 0 1
rlabel polysilicon 485 -3467 485 -3467 0 3
rlabel polysilicon 492 -3461 492 -3461 0 1
rlabel polysilicon 492 -3467 492 -3467 0 3
rlabel polysilicon 499 -3461 499 -3461 0 1
rlabel polysilicon 499 -3467 499 -3467 0 3
rlabel polysilicon 506 -3461 506 -3461 0 1
rlabel polysilicon 506 -3467 506 -3467 0 3
rlabel polysilicon 513 -3461 513 -3461 0 1
rlabel polysilicon 513 -3467 513 -3467 0 3
rlabel polysilicon 520 -3461 520 -3461 0 1
rlabel polysilicon 520 -3467 520 -3467 0 3
rlabel polysilicon 523 -3467 523 -3467 0 4
rlabel polysilicon 534 -3461 534 -3461 0 1
rlabel polysilicon 534 -3467 534 -3467 0 3
rlabel polysilicon 541 -3461 541 -3461 0 1
rlabel polysilicon 541 -3467 541 -3467 0 3
rlabel polysilicon 551 -3467 551 -3467 0 4
rlabel polysilicon 555 -3461 555 -3461 0 1
rlabel polysilicon 555 -3467 555 -3467 0 3
rlabel polysilicon 562 -3461 562 -3461 0 1
rlabel polysilicon 562 -3467 562 -3467 0 3
rlabel polysilicon 569 -3461 569 -3461 0 1
rlabel polysilicon 569 -3467 569 -3467 0 3
rlabel polysilicon 576 -3461 576 -3461 0 1
rlabel polysilicon 579 -3461 579 -3461 0 2
rlabel polysilicon 579 -3467 579 -3467 0 4
rlabel polysilicon 583 -3461 583 -3461 0 1
rlabel polysilicon 583 -3467 583 -3467 0 3
rlabel polysilicon 590 -3461 590 -3461 0 1
rlabel polysilicon 593 -3461 593 -3461 0 2
rlabel polysilicon 590 -3467 590 -3467 0 3
rlabel polysilicon 597 -3461 597 -3461 0 1
rlabel polysilicon 597 -3467 597 -3467 0 3
rlabel polysilicon 604 -3461 604 -3461 0 1
rlabel polysilicon 604 -3467 604 -3467 0 3
rlabel polysilicon 611 -3461 611 -3461 0 1
rlabel polysilicon 611 -3467 611 -3467 0 3
rlabel polysilicon 621 -3461 621 -3461 0 2
rlabel polysilicon 625 -3461 625 -3461 0 1
rlabel polysilicon 628 -3461 628 -3461 0 2
rlabel polysilicon 628 -3467 628 -3467 0 4
rlabel polysilicon 632 -3461 632 -3461 0 1
rlabel polysilicon 632 -3467 632 -3467 0 3
rlabel polysilicon 639 -3461 639 -3461 0 1
rlabel polysilicon 639 -3467 639 -3467 0 3
rlabel polysilicon 642 -3467 642 -3467 0 4
rlabel polysilicon 646 -3461 646 -3461 0 1
rlabel polysilicon 646 -3467 646 -3467 0 3
rlabel polysilicon 653 -3461 653 -3461 0 1
rlabel polysilicon 653 -3467 653 -3467 0 3
rlabel polysilicon 660 -3461 660 -3461 0 1
rlabel polysilicon 660 -3467 660 -3467 0 3
rlabel polysilicon 667 -3461 667 -3461 0 1
rlabel polysilicon 667 -3467 667 -3467 0 3
rlabel polysilicon 674 -3461 674 -3461 0 1
rlabel polysilicon 674 -3467 674 -3467 0 3
rlabel polysilicon 681 -3461 681 -3461 0 1
rlabel polysilicon 684 -3461 684 -3461 0 2
rlabel polysilicon 681 -3467 681 -3467 0 3
rlabel polysilicon 688 -3467 688 -3467 0 3
rlabel polysilicon 695 -3461 695 -3461 0 1
rlabel polysilicon 695 -3467 695 -3467 0 3
rlabel polysilicon 702 -3461 702 -3461 0 1
rlabel polysilicon 705 -3461 705 -3461 0 2
rlabel polysilicon 702 -3467 702 -3467 0 3
rlabel polysilicon 705 -3467 705 -3467 0 4
rlabel polysilicon 709 -3461 709 -3461 0 1
rlabel polysilicon 709 -3467 709 -3467 0 3
rlabel polysilicon 716 -3461 716 -3461 0 1
rlabel polysilicon 716 -3467 716 -3467 0 3
rlabel polysilicon 723 -3461 723 -3461 0 1
rlabel polysilicon 723 -3467 723 -3467 0 3
rlabel polysilicon 730 -3461 730 -3461 0 1
rlabel polysilicon 730 -3467 730 -3467 0 3
rlabel polysilicon 737 -3461 737 -3461 0 1
rlabel polysilicon 737 -3467 737 -3467 0 3
rlabel polysilicon 744 -3461 744 -3461 0 1
rlabel polysilicon 744 -3467 744 -3467 0 3
rlabel polysilicon 751 -3461 751 -3461 0 1
rlabel polysilicon 751 -3467 751 -3467 0 3
rlabel polysilicon 758 -3461 758 -3461 0 1
rlabel polysilicon 758 -3467 758 -3467 0 3
rlabel polysilicon 779 -3461 779 -3461 0 1
rlabel polysilicon 779 -3467 779 -3467 0 3
rlabel polysilicon 793 -3461 793 -3461 0 1
rlabel polysilicon 793 -3467 793 -3467 0 3
rlabel polysilicon 800 -3461 800 -3461 0 1
rlabel polysilicon 800 -3467 800 -3467 0 3
rlabel polysilicon 807 -3461 807 -3461 0 1
rlabel polysilicon 807 -3467 807 -3467 0 3
rlabel polysilicon 814 -3461 814 -3461 0 1
rlabel polysilicon 814 -3467 814 -3467 0 3
rlabel polysilicon 821 -3461 821 -3461 0 1
rlabel polysilicon 821 -3467 821 -3467 0 3
rlabel polysilicon 828 -3461 828 -3461 0 1
rlabel polysilicon 828 -3467 828 -3467 0 3
rlabel polysilicon 835 -3461 835 -3461 0 1
rlabel polysilicon 835 -3467 835 -3467 0 3
rlabel polysilicon 842 -3461 842 -3461 0 1
rlabel polysilicon 842 -3467 842 -3467 0 3
rlabel polysilicon 849 -3461 849 -3461 0 1
rlabel polysilicon 849 -3467 849 -3467 0 3
rlabel polysilicon 877 -3461 877 -3461 0 1
rlabel polysilicon 877 -3467 877 -3467 0 3
rlabel polysilicon 884 -3461 884 -3461 0 1
rlabel polysilicon 884 -3467 884 -3467 0 3
rlabel polysilicon 915 -3461 915 -3461 0 2
rlabel polysilicon 912 -3467 912 -3467 0 3
rlabel polysilicon 915 -3467 915 -3467 0 4
rlabel polysilicon 922 -3461 922 -3461 0 2
rlabel polysilicon 919 -3467 919 -3467 0 3
rlabel polysilicon 922 -3467 922 -3467 0 4
rlabel polysilicon 954 -3461 954 -3461 0 1
rlabel polysilicon 954 -3467 954 -3467 0 3
rlabel polysilicon 975 -3461 975 -3461 0 1
rlabel polysilicon 975 -3467 975 -3467 0 3
rlabel polysilicon 996 -3461 996 -3461 0 1
rlabel polysilicon 1003 -3461 1003 -3461 0 1
rlabel polysilicon 1003 -3467 1003 -3467 0 3
rlabel polysilicon 1010 -3461 1010 -3461 0 1
rlabel polysilicon 1010 -3467 1010 -3467 0 3
rlabel polysilicon 1017 -3461 1017 -3461 0 1
rlabel polysilicon 1017 -3467 1017 -3467 0 3
rlabel polysilicon 1024 -3461 1024 -3461 0 1
rlabel polysilicon 1024 -3467 1024 -3467 0 3
rlabel polysilicon 1031 -3461 1031 -3461 0 1
rlabel polysilicon 1031 -3467 1031 -3467 0 3
rlabel polysilicon 1038 -3461 1038 -3461 0 1
rlabel polysilicon 1038 -3467 1038 -3467 0 3
rlabel polysilicon 1045 -3461 1045 -3461 0 1
rlabel polysilicon 1045 -3467 1045 -3467 0 3
rlabel polysilicon 1052 -3461 1052 -3461 0 1
rlabel polysilicon 1052 -3467 1052 -3467 0 3
rlabel polysilicon 1059 -3461 1059 -3461 0 1
rlabel polysilicon 1059 -3467 1059 -3467 0 3
rlabel polysilicon 1062 -3467 1062 -3467 0 4
rlabel polysilicon 1066 -3461 1066 -3461 0 1
rlabel polysilicon 1066 -3467 1066 -3467 0 3
rlabel polysilicon 1073 -3461 1073 -3461 0 1
rlabel polysilicon 1073 -3467 1073 -3467 0 3
rlabel polysilicon 1080 -3461 1080 -3461 0 1
rlabel polysilicon 1083 -3461 1083 -3461 0 2
rlabel polysilicon 1083 -3467 1083 -3467 0 4
rlabel polysilicon 1087 -3461 1087 -3461 0 1
rlabel polysilicon 1087 -3467 1087 -3467 0 3
rlabel polysilicon 1094 -3461 1094 -3461 0 1
rlabel polysilicon 1094 -3467 1094 -3467 0 3
rlabel polysilicon 1101 -3461 1101 -3461 0 1
rlabel polysilicon 1101 -3467 1101 -3467 0 3
rlabel polysilicon 1108 -3461 1108 -3461 0 1
rlabel polysilicon 1108 -3467 1108 -3467 0 3
rlabel polysilicon 1125 -3461 1125 -3461 0 2
rlabel polysilicon 1122 -3467 1122 -3467 0 3
rlabel polysilicon 1125 -3467 1125 -3467 0 4
rlabel polysilicon 1129 -3461 1129 -3461 0 1
rlabel polysilicon 1129 -3467 1129 -3467 0 3
rlabel polysilicon 1157 -3461 1157 -3461 0 1
rlabel polysilicon 1157 -3467 1157 -3467 0 3
rlabel polysilicon 1164 -3461 1164 -3461 0 1
rlabel polysilicon 1164 -3467 1164 -3467 0 3
rlabel polysilicon 1171 -3461 1171 -3461 0 1
rlabel polysilicon 1171 -3467 1171 -3467 0 3
rlabel polysilicon 1178 -3461 1178 -3461 0 1
rlabel polysilicon 1181 -3461 1181 -3461 0 2
rlabel polysilicon 1178 -3467 1178 -3467 0 3
rlabel polysilicon 1185 -3461 1185 -3461 0 1
rlabel polysilicon 1185 -3467 1185 -3467 0 3
rlabel polysilicon 1192 -3461 1192 -3461 0 1
rlabel polysilicon 1192 -3467 1192 -3467 0 3
rlabel polysilicon 1199 -3461 1199 -3461 0 1
rlabel polysilicon 1199 -3467 1199 -3467 0 3
rlabel polysilicon 1206 -3461 1206 -3461 0 1
rlabel polysilicon 1206 -3467 1206 -3467 0 3
rlabel polysilicon 1213 -3461 1213 -3461 0 1
rlabel polysilicon 1213 -3467 1213 -3467 0 3
rlabel polysilicon 1220 -3461 1220 -3461 0 1
rlabel polysilicon 1220 -3467 1220 -3467 0 3
rlabel polysilicon 1227 -3461 1227 -3461 0 1
rlabel polysilicon 1227 -3467 1227 -3467 0 3
rlabel polysilicon 1234 -3461 1234 -3461 0 1
rlabel polysilicon 1234 -3467 1234 -3467 0 3
rlabel polysilicon 1241 -3461 1241 -3461 0 1
rlabel polysilicon 1241 -3467 1241 -3467 0 3
rlabel polysilicon 1248 -3461 1248 -3461 0 1
rlabel polysilicon 1248 -3467 1248 -3467 0 3
rlabel polysilicon 1286 -3461 1286 -3461 0 2
rlabel polysilicon 1283 -3467 1283 -3467 0 3
rlabel polysilicon 1290 -3461 1290 -3461 0 1
rlabel polysilicon 1290 -3467 1290 -3467 0 3
rlabel polysilicon 1304 -3461 1304 -3461 0 1
rlabel polysilicon 1307 -3461 1307 -3461 0 2
rlabel polysilicon 1304 -3467 1304 -3467 0 3
rlabel polysilicon 1307 -3467 1307 -3467 0 4
rlabel polysilicon 1311 -3461 1311 -3461 0 1
rlabel polysilicon 1311 -3467 1311 -3467 0 3
rlabel polysilicon 1318 -3461 1318 -3461 0 1
rlabel polysilicon 1321 -3461 1321 -3461 0 2
rlabel polysilicon 1318 -3467 1318 -3467 0 3
rlabel polysilicon 1325 -3461 1325 -3461 0 1
rlabel polysilicon 1325 -3467 1325 -3467 0 3
rlabel polysilicon 1332 -3461 1332 -3461 0 1
rlabel polysilicon 1332 -3467 1332 -3467 0 3
rlabel polysilicon 1360 -3461 1360 -3461 0 1
rlabel polysilicon 1360 -3467 1360 -3467 0 3
rlabel polysilicon 1437 -3461 1437 -3461 0 1
rlabel polysilicon 1437 -3467 1437 -3467 0 3
rlabel polysilicon 1444 -3461 1444 -3461 0 1
rlabel polysilicon 1444 -3467 1444 -3467 0 3
rlabel polysilicon 1451 -3461 1451 -3461 0 1
rlabel polysilicon 1451 -3467 1451 -3467 0 3
rlabel polysilicon 1458 -3461 1458 -3461 0 1
rlabel polysilicon 1461 -3461 1461 -3461 0 2
rlabel polysilicon 1458 -3467 1458 -3467 0 3
rlabel polysilicon 1465 -3461 1465 -3461 0 1
rlabel polysilicon 1465 -3467 1465 -3467 0 3
rlabel polysilicon 1493 -3461 1493 -3461 0 1
rlabel polysilicon 1493 -3467 1493 -3467 0 3
rlabel polysilicon 1500 -3461 1500 -3461 0 1
rlabel polysilicon 1500 -3467 1500 -3467 0 3
rlabel polysilicon 1514 -3461 1514 -3461 0 1
rlabel polysilicon 1514 -3467 1514 -3467 0 3
rlabel polysilicon 1521 -3461 1521 -3461 0 1
rlabel polysilicon 1521 -3467 1521 -3467 0 3
rlabel polysilicon 1626 -3461 1626 -3461 0 1
rlabel polysilicon 1629 -3461 1629 -3461 0 2
rlabel polysilicon 1640 -3461 1640 -3461 0 1
rlabel polysilicon 1640 -3467 1640 -3467 0 3
rlabel polysilicon 1724 -3461 1724 -3461 0 1
rlabel polysilicon 1724 -3467 1724 -3467 0 3
rlabel polysilicon 1731 -3461 1731 -3461 0 1
rlabel polysilicon 1731 -3467 1731 -3467 0 3
rlabel polysilicon 1748 -3461 1748 -3461 0 2
rlabel polysilicon 1745 -3467 1745 -3467 0 3
rlabel polysilicon 1766 -3461 1766 -3461 0 1
rlabel polysilicon 1766 -3467 1766 -3467 0 3
rlabel polysilicon 1780 -3461 1780 -3461 0 1
rlabel polysilicon 1780 -3467 1780 -3467 0 3
rlabel polysilicon 1794 -3461 1794 -3461 0 1
rlabel polysilicon 1794 -3467 1794 -3467 0 3
rlabel polysilicon 1822 -3461 1822 -3461 0 1
rlabel polysilicon 1822 -3467 1822 -3467 0 3
rlabel polysilicon 1829 -3461 1829 -3461 0 1
rlabel polysilicon 1829 -3467 1829 -3467 0 3
rlabel polysilicon 1836 -3467 1836 -3467 0 3
rlabel polysilicon 1839 -3467 1839 -3467 0 4
rlabel polysilicon 1843 -3461 1843 -3461 0 1
rlabel polysilicon 1843 -3467 1843 -3467 0 3
rlabel polysilicon 1850 -3461 1850 -3461 0 1
rlabel polysilicon 1850 -3467 1850 -3467 0 3
rlabel polysilicon 1857 -3461 1857 -3461 0 1
rlabel polysilicon 1860 -3461 1860 -3461 0 2
rlabel polysilicon 1860 -3467 1860 -3467 0 4
rlabel polysilicon 1864 -3461 1864 -3461 0 1
rlabel polysilicon 1867 -3461 1867 -3461 0 2
rlabel polysilicon 1864 -3467 1864 -3467 0 3
rlabel polysilicon 1871 -3461 1871 -3461 0 1
rlabel polysilicon 1871 -3467 1871 -3467 0 3
rlabel polysilicon 1955 -3461 1955 -3461 0 1
rlabel polysilicon 1955 -3467 1955 -3467 0 3
rlabel polysilicon 1962 -3461 1962 -3461 0 1
rlabel polysilicon 1962 -3467 1962 -3467 0 3
rlabel polysilicon 2025 -3461 2025 -3461 0 1
rlabel polysilicon 2025 -3467 2025 -3467 0 3
rlabel polysilicon 2028 -3467 2028 -3467 0 4
rlabel polysilicon 2032 -3461 2032 -3461 0 1
rlabel polysilicon 2032 -3467 2032 -3467 0 3
rlabel polysilicon 331 -3490 331 -3490 0 1
rlabel polysilicon 331 -3496 331 -3496 0 3
rlabel polysilicon 366 -3490 366 -3490 0 1
rlabel polysilicon 369 -3490 369 -3490 0 2
rlabel polysilicon 387 -3490 387 -3490 0 1
rlabel polysilicon 387 -3496 387 -3496 0 3
rlabel polysilicon 394 -3490 394 -3490 0 1
rlabel polysilicon 394 -3496 394 -3496 0 3
rlabel polysilicon 429 -3490 429 -3490 0 1
rlabel polysilicon 429 -3496 429 -3496 0 3
rlabel polysilicon 432 -3496 432 -3496 0 4
rlabel polysilicon 464 -3490 464 -3490 0 1
rlabel polysilicon 464 -3496 464 -3496 0 3
rlabel polysilicon 471 -3490 471 -3490 0 1
rlabel polysilicon 471 -3496 471 -3496 0 3
rlabel polysilicon 478 -3490 478 -3490 0 1
rlabel polysilicon 478 -3496 478 -3496 0 3
rlabel polysilicon 485 -3490 485 -3490 0 1
rlabel polysilicon 485 -3496 485 -3496 0 3
rlabel polysilicon 523 -3490 523 -3490 0 2
rlabel polysilicon 523 -3496 523 -3496 0 4
rlabel polysilicon 534 -3490 534 -3490 0 1
rlabel polysilicon 534 -3496 534 -3496 0 3
rlabel polysilicon 541 -3490 541 -3490 0 1
rlabel polysilicon 541 -3496 541 -3496 0 3
rlabel polysilicon 569 -3490 569 -3490 0 1
rlabel polysilicon 569 -3496 569 -3496 0 3
rlabel polysilicon 583 -3490 583 -3490 0 1
rlabel polysilicon 583 -3496 583 -3496 0 3
rlabel polysilicon 590 -3490 590 -3490 0 1
rlabel polysilicon 590 -3496 590 -3496 0 3
rlabel polysilicon 604 -3490 604 -3490 0 1
rlabel polysilicon 604 -3496 604 -3496 0 3
rlabel polysilicon 611 -3490 611 -3490 0 1
rlabel polysilicon 611 -3496 611 -3496 0 3
rlabel polysilicon 618 -3490 618 -3490 0 1
rlabel polysilicon 618 -3496 618 -3496 0 3
rlabel polysilicon 632 -3490 632 -3490 0 1
rlabel polysilicon 632 -3496 632 -3496 0 3
rlabel polysilicon 639 -3490 639 -3490 0 1
rlabel polysilicon 639 -3496 639 -3496 0 3
rlabel polysilicon 646 -3490 646 -3490 0 1
rlabel polysilicon 646 -3496 646 -3496 0 3
rlabel polysilicon 653 -3490 653 -3490 0 1
rlabel polysilicon 653 -3496 653 -3496 0 3
rlabel polysilicon 656 -3496 656 -3496 0 4
rlabel polysilicon 681 -3490 681 -3490 0 1
rlabel polysilicon 681 -3496 681 -3496 0 3
rlabel polysilicon 716 -3490 716 -3490 0 1
rlabel polysilicon 716 -3496 716 -3496 0 3
rlabel polysilicon 737 -3490 737 -3490 0 1
rlabel polysilicon 737 -3496 737 -3496 0 3
rlabel polysilicon 744 -3490 744 -3490 0 1
rlabel polysilicon 744 -3496 744 -3496 0 3
rlabel polysilicon 751 -3490 751 -3490 0 1
rlabel polysilicon 751 -3496 751 -3496 0 3
rlabel polysilicon 758 -3490 758 -3490 0 1
rlabel polysilicon 758 -3496 758 -3496 0 3
rlabel polysilicon 765 -3490 765 -3490 0 1
rlabel polysilicon 765 -3496 765 -3496 0 3
rlabel polysilicon 772 -3490 772 -3490 0 1
rlabel polysilicon 772 -3496 772 -3496 0 3
rlabel polysilicon 779 -3490 779 -3490 0 1
rlabel polysilicon 779 -3496 779 -3496 0 3
rlabel polysilicon 786 -3490 786 -3490 0 1
rlabel polysilicon 789 -3490 789 -3490 0 2
rlabel polysilicon 793 -3490 793 -3490 0 1
rlabel polysilicon 793 -3496 793 -3496 0 3
rlabel polysilicon 814 -3490 814 -3490 0 1
rlabel polysilicon 814 -3496 814 -3496 0 3
rlabel polysilicon 828 -3490 828 -3490 0 1
rlabel polysilicon 828 -3496 828 -3496 0 3
rlabel polysilicon 842 -3490 842 -3490 0 1
rlabel polysilicon 842 -3496 842 -3496 0 3
rlabel polysilicon 866 -3490 866 -3490 0 2
rlabel polysilicon 863 -3496 863 -3496 0 3
rlabel polysilicon 866 -3496 866 -3496 0 4
rlabel polysilicon 870 -3490 870 -3490 0 1
rlabel polysilicon 870 -3496 870 -3496 0 3
rlabel polysilicon 887 -3490 887 -3490 0 2
rlabel polysilicon 884 -3496 884 -3496 0 3
rlabel polysilicon 898 -3490 898 -3490 0 1
rlabel polysilicon 898 -3496 898 -3496 0 3
rlabel polysilicon 975 -3490 975 -3490 0 1
rlabel polysilicon 975 -3496 975 -3496 0 3
rlabel polysilicon 996 -3496 996 -3496 0 3
rlabel polysilicon 1010 -3490 1010 -3490 0 1
rlabel polysilicon 1010 -3496 1010 -3496 0 3
rlabel polysilicon 1017 -3490 1017 -3490 0 1
rlabel polysilicon 1017 -3496 1017 -3496 0 3
rlabel polysilicon 1024 -3490 1024 -3490 0 1
rlabel polysilicon 1024 -3496 1024 -3496 0 3
rlabel polysilicon 1031 -3490 1031 -3490 0 1
rlabel polysilicon 1031 -3496 1031 -3496 0 3
rlabel polysilicon 1038 -3490 1038 -3490 0 1
rlabel polysilicon 1038 -3496 1038 -3496 0 3
rlabel polysilicon 1045 -3490 1045 -3490 0 1
rlabel polysilicon 1045 -3496 1045 -3496 0 3
rlabel polysilicon 1052 -3490 1052 -3490 0 1
rlabel polysilicon 1052 -3496 1052 -3496 0 3
rlabel polysilicon 1059 -3490 1059 -3490 0 1
rlabel polysilicon 1059 -3496 1059 -3496 0 3
rlabel polysilicon 1066 -3490 1066 -3490 0 1
rlabel polysilicon 1066 -3496 1066 -3496 0 3
rlabel polysilicon 1080 -3490 1080 -3490 0 1
rlabel polysilicon 1080 -3496 1080 -3496 0 3
rlabel polysilicon 1143 -3490 1143 -3490 0 1
rlabel polysilicon 1143 -3496 1143 -3496 0 3
rlabel polysilicon 1178 -3490 1178 -3490 0 1
rlabel polysilicon 1178 -3496 1178 -3496 0 3
rlabel polysilicon 1192 -3490 1192 -3490 0 1
rlabel polysilicon 1192 -3496 1192 -3496 0 3
rlabel polysilicon 1234 -3490 1234 -3490 0 1
rlabel polysilicon 1234 -3496 1234 -3496 0 3
rlabel polysilicon 1241 -3490 1241 -3490 0 1
rlabel polysilicon 1241 -3496 1241 -3496 0 3
rlabel polysilicon 1248 -3490 1248 -3490 0 1
rlabel polysilicon 1248 -3496 1248 -3496 0 3
rlabel polysilicon 1251 -3496 1251 -3496 0 4
rlabel polysilicon 1255 -3490 1255 -3490 0 1
rlabel polysilicon 1255 -3496 1255 -3496 0 3
rlabel polysilicon 1262 -3490 1262 -3490 0 1
rlabel polysilicon 1262 -3496 1262 -3496 0 3
rlabel polysilicon 1269 -3490 1269 -3490 0 1
rlabel polysilicon 1272 -3490 1272 -3490 0 2
rlabel polysilicon 1276 -3490 1276 -3490 0 1
rlabel polysilicon 1276 -3496 1276 -3496 0 3
rlabel polysilicon 1286 -3490 1286 -3490 0 2
rlabel polysilicon 1283 -3496 1283 -3496 0 3
rlabel polysilicon 1290 -3490 1290 -3490 0 1
rlabel polysilicon 1290 -3496 1290 -3496 0 3
rlabel polysilicon 1304 -3490 1304 -3490 0 1
rlabel polysilicon 1304 -3496 1304 -3496 0 3
rlabel polysilicon 1311 -3490 1311 -3490 0 1
rlabel polysilicon 1311 -3496 1311 -3496 0 3
rlabel polysilicon 1360 -3490 1360 -3490 0 1
rlabel polysilicon 1360 -3496 1360 -3496 0 3
rlabel polysilicon 1430 -3490 1430 -3490 0 1
rlabel polysilicon 1433 -3490 1433 -3490 0 2
rlabel polysilicon 1430 -3496 1430 -3496 0 3
rlabel polysilicon 1437 -3490 1437 -3490 0 1
rlabel polysilicon 1437 -3496 1437 -3496 0 3
rlabel polysilicon 1493 -3490 1493 -3490 0 1
rlabel polysilicon 1493 -3496 1493 -3496 0 3
rlabel polysilicon 1500 -3490 1500 -3490 0 1
rlabel polysilicon 1503 -3490 1503 -3490 0 2
rlabel polysilicon 1500 -3496 1500 -3496 0 3
rlabel polysilicon 1507 -3490 1507 -3490 0 1
rlabel polysilicon 1507 -3496 1507 -3496 0 3
rlabel polysilicon 1514 -3490 1514 -3490 0 1
rlabel polysilicon 1514 -3496 1514 -3496 0 3
rlabel polysilicon 1521 -3490 1521 -3490 0 1
rlabel polysilicon 1521 -3496 1521 -3496 0 3
rlabel polysilicon 1570 -3490 1570 -3490 0 1
rlabel polysilicon 1570 -3496 1570 -3496 0 3
rlabel polysilicon 1640 -3490 1640 -3490 0 1
rlabel polysilicon 1640 -3496 1640 -3496 0 3
rlabel polysilicon 1724 -3490 1724 -3490 0 1
rlabel polysilicon 1727 -3490 1727 -3490 0 2
rlabel polysilicon 1724 -3496 1724 -3496 0 3
rlabel polysilicon 1731 -3490 1731 -3490 0 1
rlabel polysilicon 1731 -3496 1731 -3496 0 3
rlabel polysilicon 1780 -3490 1780 -3490 0 1
rlabel polysilicon 1780 -3496 1780 -3496 0 3
rlabel polysilicon 1790 -3490 1790 -3490 0 2
rlabel polysilicon 1790 -3496 1790 -3496 0 4
rlabel polysilicon 1843 -3490 1843 -3490 0 1
rlabel polysilicon 1843 -3496 1843 -3496 0 3
rlabel polysilicon 1850 -3490 1850 -3490 0 1
rlabel polysilicon 1850 -3496 1850 -3496 0 3
rlabel polysilicon 1864 -3490 1864 -3490 0 1
rlabel polysilicon 1864 -3496 1864 -3496 0 3
rlabel polysilicon 1955 -3490 1955 -3490 0 1
rlabel polysilicon 1958 -3490 1958 -3490 0 2
rlabel polysilicon 2025 -3490 2025 -3490 0 1
rlabel polysilicon 2028 -3490 2028 -3490 0 2
rlabel polysilicon 2025 -3496 2025 -3496 0 3
rlabel polysilicon 2032 -3490 2032 -3490 0 1
rlabel polysilicon 2032 -3496 2032 -3496 0 3
rlabel polysilicon 338 -3513 338 -3513 0 1
rlabel polysilicon 394 -3513 394 -3513 0 1
rlabel polysilicon 394 -3519 394 -3519 0 3
rlabel polysilicon 429 -3513 429 -3513 0 1
rlabel polysilicon 429 -3519 429 -3519 0 3
rlabel polysilicon 464 -3513 464 -3513 0 1
rlabel polysilicon 464 -3519 464 -3519 0 3
rlabel polysilicon 478 -3513 478 -3513 0 1
rlabel polysilicon 478 -3519 478 -3519 0 3
rlabel polysilicon 541 -3513 541 -3513 0 1
rlabel polysilicon 541 -3519 541 -3519 0 3
rlabel polysilicon 548 -3513 548 -3513 0 1
rlabel polysilicon 548 -3519 548 -3519 0 3
rlabel polysilicon 576 -3513 576 -3513 0 1
rlabel polysilicon 576 -3519 576 -3519 0 3
rlabel polysilicon 583 -3513 583 -3513 0 1
rlabel polysilicon 583 -3519 583 -3519 0 3
rlabel polysilicon 604 -3513 604 -3513 0 1
rlabel polysilicon 604 -3519 604 -3519 0 3
rlabel polysilicon 611 -3513 611 -3513 0 1
rlabel polysilicon 611 -3519 611 -3519 0 3
rlabel polysilicon 618 -3513 618 -3513 0 1
rlabel polysilicon 618 -3519 618 -3519 0 3
rlabel polysilicon 625 -3513 625 -3513 0 1
rlabel polysilicon 625 -3519 625 -3519 0 3
rlabel polysilicon 632 -3513 632 -3513 0 1
rlabel polysilicon 632 -3519 632 -3519 0 3
rlabel polysilicon 639 -3513 639 -3513 0 1
rlabel polysilicon 639 -3519 639 -3519 0 3
rlabel polysilicon 709 -3513 709 -3513 0 1
rlabel polysilicon 709 -3519 709 -3519 0 3
rlabel polysilicon 730 -3513 730 -3513 0 1
rlabel polysilicon 730 -3519 730 -3519 0 3
rlabel polysilicon 737 -3513 737 -3513 0 1
rlabel polysilicon 737 -3519 737 -3519 0 3
rlabel polysilicon 744 -3513 744 -3513 0 1
rlabel polysilicon 744 -3519 744 -3519 0 3
rlabel polysilicon 751 -3513 751 -3513 0 1
rlabel polysilicon 751 -3519 751 -3519 0 3
rlabel polysilicon 758 -3513 758 -3513 0 1
rlabel polysilicon 758 -3519 758 -3519 0 3
rlabel polysilicon 765 -3513 765 -3513 0 1
rlabel polysilicon 765 -3519 765 -3519 0 3
rlabel polysilicon 775 -3513 775 -3513 0 2
rlabel polysilicon 772 -3519 772 -3519 0 3
rlabel polysilicon 775 -3519 775 -3519 0 4
rlabel polysilicon 779 -3513 779 -3513 0 1
rlabel polysilicon 779 -3519 779 -3519 0 3
rlabel polysilicon 789 -3513 789 -3513 0 2
rlabel polysilicon 786 -3519 786 -3519 0 3
rlabel polysilicon 789 -3519 789 -3519 0 4
rlabel polysilicon 793 -3513 793 -3513 0 1
rlabel polysilicon 793 -3519 793 -3519 0 3
rlabel polysilicon 800 -3513 800 -3513 0 1
rlabel polysilicon 800 -3519 800 -3519 0 3
rlabel polysilicon 810 -3513 810 -3513 0 2
rlabel polysilicon 810 -3519 810 -3519 0 4
rlabel polysilicon 891 -3513 891 -3513 0 1
rlabel polysilicon 891 -3519 891 -3519 0 3
rlabel polysilicon 968 -3513 968 -3513 0 1
rlabel polysilicon 968 -3519 968 -3519 0 3
rlabel polysilicon 1003 -3513 1003 -3513 0 1
rlabel polysilicon 1003 -3519 1003 -3519 0 3
rlabel polysilicon 1010 -3513 1010 -3513 0 1
rlabel polysilicon 1010 -3519 1010 -3519 0 3
rlabel polysilicon 1017 -3513 1017 -3513 0 1
rlabel polysilicon 1017 -3519 1017 -3519 0 3
rlabel polysilicon 1024 -3513 1024 -3513 0 1
rlabel polysilicon 1024 -3519 1024 -3519 0 3
rlabel polysilicon 1031 -3513 1031 -3513 0 1
rlabel polysilicon 1031 -3519 1031 -3519 0 3
rlabel polysilicon 1038 -3513 1038 -3513 0 1
rlabel polysilicon 1038 -3519 1038 -3519 0 3
rlabel polysilicon 1045 -3513 1045 -3513 0 1
rlabel polysilicon 1052 -3513 1052 -3513 0 1
rlabel polysilicon 1052 -3519 1052 -3519 0 3
rlabel polysilicon 1059 -3513 1059 -3513 0 1
rlabel polysilicon 1062 -3513 1062 -3513 0 2
rlabel polysilicon 1059 -3519 1059 -3519 0 3
rlabel polysilicon 1066 -3513 1066 -3513 0 1
rlabel polysilicon 1066 -3519 1066 -3519 0 3
rlabel polysilicon 1122 -3513 1122 -3513 0 1
rlabel polysilicon 1122 -3519 1122 -3519 0 3
rlabel polysilicon 1150 -3513 1150 -3513 0 1
rlabel polysilicon 1150 -3519 1150 -3519 0 3
rlabel polysilicon 1160 -3513 1160 -3513 0 2
rlabel polysilicon 1157 -3519 1157 -3519 0 3
rlabel polysilicon 1160 -3519 1160 -3519 0 4
rlabel polysilicon 1206 -3513 1206 -3513 0 1
rlabel polysilicon 1206 -3519 1206 -3519 0 3
rlabel polysilicon 1234 -3513 1234 -3513 0 1
rlabel polysilicon 1234 -3519 1234 -3519 0 3
rlabel polysilicon 1360 -3513 1360 -3513 0 1
rlabel polysilicon 1360 -3519 1360 -3519 0 3
rlabel polysilicon 1367 -3513 1367 -3513 0 1
rlabel polysilicon 1367 -3519 1367 -3519 0 3
rlabel polysilicon 1507 -3513 1507 -3513 0 1
rlabel polysilicon 1507 -3519 1507 -3519 0 3
rlabel polysilicon 1510 -3519 1510 -3519 0 4
rlabel polysilicon 1514 -3513 1514 -3513 0 1
rlabel polysilicon 1514 -3519 1514 -3519 0 3
rlabel polysilicon 1521 -3513 1521 -3513 0 1
rlabel polysilicon 1521 -3519 1521 -3519 0 3
rlabel polysilicon 1612 -3513 1612 -3513 0 1
rlabel polysilicon 1612 -3519 1612 -3519 0 3
rlabel polysilicon 1640 -3513 1640 -3513 0 1
rlabel polysilicon 1640 -3519 1640 -3519 0 3
rlabel polysilicon 1850 -3513 1850 -3513 0 1
rlabel polysilicon 1850 -3519 1850 -3519 0 3
rlabel polysilicon 1857 -3513 1857 -3513 0 1
rlabel polysilicon 1860 -3513 1860 -3513 0 2
rlabel polysilicon 1857 -3519 1857 -3519 0 3
rlabel polysilicon 2025 -3513 2025 -3513 0 1
rlabel polysilicon 2025 -3519 2025 -3519 0 3
rlabel polysilicon 2032 -3513 2032 -3513 0 1
rlabel polysilicon 2032 -3519 2032 -3519 0 3
rlabel polysilicon 394 -3532 394 -3532 0 1
rlabel polysilicon 394 -3538 394 -3538 0 3
rlabel polysilicon 408 -3532 408 -3532 0 1
rlabel polysilicon 408 -3538 408 -3538 0 3
rlabel polysilicon 464 -3532 464 -3532 0 1
rlabel polysilicon 464 -3538 464 -3538 0 3
rlabel polysilicon 471 -3538 471 -3538 0 3
rlabel polysilicon 474 -3538 474 -3538 0 4
rlabel polysilicon 478 -3532 478 -3532 0 1
rlabel polysilicon 478 -3538 478 -3538 0 3
rlabel polysilicon 541 -3532 541 -3532 0 1
rlabel polysilicon 541 -3538 541 -3538 0 3
rlabel polysilicon 548 -3532 548 -3532 0 1
rlabel polysilicon 548 -3538 548 -3538 0 3
rlabel polysilicon 576 -3532 576 -3532 0 1
rlabel polysilicon 576 -3538 576 -3538 0 3
rlabel polysilicon 583 -3532 583 -3532 0 1
rlabel polysilicon 583 -3538 583 -3538 0 3
rlabel polysilicon 604 -3532 604 -3532 0 1
rlabel polysilicon 604 -3538 604 -3538 0 3
rlabel polysilicon 611 -3532 611 -3532 0 1
rlabel polysilicon 611 -3538 611 -3538 0 3
rlabel polysilicon 618 -3532 618 -3532 0 1
rlabel polysilicon 618 -3538 618 -3538 0 3
rlabel polysilicon 625 -3532 625 -3532 0 1
rlabel polysilicon 632 -3532 632 -3532 0 1
rlabel polysilicon 635 -3532 635 -3532 0 2
rlabel polysilicon 635 -3538 635 -3538 0 4
rlabel polysilicon 639 -3532 639 -3532 0 1
rlabel polysilicon 639 -3538 639 -3538 0 3
rlabel polysilicon 646 -3532 646 -3532 0 1
rlabel polysilicon 646 -3538 646 -3538 0 3
rlabel polysilicon 709 -3532 709 -3532 0 1
rlabel polysilicon 709 -3538 709 -3538 0 3
rlabel polysilicon 716 -3532 716 -3532 0 1
rlabel polysilicon 716 -3538 716 -3538 0 3
rlabel polysilicon 723 -3532 723 -3532 0 1
rlabel polysilicon 723 -3538 723 -3538 0 3
rlabel polysilicon 730 -3532 730 -3532 0 1
rlabel polysilicon 730 -3538 730 -3538 0 3
rlabel polysilicon 740 -3532 740 -3532 0 2
rlabel polysilicon 740 -3538 740 -3538 0 4
rlabel polysilicon 744 -3532 744 -3532 0 1
rlabel polysilicon 744 -3538 744 -3538 0 3
rlabel polysilicon 765 -3532 765 -3532 0 1
rlabel polysilicon 765 -3538 765 -3538 0 3
rlabel polysilicon 786 -3532 786 -3532 0 1
rlabel polysilicon 786 -3538 786 -3538 0 3
rlabel polysilicon 793 -3532 793 -3532 0 1
rlabel polysilicon 793 -3538 793 -3538 0 3
rlabel polysilicon 926 -3532 926 -3532 0 1
rlabel polysilicon 926 -3538 926 -3538 0 3
rlabel polysilicon 971 -3532 971 -3532 0 2
rlabel polysilicon 968 -3538 968 -3538 0 3
rlabel polysilicon 1010 -3532 1010 -3532 0 1
rlabel polysilicon 1010 -3538 1010 -3538 0 3
rlabel polysilicon 1024 -3532 1024 -3532 0 1
rlabel polysilicon 1027 -3532 1027 -3532 0 2
rlabel polysilicon 1027 -3538 1027 -3538 0 4
rlabel polysilicon 1031 -3532 1031 -3532 0 1
rlabel polysilicon 1031 -3538 1031 -3538 0 3
rlabel polysilicon 1038 -3532 1038 -3532 0 1
rlabel polysilicon 1038 -3538 1038 -3538 0 3
rlabel polysilicon 1045 -3538 1045 -3538 0 3
rlabel polysilicon 1059 -3532 1059 -3532 0 1
rlabel polysilicon 1059 -3538 1059 -3538 0 3
rlabel polysilicon 1066 -3532 1066 -3532 0 1
rlabel polysilicon 1066 -3538 1066 -3538 0 3
rlabel polysilicon 1213 -3532 1213 -3532 0 1
rlabel polysilicon 1213 -3538 1213 -3538 0 3
rlabel polysilicon 1223 -3532 1223 -3532 0 2
rlabel polysilicon 1223 -3538 1223 -3538 0 4
rlabel polysilicon 1507 -3532 1507 -3532 0 1
rlabel polysilicon 1510 -3532 1510 -3532 0 2
rlabel polysilicon 1507 -3538 1507 -3538 0 3
rlabel polysilicon 1514 -3532 1514 -3532 0 1
rlabel polysilicon 1514 -3538 1514 -3538 0 3
rlabel polysilicon 1521 -3532 1521 -3532 0 1
rlabel polysilicon 1521 -3538 1521 -3538 0 3
rlabel polysilicon 1633 -3532 1633 -3532 0 1
rlabel polysilicon 1633 -3538 1633 -3538 0 3
rlabel polysilicon 1640 -3532 1640 -3532 0 1
rlabel polysilicon 1640 -3538 1640 -3538 0 3
rlabel polysilicon 2025 -3532 2025 -3532 0 1
rlabel polysilicon 2025 -3538 2025 -3538 0 3
rlabel polysilicon 2032 -3532 2032 -3532 0 1
rlabel polysilicon 2032 -3538 2032 -3538 0 3
rlabel polysilicon 401 -3547 401 -3547 0 1
rlabel polysilicon 401 -3553 401 -3553 0 3
rlabel polysilicon 408 -3547 408 -3547 0 1
rlabel polysilicon 541 -3547 541 -3547 0 1
rlabel polysilicon 541 -3553 541 -3553 0 3
rlabel polysilicon 548 -3553 548 -3553 0 3
rlabel polysilicon 551 -3553 551 -3553 0 4
rlabel polysilicon 555 -3547 555 -3547 0 1
rlabel polysilicon 555 -3553 555 -3553 0 3
rlabel polysilicon 583 -3547 583 -3547 0 1
rlabel polysilicon 586 -3553 586 -3553 0 4
rlabel polysilicon 590 -3547 590 -3547 0 1
rlabel polysilicon 590 -3553 590 -3553 0 3
rlabel polysilicon 604 -3547 604 -3547 0 1
rlabel polysilicon 604 -3553 604 -3553 0 3
rlabel polysilicon 607 -3553 607 -3553 0 4
rlabel polysilicon 611 -3547 611 -3547 0 1
rlabel polysilicon 611 -3553 611 -3553 0 3
rlabel polysilicon 618 -3547 618 -3547 0 1
rlabel polysilicon 618 -3553 618 -3553 0 3
rlabel polysilicon 646 -3547 646 -3547 0 1
rlabel polysilicon 646 -3553 646 -3553 0 3
rlabel polysilicon 702 -3547 702 -3547 0 1
rlabel polysilicon 702 -3553 702 -3553 0 3
rlabel polysilicon 716 -3547 716 -3547 0 1
rlabel polysilicon 716 -3553 716 -3553 0 3
rlabel polysilicon 723 -3547 723 -3547 0 1
rlabel polysilicon 723 -3553 723 -3553 0 3
rlabel polysilicon 730 -3547 730 -3547 0 1
rlabel polysilicon 730 -3553 730 -3553 0 3
rlabel polysilicon 758 -3547 758 -3547 0 1
rlabel polysilicon 758 -3553 758 -3553 0 3
rlabel polysilicon 789 -3547 789 -3547 0 2
rlabel polysilicon 789 -3553 789 -3553 0 4
rlabel polysilicon 793 -3547 793 -3547 0 1
rlabel polysilicon 793 -3553 793 -3553 0 3
rlabel polysilicon 1020 -3547 1020 -3547 0 2
rlabel polysilicon 1017 -3553 1017 -3553 0 3
rlabel polysilicon 1038 -3547 1038 -3547 0 1
rlabel polysilicon 1038 -3553 1038 -3553 0 3
rlabel polysilicon 1059 -3547 1059 -3547 0 1
rlabel polysilicon 1059 -3553 1059 -3553 0 3
rlabel polysilicon 1507 -3547 1507 -3547 0 1
rlabel polysilicon 1507 -3553 1507 -3553 0 3
rlabel polysilicon 1514 -3547 1514 -3547 0 1
rlabel polysilicon 1514 -3553 1514 -3553 0 3
rlabel polysilicon 1521 -3547 1521 -3547 0 1
rlabel polysilicon 1521 -3553 1521 -3553 0 3
rlabel polysilicon 1640 -3547 1640 -3547 0 1
rlabel polysilicon 1640 -3553 1640 -3553 0 3
rlabel polysilicon 1647 -3547 1647 -3547 0 1
rlabel polysilicon 1647 -3553 1647 -3553 0 3
rlabel polysilicon 2025 -3547 2025 -3547 0 1
rlabel polysilicon 2025 -3553 2025 -3553 0 3
rlabel polysilicon 2032 -3547 2032 -3547 0 1
rlabel polysilicon 2032 -3553 2032 -3553 0 3
rlabel polysilicon 401 -3562 401 -3562 0 1
rlabel polysilicon 401 -3568 401 -3568 0 3
rlabel polysilicon 408 -3568 408 -3568 0 3
rlabel polysilicon 604 -3562 604 -3562 0 1
rlabel polysilicon 607 -3562 607 -3562 0 2
rlabel polysilicon 604 -3568 604 -3568 0 3
rlabel polysilicon 611 -3562 611 -3562 0 1
rlabel polysilicon 611 -3568 611 -3568 0 3
rlabel polysilicon 618 -3562 618 -3562 0 1
rlabel polysilicon 618 -3568 618 -3568 0 3
rlabel polysilicon 649 -3562 649 -3562 0 2
rlabel polysilicon 702 -3562 702 -3562 0 1
rlabel polysilicon 702 -3568 702 -3568 0 3
rlabel polysilicon 716 -3562 716 -3562 0 1
rlabel polysilicon 716 -3568 716 -3568 0 3
rlabel polysilicon 723 -3562 723 -3562 0 1
rlabel polysilicon 723 -3568 723 -3568 0 3
rlabel polysilicon 730 -3562 730 -3562 0 1
rlabel polysilicon 730 -3568 730 -3568 0 3
rlabel polysilicon 758 -3562 758 -3562 0 1
rlabel polysilicon 758 -3568 758 -3568 0 3
rlabel polysilicon 1062 -3568 1062 -3568 0 4
rlabel polysilicon 1066 -3562 1066 -3562 0 1
rlabel polysilicon 1066 -3568 1066 -3568 0 3
rlabel polysilicon 1514 -3562 1514 -3562 0 1
rlabel polysilicon 1517 -3562 1517 -3562 0 2
rlabel polysilicon 1514 -3568 1514 -3568 0 3
rlabel polysilicon 1521 -3562 1521 -3562 0 1
rlabel polysilicon 1521 -3568 1521 -3568 0 3
rlabel polysilicon 1640 -3562 1640 -3562 0 1
rlabel polysilicon 1640 -3568 1640 -3568 0 3
rlabel polysilicon 1647 -3562 1647 -3562 0 1
rlabel polysilicon 1647 -3568 1647 -3568 0 3
rlabel polysilicon 2025 -3562 2025 -3562 0 1
rlabel polysilicon 2028 -3562 2028 -3562 0 2
rlabel polysilicon 401 -3577 401 -3577 0 1
rlabel polysilicon 401 -3583 401 -3583 0 3
rlabel polysilicon 408 -3577 408 -3577 0 1
rlabel polysilicon 408 -3583 408 -3583 0 3
rlabel polysilicon 604 -3577 604 -3577 0 1
rlabel polysilicon 604 -3583 604 -3583 0 3
rlabel polysilicon 611 -3577 611 -3577 0 1
rlabel polysilicon 611 -3583 611 -3583 0 3
rlabel polysilicon 618 -3577 618 -3577 0 1
rlabel polysilicon 618 -3583 618 -3583 0 3
rlabel polysilicon 702 -3577 702 -3577 0 1
rlabel polysilicon 702 -3583 702 -3583 0 3
rlabel polysilicon 716 -3577 716 -3577 0 1
rlabel polysilicon 716 -3583 716 -3583 0 3
rlabel polysilicon 723 -3577 723 -3577 0 1
rlabel polysilicon 723 -3583 723 -3583 0 3
rlabel polysilicon 730 -3577 730 -3577 0 1
rlabel polysilicon 730 -3583 730 -3583 0 3
rlabel polysilicon 758 -3577 758 -3577 0 1
rlabel polysilicon 758 -3583 758 -3583 0 3
rlabel polysilicon 1640 -3577 1640 -3577 0 1
rlabel polysilicon 1640 -3583 1640 -3583 0 3
rlabel polysilicon 1647 -3577 1647 -3577 0 1
rlabel polysilicon 1647 -3583 1647 -3583 0 3
rlabel polysilicon 394 -3590 394 -3590 0 1
rlabel polysilicon 394 -3596 394 -3596 0 3
rlabel polysilicon 401 -3590 401 -3590 0 1
rlabel polysilicon 401 -3596 401 -3596 0 3
rlabel polysilicon 604 -3590 604 -3590 0 1
rlabel polysilicon 604 -3596 604 -3596 0 3
rlabel polysilicon 611 -3590 611 -3590 0 1
rlabel polysilicon 611 -3596 611 -3596 0 3
rlabel polysilicon 621 -3590 621 -3590 0 2
rlabel polysilicon 702 -3590 702 -3590 0 1
rlabel polysilicon 702 -3596 702 -3596 0 3
rlabel polysilicon 723 -3590 723 -3590 0 1
rlabel polysilicon 726 -3590 726 -3590 0 2
rlabel polysilicon 723 -3596 723 -3596 0 3
rlabel polysilicon 730 -3590 730 -3590 0 1
rlabel polysilicon 730 -3596 730 -3596 0 3
rlabel polysilicon 758 -3590 758 -3590 0 1
rlabel polysilicon 758 -3596 758 -3596 0 3
rlabel polysilicon 1640 -3590 1640 -3590 0 1
rlabel polysilicon 1640 -3596 1640 -3596 0 3
rlabel polysilicon 1647 -3590 1647 -3590 0 1
rlabel polysilicon 1647 -3596 1647 -3596 0 3
rlabel polysilicon 394 -3601 394 -3601 0 1
rlabel polysilicon 394 -3607 394 -3607 0 3
rlabel polysilicon 401 -3601 401 -3601 0 1
rlabel polysilicon 401 -3607 401 -3607 0 3
rlabel polysilicon 604 -3601 604 -3601 0 1
rlabel polysilicon 604 -3607 604 -3607 0 3
rlabel polysilicon 611 -3601 611 -3601 0 1
rlabel polysilicon 611 -3607 611 -3607 0 3
rlabel polysilicon 702 -3601 702 -3601 0 1
rlabel polysilicon 705 -3607 705 -3607 0 4
rlabel polysilicon 758 -3601 758 -3601 0 1
rlabel polysilicon 758 -3607 758 -3607 0 3
rlabel polysilicon 1640 -3601 1640 -3601 0 1
rlabel polysilicon 1640 -3607 1640 -3607 0 3
rlabel polysilicon 1647 -3601 1647 -3601 0 1
rlabel polysilicon 1647 -3607 1647 -3607 0 3
rlabel polysilicon 394 -3612 394 -3612 0 1
rlabel polysilicon 394 -3618 394 -3618 0 3
rlabel polysilicon 401 -3612 401 -3612 0 1
rlabel polysilicon 401 -3618 401 -3618 0 3
rlabel polysilicon 604 -3612 604 -3612 0 1
rlabel polysilicon 604 -3618 604 -3618 0 3
rlabel polysilicon 611 -3612 611 -3612 0 1
rlabel polysilicon 611 -3618 611 -3618 0 3
rlabel polysilicon 695 -3612 695 -3612 0 1
rlabel polysilicon 695 -3618 695 -3618 0 3
rlabel polysilicon 758 -3612 758 -3612 0 1
rlabel polysilicon 758 -3618 758 -3618 0 3
rlabel polysilicon 1643 -3612 1643 -3612 0 2
rlabel polysilicon 1640 -3618 1640 -3618 0 3
rlabel polysilicon 1647 -3612 1647 -3612 0 1
rlabel polysilicon 1647 -3618 1647 -3618 0 3
rlabel polysilicon 394 -3623 394 -3623 0 1
rlabel polysilicon 394 -3629 394 -3629 0 3
rlabel polysilicon 401 -3623 401 -3623 0 1
rlabel polysilicon 401 -3629 401 -3629 0 3
rlabel polysilicon 604 -3623 604 -3623 0 1
rlabel polysilicon 604 -3629 604 -3629 0 3
rlabel polysilicon 611 -3623 611 -3623 0 1
rlabel polysilicon 611 -3629 611 -3629 0 3
rlabel polysilicon 695 -3623 695 -3623 0 1
rlabel polysilicon 695 -3629 695 -3629 0 3
rlabel polysilicon 761 -3629 761 -3629 0 4
rlabel polysilicon 765 -3623 765 -3623 0 1
rlabel polysilicon 765 -3629 765 -3629 0 3
rlabel polysilicon 394 -3634 394 -3634 0 1
rlabel polysilicon 394 -3640 394 -3640 0 3
rlabel polysilicon 401 -3634 401 -3634 0 1
rlabel polysilicon 401 -3640 401 -3640 0 3
rlabel polysilicon 604 -3634 604 -3634 0 1
rlabel polysilicon 604 -3640 604 -3640 0 3
rlabel polysilicon 611 -3634 611 -3634 0 1
rlabel polysilicon 611 -3640 611 -3640 0 3
rlabel polysilicon 695 -3634 695 -3634 0 1
rlabel polysilicon 695 -3640 695 -3640 0 3
rlabel polysilicon 394 -3645 394 -3645 0 1
rlabel polysilicon 394 -3651 394 -3651 0 3
rlabel polysilicon 401 -3645 401 -3645 0 1
rlabel polysilicon 401 -3651 401 -3651 0 3
rlabel polysilicon 604 -3645 604 -3645 0 1
rlabel polysilicon 604 -3651 604 -3651 0 3
rlabel polysilicon 611 -3645 611 -3645 0 1
rlabel polysilicon 611 -3651 611 -3651 0 3
rlabel polysilicon 695 -3645 695 -3645 0 1
rlabel polysilicon 695 -3651 695 -3651 0 3
rlabel polysilicon 394 -3660 394 -3660 0 1
rlabel polysilicon 397 -3666 397 -3666 0 4
rlabel polysilicon 401 -3660 401 -3660 0 1
rlabel polysilicon 401 -3666 401 -3666 0 3
rlabel polysilicon 604 -3660 604 -3660 0 1
rlabel polysilicon 604 -3666 604 -3666 0 3
rlabel polysilicon 611 -3660 611 -3660 0 1
rlabel polysilicon 611 -3666 611 -3666 0 3
rlabel polysilicon 698 -3660 698 -3660 0 2
rlabel metal2 254 1 254 1 0 net=5879
rlabel metal2 485 1 485 1 0 net=3145
rlabel metal2 635 1 635 1 0 net=8547
rlabel metal2 796 1 796 1 0 net=12633
rlabel metal2 824 1 824 1 0 net=12941
rlabel metal2 968 1 968 1 0 net=9893
rlabel metal2 352 -1 352 -1 0 net=2965
rlabel metal2 576 -1 576 -1 0 net=4031
rlabel metal2 688 -1 688 -1 0 net=3723
rlabel metal2 800 -1 800 -1 0 net=13789
rlabel metal2 978 -1 978 -1 0 net=9101
rlabel metal2 1038 -1 1038 -1 0 net=4921
rlabel metal2 397 -3 397 -3 0 net=6197
rlabel metal2 555 -3 555 -3 0 net=11131
rlabel metal2 604 -3 604 -3 0 net=2837
rlabel metal2 863 -3 863 -3 0 net=5933
rlabel metal2 1073 -3 1073 -3 0 net=14095
rlabel metal2 415 -5 415 -5 0 net=7257
rlabel metal2 611 -5 611 -5 0 net=6261
rlabel metal2 639 -5 639 -5 0 net=1689
rlabel metal2 884 -5 884 -5 0 net=11987
rlabel metal2 1094 -5 1094 -5 0 net=6981
rlabel metal2 618 -7 618 -7 0 net=2401
rlabel metal2 646 -9 646 -9 0 net=11601
rlabel metal2 709 -9 709 -9 0 net=12051
rlabel metal2 663 -11 663 -11 0 net=8953
rlabel metal2 716 -13 716 -13 0 net=9603
rlabel metal2 828 -13 828 -13 0 net=5141
rlabel metal2 730 -15 730 -15 0 net=11751
rlabel metal2 810 -15 810 -15 0 net=8899
rlabel metal2 835 -17 835 -17 0 net=6523
rlabel metal2 184 -28 184 -28 0 net=3945
rlabel metal2 240 -28 240 -28 0 net=11791
rlabel metal2 404 -28 404 -28 0 net=4111
rlabel metal2 492 -28 492 -28 0 net=2403
rlabel metal2 646 -28 646 -28 0 net=11603
rlabel metal2 737 -28 737 -28 0 net=10573
rlabel metal2 765 -28 765 -28 0 net=5143
rlabel metal2 842 -28 842 -28 0 net=11553
rlabel metal2 1234 -28 1234 -28 0 net=12687
rlabel metal2 1437 -28 1437 -28 0 net=13273
rlabel metal2 1629 -28 1629 -28 0 net=13617
rlabel metal2 198 -30 198 -30 0 net=5881
rlabel metal2 275 -30 275 -30 0 net=4651
rlabel metal2 317 -30 317 -30 0 net=6863
rlabel metal2 667 -30 667 -30 0 net=2867
rlabel metal2 744 -30 744 -30 0 net=4337
rlabel metal2 870 -30 870 -30 0 net=8900
rlabel metal2 908 -30 908 -30 0 net=9349
rlabel metal2 961 -30 961 -30 0 net=12943
rlabel metal2 1066 -30 1066 -30 0 net=6595
rlabel metal2 1108 -30 1108 -30 0 net=8171
rlabel metal2 1206 -30 1206 -30 0 net=9895
rlabel metal2 1321 -30 1321 -30 0 net=14131
rlabel metal2 1440 -30 1440 -30 0 net=14717
rlabel metal2 296 -32 296 -32 0 net=2967
rlabel metal2 355 -32 355 -32 0 net=3353
rlabel metal2 471 -32 471 -32 0 net=5577
rlabel metal2 618 -32 618 -32 0 net=6263
rlabel metal2 660 -32 660 -32 0 net=4097
rlabel metal2 702 -32 702 -32 0 net=7649
rlabel metal2 828 -32 828 -32 0 net=4923
rlabel metal2 1087 -32 1087 -32 0 net=11989
rlabel metal2 394 -34 394 -34 0 net=3147
rlabel metal2 499 -34 499 -34 0 net=1691
rlabel metal2 677 -34 677 -34 0 net=7361
rlabel metal2 978 -34 978 -34 0 net=13487
rlabel metal2 1010 -34 1010 -34 0 net=6983
rlabel metal2 1132 -34 1132 -34 0 net=13815
rlabel metal2 415 -36 415 -36 0 net=7259
rlabel metal2 432 -36 432 -36 0 net=6245
rlabel metal2 611 -36 611 -36 0 net=4709
rlabel metal2 702 -36 702 -36 0 net=9605
rlabel metal2 751 -36 751 -36 0 net=4883
rlabel metal2 912 -36 912 -36 0 net=9677
rlabel metal2 1073 -36 1073 -36 0 net=14097
rlabel metal2 1094 -36 1094 -36 0 net=4095
rlabel metal2 422 -38 422 -38 0 net=1681
rlabel metal2 485 -38 485 -38 0 net=2839
rlabel metal2 639 -38 639 -38 0 net=4449
rlabel metal2 716 -38 716 -38 0 net=7301
rlabel metal2 842 -38 842 -38 0 net=6379
rlabel metal2 926 -38 926 -38 0 net=7389
rlabel metal2 506 -40 506 -40 0 net=3653
rlabel metal2 856 -40 856 -40 0 net=8233
rlabel metal2 520 -42 520 -42 0 net=4033
rlabel metal2 583 -42 583 -42 0 net=11133
rlabel metal2 653 -42 653 -42 0 net=11809
rlabel metal2 982 -42 982 -42 0 net=9103
rlabel metal2 534 -44 534 -44 0 net=3725
rlabel metal2 768 -44 768 -44 0 net=9611
rlabel metal2 870 -44 870 -44 0 net=5935
rlabel metal2 982 -44 982 -44 0 net=7921
rlabel metal2 548 -46 548 -46 0 net=6199
rlabel metal2 604 -46 604 -46 0 net=3643
rlabel metal2 989 -46 989 -46 0 net=8955
rlabel metal2 548 -48 548 -48 0 net=3487
rlabel metal2 583 -48 583 -48 0 net=13059
rlabel metal2 1024 -48 1024 -48 0 net=14471
rlabel metal2 569 -50 569 -50 0 net=6637
rlabel metal2 793 -50 793 -50 0 net=6525
rlabel metal2 849 -50 849 -50 0 net=12619
rlabel metal2 569 -52 569 -52 0 net=1829
rlabel metal2 688 -52 688 -52 0 net=12053
rlabel metal2 772 -52 772 -52 0 net=8549
rlabel metal2 849 -52 849 -52 0 net=9569
rlabel metal2 709 -54 709 -54 0 net=11753
rlabel metal2 772 -54 772 -54 0 net=5587
rlabel metal2 877 -54 877 -54 0 net=9789
rlabel metal2 730 -56 730 -56 0 net=8685
rlabel metal2 800 -58 800 -58 0 net=11641
rlabel metal2 807 -60 807 -60 0 net=12635
rlabel metal2 887 -60 887 -60 0 net=8813
rlabel metal2 681 -62 681 -62 0 net=6875
rlabel metal2 891 -62 891 -62 0 net=13791
rlabel metal2 565 -64 565 -64 0 net=10689
rlabel metal2 803 -64 803 -64 0 net=12131
rlabel metal2 915 -64 915 -64 0 net=8363
rlabel metal2 58 -75 58 -75 0 net=5105
rlabel metal2 530 -75 530 -75 0 net=9743
rlabel metal2 1290 -75 1290 -75 0 net=9897
rlabel metal2 1332 -75 1332 -75 0 net=14133
rlabel metal2 1486 -75 1486 -75 0 net=13275
rlabel metal2 1633 -75 1633 -75 0 net=13619
rlabel metal2 1759 -75 1759 -75 0 net=14719
rlabel metal2 65 -77 65 -77 0 net=10195
rlabel metal2 233 -77 233 -77 0 net=9801
rlabel metal2 852 -77 852 -77 0 net=12869
rlabel metal2 1157 -77 1157 -77 0 net=10873
rlabel metal2 1171 -77 1171 -77 0 net=6283
rlabel metal2 1360 -77 1360 -77 0 net=12689
rlabel metal2 72 -79 72 -79 0 net=7489
rlabel metal2 404 -79 404 -79 0 net=3759
rlabel metal2 450 -79 450 -79 0 net=4035
rlabel metal2 555 -79 555 -79 0 net=4099
rlabel metal2 674 -79 674 -79 0 net=11754
rlabel metal2 740 -79 740 -79 0 net=14177
rlabel metal2 79 -81 79 -81 0 net=4825
rlabel metal2 359 -81 359 -81 0 net=1683
rlabel metal2 429 -81 429 -81 0 net=3645
rlabel metal2 625 -81 625 -81 0 net=4925
rlabel metal2 835 -81 835 -81 0 net=8551
rlabel metal2 919 -81 919 -81 0 net=11643
rlabel metal2 943 -81 943 -81 0 net=8665
rlabel metal2 1321 -81 1321 -81 0 net=13699
rlabel metal2 86 -83 86 -83 0 net=10547
rlabel metal2 282 -83 282 -83 0 net=1693
rlabel metal2 513 -83 513 -83 0 net=3309
rlabel metal2 562 -83 562 -83 0 net=6415
rlabel metal2 653 -83 653 -83 0 net=5145
rlabel metal2 786 -83 786 -83 0 net=7651
rlabel metal2 856 -83 856 -83 0 net=10983
rlabel metal2 1125 -83 1125 -83 0 net=13097
rlabel metal2 93 -85 93 -85 0 net=5579
rlabel metal2 478 -85 478 -85 0 net=4113
rlabel metal2 478 -85 478 -85 0 net=4113
rlabel metal2 499 -85 499 -85 0 net=4437
rlabel metal2 541 -85 541 -85 0 net=4711
rlabel metal2 660 -85 660 -85 0 net=4885
rlabel metal2 779 -85 779 -85 0 net=6639
rlabel metal2 856 -85 856 -85 0 net=6985
rlabel metal2 1031 -85 1031 -85 0 net=9105
rlabel metal2 1031 -85 1031 -85 0 net=9105
rlabel metal2 1038 -85 1038 -85 0 net=8235
rlabel metal2 1115 -85 1115 -85 0 net=8173
rlabel metal2 1178 -85 1178 -85 0 net=11991
rlabel metal2 100 -87 100 -87 0 net=7511
rlabel metal2 604 -87 604 -87 0 net=6265
rlabel metal2 702 -87 702 -87 0 net=9607
rlabel metal2 863 -87 863 -87 0 net=9613
rlabel metal2 919 -87 919 -87 0 net=8365
rlabel metal2 975 -87 975 -87 0 net=7363
rlabel metal2 107 -89 107 -89 0 net=3947
rlabel metal2 191 -89 191 -89 0 net=11793
rlabel metal2 247 -89 247 -89 0 net=4179
rlabel metal2 471 -89 471 -89 0 net=843
rlabel metal2 989 -89 989 -89 0 net=13793
rlabel metal2 1213 -89 1213 -89 0 net=13817
rlabel metal2 114 -91 114 -91 0 net=7183
rlabel metal2 240 -91 240 -91 0 net=4653
rlabel metal2 296 -91 296 -91 0 net=2969
rlabel metal2 338 -91 338 -91 0 net=7583
rlabel metal2 702 -91 702 -91 0 net=5937
rlabel metal2 898 -91 898 -91 0 net=10853
rlabel metal2 1220 -91 1220 -91 0 net=11555
rlabel metal2 124 -93 124 -93 0 net=4861
rlabel metal2 310 -93 310 -93 0 net=3117
rlabel metal2 345 -93 345 -93 0 net=2157
rlabel metal2 576 -93 576 -93 0 net=4451
rlabel metal2 709 -93 709 -93 0 net=7303
rlabel metal2 751 -93 751 -93 0 net=5067
rlabel metal2 1237 -93 1237 -93 0 net=13073
rlabel metal2 128 -95 128 -95 0 net=5303
rlabel metal2 590 -95 590 -95 0 net=6247
rlabel metal2 618 -95 618 -95 0 net=5133
rlabel metal2 961 -95 961 -95 0 net=11811
rlabel metal2 1227 -95 1227 -95 0 net=13857
rlabel metal2 135 -97 135 -97 0 net=3655
rlabel metal2 583 -97 583 -97 0 net=6201
rlabel metal2 639 -97 639 -97 0 net=3059
rlabel metal2 863 -97 863 -97 0 net=9791
rlabel metal2 954 -97 954 -97 0 net=9393
rlabel metal2 999 -97 999 -97 0 net=4096
rlabel metal2 1101 -97 1101 -97 0 net=6597
rlabel metal2 149 -99 149 -99 0 net=2527
rlabel metal2 366 -99 366 -99 0 net=1831
rlabel metal2 758 -99 758 -99 0 net=10575
rlabel metal2 933 -99 933 -99 0 net=13061
rlabel metal2 1118 -99 1118 -99 0 net=12949
rlabel metal2 152 -101 152 -101 0 net=1815
rlabel metal2 310 -101 310 -101 0 net=4577
rlabel metal2 870 -101 870 -101 0 net=7923
rlabel metal2 996 -101 996 -101 0 net=13577
rlabel metal2 156 -103 156 -103 0 net=6865
rlabel metal2 380 -103 380 -103 0 net=2405
rlabel metal2 730 -103 730 -103 0 net=8687
rlabel metal2 779 -103 779 -103 0 net=2889
rlabel metal2 912 -103 912 -103 0 net=9571
rlabel metal2 1003 -103 1003 -103 0 net=13489
rlabel metal2 163 -105 163 -105 0 net=3779
rlabel metal2 789 -105 789 -105 0 net=531
rlabel metal2 803 -105 803 -105 0 net=9931
rlabel metal2 968 -105 968 -105 0 net=9679
rlabel metal2 1027 -105 1027 -105 0 net=5087
rlabel metal2 170 -107 170 -107 0 net=3801
rlabel metal2 411 -107 411 -107 0 net=7260
rlabel metal2 422 -107 422 -107 0 net=3489
rlabel metal2 807 -107 807 -107 0 net=12637
rlabel metal2 1010 -107 1010 -107 0 net=4551
rlabel metal2 177 -109 177 -109 0 net=3727
rlabel metal2 548 -109 548 -109 0 net=4339
rlabel metal2 807 -109 807 -109 0 net=7391
rlabel metal2 933 -109 933 -109 0 net=14433
rlabel metal2 184 -111 184 -111 0 net=4169
rlabel metal2 744 -111 744 -111 0 net=6381
rlabel metal2 947 -111 947 -111 0 net=9351
rlabel metal2 1017 -111 1017 -111 0 net=8957
rlabel metal2 1073 -111 1073 -111 0 net=14473
rlabel metal2 198 -113 198 -113 0 net=5883
rlabel metal2 229 -113 229 -113 0 net=2503
rlabel metal2 373 -113 373 -113 0 net=5993
rlabel metal2 814 -113 814 -113 0 net=6877
rlabel metal2 912 -113 912 -113 0 net=10533
rlabel metal2 1024 -113 1024 -113 0 net=9169
rlabel metal2 1080 -113 1080 -113 0 net=12621
rlabel metal2 198 -115 198 -115 0 net=3819
rlabel metal2 492 -115 492 -115 0 net=4483
rlabel metal2 891 -115 891 -115 0 net=12133
rlabel metal2 1087 -115 1087 -115 0 net=14099
rlabel metal2 205 -117 205 -117 0 net=1991
rlabel metal2 534 -117 534 -117 0 net=5283
rlabel metal2 1087 -117 1087 -117 0 net=10615
rlabel metal2 212 -119 212 -119 0 net=2453
rlabel metal2 390 -119 390 -119 0 net=2069
rlabel metal2 597 -119 597 -119 0 net=13467
rlabel metal2 1038 -119 1038 -119 0 net=8729
rlabel metal2 261 -121 261 -121 0 net=984
rlabel metal2 681 -121 681 -121 0 net=10691
rlabel metal2 1045 -121 1045 -121 0 net=12945
rlabel metal2 275 -123 275 -123 0 net=3149
rlabel metal2 401 -123 401 -123 0 net=2841
rlabel metal2 646 -123 646 -123 0 net=11135
rlabel metal2 1052 -123 1052 -123 0 net=8815
rlabel metal2 296 -125 296 -125 0 net=3903
rlabel metal2 688 -125 688 -125 0 net=12055
rlabel metal2 142 -127 142 -127 0 net=7067
rlabel metal2 723 -127 723 -127 0 net=11605
rlabel metal2 394 -129 394 -129 0 net=3569
rlabel metal2 408 -131 408 -131 0 net=6467
rlabel metal2 723 -131 723 -131 0 net=6527
rlabel metal2 121 -133 121 -133 0 net=8889
rlabel metal2 415 -135 415 -135 0 net=3355
rlabel metal2 485 -135 485 -135 0 net=2869
rlabel metal2 446 -137 446 -137 0 net=3987
rlabel metal2 667 -137 667 -137 0 net=5589
rlabel metal2 457 -139 457 -139 0 net=2271
rlabel metal2 565 -139 565 -139 0 net=7975
rlabel metal2 772 -139 772 -139 0 net=9833
rlabel metal2 460 -141 460 -141 0 net=4687
rlabel metal2 16 -152 16 -152 0 net=7105
rlabel metal2 282 -152 282 -152 0 net=1695
rlabel metal2 408 -152 408 -152 0 net=6468
rlabel metal2 768 -152 768 -152 0 net=12419
rlabel metal2 1353 -152 1353 -152 0 net=11557
rlabel metal2 1374 -152 1374 -152 0 net=14135
rlabel metal2 1507 -152 1507 -152 0 net=13075
rlabel metal2 1640 -152 1640 -152 0 net=13621
rlabel metal2 1885 -152 1885 -152 0 net=14721
rlabel metal2 23 -154 23 -154 0 net=3949
rlabel metal2 114 -154 114 -154 0 net=7184
rlabel metal2 240 -154 240 -154 0 net=4654
rlabel metal2 282 -154 282 -154 0 net=2971
rlabel metal2 345 -154 345 -154 0 net=2158
rlabel metal2 541 -154 541 -154 0 net=4712
rlabel metal2 611 -154 611 -154 0 net=6248
rlabel metal2 803 -154 803 -154 0 net=11644
rlabel metal2 950 -154 950 -154 0 net=12923
rlabel metal2 1423 -154 1423 -154 0 net=12691
rlabel metal2 1514 -154 1514 -154 0 net=13277
rlabel metal2 1566 -154 1566 -154 0 net=9263
rlabel metal2 1615 -154 1615 -154 0 net=13759
rlabel metal2 37 -156 37 -156 0 net=9995
rlabel metal2 289 -156 289 -156 0 net=1817
rlabel metal2 289 -156 289 -156 0 net=1817
rlabel metal2 331 -156 331 -156 0 net=3357
rlabel metal2 422 -156 422 -156 0 net=3491
rlabel metal2 450 -156 450 -156 0 net=4036
rlabel metal2 541 -156 541 -156 0 net=4101
rlabel metal2 590 -156 590 -156 0 net=3989
rlabel metal2 684 -156 684 -156 0 net=7349
rlabel metal2 1013 -156 1013 -156 0 net=13515
rlabel metal2 1542 -156 1542 -156 0 net=9069
rlabel metal2 44 -158 44 -158 0 net=7491
rlabel metal2 86 -158 86 -158 0 net=10548
rlabel metal2 814 -158 814 -158 0 net=12057
rlabel metal2 1076 -158 1076 -158 0 net=10616
rlabel metal2 1276 -158 1276 -158 0 net=6599
rlabel metal2 51 -160 51 -160 0 net=4827
rlabel metal2 93 -160 93 -160 0 net=5581
rlabel metal2 649 -160 649 -160 0 net=12134
rlabel metal2 1090 -160 1090 -160 0 net=13881
rlabel metal2 72 -162 72 -162 0 net=1833
rlabel metal2 380 -162 380 -162 0 net=2407
rlabel metal2 429 -162 429 -162 0 net=3647
rlabel metal2 467 -162 467 -162 0 net=10692
rlabel metal2 1073 -162 1073 -162 0 net=10123
rlabel metal2 1283 -162 1283 -162 0 net=7365
rlabel metal2 79 -164 79 -164 0 net=3183
rlabel metal2 100 -164 100 -164 0 net=7512
rlabel metal2 128 -164 128 -164 0 net=5304
rlabel metal2 163 -164 163 -164 0 net=3781
rlabel metal2 240 -164 240 -164 0 net=13441
rlabel metal2 100 -166 100 -166 0 net=8683
rlabel metal2 618 -166 618 -166 0 net=5135
rlabel metal2 737 -166 737 -166 0 net=4553
rlabel metal2 1073 -166 1073 -166 0 net=8237
rlabel metal2 1129 -166 1129 -166 0 net=12947
rlabel metal2 107 -168 107 -168 0 net=2071
rlabel metal2 621 -168 621 -168 0 net=6887
rlabel metal2 814 -168 814 -168 0 net=4201
rlabel metal2 849 -168 849 -168 0 net=9802
rlabel metal2 975 -168 975 -168 0 net=11827
rlabel metal2 1290 -168 1290 -168 0 net=8667
rlabel metal2 117 -170 117 -170 0 net=6889
rlabel metal2 849 -170 849 -170 0 net=6879
rlabel metal2 884 -170 884 -170 0 net=9615
rlabel metal2 1122 -170 1122 -170 0 net=10985
rlabel metal2 1304 -170 1304 -170 0 net=13819
rlabel metal2 121 -172 121 -172 0 net=2947
rlabel metal2 226 -172 226 -172 0 net=4251
rlabel metal2 856 -172 856 -172 0 net=6987
rlabel metal2 887 -172 887 -172 0 net=4688
rlabel metal2 1311 -172 1311 -172 0 net=13859
rlabel metal2 128 -174 128 -174 0 net=8069
rlabel metal2 275 -174 275 -174 0 net=3151
rlabel metal2 450 -174 450 -174 0 net=4115
rlabel metal2 492 -174 492 -174 0 net=4485
rlabel metal2 667 -174 667 -174 0 net=5591
rlabel metal2 870 -174 870 -174 0 net=7925
rlabel metal2 1059 -174 1059 -174 0 net=9171
rlabel metal2 1136 -174 1136 -174 0 net=12871
rlabel metal2 65 -176 65 -176 0 net=10197
rlabel metal2 275 -176 275 -176 0 net=1685
rlabel metal2 366 -176 366 -176 0 net=4591
rlabel metal2 905 -176 905 -176 0 net=8553
rlabel metal2 989 -176 989 -176 0 net=9395
rlabel metal2 1150 -176 1150 -176 0 net=11813
rlabel metal2 1318 -176 1318 -176 0 net=13099
rlabel metal2 135 -178 135 -178 0 net=3657
rlabel metal2 338 -178 338 -178 0 net=7585
rlabel metal2 513 -178 513 -178 0 net=3311
rlabel metal2 569 -178 569 -178 0 net=6481
rlabel metal2 961 -178 961 -178 0 net=11865
rlabel metal2 1325 -178 1325 -178 0 net=14179
rlabel metal2 142 -180 142 -180 0 net=2455
rlabel metal2 243 -180 243 -180 0 net=616
rlabel metal2 296 -180 296 -180 0 net=3905
rlabel metal2 345 -180 345 -180 0 net=2871
rlabel metal2 513 -180 513 -180 0 net=3881
rlabel metal2 705 -180 705 -180 0 net=12301
rlabel metal2 1325 -180 1325 -180 0 net=8945
rlabel metal2 1360 -180 1360 -180 0 net=13701
rlabel metal2 145 -182 145 -182 0 net=6866
rlabel metal2 163 -182 163 -182 0 net=4987
rlabel metal2 401 -182 401 -182 0 net=2843
rlabel metal2 471 -182 471 -182 0 net=2623
rlabel metal2 1017 -182 1017 -182 0 net=8959
rlabel metal2 1164 -182 1164 -182 0 net=13491
rlabel metal2 149 -184 149 -184 0 net=7977
rlabel metal2 786 -184 786 -184 0 net=7653
rlabel metal2 919 -184 919 -184 0 net=8367
rlabel metal2 1080 -184 1080 -184 0 net=8175
rlabel metal2 1171 -184 1171 -184 0 net=12591
rlabel metal2 156 -186 156 -186 0 net=14497
rlabel metal2 170 -188 170 -188 0 net=3803
rlabel metal2 520 -188 520 -188 0 net=1156
rlabel metal2 1003 -188 1003 -188 0 net=12639
rlabel metal2 177 -190 177 -190 0 net=3729
rlabel metal2 373 -190 373 -190 0 net=5995
rlabel metal2 709 -190 709 -190 0 net=7305
rlabel metal2 912 -190 912 -190 0 net=10535
rlabel metal2 954 -190 954 -190 0 net=9933
rlabel metal2 1171 -190 1171 -190 0 net=10063
rlabel metal2 177 -192 177 -192 0 net=3761
rlabel metal2 520 -192 520 -192 0 net=9165
rlabel metal2 968 -192 968 -192 0 net=9681
rlabel metal2 1174 -192 1174 -192 0 net=9744
rlabel metal2 58 -194 58 -194 0 net=5106
rlabel metal2 527 -194 527 -194 0 net=11606
rlabel metal2 1094 -194 1094 -194 0 net=13579
rlabel metal2 58 -196 58 -196 0 net=4629
rlabel metal2 184 -196 184 -196 0 net=4170
rlabel metal2 310 -196 310 -196 0 net=4579
rlabel metal2 506 -196 506 -196 0 net=2273
rlabel metal2 534 -196 534 -196 0 net=5285
rlabel metal2 758 -196 758 -196 0 net=8689
rlabel metal2 793 -196 793 -196 0 net=8891
rlabel metal2 1017 -196 1017 -196 0 net=9221
rlabel metal2 1178 -196 1178 -196 0 net=12623
rlabel metal2 170 -198 170 -198 0 net=3893
rlabel metal2 317 -198 317 -198 0 net=2505
rlabel metal2 394 -198 394 -198 0 net=3571
rlabel metal2 555 -198 555 -198 0 net=2891
rlabel metal2 821 -198 821 -198 0 net=6641
rlabel metal2 1038 -198 1038 -198 0 net=8731
rlabel metal2 1094 -198 1094 -198 0 net=12211
rlabel metal2 1185 -198 1185 -198 0 net=12951
rlabel metal2 184 -200 184 -200 0 net=3751
rlabel metal2 674 -200 674 -200 0 net=8311
rlabel metal2 1038 -200 1038 -200 0 net=9337
rlabel metal2 194 -202 194 -202 0 net=10919
rlabel metal2 1101 -202 1101 -202 0 net=13063
rlabel metal2 198 -204 198 -204 0 net=3821
rlabel metal2 660 -204 660 -204 0 net=4887
rlabel metal2 688 -204 688 -204 0 net=7069
rlabel metal2 1066 -204 1066 -204 0 net=8817
rlabel metal2 1143 -204 1143 -204 0 net=6285
rlabel metal2 30 -206 30 -206 0 net=12453
rlabel metal2 212 -206 212 -206 0 net=10137
rlabel metal2 898 -206 898 -206 0 net=10577
rlabel metal2 1192 -206 1192 -206 0 net=13795
rlabel metal2 219 -208 219 -208 0 net=5885
rlabel metal2 324 -208 324 -208 0 net=3119
rlabel metal2 401 -208 401 -208 0 net=3061
rlabel metal2 698 -208 698 -208 0 net=9911
rlabel metal2 1199 -208 1199 -208 0 net=14435
rlabel metal2 219 -210 219 -210 0 net=4439
rlabel metal2 548 -210 548 -210 0 net=4341
rlabel metal2 709 -210 709 -210 0 net=5088
rlabel metal2 1241 -210 1241 -210 0 net=9899
rlabel metal2 247 -212 247 -212 0 net=4180
rlabel metal2 1031 -212 1031 -212 0 net=9107
rlabel metal2 1157 -212 1157 -212 0 net=10875
rlabel metal2 1255 -212 1255 -212 0 net=11993
rlabel metal2 89 -214 89 -214 0 net=5085
rlabel metal2 324 -214 324 -214 0 net=2359
rlabel metal2 1269 -214 1269 -214 0 net=6503
rlabel metal2 352 -216 352 -216 0 net=2529
rlabel metal2 499 -216 499 -216 0 net=5069
rlabel metal2 758 -216 758 -216 0 net=7151
rlabel metal2 1199 -216 1199 -216 0 net=11309
rlabel metal2 352 -218 352 -218 0 net=4161
rlabel metal2 548 -218 548 -218 0 net=5567
rlabel metal2 996 -218 996 -218 0 net=9353
rlabel metal2 1202 -218 1202 -218 0 net=12343
rlabel metal2 523 -220 523 -220 0 net=11136
rlabel metal2 863 -220 863 -220 0 net=9793
rlabel metal2 1045 -220 1045 -220 0 net=9835
rlabel metal2 1206 -220 1206 -220 0 net=14101
rlabel metal2 583 -222 583 -222 0 net=6203
rlabel metal2 765 -222 765 -222 0 net=7327
rlabel metal2 1213 -222 1213 -222 0 net=10855
rlabel metal2 576 -224 576 -224 0 net=4453
rlabel metal2 604 -224 604 -224 0 net=6267
rlabel metal2 702 -224 702 -224 0 net=5939
rlabel metal2 891 -224 891 -224 0 net=13469
rlabel metal2 303 -226 303 -226 0 net=4863
rlabel metal2 632 -226 632 -226 0 net=6417
rlabel metal2 982 -226 982 -226 0 net=9573
rlabel metal2 1216 -226 1216 -226 0 net=12335
rlabel metal2 205 -228 205 -228 0 net=1993
rlabel metal2 576 -228 576 -228 0 net=7021
rlabel metal2 744 -228 744 -228 0 net=6383
rlabel metal2 807 -228 807 -228 0 net=7393
rlabel metal2 936 -228 936 -228 0 net=8693
rlabel metal2 1003 -228 1003 -228 0 net=5641
rlabel metal2 1220 -228 1220 -228 0 net=14475
rlabel metal2 439 -230 439 -230 0 net=11607
rlabel metal2 1255 -230 1255 -230 0 net=8499
rlabel metal2 625 -232 625 -232 0 net=4927
rlabel metal2 639 -232 639 -232 0 net=4705
rlabel metal2 779 -232 779 -232 0 net=7721
rlabel metal2 191 -234 191 -234 0 net=11795
rlabel metal2 653 -234 653 -234 0 net=5147
rlabel metal2 807 -234 807 -234 0 net=7751
rlabel metal2 135 -236 135 -236 0 net=6323
rlabel metal2 835 -236 835 -236 0 net=10971
rlabel metal2 800 -238 800 -238 0 net=6919
rlabel metal2 800 -240 800 -240 0 net=9609
rlabel metal2 723 -242 723 -242 0 net=6529
rlabel metal2 534 -244 534 -244 0 net=6429
rlabel metal2 16 -255 16 -255 0 net=7106
rlabel metal2 198 -255 198 -255 0 net=3907
rlabel metal2 366 -255 366 -255 0 net=4592
rlabel metal2 761 -255 761 -255 0 net=1008
rlabel metal2 992 -255 992 -255 0 net=12559
rlabel metal2 1612 -255 1612 -255 0 net=3741
rlabel metal2 16 -257 16 -257 0 net=7979
rlabel metal2 156 -257 156 -257 0 net=1499
rlabel metal2 618 -257 618 -257 0 net=9610
rlabel metal2 810 -257 810 -257 0 net=14303
rlabel metal2 1815 -257 1815 -257 0 net=9071
rlabel metal2 1941 -257 1941 -257 0 net=14723
rlabel metal2 44 -259 44 -259 0 net=7492
rlabel metal2 240 -259 240 -259 0 net=1304
rlabel metal2 338 -259 338 -259 0 net=2409
rlabel metal2 432 -259 432 -259 0 net=981
rlabel metal2 828 -259 828 -259 0 net=6530
rlabel metal2 880 -259 880 -259 0 net=13796
rlabel metal2 1542 -259 1542 -259 0 net=12567
rlabel metal2 1615 -259 1615 -259 0 net=12885
rlabel metal2 1668 -259 1668 -259 0 net=13623
rlabel metal2 1962 -259 1962 -259 0 net=12541
rlabel metal2 23 -261 23 -261 0 net=3950
rlabel metal2 247 -261 247 -261 0 net=5086
rlabel metal2 439 -261 439 -261 0 net=648
rlabel metal2 653 -261 653 -261 0 net=6325
rlabel metal2 891 -261 891 -261 0 net=12787
rlabel metal2 23 -263 23 -263 0 net=9997
rlabel metal2 54 -263 54 -263 0 net=13442
rlabel metal2 1514 -263 1514 -263 0 net=14499
rlabel metal2 37 -265 37 -265 0 net=2845
rlabel metal2 422 -265 422 -265 0 net=3823
rlabel metal2 709 -265 709 -265 0 net=9794
rlabel metal2 1083 -265 1083 -265 0 net=12989
rlabel metal2 65 -267 65 -267 0 net=8071
rlabel metal2 149 -267 149 -267 0 net=3895
rlabel metal2 187 -267 187 -267 0 net=10198
rlabel metal2 268 -267 268 -267 0 net=1994
rlabel metal2 310 -267 310 -267 0 net=8694
rlabel metal2 996 -267 996 -267 0 net=14347
rlabel metal2 86 -269 86 -269 0 net=3185
rlabel metal2 114 -269 114 -269 0 net=2457
rlabel metal2 156 -269 156 -269 0 net=4929
rlabel metal2 709 -269 709 -269 0 net=4203
rlabel metal2 828 -269 828 -269 0 net=6881
rlabel metal2 856 -269 856 -269 0 net=7307
rlabel metal2 1010 -269 1010 -269 0 net=13797
rlabel metal2 58 -271 58 -271 0 net=4631
rlabel metal2 233 -271 233 -271 0 net=3783
rlabel metal2 422 -271 422 -271 0 net=3649
rlabel metal2 506 -271 506 -271 0 net=3573
rlabel metal2 534 -271 534 -271 0 net=12058
rlabel metal2 954 -271 954 -271 0 net=7071
rlabel metal2 1094 -271 1094 -271 0 net=12213
rlabel metal2 1552 -271 1552 -271 0 net=13507
rlabel metal2 58 -273 58 -273 0 net=5149
rlabel metal2 772 -273 772 -273 0 net=5593
rlabel metal2 856 -273 856 -273 0 net=8187
rlabel metal2 1010 -273 1010 -273 0 net=9223
rlabel metal2 1020 -273 1020 -273 0 net=12948
rlabel metal2 1465 -273 1465 -273 0 net=13883
rlabel metal2 93 -275 93 -275 0 net=8684
rlabel metal2 128 -275 128 -275 0 net=3659
rlabel metal2 268 -275 268 -275 0 net=2625
rlabel metal2 506 -275 506 -275 0 net=7723
rlabel metal2 863 -275 863 -275 0 net=5941
rlabel metal2 954 -275 954 -275 0 net=5643
rlabel metal2 1101 -275 1101 -275 0 net=8819
rlabel metal2 1227 -275 1227 -275 0 net=12303
rlabel metal2 100 -277 100 -277 0 net=3763
rlabel metal2 205 -277 205 -277 0 net=7269
rlabel metal2 842 -277 842 -277 0 net=6419
rlabel metal2 894 -277 894 -277 0 net=14476
rlabel metal2 1556 -277 1556 -277 0 net=13279
rlabel metal2 72 -279 72 -279 0 net=1835
rlabel metal2 191 -279 191 -279 0 net=5931
rlabel metal2 219 -279 219 -279 0 net=4441
rlabel metal2 555 -279 555 -279 0 net=2893
rlabel metal2 628 -279 628 -279 0 net=7735
rlabel metal2 1153 -279 1153 -279 0 net=13151
rlabel metal2 72 -281 72 -281 0 net=6921
rlabel metal2 926 -281 926 -281 0 net=7351
rlabel metal2 1178 -281 1178 -281 0 net=11849
rlabel metal2 1591 -281 1591 -281 0 net=14181
rlabel metal2 107 -283 107 -283 0 net=2073
rlabel metal2 275 -283 275 -283 0 net=1686
rlabel metal2 471 -283 471 -283 0 net=4581
rlabel metal2 513 -283 513 -283 0 net=3883
rlabel metal2 667 -283 667 -283 0 net=5997
rlabel metal2 947 -283 947 -283 0 net=9167
rlabel metal2 1262 -283 1262 -283 0 net=13471
rlabel metal2 107 -285 107 -285 0 net=3157
rlabel metal2 219 -285 219 -285 0 net=4253
rlabel metal2 233 -285 233 -285 0 net=5871
rlabel metal2 947 -285 947 -285 0 net=6855
rlabel metal2 1626 -285 1626 -285 0 net=13077
rlabel metal2 135 -287 135 -287 0 net=3195
rlabel metal2 310 -287 310 -287 0 net=4117
rlabel metal2 548 -287 548 -287 0 net=5569
rlabel metal2 569 -287 569 -287 0 net=6483
rlabel metal2 968 -287 968 -287 0 net=8313
rlabel metal2 1213 -287 1213 -287 0 net=12659
rlabel metal2 1633 -287 1633 -287 0 net=13761
rlabel metal2 30 -289 30 -289 0 net=12455
rlabel metal2 548 -289 548 -289 0 net=3427
rlabel metal2 1122 -289 1122 -289 0 net=8961
rlabel metal2 1276 -289 1276 -289 0 net=11829
rlabel metal2 30 -291 30 -291 0 net=4829
rlabel metal2 138 -291 138 -291 0 net=11547
rlabel metal2 226 -291 226 -291 0 net=4163
rlabel metal2 394 -291 394 -291 0 net=3121
rlabel metal2 611 -291 611 -291 0 net=6891
rlabel metal2 975 -291 975 -291 0 net=8555
rlabel metal2 1136 -291 1136 -291 0 net=9397
rlabel metal2 1297 -291 1297 -291 0 net=11995
rlabel metal2 47 -293 47 -293 0 net=1136
rlabel metal2 138 -293 138 -293 0 net=1935
rlabel metal2 394 -293 394 -293 0 net=2149
rlabel metal2 611 -293 611 -293 0 net=3991
rlabel metal2 702 -293 702 -293 0 net=9471
rlabel metal2 1318 -293 1318 -293 0 net=12337
rlabel metal2 89 -295 89 -295 0 net=6821
rlabel metal2 688 -295 688 -295 0 net=6269
rlabel metal2 723 -295 723 -295 0 net=6431
rlabel metal2 919 -295 919 -295 0 net=10537
rlabel metal2 1328 -295 1328 -295 0 net=14033
rlabel metal2 243 -297 243 -297 0 net=4875
rlabel metal2 429 -297 429 -297 0 net=3153
rlabel metal2 576 -297 576 -297 0 net=7023
rlabel metal2 1108 -297 1108 -297 0 net=9617
rlabel metal2 1353 -297 1353 -297 0 net=12625
rlabel metal2 247 -299 247 -299 0 net=1599
rlabel metal2 576 -299 576 -299 0 net=3077
rlabel metal2 1024 -299 1024 -299 0 net=7927
rlabel metal2 1360 -299 1360 -299 0 net=12641
rlabel metal2 254 -301 254 -301 0 net=2347
rlabel metal2 275 -301 275 -301 0 net=2361
rlabel metal2 345 -301 345 -301 0 net=2873
rlabel metal2 597 -301 597 -301 0 net=4487
rlabel metal2 723 -301 723 -301 0 net=7153
rlabel metal2 772 -301 772 -301 0 net=12555
rlabel metal2 282 -303 282 -303 0 net=2973
rlabel metal2 660 -303 660 -303 0 net=4343
rlabel metal2 730 -303 730 -303 0 net=6888
rlabel metal2 1171 -303 1171 -303 0 net=10065
rlabel metal2 1374 -303 1374 -303 0 net=8669
rlabel metal2 135 -305 135 -305 0 net=1707
rlabel metal2 289 -305 289 -305 0 net=1819
rlabel metal2 660 -305 660 -305 0 net=4069
rlabel metal2 1381 -305 1381 -305 0 net=11311
rlabel metal2 1472 -305 1472 -305 0 net=13861
rlabel metal2 289 -307 289 -307 0 net=1697
rlabel metal2 401 -307 401 -307 0 net=3063
rlabel metal2 716 -307 716 -307 0 net=5287
rlabel metal2 786 -307 786 -307 0 net=8691
rlabel metal2 1185 -307 1185 -307 0 net=10579
rlabel metal2 1388 -307 1388 -307 0 net=12593
rlabel metal2 296 -309 296 -309 0 net=5071
rlabel metal2 646 -309 646 -309 0 net=5583
rlabel metal2 786 -309 786 -309 0 net=1611
rlabel metal2 1073 -309 1073 -309 0 net=8239
rlabel metal2 1185 -309 1185 -309 0 net=8947
rlabel metal2 1395 -309 1395 -309 0 net=12873
rlabel metal2 212 -311 212 -311 0 net=5673
rlabel metal2 1073 -311 1073 -311 0 net=6504
rlabel metal2 1402 -311 1402 -311 0 net=12925
rlabel metal2 299 -313 299 -313 0 net=7752
rlabel metal2 1076 -313 1076 -313 0 net=10885
rlabel metal2 1409 -313 1409 -313 0 net=12953
rlabel metal2 324 -315 324 -315 0 net=4103
rlabel metal2 1157 -315 1157 -315 0 net=9837
rlabel metal2 1311 -315 1311 -315 0 net=10857
rlabel metal2 1416 -315 1416 -315 0 net=13065
rlabel metal2 331 -317 331 -317 0 net=3359
rlabel metal2 933 -317 933 -317 0 net=10921
rlabel metal2 1423 -317 1423 -317 0 net=13493
rlabel metal2 331 -319 331 -319 0 net=2639
rlabel metal2 870 -319 870 -319 0 net=6643
rlabel metal2 1104 -319 1104 -319 0 net=9701
rlabel metal2 1430 -319 1430 -319 0 net=13517
rlabel metal2 345 -321 345 -321 0 net=2275
rlabel metal2 632 -321 632 -321 0 net=8489
rlabel metal2 1157 -321 1157 -321 0 net=8501
rlabel metal2 1437 -321 1437 -321 0 net=13101
rlabel metal2 79 -323 79 -323 0 net=3579
rlabel metal2 712 -323 712 -323 0 net=10223
rlabel metal2 1444 -323 1444 -323 0 net=13821
rlabel metal2 79 -325 79 -325 0 net=4989
rlabel metal2 352 -325 352 -325 0 net=5209
rlabel metal2 1164 -325 1164 -325 0 net=9935
rlabel metal2 1451 -325 1451 -325 0 net=11437
rlabel metal2 163 -327 163 -327 0 net=342
rlabel metal2 359 -327 359 -327 0 net=3731
rlabel metal2 1017 -327 1017 -327 0 net=10915
rlabel metal2 1192 -327 1192 -327 0 net=9913
rlabel metal2 1472 -327 1472 -327 0 net=9265
rlabel metal2 359 -329 359 -329 0 net=2139
rlabel metal2 1066 -329 1066 -329 0 net=9109
rlabel metal2 1206 -329 1206 -329 0 net=10973
rlabel metal2 1486 -329 1486 -329 0 net=14437
rlabel metal2 117 -331 117 -331 0 net=8133
rlabel metal2 1087 -331 1087 -331 0 net=9355
rlabel metal2 1220 -331 1220 -331 0 net=11609
rlabel metal2 1493 -331 1493 -331 0 net=12693
rlabel metal2 380 -333 380 -333 0 net=2531
rlabel metal2 443 -333 443 -333 0 net=3493
rlabel metal2 961 -333 961 -333 0 net=8893
rlabel metal2 1234 -333 1234 -333 0 net=10877
rlabel metal2 1500 -333 1500 -333 0 net=14137
rlabel metal2 373 -335 373 -335 0 net=2507
rlabel metal2 443 -335 443 -335 0 net=7586
rlabel metal2 765 -335 765 -335 0 net=7329
rlabel metal2 1038 -335 1038 -335 0 net=9339
rlabel metal2 1248 -335 1248 -335 0 net=10125
rlabel metal2 1479 -335 1479 -335 0 net=14103
rlabel metal2 1563 -335 1563 -335 0 net=12497
rlabel metal2 373 -337 373 -337 0 net=5773
rlabel metal2 1038 -337 1038 -337 0 net=6721
rlabel metal2 1248 -337 1248 -337 0 net=7367
rlabel metal2 478 -339 478 -339 0 net=12095
rlabel metal2 639 -341 639 -341 0 net=4707
rlabel metal2 1129 -341 1129 -341 0 net=9173
rlabel metal2 1283 -341 1283 -341 0 net=11815
rlabel metal2 639 -343 639 -343 0 net=5137
rlabel metal2 1045 -343 1045 -343 0 net=9575
rlabel metal2 1290 -343 1290 -343 0 net=10987
rlabel metal2 695 -345 695 -345 0 net=4555
rlabel metal2 877 -345 877 -345 0 net=6989
rlabel metal2 1052 -345 1052 -345 0 net=8733
rlabel metal2 1150 -345 1150 -345 0 net=6601
rlabel metal2 604 -347 604 -347 0 net=4865
rlabel metal2 877 -347 877 -347 0 net=10695
rlabel metal2 1458 -347 1458 -347 0 net=13703
rlabel metal2 317 -349 317 -349 0 net=5887
rlabel metal2 625 -349 625 -349 0 net=11797
rlabel metal2 121 -351 121 -351 0 net=2949
rlabel metal2 401 -351 401 -351 0 net=411
rlabel metal2 898 -351 898 -351 0 net=7395
rlabel metal2 1304 -351 1304 -351 0 net=11867
rlabel metal2 121 -353 121 -353 0 net=4455
rlabel metal2 898 -353 898 -353 0 net=6287
rlabel metal2 1339 -353 1339 -353 0 net=12345
rlabel metal2 492 -355 492 -355 0 net=3805
rlabel metal2 1024 -355 1024 -355 0 net=9657
rlabel metal2 1346 -355 1346 -355 0 net=12421
rlabel metal2 492 -357 492 -357 0 net=3313
rlabel metal2 821 -357 821 -357 0 net=10139
rlabel metal2 1367 -357 1367 -357 0 net=11559
rlabel metal2 184 -359 184 -359 0 net=3753
rlabel metal2 751 -359 751 -359 0 net=6205
rlabel metal2 1059 -359 1059 -359 0 net=8369
rlabel metal2 1181 -359 1181 -359 0 net=10659
rlabel metal2 674 -361 674 -361 0 net=4889
rlabel metal2 905 -361 905 -361 0 net=7655
rlabel metal2 1115 -361 1115 -361 0 net=9683
rlabel metal2 467 -363 467 -363 0 net=4771
rlabel metal2 793 -363 793 -363 0 net=6385
rlabel metal2 1080 -363 1080 -363 0 net=8177
rlabel metal2 1241 -363 1241 -363 0 net=9901
rlabel metal2 793 -365 793 -365 0 net=13580
rlabel metal2 835 -367 835 -367 0 net=11889
rlabel metal2 887 -369 887 -369 0 net=11001
rlabel metal2 16 -380 16 -380 0 net=7980
rlabel metal2 625 -380 625 -380 0 net=6270
rlabel metal2 758 -380 758 -380 0 net=9618
rlabel metal2 1353 -380 1353 -380 0 net=14453
rlabel metal2 1958 -380 1958 -380 0 net=13695
rlabel metal2 2193 -380 2193 -380 0 net=12543
rlabel metal2 23 -382 23 -382 0 net=9998
rlabel metal2 751 -382 751 -382 0 net=4891
rlabel metal2 761 -382 761 -382 0 net=5523
rlabel metal2 810 -382 810 -382 0 net=6882
rlabel metal2 845 -382 845 -382 0 net=13472
rlabel metal2 1766 -382 1766 -382 0 net=13508
rlabel metal2 1969 -382 1969 -382 0 net=3743
rlabel metal2 23 -384 23 -384 0 net=8421
rlabel metal2 51 -384 51 -384 0 net=4991
rlabel metal2 96 -384 96 -384 0 net=1200
rlabel metal2 1185 -384 1185 -384 0 net=8949
rlabel metal2 1353 -384 1353 -384 0 net=9267
rlabel metal2 1528 -384 1528 -384 0 net=11997
rlabel metal2 1528 -384 1528 -384 0 net=11997
rlabel metal2 1591 -384 1591 -384 0 net=12557
rlabel metal2 1773 -384 1773 -384 0 net=13823
rlabel metal2 1927 -384 1927 -384 0 net=9073
rlabel metal2 2004 -384 2004 -384 0 net=14035
rlabel metal2 37 -386 37 -386 0 net=2846
rlabel metal2 495 -386 495 -386 0 net=3754
rlabel metal2 600 -386 600 -386 0 net=8692
rlabel metal2 1167 -386 1167 -386 0 net=12874
rlabel metal2 1710 -386 1710 -386 0 net=13153
rlabel metal2 1976 -386 1976 -386 0 net=12539
rlabel metal2 2011 -386 2011 -386 0 net=14777
rlabel metal2 44 -388 44 -388 0 net=2479
rlabel metal2 478 -388 478 -388 0 net=8188
rlabel metal2 971 -388 971 -388 0 net=13494
rlabel metal2 1794 -388 1794 -388 0 net=13885
rlabel metal2 1983 -388 1983 -388 0 net=14725
rlabel metal2 61 -390 61 -390 0 net=1600
rlabel metal2 345 -390 345 -390 0 net=2277
rlabel metal2 499 -390 499 -390 0 net=3361
rlabel metal2 499 -390 499 -390 0 net=3361
rlabel metal2 513 -390 513 -390 0 net=3065
rlabel metal2 625 -390 625 -390 0 net=6327
rlabel metal2 978 -390 978 -390 0 net=10140
rlabel metal2 1356 -390 1356 -390 0 net=11610
rlabel metal2 1440 -390 1440 -390 0 net=14647
rlabel metal2 65 -392 65 -392 0 net=8073
rlabel metal2 65 -392 65 -392 0 net=8073
rlabel metal2 72 -392 72 -392 0 net=6923
rlabel metal2 163 -392 163 -392 0 net=14304
rlabel metal2 1808 -392 1808 -392 0 net=14139
rlabel metal2 16 -394 16 -394 0 net=5309
rlabel metal2 170 -394 170 -394 0 net=11548
rlabel metal2 222 -394 222 -394 0 net=3824
rlabel metal2 635 -394 635 -394 0 net=11645
rlabel metal2 1612 -394 1612 -394 0 net=14305
rlabel metal2 72 -396 72 -396 0 net=3187
rlabel metal2 173 -396 173 -396 0 net=5932
rlabel metal2 233 -396 233 -396 0 net=5873
rlabel metal2 765 -396 765 -396 0 net=4708
rlabel metal2 978 -396 978 -396 0 net=8894
rlabel metal2 1125 -396 1125 -396 0 net=13189
rlabel metal2 30 -398 30 -398 0 net=4830
rlabel metal2 247 -398 247 -398 0 net=5775
rlabel metal2 401 -398 401 -398 0 net=7724
rlabel metal2 513 -398 513 -398 0 net=4489
rlabel metal2 702 -398 702 -398 0 net=6351
rlabel metal2 1017 -398 1017 -398 0 net=13798
rlabel metal2 1815 -398 1815 -398 0 net=14183
rlabel metal2 79 -400 79 -400 0 net=3993
rlabel metal2 646 -400 646 -400 0 net=6433
rlabel metal2 982 -400 982 -400 0 net=8314
rlabel metal2 1136 -400 1136 -400 0 net=7369
rlabel metal2 1262 -400 1262 -400 0 net=9473
rlabel metal2 1360 -400 1360 -400 0 net=10067
rlabel metal2 1493 -400 1493 -400 0 net=11817
rlabel metal2 1633 -400 1633 -400 0 net=12695
rlabel metal2 1787 -400 1787 -400 0 net=13863
rlabel metal2 1836 -400 1836 -400 0 net=14439
rlabel metal2 86 -402 86 -402 0 net=4877
rlabel metal2 443 -402 443 -402 0 net=5207
rlabel metal2 527 -402 527 -402 0 net=3580
rlabel metal2 1020 -402 1020 -402 0 net=10927
rlabel metal2 1360 -402 1360 -402 0 net=12097
rlabel metal2 1549 -402 1549 -402 0 net=12215
rlabel metal2 1654 -402 1654 -402 0 net=13281
rlabel metal2 121 -404 121 -404 0 net=4457
rlabel metal2 212 -404 212 -404 0 net=5675
rlabel metal2 527 -404 527 -404 0 net=3429
rlabel metal2 667 -404 667 -404 0 net=4344
rlabel metal2 793 -404 793 -404 0 net=12642
rlabel metal2 1745 -404 1745 -404 0 net=13763
rlabel metal2 114 -406 114 -406 0 net=2459
rlabel metal2 156 -406 156 -406 0 net=4931
rlabel metal2 849 -406 849 -406 0 net=5999
rlabel metal2 1024 -406 1024 -406 0 net=12755
rlabel metal2 1843 -406 1843 -406 0 net=14501
rlabel metal2 156 -408 156 -408 0 net=9321
rlabel metal2 219 -408 219 -408 0 net=4255
rlabel metal2 674 -408 674 -408 0 net=4773
rlabel metal2 852 -408 852 -408 0 net=8556
rlabel metal2 1129 -408 1129 -408 0 net=8735
rlabel metal2 1388 -408 1388 -408 0 net=9915
rlabel metal2 1500 -408 1500 -408 0 net=14105
rlabel metal2 149 -410 149 -410 0 net=3897
rlabel metal2 226 -410 226 -410 0 net=4165
rlabel metal2 674 -410 674 -410 0 net=4205
rlabel metal2 716 -410 716 -410 0 net=5585
rlabel metal2 856 -410 856 -410 0 net=5813
rlabel metal2 1027 -410 1027 -410 0 net=14477
rlabel metal2 149 -412 149 -412 0 net=2885
rlabel metal2 541 -412 541 -412 0 net=3495
rlabel metal2 653 -412 653 -412 0 net=3885
rlabel metal2 730 -412 730 -412 0 net=5289
rlabel metal2 863 -412 863 -412 0 net=6420
rlabel metal2 1031 -412 1031 -412 0 net=7073
rlabel metal2 1164 -412 1164 -412 0 net=10917
rlabel metal2 1563 -412 1563 -412 0 net=12347
rlabel metal2 1661 -412 1661 -412 0 net=12887
rlabel metal2 187 -414 187 -414 0 net=12649
rlabel metal2 226 -416 226 -416 0 net=3817
rlabel metal2 345 -416 345 -416 0 net=3155
rlabel metal2 541 -416 541 -416 0 net=2327
rlabel metal2 653 -416 653 -416 0 net=11868
rlabel metal2 1507 -416 1507 -416 0 net=11831
rlabel metal2 1570 -416 1570 -416 0 net=13705
rlabel metal2 240 -418 240 -418 0 net=2627
rlabel metal2 359 -418 359 -418 0 net=2140
rlabel metal2 548 -418 548 -418 0 net=2875
rlabel metal2 681 -418 681 -418 0 net=6823
rlabel metal2 1059 -418 1059 -418 0 net=7657
rlabel metal2 1178 -418 1178 -418 0 net=9659
rlabel metal2 1311 -418 1311 -418 0 net=9703
rlabel metal2 1402 -418 1402 -418 0 net=10859
rlabel metal2 1584 -418 1584 -418 0 net=12499
rlabel metal2 1724 -418 1724 -418 0 net=13519
rlabel metal2 166 -420 166 -420 0 net=1977
rlabel metal2 373 -420 373 -420 0 net=2975
rlabel metal2 471 -420 471 -420 0 net=4583
rlabel metal2 688 -420 688 -420 0 net=4345
rlabel metal2 968 -420 968 -420 0 net=6893
rlabel metal2 1073 -420 1073 -420 0 net=13499
rlabel metal2 100 -422 100 -422 0 net=3765
rlabel metal2 457 -422 457 -422 0 net=3123
rlabel metal2 730 -422 730 -422 0 net=4537
rlabel metal2 1076 -422 1076 -422 0 net=12304
rlabel metal2 1668 -422 1668 -422 0 net=12927
rlabel metal2 100 -424 100 -424 0 net=3575
rlabel metal2 744 -424 744 -424 0 net=9307
rlabel metal2 1328 -424 1328 -424 0 net=12235
rlabel metal2 1675 -424 1675 -424 0 net=12955
rlabel metal2 166 -426 166 -426 0 net=2640
rlabel metal2 401 -426 401 -426 0 net=1821
rlabel metal2 737 -426 737 -426 0 net=4867
rlabel metal2 779 -426 779 -426 0 net=7271
rlabel metal2 1080 -426 1080 -426 0 net=9168
rlabel metal2 1332 -426 1332 -426 0 net=9937
rlabel metal2 1409 -426 1409 -426 0 net=10879
rlabel metal2 1556 -426 1556 -426 0 net=12339
rlabel metal2 1682 -426 1682 -426 0 net=14349
rlabel metal2 212 -428 212 -428 0 net=7213
rlabel metal2 1083 -428 1083 -428 0 net=12185
rlabel metal2 1689 -428 1689 -428 0 net=12991
rlabel metal2 268 -430 268 -430 0 net=6387
rlabel metal2 968 -430 968 -430 0 net=12217
rlabel metal2 1703 -430 1703 -430 0 net=13103
rlabel metal2 296 -432 296 -432 0 net=5073
rlabel metal2 803 -432 803 -432 0 net=6391
rlabel metal2 1367 -432 1367 -432 0 net=10661
rlabel metal2 1486 -432 1486 -432 0 net=11561
rlabel metal2 1619 -432 1619 -432 0 net=12595
rlabel metal2 296 -434 296 -434 0 net=1613
rlabel metal2 807 -434 807 -434 0 net=5093
rlabel metal2 1192 -434 1192 -434 0 net=9111
rlabel metal2 1437 -434 1437 -434 0 net=10127
rlabel metal2 1514 -434 1514 -434 0 net=11851
rlabel metal2 1626 -434 1626 -434 0 net=12627
rlabel metal2 303 -436 303 -436 0 net=3197
rlabel metal2 632 -436 632 -436 0 net=5247
rlabel metal2 842 -436 842 -436 0 net=10029
rlabel metal2 1423 -436 1423 -436 0 net=10975
rlabel metal2 1521 -436 1521 -436 0 net=11891
rlabel metal2 1640 -436 1640 -436 0 net=12789
rlabel metal2 1731 -436 1731 -436 0 net=13625
rlabel metal2 177 -438 177 -438 0 net=1837
rlabel metal2 310 -438 310 -438 0 net=4119
rlabel metal2 632 -438 632 -438 0 net=167
rlabel metal2 887 -438 887 -438 0 net=12031
rlabel metal2 1717 -438 1717 -438 0 net=13079
rlabel metal2 177 -440 177 -440 0 net=2411
rlabel metal2 408 -440 408 -440 0 net=3785
rlabel metal2 719 -440 719 -440 0 net=10343
rlabel metal2 1444 -440 1444 -440 0 net=10989
rlabel metal2 1577 -440 1577 -440 0 net=12423
rlabel metal2 107 -442 107 -442 0 net=3159
rlabel metal2 415 -442 415 -442 0 net=5139
rlabel metal2 775 -442 775 -442 0 net=10147
rlabel metal2 1451 -442 1451 -442 0 net=11439
rlabel metal2 1598 -442 1598 -442 0 net=12561
rlabel metal2 107 -444 107 -444 0 net=2363
rlabel metal2 310 -444 310 -444 0 net=1937
rlabel metal2 429 -444 429 -444 0 net=2895
rlabel metal2 814 -444 814 -444 0 net=5595
rlabel metal2 870 -444 870 -444 0 net=8491
rlabel metal2 1241 -444 1241 -444 0 net=11003
rlabel metal2 1605 -444 1605 -444 0 net=12569
rlabel metal2 2 -446 2 -446 0 net=3233
rlabel metal2 821 -446 821 -446 0 net=6207
rlabel metal2 905 -446 905 -446 0 net=5943
rlabel metal2 1010 -446 1010 -446 0 net=9225
rlabel metal2 1255 -446 1255 -446 0 net=10225
rlabel metal2 1458 -446 1458 -446 0 net=11799
rlabel metal2 58 -448 58 -448 0 net=5151
rlabel metal2 870 -448 870 -448 0 net=7647
rlabel metal2 1083 -448 1083 -448 0 net=10886
rlabel metal2 1465 -448 1465 -448 0 net=11313
rlabel metal2 128 -450 128 -450 0 net=3661
rlabel metal2 450 -450 450 -450 0 net=12457
rlabel metal2 128 -452 128 -452 0 net=4633
rlabel metal2 198 -452 198 -452 0 net=3909
rlabel metal2 695 -452 695 -452 0 net=4557
rlabel metal2 940 -452 940 -452 0 net=6603
rlabel metal2 1181 -452 1181 -452 0 net=10291
rlabel metal2 1486 -452 1486 -452 0 net=8671
rlabel metal2 142 -454 142 -454 0 net=6485
rlabel metal2 1010 -454 1010 -454 0 net=6723
rlabel metal2 1066 -454 1066 -454 0 net=8135
rlabel metal2 1220 -454 1220 -454 0 net=9341
rlabel metal2 1318 -454 1318 -454 0 net=10539
rlabel metal2 1696 -454 1696 -454 0 net=13067
rlabel metal2 184 -456 184 -456 0 net=4447
rlabel metal2 726 -456 726 -456 0 net=8749
rlabel metal2 1269 -456 1269 -456 0 net=9839
rlabel metal2 1535 -456 1535 -456 0 net=12661
rlabel metal2 184 -458 184 -458 0 net=3079
rlabel metal2 1038 -458 1038 -458 0 net=7397
rlabel metal2 1066 -458 1066 -458 0 net=7165
rlabel metal2 198 -460 198 -460 0 net=5211
rlabel metal2 450 -460 450 -460 0 net=7155
rlabel metal2 898 -460 898 -460 0 net=6289
rlabel metal2 1101 -460 1101 -460 0 net=11689
rlabel metal2 219 -462 219 -462 0 net=6497
rlabel metal2 1045 -462 1045 -462 0 net=6991
rlabel metal2 1108 -462 1108 -462 0 net=7929
rlabel metal2 1199 -462 1199 -462 0 net=8821
rlabel metal2 1283 -462 1283 -462 0 net=9577
rlabel metal2 1416 -462 1416 -462 0 net=10923
rlabel metal2 275 -464 275 -464 0 net=2533
rlabel metal2 576 -464 576 -464 0 net=5889
rlabel metal2 723 -464 723 -464 0 net=10580
rlabel metal2 289 -466 289 -466 0 net=1699
rlabel metal2 583 -466 583 -466 0 net=3807
rlabel metal2 849 -466 849 -466 0 net=10173
rlabel metal2 1339 -466 1339 -466 0 net=9903
rlabel metal2 282 -468 282 -468 0 net=1709
rlabel metal2 317 -468 317 -468 0 net=2951
rlabel metal2 583 -468 583 -468 0 net=3013
rlabel metal2 898 -468 898 -468 0 net=5645
rlabel metal2 961 -468 961 -468 0 net=7331
rlabel metal2 1115 -468 1115 -468 0 net=8179
rlabel metal2 1276 -468 1276 -468 0 net=9399
rlabel metal2 1374 -468 1374 -468 0 net=10697
rlabel metal2 254 -470 254 -470 0 net=2349
rlabel metal2 317 -470 317 -470 0 net=1971
rlabel metal2 740 -470 740 -470 0 net=7685
rlabel metal2 1171 -470 1171 -470 0 net=8241
rlabel metal2 1206 -470 1206 -470 0 net=9357
rlabel metal2 254 -472 254 -472 0 net=3733
rlabel metal2 863 -472 863 -472 0 net=5741
rlabel metal2 992 -472 992 -472 0 net=8625
rlabel metal2 1213 -472 1213 -472 0 net=8963
rlabel metal2 1304 -472 1304 -472 0 net=9685
rlabel metal2 324 -474 324 -474 0 net=4104
rlabel metal2 919 -474 919 -474 0 net=7025
rlabel metal2 1143 -474 1143 -474 0 net=8371
rlabel metal2 1234 -474 1234 -474 0 net=9175
rlabel metal2 324 -476 324 -476 0 net=3651
rlabel metal2 464 -476 464 -476 0 net=3771
rlabel metal2 919 -476 919 -476 0 net=6949
rlabel metal2 1094 -476 1094 -476 0 net=7353
rlabel metal2 1157 -476 1157 -476 0 net=8503
rlabel metal2 331 -478 331 -478 0 net=2509
rlabel metal2 422 -478 422 -478 0 net=4443
rlabel metal2 947 -478 947 -478 0 net=6857
rlabel metal2 975 -478 975 -478 0 net=8265
rlabel metal2 93 -480 93 -480 0 net=8105
rlabel metal2 933 -480 933 -480 0 net=6645
rlabel metal2 989 -480 989 -480 0 net=14293
rlabel metal2 93 -482 93 -482 0 net=5565
rlabel metal2 933 -482 933 -482 0 net=11137
rlabel metal2 338 -484 338 -484 0 net=2151
rlabel metal2 996 -484 996 -484 0 net=7309
rlabel metal2 261 -486 261 -486 0 net=2075
rlabel metal2 835 -486 835 -486 0 net=3705
rlabel metal2 1003 -486 1003 -486 0 net=7737
rlabel metal2 261 -488 261 -488 0 net=4071
rlabel metal2 54 -490 54 -490 0 net=4369
rlabel metal2 352 -492 352 -492 0 net=3629
rlabel metal2 555 -494 555 -494 0 net=5571
rlabel metal2 492 -496 492 -496 0 net=3315
rlabel metal2 492 -498 492 -498 0 net=7981
rlabel metal2 30 -509 30 -509 0 net=3189
rlabel metal2 93 -509 93 -509 0 net=5566
rlabel metal2 205 -509 205 -509 0 net=4458
rlabel metal2 737 -509 737 -509 0 net=12216
rlabel metal2 1682 -509 1682 -509 0 net=14351
rlabel metal2 2214 -509 2214 -509 0 net=8359
rlabel metal2 37 -511 37 -511 0 net=6435
rlabel metal2 656 -511 656 -511 0 net=4448
rlabel metal2 723 -511 723 -511 0 net=5586
rlabel metal2 814 -511 814 -511 0 net=5153
rlabel metal2 814 -511 814 -511 0 net=5153
rlabel metal2 824 -511 824 -511 0 net=7658
rlabel metal2 1146 -511 1146 -511 0 net=10698
rlabel metal2 1535 -511 1535 -511 0 net=10925
rlabel metal2 2039 -511 2039 -511 0 net=14727
rlabel metal2 2263 -511 2263 -511 0 net=14037
rlabel metal2 44 -513 44 -513 0 net=2481
rlabel metal2 215 -513 215 -513 0 net=12650
rlabel metal2 1836 -513 1836 -513 0 net=13105
rlabel metal2 2014 -513 2014 -513 0 net=3615
rlabel metal2 2284 -513 2284 -513 0 net=12545
rlabel metal2 44 -515 44 -515 0 net=6461
rlabel metal2 170 -515 170 -515 0 net=7156
rlabel metal2 541 -515 541 -515 0 net=2329
rlabel metal2 635 -515 635 -515 0 net=4781
rlabel metal2 842 -515 842 -515 0 net=5597
rlabel metal2 898 -515 898 -515 0 net=5646
rlabel metal2 982 -515 982 -515 0 net=12558
rlabel metal2 1864 -515 1864 -515 0 net=13283
rlabel metal2 2088 -515 2088 -515 0 net=3744
rlabel metal2 128 -517 128 -517 0 net=4635
rlabel metal2 128 -517 128 -517 0 net=4635
rlabel metal2 135 -517 135 -517 0 net=6925
rlabel metal2 751 -517 751 -517 0 net=5875
rlabel metal2 786 -517 786 -517 0 net=5249
rlabel metal2 849 -517 849 -517 0 net=6950
rlabel metal2 975 -517 975 -517 0 net=11621
rlabel metal2 1864 -517 1864 -517 0 net=12411
rlabel metal2 1983 -517 1983 -517 0 net=14649
rlabel metal2 75 -519 75 -519 0 net=5781
rlabel metal2 985 -519 985 -519 0 net=11655
rlabel metal2 1794 -519 1794 -519 0 net=12957
rlabel metal2 1990 -519 1990 -519 0 net=12540
rlabel metal2 2116 -519 2116 -519 0 net=13697
rlabel metal2 114 -521 114 -521 0 net=6169
rlabel metal2 992 -521 992 -521 0 net=8266
rlabel metal2 1269 -521 1269 -521 0 net=8823
rlabel metal2 1472 -521 1472 -521 0 net=9917
rlabel metal2 1612 -521 1612 -521 0 net=11819
rlabel metal2 1808 -521 1808 -521 0 net=12993
rlabel metal2 2116 -521 2116 -521 0 net=14359
rlabel metal2 114 -523 114 -523 0 net=2511
rlabel metal2 380 -523 380 -523 0 net=8106
rlabel metal2 996 -523 996 -523 0 net=3706
rlabel metal2 1164 -523 1164 -523 0 net=14291
rlabel metal2 2144 -523 2144 -523 0 net=14779
rlabel metal2 138 -525 138 -525 0 net=5709
rlabel metal2 940 -525 940 -525 0 net=6605
rlabel metal2 1003 -525 1003 -525 0 net=14106
rlabel metal2 1871 -525 1871 -525 0 net=13501
rlabel metal2 163 -527 163 -527 0 net=2393
rlabel metal2 723 -527 723 -527 0 net=7333
rlabel metal2 1167 -527 1167 -527 0 net=12098
rlabel metal2 1395 -527 1395 -527 0 net=9841
rlabel metal2 1619 -527 1619 -527 0 net=11853
rlabel metal2 1878 -527 1878 -527 0 net=13521
rlabel metal2 205 -529 205 -529 0 net=9308
rlabel metal2 1290 -529 1290 -529 0 net=9113
rlabel metal2 1479 -529 1479 -529 0 net=10663
rlabel metal2 1633 -529 1633 -529 0 net=10523
rlabel metal2 219 -531 219 -531 0 net=13909
rlabel metal2 219 -533 219 -533 0 net=2387
rlabel metal2 660 -533 660 -533 0 net=4370
rlabel metal2 1017 -533 1017 -533 0 net=6825
rlabel metal2 1192 -533 1192 -533 0 net=8137
rlabel metal2 1290 -533 1290 -533 0 net=9579
rlabel metal2 1479 -533 1479 -533 0 net=7565
rlabel metal2 79 -535 79 -535 0 net=3995
rlabel metal2 702 -535 702 -535 0 net=6353
rlabel metal2 1024 -535 1024 -535 0 net=9475
rlabel metal2 1367 -535 1367 -535 0 net=8673
rlabel metal2 1640 -535 1640 -535 0 net=12033
rlabel metal2 1885 -535 1885 -535 0 net=13627
rlabel metal2 222 -537 222 -537 0 net=2350
rlabel metal2 296 -537 296 -537 0 net=1615
rlabel metal2 296 -537 296 -537 0 net=1615
rlabel metal2 310 -537 310 -537 0 net=1938
rlabel metal2 716 -537 716 -537 0 net=5107
rlabel metal2 730 -537 730 -537 0 net=4539
rlabel metal2 1031 -537 1031 -537 0 net=6895
rlabel metal2 1136 -537 1136 -537 0 net=7371
rlabel metal2 1227 -537 1227 -537 0 net=8493
rlabel metal2 1493 -537 1493 -537 0 net=10861
rlabel metal2 1661 -537 1661 -537 0 net=12187
rlabel metal2 103 -539 103 -539 0 net=9907
rlabel metal2 1710 -539 1710 -539 0 net=12501
rlabel metal2 1892 -539 1892 -539 0 net=13765
rlabel metal2 1892 -539 1892 -539 0 net=13765
rlabel metal2 1899 -539 1899 -539 0 net=13825
rlabel metal2 226 -541 226 -541 0 net=3818
rlabel metal2 240 -541 240 -541 0 net=2629
rlabel metal2 324 -541 324 -541 0 net=3652
rlabel metal2 534 -541 534 -541 0 net=779
rlabel metal2 1255 -541 1255 -541 0 net=8751
rlabel metal2 1717 -541 1717 -541 0 net=12563
rlabel metal2 1906 -541 1906 -541 0 net=13887
rlabel metal2 65 -543 65 -543 0 net=8075
rlabel metal2 233 -543 233 -543 0 net=11121
rlabel metal2 1731 -543 1731 -543 0 net=12571
rlabel metal2 9 -545 9 -545 0 net=4177
rlabel metal2 72 -545 72 -545 0 net=1703
rlabel metal2 254 -545 254 -545 0 net=3735
rlabel metal2 600 -545 600 -545 0 net=133
rlabel metal2 1570 -545 1570 -545 0 net=11315
rlabel metal2 1738 -545 1738 -545 0 net=12597
rlabel metal2 1913 -545 1913 -545 0 net=14141
rlabel metal2 9 -547 9 -547 0 net=5213
rlabel metal2 233 -547 233 -547 0 net=2897
rlabel metal2 450 -547 450 -547 0 net=4491
rlabel metal2 541 -547 541 -547 0 net=1803
rlabel metal2 751 -547 751 -547 0 net=5945
rlabel metal2 947 -547 947 -547 0 net=6647
rlabel metal2 1034 -547 1034 -547 0 net=14440
rlabel metal2 1941 -547 1941 -547 0 net=14307
rlabel metal2 107 -549 107 -549 0 net=2365
rlabel metal2 282 -549 282 -549 0 net=1701
rlabel metal2 394 -549 394 -549 0 net=2076
rlabel metal2 1062 -549 1062 -549 0 net=13237
rlabel metal2 16 -551 16 -551 0 net=5311
rlabel metal2 177 -551 177 -551 0 net=2413
rlabel metal2 317 -551 317 -551 0 net=1973
rlabel metal2 331 -551 331 -551 0 net=4689
rlabel metal2 565 -551 565 -551 0 net=9226
rlabel metal2 1262 -551 1262 -551 0 net=7867
rlabel metal2 1962 -551 1962 -551 0 net=14479
rlabel metal2 16 -553 16 -553 0 net=9323
rlabel metal2 177 -553 177 -553 0 net=4427
rlabel metal2 891 -553 891 -553 0 net=6001
rlabel metal2 978 -553 978 -553 0 net=11355
rlabel metal2 1759 -553 1759 -553 0 net=12697
rlabel metal2 1948 -553 1948 -553 0 net=14455
rlabel metal2 93 -555 93 -555 0 net=3641
rlabel metal2 569 -555 569 -555 0 net=4120
rlabel metal2 611 -555 611 -555 0 net=4167
rlabel metal2 786 -555 786 -555 0 net=10449
rlabel metal2 1675 -555 1675 -555 0 net=12341
rlabel metal2 1920 -555 1920 -555 0 net=14185
rlabel metal2 1969 -555 1969 -555 0 net=14503
rlabel metal2 121 -557 121 -557 0 net=2461
rlabel metal2 303 -557 303 -557 0 net=1839
rlabel metal2 345 -557 345 -557 0 net=3156
rlabel metal2 492 -557 492 -557 0 net=3067
rlabel metal2 569 -557 569 -557 0 net=4869
rlabel metal2 835 -557 835 -557 0 net=5573
rlabel metal2 905 -557 905 -557 0 net=6859
rlabel metal2 1031 -557 1031 -557 0 net=7763
rlabel metal2 1283 -557 1283 -557 0 net=10175
rlabel metal2 1591 -557 1591 -557 0 net=11647
rlabel metal2 1773 -557 1773 -557 0 net=12757
rlabel metal2 1976 -557 1976 -557 0 net=9074
rlabel metal2 121 -559 121 -559 0 net=2877
rlabel metal2 604 -559 604 -559 0 net=3809
rlabel metal2 621 -559 621 -559 0 net=7648
rlabel metal2 877 -559 877 -559 0 net=6209
rlabel metal2 1297 -559 1297 -559 0 net=8951
rlabel metal2 1696 -559 1696 -559 0 net=12663
rlabel metal2 100 -561 100 -561 0 net=3577
rlabel metal2 649 -561 649 -561 0 net=12135
rlabel metal2 1927 -561 1927 -561 0 net=14295
rlabel metal2 100 -563 100 -563 0 net=3910
rlabel metal2 688 -563 688 -563 0 net=4346
rlabel metal2 985 -563 985 -563 0 net=11063
rlabel metal2 1703 -563 1703 -563 0 net=12459
rlabel metal2 61 -565 61 -565 0 net=4105
rlabel metal2 793 -565 793 -565 0 net=5291
rlabel metal2 1073 -565 1073 -565 0 net=7273
rlabel metal2 1150 -565 1150 -565 0 net=7931
rlabel metal2 1297 -565 1297 -565 0 net=13706
rlabel metal2 1829 -565 1829 -565 0 net=13081
rlabel metal2 2 -567 2 -567 0 net=3234
rlabel metal2 303 -567 303 -567 0 net=3431
rlabel metal2 639 -567 639 -567 0 net=3887
rlabel metal2 793 -567 793 -567 0 net=4775
rlabel metal2 852 -567 852 -567 0 net=7398
rlabel metal2 1080 -567 1080 -567 0 net=9699
rlabel metal2 1724 -567 1724 -567 0 net=12791
rlabel metal2 250 -569 250 -569 0 net=6681
rlabel metal2 1083 -569 1083 -569 0 net=12928
rlabel metal2 338 -571 338 -571 0 net=2153
rlabel metal2 366 -571 366 -571 0 net=3663
rlabel metal2 387 -571 387 -571 0 net=4969
rlabel metal2 436 -571 436 -571 0 net=3767
rlabel metal2 709 -571 709 -571 0 net=4893
rlabel metal2 765 -571 765 -571 0 net=4933
rlabel metal2 863 -571 863 -571 0 net=5743
rlabel metal2 971 -571 971 -571 0 net=11195
rlabel metal2 1745 -571 1745 -571 0 net=12629
rlabel metal2 142 -573 142 -573 0 net=6487
rlabel metal2 821 -573 821 -573 0 net=4559
rlabel metal2 863 -573 863 -573 0 net=12219
rlabel metal2 1703 -573 1703 -573 0 net=13069
rlabel metal2 142 -575 142 -575 0 net=1823
rlabel metal2 408 -575 408 -575 0 net=3161
rlabel metal2 527 -575 527 -575 0 net=3317
rlabel metal2 695 -575 695 -575 0 net=3849
rlabel metal2 954 -575 954 -575 0 net=10007
rlabel metal2 1780 -575 1780 -575 0 net=12889
rlabel metal2 117 -577 117 -577 0 net=6153
rlabel metal2 415 -577 415 -577 0 net=5140
rlabel metal2 856 -577 856 -577 0 net=5815
rlabel metal2 1010 -577 1010 -577 0 net=6725
rlabel metal2 1094 -577 1094 -577 0 net=7311
rlabel metal2 1216 -577 1216 -577 0 net=13005
rlabel metal2 275 -579 275 -579 0 net=2535
rlabel metal2 422 -579 422 -579 0 net=4445
rlabel metal2 495 -579 495 -579 0 net=1358
rlabel metal2 758 -579 758 -579 0 net=5075
rlabel metal2 800 -579 800 -579 0 net=5525
rlabel metal2 1010 -579 1010 -579 0 net=12905
rlabel metal2 86 -581 86 -581 0 net=4879
rlabel metal2 1094 -581 1094 -581 0 net=10851
rlabel metal2 86 -583 86 -583 0 net=3631
rlabel metal2 359 -583 359 -583 0 net=1979
rlabel metal2 506 -583 506 -583 0 net=5208
rlabel metal2 586 -583 586 -583 0 net=10461
rlabel metal2 58 -585 58 -585 0 net=2177
rlabel metal2 359 -585 359 -585 0 net=2279
rlabel metal2 555 -585 555 -585 0 net=4585
rlabel metal2 1101 -585 1101 -585 0 net=6993
rlabel metal2 1220 -585 1220 -585 0 net=8181
rlabel metal2 1325 -585 1325 -585 0 net=10929
rlabel metal2 23 -587 23 -587 0 net=8423
rlabel metal2 1332 -587 1332 -587 0 net=6392
rlabel metal2 23 -589 23 -589 0 net=4993
rlabel metal2 275 -589 275 -589 0 net=2953
rlabel metal2 471 -589 471 -589 0 net=3125
rlabel metal2 674 -589 674 -589 0 net=4207
rlabel metal2 1080 -589 1080 -589 0 net=6977
rlabel metal2 1199 -589 1199 -589 0 net=8243
rlabel metal2 1234 -589 1234 -589 0 net=8505
rlabel metal2 1353 -589 1353 -589 0 net=9269
rlabel metal2 1465 -589 1465 -589 0 net=10541
rlabel metal2 51 -591 51 -591 0 net=6329
rlabel metal2 667 -591 667 -591 0 net=4257
rlabel metal2 681 -591 681 -591 0 net=4077
rlabel metal2 1248 -591 1248 -591 0 net=8737
rlabel metal2 1416 -591 1416 -591 0 net=9905
rlabel metal2 1850 -591 1850 -591 0 net=13155
rlabel metal2 135 -593 135 -593 0 net=4759
rlabel metal2 464 -593 464 -593 0 net=3773
rlabel metal2 1157 -593 1157 -593 0 net=7739
rlabel metal2 1318 -593 1318 -593 0 net=9359
rlabel metal2 1500 -593 1500 -593 0 net=10881
rlabel metal2 184 -595 184 -595 0 net=3081
rlabel metal2 576 -595 576 -595 0 net=5891
rlabel metal2 1087 -595 1087 -595 0 net=7075
rlabel metal2 1311 -595 1311 -595 0 net=9343
rlabel metal2 1402 -595 1402 -595 0 net=9939
rlabel metal2 1521 -595 1521 -595 0 net=10991
rlabel metal2 184 -597 184 -597 0 net=4073
rlabel metal2 289 -597 289 -597 0 net=1711
rlabel metal2 576 -597 576 -597 0 net=3497
rlabel metal2 618 -597 618 -597 0 net=7713
rlabel metal2 1304 -597 1304 -597 0 net=9177
rlabel metal2 1416 -597 1416 -597 0 net=10049
rlabel metal2 149 -599 149 -599 0 net=2887
rlabel metal2 289 -599 289 -599 0 net=4065
rlabel metal2 1206 -599 1206 -599 0 net=8373
rlabel metal2 1430 -599 1430 -599 0 net=10069
rlabel metal2 1528 -599 1528 -599 0 net=11999
rlabel metal2 1857 -599 1857 -599 0 net=13191
rlabel metal2 149 -601 149 -601 0 net=5777
rlabel metal2 338 -601 338 -601 0 net=2483
rlabel metal2 1115 -601 1115 -601 0 net=7687
rlabel metal2 1440 -601 1440 -601 0 net=12161
rlabel metal2 79 -603 79 -603 0 net=8115
rlabel metal2 366 -603 366 -603 0 net=4151
rlabel metal2 912 -603 912 -603 0 net=8317
rlabel metal2 1528 -603 1528 -603 0 net=11441
rlabel metal2 1598 -603 1598 -603 0 net=11691
rlabel metal2 373 -605 373 -605 0 net=2977
rlabel metal2 590 -605 590 -605 0 net=5327
rlabel metal2 929 -605 929 -605 0 net=6539
rlabel metal2 1178 -605 1178 -605 0 net=9661
rlabel metal2 1458 -605 1458 -605 0 net=10293
rlabel metal2 1605 -605 1605 -605 0 net=11801
rlabel metal2 191 -607 191 -607 0 net=3899
rlabel metal2 394 -607 394 -607 0 net=3363
rlabel metal2 807 -607 807 -607 0 net=5095
rlabel metal2 933 -607 933 -607 0 net=5785
rlabel metal2 1045 -607 1045 -607 0 net=7027
rlabel metal2 1143 -607 1143 -607 0 net=7355
rlabel metal2 1388 -607 1388 -607 0 net=9705
rlabel metal2 1507 -607 1507 -607 0 net=10129
rlabel metal2 1668 -607 1668 -607 0 net=12237
rlabel metal2 173 -609 173 -609 0 net=2487
rlabel metal2 443 -609 443 -609 0 net=5677
rlabel metal2 926 -609 926 -609 0 net=6499
rlabel metal2 1143 -609 1143 -609 0 net=13864
rlabel metal2 443 -611 443 -611 0 net=3787
rlabel metal2 926 -611 926 -611 0 net=10918
rlabel metal2 1549 -611 1549 -611 0 net=11833
rlabel metal2 485 -613 485 -613 0 net=3199
rlabel metal2 1202 -613 1202 -613 0 net=10103
rlabel metal2 1626 -613 1626 -613 0 net=11893
rlabel metal2 485 -615 485 -615 0 net=3015
rlabel metal2 1276 -615 1276 -615 0 net=8965
rlabel metal2 1423 -615 1423 -615 0 net=10345
rlabel metal2 1668 -615 1668 -615 0 net=12425
rlabel metal2 499 -617 499 -617 0 net=4059
rlabel metal2 1185 -617 1185 -617 0 net=7983
rlabel metal2 1339 -617 1339 -617 0 net=9401
rlabel metal2 1444 -617 1444 -617 0 net=10149
rlabel metal2 1556 -617 1556 -617 0 net=11005
rlabel metal2 583 -619 583 -619 0 net=12348
rlabel metal2 1059 -621 1059 -621 0 net=7215
rlabel metal2 1381 -621 1381 -621 0 net=9687
rlabel metal2 1451 -621 1451 -621 0 net=10227
rlabel metal2 1059 -623 1059 -623 0 net=14763
rlabel metal2 1066 -625 1066 -625 0 net=7167
rlabel metal2 1507 -625 1507 -625 0 net=10977
rlabel metal2 1556 -625 1556 -625 0 net=11139
rlabel metal2 1584 -625 1584 -625 0 net=11563
rlabel metal2 1052 -627 1052 -627 0 net=6291
rlabel metal2 1171 -627 1171 -627 0 net=8627
rlabel metal2 1409 -627 1409 -627 0 net=10031
rlabel metal2 1563 -627 1563 -627 0 net=7239
rlabel metal2 268 -629 268 -629 0 net=6389
rlabel metal2 1199 -629 1199 -629 0 net=10009
rlabel metal2 1409 -629 1409 -629 0 net=8901
rlabel metal2 268 -631 268 -631 0 net=2117
rlabel metal2 915 -631 915 -631 0 net=8695
rlabel metal2 1489 -631 1489 -631 0 net=10199
rlabel metal2 2 -642 2 -642 0 net=2879
rlabel metal2 131 -642 131 -642 0 net=14292
rlabel metal2 2144 -642 2144 -642 0 net=14505
rlabel metal2 2326 -642 2326 -642 0 net=12547
rlabel metal2 2361 -642 2361 -642 0 net=14039
rlabel metal2 44 -644 44 -644 0 net=6462
rlabel metal2 1300 -644 1300 -644 0 net=14142
rlabel metal2 2137 -644 2137 -644 0 net=14729
rlabel metal2 2193 -644 2193 -644 0 net=13698
rlabel metal2 2214 -644 2214 -644 0 net=14323
rlabel metal2 2291 -644 2291 -644 0 net=8361
rlabel metal2 47 -646 47 -646 0 net=4178
rlabel metal2 68 -646 68 -646 0 net=574
rlabel metal2 807 -646 807 -646 0 net=6896
rlabel metal2 1143 -646 1143 -646 0 net=8952
rlabel metal2 1703 -646 1703 -646 0 net=13071
rlabel metal2 12 -648 12 -648 0 net=1424
rlabel metal2 72 -648 72 -648 0 net=10462
rlabel metal2 1843 -648 1843 -648 0 net=12137
rlabel metal2 51 -650 51 -650 0 net=6330
rlabel metal2 940 -650 940 -650 0 net=12342
rlabel metal2 1955 -650 1955 -650 0 net=14187
rlabel metal2 51 -652 51 -652 0 net=4079
rlabel metal2 698 -652 698 -652 0 net=5853
rlabel metal2 1010 -652 1010 -652 0 net=14352
rlabel metal2 2158 -652 2158 -652 0 net=14651
rlabel metal2 58 -654 58 -654 0 net=10852
rlabel metal2 1885 -654 1885 -654 0 net=13083
rlabel metal2 2200 -654 2200 -654 0 net=14780
rlabel metal2 72 -656 72 -656 0 net=6355
rlabel metal2 1059 -656 1059 -656 0 net=10228
rlabel metal2 1885 -656 1885 -656 0 net=12891
rlabel metal2 2004 -656 2004 -656 0 net=13107
rlabel metal2 82 -658 82 -658 0 net=1144
rlabel metal2 1059 -658 1059 -658 0 net=6727
rlabel metal2 1083 -658 1083 -658 0 net=9360
rlabel metal2 1486 -658 1486 -658 0 net=14456
rlabel metal2 16 -660 16 -660 0 net=9325
rlabel metal2 1094 -660 1094 -660 0 net=14764
rlabel metal2 93 -662 93 -662 0 net=3642
rlabel metal2 618 -662 618 -662 0 net=5679
rlabel metal2 957 -662 957 -662 0 net=6390
rlabel metal2 1062 -662 1062 -662 0 net=3616
rlabel metal2 93 -664 93 -664 0 net=1825
rlabel metal2 145 -664 145 -664 0 net=1058
rlabel metal2 1052 -664 1052 -664 0 net=6827
rlabel metal2 1150 -664 1150 -664 0 net=13483
rlabel metal2 75 -666 75 -666 0 net=211
rlabel metal2 1136 -666 1136 -666 0 net=6995
rlabel metal2 1174 -666 1174 -666 0 net=14561
rlabel metal2 135 -668 135 -668 0 net=11802
rlabel metal2 1857 -668 1857 -668 0 net=12239
rlabel metal2 2011 -668 2011 -668 0 net=13157
rlabel metal2 170 -670 170 -670 0 net=2631
rlabel metal2 401 -670 401 -670 0 net=6155
rlabel metal2 1101 -670 1101 -670 0 net=6979
rlabel metal2 1178 -670 1178 -670 0 net=7356
rlabel metal2 1216 -670 1216 -670 0 net=13888
rlabel metal2 2116 -670 2116 -670 0 net=14361
rlabel metal2 173 -672 173 -672 0 net=12460
rlabel metal2 1983 -672 1983 -672 0 net=12959
rlabel metal2 2123 -672 2123 -672 0 net=14481
rlabel metal2 187 -674 187 -674 0 net=4168
rlabel metal2 733 -674 733 -674 0 net=13297
rlabel metal2 205 -676 205 -676 0 net=7168
rlabel metal2 1493 -676 1493 -676 0 net=9909
rlabel metal2 1717 -676 1717 -676 0 net=11123
rlabel metal2 1864 -676 1864 -676 0 net=12413
rlabel metal2 2018 -676 2018 -676 0 net=13193
rlabel metal2 212 -678 212 -678 0 net=2482
rlabel metal2 765 -678 765 -678 0 net=6489
rlabel metal2 1101 -678 1101 -678 0 net=5467
rlabel metal2 1199 -678 1199 -678 0 net=12083
rlabel metal2 1990 -678 1990 -678 0 net=12995
rlabel metal2 191 -680 191 -680 0 net=2489
rlabel metal2 236 -680 236 -680 0 net=9005
rlabel metal2 1213 -680 1213 -680 0 net=8902
rlabel metal2 1430 -680 1430 -680 0 net=9663
rlabel metal2 1605 -680 1605 -680 0 net=10347
rlabel metal2 1738 -680 1738 -680 0 net=11357
rlabel metal2 1892 -680 1892 -680 0 net=13767
rlabel metal2 1892 -680 1892 -680 0 net=13767
rlabel metal2 1990 -680 1990 -680 0 net=13629
rlabel metal2 2074 -680 2074 -680 0 net=13827
rlabel metal2 149 -682 149 -682 0 net=5779
rlabel metal2 247 -682 247 -682 0 net=1841
rlabel metal2 366 -682 366 -682 0 net=4153
rlabel metal2 800 -682 800 -682 0 net=4881
rlabel metal2 824 -682 824 -682 0 net=14363
rlabel metal2 30 -684 30 -684 0 net=3191
rlabel metal2 366 -684 366 -684 0 net=4783
rlabel metal2 849 -684 849 -684 0 net=12220
rlabel metal2 891 -684 891 -684 0 net=5575
rlabel metal2 929 -684 929 -684 0 net=11957
rlabel metal2 1962 -684 1962 -684 0 net=12793
rlabel metal2 2081 -684 2081 -684 0 net=13911
rlabel metal2 9 -686 9 -686 0 net=5215
rlabel metal2 877 -686 877 -686 0 net=5329
rlabel metal2 1080 -686 1080 -686 0 net=10633
rlabel metal2 1752 -686 1752 -686 0 net=11623
rlabel metal2 2088 -686 2088 -686 0 net=14297
rlabel metal2 19 -688 19 -688 0 net=11803
rlabel metal2 2095 -688 2095 -688 0 net=14309
rlabel metal2 30 -690 30 -690 0 net=6437
rlabel metal2 149 -690 149 -690 0 net=2925
rlabel metal2 1080 -690 1080 -690 0 net=6541
rlabel metal2 1129 -690 1129 -690 0 net=7275
rlabel metal2 1360 -690 1360 -690 0 net=8753
rlabel metal2 1549 -690 1549 -690 0 net=10151
rlabel metal2 1759 -690 1759 -690 0 net=11649
rlabel metal2 37 -692 37 -692 0 net=7335
rlabel metal2 730 -692 730 -692 0 net=7383
rlabel metal2 1556 -692 1556 -692 0 net=11141
rlabel metal2 1976 -692 1976 -692 0 net=12907
rlabel metal2 261 -694 261 -694 0 net=2888
rlabel metal2 401 -694 401 -694 0 net=4587
rlabel metal2 562 -694 562 -694 0 net=5893
rlabel metal2 681 -694 681 -694 0 net=9700
rlabel metal2 1794 -694 1794 -694 0 net=11821
rlabel metal2 1997 -694 1997 -694 0 net=13007
rlabel metal2 156 -696 156 -696 0 net=2463
rlabel metal2 282 -696 282 -696 0 net=1702
rlabel metal2 590 -696 590 -696 0 net=4803
rlabel metal2 702 -696 702 -696 0 net=8319
rlabel metal2 1360 -696 1360 -696 0 net=9906
rlabel metal2 1829 -696 1829 -696 0 net=12001
rlabel metal2 2025 -696 2025 -696 0 net=13239
rlabel metal2 128 -698 128 -698 0 net=4637
rlabel metal2 240 -698 240 -698 0 net=1705
rlabel metal2 310 -698 310 -698 0 net=3127
rlabel metal2 523 -698 523 -698 0 net=8991
rlabel metal2 1507 -698 1507 -698 0 net=10979
rlabel metal2 1829 -698 1829 -698 0 net=12699
rlabel metal2 2039 -698 2039 -698 0 net=12188
rlabel metal2 114 -700 114 -700 0 net=2513
rlabel metal2 324 -700 324 -700 0 net=1975
rlabel metal2 548 -700 548 -700 0 net=3578
rlabel metal2 569 -700 569 -700 0 net=4871
rlabel metal2 814 -700 814 -700 0 net=5155
rlabel metal2 852 -700 852 -700 0 net=10008
rlabel metal2 1808 -700 1808 -700 0 net=11855
rlabel metal2 2046 -700 2046 -700 0 net=13285
rlabel metal2 86 -702 86 -702 0 net=3633
rlabel metal2 324 -702 324 -702 0 net=3083
rlabel metal2 492 -702 492 -702 0 net=3068
rlabel metal2 737 -702 737 -702 0 net=6927
rlabel metal2 737 -702 737 -702 0 net=6927
rlabel metal2 744 -702 744 -702 0 net=13581
rlabel metal2 5 -704 5 -704 0 net=2597
rlabel metal2 415 -704 415 -704 0 net=2119
rlabel metal2 492 -704 492 -704 0 net=3851
rlabel metal2 747 -704 747 -704 0 net=12572
rlabel metal2 408 -706 408 -706 0 net=2537
rlabel metal2 429 -706 429 -706 0 net=3513
rlabel metal2 590 -706 590 -706 0 net=8895
rlabel metal2 1584 -706 1584 -706 0 net=10201
rlabel metal2 1836 -706 1836 -706 0 net=12035
rlabel metal2 2053 -706 2053 -706 0 net=13503
rlabel metal2 303 -708 303 -708 0 net=3433
rlabel metal2 422 -708 422 -708 0 net=1981
rlabel metal2 432 -708 432 -708 0 net=3774
rlabel metal2 639 -708 639 -708 0 net=3889
rlabel metal2 1850 -708 1850 -708 0 net=12163
rlabel metal2 2060 -708 2060 -708 0 net=13523
rlabel metal2 100 -710 100 -710 0 net=10183
rlabel metal2 646 -710 646 -710 0 net=6210
rlabel metal2 1248 -710 1248 -710 0 net=7741
rlabel metal2 1871 -710 1871 -710 0 net=12503
rlabel metal2 100 -712 100 -712 0 net=2367
rlabel metal2 219 -712 219 -712 0 net=2389
rlabel metal2 422 -712 422 -712 0 net=7185
rlabel metal2 1248 -712 1248 -712 0 net=9707
rlabel metal2 1528 -712 1528 -712 0 net=11443
rlabel metal2 1878 -712 1878 -712 0 net=12565
rlabel metal2 163 -714 163 -714 0 net=2395
rlabel metal2 443 -714 443 -714 0 net=3789
rlabel metal2 604 -714 604 -714 0 net=3769
rlabel metal2 653 -714 653 -714 0 net=3996
rlabel metal2 814 -714 814 -714 0 net=5293
rlabel metal2 947 -714 947 -714 0 net=5744
rlabel metal2 1136 -714 1136 -714 0 net=10653
rlabel metal2 1899 -714 1899 -714 0 net=12599
rlabel metal2 163 -716 163 -716 0 net=3017
rlabel metal2 534 -716 534 -716 0 net=3263
rlabel metal2 576 -716 576 -716 0 net=3499
rlabel metal2 611 -716 611 -716 0 net=3811
rlabel metal2 660 -716 660 -716 0 net=14071
rlabel metal2 23 -718 23 -718 0 net=4995
rlabel metal2 583 -718 583 -718 0 net=8333
rlabel metal2 996 -718 996 -718 0 net=6607
rlabel metal2 1097 -718 1097 -718 0 net=9227
rlabel metal2 1598 -718 1598 -718 0 net=10295
rlabel metal2 1724 -718 1724 -718 0 net=11197
rlabel metal2 1920 -718 1920 -718 0 net=12631
rlabel metal2 23 -720 23 -720 0 net=5977
rlabel metal2 772 -720 772 -720 0 net=4209
rlabel metal2 793 -720 793 -720 0 net=4777
rlabel metal2 989 -720 989 -720 0 net=4541
rlabel metal2 1045 -720 1045 -720 0 net=6501
rlabel metal2 1598 -720 1598 -720 0 net=10993
rlabel metal2 1689 -720 1689 -720 0 net=11007
rlabel metal2 1920 -720 1920 -720 0 net=12759
rlabel metal2 289 -722 289 -722 0 net=4067
rlabel metal2 663 -722 663 -722 0 net=4894
rlabel metal2 758 -722 758 -722 0 net=5077
rlabel metal2 856 -722 856 -722 0 net=5527
rlabel metal2 856 -722 856 -722 0 net=5527
rlabel metal2 1045 -722 1045 -722 0 net=6293
rlabel metal2 1143 -722 1143 -722 0 net=12965
rlabel metal2 184 -724 184 -724 0 net=4075
rlabel metal2 779 -724 779 -724 0 net=7029
rlabel metal2 1192 -724 1192 -724 0 net=7373
rlabel metal2 1255 -724 1255 -724 0 net=7933
rlabel metal2 1367 -724 1367 -724 0 net=8675
rlabel metal2 1437 -724 1437 -724 0 net=9271
rlabel metal2 1570 -724 1570 -724 0 net=10177
rlabel metal2 1731 -724 1731 -724 0 net=11317
rlabel metal2 1934 -724 1934 -724 0 net=12665
rlabel metal2 184 -726 184 -726 0 net=5108
rlabel metal2 898 -726 898 -726 0 net=5711
rlabel metal2 1171 -726 1171 -726 0 net=8697
rlabel metal2 1577 -726 1577 -726 0 net=10131
rlabel metal2 1766 -726 1766 -726 0 net=11657
rlabel metal2 177 -728 177 -728 0 net=4429
rlabel metal2 898 -728 898 -728 0 net=5397
rlabel metal2 1171 -728 1171 -728 0 net=8601
rlabel metal2 1423 -728 1423 -728 0 net=9403
rlabel metal2 1605 -728 1605 -728 0 net=10863
rlabel metal2 1647 -728 1647 -728 0 net=10883
rlabel metal2 1801 -728 1801 -728 0 net=11835
rlabel metal2 58 -730 58 -730 0 net=3601
rlabel metal2 1234 -730 1234 -730 0 net=7715
rlabel metal2 1290 -730 1290 -730 0 net=9581
rlabel metal2 1612 -730 1612 -730 0 net=10451
rlabel metal2 1815 -730 1815 -730 0 net=11895
rlabel metal2 177 -732 177 -732 0 net=8139
rlabel metal2 1339 -732 1339 -732 0 net=8629
rlabel metal2 1444 -732 1444 -732 0 net=9689
rlabel metal2 219 -734 219 -734 0 net=9783
rlabel metal2 1619 -734 1619 -734 0 net=10665
rlabel metal2 250 -736 250 -736 0 net=7249
rlabel metal2 1206 -736 1206 -736 0 net=7689
rlabel metal2 1353 -736 1353 -736 0 net=8739
rlabel metal2 1472 -736 1472 -736 0 net=9843
rlabel metal2 1633 -736 1633 -736 0 net=10525
rlabel metal2 142 -738 142 -738 0 net=8903
rlabel metal2 1500 -738 1500 -738 0 net=9941
rlabel metal2 1654 -738 1654 -738 0 net=11565
rlabel metal2 205 -740 205 -740 0 net=9035
rlabel metal2 1514 -740 1514 -740 0 net=10033
rlabel metal2 1668 -740 1668 -740 0 net=12427
rlabel metal2 289 -742 289 -742 0 net=4061
rlabel metal2 537 -742 537 -742 0 net=9157
rlabel metal2 1024 -742 1024 -742 0 net=9477
rlabel metal2 1696 -742 1696 -742 0 net=11065
rlabel metal2 373 -744 373 -744 0 net=3901
rlabel metal2 352 -746 352 -746 0 net=2179
rlabel metal2 380 -746 380 -746 0 net=3665
rlabel metal2 611 -746 611 -746 0 net=4107
rlabel metal2 726 -746 726 -746 0 net=8193
rlabel metal2 1370 -746 1370 -746 0 net=11253
rlabel metal2 254 -748 254 -748 0 net=2415
rlabel metal2 394 -748 394 -748 0 net=3365
rlabel metal2 632 -748 632 -748 0 net=2331
rlabel metal2 674 -748 674 -748 0 net=4259
rlabel metal2 1017 -748 1017 -748 0 net=6649
rlabel metal2 1038 -748 1038 -748 0 net=6683
rlabel metal2 1185 -748 1185 -748 0 net=7217
rlabel metal2 1241 -748 1241 -748 0 net=7765
rlabel metal2 1374 -748 1374 -748 0 net=8825
rlabel metal2 1514 -748 1514 -748 0 net=10071
rlabel metal2 1535 -748 1535 -748 0 net=9919
rlabel metal2 254 -750 254 -750 0 net=3201
rlabel metal2 597 -750 597 -750 0 net=3737
rlabel metal2 688 -750 688 -750 0 net=7313
rlabel metal2 1185 -750 1185 -750 0 net=7241
rlabel metal2 331 -752 331 -752 0 net=4691
rlabel metal2 387 -752 387 -752 0 net=4971
rlabel metal2 968 -752 968 -752 0 net=6003
rlabel metal2 1094 -752 1094 -752 0 net=9235
rlabel metal2 1346 -752 1346 -752 0 net=8495
rlabel metal2 1535 -752 1535 -752 0 net=11405
rlabel metal2 275 -754 275 -754 0 net=2955
rlabel metal2 387 -754 387 -754 0 net=2979
rlabel metal2 499 -754 499 -754 0 net=3163
rlabel metal2 933 -754 933 -754 0 net=5787
rlabel metal2 975 -754 975 -754 0 net=6171
rlabel metal2 1139 -754 1139 -754 0 net=12023
rlabel metal2 1381 -754 1381 -754 0 net=10011
rlabel metal2 275 -756 275 -756 0 net=1617
rlabel metal2 359 -756 359 -756 0 net=2281
rlabel metal2 513 -756 513 -756 0 net=5783
rlabel metal2 954 -756 954 -756 0 net=5817
rlabel metal2 1153 -756 1153 -756 0 net=7485
rlabel metal2 1283 -756 1283 -756 0 net=8183
rlabel metal2 1395 -756 1395 -756 0 net=9115
rlabel metal2 1538 -756 1538 -756 0 net=7515
rlabel metal2 208 -758 208 -758 0 net=5183
rlabel metal2 1157 -758 1157 -758 0 net=7077
rlabel metal2 1206 -758 1206 -758 0 net=8244
rlabel metal2 1311 -758 1311 -758 0 net=8375
rlabel metal2 1395 -758 1395 -758 0 net=9179
rlabel metal2 1542 -758 1542 -758 0 net=10105
rlabel metal2 44 -760 44 -760 0 net=9253
rlabel metal2 135 -762 135 -762 0 net=4467
rlabel metal2 296 -762 296 -762 0 net=1805
rlabel metal2 786 -762 786 -762 0 net=7315
rlabel metal2 961 -762 961 -762 0 net=5877
rlabel metal2 1318 -762 1318 -762 0 net=9345
rlabel metal2 345 -764 345 -764 0 net=2154
rlabel metal2 443 -764 443 -764 0 net=3319
rlabel metal2 810 -764 810 -764 0 net=10743
rlabel metal2 79 -766 79 -766 0 net=8117
rlabel metal2 884 -766 884 -766 0 net=5599
rlabel metal2 1157 -766 1157 -766 0 net=10926
rlabel metal2 79 -768 79 -768 0 net=10899
rlabel metal2 905 -768 905 -768 0 net=6861
rlabel metal2 1209 -768 1209 -768 0 net=12513
rlabel metal2 107 -770 107 -770 0 net=5313
rlabel metal2 1220 -770 1220 -770 0 net=13723
rlabel metal2 107 -772 107 -772 0 net=6715
rlabel metal2 1262 -772 1262 -772 0 net=7869
rlabel metal2 268 -774 268 -774 0 net=5427
rlabel metal2 268 -776 268 -776 0 net=2485
rlabel metal2 345 -776 345 -776 0 net=3675
rlabel metal2 821 -776 821 -776 0 net=4561
rlabel metal2 880 -776 880 -776 0 net=7627
rlabel metal2 338 -778 338 -778 0 net=5947
rlabel metal2 828 -778 828 -778 0 net=4935
rlabel metal2 450 -780 450 -780 0 net=4493
rlabel metal2 751 -780 751 -780 0 net=10050
rlabel metal2 128 -782 128 -782 0 net=8603
rlabel metal2 233 -784 233 -784 0 net=2899
rlabel metal2 457 -784 457 -784 0 net=4761
rlabel metal2 828 -784 828 -784 0 net=10542
rlabel metal2 233 -786 233 -786 0 net=4241
rlabel metal2 457 -786 457 -786 0 net=5251
rlabel metal2 1787 -786 1787 -786 0 net=11693
rlabel metal2 471 -788 471 -788 0 net=1713
rlabel metal2 842 -788 842 -788 0 net=5097
rlabel metal2 1661 -788 1661 -788 0 net=10931
rlabel metal2 471 -790 471 -790 0 net=6063
rlabel metal2 1276 -790 1276 -790 0 net=7985
rlabel metal2 520 -792 520 -792 0 net=8007
rlabel metal2 912 -794 912 -794 0 net=3861
rlabel metal2 1276 -796 1276 -796 0 net=7567
rlabel metal2 1297 -798 1297 -798 0 net=8507
rlabel metal2 1388 -798 1388 -798 0 net=8967
rlabel metal2 1325 -800 1325 -800 0 net=8425
rlabel metal2 226 -802 226 -802 0 net=8077
rlabel metal2 1332 -802 1332 -802 0 net=11661
rlabel metal2 226 -804 226 -804 0 net=4225
rlabel metal2 436 -806 436 -806 0 net=4446
rlabel metal2 222 -808 222 -808 0 net=2653
rlabel metal2 9 -819 9 -819 0 net=9910
rlabel metal2 1661 -819 1661 -819 0 net=7987
rlabel metal2 2403 -819 2403 -819 0 net=14041
rlabel metal2 9 -821 9 -821 0 net=1827
rlabel metal2 103 -821 103 -821 0 net=4692
rlabel metal2 457 -821 457 -821 0 net=5252
rlabel metal2 614 -821 614 -821 0 net=4068
rlabel metal2 674 -821 674 -821 0 net=3738
rlabel metal2 782 -821 782 -821 0 net=5156
rlabel metal2 898 -821 898 -821 0 net=5399
rlabel metal2 898 -821 898 -821 0 net=5399
rlabel metal2 947 -821 947 -821 0 net=8334
rlabel metal2 1332 -821 1332 -821 0 net=8631
rlabel metal2 1538 -821 1538 -821 0 net=11650
rlabel metal2 2326 -821 2326 -821 0 net=8362
rlabel metal2 2343 -821 2343 -821 0 net=14217
rlabel metal2 16 -823 16 -823 0 net=5780
rlabel metal2 212 -823 212 -823 0 net=2491
rlabel metal2 212 -823 212 -823 0 net=2491
rlabel metal2 222 -823 222 -823 0 net=13912
rlabel metal2 2277 -823 2277 -823 0 net=14325
rlabel metal2 2347 -823 2347 -823 0 net=12549
rlabel metal2 16 -825 16 -825 0 net=8079
rlabel metal2 1335 -825 1335 -825 0 net=8496
rlabel metal2 1598 -825 1598 -825 0 net=10995
rlabel metal2 1626 -825 1626 -825 0 net=10035
rlabel metal2 1661 -825 1661 -825 0 net=11067
rlabel metal2 1934 -825 1934 -825 0 net=11837
rlabel metal2 1934 -825 1934 -825 0 net=11837
rlabel metal2 2095 -825 2095 -825 0 net=13159
rlabel metal2 2277 -825 2277 -825 0 net=10379
rlabel metal2 2347 -825 2347 -825 0 net=8933
rlabel metal2 44 -827 44 -827 0 net=3902
rlabel metal2 1815 -827 1815 -827 0 net=11567
rlabel metal2 2151 -827 2151 -827 0 net=13299
rlabel metal2 44 -829 44 -829 0 net=5681
rlabel metal2 947 -829 947 -829 0 net=5789
rlabel metal2 989 -829 989 -829 0 net=9159
rlabel metal2 1598 -829 1598 -829 0 net=10349
rlabel metal2 1878 -829 1878 -829 0 net=11857
rlabel metal2 1990 -829 1990 -829 0 net=13631
rlabel metal2 58 -831 58 -831 0 net=3602
rlabel metal2 817 -831 817 -831 0 net=8602
rlabel metal2 1899 -831 1899 -831 0 net=11659
rlabel metal2 58 -833 58 -833 0 net=4469
rlabel metal2 142 -833 142 -833 0 net=6135
rlabel metal2 254 -833 254 -833 0 net=3203
rlabel metal2 635 -833 635 -833 0 net=5576
rlabel metal2 989 -833 989 -833 0 net=6035
rlabel metal2 1136 -833 1136 -833 0 net=9690
rlabel metal2 1941 -833 1941 -833 0 net=12085
rlabel metal2 79 -835 79 -835 0 net=2464
rlabel metal2 282 -835 282 -835 0 net=1706
rlabel metal2 422 -835 422 -835 0 net=7187
rlabel metal2 870 -835 870 -835 0 net=4779
rlabel metal2 996 -835 996 -835 0 net=4542
rlabel metal2 1248 -835 1248 -835 0 net=9709
rlabel metal2 1605 -835 1605 -835 0 net=10865
rlabel metal2 1983 -835 1983 -835 0 net=12505
rlabel metal2 72 -837 72 -837 0 net=6357
rlabel metal2 1020 -837 1020 -837 0 net=6502
rlabel metal2 1573 -837 1573 -837 0 net=12843
rlabel metal2 72 -839 72 -839 0 net=4805
rlabel metal2 681 -839 681 -839 0 net=4431
rlabel metal2 821 -839 821 -839 0 net=4563
rlabel metal2 926 -839 926 -839 0 net=7251
rlabel metal2 1195 -839 1195 -839 0 net=12960
rlabel metal2 79 -841 79 -841 0 net=3085
rlabel metal2 352 -841 352 -841 0 net=3165
rlabel metal2 506 -841 506 -841 0 net=1976
rlabel metal2 772 -841 772 -841 0 net=4211
rlabel metal2 1010 -841 1010 -841 0 net=13205
rlabel metal2 121 -843 121 -843 0 net=2486
rlabel metal2 282 -843 282 -843 0 net=2421
rlabel metal2 1174 -843 1174 -843 0 net=10884
rlabel metal2 47 -845 47 -845 0 net=10425
rlabel metal2 128 -847 128 -847 0 net=5894
rlabel metal2 646 -847 646 -847 0 net=1714
rlabel metal2 1010 -847 1010 -847 0 net=6609
rlabel metal2 1094 -847 1094 -847 0 net=6980
rlabel metal2 1129 -847 1129 -847 0 net=13072
rlabel metal2 128 -849 128 -849 0 net=4757
rlabel metal2 1045 -849 1045 -849 0 net=6295
rlabel metal2 1094 -849 1094 -849 0 net=5469
rlabel metal2 1111 -849 1111 -849 0 net=12566
rlabel metal2 2235 -849 2235 -849 0 net=14365
rlabel metal2 145 -851 145 -851 0 net=4872
rlabel metal2 828 -851 828 -851 0 net=7441
rlabel metal2 1136 -851 1136 -851 0 net=7375
rlabel metal2 1248 -851 1248 -851 0 net=8427
rlabel metal2 1402 -851 1402 -851 0 net=7871
rlabel metal2 1430 -851 1430 -851 0 net=8677
rlabel metal2 170 -853 170 -853 0 net=2633
rlabel metal2 205 -853 205 -853 0 net=10491
rlabel metal2 170 -855 170 -855 0 net=2351
rlabel metal2 296 -855 296 -855 0 net=1806
rlabel metal2 646 -855 646 -855 0 net=7717
rlabel metal2 1272 -855 1272 -855 0 net=11142
rlabel metal2 184 -857 184 -857 0 net=4062
rlabel metal2 310 -857 310 -857 0 net=3128
rlabel metal2 422 -857 422 -857 0 net=3093
rlabel metal2 1139 -857 1139 -857 0 net=7486
rlabel metal2 1255 -857 1255 -857 0 net=8195
rlabel metal2 1360 -857 1360 -857 0 net=14506
rlabel metal2 184 -859 184 -859 0 net=4076
rlabel metal2 775 -859 775 -859 0 net=5659
rlabel metal2 1143 -859 1143 -859 0 net=11624
rlabel metal2 198 -861 198 -861 0 net=2397
rlabel metal2 310 -861 310 -861 0 net=2901
rlabel metal2 457 -861 457 -861 0 net=3791
rlabel metal2 562 -861 562 -861 0 net=3265
rlabel metal2 653 -861 653 -861 0 net=6651
rlabel metal2 1045 -861 1045 -861 0 net=6729
rlabel metal2 1101 -861 1101 -861 0 net=7243
rlabel metal2 1206 -861 1206 -861 0 net=7742
rlabel metal2 1969 -861 1969 -861 0 net=12241
rlabel metal2 2074 -861 2074 -861 0 net=13085
rlabel metal2 156 -863 156 -863 0 net=4639
rlabel metal2 205 -863 205 -863 0 net=2817
rlabel metal2 254 -863 254 -863 0 net=3109
rlabel metal2 527 -863 527 -863 0 net=8119
rlabel metal2 1209 -863 1209 -863 0 net=12996
rlabel metal2 2130 -863 2130 -863 0 net=13241
rlabel metal2 156 -865 156 -865 0 net=3321
rlabel metal2 478 -865 478 -865 0 net=2283
rlabel metal2 527 -865 527 -865 0 net=4882
rlabel metal2 828 -865 828 -865 0 net=3890
rlabel metal2 2004 -865 2004 -865 0 net=12667
rlabel metal2 2123 -865 2123 -865 0 net=14731
rlabel metal2 163 -867 163 -867 0 net=3019
rlabel metal2 478 -867 478 -867 0 net=3473
rlabel metal2 807 -867 807 -867 0 net=6543
rlabel metal2 1143 -867 1143 -867 0 net=6131
rlabel metal2 1220 -867 1220 -867 0 net=12632
rlabel metal2 2102 -867 2102 -867 0 net=12967
rlabel metal2 163 -869 163 -869 0 net=2957
rlabel metal2 359 -869 359 -869 0 net=6659
rlabel metal2 667 -869 667 -869 0 net=3891
rlabel metal2 187 -871 187 -871 0 net=11493
rlabel metal2 1787 -871 1787 -871 0 net=10933
rlabel metal2 2102 -871 2102 -871 0 net=13195
rlabel metal2 219 -873 219 -873 0 net=7861
rlabel metal2 957 -873 957 -873 0 net=12651
rlabel metal2 1556 -873 1556 -873 0 net=10013
rlabel metal2 1654 -873 1654 -873 0 net=10655
rlabel metal2 1787 -873 1787 -873 0 net=12701
rlabel metal2 2053 -873 2053 -873 0 net=12909
rlabel metal2 233 -875 233 -875 0 net=2391
rlabel metal2 317 -875 317 -875 0 net=3193
rlabel metal2 317 -875 317 -875 0 net=3193
rlabel metal2 324 -875 324 -875 0 net=2181
rlabel metal2 387 -875 387 -875 0 net=2981
rlabel metal2 492 -875 492 -875 0 net=3853
rlabel metal2 1024 -875 1024 -875 0 net=9229
rlabel metal2 1605 -875 1605 -875 0 net=10133
rlabel metal2 1682 -875 1682 -875 0 net=10153
rlabel metal2 1829 -875 1829 -875 0 net=11695
rlabel metal2 100 -877 100 -877 0 net=2368
rlabel metal2 408 -877 408 -877 0 net=3435
rlabel metal2 688 -877 688 -877 0 net=7314
rlabel metal2 737 -877 737 -877 0 net=6929
rlabel metal2 1055 -877 1055 -877 0 net=11804
rlabel metal2 100 -879 100 -879 0 net=1209
rlabel metal2 1080 -879 1080 -879 0 net=7079
rlabel metal2 1185 -879 1185 -879 0 net=7517
rlabel metal2 1871 -879 1871 -879 0 net=11445
rlabel metal2 121 -881 121 -881 0 net=3027
rlabel metal2 408 -881 408 -881 0 net=2539
rlabel metal2 436 -881 436 -881 0 net=2655
rlabel metal2 513 -881 513 -881 0 net=5784
rlabel metal2 723 -881 723 -881 0 net=6157
rlabel metal2 1146 -881 1146 -881 0 net=1111
rlabel metal2 1647 -881 1647 -881 0 net=10635
rlabel metal2 1745 -881 1745 -881 0 net=11255
rlabel metal2 1913 -881 1913 -881 0 net=12003
rlabel metal2 2081 -881 2081 -881 0 net=13109
rlabel metal2 2 -883 2 -883 0 net=2881
rlabel metal2 492 -883 492 -883 0 net=4155
rlabel metal2 1031 -883 1031 -883 0 net=5713
rlabel metal2 1157 -883 1157 -883 0 net=14362
rlabel metal2 2 -885 2 -885 0 net=8141
rlabel metal2 247 -885 247 -885 0 net=1843
rlabel metal2 359 -885 359 -885 0 net=2417
rlabel metal2 499 -885 499 -885 0 net=2769
rlabel metal2 534 -885 534 -885 0 net=3367
rlabel metal2 688 -885 688 -885 0 net=4261
rlabel metal2 737 -885 737 -885 0 net=5315
rlabel metal2 954 -885 954 -885 0 net=14759
rlabel metal2 65 -887 65 -887 0 net=12191
rlabel metal2 2144 -887 2144 -887 0 net=13287
rlabel metal2 65 -889 65 -889 0 net=4243
rlabel metal2 464 -889 464 -889 0 net=2121
rlabel metal2 541 -889 541 -889 0 net=4763
rlabel metal2 698 -889 698 -889 0 net=5184
rlabel metal2 1052 -889 1052 -889 0 net=6829
rlabel metal2 1157 -889 1157 -889 0 net=7277
rlabel metal2 1213 -889 1213 -889 0 net=13828
rlabel metal2 86 -891 86 -891 0 net=2599
rlabel metal2 401 -891 401 -891 0 net=4589
rlabel metal2 513 -891 513 -891 0 net=4973
rlabel metal2 702 -891 702 -891 0 net=8320
rlabel metal2 1199 -891 1199 -891 0 net=7569
rlabel metal2 1286 -891 1286 -891 0 net=9729
rlabel metal2 1682 -891 1682 -891 0 net=10203
rlabel metal2 1738 -891 1738 -891 0 net=11407
rlabel metal2 2172 -891 2172 -891 0 net=13525
rlabel metal2 2207 -891 2207 -891 0 net=13583
rlabel metal2 86 -893 86 -893 0 net=4785
rlabel metal2 380 -893 380 -893 0 net=4109
rlabel metal2 702 -893 702 -893 0 net=4937
rlabel metal2 905 -893 905 -893 0 net=5428
rlabel metal2 1125 -893 1125 -893 0 net=11577
rlabel metal2 2193 -893 2193 -893 0 net=14073
rlabel metal2 107 -895 107 -895 0 net=6717
rlabel metal2 919 -895 919 -895 0 net=6685
rlabel metal2 1164 -895 1164 -895 0 net=7691
rlabel metal2 1290 -895 1290 -895 0 net=7767
rlabel metal2 1395 -895 1395 -895 0 net=9181
rlabel metal2 1766 -895 1766 -895 0 net=14653
rlabel metal2 107 -897 107 -897 0 net=2515
rlabel metal2 247 -897 247 -897 0 net=6005
rlabel metal2 1038 -897 1038 -897 0 net=6173
rlabel metal2 1171 -897 1171 -897 0 net=13504
rlabel metal2 2207 -897 2207 -897 0 net=14299
rlabel metal2 51 -899 51 -899 0 net=4081
rlabel metal2 261 -899 261 -899 0 net=10901
rlabel metal2 765 -899 765 -899 0 net=5295
rlabel metal2 1192 -899 1192 -899 0 net=8979
rlabel metal2 1290 -899 1290 -899 0 net=8185
rlabel metal2 1353 -899 1353 -899 0 net=9583
rlabel metal2 1794 -899 1794 -899 0 net=10981
rlabel metal2 1892 -899 1892 -899 0 net=13769
rlabel metal2 51 -901 51 -901 0 net=5319
rlabel metal2 639 -901 639 -901 0 net=10185
rlabel metal2 2018 -901 2018 -901 0 net=12429
rlabel metal2 124 -903 124 -903 0 net=11883
rlabel metal2 1794 -903 1794 -903 0 net=11663
rlabel metal2 2018 -903 2018 -903 0 net=12795
rlabel metal2 2186 -903 2186 -903 0 net=13485
rlabel metal2 149 -905 149 -905 0 net=2927
rlabel metal2 541 -905 541 -905 0 net=4331
rlabel metal2 618 -905 618 -905 0 net=3770
rlabel metal2 786 -905 786 -905 0 net=7317
rlabel metal2 1213 -905 1213 -905 0 net=7879
rlabel metal2 1304 -905 1304 -905 0 net=7935
rlabel metal2 30 -907 30 -907 0 net=6439
rlabel metal2 796 -907 796 -907 0 net=3915
rlabel metal2 1220 -907 1220 -907 0 net=7219
rlabel metal2 1241 -907 1241 -907 0 net=11008
rlabel metal2 1843 -907 1843 -907 0 net=12601
rlabel metal2 2067 -907 2067 -907 0 net=13009
rlabel metal2 2200 -907 2200 -907 0 net=14189
rlabel metal2 30 -909 30 -909 0 net=3595
rlabel metal2 180 -909 180 -909 0 net=5167
rlabel metal2 716 -909 716 -909 0 net=11543
rlabel metal2 1906 -909 1906 -909 0 net=11959
rlabel metal2 2039 -909 2039 -909 0 net=14483
rlabel metal2 135 -911 135 -911 0 net=13217
rlabel metal2 2214 -911 2214 -911 0 net=13725
rlabel metal2 149 -913 149 -913 0 net=1553
rlabel metal2 1223 -913 1223 -913 0 net=14275
rlabel metal2 1955 -913 1955 -913 0 net=12165
rlabel metal2 2214 -913 2214 -913 0 net=14311
rlabel metal2 226 -915 226 -915 0 net=4227
rlabel metal2 814 -915 814 -915 0 net=5878
rlabel metal2 1325 -915 1325 -915 0 net=8605
rlabel metal2 1535 -915 1535 -915 0 net=13867
rlabel metal2 2270 -915 2270 -915 0 net=14563
rlabel metal2 226 -917 226 -917 0 net=1513
rlabel metal2 1178 -917 1178 -917 0 net=9007
rlabel metal2 1493 -917 1493 -917 0 net=7385
rlabel metal2 23 -919 23 -919 0 net=5979
rlabel metal2 1122 -919 1122 -919 0 net=7405
rlabel metal2 1227 -919 1227 -919 0 net=7629
rlabel metal2 1304 -919 1304 -919 0 net=8741
rlabel metal2 1493 -919 1493 -919 0 net=9273
rlabel metal2 1584 -919 1584 -919 0 net=9921
rlabel metal2 1997 -919 1997 -919 0 net=12515
rlabel metal2 23 -921 23 -921 0 net=3635
rlabel metal2 268 -921 268 -921 0 net=14163
rlabel metal2 114 -923 114 -923 0 net=4997
rlabel metal2 593 -923 593 -923 0 net=188
rlabel metal2 1234 -923 1234 -923 0 net=8699
rlabel metal2 1535 -923 1535 -923 0 net=9785
rlabel metal2 1633 -923 1633 -923 0 net=10297
rlabel metal2 1857 -923 1857 -923 0 net=11359
rlabel metal2 275 -925 275 -925 0 net=1619
rlabel metal2 345 -925 345 -925 0 net=3677
rlabel metal2 1262 -925 1262 -925 0 net=8509
rlabel metal2 1311 -925 1311 -925 0 net=14639
rlabel metal2 275 -927 275 -927 0 net=1983
rlabel metal2 485 -927 485 -927 0 net=3515
rlabel metal2 597 -927 597 -927 0 net=3501
rlabel metal2 684 -927 684 -927 0 net=8583
rlabel metal2 1339 -927 1339 -927 0 net=9237
rlabel metal2 1549 -927 1549 -927 0 net=9347
rlabel metal2 1612 -927 1612 -927 0 net=9845
rlabel metal2 1710 -927 1710 -927 0 net=11125
rlabel metal2 1857 -927 1857 -927 0 net=12893
rlabel metal2 345 -929 345 -929 0 net=2333
rlabel metal2 1283 -929 1283 -929 0 net=10745
rlabel metal2 1563 -929 1563 -929 0 net=10107
rlabel metal2 1822 -929 1822 -929 0 net=11199
rlabel metal2 1885 -929 1885 -929 0 net=11897
rlabel metal2 19 -931 19 -931 0 net=11773
rlabel metal2 331 -933 331 -933 0 net=3129
rlabel metal2 1339 -933 1339 -933 0 net=8755
rlabel metal2 1500 -933 1500 -933 0 net=9037
rlabel metal2 366 -935 366 -935 0 net=4515
rlabel metal2 1500 -935 1500 -935 0 net=9479
rlabel metal2 1619 -935 1619 -935 0 net=10453
rlabel metal2 401 -937 401 -937 0 net=3825
rlabel metal2 1059 -937 1059 -937 0 net=12141
rlabel metal2 187 -939 187 -939 0 net=6211
rlabel metal2 1318 -939 1318 -939 0 net=8009
rlabel metal2 1577 -939 1577 -939 0 net=12349
rlabel metal2 429 -941 429 -941 0 net=2689
rlabel metal2 1318 -941 1318 -941 0 net=9117
rlabel metal2 1724 -941 1724 -941 0 net=11319
rlabel metal2 604 -943 604 -943 0 net=5099
rlabel metal2 1346 -943 1346 -943 0 net=7261
rlabel metal2 1507 -943 1507 -943 0 net=9665
rlabel metal2 1850 -943 1850 -943 0 net=11823
rlabel metal2 660 -945 660 -945 0 net=3863
rlabel metal2 1360 -945 1360 -945 0 net=8377
rlabel metal2 1591 -945 1591 -945 0 net=10179
rlabel metal2 1927 -945 1927 -945 0 net=12037
rlabel metal2 744 -947 744 -947 0 net=10673
rlabel metal2 1976 -947 1976 -947 0 net=12415
rlabel metal2 744 -949 744 -949 0 net=5079
rlabel metal2 842 -949 842 -949 0 net=5601
rlabel metal2 1363 -949 1363 -949 0 net=13329
rlabel metal2 555 -951 555 -951 0 net=3707
rlabel metal2 1367 -951 1367 -951 0 net=10666
rlabel metal2 1920 -951 1920 -951 0 net=12761
rlabel metal2 793 -953 793 -953 0 net=6862
rlabel metal2 1017 -953 1017 -953 0 net=11465
rlabel metal2 856 -955 856 -955 0 net=5529
rlabel metal2 961 -955 961 -955 0 net=5855
rlabel metal2 1367 -955 1367 -955 0 net=8827
rlabel metal2 856 -957 856 -957 0 net=5331
rlabel metal2 982 -957 982 -957 0 net=6491
rlabel metal2 1370 -957 1370 -957 0 net=13427
rlabel metal2 471 -959 471 -959 0 net=6065
rlabel metal2 1374 -959 1374 -959 0 net=12025
rlabel metal2 471 -961 471 -961 0 net=3667
rlabel metal2 586 -961 586 -961 0 net=7085
rlabel metal2 1374 -961 1374 -961 0 net=8969
rlabel metal2 576 -963 576 -963 0 net=3813
rlabel metal2 1381 -963 1381 -963 0 net=8993
rlabel metal2 625 -965 625 -965 0 net=12903
rlabel metal2 1458 -967 1458 -967 0 net=9255
rlabel metal2 1479 -969 1479 -969 0 net=9405
rlabel metal2 1486 -971 1486 -971 0 net=10527
rlabel metal2 1465 -973 1465 -973 0 net=8897
rlabel metal2 1465 -975 1465 -975 0 net=8905
rlabel metal2 1542 -975 1542 -975 0 net=9943
rlabel metal2 1073 -977 1073 -977 0 net=9327
rlabel metal2 1514 -977 1514 -977 0 net=10073
rlabel metal2 779 -979 779 -979 0 net=7031
rlabel metal2 1514 -979 1514 -979 0 net=14531
rlabel metal2 1570 -981 1570 -981 0 net=12138
rlabel metal2 751 -983 751 -983 0 net=10839
rlabel metal2 37 -985 37 -985 0 net=7337
rlabel metal2 37 -987 37 -987 0 net=5819
rlabel metal2 975 -989 975 -989 0 net=6997
rlabel metal2 730 -991 730 -991 0 net=4495
rlabel metal2 730 -993 730 -993 0 net=5217
rlabel metal2 338 -995 338 -995 0 net=5949
rlabel metal2 338 -997 338 -997 0 net=2319
rlabel metal2 9 -1008 9 -1008 0 net=1828
rlabel metal2 772 -1008 772 -1008 0 net=12968
rlabel metal2 2284 -1008 2284 -1008 0 net=14641
rlabel metal2 2375 -1008 2375 -1008 0 net=12551
rlabel metal2 9 -1010 9 -1010 0 net=4471
rlabel metal2 93 -1010 93 -1010 0 net=13726
rlabel metal2 2298 -1010 2298 -1010 0 net=14761
rlabel metal2 2382 -1010 2382 -1010 0 net=6243
rlabel metal2 2403 -1010 2403 -1010 0 net=14219
rlabel metal2 16 -1012 16 -1012 0 net=8081
rlabel metal2 93 -1012 93 -1012 0 net=5603
rlabel metal2 884 -1012 884 -1012 0 net=3917
rlabel metal2 936 -1012 936 -1012 0 net=7768
rlabel metal2 1409 -1012 1409 -1012 0 net=7873
rlabel metal2 1409 -1012 1409 -1012 0 net=7873
rlabel metal2 1507 -1012 1507 -1012 0 net=9667
rlabel metal2 1703 -1012 1703 -1012 0 net=14277
rlabel metal2 2368 -1012 2368 -1012 0 net=8935
rlabel metal2 2417 -1012 2417 -1012 0 net=14043
rlabel metal2 16 -1014 16 -1014 0 net=3131
rlabel metal2 345 -1014 345 -1014 0 net=2334
rlabel metal2 1020 -1014 1020 -1014 0 net=13486
rlabel metal2 103 -1016 103 -1016 0 net=4496
rlabel metal2 1174 -1016 1174 -1016 0 net=10982
rlabel metal2 2123 -1016 2123 -1016 0 net=14733
rlabel metal2 110 -1018 110 -1018 0 net=3194
rlabel metal2 324 -1018 324 -1018 0 net=2183
rlabel metal2 345 -1018 345 -1018 0 net=2983
rlabel metal2 590 -1018 590 -1018 0 net=3204
rlabel metal2 646 -1018 646 -1018 0 net=7718
rlabel metal2 964 -1018 964 -1018 0 net=13584
rlabel metal2 117 -1020 117 -1020 0 net=8010
rlabel metal2 1514 -1020 1514 -1020 0 net=10204
rlabel metal2 1689 -1020 1689 -1020 0 net=10675
rlabel metal2 1787 -1020 1787 -1020 0 net=12703
rlabel metal2 2165 -1020 2165 -1020 0 net=13429
rlabel metal2 128 -1022 128 -1022 0 net=4758
rlabel metal2 793 -1022 793 -1022 0 net=5660
rlabel metal2 1122 -1022 1122 -1022 0 net=8378
rlabel metal2 1514 -1022 1514 -1022 0 net=9787
rlabel metal2 1570 -1022 1570 -1022 0 net=9595
rlabel metal2 1570 -1022 1570 -1022 0 net=9595
rlabel metal2 1710 -1022 1710 -1022 0 net=11127
rlabel metal2 1801 -1022 1801 -1022 0 net=10492
rlabel metal2 128 -1024 128 -1024 0 net=10903
rlabel metal2 268 -1024 268 -1024 0 net=3475
rlabel metal2 590 -1024 590 -1024 0 net=3892
rlabel metal2 733 -1024 733 -1024 0 net=14164
rlabel metal2 86 -1026 86 -1026 0 net=4787
rlabel metal2 779 -1026 779 -1026 0 net=11660
rlabel metal2 2102 -1026 2102 -1026 0 net=13197
rlabel metal2 86 -1028 86 -1028 0 net=901
rlabel metal2 138 -1028 138 -1028 0 net=10186
rlabel metal2 1962 -1028 1962 -1028 0 net=12193
rlabel metal2 2172 -1028 2172 -1028 0 net=13527
rlabel metal2 135 -1030 135 -1030 0 net=11200
rlabel metal2 1836 -1030 1836 -1030 0 net=11775
rlabel metal2 1962 -1030 1962 -1030 0 net=12797
rlabel metal2 2130 -1030 2130 -1030 0 net=13243
rlabel metal2 177 -1032 177 -1032 0 net=12904
rlabel metal2 23 -1034 23 -1034 0 net=3637
rlabel metal2 180 -1034 180 -1034 0 net=4590
rlabel metal2 478 -1034 478 -1034 0 net=3517
rlabel metal2 611 -1034 611 -1034 0 net=10840
rlabel metal2 23 -1036 23 -1036 0 net=5683
rlabel metal2 100 -1036 100 -1036 0 net=14457
rlabel metal2 44 -1038 44 -1038 0 net=4083
rlabel metal2 261 -1038 261 -1038 0 net=1985
rlabel metal2 310 -1038 310 -1038 0 net=2902
rlabel metal2 919 -1038 919 -1038 0 net=6687
rlabel metal2 919 -1038 919 -1038 0 net=6687
rlabel metal2 940 -1038 940 -1038 0 net=4780
rlabel metal2 1024 -1038 1024 -1038 0 net=9231
rlabel metal2 1517 -1038 1517 -1038 0 net=13770
rlabel metal2 184 -1040 184 -1040 0 net=3111
rlabel metal2 271 -1040 271 -1040 0 net=4831
rlabel metal2 793 -1040 793 -1040 0 net=5333
rlabel metal2 863 -1040 863 -1040 0 net=5951
rlabel metal2 891 -1040 891 -1040 0 net=6067
rlabel metal2 975 -1040 975 -1040 0 net=6999
rlabel metal2 1125 -1040 1125 -1040 0 net=11446
rlabel metal2 2158 -1040 2158 -1040 0 net=13331
rlabel metal2 138 -1042 138 -1042 0 net=13179
rlabel metal2 187 -1044 187 -1044 0 net=10380
rlabel metal2 191 -1046 191 -1046 0 net=2635
rlabel metal2 324 -1046 324 -1046 0 net=4433
rlabel metal2 723 -1046 723 -1046 0 net=6159
rlabel metal2 989 -1046 989 -1046 0 net=6036
rlabel metal2 1041 -1046 1041 -1046 0 net=12273
rlabel metal2 2067 -1046 2067 -1046 0 net=13011
rlabel metal2 2200 -1046 2200 -1046 0 net=14191
rlabel metal2 170 -1048 170 -1048 0 net=2353
rlabel metal2 205 -1048 205 -1048 0 net=2819
rlabel metal2 366 -1048 366 -1048 0 net=4517
rlabel metal2 625 -1048 625 -1048 0 net=8898
rlabel metal2 1738 -1048 1738 -1048 0 net=11409
rlabel metal2 1843 -1048 1843 -1048 0 net=12603
rlabel metal2 2200 -1048 2200 -1048 0 net=14533
rlabel metal2 121 -1050 121 -1050 0 net=3029
rlabel metal2 219 -1050 219 -1050 0 net=6653
rlabel metal2 660 -1050 660 -1050 0 net=3865
rlabel metal2 730 -1050 730 -1050 0 net=5219
rlabel metal2 863 -1050 863 -1050 0 net=11413
rlabel metal2 1710 -1050 1710 -1050 0 net=7989
rlabel metal2 121 -1052 121 -1052 0 net=2419
rlabel metal2 366 -1052 366 -1052 0 net=2857
rlabel metal2 1181 -1052 1181 -1052 0 net=10036
rlabel metal2 1745 -1052 1745 -1052 0 net=11257
rlabel metal2 1843 -1052 1843 -1052 0 net=11825
rlabel metal2 1864 -1052 1864 -1052 0 net=11579
rlabel metal2 2186 -1052 2186 -1052 0 net=13869
rlabel metal2 145 -1054 145 -1054 0 net=62
rlabel metal2 796 -1054 796 -1054 0 net=5530
rlabel metal2 996 -1054 996 -1054 0 net=6358
rlabel metal2 1234 -1054 1234 -1054 0 net=8701
rlabel metal2 1437 -1054 1437 -1054 0 net=10747
rlabel metal2 1815 -1054 1815 -1054 0 net=11569
rlabel metal2 1871 -1054 1871 -1054 0 net=11961
rlabel metal2 1983 -1054 1983 -1054 0 net=12507
rlabel metal2 170 -1056 170 -1056 0 net=2449
rlabel metal2 380 -1056 380 -1056 0 net=4110
rlabel metal2 817 -1056 817 -1056 0 net=9038
rlabel metal2 1675 -1056 1675 -1056 0 net=11885
rlabel metal2 1955 -1056 1955 -1056 0 net=12167
rlabel metal2 2004 -1056 2004 -1056 0 net=12669
rlabel metal2 2186 -1056 2186 -1056 0 net=13303
rlabel metal2 79 -1058 79 -1058 0 net=3087
rlabel metal2 387 -1058 387 -1058 0 net=2641
rlabel metal2 831 -1058 831 -1058 0 net=11360
rlabel metal2 2039 -1058 2039 -1058 0 net=14485
rlabel metal2 79 -1060 79 -1060 0 net=4999
rlabel metal2 222 -1060 222 -1060 0 net=3678
rlabel metal2 639 -1060 639 -1060 0 net=4229
rlabel metal2 775 -1060 775 -1060 0 net=3854
rlabel metal2 982 -1060 982 -1060 0 net=6493
rlabel metal2 1003 -1060 1003 -1060 0 net=7087
rlabel metal2 1192 -1060 1192 -1060 0 net=8678
rlabel metal2 30 -1062 30 -1062 0 net=3597
rlabel metal2 646 -1062 646 -1062 0 net=5169
rlabel metal2 835 -1062 835 -1062 0 net=7319
rlabel metal2 1136 -1062 1136 -1062 0 net=7377
rlabel metal2 1157 -1062 1157 -1062 0 net=7279
rlabel metal2 1234 -1062 1234 -1062 0 net=11515
rlabel metal2 1878 -1062 1878 -1062 0 net=11859
rlabel metal2 30 -1064 30 -1064 0 net=8873
rlabel metal2 835 -1064 835 -1064 0 net=5791
rlabel metal2 968 -1064 968 -1064 0 net=7033
rlabel metal2 1129 -1064 1129 -1064 0 net=7442
rlabel metal2 1237 -1064 1237 -1064 0 net=8186
rlabel metal2 1307 -1064 1307 -1064 0 net=12221
rlabel metal2 2011 -1064 2011 -1064 0 net=12763
rlabel metal2 65 -1066 65 -1066 0 net=4245
rlabel metal2 660 -1066 660 -1066 0 net=6931
rlabel metal2 842 -1066 842 -1066 0 net=4565
rlabel metal2 877 -1066 877 -1066 0 net=5981
rlabel metal2 947 -1066 947 -1066 0 net=14049
rlabel metal2 65 -1068 65 -1068 0 net=3669
rlabel metal2 485 -1068 485 -1068 0 net=2123
rlabel metal2 597 -1068 597 -1068 0 net=3503
rlabel metal2 635 -1068 635 -1068 0 net=6671
rlabel metal2 1087 -1068 1087 -1068 0 net=6297
rlabel metal2 1136 -1068 1136 -1068 0 net=9329
rlabel metal2 1479 -1068 1479 -1068 0 net=9407
rlabel metal2 1542 -1068 1542 -1068 0 net=9945
rlabel metal2 1633 -1068 1633 -1068 0 net=10299
rlabel metal2 1815 -1068 1815 -1068 0 net=11157
rlabel metal2 226 -1070 226 -1070 0 net=1515
rlabel metal2 513 -1070 513 -1070 0 net=4975
rlabel metal2 891 -1070 891 -1070 0 net=5401
rlabel metal2 1003 -1070 1003 -1070 0 net=6363
rlabel metal2 1045 -1070 1045 -1070 0 net=6731
rlabel metal2 1241 -1070 1241 -1070 0 net=10934
rlabel metal2 51 -1072 51 -1072 0 net=5321
rlabel metal2 534 -1072 534 -1072 0 net=2083
rlabel metal2 1272 -1072 1272 -1072 0 net=12387
rlabel metal2 2039 -1072 2039 -1072 0 net=12359
rlabel metal2 51 -1074 51 -1074 0 net=6137
rlabel metal2 212 -1074 212 -1074 0 net=2493
rlabel metal2 240 -1074 240 -1074 0 net=3245
rlabel metal2 597 -1074 597 -1074 0 net=5809
rlabel metal2 1223 -1074 1223 -1074 0 net=7621
rlabel metal2 1244 -1074 1244 -1074 0 net=14237
rlabel metal2 142 -1076 142 -1076 0 net=6909
rlabel metal2 1010 -1076 1010 -1076 0 net=6611
rlabel metal2 1055 -1076 1055 -1076 0 net=9348
rlabel metal2 1598 -1076 1598 -1076 0 net=10351
rlabel metal2 1829 -1076 1829 -1076 0 net=11697
rlabel metal2 1878 -1076 1878 -1076 0 net=12039
rlabel metal2 1941 -1076 1941 -1076 0 net=12087
rlabel metal2 1969 -1076 1969 -1076 0 net=12243
rlabel metal2 2207 -1076 2207 -1076 0 net=14301
rlabel metal2 198 -1078 198 -1078 0 net=4641
rlabel metal2 254 -1078 254 -1078 0 net=4333
rlabel metal2 681 -1078 681 -1078 0 net=3069
rlabel metal2 1017 -1078 1017 -1078 0 net=6175
rlabel metal2 1248 -1078 1248 -1078 0 net=8429
rlabel metal2 1374 -1078 1374 -1078 0 net=8971
rlabel metal2 1486 -1078 1486 -1078 0 net=10529
rlabel metal2 1927 -1078 1927 -1078 0 net=14075
rlabel metal2 198 -1080 198 -1080 0 net=6545
rlabel metal2 877 -1080 877 -1080 0 net=7753
rlabel metal2 1283 -1080 1283 -1080 0 net=12430
rlabel metal2 275 -1082 275 -1082 0 net=2883
rlabel metal2 429 -1082 429 -1082 0 net=2690
rlabel metal2 1500 -1082 1500 -1082 0 net=9481
rlabel metal2 1580 -1082 1580 -1082 0 net=11881
rlabel metal2 1997 -1082 1997 -1082 0 net=12517
rlabel metal2 2109 -1082 2109 -1082 0 net=13207
rlabel metal2 2235 -1082 2235 -1082 0 net=14367
rlabel metal2 359 -1084 359 -1084 0 net=5829
rlabel metal2 443 -1084 443 -1084 0 net=2771
rlabel metal2 541 -1084 541 -1084 0 net=5101
rlabel metal2 607 -1084 607 -1084 0 net=13315
rlabel metal2 114 -1086 114 -1086 0 net=4365
rlabel metal2 604 -1086 604 -1086 0 net=854
rlabel metal2 1059 -1086 1059 -1086 0 net=6133
rlabel metal2 1227 -1086 1227 -1086 0 net=7631
rlabel metal2 1286 -1086 1286 -1086 0 net=10154
rlabel metal2 1808 -1086 1808 -1086 0 net=11545
rlabel metal2 2151 -1086 2151 -1086 0 net=13301
rlabel metal2 401 -1088 401 -1088 0 net=3827
rlabel metal2 415 -1088 415 -1088 0 net=2657
rlabel metal2 695 -1088 695 -1088 0 net=6213
rlabel metal2 1080 -1088 1080 -1088 0 net=7081
rlabel metal2 1213 -1088 1213 -1088 0 net=7881
rlabel metal2 1314 -1088 1314 -1088 0 net=10074
rlabel metal2 1654 -1088 1654 -1088 0 net=10657
rlabel metal2 1857 -1088 1857 -1088 0 net=12895
rlabel metal2 401 -1090 401 -1090 0 net=2541
rlabel metal2 429 -1090 429 -1090 0 net=10426
rlabel metal2 1794 -1090 1794 -1090 0 net=11665
rlabel metal2 2095 -1090 2095 -1090 0 net=13161
rlabel metal2 408 -1092 408 -1092 0 net=3815
rlabel metal2 688 -1092 688 -1092 0 net=4263
rlabel metal2 702 -1092 702 -1092 0 net=4939
rlabel metal2 898 -1092 898 -1092 0 net=5471
rlabel metal2 1101 -1092 1101 -1092 0 net=7245
rlabel metal2 1213 -1092 1213 -1092 0 net=9691
rlabel metal2 2 -1094 2 -1094 0 net=8143
rlabel metal2 709 -1094 709 -1094 0 net=7253
rlabel metal2 1031 -1094 1031 -1094 0 net=5715
rlabel metal2 1318 -1094 1318 -1094 0 net=9119
rlabel metal2 1556 -1094 1556 -1094 0 net=10015
rlabel metal2 1696 -1094 1696 -1094 0 net=10867
rlabel metal2 2025 -1094 2025 -1094 0 net=12845
rlabel metal2 72 -1096 72 -1096 0 net=4807
rlabel metal2 737 -1096 737 -1096 0 net=5317
rlabel metal2 1325 -1096 1325 -1096 0 net=8607
rlabel metal2 1381 -1096 1381 -1096 0 net=8995
rlabel metal2 1598 -1096 1598 -1096 0 net=10135
rlabel metal2 1717 -1096 1717 -1096 0 net=10997
rlabel metal2 1899 -1096 1899 -1096 0 net=12351
rlabel metal2 37 -1098 37 -1098 0 net=5821
rlabel metal2 89 -1098 89 -1098 0 net=8159
rlabel metal2 1185 -1098 1185 -1098 0 net=7519
rlabel metal2 1717 -1098 1717 -1098 0 net=11467
rlabel metal2 1899 -1098 1899 -1098 0 net=10091
rlabel metal2 37 -1100 37 -1100 0 net=5051
rlabel metal2 751 -1100 751 -1100 0 net=7339
rlabel metal2 905 -1100 905 -1100 0 net=6719
rlabel metal2 1066 -1100 1066 -1100 0 net=6831
rlabel metal2 1185 -1100 1185 -1100 0 net=7571
rlabel metal2 1206 -1100 1206 -1100 0 net=8121
rlabel metal2 1335 -1100 1335 -1100 0 net=7386
rlabel metal2 247 -1102 247 -1102 0 net=6007
rlabel metal2 961 -1102 961 -1102 0 net=5857
rlabel metal2 1178 -1102 1178 -1102 0 net=7407
rlabel metal2 1255 -1102 1255 -1102 0 net=8197
rlabel metal2 1367 -1102 1367 -1102 0 net=8829
rlabel metal2 1395 -1102 1395 -1102 0 net=10821
rlabel metal2 2214 -1102 2214 -1102 0 net=14313
rlabel metal2 163 -1104 163 -1104 0 net=2959
rlabel metal2 373 -1104 373 -1104 0 net=164
rlabel metal2 1195 -1104 1195 -1104 0 net=9501
rlabel metal2 1724 -1104 1724 -1104 0 net=11321
rlabel metal2 2116 -1104 2116 -1104 0 net=13219
rlabel metal2 2270 -1104 2270 -1104 0 net=14565
rlabel metal2 163 -1106 163 -1106 0 net=2321
rlabel metal2 352 -1106 352 -1106 0 net=3167
rlabel metal2 390 -1106 390 -1106 0 net=5895
rlabel metal2 772 -1106 772 -1106 0 net=9957
rlabel metal2 2053 -1106 2053 -1106 0 net=12911
rlabel metal2 233 -1108 233 -1108 0 net=2392
rlabel metal2 1052 -1108 1052 -1108 0 net=11219
rlabel metal2 2053 -1108 2053 -1108 0 net=12283
rlabel metal2 233 -1110 233 -1110 0 net=2601
rlabel metal2 450 -1110 450 -1110 0 net=3021
rlabel metal2 506 -1110 506 -1110 0 net=10545
rlabel metal2 107 -1112 107 -1112 0 net=2517
rlabel metal2 450 -1112 450 -1112 0 net=4157
rlabel metal2 548 -1112 548 -1112 0 net=3437
rlabel metal2 674 -1112 674 -1112 0 net=4765
rlabel metal2 786 -1112 786 -1112 0 net=6441
rlabel metal2 1199 -1112 1199 -1112 0 net=14654
rlabel metal2 107 -1114 107 -1114 0 net=14326
rlabel metal2 338 -1116 338 -1116 0 net=2285
rlabel metal2 569 -1116 569 -1116 0 net=6661
rlabel metal2 1220 -1116 1220 -1116 0 net=7221
rlabel metal2 1262 -1116 1262 -1116 0 net=8511
rlabel metal2 1402 -1116 1402 -1116 0 net=12653
rlabel metal2 352 -1118 352 -1118 0 net=4347
rlabel metal2 905 -1118 905 -1118 0 net=10557
rlabel metal2 1766 -1118 1766 -1118 0 net=11495
rlabel metal2 422 -1120 422 -1120 0 net=3095
rlabel metal2 674 -1120 674 -1120 0 net=3625
rlabel metal2 1220 -1120 1220 -1120 0 net=13509
rlabel metal2 100 -1122 100 -1122 0 net=8497
rlabel metal2 436 -1122 436 -1122 0 net=2929
rlabel metal2 520 -1122 520 -1122 0 net=3369
rlabel metal2 744 -1122 744 -1122 0 net=5081
rlabel metal2 800 -1122 800 -1122 0 net=7863
rlabel metal2 1297 -1122 1297 -1122 0 net=8585
rlabel metal2 1423 -1122 1423 -1122 0 net=9161
rlabel metal2 1549 -1122 1549 -1122 0 net=10761
rlabel metal2 1661 -1122 1661 -1122 0 net=11069
rlabel metal2 289 -1124 289 -1124 0 net=2399
rlabel metal2 800 -1124 800 -1124 0 net=4213
rlabel metal2 1164 -1124 1164 -1124 0 net=7693
rlabel metal2 1297 -1124 1297 -1124 0 net=7937
rlabel metal2 289 -1126 289 -1126 0 net=1621
rlabel metal2 436 -1126 436 -1126 0 net=2691
rlabel metal2 821 -1126 821 -1126 0 net=12139
rlabel metal2 296 -1128 296 -1128 0 net=1845
rlabel metal2 457 -1128 457 -1128 0 net=3793
rlabel metal2 555 -1128 555 -1128 0 net=3709
rlabel metal2 1164 -1128 1164 -1128 0 net=9846
rlabel metal2 1619 -1128 1619 -1128 0 net=10455
rlabel metal2 282 -1130 282 -1130 0 net=2423
rlabel metal2 555 -1130 555 -1130 0 net=3267
rlabel metal2 1304 -1130 1304 -1130 0 net=8743
rlabel metal2 1416 -1130 1416 -1130 0 net=9009
rlabel metal2 1430 -1130 1430 -1130 0 net=9183
rlabel metal2 1584 -1130 1584 -1130 0 net=9923
rlabel metal2 149 -1132 149 -1132 0 net=1555
rlabel metal2 1304 -1132 1304 -1132 0 net=11838
rlabel metal2 149 -1134 149 -1134 0 net=6973
rlabel metal2 1311 -1134 1311 -1134 0 net=14491
rlabel metal2 156 -1136 156 -1136 0 net=3323
rlabel metal2 1311 -1136 1311 -1136 0 net=8757
rlabel metal2 1398 -1136 1398 -1136 0 net=14655
rlabel metal2 96 -1138 96 -1138 0 net=2041
rlabel metal2 824 -1138 824 -1138 0 net=8379
rlabel metal2 1430 -1138 1430 -1138 0 net=9711
rlabel metal2 1528 -1138 1528 -1138 0 net=9731
rlabel metal2 1591 -1138 1591 -1138 0 net=10181
rlabel metal2 1934 -1138 1934 -1138 0 net=13111
rlabel metal2 632 -1140 632 -1140 0 net=9851
rlabel metal2 2081 -1140 2081 -1140 0 net=13633
rlabel metal2 632 -1142 632 -1142 0 net=4381
rlabel metal2 1444 -1142 1444 -1142 0 net=9239
rlabel metal2 2144 -1142 2144 -1142 0 net=13289
rlabel metal2 1458 -1144 1458 -1144 0 net=9257
rlabel metal2 2074 -1144 2074 -1144 0 net=13087
rlabel metal2 1276 -1146 1276 -1146 0 net=8981
rlabel metal2 1493 -1146 1493 -1146 0 net=9275
rlabel metal2 1976 -1146 1976 -1146 0 net=12417
rlabel metal2 828 -1148 828 -1148 0 net=7837
rlabel metal2 1465 -1148 1465 -1148 0 net=8907
rlabel metal2 1948 -1148 1948 -1148 0 net=12143
rlabel metal2 765 -1150 765 -1150 0 net=5297
rlabel metal2 1465 -1150 1465 -1150 0 net=10637
rlabel metal2 1920 -1150 1920 -1150 0 net=12027
rlabel metal2 765 -1152 765 -1152 0 net=7189
rlabel metal2 1563 -1152 1563 -1152 0 net=10109
rlabel metal2 1913 -1152 1913 -1152 0 net=12005
rlabel metal2 849 -1154 849 -1154 0 net=8779
rlabel metal2 1885 -1154 1885 -1154 0 net=11899
rlabel metal2 1353 -1156 1353 -1156 0 net=9585
rlabel metal2 1741 -1156 1741 -1156 0 net=11755
rlabel metal2 1346 -1158 1346 -1158 0 net=7263
rlabel metal2 1332 -1160 1332 -1160 0 net=8633
rlabel metal2 957 -1162 957 -1162 0 net=1458
rlabel metal2 957 -1164 957 -1164 0 net=10141
rlabel metal2 5 -1175 5 -1175 0 net=709
rlabel metal2 485 -1175 485 -1175 0 net=2124
rlabel metal2 656 -1175 656 -1175 0 net=9788
rlabel metal2 1549 -1175 1549 -1175 0 net=13198
rlabel metal2 2298 -1175 2298 -1175 0 net=14279
rlabel metal2 19 -1177 19 -1177 0 net=8874
rlabel metal2 89 -1177 89 -1177 0 net=5220
rlabel metal2 866 -1177 866 -1177 0 net=6720
rlabel metal2 1041 -1177 1041 -1177 0 net=14209
rlabel metal2 23 -1179 23 -1179 0 net=5684
rlabel metal2 842 -1179 842 -1179 0 net=4567
rlabel metal2 880 -1179 880 -1179 0 net=10658
rlabel metal2 1906 -1179 1906 -1179 0 net=11887
rlabel metal2 23 -1181 23 -1181 0 net=4519
rlabel metal2 667 -1181 667 -1181 0 net=4789
rlabel metal2 905 -1181 905 -1181 0 net=6009
rlabel metal2 947 -1181 947 -1181 0 net=527
rlabel metal2 1447 -1181 1447 -1181 0 net=14486
rlabel metal2 2368 -1181 2368 -1181 0 net=14735
rlabel metal2 30 -1183 30 -1183 0 net=3103
rlabel metal2 751 -1183 751 -1183 0 net=4767
rlabel metal2 912 -1183 912 -1183 0 net=5983
rlabel metal2 1048 -1183 1048 -1183 0 net=7320
rlabel metal2 1157 -1183 1157 -1183 0 net=12508
rlabel metal2 2277 -1183 2277 -1183 0 net=14193
rlabel metal2 100 -1185 100 -1185 0 net=8498
rlabel metal2 947 -1185 947 -1185 0 net=8161
rlabel metal2 1104 -1185 1104 -1185 0 net=14613
rlabel metal2 100 -1187 100 -1187 0 net=2961
rlabel metal2 254 -1187 254 -1187 0 net=4335
rlabel metal2 950 -1187 950 -1187 0 net=9120
rlabel metal2 1458 -1187 1458 -1187 0 net=8983
rlabel metal2 1552 -1187 1552 -1187 0 net=10136
rlabel metal2 1605 -1187 1605 -1187 0 net=10763
rlabel metal2 1927 -1187 1927 -1187 0 net=14077
rlabel metal2 121 -1189 121 -1189 0 net=2420
rlabel metal2 513 -1189 513 -1189 0 net=5323
rlabel metal2 667 -1189 667 -1189 0 net=7755
rlabel metal2 1307 -1189 1307 -1189 0 net=1450
rlabel metal2 2431 -1189 2431 -1189 0 net=12553
rlabel metal2 124 -1191 124 -1191 0 net=5318
rlabel metal2 1335 -1191 1335 -1191 0 net=14302
rlabel metal2 2354 -1191 2354 -1191 0 net=14657
rlabel metal2 128 -1193 128 -1193 0 net=10905
rlabel metal2 1969 -1193 1969 -1193 0 net=11546
rlabel metal2 2438 -1193 2438 -1193 0 net=14221
rlabel metal2 128 -1195 128 -1195 0 net=3477
rlabel metal2 275 -1195 275 -1195 0 net=2884
rlabel metal2 796 -1195 796 -1195 0 net=7034
rlabel metal2 982 -1195 982 -1195 0 net=6215
rlabel metal2 1115 -1195 1115 -1195 0 net=7247
rlabel metal2 1339 -1195 1339 -1195 0 net=8381
rlabel metal2 1500 -1195 1500 -1195 0 net=9241
rlabel metal2 1605 -1195 1605 -1195 0 net=9925
rlabel metal2 1745 -1195 1745 -1195 0 net=11259
rlabel metal2 2060 -1195 2060 -1195 0 net=12655
rlabel metal2 2284 -1195 2284 -1195 0 net=14239
rlabel metal2 138 -1197 138 -1197 0 net=2400
rlabel metal2 590 -1197 590 -1197 0 net=11158
rlabel metal2 1857 -1197 1857 -1197 0 net=11667
rlabel metal2 2095 -1197 2095 -1197 0 net=12847
rlabel metal2 2305 -1197 2305 -1197 0 net=14315
rlabel metal2 208 -1199 208 -1199 0 net=56
rlabel metal2 751 -1199 751 -1199 0 net=5953
rlabel metal2 992 -1199 992 -1199 0 net=13969
rlabel metal2 37 -1201 37 -1201 0 net=5053
rlabel metal2 1003 -1201 1003 -1201 0 net=10530
rlabel metal2 1962 -1201 1962 -1201 0 net=12799
rlabel metal2 2312 -1201 2312 -1201 0 net=14369
rlabel metal2 37 -1203 37 -1203 0 net=4809
rlabel metal2 758 -1203 758 -1203 0 net=12121
rlabel metal2 1521 -1203 1521 -1203 0 net=9259
rlabel metal2 1668 -1203 1668 -1203 0 net=10353
rlabel metal2 2109 -1203 2109 -1203 0 net=12897
rlabel metal2 2319 -1203 2319 -1203 0 net=14459
rlabel metal2 268 -1205 268 -1205 0 net=14762
rlabel metal2 2424 -1205 2424 -1205 0 net=14045
rlabel metal2 275 -1207 275 -1207 0 net=1507
rlabel metal2 310 -1209 310 -1209 0 net=2637
rlabel metal2 1003 -1209 1003 -1209 0 net=13510
rlabel metal2 2333 -1209 2333 -1209 0 net=14567
rlabel metal2 72 -1211 72 -1211 0 net=5823
rlabel metal2 380 -1211 380 -1211 0 net=3089
rlabel metal2 436 -1211 436 -1211 0 net=2693
rlabel metal2 527 -1211 527 -1211 0 net=3247
rlabel metal2 604 -1211 604 -1211 0 net=7811
rlabel metal2 828 -1211 828 -1211 0 net=5299
rlabel metal2 1010 -1211 1010 -1211 0 net=6443
rlabel metal2 1164 -1211 1164 -1211 0 net=6244
rlabel metal2 72 -1213 72 -1213 0 net=2773
rlabel metal2 485 -1213 485 -1213 0 net=3795
rlabel metal2 555 -1213 555 -1213 0 net=3269
rlabel metal2 642 -1213 642 -1213 0 net=10647
rlabel metal2 1920 -1213 1920 -1213 0 net=12007
rlabel metal2 2116 -1213 2116 -1213 0 net=12913
rlabel metal2 2340 -1213 2340 -1213 0 net=14643
rlabel metal2 9 -1215 9 -1215 0 net=4473
rlabel metal2 569 -1215 569 -1215 0 net=3097
rlabel metal2 702 -1215 702 -1215 0 net=1861
rlabel metal2 1038 -1215 1038 -1215 0 net=6613
rlabel metal2 1167 -1215 1167 -1215 0 net=14765
rlabel metal2 9 -1217 9 -1217 0 net=5273
rlabel metal2 219 -1217 219 -1217 0 net=6655
rlabel metal2 1178 -1217 1178 -1217 0 net=11826
rlabel metal2 1934 -1217 1934 -1217 0 net=13113
rlabel metal2 16 -1219 16 -1219 0 net=3133
rlabel metal2 499 -1219 499 -1219 0 net=4367
rlabel metal2 758 -1219 758 -1219 0 net=5083
rlabel metal2 800 -1219 800 -1219 0 net=4214
rlabel metal2 1045 -1219 1045 -1219 0 net=6463
rlabel metal2 1185 -1219 1185 -1219 0 net=7573
rlabel metal2 1370 -1219 1370 -1219 0 net=12604
rlabel metal2 2116 -1219 2116 -1219 0 net=14051
rlabel metal2 65 -1221 65 -1221 0 net=3671
rlabel metal2 772 -1221 772 -1221 0 net=4501
rlabel metal2 772 -1221 772 -1221 0 net=4501
rlabel metal2 800 -1221 800 -1221 0 net=2781
rlabel metal2 1045 -1221 1045 -1221 0 net=5717
rlabel metal2 1192 -1221 1192 -1221 0 net=7281
rlabel metal2 1311 -1221 1311 -1221 0 net=8759
rlabel metal2 1563 -1221 1563 -1221 0 net=9587
rlabel metal2 65 -1223 65 -1223 0 net=5001
rlabel metal2 114 -1223 114 -1223 0 net=10221
rlabel metal2 2144 -1223 2144 -1223 0 net=13089
rlabel metal2 114 -1225 114 -1225 0 net=5171
rlabel metal2 807 -1225 807 -1225 0 net=4941
rlabel metal2 852 -1225 852 -1225 0 net=10163
rlabel metal2 1815 -1225 1815 -1225 0 net=11777
rlabel metal2 1948 -1225 1948 -1225 0 net=12029
rlabel metal2 2151 -1225 2151 -1225 0 net=13163
rlabel metal2 135 -1227 135 -1227 0 net=3071
rlabel metal2 789 -1227 789 -1227 0 net=11167
rlabel metal2 1955 -1227 1955 -1227 0 net=12089
rlabel metal2 2158 -1227 2158 -1227 0 net=13181
rlabel metal2 191 -1229 191 -1229 0 net=2355
rlabel metal2 373 -1229 373 -1229 0 net=3169
rlabel metal2 506 -1229 506 -1229 0 net=14059
rlabel metal2 191 -1231 191 -1231 0 net=2643
rlabel metal2 408 -1231 408 -1231 0 net=3816
rlabel metal2 646 -1231 646 -1231 0 net=6733
rlabel metal2 1192 -1231 1192 -1231 0 net=7695
rlabel metal2 1283 -1231 1283 -1231 0 net=7865
rlabel metal2 1570 -1231 1570 -1231 0 net=9597
rlabel metal2 1731 -1231 1731 -1231 0 net=10749
rlabel metal2 1955 -1231 1955 -1231 0 net=12671
rlabel metal2 2088 -1231 2088 -1231 0 net=12765
rlabel metal2 198 -1233 198 -1233 0 net=6547
rlabel metal2 1234 -1233 1234 -1233 0 net=13655
rlabel metal2 149 -1235 149 -1235 0 net=6975
rlabel metal2 1255 -1235 1255 -1235 0 net=7223
rlabel metal2 1283 -1235 1283 -1235 0 net=7265
rlabel metal2 1381 -1235 1381 -1235 0 net=8831
rlabel metal2 1416 -1235 1416 -1235 0 net=8781
rlabel metal2 1591 -1235 1591 -1235 0 net=9853
rlabel metal2 1738 -1235 1738 -1235 0 net=12963
rlabel metal2 145 -1237 145 -1237 0 net=6469
rlabel metal2 198 -1237 198 -1237 0 net=8431
rlabel metal2 1381 -1237 1381 -1237 0 net=10182
rlabel metal2 1633 -1237 1633 -1237 0 net=9959
rlabel metal2 1741 -1237 1741 -1237 0 net=11685
rlabel metal2 2172 -1237 2172 -1237 0 net=13245
rlabel metal2 233 -1239 233 -1239 0 net=2603
rlabel metal2 422 -1239 422 -1239 0 net=10546
rlabel metal2 1885 -1239 1885 -1239 0 net=11757
rlabel metal2 2179 -1239 2179 -1239 0 net=13291
rlabel metal2 226 -1241 226 -1241 0 net=2495
rlabel metal2 261 -1241 261 -1241 0 net=1987
rlabel metal2 436 -1241 436 -1241 0 net=3627
rlabel metal2 681 -1241 681 -1241 0 net=3711
rlabel metal2 807 -1241 807 -1241 0 net=5199
rlabel metal2 1332 -1241 1332 -1241 0 net=11293
rlabel metal2 1983 -1241 1983 -1241 0 net=12169
rlabel metal2 2186 -1241 2186 -1241 0 net=13305
rlabel metal2 261 -1243 261 -1243 0 net=1761
rlabel metal2 1059 -1243 1059 -1243 0 net=6134
rlabel metal2 1241 -1243 1241 -1243 0 net=7623
rlabel metal2 1384 -1243 1384 -1243 0 net=13208
rlabel metal2 2221 -1243 2221 -1243 0 net=13333
rlabel metal2 303 -1245 303 -1245 0 net=2425
rlabel metal2 380 -1245 380 -1245 0 net=3829
rlabel metal2 506 -1245 506 -1245 0 net=4231
rlabel metal2 744 -1245 744 -1245 0 net=6099
rlabel metal2 961 -1245 961 -1245 0 net=9367
rlabel metal2 1654 -1245 1654 -1245 0 net=10143
rlabel metal2 1990 -1245 1990 -1245 0 net=12195
rlabel metal2 2193 -1245 2193 -1245 0 net=13317
rlabel metal2 229 -1247 229 -1247 0 net=1995
rlabel metal2 527 -1247 527 -1247 0 net=3325
rlabel metal2 877 -1247 877 -1247 0 net=11869
rlabel metal2 2200 -1247 2200 -1247 0 net=14535
rlabel metal2 303 -1249 303 -1249 0 net=2085
rlabel metal2 548 -1249 548 -1249 0 net=2241
rlabel metal2 1206 -1249 1206 -1249 0 net=7409
rlabel metal2 1325 -1249 1325 -1249 0 net=8199
rlabel metal2 1416 -1249 1416 -1249 0 net=12704
rlabel metal2 2137 -1249 2137 -1249 0 net=11581
rlabel metal2 2228 -1249 2228 -1249 0 net=13431
rlabel metal2 331 -1251 331 -1251 0 net=2185
rlabel metal2 520 -1251 520 -1251 0 net=3371
rlabel metal2 562 -1251 562 -1251 0 net=3324
rlabel metal2 891 -1251 891 -1251 0 net=5403
rlabel metal2 975 -1251 975 -1251 0 net=6161
rlabel metal2 1073 -1251 1073 -1251 0 net=6673
rlabel metal2 1241 -1251 1241 -1251 0 net=7633
rlabel metal2 1255 -1251 1255 -1251 0 net=8703
rlabel metal2 1423 -1251 1423 -1251 0 net=9011
rlabel metal2 1591 -1251 1591 -1251 0 net=11221
rlabel metal2 1759 -1251 1759 -1251 0 net=10869
rlabel metal2 2004 -1251 2004 -1251 0 net=12223
rlabel metal2 2242 -1251 2242 -1251 0 net=13529
rlabel metal2 205 -1253 205 -1253 0 net=3031
rlabel metal2 562 -1253 562 -1253 0 net=4247
rlabel metal2 660 -1253 660 -1253 0 net=6933
rlabel metal2 1276 -1253 1276 -1253 0 net=7839
rlabel metal2 1447 -1253 1447 -1253 0 net=11860
rlabel metal2 2249 -1253 2249 -1253 0 net=13871
rlabel metal2 205 -1255 205 -1255 0 net=12418
rlabel metal2 282 -1257 282 -1257 0 net=1557
rlabel metal2 607 -1257 607 -1257 0 net=4976
rlabel metal2 863 -1257 863 -1257 0 net=12493
rlabel metal2 282 -1259 282 -1259 0 net=1517
rlabel metal2 541 -1259 541 -1259 0 net=5103
rlabel metal2 898 -1259 898 -1259 0 net=5473
rlabel metal2 985 -1259 985 -1259 0 net=9891
rlabel metal2 2004 -1259 2004 -1259 0 net=13013
rlabel metal2 93 -1261 93 -1261 0 net=5605
rlabel metal2 919 -1261 919 -1261 0 net=6689
rlabel metal2 1276 -1261 1276 -1261 0 net=7939
rlabel metal2 1367 -1261 1367 -1261 0 net=8513
rlabel metal2 1451 -1261 1451 -1261 0 net=7521
rlabel metal2 1703 -1261 1703 -1261 0 net=10677
rlabel metal2 1913 -1261 1913 -1261 0 net=11901
rlabel metal2 86 -1263 86 -1263 0 net=3937
rlabel metal2 110 -1263 110 -1263 0 net=9721
rlabel metal2 1752 -1263 1752 -1263 0 net=10823
rlabel metal2 2018 -1263 2018 -1263 0 net=12275
rlabel metal2 86 -1265 86 -1265 0 net=5811
rlabel metal2 632 -1265 632 -1265 0 net=4382
rlabel metal2 709 -1265 709 -1265 0 net=7255
rlabel metal2 954 -1265 954 -1265 0 net=896
rlabel metal2 1073 -1265 1073 -1265 0 net=5305
rlabel metal2 1325 -1265 1325 -1265 0 net=7497
rlabel metal2 1402 -1265 1402 -1265 0 net=8745
rlabel metal2 44 -1267 44 -1267 0 net=4085
rlabel metal2 723 -1267 723 -1267 0 net=11882
rlabel metal2 2032 -1267 2032 -1267 0 net=12389
rlabel metal2 44 -1269 44 -1269 0 net=4435
rlabel metal2 464 -1269 464 -1269 0 net=5793
rlabel metal2 1080 -1269 1080 -1269 0 net=6833
rlabel metal2 1402 -1269 1402 -1269 0 net=7875
rlabel metal2 1507 -1269 1507 -1269 0 net=9233
rlabel metal2 1766 -1269 1766 -1269 0 net=11497
rlabel metal2 2039 -1269 2039 -1269 0 net=12361
rlabel metal2 243 -1271 243 -1271 0 net=4037
rlabel metal2 541 -1271 541 -1271 0 net=3599
rlabel metal2 625 -1271 625 -1271 0 net=3505
rlabel metal2 639 -1271 639 -1271 0 net=13747
rlabel metal2 597 -1273 597 -1273 0 net=3745
rlabel metal2 989 -1273 989 -1273 0 net=6911
rlabel metal2 1143 -1273 1143 -1273 0 net=7083
rlabel metal2 1528 -1273 1528 -1273 0 net=9277
rlabel metal2 1626 -1273 1626 -1273 0 net=9947
rlabel metal2 1773 -1273 1773 -1273 0 net=10999
rlabel metal2 2046 -1273 2046 -1273 0 net=12519
rlabel metal2 142 -1275 142 -1275 0 net=11651
rlabel metal2 2053 -1275 2053 -1275 0 net=12285
rlabel metal2 142 -1277 142 -1277 0 net=2375
rlabel metal2 1136 -1277 1136 -1277 0 net=9331
rlabel metal2 1640 -1277 1640 -1277 0 net=10017
rlabel metal2 1780 -1277 1780 -1277 0 net=11071
rlabel metal2 2011 -1277 2011 -1277 0 net=12245
rlabel metal2 618 -1279 618 -1279 0 net=3395
rlabel metal2 1227 -1279 1227 -1279 0 net=7883
rlabel metal2 1535 -1279 1535 -1279 0 net=9409
rlabel metal2 1647 -1279 1647 -1279 0 net=10111
rlabel metal2 1780 -1279 1780 -1279 0 net=12145
rlabel metal2 625 -1281 625 -1281 0 net=4833
rlabel metal2 996 -1281 996 -1281 0 net=6495
rlabel metal2 1143 -1281 1143 -1281 0 net=6583
rlabel metal2 1171 -1281 1171 -1281 0 net=7089
rlabel metal2 1237 -1281 1237 -1281 0 net=9415
rlabel metal2 1661 -1281 1661 -1281 0 net=10457
rlabel metal2 1850 -1281 1850 -1281 0 net=11571
rlabel metal2 660 -1283 660 -1283 0 net=5421
rlabel metal2 996 -1283 996 -1283 0 net=10089
rlabel metal2 688 -1285 688 -1285 0 net=8144
rlabel metal2 999 -1285 999 -1285 0 net=6765
rlabel metal2 1311 -1285 1311 -1285 0 net=7425
rlabel metal2 1542 -1285 1542 -1285 0 net=9483
rlabel metal2 1717 -1285 1717 -1285 0 net=11469
rlabel metal2 688 -1287 688 -1287 0 net=3307
rlabel metal2 1052 -1287 1052 -1287 0 net=6663
rlabel metal2 1391 -1287 1391 -1287 0 net=1
rlabel metal2 1556 -1287 1556 -1287 0 net=9503
rlabel metal2 1787 -1287 1787 -1287 0 net=11129
rlabel metal2 765 -1289 765 -1289 0 net=7191
rlabel metal2 1430 -1289 1430 -1289 0 net=9713
rlabel metal2 1808 -1289 1808 -1289 0 net=11323
rlabel metal2 695 -1291 695 -1291 0 net=4265
rlabel metal2 1024 -1291 1024 -1291 0 net=6365
rlabel metal2 1150 -1291 1150 -1291 0 net=7379
rlabel metal2 1430 -1291 1430 -1291 0 net=11201
rlabel metal2 695 -1293 695 -1293 0 net=6069
rlabel metal2 1024 -1293 1024 -1293 0 net=5859
rlabel metal2 1108 -1293 1108 -1293 0 net=7000
rlabel metal2 1213 -1293 1213 -1293 0 net=9693
rlabel metal2 1836 -1293 1836 -1293 0 net=11517
rlabel metal2 51 -1295 51 -1295 0 net=6139
rlabel metal2 1108 -1295 1108 -1295 0 net=6299
rlabel metal2 1153 -1295 1153 -1295 0 net=10419
rlabel metal2 1850 -1295 1850 -1295 0 net=10463
rlabel metal2 51 -1297 51 -1297 0 net=8083
rlabel metal2 450 -1297 450 -1297 0 net=4159
rlabel metal2 1213 -1297 1213 -1297 0 net=13220
rlabel metal2 58 -1299 58 -1299 0 net=5277
rlabel metal2 450 -1299 450 -1299 0 net=3439
rlabel metal2 1017 -1299 1017 -1299 0 net=6177
rlabel metal2 1444 -1299 1444 -1299 0 net=8885
rlabel metal2 1556 -1299 1556 -1299 0 net=8937
rlabel metal2 352 -1301 352 -1301 0 net=4349
rlabel metal2 933 -1301 933 -1301 0 net=3919
rlabel metal2 1479 -1301 1479 -1301 0 net=9163
rlabel metal2 2025 -1301 2025 -1301 0 net=12353
rlabel metal2 352 -1303 352 -1303 0 net=2543
rlabel metal2 793 -1303 793 -1303 0 net=5335
rlabel metal2 1013 -1303 1013 -1303 0 net=11509
rlabel metal2 2081 -1303 2081 -1303 0 net=13635
rlabel metal2 394 -1305 394 -1305 0 net=2519
rlabel metal2 761 -1305 761 -1305 0 net=11741
rlabel metal2 212 -1307 212 -1307 0 net=4643
rlabel metal2 793 -1307 793 -1307 0 net=12140
rlabel metal2 212 -1309 212 -1309 0 net=2659
rlabel metal2 1395 -1309 1395 -1309 0 net=8587
rlabel metal2 1493 -1309 1493 -1309 0 net=8909
rlabel metal2 1577 -1309 1577 -1309 0 net=9669
rlabel metal2 1864 -1309 1864 -1309 0 net=11699
rlabel metal2 170 -1311 170 -1311 0 net=2451
rlabel metal2 1006 -1311 1006 -1311 0 net=10531
rlabel metal2 1871 -1311 1871 -1311 0 net=11963
rlabel metal2 107 -1313 107 -1313 0 net=9565
rlabel metal2 1346 -1313 1346 -1313 0 net=8635
rlabel metal2 1584 -1313 1584 -1313 0 net=9733
rlabel metal2 1878 -1313 1878 -1313 0 net=12041
rlabel metal2 170 -1315 170 -1315 0 net=5897
rlabel metal2 1395 -1315 1395 -1315 0 net=8973
rlabel metal2 1465 -1315 1465 -1315 0 net=10639
rlabel metal2 247 -1317 247 -1317 0 net=7591
rlabel metal2 1472 -1317 1472 -1317 0 net=8997
rlabel metal2 1675 -1317 1675 -1317 0 net=10301
rlabel metal2 716 -1319 716 -1319 0 net=3867
rlabel metal2 779 -1319 779 -1319 0 net=8515
rlabel metal2 1472 -1319 1472 -1319 0 net=7991
rlabel metal2 359 -1321 359 -1321 0 net=5831
rlabel metal2 1318 -1321 1318 -1321 0 net=8123
rlabel metal2 1486 -1321 1486 -1321 0 net=9185
rlabel metal2 1675 -1321 1675 -1321 0 net=13302
rlabel metal2 163 -1323 163 -1323 0 net=2323
rlabel metal2 1202 -1323 1202 -1323 0 net=7463
rlabel metal2 1374 -1323 1374 -1323 0 net=8609
rlabel metal2 1510 -1323 1510 -1323 0 net=12433
rlabel metal2 156 -1325 156 -1325 0 net=2043
rlabel metal2 177 -1325 177 -1325 0 net=3639
rlabel metal2 1682 -1325 1682 -1325 0 net=10559
rlabel metal2 156 -1327 156 -1327 0 net=6939
rlabel metal2 1682 -1327 1682 -1327 0 net=14493
rlabel metal2 177 -1329 177 -1329 0 net=3113
rlabel metal2 240 -1329 240 -1329 0 net=1847
rlabel metal2 1689 -1329 1689 -1329 0 net=11415
rlabel metal2 184 -1331 184 -1331 0 net=1623
rlabel metal2 296 -1331 296 -1331 0 net=3519
rlabel metal2 1101 -1331 1101 -1331 0 net=9641
rlabel metal2 1710 -1331 1710 -1331 0 net=10093
rlabel metal2 289 -1333 289 -1333 0 net=3023
rlabel metal2 1822 -1333 1822 -1333 0 net=11411
rlabel metal2 317 -1335 317 -1335 0 net=2821
rlabel metal2 828 -1335 828 -1335 0 net=10317
rlabel metal2 1899 -1335 1899 -1335 0 net=10717
rlabel metal2 317 -1337 317 -1337 0 net=3239
rlabel metal2 366 -1339 366 -1339 0 net=2859
rlabel metal2 345 -1341 345 -1341 0 net=2985
rlabel metal2 345 -1343 345 -1343 0 net=2931
rlabel metal2 338 -1345 338 -1345 0 net=2287
rlabel metal2 121 -1347 121 -1347 0 net=4593
rlabel metal2 2 -1358 2 -1358 0 net=744
rlabel metal2 880 -1358 880 -1358 0 net=6496
rlabel metal2 1150 -1358 1150 -1358 0 net=12656
rlabel metal2 2343 -1358 2343 -1358 0 net=12554
rlabel metal2 26 -1360 26 -1360 0 net=8998
rlabel metal2 1794 -1360 1794 -1360 0 net=10145
rlabel metal2 2263 -1360 2263 -1360 0 net=13293
rlabel metal2 37 -1362 37 -1362 0 net=4810
rlabel metal2 996 -1362 996 -1362 0 net=9714
rlabel metal2 1794 -1362 1794 -1362 0 net=10465
rlabel metal2 2361 -1362 2361 -1362 0 net=13873
rlabel metal2 40 -1364 40 -1364 0 net=9892
rlabel metal2 44 -1366 44 -1366 0 net=4436
rlabel metal2 208 -1366 208 -1366 0 net=3628
rlabel metal2 464 -1366 464 -1366 0 net=5794
rlabel metal2 943 -1366 943 -1366 0 net=9164
rlabel metal2 1983 -1366 1983 -1366 0 net=13307
rlabel metal2 44 -1368 44 -1368 0 net=5812
rlabel metal2 89 -1368 89 -1368 0 net=2638
rlabel metal2 989 -1368 989 -1368 0 net=6445
rlabel metal2 1129 -1368 1129 -1368 0 net=6179
rlabel metal2 1129 -1368 1129 -1368 0 net=6179
rlabel metal2 1136 -1368 1136 -1368 0 net=7697
rlabel metal2 1213 -1368 1213 -1368 0 net=8938
rlabel metal2 1577 -1368 1577 -1368 0 net=9927
rlabel metal2 1717 -1368 1717 -1368 0 net=10019
rlabel metal2 1850 -1368 1850 -1368 0 net=10825
rlabel metal2 1976 -1368 1976 -1368 0 net=11573
rlabel metal2 2368 -1368 2368 -1368 0 net=13971
rlabel metal2 54 -1370 54 -1370 0 net=1015
rlabel metal2 93 -1370 93 -1370 0 net=3938
rlabel metal2 163 -1370 163 -1370 0 net=2045
rlabel metal2 163 -1370 163 -1370 0 net=2045
rlabel metal2 170 -1370 170 -1370 0 net=5899
rlabel metal2 282 -1370 282 -1370 0 net=1519
rlabel metal2 282 -1370 282 -1370 0 net=1519
rlabel metal2 317 -1370 317 -1370 0 net=3241
rlabel metal2 499 -1370 499 -1370 0 net=3170
rlabel metal2 642 -1370 642 -1370 0 net=8557
rlabel metal2 996 -1370 996 -1370 0 net=8761
rlabel metal2 1507 -1370 1507 -1370 0 net=10113
rlabel metal2 1913 -1370 1913 -1370 0 net=11295
rlabel metal2 2431 -1370 2431 -1370 0 net=14223
rlabel metal2 58 -1372 58 -1372 0 net=5279
rlabel metal2 72 -1372 72 -1372 0 net=2774
rlabel metal2 831 -1372 831 -1372 0 net=6010
rlabel metal2 957 -1372 957 -1372 0 net=8514
rlabel metal2 1426 -1372 1426 -1372 0 net=10532
rlabel metal2 1962 -1372 1962 -1372 0 net=11519
rlabel metal2 58 -1374 58 -1374 0 net=5003
rlabel metal2 79 -1374 79 -1374 0 net=6941
rlabel metal2 170 -1374 170 -1374 0 net=2095
rlabel metal2 240 -1374 240 -1374 0 net=1848
rlabel metal2 646 -1374 646 -1374 0 net=6734
rlabel metal2 982 -1374 982 -1374 0 net=14487
rlabel metal2 82 -1376 82 -1376 0 net=9234
rlabel metal2 1766 -1376 1766 -1376 0 net=12009
rlabel metal2 93 -1378 93 -1378 0 net=3521
rlabel metal2 317 -1378 317 -1378 0 net=1733
rlabel metal2 891 -1378 891 -1378 0 net=9588
rlabel metal2 107 -1380 107 -1380 0 net=9566
rlabel metal2 646 -1380 646 -1380 0 net=3099
rlabel metal2 681 -1380 681 -1380 0 net=3712
rlabel metal2 1006 -1380 1006 -1380 0 net=539
rlabel metal2 1472 -1380 1472 -1380 0 net=7993
rlabel metal2 1773 -1380 1773 -1380 0 net=10319
rlabel metal2 1864 -1380 1864 -1380 0 net=10871
rlabel metal2 2109 -1380 2109 -1380 0 net=12277
rlabel metal2 2529 -1380 2529 -1380 0 net=14659
rlabel metal2 110 -1382 110 -1382 0 net=9694
rlabel metal2 1797 -1382 1797 -1382 0 net=1
rlabel metal2 2193 -1382 2193 -1382 0 net=12849
rlabel metal2 2340 -1382 2340 -1382 0 net=6345
rlabel metal2 117 -1384 117 -1384 0 net=1153
rlabel metal2 226 -1384 226 -1384 0 net=3640
rlabel metal2 1430 -1384 1430 -1384 0 net=10560
rlabel metal2 2200 -1384 2200 -1384 0 net=11583
rlabel metal2 121 -1386 121 -1386 0 net=6976
rlabel metal2 1251 -1386 1251 -1386 0 net=11412
rlabel metal2 107 -1388 107 -1388 0 net=2175
rlabel metal2 128 -1388 128 -1388 0 net=3479
rlabel metal2 681 -1388 681 -1388 0 net=3869
rlabel metal2 772 -1388 772 -1388 0 net=4502
rlabel metal2 796 -1388 796 -1388 0 net=4336
rlabel metal2 954 -1388 954 -1388 0 net=5475
rlabel metal2 982 -1388 982 -1388 0 net=5307
rlabel metal2 1087 -1388 1087 -1388 0 net=6549
rlabel metal2 1213 -1388 1213 -1388 0 net=7091
rlabel metal2 1234 -1388 1234 -1388 0 net=7411
rlabel metal2 1332 -1388 1332 -1388 0 net=8201
rlabel metal2 1472 -1388 1472 -1388 0 net=8611
rlabel metal2 1500 -1388 1500 -1388 0 net=12964
rlabel metal2 128 -1390 128 -1390 0 net=5499
rlabel metal2 1013 -1390 1013 -1390 0 net=9948
rlabel metal2 1787 -1390 1787 -1390 0 net=10421
rlabel metal2 1871 -1390 1871 -1390 0 net=11073
rlabel metal2 2200 -1390 2200 -1390 0 net=14371
rlabel metal2 226 -1392 226 -1392 0 net=3797
rlabel metal2 516 -1392 516 -1392 0 net=3672
rlabel metal2 723 -1392 723 -1392 0 net=5661
rlabel metal2 1104 -1392 1104 -1392 0 net=842
rlabel metal2 1759 -1392 1759 -1392 0 net=11779
rlabel metal2 1822 -1392 1822 -1392 0 net=10751
rlabel metal2 1934 -1392 1934 -1392 0 net=11417
rlabel metal2 2270 -1392 2270 -1392 0 net=13335
rlabel metal2 2508 -1392 2508 -1392 0 net=14537
rlabel metal2 229 -1394 229 -1394 0 net=11341
rlabel metal2 1997 -1394 1997 -1394 0 net=11701
rlabel metal2 2116 -1394 2116 -1394 0 net=14053
rlabel metal2 2522 -1394 2522 -1394 0 net=14615
rlabel metal2 240 -1396 240 -1396 0 net=5955
rlabel metal2 772 -1396 772 -1396 0 net=4769
rlabel metal2 880 -1396 880 -1396 0 net=7256
rlabel metal2 1038 -1396 1038 -1396 0 net=7084
rlabel metal2 1370 -1396 1370 -1396 0 net=14225
rlabel metal2 2543 -1396 2543 -1396 0 net=14767
rlabel metal2 254 -1398 254 -1398 0 net=3308
rlabel metal2 726 -1398 726 -1398 0 net=1347
rlabel metal2 891 -1398 891 -1398 0 net=5405
rlabel metal2 1031 -1398 1031 -1398 0 net=5985
rlabel metal2 1041 -1398 1041 -1398 0 net=8746
rlabel metal2 254 -1400 254 -1400 0 net=3397
rlabel metal2 688 -1400 688 -1400 0 net=5084
rlabel metal2 779 -1400 779 -1400 0 net=10640
rlabel metal2 2165 -1400 2165 -1400 0 net=12767
rlabel metal2 296 -1402 296 -1402 0 net=2003
rlabel metal2 898 -1402 898 -1402 0 net=5607
rlabel metal2 1066 -1402 1066 -1402 0 net=4160
rlabel metal2 1115 -1402 1115 -1402 0 net=7381
rlabel metal2 1304 -1402 1304 -1402 0 net=7523
rlabel metal2 1482 -1402 1482 -1402 0 net=11902
rlabel metal2 2256 -1402 2256 -1402 0 net=13247
rlabel metal2 16 -1404 16 -1404 0 net=5545
rlabel metal2 1510 -1404 1510 -1404 0 net=11130
rlabel metal2 16 -1406 16 -1406 0 net=12309
rlabel metal2 2123 -1406 2123 -1406 0 net=12287
rlabel metal2 2277 -1406 2277 -1406 0 net=13657
rlabel metal2 310 -1408 310 -1408 0 net=5825
rlabel metal2 618 -1408 618 -1408 0 net=1863
rlabel metal2 730 -1408 730 -1408 0 net=4368
rlabel metal2 758 -1408 758 -1408 0 net=4943
rlabel metal2 905 -1408 905 -1408 0 net=11929
rlabel metal2 2207 -1408 2207 -1408 0 net=14061
rlabel metal2 184 -1410 184 -1410 0 net=1625
rlabel metal2 387 -1410 387 -1410 0 net=2187
rlabel metal2 387 -1410 387 -1410 0 net=2187
rlabel metal2 408 -1410 408 -1410 0 net=2604
rlabel metal2 866 -1410 866 -1410 0 net=11964
rlabel metal2 2410 -1410 2410 -1410 0 net=14079
rlabel metal2 184 -1412 184 -1412 0 net=1509
rlabel metal2 366 -1412 366 -1412 0 net=2987
rlabel metal2 415 -1412 415 -1412 0 net=2452
rlabel metal2 642 -1412 642 -1412 0 net=13847
rlabel metal2 2445 -1412 2445 -1412 0 net=14281
rlabel metal2 257 -1414 257 -1414 0 net=4597
rlabel metal2 422 -1414 422 -1414 0 net=1988
rlabel metal2 702 -1414 702 -1414 0 net=6675
rlabel metal2 1227 -1414 1227 -1414 0 net=7193
rlabel metal2 1258 -1414 1258 -1414 0 net=10090
rlabel metal2 219 -1416 219 -1416 0 net=2357
rlabel metal2 429 -1416 429 -1416 0 net=3091
rlabel metal2 730 -1416 730 -1416 0 net=8727
rlabel metal2 1384 -1416 1384 -1416 0 net=9765
rlabel metal2 1682 -1416 1682 -1416 0 net=14495
rlabel metal2 19 -1418 19 -1418 0 net=7443
rlabel metal2 436 -1418 436 -1418 0 net=7427
rlabel metal2 1332 -1418 1332 -1418 0 net=7625
rlabel metal2 1556 -1418 1556 -1418 0 net=9187
rlabel metal2 1591 -1418 1591 -1418 0 net=11223
rlabel metal2 2172 -1418 2172 -1418 0 net=12495
rlabel metal2 149 -1420 149 -1420 0 net=6471
rlabel metal2 247 -1420 247 -1420 0 net=9817
rlabel metal2 1780 -1420 1780 -1420 0 net=12147
rlabel metal2 2242 -1420 2242 -1420 0 net=13165
rlabel metal2 149 -1422 149 -1422 0 net=4267
rlabel metal2 789 -1422 789 -1422 0 net=14427
rlabel metal2 247 -1424 247 -1424 0 net=2545
rlabel metal2 366 -1424 366 -1424 0 net=2289
rlabel metal2 506 -1424 506 -1424 0 net=4233
rlabel metal2 765 -1424 765 -1424 0 net=6665
rlabel metal2 1178 -1424 1178 -1424 0 net=7283
rlabel metal2 1297 -1424 1297 -1424 0 net=7499
rlabel metal2 1353 -1424 1353 -1424 0 net=8637
rlabel metal2 1584 -1424 1584 -1424 0 net=10679
rlabel metal2 142 -1426 142 -1426 0 net=2377
rlabel metal2 1311 -1426 1311 -1426 0 net=7575
rlabel metal2 1591 -1426 1591 -1426 0 net=9369
rlabel metal2 1780 -1426 1780 -1426 0 net=10355
rlabel metal2 1836 -1426 1836 -1426 0 net=10719
rlabel metal2 142 -1428 142 -1428 0 net=2113
rlabel metal2 1003 -1428 1003 -1428 0 net=7607
rlabel metal2 1605 -1428 1605 -1428 0 net=9417
rlabel metal2 1815 -1428 1815 -1428 0 net=10649
rlabel metal2 1878 -1428 1878 -1428 0 net=12673
rlabel metal2 275 -1430 275 -1430 0 net=2325
rlabel metal2 471 -1430 471 -1430 0 net=2861
rlabel metal2 541 -1430 541 -1430 0 net=3600
rlabel metal2 1024 -1430 1024 -1430 0 net=5861
rlabel metal2 1150 -1430 1150 -1430 0 net=6690
rlabel metal2 1241 -1430 1241 -1430 0 net=7635
rlabel metal2 1619 -1430 1619 -1430 0 net=9279
rlabel metal2 1857 -1430 1857 -1430 0 net=10907
rlabel metal2 1955 -1430 1955 -1430 0 net=11511
rlabel metal2 289 -1432 289 -1432 0 net=3025
rlabel metal2 541 -1432 541 -1432 0 net=2937
rlabel metal2 1489 -1432 1489 -1432 0 net=9489
rlabel metal2 1633 -1432 1633 -1432 0 net=9599
rlabel metal2 1885 -1432 1885 -1432 0 net=11169
rlabel metal2 2025 -1432 2025 -1432 0 net=11871
rlabel metal2 289 -1434 289 -1434 0 net=2243
rlabel metal2 555 -1434 555 -1434 0 net=4475
rlabel metal2 814 -1434 814 -1434 0 net=5104
rlabel metal2 1153 -1434 1153 -1434 0 net=13385
rlabel metal2 135 -1436 135 -1436 0 net=3073
rlabel metal2 716 -1436 716 -1436 0 net=5833
rlabel metal2 1010 -1436 1010 -1436 0 net=6367
rlabel metal2 1059 -1436 1059 -1436 0 net=6163
rlabel metal2 1185 -1436 1185 -1436 0 net=6835
rlabel metal2 1241 -1436 1241 -1436 0 net=7225
rlabel metal2 1283 -1436 1283 -1436 0 net=7267
rlabel metal2 1647 -1436 1647 -1436 0 net=9643
rlabel metal2 1899 -1436 1899 -1436 0 net=12197
rlabel metal2 135 -1438 135 -1438 0 net=7757
rlabel metal2 716 -1438 716 -1438 0 net=4013
rlabel metal2 835 -1438 835 -1438 0 net=6883
rlabel metal2 1206 -1438 1206 -1438 0 net=6935
rlabel metal2 1248 -1438 1248 -1438 0 net=13647
rlabel metal2 250 -1440 250 -1440 0 net=7107
rlabel metal2 1255 -1440 1255 -1440 0 net=8705
rlabel metal2 1668 -1440 1668 -1440 0 net=9735
rlabel metal2 1927 -1440 1927 -1440 0 net=13015
rlabel metal2 2067 -1440 2067 -1440 0 net=11687
rlabel metal2 261 -1442 261 -1442 0 net=1763
rlabel metal2 677 -1442 677 -1442 0 net=559
rlabel metal2 1262 -1442 1262 -1442 0 net=7248
rlabel metal2 1283 -1442 1283 -1442 0 net=11000
rlabel metal2 1948 -1442 1948 -1442 0 net=11499
rlabel metal2 261 -1444 261 -1444 0 net=3033
rlabel metal2 674 -1444 674 -1444 0 net=7387
rlabel metal2 1381 -1444 1381 -1444 0 net=9847
rlabel metal2 1941 -1444 1941 -1444 0 net=11471
rlabel metal2 2018 -1444 2018 -1444 0 net=11759
rlabel metal2 9 -1446 9 -1446 0 net=5275
rlabel metal2 674 -1446 674 -1446 0 net=3537
rlabel metal2 737 -1446 737 -1446 0 net=12325
rlabel metal2 9 -1448 9 -1448 0 net=4609
rlabel metal2 1381 -1448 1381 -1448 0 net=7841
rlabel metal2 1503 -1448 1503 -1448 0 net=10037
rlabel metal2 1969 -1448 1969 -1448 0 net=11203
rlabel metal2 303 -1450 303 -1450 0 net=2087
rlabel metal2 450 -1450 450 -1450 0 net=3441
rlabel metal2 744 -1450 744 -1450 0 net=6101
rlabel metal2 1388 -1450 1388 -1450 0 net=7877
rlabel metal2 1514 -1450 1514 -1450 0 net=12123
rlabel metal2 2088 -1450 2088 -1450 0 net=12225
rlabel metal2 177 -1452 177 -1452 0 net=3115
rlabel metal2 352 -1452 352 -1452 0 net=2427
rlabel metal2 450 -1452 450 -1452 0 net=3747
rlabel metal2 709 -1452 709 -1452 0 net=4087
rlabel metal2 786 -1452 786 -1452 0 net=10953
rlabel metal2 177 -1454 177 -1454 0 net=2645
rlabel metal2 271 -1454 271 -1454 0 net=3739
rlabel metal2 786 -1454 786 -1454 0 net=8163
rlabel metal2 1024 -1454 1024 -1454 0 net=6657
rlabel metal2 1276 -1454 1276 -1454 0 net=7941
rlabel metal2 1969 -1454 1969 -1454 0 net=11669
rlabel metal2 191 -1456 191 -1456 0 net=2933
rlabel metal2 373 -1456 373 -1456 0 net=2521
rlabel metal2 443 -1456 443 -1456 0 net=3135
rlabel metal2 660 -1456 660 -1456 0 net=5423
rlabel metal2 1031 -1456 1031 -1456 0 net=5957
rlabel metal2 1157 -1456 1157 -1456 0 net=6615
rlabel metal2 2004 -1456 2004 -1456 0 net=12521
rlabel metal2 331 -1458 331 -1458 0 net=1559
rlabel metal2 401 -1458 401 -1458 0 net=1715
rlabel metal2 2011 -1458 2011 -1458 0 net=11743
rlabel metal2 2249 -1458 2249 -1458 0 net=13183
rlabel metal2 331 -1460 331 -1460 0 net=3271
rlabel metal2 632 -1460 632 -1460 0 net=3507
rlabel metal2 814 -1460 814 -1460 0 net=5301
rlabel metal2 940 -1460 940 -1460 0 net=6141
rlabel metal2 1122 -1460 1122 -1460 0 net=6465
rlabel metal2 2060 -1460 2060 -1460 0 net=12091
rlabel metal2 2347 -1460 2347 -1460 0 net=13749
rlabel metal2 114 -1462 114 -1462 0 net=5173
rlabel metal2 828 -1462 828 -1462 0 net=9261
rlabel metal2 2081 -1462 2081 -1462 0 net=12171
rlabel metal2 2417 -1462 2417 -1462 0 net=14211
rlabel metal2 51 -1464 51 -1464 0 net=8084
rlabel metal2 443 -1464 443 -1464 0 net=2445
rlabel metal2 835 -1464 835 -1464 0 net=4791
rlabel metal2 856 -1464 856 -1464 0 net=4569
rlabel metal2 912 -1464 912 -1464 0 net=3973
rlabel metal2 1612 -1464 1612 -1464 0 net=9485
rlabel metal2 2151 -1464 2151 -1464 0 net=12391
rlabel metal2 2473 -1464 2473 -1464 0 net=14461
rlabel metal2 51 -1466 51 -1466 0 net=4811
rlabel metal2 870 -1466 870 -1466 0 net=5055
rlabel metal2 919 -1466 919 -1466 0 net=3921
rlabel metal2 1122 -1466 1122 -1466 0 net=6585
rlabel metal2 1157 -1466 1157 -1466 0 net=11888
rlabel metal2 2515 -1466 2515 -1466 0 net=14569
rlabel metal2 471 -1468 471 -1468 0 net=2783
rlabel metal2 884 -1468 884 -1468 0 net=7866
rlabel metal2 1654 -1468 1654 -1468 0 net=9671
rlabel metal2 2158 -1468 2158 -1468 0 net=12435
rlabel metal2 2452 -1468 2452 -1468 0 net=14317
rlabel metal2 2536 -1468 2536 -1468 0 net=14645
rlabel metal2 338 -1470 338 -1470 0 net=4595
rlabel metal2 926 -1470 926 -1470 0 net=5337
rlabel metal2 940 -1470 940 -1470 0 net=13799
rlabel metal2 2375 -1470 2375 -1470 0 net=13319
rlabel metal2 205 -1472 205 -1472 0 net=5381
rlabel metal2 1017 -1472 1017 -1472 0 net=12030
rlabel metal2 2228 -1472 2228 -1472 0 net=13091
rlabel metal2 338 -1474 338 -1474 0 net=1997
rlabel metal2 478 -1474 478 -1474 0 net=2823
rlabel metal2 562 -1474 562 -1474 0 net=4249
rlabel metal2 877 -1474 877 -1474 0 net=13979
rlabel metal2 23 -1476 23 -1476 0 net=4521
rlabel metal2 625 -1476 625 -1476 0 net=4835
rlabel metal2 1143 -1476 1143 -1476 0 net=8783
rlabel metal2 1563 -1476 1563 -1476 0 net=9243
rlabel metal2 1696 -1476 1696 -1476 0 net=9855
rlabel metal2 1990 -1476 1990 -1476 0 net=11325
rlabel metal2 2312 -1476 2312 -1476 0 net=13531
rlabel metal2 2 -1478 2 -1478 0 net=2337
rlabel metal2 793 -1478 793 -1478 0 net=10081
rlabel metal2 1990 -1478 1990 -1478 0 net=12899
rlabel metal2 2396 -1478 2396 -1478 0 net=14195
rlabel metal2 23 -1480 23 -1480 0 net=10222
rlabel metal2 2144 -1480 2144 -1480 0 net=12363
rlabel metal2 2284 -1480 2284 -1480 0 net=12801
rlabel metal2 156 -1482 156 -1482 0 net=3051
rlabel metal2 1160 -1482 1160 -1482 0 net=8399
rlabel metal2 1486 -1482 1486 -1482 0 net=14523
rlabel metal2 380 -1484 380 -1484 0 net=3831
rlabel metal2 485 -1484 485 -1484 0 net=2695
rlabel metal2 1164 -1484 1164 -1484 0 net=6767
rlabel metal2 1521 -1484 1521 -1484 0 net=8911
rlabel metal2 1598 -1484 1598 -1484 0 net=9411
rlabel metal2 2046 -1484 2046 -1484 0 net=11653
rlabel metal2 2284 -1484 2284 -1484 0 net=14737
rlabel metal2 47 -1486 47 -1486 0 net=1130
rlabel metal2 1080 -1486 1080 -1486 0 net=6913
rlabel metal2 1367 -1486 1367 -1486 0 net=9589
rlabel metal2 2046 -1486 2046 -1486 0 net=12043
rlabel metal2 2298 -1486 2298 -1486 0 net=13433
rlabel metal2 212 -1488 212 -1488 0 net=2661
rlabel metal2 394 -1488 394 -1488 0 net=4645
rlabel metal2 821 -1488 821 -1488 0 net=7813
rlabel metal2 1542 -1488 1542 -1488 0 net=8985
rlabel metal2 2053 -1488 2053 -1488 0 net=12247
rlabel metal2 2137 -1488 2137 -1488 0 net=12355
rlabel metal2 2389 -1488 2389 -1488 0 net=14047
rlabel metal2 212 -1490 212 -1490 0 net=5201
rlabel metal2 1080 -1490 1080 -1490 0 net=6217
rlabel metal2 1549 -1490 1549 -1490 0 net=9013
rlabel metal2 1801 -1490 1801 -1490 0 net=10165
rlabel metal2 2214 -1490 2214 -1490 0 net=12915
rlabel metal2 2438 -1490 2438 -1490 0 net=14241
rlabel metal2 37 -1492 37 -1492 0 net=14515
rlabel metal2 394 -1494 394 -1494 0 net=3373
rlabel metal2 807 -1494 807 -1494 0 net=7825
rlabel metal2 1535 -1494 1535 -1494 0 net=8887
rlabel metal2 324 -1496 324 -1496 0 net=4039
rlabel metal2 1094 -1496 1094 -1496 0 net=6301
rlabel metal2 1395 -1496 1395 -1496 0 net=8975
rlabel metal2 1570 -1496 1570 -1496 0 net=9333
rlabel metal2 1801 -1496 1801 -1496 0 net=10459
rlabel metal2 324 -1498 324 -1498 0 net=5325
rlabel metal2 1045 -1498 1045 -1498 0 net=5719
rlabel metal2 1395 -1498 1395 -1498 0 net=7885
rlabel metal2 1626 -1498 1626 -1498 0 net=9505
rlabel metal2 1843 -1498 1843 -1498 0 net=10765
rlabel metal2 583 -1500 583 -1500 0 net=3249
rlabel metal2 695 -1500 695 -1500 0 net=6071
rlabel metal2 1409 -1500 1409 -1500 0 net=8833
rlabel metal2 1661 -1500 1661 -1500 0 net=9723
rlabel metal2 1745 -1500 1745 -1500 0 net=11261
rlabel metal2 30 -1502 30 -1502 0 net=3105
rlabel metal2 639 -1502 639 -1502 0 net=13409
rlabel metal2 1703 -1502 1703 -1502 0 net=9961
rlabel metal2 1745 -1502 1745 -1502 0 net=10303
rlabel metal2 30 -1504 30 -1504 0 net=3327
rlabel metal2 1416 -1504 1416 -1504 0 net=10493
rlabel metal2 100 -1506 100 -1506 0 net=2963
rlabel metal2 1416 -1506 1416 -1506 0 net=8125
rlabel metal2 1710 -1506 1710 -1506 0 net=10095
rlabel metal2 100 -1508 100 -1508 0 net=8433
rlabel metal2 233 -1508 233 -1508 0 net=2497
rlabel metal2 1437 -1508 1437 -1508 0 net=8383
rlabel metal2 72 -1510 72 -1510 0 net=7719
rlabel metal2 576 -1510 576 -1510 0 net=4351
rlabel metal2 198 -1512 198 -1512 0 net=6807
rlabel metal2 1458 -1512 1458 -1512 0 net=8517
rlabel metal2 576 -1514 576 -1514 0 net=1547
rlabel metal2 1465 -1514 1465 -1514 0 net=8589
rlabel metal2 1318 -1516 1318 -1516 0 net=7464
rlabel metal2 1318 -1518 1318 -1518 0 net=7593
rlabel metal2 1346 -1520 1346 -1520 0 net=13114
rlabel metal2 2319 -1522 2319 -1522 0 net=13637
rlabel metal2 1678 -1524 1678 -1524 0 net=12829
rlabel metal2 16 -1535 16 -1535 0 net=10819
rlabel metal2 93 -1535 93 -1535 0 net=3522
rlabel metal2 229 -1535 229 -1535 0 net=4352
rlabel metal2 1836 -1535 1836 -1535 0 net=10721
rlabel metal2 1836 -1535 1836 -1535 0 net=10721
rlabel metal2 1885 -1535 1885 -1535 0 net=11171
rlabel metal2 1885 -1535 1885 -1535 0 net=11171
rlabel metal2 2389 -1535 2389 -1535 0 net=14048
rlabel metal2 2431 -1535 2431 -1535 0 net=14224
rlabel metal2 23 -1537 23 -1537 0 net=2824
rlabel metal2 583 -1537 583 -1537 0 net=3106
rlabel metal2 807 -1537 807 -1537 0 net=7626
rlabel metal2 1360 -1537 1360 -1537 0 net=7268
rlabel metal2 1479 -1537 1479 -1537 0 net=11574
rlabel metal2 2284 -1537 2284 -1537 0 net=14739
rlabel metal2 23 -1539 23 -1539 0 net=6421
rlabel metal2 642 -1539 642 -1539 0 net=3740
rlabel metal2 719 -1539 719 -1539 0 net=8888
rlabel metal2 40 -1541 40 -1541 0 net=9262
rlabel metal2 859 -1541 859 -1541 0 net=8706
rlabel metal2 1496 -1541 1496 -1541 0 net=14646
rlabel metal2 44 -1543 44 -1543 0 net=7997
rlabel metal2 58 -1543 58 -1543 0 net=5005
rlabel metal2 58 -1543 58 -1543 0 net=5005
rlabel metal2 72 -1543 72 -1543 0 net=7720
rlabel metal2 943 -1543 943 -1543 0 net=9590
rlabel metal2 1710 -1543 1710 -1543 0 net=10753
rlabel metal2 1976 -1543 1976 -1543 0 net=12227
rlabel metal2 2284 -1543 2284 -1543 0 net=14213
rlabel metal2 44 -1545 44 -1545 0 net=8435
rlabel metal2 107 -1545 107 -1545 0 net=4135
rlabel metal2 821 -1545 821 -1545 0 net=10146
rlabel metal2 2305 -1545 2305 -1545 0 net=14243
rlabel metal2 47 -1547 47 -1547 0 net=2358
rlabel metal2 481 -1547 481 -1547 0 net=2964
rlabel metal2 583 -1547 583 -1547 0 net=3509
rlabel metal2 691 -1547 691 -1547 0 net=5302
rlabel metal2 821 -1547 821 -1547 0 net=8785
rlabel metal2 1150 -1547 1150 -1547 0 net=10680
rlabel metal2 1822 -1547 1822 -1547 0 net=11263
rlabel metal2 1990 -1547 1990 -1547 0 net=12901
rlabel metal2 2340 -1547 2340 -1547 0 net=11584
rlabel metal2 30 -1549 30 -1549 0 net=3329
rlabel metal2 527 -1549 527 -1549 0 net=4477
rlabel metal2 793 -1549 793 -1549 0 net=6447
rlabel metal2 1076 -1549 1076 -1549 0 net=12830
rlabel metal2 30 -1551 30 -1551 0 net=1521
rlabel metal2 310 -1551 310 -1551 0 net=1627
rlabel metal2 310 -1551 310 -1551 0 net=1627
rlabel metal2 366 -1551 366 -1551 0 net=2291
rlabel metal2 590 -1551 590 -1551 0 net=5826
rlabel metal2 625 -1551 625 -1551 0 net=10166
rlabel metal2 2403 -1551 2403 -1551 0 net=14571
rlabel metal2 51 -1553 51 -1553 0 net=3116
rlabel metal2 366 -1553 366 -1553 0 net=2989
rlabel metal2 590 -1553 590 -1553 0 net=1865
rlabel metal2 625 -1553 625 -1553 0 net=4837
rlabel metal2 880 -1553 880 -1553 0 net=6616
rlabel metal2 1538 -1553 1538 -1553 0 net=12288
rlabel metal2 51 -1555 51 -1555 0 net=5281
rlabel metal2 72 -1555 72 -1555 0 net=3035
rlabel metal2 268 -1555 268 -1555 0 net=5900
rlabel metal2 814 -1555 814 -1555 0 net=5987
rlabel metal2 1090 -1555 1090 -1555 0 net=14080
rlabel metal2 2 -1557 2 -1557 0 net=2339
rlabel metal2 268 -1557 268 -1557 0 net=5663
rlabel metal2 730 -1557 730 -1557 0 net=8728
rlabel metal2 1038 -1557 1038 -1557 0 net=7109
rlabel metal2 1248 -1557 1248 -1557 0 net=13750
rlabel metal2 65 -1559 65 -1559 0 net=7445
rlabel metal2 597 -1559 597 -1559 0 net=3137
rlabel metal2 597 -1559 597 -1559 0 net=3137
rlabel metal2 604 -1559 604 -1559 0 net=6937
rlabel metal2 1220 -1559 1220 -1559 0 net=7577
rlabel metal2 1332 -1559 1332 -1559 0 net=9419
rlabel metal2 1878 -1559 1878 -1559 0 net=12675
rlabel metal2 2123 -1559 2123 -1559 0 net=13167
rlabel metal2 2347 -1559 2347 -1559 0 net=14463
rlabel metal2 79 -1561 79 -1561 0 net=6943
rlabel metal2 723 -1561 723 -1561 0 net=6165
rlabel metal2 1094 -1561 1094 -1561 0 net=6303
rlabel metal2 1094 -1561 1094 -1561 0 net=6303
rlabel metal2 1129 -1561 1129 -1561 0 net=6181
rlabel metal2 1248 -1561 1248 -1561 0 net=7887
rlabel metal2 1402 -1561 1402 -1561 0 net=7943
rlabel metal2 79 -1563 79 -1563 0 net=3799
rlabel metal2 233 -1563 233 -1563 0 net=5276
rlabel metal2 646 -1563 646 -1563 0 net=3101
rlabel metal2 698 -1563 698 -1563 0 net=14375
rlabel metal2 100 -1565 100 -1565 0 net=2785
rlabel metal2 520 -1565 520 -1565 0 net=3871
rlabel metal2 702 -1565 702 -1565 0 net=6677
rlabel metal2 887 -1565 887 -1565 0 net=6658
rlabel metal2 1066 -1565 1066 -1565 0 net=6809
rlabel metal2 1192 -1565 1192 -1565 0 net=6550
rlabel metal2 1255 -1565 1255 -1565 0 net=7501
rlabel metal2 1311 -1565 1311 -1565 0 net=8519
rlabel metal2 1479 -1565 1479 -1565 0 net=8913
rlabel metal2 1584 -1565 1584 -1565 0 net=9767
rlabel metal2 1878 -1565 1878 -1565 0 net=11671
rlabel metal2 1990 -1565 1990 -1565 0 net=12093
rlabel metal2 2095 -1565 2095 -1565 0 net=11205
rlabel metal2 37 -1567 37 -1567 0 net=7095
rlabel metal2 1111 -1567 1111 -1567 0 net=10407
rlabel metal2 1906 -1567 1906 -1567 0 net=11761
rlabel metal2 2032 -1567 2032 -1567 0 net=12365
rlabel metal2 37 -1569 37 -1569 0 net=9487
rlabel metal2 1955 -1569 1955 -1569 0 net=11513
rlabel metal2 2095 -1569 2095 -1569 0 net=12917
rlabel metal2 121 -1571 121 -1571 0 net=2176
rlabel metal2 471 -1571 471 -1571 0 net=2863
rlabel metal2 534 -1571 534 -1571 0 net=4041
rlabel metal2 702 -1571 702 -1571 0 net=4235
rlabel metal2 779 -1571 779 -1571 0 net=5057
rlabel metal2 898 -1571 898 -1571 0 net=4570
rlabel metal2 961 -1571 961 -1571 0 net=12496
rlabel metal2 2214 -1571 2214 -1571 0 net=13649
rlabel metal2 114 -1573 114 -1573 0 net=4723
rlabel metal2 824 -1573 824 -1573 0 net=6145
rlabel metal2 898 -1573 898 -1573 0 net=6369
rlabel metal2 1129 -1573 1129 -1573 0 net=7413
rlabel metal2 1283 -1573 1283 -1573 0 net=7525
rlabel metal2 1360 -1573 1360 -1573 0 net=10872
rlabel metal2 1955 -1573 1955 -1573 0 net=12125
rlabel metal2 2172 -1573 2172 -1573 0 net=13387
rlabel metal2 2326 -1573 2326 -1573 0 net=14283
rlabel metal2 114 -1575 114 -1575 0 net=2159
rlabel metal2 212 -1575 212 -1575 0 net=5203
rlabel metal2 737 -1575 737 -1575 0 net=7388
rlabel metal2 1297 -1575 1297 -1575 0 net=8639
rlabel metal2 1395 -1575 1395 -1575 0 net=9281
rlabel metal2 1864 -1575 1864 -1575 0 net=11473
rlabel metal2 1969 -1575 1969 -1575 0 net=12173
rlabel metal2 2291 -1575 2291 -1575 0 net=13875
rlabel metal2 2445 -1575 2445 -1575 0 net=14769
rlabel metal2 121 -1577 121 -1577 0 net=3975
rlabel metal2 964 -1577 964 -1577 0 net=8189
rlabel metal2 1423 -1577 1423 -1577 0 net=10460
rlabel metal2 1829 -1577 1829 -1577 0 net=11521
rlabel metal2 2067 -1577 2067 -1577 0 net=12437
rlabel metal2 2361 -1577 2361 -1577 0 net=14517
rlabel metal2 128 -1579 128 -1579 0 net=5501
rlabel metal2 163 -1579 163 -1579 0 net=2047
rlabel metal2 163 -1579 163 -1579 0 net=2047
rlabel metal2 198 -1579 198 -1579 0 net=14496
rlabel metal2 128 -1581 128 -1581 0 net=3539
rlabel metal2 849 -1581 849 -1581 0 net=3923
rlabel metal2 989 -1581 989 -1581 0 net=6587
rlabel metal2 1143 -1581 1143 -1581 0 net=7285
rlabel metal2 1192 -1581 1192 -1581 0 net=7609
rlabel metal2 1353 -1581 1353 -1581 0 net=9015
rlabel metal2 1605 -1581 1605 -1581 0 net=9601
rlabel metal2 1766 -1581 1766 -1581 0 net=12011
rlabel metal2 1962 -1581 1962 -1581 0 net=12149
rlabel metal2 2081 -1581 2081 -1581 0 net=12851
rlabel metal2 2494 -1581 2494 -1581 0 net=14617
rlabel metal2 184 -1583 184 -1583 0 net=1511
rlabel metal2 212 -1583 212 -1583 0 net=1548
rlabel metal2 593 -1583 593 -1583 0 net=13209
rlabel metal2 2193 -1583 2193 -1583 0 net=13435
rlabel metal2 177 -1585 177 -1585 0 net=2647
rlabel metal2 219 -1585 219 -1585 0 net=6473
rlabel metal2 1122 -1585 1122 -1585 0 net=6617
rlabel metal2 2074 -1585 2074 -1585 0 net=12769
rlabel metal2 2298 -1585 2298 -1585 0 net=14227
rlabel metal2 135 -1587 135 -1587 0 net=7759
rlabel metal2 226 -1587 226 -1587 0 net=7035
rlabel metal2 1153 -1587 1153 -1587 0 net=8679
rlabel metal2 1286 -1587 1286 -1587 0 net=12159
rlabel metal2 2165 -1587 2165 -1587 0 net=13337
rlabel metal2 135 -1589 135 -1589 0 net=6103
rlabel metal2 1157 -1589 1157 -1589 0 net=11654
rlabel metal2 2270 -1589 2270 -1589 0 net=13533
rlabel metal2 233 -1591 233 -1591 0 net=2498
rlabel metal2 800 -1591 800 -1591 0 net=4596
rlabel metal2 236 -1593 236 -1593 0 net=4646
rlabel metal2 506 -1593 506 -1593 0 net=2939
rlabel metal2 667 -1593 667 -1593 0 net=3443
rlabel metal2 870 -1593 870 -1593 0 net=6073
rlabel metal2 1157 -1593 1157 -1593 0 net=7827
rlabel metal2 1423 -1593 1423 -1593 0 net=9491
rlabel metal2 1633 -1593 1633 -1593 0 net=10097
rlabel metal2 1766 -1593 1766 -1593 0 net=11343
rlabel metal2 2221 -1593 2221 -1593 0 net=13659
rlabel metal2 2312 -1593 2312 -1593 0 net=14055
rlabel metal2 240 -1595 240 -1595 0 net=5956
rlabel metal2 1045 -1595 1045 -1595 0 net=5721
rlabel metal2 1160 -1595 1160 -1595 0 net=2378
rlabel metal2 1304 -1595 1304 -1595 0 net=8385
rlabel metal2 1458 -1595 1458 -1595 0 net=10321
rlabel metal2 2277 -1595 2277 -1595 0 net=14197
rlabel metal2 156 -1597 156 -1597 0 net=3053
rlabel metal2 247 -1597 247 -1597 0 net=2547
rlabel metal2 415 -1597 415 -1597 0 net=4599
rlabel metal2 828 -1597 828 -1597 0 net=2729
rlabel metal2 1171 -1597 1171 -1597 0 net=8127
rlabel metal2 1486 -1597 1486 -1597 0 net=9245
rlabel metal2 1612 -1597 1612 -1597 0 net=10467
rlabel metal2 2382 -1597 2382 -1597 0 net=14539
rlabel metal2 156 -1599 156 -1599 0 net=2097
rlabel metal2 275 -1599 275 -1599 0 net=2326
rlabel metal2 464 -1599 464 -1599 0 net=3243
rlabel metal2 667 -1599 667 -1599 0 net=5383
rlabel metal2 954 -1599 954 -1599 0 net=5476
rlabel metal2 1325 -1599 1325 -1599 0 net=8401
rlabel metal2 1489 -1599 1489 -1599 0 net=11326
rlabel metal2 2396 -1599 2396 -1599 0 net=14489
rlabel metal2 117 -1601 117 -1601 0 net=4303
rlabel metal2 478 -1601 478 -1601 0 net=3026
rlabel metal2 516 -1601 516 -1601 0 net=7179
rlabel metal2 1178 -1601 1178 -1601 0 net=7093
rlabel metal2 1265 -1601 1265 -1601 0 net=11113
rlabel metal2 1794 -1601 1794 -1601 0 net=11225
rlabel metal2 2235 -1601 2235 -1601 0 net=13849
rlabel metal2 149 -1603 149 -1603 0 net=4269
rlabel metal2 674 -1603 674 -1603 0 net=5407
rlabel metal2 905 -1603 905 -1603 0 net=5546
rlabel metal2 1493 -1603 1493 -1603 0 net=11039
rlabel metal2 1738 -1603 1738 -1603 0 net=10423
rlabel metal2 1892 -1603 1892 -1603 0 net=11703
rlabel metal2 2207 -1603 2207 -1603 0 net=14063
rlabel metal2 86 -1605 86 -1605 0 net=2825
rlabel metal2 170 -1605 170 -1605 0 net=3399
rlabel metal2 275 -1605 275 -1605 0 net=2005
rlabel metal2 303 -1605 303 -1605 0 net=1717
rlabel metal2 429 -1605 429 -1605 0 net=2447
rlabel metal2 695 -1605 695 -1605 0 net=4770
rlabel metal2 891 -1605 891 -1605 0 net=5609
rlabel metal2 982 -1605 982 -1605 0 net=5308
rlabel metal2 1213 -1605 1213 -1605 0 net=7995
rlabel metal2 1759 -1605 1759 -1605 0 net=11781
rlabel metal2 1983 -1605 1983 -1605 0 net=13309
rlabel metal2 86 -1607 86 -1607 0 net=2115
rlabel metal2 250 -1607 250 -1607 0 net=9807
rlabel metal2 1503 -1607 1503 -1607 0 net=12802
rlabel metal2 142 -1609 142 -1609 0 net=3713
rlabel metal2 772 -1609 772 -1609 0 net=4813
rlabel metal2 905 -1609 905 -1609 0 net=7843
rlabel metal2 1416 -1609 1416 -1609 0 net=8591
rlabel metal2 1507 -1609 1507 -1609 0 net=10115
rlabel metal2 1752 -1609 1752 -1609 0 net=11075
rlabel metal2 1997 -1609 1997 -1609 0 net=12249
rlabel metal2 110 -1611 110 -1611 0 net=190
rlabel metal2 1514 -1611 1514 -1611 0 net=9819
rlabel metal2 1759 -1611 1759 -1611 0 net=12199
rlabel metal2 2102 -1611 2102 -1611 0 net=13639
rlabel metal2 205 -1613 205 -1613 0 net=9309
rlabel metal2 1444 -1613 1444 -1613 0 net=9413
rlabel metal2 1787 -1613 1787 -1613 0 net=12279
rlabel metal2 2319 -1613 2319 -1613 0 net=14661
rlabel metal2 205 -1615 205 -1615 0 net=3481
rlabel metal2 842 -1615 842 -1615 0 net=5339
rlabel metal2 933 -1615 933 -1615 0 net=7382
rlabel metal2 1234 -1615 1234 -1615 0 net=7967
rlabel metal2 1531 -1615 1531 -1615 0 net=13321
rlabel metal2 254 -1617 254 -1617 0 net=7055
rlabel metal2 1276 -1617 1276 -1617 0 net=6466
rlabel metal2 1549 -1617 1549 -1617 0 net=9737
rlabel metal2 1815 -1617 1815 -1617 0 net=10651
rlabel metal2 282 -1619 282 -1619 0 net=2523
rlabel metal2 380 -1619 380 -1619 0 net=2663
rlabel metal2 380 -1619 380 -1619 0 net=2663
rlabel metal2 387 -1619 387 -1619 0 net=2189
rlabel metal2 912 -1619 912 -1619 0 net=9335
rlabel metal2 1668 -1619 1668 -1619 0 net=10357
rlabel metal2 1871 -1619 1871 -1619 0 net=11501
rlabel metal2 96 -1621 96 -1621 0 net=9869
rlabel metal2 1899 -1621 1899 -1621 0 net=11745
rlabel metal2 296 -1623 296 -1623 0 net=3251
rlabel metal2 919 -1623 919 -1623 0 net=5959
rlabel metal2 1034 -1623 1034 -1623 0 net=10075
rlabel metal2 1927 -1623 1927 -1623 0 net=13017
rlabel metal2 338 -1625 338 -1625 0 net=1999
rlabel metal2 436 -1625 436 -1625 0 net=7429
rlabel metal2 954 -1625 954 -1625 0 net=6143
rlabel metal2 1115 -1625 1115 -1625 0 net=7699
rlabel metal2 1258 -1625 1258 -1625 0 net=11235
rlabel metal2 1927 -1625 1927 -1625 0 net=11873
rlabel metal2 338 -1627 338 -1627 0 net=1561
rlabel metal2 352 -1627 352 -1627 0 net=2429
rlabel metal2 436 -1627 436 -1627 0 net=6735
rlabel metal2 1563 -1627 1563 -1627 0 net=9857
rlabel metal2 1948 -1627 1948 -1627 0 net=12045
rlabel metal2 289 -1629 289 -1629 0 net=2245
rlabel metal2 373 -1629 373 -1629 0 net=3833
rlabel metal2 562 -1629 562 -1629 0 net=4523
rlabel metal2 926 -1629 926 -1629 0 net=6885
rlabel metal2 1136 -1629 1136 -1629 0 net=7595
rlabel metal2 1349 -1629 1349 -1629 0 net=10403
rlabel metal2 1689 -1629 1689 -1629 0 net=9849
rlabel metal2 2004 -1629 2004 -1629 0 net=12523
rlabel metal2 2025 -1629 2025 -1629 0 net=12327
rlabel metal2 191 -1631 191 -1631 0 net=2935
rlabel metal2 317 -1631 317 -1631 0 net=1735
rlabel metal2 387 -1631 387 -1631 0 net=5835
rlabel metal2 1059 -1631 1059 -1631 0 net=5863
rlabel metal2 1262 -1631 1262 -1631 0 net=11173
rlabel metal2 2004 -1631 2004 -1631 0 net=12311
rlabel metal2 2130 -1631 2130 -1631 0 net=13185
rlabel metal2 191 -1633 191 -1633 0 net=6815
rlabel metal2 975 -1633 975 -1633 0 net=6219
rlabel metal2 1101 -1633 1101 -1633 0 net=7195
rlabel metal2 1276 -1633 1276 -1633 0 net=7911
rlabel metal2 1689 -1633 1689 -1633 0 net=10495
rlabel metal2 2046 -1633 2046 -1633 0 net=12357
rlabel metal2 2249 -1633 2249 -1633 0 net=14429
rlabel metal2 194 -1635 194 -1635 0 net=605
rlabel metal2 1318 -1635 1318 -1635 0 net=9673
rlabel metal2 1808 -1635 1808 -1635 0 net=11688
rlabel metal2 317 -1637 317 -1637 0 net=2089
rlabel metal2 394 -1637 394 -1637 0 net=3374
rlabel metal2 968 -1637 968 -1637 0 net=8559
rlabel metal2 1293 -1637 1293 -1637 0 net=10167
rlabel metal2 2116 -1637 2116 -1637 0 net=13093
rlabel metal2 324 -1639 324 -1639 0 net=5326
rlabel metal2 548 -1639 548 -1639 0 net=3075
rlabel metal2 639 -1639 639 -1639 0 net=13320
rlabel metal2 324 -1641 324 -1641 0 net=1765
rlabel metal2 856 -1641 856 -1641 0 net=4250
rlabel metal2 982 -1641 982 -1641 0 net=6769
rlabel metal2 1374 -1641 1374 -1641 0 net=8977
rlabel metal2 2137 -1641 2137 -1641 0 net=13981
rlabel metal2 331 -1643 331 -1643 0 net=3273
rlabel metal2 394 -1643 394 -1643 0 net=5175
rlabel metal2 653 -1643 653 -1643 0 net=6051
rlabel metal2 1003 -1643 1003 -1643 0 net=6837
rlabel metal2 1500 -1643 1500 -1643 0 net=9507
rlabel metal2 2200 -1643 2200 -1643 0 net=14373
rlabel metal2 331 -1645 331 -1645 0 net=2697
rlabel metal2 548 -1645 548 -1645 0 net=4945
rlabel metal2 1073 -1645 1073 -1645 0 net=10954
rlabel metal2 2200 -1645 2200 -1645 0 net=13295
rlabel metal2 180 -1647 180 -1647 0 net=13235
rlabel metal2 2228 -1647 2228 -1647 0 net=13801
rlabel metal2 443 -1649 443 -1649 0 net=5841
rlabel metal2 1468 -1649 1468 -1649 0 net=14143
rlabel metal2 2333 -1649 2333 -1649 0 net=14319
rlabel metal2 450 -1651 450 -1651 0 net=3749
rlabel metal2 758 -1651 758 -1651 0 net=4793
rlabel metal2 996 -1651 996 -1651 0 net=8763
rlabel metal2 1430 -1651 1430 -1651 0 net=8203
rlabel metal2 450 -1653 450 -1653 0 net=4571
rlabel metal2 765 -1653 765 -1653 0 net=6667
rlabel metal2 1080 -1653 1080 -1653 0 net=6915
rlabel metal2 1430 -1653 1430 -1653 0 net=9189
rlabel metal2 1626 -1653 1626 -1653 0 net=10083
rlabel metal2 485 -1655 485 -1655 0 net=4015
rlabel metal2 765 -1655 765 -1655 0 net=4669
rlabel metal2 1164 -1655 1164 -1655 0 net=7815
rlabel metal2 1528 -1655 1528 -1655 0 net=13411
rlabel metal2 513 -1657 513 -1657 0 net=6963
rlabel metal2 1087 -1657 1087 -1657 0 net=7169
rlabel metal2 1367 -1657 1367 -1657 0 net=8613
rlabel metal2 1535 -1657 1535 -1657 0 net=12729
rlabel metal2 513 -1659 513 -1659 0 net=2379
rlabel metal2 786 -1659 786 -1659 0 net=8165
rlabel metal2 1388 -1659 1388 -1659 0 net=7878
rlabel metal2 1556 -1659 1556 -1659 0 net=10039
rlabel metal2 866 -1661 866 -1661 0 net=10417
rlabel metal2 555 -1663 555 -1663 0 net=3205
rlabel metal2 569 -1665 569 -1665 0 net=3092
rlabel metal2 1185 -1665 1185 -1665 0 net=7227
rlabel metal2 1388 -1665 1388 -1665 0 net=8987
rlabel metal2 1724 -1665 1724 -1665 0 net=10827
rlabel metal2 569 -1667 569 -1667 0 net=1573
rlabel metal2 1241 -1667 1241 -1667 0 net=7637
rlabel metal2 1472 -1667 1472 -1667 0 net=9725
rlabel metal2 1850 -1667 1850 -1667 0 net=11419
rlabel metal2 688 -1669 688 -1669 0 net=4089
rlabel metal2 863 -1669 863 -1669 0 net=5425
rlabel metal2 1339 -1669 1339 -1669 0 net=8835
rlabel metal2 1542 -1669 1542 -1669 0 net=9645
rlabel metal2 1661 -1669 1661 -1669 0 net=10305
rlabel metal2 1934 -1669 1934 -1669 0 net=11931
rlabel metal2 9 -1671 9 -1671 0 net=4611
rlabel metal2 947 -1671 947 -1671 0 net=6347
rlabel metal2 93 -1673 93 -1673 0 net=12477
rlabel metal2 1409 -1675 1409 -1675 0 net=9371
rlabel metal2 1745 -1675 1745 -1675 0 net=10909
rlabel metal2 1510 -1677 1510 -1677 0 net=11453
rlabel metal2 1577 -1679 1577 -1679 0 net=9929
rlabel metal2 1577 -1681 1577 -1681 0 net=9963
rlabel metal2 1591 -1683 1591 -1683 0 net=10021
rlabel metal2 1703 -1685 1703 -1685 0 net=4383
rlabel metal2 1717 -1687 1717 -1687 0 net=10767
rlabel metal2 1843 -1689 1843 -1689 0 net=11297
rlabel metal2 1913 -1691 1913 -1691 0 net=12393
rlabel metal2 2151 -1693 2151 -1693 0 net=13249
rlabel metal2 2256 -1695 2256 -1695 0 net=13973
rlabel metal2 2368 -1697 2368 -1697 0 net=14525
rlabel metal2 2 -1708 2 -1708 0 net=5837
rlabel metal2 422 -1708 422 -1708 0 net=3331
rlabel metal2 422 -1708 422 -1708 0 net=3331
rlabel metal2 429 -1708 429 -1708 0 net=2448
rlabel metal2 1549 -1708 1549 -1708 0 net=9739
rlabel metal2 1549 -1708 1549 -1708 0 net=9739
rlabel metal2 1629 -1708 1629 -1708 0 net=12358
rlabel metal2 2389 -1708 2389 -1708 0 net=14741
rlabel metal2 2445 -1708 2445 -1708 0 net=14771
rlabel metal2 2469 -1708 2469 -1708 0 net=14618
rlabel metal2 9 -1710 9 -1710 0 net=4137
rlabel metal2 142 -1710 142 -1710 0 net=3715
rlabel metal2 163 -1710 163 -1710 0 net=2049
rlabel metal2 163 -1710 163 -1710 0 net=2049
rlabel metal2 187 -1710 187 -1710 0 net=147
rlabel metal2 1276 -1710 1276 -1710 0 net=4384
rlabel metal2 16 -1712 16 -1712 0 net=10820
rlabel metal2 649 -1712 649 -1712 0 net=716
rlabel metal2 1017 -1712 1017 -1712 0 net=9602
rlabel metal2 1640 -1712 1640 -1712 0 net=10117
rlabel metal2 1640 -1712 1640 -1712 0 net=10117
rlabel metal2 1664 -1712 1664 -1712 0 net=14056
rlabel metal2 2347 -1712 2347 -1712 0 net=14465
rlabel metal2 16 -1714 16 -1714 0 net=6839
rlabel metal2 1020 -1714 1020 -1714 0 net=7610
rlabel metal2 1206 -1714 1206 -1714 0 net=6182
rlabel metal2 1293 -1714 1293 -1714 0 net=13534
rlabel metal2 2389 -1714 2389 -1714 0 net=13035
rlabel metal2 23 -1716 23 -1716 0 net=6423
rlabel metal2 23 -1716 23 -1716 0 net=6423
rlabel metal2 30 -1716 30 -1716 0 net=1522
rlabel metal2 919 -1716 919 -1716 0 net=5961
rlabel metal2 919 -1716 919 -1716 0 net=5961
rlabel metal2 989 -1716 989 -1716 0 net=6589
rlabel metal2 1031 -1716 1031 -1716 0 net=8190
rlabel metal2 1437 -1716 1437 -1716 0 net=10424
rlabel metal2 1801 -1716 1801 -1716 0 net=12160
rlabel metal2 30 -1718 30 -1718 0 net=2699
rlabel metal2 446 -1718 446 -1718 0 net=2190
rlabel metal2 821 -1718 821 -1718 0 net=8786
rlabel metal2 1108 -1718 1108 -1718 0 net=7944
rlabel metal2 37 -1720 37 -1720 0 net=9488
rlabel metal2 107 -1720 107 -1720 0 net=3835
rlabel metal2 394 -1720 394 -1720 0 net=5177
rlabel metal2 821 -1720 821 -1720 0 net=2909
rlabel metal2 1367 -1720 1367 -1720 0 net=8615
rlabel metal2 1440 -1720 1440 -1720 0 net=13876
rlabel metal2 2361 -1720 2361 -1720 0 net=14519
rlabel metal2 37 -1722 37 -1722 0 net=5843
rlabel metal2 457 -1722 457 -1722 0 net=2731
rlabel metal2 835 -1722 835 -1722 0 net=6668
rlabel metal2 961 -1722 961 -1722 0 net=6475
rlabel metal2 1059 -1722 1059 -1722 0 net=5865
rlabel metal2 1111 -1722 1111 -1722 0 net=11172
rlabel metal2 1997 -1722 1997 -1722 0 net=12251
rlabel metal2 2228 -1722 2228 -1722 0 net=13803
rlabel metal2 2305 -1722 2305 -1722 0 net=14245
rlabel metal2 47 -1724 47 -1724 0 net=5282
rlabel metal2 65 -1724 65 -1724 0 net=7446
rlabel metal2 194 -1724 194 -1724 0 net=7196
rlabel metal2 1129 -1724 1129 -1724 0 net=7415
rlabel metal2 1129 -1724 1129 -1724 0 net=7415
rlabel metal2 1153 -1724 1153 -1724 0 net=9850
rlabel metal2 1706 -1724 1706 -1724 0 net=14374
rlabel metal2 51 -1726 51 -1726 0 net=3055
rlabel metal2 247 -1726 247 -1726 0 net=3244
rlabel metal2 548 -1726 548 -1726 0 net=4946
rlabel metal2 870 -1726 870 -1726 0 net=6075
rlabel metal2 989 -1726 989 -1726 0 net=7037
rlabel metal2 1059 -1726 1059 -1726 0 net=9373
rlabel metal2 1440 -1726 1440 -1726 0 net=10427
rlabel metal2 1836 -1726 1836 -1726 0 net=10722
rlabel metal2 58 -1728 58 -1728 0 net=5007
rlabel metal2 86 -1728 86 -1728 0 net=2116
rlabel metal2 198 -1728 198 -1728 0 net=1512
rlabel metal2 1192 -1728 1192 -1728 0 net=7527
rlabel metal2 1293 -1728 1293 -1728 0 net=9414
rlabel metal2 1458 -1728 1458 -1728 0 net=10323
rlabel metal2 2039 -1728 2039 -1728 0 net=12479
rlabel metal2 2228 -1728 2228 -1728 0 net=14663
rlabel metal2 58 -1730 58 -1730 0 net=6371
rlabel metal2 957 -1730 957 -1730 0 net=10783
rlabel metal2 1468 -1730 1468 -1730 0 net=14490
rlabel metal2 86 -1732 86 -1732 0 net=6105
rlabel metal2 142 -1732 142 -1732 0 net=1947
rlabel metal2 460 -1732 460 -1732 0 net=3750
rlabel metal2 653 -1732 653 -1732 0 net=6053
rlabel metal2 870 -1732 870 -1732 0 net=5611
rlabel metal2 1003 -1732 1003 -1732 0 net=6305
rlabel metal2 1143 -1732 1143 -1732 0 net=7287
rlabel metal2 1209 -1732 1209 -1732 0 net=8978
rlabel metal2 1388 -1732 1388 -1732 0 net=8989
rlabel metal2 1468 -1732 1468 -1732 0 net=13813
rlabel metal2 44 -1734 44 -1734 0 net=8437
rlabel metal2 1493 -1734 1493 -1734 0 net=9930
rlabel metal2 1696 -1734 1696 -1734 0 net=12013
rlabel metal2 2039 -1734 2039 -1734 0 net=13983
rlabel metal2 2235 -1734 2235 -1734 0 net=13851
rlabel metal2 93 -1736 93 -1736 0 net=6886
rlabel metal2 1143 -1736 1143 -1736 0 net=7047
rlabel metal2 1213 -1736 1213 -1736 0 net=7996
rlabel metal2 1325 -1736 1325 -1736 0 net=8403
rlabel metal2 1493 -1736 1493 -1736 0 net=10023
rlabel metal2 1647 -1736 1647 -1736 0 net=10061
rlabel metal2 1815 -1736 1815 -1736 0 net=11237
rlabel metal2 1850 -1736 1850 -1736 0 net=11421
rlabel metal2 1941 -1736 1941 -1736 0 net=13323
rlabel metal2 2179 -1736 2179 -1736 0 net=13413
rlabel metal2 2242 -1736 2242 -1736 0 net=11207
rlabel metal2 2284 -1736 2284 -1736 0 net=14215
rlabel metal2 93 -1738 93 -1738 0 net=2665
rlabel metal2 429 -1738 429 -1738 0 net=7957
rlabel metal2 1171 -1738 1171 -1738 0 net=8129
rlabel metal2 1360 -1738 1360 -1738 0 net=13310
rlabel metal2 2221 -1738 2221 -1738 0 net=13661
rlabel metal2 135 -1740 135 -1740 0 net=3483
rlabel metal2 212 -1740 212 -1740 0 net=5426
rlabel metal2 884 -1740 884 -1740 0 net=6679
rlabel metal2 1164 -1740 1164 -1740 0 net=7817
rlabel metal2 1213 -1740 1213 -1740 0 net=7639
rlabel metal2 1255 -1740 1255 -1740 0 net=7503
rlabel metal2 1255 -1740 1255 -1740 0 net=7503
rlabel metal2 1262 -1740 1262 -1740 0 net=11514
rlabel metal2 2081 -1740 2081 -1740 0 net=12853
rlabel metal2 2151 -1740 2151 -1740 0 net=13251
rlabel metal2 2263 -1740 2263 -1740 0 net=14145
rlabel metal2 100 -1742 100 -1742 0 net=2787
rlabel metal2 212 -1742 212 -1742 0 net=4795
rlabel metal2 765 -1742 765 -1742 0 net=4671
rlabel metal2 765 -1742 765 -1742 0 net=4671
rlabel metal2 793 -1742 793 -1742 0 net=6449
rlabel metal2 1220 -1742 1220 -1742 0 net=7579
rlabel metal2 1220 -1742 1220 -1742 0 net=7579
rlabel metal2 1227 -1742 1227 -1742 0 net=8561
rlabel metal2 1500 -1742 1500 -1742 0 net=9509
rlabel metal2 1500 -1742 1500 -1742 0 net=9509
rlabel metal2 1510 -1742 1510 -1742 0 net=13296
rlabel metal2 198 -1744 198 -1744 0 net=2990
rlabel metal2 373 -1744 373 -1744 0 net=8315
rlabel metal2 579 -1744 579 -1744 0 net=10707
rlabel metal2 1745 -1744 1745 -1744 0 net=10911
rlabel metal2 226 -1746 226 -1746 0 net=9336
rlabel metal2 940 -1746 940 -1746 0 net=7431
rlabel metal2 1185 -1746 1185 -1746 0 net=7229
rlabel metal2 1241 -1746 1241 -1746 0 net=8521
rlabel metal2 1353 -1746 1353 -1746 0 net=9017
rlabel metal2 1528 -1746 1528 -1746 0 net=14572
rlabel metal2 229 -1748 229 -1748 0 net=3581
rlabel metal2 1248 -1748 1248 -1748 0 net=7889
rlabel metal2 1283 -1748 1283 -1748 0 net=7913
rlabel metal2 1528 -1748 1528 -1748 0 net=9647
rlabel metal2 1556 -1748 1556 -1748 0 net=10041
rlabel metal2 1724 -1748 1724 -1748 0 net=10829
rlabel metal2 1759 -1748 1759 -1748 0 net=12201
rlabel metal2 2102 -1748 2102 -1748 0 net=13641
rlabel metal2 2333 -1748 2333 -1748 0 net=14321
rlabel metal2 124 -1750 124 -1750 0 net=9619
rlabel metal2 1531 -1750 1531 -1750 0 net=14081
rlabel metal2 236 -1752 236 -1752 0 net=6144
rlabel metal2 1052 -1752 1052 -1752 0 net=7181
rlabel metal2 1297 -1752 1297 -1752 0 net=8641
rlabel metal2 1535 -1752 1535 -1752 0 net=12902
rlabel metal2 2130 -1752 2130 -1752 0 net=13187
rlabel metal2 240 -1754 240 -1754 0 net=2611
rlabel metal2 1234 -1754 1234 -1754 0 net=7969
rlabel metal2 1304 -1754 1304 -1754 0 net=8387
rlabel metal2 1535 -1754 1535 -1754 0 net=10469
rlabel metal2 1619 -1754 1619 -1754 0 net=11041
rlabel metal2 1773 -1754 1773 -1754 0 net=11115
rlabel metal2 1850 -1754 1850 -1754 0 net=14064
rlabel metal2 254 -1756 254 -1756 0 net=7057
rlabel metal2 254 -1756 254 -1756 0 net=7057
rlabel metal2 289 -1756 289 -1756 0 net=2936
rlabel metal2 702 -1756 702 -1756 0 net=4237
rlabel metal2 702 -1756 702 -1756 0 net=4237
rlabel metal2 716 -1756 716 -1756 0 net=11507
rlabel metal2 2165 -1756 2165 -1756 0 net=13339
rlabel metal2 2298 -1756 2298 -1756 0 net=14229
rlabel metal2 289 -1758 289 -1758 0 net=1767
rlabel metal2 331 -1758 331 -1758 0 net=2381
rlabel metal2 520 -1758 520 -1758 0 net=3873
rlabel metal2 653 -1758 653 -1758 0 net=4601
rlabel metal2 744 -1758 744 -1758 0 net=4613
rlabel metal2 1157 -1758 1157 -1758 0 net=7829
rlabel metal2 1290 -1758 1290 -1758 0 net=13115
rlabel metal2 2179 -1758 2179 -1758 0 net=14541
rlabel metal2 303 -1760 303 -1760 0 net=1719
rlabel metal2 303 -1760 303 -1760 0 net=1719
rlabel metal2 324 -1760 324 -1760 0 net=1867
rlabel metal2 618 -1760 618 -1760 0 net=6817
rlabel metal2 1115 -1760 1115 -1760 0 net=7701
rlabel metal2 1304 -1760 1304 -1760 0 net=13379
rlabel metal2 1808 -1760 1808 -1760 0 net=12395
rlabel metal2 2053 -1760 2053 -1760 0 net=12677
rlabel metal2 2151 -1760 2151 -1760 0 net=13023
rlabel metal2 121 -1762 121 -1762 0 net=3977
rlabel metal2 660 -1762 660 -1762 0 net=3102
rlabel metal2 744 -1762 744 -1762 0 net=7845
rlabel metal2 912 -1762 912 -1762 0 net=5723
rlabel metal2 1496 -1762 1496 -1762 0 net=12189
rlabel metal2 2340 -1762 2340 -1762 0 net=14377
rlabel metal2 79 -1764 79 -1764 0 net=3800
rlabel metal2 345 -1764 345 -1764 0 net=1737
rlabel metal2 387 -1764 387 -1764 0 net=4125
rlabel metal2 520 -1764 520 -1764 0 net=4525
rlabel metal2 667 -1764 667 -1764 0 net=5385
rlabel metal2 849 -1764 849 -1764 0 net=3925
rlabel metal2 891 -1764 891 -1764 0 net=10652
rlabel metal2 2004 -1764 2004 -1764 0 net=12313
rlabel metal2 79 -1766 79 -1766 0 net=5665
rlabel metal2 275 -1766 275 -1766 0 net=2007
rlabel metal2 352 -1766 352 -1766 0 net=2247
rlabel metal2 436 -1766 436 -1766 0 net=6737
rlabel metal2 548 -1766 548 -1766 0 net=6349
rlabel metal2 954 -1766 954 -1766 0 net=968
rlabel metal2 1556 -1766 1556 -1766 0 net=10085
rlabel metal2 1724 -1766 1724 -1766 0 net=11503
rlabel metal2 1934 -1766 1934 -1766 0 net=11933
rlabel metal2 2025 -1766 2025 -1766 0 net=12329
rlabel metal2 2249 -1766 2249 -1766 0 net=14431
rlabel metal2 149 -1768 149 -1768 0 net=2827
rlabel metal2 443 -1768 443 -1768 0 net=9771
rlabel metal2 1563 -1768 1563 -1768 0 net=9859
rlabel metal2 1598 -1768 1598 -1768 0 net=10077
rlabel metal2 1619 -1768 1619 -1768 0 net=10769
rlabel metal2 1773 -1768 1773 -1768 0 net=11747
rlabel metal2 1955 -1768 1955 -1768 0 net=12127
rlabel metal2 2042 -1768 2042 -1768 0 net=1
rlabel metal2 149 -1770 149 -1770 0 net=2649
rlabel metal2 268 -1770 268 -1770 0 net=1563
rlabel metal2 352 -1770 352 -1770 0 net=2549
rlabel metal2 481 -1770 481 -1770 0 net=8043
rlabel metal2 1465 -1770 1465 -1770 0 net=10741
rlabel metal2 1969 -1770 1969 -1770 0 net=12175
rlabel metal2 114 -1772 114 -1772 0 net=2161
rlabel metal2 359 -1772 359 -1772 0 net=3275
rlabel metal2 408 -1772 408 -1772 0 net=2431
rlabel metal2 492 -1772 492 -1772 0 net=4271
rlabel metal2 667 -1772 667 -1772 0 net=4043
rlabel metal2 695 -1772 695 -1772 0 net=13311
rlabel metal2 114 -1774 114 -1774 0 net=9493
rlabel metal2 1465 -1774 1465 -1774 0 net=10418
rlabel metal2 1787 -1774 1787 -1774 0 net=12281
rlabel metal2 275 -1776 275 -1776 0 net=2525
rlabel metal2 317 -1776 317 -1776 0 net=2091
rlabel metal2 415 -1776 415 -1776 0 net=3139
rlabel metal2 646 -1776 646 -1776 0 net=5205
rlabel metal2 968 -1776 968 -1776 0 net=11485
rlabel metal2 1927 -1776 1927 -1776 0 net=11875
rlabel metal2 1976 -1776 1976 -1776 0 net=12229
rlabel metal2 282 -1778 282 -1778 0 net=1575
rlabel metal2 590 -1778 590 -1778 0 net=4091
rlabel metal2 695 -1778 695 -1778 0 net=4573
rlabel metal2 733 -1778 733 -1778 0 net=6964
rlabel metal2 1045 -1778 1045 -1778 0 net=6811
rlabel metal2 1269 -1778 1269 -1778 0 net=8681
rlabel metal2 1479 -1778 1479 -1778 0 net=8915
rlabel metal2 1843 -1778 1843 -1778 0 net=11299
rlabel metal2 1878 -1778 1878 -1778 0 net=11673
rlabel metal2 1976 -1778 1976 -1778 0 net=13389
rlabel metal2 219 -1780 219 -1780 0 net=7761
rlabel metal2 1276 -1780 1276 -1780 0 net=11393
rlabel metal2 2123 -1780 2123 -1780 0 net=13169
rlabel metal2 191 -1782 191 -1782 0 net=3043
rlabel metal2 296 -1782 296 -1782 0 net=3253
rlabel metal2 674 -1782 674 -1782 0 net=5409
rlabel metal2 863 -1782 863 -1782 0 net=5623
rlabel metal2 1563 -1782 1563 -1782 0 net=11227
rlabel metal2 1857 -1782 1857 -1782 0 net=11455
rlabel metal2 2074 -1782 2074 -1782 0 net=12771
rlabel metal2 191 -1784 191 -1784 0 net=4017
rlabel metal2 492 -1784 492 -1784 0 net=2941
rlabel metal2 516 -1784 516 -1784 0 net=5647
rlabel metal2 1472 -1784 1472 -1784 0 net=9727
rlabel metal2 2074 -1784 2074 -1784 0 net=14285
rlabel metal2 261 -1786 261 -1786 0 net=2341
rlabel metal2 310 -1786 310 -1786 0 net=1629
rlabel metal2 453 -1786 453 -1786 0 net=4145
rlabel metal2 716 -1786 716 -1786 0 net=4725
rlabel metal2 758 -1786 758 -1786 0 net=6771
rlabel metal2 1430 -1786 1430 -1786 0 net=9191
rlabel metal2 1479 -1786 1479 -1786 0 net=9247
rlabel metal2 1507 -1786 1507 -1786 0 net=12094
rlabel metal2 2116 -1786 2116 -1786 0 net=13095
rlabel metal2 250 -1788 250 -1788 0 net=5351
rlabel metal2 310 -1788 310 -1788 0 net=4479
rlabel metal2 562 -1788 562 -1788 0 net=3076
rlabel metal2 625 -1788 625 -1788 0 net=4839
rlabel metal2 779 -1788 779 -1788 0 net=5059
rlabel metal2 877 -1788 877 -1788 0 net=6147
rlabel metal2 971 -1788 971 -1788 0 net=12831
rlabel metal2 100 -1790 100 -1790 0 net=1687
rlabel metal2 576 -1790 576 -1790 0 net=5531
rlabel metal2 803 -1790 803 -1790 0 net=5757
rlabel metal2 898 -1790 898 -1790 0 net=3877
rlabel metal2 1332 -1790 1332 -1790 0 net=9421
rlabel metal2 1570 -1790 1570 -1790 0 net=9871
rlabel metal2 1675 -1790 1675 -1790 0 net=10409
rlabel metal2 1948 -1790 1948 -1790 0 net=12047
rlabel metal2 2060 -1790 2060 -1790 0 net=12731
rlabel metal2 128 -1792 128 -1792 0 net=3541
rlabel metal2 625 -1792 625 -1792 0 net=5651
rlabel metal2 674 -1792 674 -1792 0 net=6945
rlabel metal2 719 -1792 719 -1792 0 net=11327
rlabel metal2 1346 -1792 1346 -1792 0 net=8765
rlabel metal2 1451 -1792 1451 -1792 0 net=9809
rlabel metal2 1661 -1792 1661 -1792 0 net=10307
rlabel metal2 1717 -1792 1717 -1792 0 net=12643
rlabel metal2 1920 -1792 1920 -1792 0 net=11783
rlabel metal2 2032 -1792 2032 -1792 0 net=12367
rlabel metal2 128 -1794 128 -1794 0 net=4215
rlabel metal2 464 -1794 464 -1794 0 net=4305
rlabel metal2 723 -1794 723 -1794 0 net=6167
rlabel metal2 1199 -1794 1199 -1794 0 net=8167
rlabel metal2 1346 -1794 1346 -1794 0 net=9965
rlabel metal2 1752 -1794 1752 -1794 0 net=11077
rlabel metal2 1822 -1794 1822 -1794 0 net=11265
rlabel metal2 1892 -1794 1892 -1794 0 net=11705
rlabel metal2 2032 -1794 2032 -1794 0 net=13771
rlabel metal2 177 -1796 177 -1796 0 net=5185
rlabel metal2 730 -1796 730 -1796 0 net=9567
rlabel metal2 1892 -1796 1892 -1796 0 net=12919
rlabel metal2 170 -1798 170 -1798 0 net=3401
rlabel metal2 201 -1798 201 -1798 0 net=7001
rlabel metal2 905 -1798 905 -1798 0 net=14403
rlabel metal2 156 -1800 156 -1800 0 net=2099
rlabel metal2 215 -1800 215 -1800 0 net=10549
rlabel metal2 2011 -1800 2011 -1800 0 net=12525
rlabel metal2 233 -1802 233 -1802 0 net=4459
rlabel metal2 499 -1802 499 -1802 0 net=2293
rlabel metal2 604 -1802 604 -1802 0 net=6938
rlabel metal2 933 -1802 933 -1802 0 net=11017
rlabel metal2 464 -1804 464 -1804 0 net=2865
rlabel metal2 478 -1804 478 -1804 0 net=4021
rlabel metal2 611 -1804 611 -1804 0 net=9021
rlabel metal2 1577 -1804 1577 -1804 0 net=9769
rlabel metal2 1962 -1804 1962 -1804 0 net=12151
rlabel metal2 72 -1806 72 -1806 0 net=3037
rlabel metal2 499 -1806 499 -1806 0 net=3207
rlabel metal2 936 -1806 936 -1806 0 net=6249
rlabel metal2 1024 -1806 1024 -1806 0 net=7097
rlabel metal2 1514 -1806 1514 -1806 0 net=9821
rlabel metal2 1710 -1806 1710 -1806 0 net=10755
rlabel metal2 72 -1808 72 -1808 0 net=2001
rlabel metal2 506 -1808 506 -1808 0 net=5989
rlabel metal2 940 -1808 940 -1808 0 net=13236
rlabel metal2 184 -1810 184 -1810 0 net=9981
rlabel metal2 541 -1810 541 -1810 0 net=7999
rlabel metal2 975 -1810 975 -1810 0 net=6221
rlabel metal2 1024 -1810 1024 -1810 0 net=9675
rlabel metal2 1381 -1810 1381 -1810 0 net=9311
rlabel metal2 1689 -1810 1689 -1810 0 net=10497
rlabel metal2 2186 -1810 2186 -1810 0 net=13931
rlabel metal2 401 -1812 401 -1812 0 net=3511
rlabel metal2 814 -1812 814 -1812 0 net=5341
rlabel metal2 975 -1812 975 -1812 0 net=7111
rlabel metal2 1136 -1812 1136 -1812 0 net=7597
rlabel metal2 1437 -1812 1437 -1812 0 net=10381
rlabel metal2 541 -1814 541 -1814 0 net=4815
rlabel metal2 786 -1814 786 -1814 0 net=5503
rlabel metal2 859 -1814 859 -1814 0 net=6553
rlabel metal2 1136 -1814 1136 -1814 0 net=7094
rlabel metal2 1318 -1814 1318 -1814 0 net=8837
rlabel metal2 555 -1816 555 -1816 0 net=3463
rlabel metal2 583 -1818 583 -1818 0 net=7599
rlabel metal2 772 -1818 772 -1818 0 net=3445
rlabel metal2 1178 -1818 1178 -1818 0 net=11143
rlabel metal2 786 -1820 786 -1820 0 net=7171
rlabel metal2 1339 -1820 1339 -1820 0 net=8205
rlabel metal2 800 -1822 800 -1822 0 net=12438
rlabel metal2 2193 -1822 2193 -1822 0 net=13437
rlabel metal2 1087 -1824 1087 -1824 0 net=6619
rlabel metal2 2067 -1824 2067 -1824 0 net=13975
rlabel metal2 1080 -1826 1080 -1826 0 net=6917
rlabel metal2 2144 -1826 2144 -1826 0 net=13211
rlabel metal2 2256 -1826 2256 -1826 0 net=13443
rlabel metal2 1080 -1828 1080 -1828 0 net=6695
rlabel metal2 2109 -1828 2109 -1828 0 net=13019
rlabel metal2 2368 -1828 2368 -1828 0 net=14527
rlabel metal2 1682 -1830 1682 -1830 0 net=10405
rlabel metal2 2277 -1830 2277 -1830 0 net=14199
rlabel metal2 1668 -1832 1668 -1832 0 net=10359
rlabel metal2 2214 -1832 2214 -1832 0 net=13651
rlabel metal2 1654 -1834 1654 -1834 0 net=10169
rlabel metal2 1906 -1834 1906 -1834 0 net=11763
rlabel metal2 1633 -1836 1633 -1836 0 net=10099
rlabel metal2 1864 -1836 1864 -1836 0 net=11475
rlabel metal2 1633 -1838 1633 -1838 0 net=11345
rlabel metal2 1766 -1840 1766 -1840 0 net=11523
rlabel metal2 1780 -1842 1780 -1842 0 net=11175
rlabel metal2 1395 -1844 1395 -1844 0 net=9283
rlabel metal2 1395 -1846 1395 -1846 0 net=8593
rlabel metal2 1416 -1848 1416 -1848 0 net=8839
rlabel metal2 30 -1859 30 -1859 0 net=2700
rlabel metal2 618 -1859 618 -1859 0 net=3978
rlabel metal2 1206 -1859 1206 -1859 0 net=10331
rlabel metal2 1636 -1859 1636 -1859 0 net=14200
rlabel metal2 30 -1861 30 -1861 0 net=2651
rlabel metal2 163 -1861 163 -1861 0 net=2051
rlabel metal2 163 -1861 163 -1861 0 net=2051
rlabel metal2 184 -1861 184 -1861 0 net=10410
rlabel metal2 2186 -1861 2186 -1861 0 net=13933
rlabel metal2 2186 -1861 2186 -1861 0 net=13933
rlabel metal2 2270 -1861 2270 -1861 0 net=11208
rlabel metal2 37 -1863 37 -1863 0 net=5845
rlabel metal2 632 -1863 632 -1863 0 net=860
rlabel metal2 1307 -1863 1307 -1863 0 net=10062
rlabel metal2 1664 -1863 1664 -1863 0 net=10406
rlabel metal2 2319 -1863 2319 -1863 0 net=13814
rlabel metal2 37 -1865 37 -1865 0 net=4019
rlabel metal2 194 -1865 194 -1865 0 net=395
rlabel metal2 635 -1865 635 -1865 0 net=7098
rlabel metal2 1206 -1865 1206 -1865 0 net=7581
rlabel metal2 1241 -1865 1241 -1865 0 net=8523
rlabel metal2 1276 -1865 1276 -1865 0 net=10756
rlabel metal2 2109 -1865 2109 -1865 0 net=13653
rlabel metal2 2319 -1865 2319 -1865 0 net=14521
rlabel metal2 47 -1867 47 -1867 0 net=10912
rlabel metal2 2368 -1867 2368 -1867 0 net=14467
rlabel metal2 72 -1869 72 -1869 0 net=2002
rlabel metal2 814 -1869 814 -1869 0 net=5343
rlabel metal2 814 -1869 814 -1869 0 net=5343
rlabel metal2 835 -1869 835 -1869 0 net=5387
rlabel metal2 835 -1869 835 -1869 0 net=5387
rlabel metal2 852 -1869 852 -1869 0 net=7598
rlabel metal2 1437 -1869 1437 -1869 0 net=13252
rlabel metal2 2410 -1869 2410 -1869 0 net=14773
rlabel metal2 72 -1871 72 -1871 0 net=4217
rlabel metal2 131 -1871 131 -1871 0 net=13929
rlabel metal2 89 -1873 89 -1873 0 net=9568
rlabel metal2 1734 -1873 1734 -1873 0 net=13438
rlabel metal2 100 -1875 100 -1875 0 net=1688
rlabel metal2 215 -1875 215 -1875 0 net=887
rlabel metal2 1332 -1875 1332 -1875 0 net=8169
rlabel metal2 1363 -1875 1363 -1875 0 net=10742
rlabel metal2 1962 -1875 1962 -1875 0 net=12049
rlabel metal2 2067 -1875 2067 -1875 0 net=13977
rlabel metal2 100 -1877 100 -1877 0 net=8682
rlabel metal2 1468 -1877 1468 -1877 0 net=13188
rlabel metal2 2221 -1877 2221 -1877 0 net=13663
rlabel metal2 107 -1879 107 -1879 0 net=3836
rlabel metal2 548 -1879 548 -1879 0 net=6350
rlabel metal2 1475 -1879 1475 -1879 0 net=12176
rlabel metal2 2256 -1879 2256 -1879 0 net=13445
rlabel metal2 107 -1881 107 -1881 0 net=3485
rlabel metal2 142 -1881 142 -1881 0 net=1948
rlabel metal2 1164 -1881 1164 -1881 0 net=7433
rlabel metal2 1241 -1881 1241 -1881 0 net=8131
rlabel metal2 1332 -1881 1332 -1881 0 net=8207
rlabel metal2 1353 -1881 1353 -1881 0 net=8389
rlabel metal2 1489 -1881 1489 -1881 0 net=9770
rlabel metal2 1622 -1881 1622 -1881 0 net=11674
rlabel metal2 2067 -1881 2067 -1881 0 net=12773
rlabel metal2 2249 -1881 2249 -1881 0 net=13805
rlabel metal2 103 -1883 103 -1883 0 net=4675
rlabel metal2 142 -1883 142 -1883 0 net=2249
rlabel metal2 401 -1883 401 -1883 0 net=3512
rlabel metal2 688 -1883 688 -1883 0 net=4146
rlabel metal2 737 -1883 737 -1883 0 net=9676
rlabel metal2 1059 -1883 1059 -1883 0 net=9375
rlabel metal2 1094 -1883 1094 -1883 0 net=3582
rlabel metal2 1773 -1883 1773 -1883 0 net=11749
rlabel metal2 2256 -1883 2256 -1883 0 net=13853
rlabel metal2 16 -1885 16 -1885 0 net=6841
rlabel metal2 1136 -1885 1136 -1885 0 net=11018
rlabel metal2 16 -1887 16 -1887 0 net=2551
rlabel metal2 373 -1887 373 -1887 0 net=8316
rlabel metal2 611 -1887 611 -1887 0 net=4307
rlabel metal2 688 -1887 688 -1887 0 net=7173
rlabel metal2 894 -1887 894 -1887 0 net=10324
rlabel metal2 124 -1889 124 -1889 0 net=6168
rlabel metal2 1129 -1889 1129 -1889 0 net=7417
rlabel metal2 1150 -1889 1150 -1889 0 net=7289
rlabel metal2 1209 -1889 1209 -1889 0 net=13312
rlabel metal2 128 -1891 128 -1891 0 net=6680
rlabel metal2 1080 -1891 1080 -1891 0 net=6697
rlabel metal2 1129 -1891 1129 -1891 0 net=5547
rlabel metal2 1164 -1891 1164 -1891 0 net=8990
rlabel metal2 1507 -1891 1507 -1891 0 net=13036
rlabel metal2 184 -1893 184 -1893 0 net=3045
rlabel metal2 233 -1893 233 -1893 0 net=13127
rlabel metal2 2228 -1893 2228 -1893 0 net=14665
rlabel metal2 177 -1895 177 -1895 0 net=3403
rlabel metal2 250 -1895 250 -1895 0 net=8766
rlabel metal2 1440 -1895 1440 -1895 0 net=14069
rlabel metal2 177 -1897 177 -1897 0 net=5353
rlabel metal2 275 -1897 275 -1897 0 net=2526
rlabel metal2 446 -1897 446 -1897 0 net=2866
rlabel metal2 478 -1897 478 -1897 0 net=9982
rlabel metal2 905 -1897 905 -1897 0 net=10079
rlabel metal2 1633 -1897 1633 -1897 0 net=11347
rlabel metal2 2032 -1897 2032 -1897 0 net=13773
rlabel metal2 205 -1899 205 -1899 0 net=2789
rlabel metal2 401 -1899 401 -1899 0 net=2141
rlabel metal2 646 -1899 646 -1899 0 net=7762
rlabel metal2 1290 -1899 1290 -1899 0 net=7971
rlabel metal2 1304 -1899 1304 -1899 0 net=13545
rlabel metal2 205 -1901 205 -1901 0 net=1577
rlabel metal2 303 -1901 303 -1901 0 net=1721
rlabel metal2 373 -1901 373 -1901 0 net=2911
rlabel metal2 908 -1901 908 -1901 0 net=5206
rlabel metal2 957 -1901 957 -1901 0 net=9728
rlabel metal2 1853 -1901 1853 -1901 0 net=14432
rlabel metal2 51 -1903 51 -1903 0 net=3057
rlabel metal2 303 -1903 303 -1903 0 net=3717
rlabel metal2 464 -1903 464 -1903 0 net=3543
rlabel metal2 541 -1903 541 -1903 0 net=4817
rlabel metal2 744 -1903 744 -1903 0 net=7847
rlabel metal2 1339 -1903 1339 -1903 0 net=8405
rlabel metal2 1381 -1903 1381 -1903 0 net=8841
rlabel metal2 1430 -1903 1430 -1903 0 net=9023
rlabel metal2 1458 -1903 1458 -1903 0 net=9193
rlabel metal2 1507 -1903 1507 -1903 0 net=9823
rlabel metal2 1605 -1903 1605 -1903 0 net=10043
rlabel metal2 1647 -1903 1647 -1903 0 net=12315
rlabel metal2 1864 -1903 1864 -1903 0 net=14322
rlabel metal2 51 -1905 51 -1905 0 net=9967
rlabel metal2 1664 -1905 1664 -1905 0 net=14216
rlabel metal2 2403 -1905 2403 -1905 0 net=14743
rlabel metal2 219 -1907 219 -1907 0 net=9621
rlabel metal2 1528 -1907 1528 -1907 0 net=9649
rlabel metal2 1528 -1907 1528 -1907 0 net=9649
rlabel metal2 1577 -1907 1577 -1907 0 net=9861
rlabel metal2 1773 -1907 1773 -1907 0 net=11145
rlabel metal2 1843 -1907 1843 -1907 0 net=12481
rlabel metal2 226 -1909 226 -1909 0 net=14507
rlabel metal2 170 -1911 170 -1911 0 net=2101
rlabel metal2 261 -1911 261 -1911 0 net=1565
rlabel metal2 275 -1911 275 -1911 0 net=3609
rlabel metal2 562 -1911 562 -1911 0 net=6818
rlabel metal2 1167 -1911 1167 -1911 0 net=14357
rlabel metal2 156 -1913 156 -1913 0 net=5237
rlabel metal2 394 -1913 394 -1913 0 net=3277
rlabel metal2 565 -1913 565 -1913 0 net=4614
rlabel metal2 1059 -1913 1059 -1913 0 net=9966
rlabel metal2 1353 -1913 1353 -1913 0 net=8617
rlabel metal2 1416 -1913 1416 -1913 0 net=9511
rlabel metal2 1584 -1913 1584 -1913 0 net=10771
rlabel metal2 1822 -1913 1822 -1913 0 net=11239
rlabel metal2 1850 -1913 1850 -1913 0 net=11395
rlabel metal2 1934 -1913 1934 -1913 0 net=11877
rlabel metal2 2032 -1913 2032 -1913 0 net=13021
rlabel metal2 170 -1915 170 -1915 0 net=11508
rlabel metal2 173 -1917 173 -1917 0 net=13353
rlabel metal2 229 -1919 229 -1919 0 net=11371
rlabel metal2 1864 -1919 1864 -1919 0 net=11457
rlabel metal2 1941 -1919 1941 -1919 0 net=13325
rlabel metal2 240 -1921 240 -1921 0 net=2613
rlabel metal2 422 -1921 422 -1921 0 net=3333
rlabel metal2 569 -1921 569 -1921 0 net=2294
rlabel metal2 744 -1921 744 -1921 0 net=5179
rlabel metal2 821 -1921 821 -1921 0 net=8091
rlabel metal2 943 -1921 943 -1921 0 net=7182
rlabel metal2 1227 -1921 1227 -1921 0 net=7231
rlabel metal2 1346 -1921 1346 -1921 0 net=9811
rlabel metal2 1591 -1921 1591 -1921 0 net=9285
rlabel metal2 1878 -1921 1878 -1921 0 net=11487
rlabel metal2 1941 -1921 1941 -1921 0 net=11935
rlabel metal2 2081 -1921 2081 -1921 0 net=12855
rlabel metal2 2 -1923 2 -1923 0 net=5839
rlabel metal2 422 -1923 422 -1923 0 net=6691
rlabel metal2 646 -1923 646 -1923 0 net=5625
rlabel metal2 919 -1923 919 -1923 0 net=5963
rlabel metal2 957 -1923 957 -1923 0 net=13865
rlabel metal2 2 -1925 2 -1925 0 net=2191
rlabel metal2 807 -1925 807 -1925 0 net=6451
rlabel metal2 1024 -1925 1024 -1925 0 net=6271
rlabel metal2 1444 -1925 1444 -1925 0 net=10785
rlabel metal2 1780 -1925 1780 -1925 0 net=11177
rlabel metal2 1899 -1925 1899 -1925 0 net=11537
rlabel metal2 159 -1927 159 -1927 0 net=6255
rlabel metal2 1038 -1927 1038 -1927 0 net=6555
rlabel metal2 1178 -1927 1178 -1927 0 net=12282
rlabel metal2 9 -1929 9 -1929 0 net=4138
rlabel metal2 429 -1929 429 -1929 0 net=3209
rlabel metal2 506 -1929 506 -1929 0 net=5990
rlabel metal2 863 -1929 863 -1929 0 net=7113
rlabel metal2 978 -1929 978 -1929 0 net=206
rlabel metal2 1913 -1929 1913 -1929 0 net=11785
rlabel metal2 1955 -1929 1955 -1929 0 net=12153
rlabel metal2 2074 -1929 2074 -1929 0 net=14287
rlabel metal2 9 -1931 9 -1931 0 net=12431
rlabel metal2 324 -1931 324 -1931 0 net=1869
rlabel metal2 506 -1931 506 -1931 0 net=5759
rlabel metal2 919 -1931 919 -1931 0 net=6918
rlabel metal2 1178 -1931 1178 -1931 0 net=9555
rlabel metal2 1696 -1931 1696 -1931 0 net=12015
rlabel metal2 1969 -1931 1969 -1931 0 net=12129
rlabel metal2 2011 -1931 2011 -1931 0 net=12369
rlabel metal2 2074 -1931 2074 -1931 0 net=12833
rlabel metal2 2137 -1931 2137 -1931 0 net=13213
rlabel metal2 58 -1933 58 -1933 0 net=6373
rlabel metal2 1062 -1933 1062 -1933 0 net=12190
rlabel metal2 23 -1935 23 -1935 0 net=6425
rlabel metal2 198 -1935 198 -1935 0 net=6307
rlabel metal2 1066 -1935 1066 -1935 0 net=5648
rlabel metal2 1696 -1935 1696 -1935 0 net=10429
rlabel metal2 1983 -1935 1983 -1935 0 net=12231
rlabel metal2 2060 -1935 2060 -1935 0 net=12733
rlabel metal2 2130 -1935 2130 -1935 0 net=13171
rlabel metal2 2298 -1935 2298 -1935 0 net=14083
rlabel metal2 23 -1937 23 -1937 0 net=9495
rlabel metal2 324 -1937 324 -1937 0 net=1807
rlabel metal2 1472 -1937 1472 -1937 0 net=2039
rlabel metal2 114 -1939 114 -1939 0 net=6773
rlabel metal2 828 -1939 828 -1939 0 net=6055
rlabel metal2 926 -1939 926 -1939 0 net=7959
rlabel metal2 1367 -1939 1367 -1939 0 net=8643
rlabel metal2 1444 -1939 1444 -1939 0 net=9249
rlabel metal2 1486 -1939 1486 -1939 0 net=9423
rlabel metal2 1703 -1939 1703 -1939 0 net=11423
rlabel metal2 1892 -1939 1892 -1939 0 net=12921
rlabel metal2 2312 -1939 2312 -1939 0 net=14147
rlabel metal2 432 -1941 432 -1941 0 net=6331
rlabel metal2 674 -1941 674 -1941 0 net=6947
rlabel metal2 695 -1941 695 -1941 0 net=4575
rlabel metal2 1066 -1941 1066 -1941 0 net=5867
rlabel metal2 1185 -1941 1185 -1941 0 net=8838
rlabel metal2 1335 -1941 1335 -1941 0 net=1
rlabel metal2 1451 -1941 1451 -1941 0 net=9873
rlabel metal2 1724 -1941 1724 -1941 0 net=11505
rlabel metal2 2347 -1941 2347 -1941 0 net=14379
rlabel metal2 191 -1943 191 -1943 0 net=5477
rlabel metal2 702 -1943 702 -1943 0 net=4238
rlabel metal2 961 -1943 961 -1943 0 net=6077
rlabel metal2 961 -1943 961 -1943 0 net=6077
rlabel metal2 975 -1943 975 -1943 0 net=10550
rlabel metal2 1766 -1943 1766 -1943 0 net=11525
rlabel metal2 1892 -1943 1892 -1943 0 net=13117
rlabel metal2 2179 -1943 2179 -1943 0 net=14543
rlabel metal2 450 -1945 450 -1945 0 net=4093
rlabel metal2 660 -1945 660 -1945 0 net=4273
rlabel metal2 702 -1945 702 -1945 0 net=6251
rlabel metal2 1073 -1945 1073 -1945 0 net=6515
rlabel metal2 1976 -1945 1976 -1945 0 net=13391
rlabel metal2 2179 -1945 2179 -1945 0 net=13415
rlabel metal2 121 -1947 121 -1947 0 net=9519
rlabel metal2 709 -1947 709 -1947 0 net=5187
rlabel metal2 982 -1947 982 -1947 0 net=6223
rlabel metal2 1087 -1947 1087 -1947 0 net=6621
rlabel metal2 1125 -1947 1125 -1947 0 net=11191
rlabel metal2 2004 -1947 2004 -1947 0 net=12331
rlabel metal2 86 -1949 86 -1949 0 net=6107
rlabel metal2 1111 -1949 1111 -1949 0 net=13449
rlabel metal2 121 -1951 121 -1951 0 net=2343
rlabel metal2 443 -1951 443 -1951 0 net=6703
rlabel metal2 1227 -1951 1227 -1951 0 net=13775
rlabel metal2 296 -1953 296 -1953 0 net=2093
rlabel metal2 443 -1953 443 -1953 0 net=3465
rlabel metal2 590 -1953 590 -1953 0 net=3673
rlabel metal2 772 -1953 772 -1953 0 net=3446
rlabel metal2 1248 -1953 1248 -1953 0 net=11329
rlabel metal2 2053 -1953 2053 -1953 0 net=12679
rlabel metal2 289 -1955 289 -1955 0 net=1769
rlabel metal2 653 -1955 653 -1955 0 net=4603
rlabel metal2 723 -1955 723 -1955 0 net=4823
rlabel metal2 772 -1955 772 -1955 0 net=5115
rlabel metal2 926 -1955 926 -1955 0 net=6813
rlabel metal2 1213 -1955 1213 -1955 0 net=7641
rlabel metal2 1395 -1955 1395 -1955 0 net=8595
rlabel metal2 1465 -1955 1465 -1955 0 net=9391
rlabel metal2 1654 -1955 1654 -1955 0 net=10101
rlabel metal2 1752 -1955 1752 -1955 0 net=11043
rlabel metal2 1766 -1955 1766 -1955 0 net=11117
rlabel metal2 2102 -1955 2102 -1955 0 net=13025
rlabel metal2 289 -1957 289 -1957 0 net=1589
rlabel metal2 933 -1957 933 -1957 0 net=8001
rlabel metal2 1360 -1957 1360 -1957 0 net=9019
rlabel metal2 1486 -1957 1486 -1957 0 net=11839
rlabel metal2 2151 -1957 2151 -1957 0 net=13341
rlabel metal2 359 -1959 359 -1959 0 net=2829
rlabel metal2 478 -1959 478 -1959 0 net=4023
rlabel metal2 653 -1959 653 -1959 0 net=5505
rlabel metal2 849 -1959 849 -1959 0 net=3879
rlabel metal2 933 -1959 933 -1959 0 net=5917
rlabel metal2 436 -1961 436 -1961 0 net=3255
rlabel metal2 604 -1961 604 -1961 0 net=4841
rlabel metal2 842 -1961 842 -1961 0 net=5411
rlabel metal2 1017 -1961 1017 -1961 0 net=6591
rlabel metal2 1213 -1961 1213 -1961 0 net=7831
rlabel metal2 1279 -1961 1279 -1961 0 net=11289
rlabel metal2 310 -1963 310 -1963 0 net=4481
rlabel metal2 1234 -1963 1234 -1963 0 net=8045
rlabel metal2 1360 -1963 1360 -1963 0 net=12997
rlabel metal2 310 -1965 310 -1965 0 net=1631
rlabel metal2 485 -1965 485 -1965 0 net=4461
rlabel metal2 576 -1965 576 -1965 0 net=5533
rlabel metal2 1297 -1965 1297 -1965 0 net=13473
rlabel metal2 212 -1967 212 -1967 0 net=4797
rlabel metal2 485 -1967 485 -1967 0 net=2943
rlabel metal2 513 -1967 513 -1967 0 net=697
rlabel metal2 1311 -1967 1311 -1967 0 net=7945
rlabel metal2 1675 -1967 1675 -1967 0 net=10309
rlabel metal2 1801 -1967 1801 -1967 0 net=13381
rlabel metal2 149 -1969 149 -1969 0 net=3171
rlabel metal2 247 -1969 247 -1969 0 net=5729
rlabel metal2 534 -1969 534 -1969 0 net=6739
rlabel metal2 625 -1969 625 -1969 0 net=5653
rlabel metal2 1549 -1969 1549 -1969 0 net=9741
rlabel metal2 1654 -1969 1654 -1969 0 net=10831
rlabel metal2 1801 -1969 1801 -1969 0 net=11267
rlabel metal2 86 -1971 86 -1971 0 net=9361
rlabel metal2 387 -1971 387 -1971 0 net=4127
rlabel metal2 576 -1971 576 -1971 0 net=5061
rlabel metal2 1524 -1971 1524 -1971 0 net=10887
rlabel metal2 93 -1973 93 -1973 0 net=2667
rlabel metal2 716 -1973 716 -1973 0 net=4727
rlabel metal2 751 -1973 751 -1973 0 net=4947
rlabel metal2 1535 -1973 1535 -1973 0 net=10471
rlabel metal2 93 -1975 93 -1975 0 net=2163
rlabel metal2 387 -1975 387 -1975 0 net=3141
rlabel metal2 457 -1975 457 -1975 0 net=2733
rlabel metal2 639 -1975 639 -1975 0 net=3875
rlabel metal2 793 -1975 793 -1975 0 net=5481
rlabel metal2 1549 -1975 1549 -1975 0 net=12314
rlabel metal2 79 -1977 79 -1977 0 net=5667
rlabel metal2 828 -1977 828 -1977 0 net=14333
rlabel metal2 79 -1979 79 -1979 0 net=4749
rlabel metal2 870 -1979 870 -1979 0 net=5613
rlabel metal2 1052 -1979 1052 -1979 0 net=8145
rlabel metal2 1661 -1979 1661 -1979 0 net=13096
rlabel metal2 254 -1981 254 -1981 0 net=7059
rlabel metal2 870 -1981 870 -1981 0 net=5725
rlabel metal2 1675 -1981 1675 -1981 0 net=10361
rlabel metal2 2326 -1981 2326 -1981 0 net=14247
rlabel metal2 44 -1983 44 -1983 0 net=5761
rlabel metal2 331 -1983 331 -1983 0 net=2383
rlabel metal2 345 -1983 345 -1983 0 net=2009
rlabel metal2 583 -1983 583 -1983 0 net=7601
rlabel metal2 1682 -1983 1682 -1983 0 net=10383
rlabel metal2 2361 -1983 2361 -1983 0 net=14405
rlabel metal2 44 -1985 44 -1985 0 net=5009
rlabel metal2 331 -1985 331 -1985 0 net=7891
rlabel metal2 1689 -1985 1689 -1985 0 net=10499
rlabel metal2 1787 -1985 1787 -1985 0 net=8917
rlabel metal2 65 -1987 65 -1987 0 net=8439
rlabel metal2 1563 -1987 1563 -1987 0 net=11229
rlabel metal2 345 -1989 345 -1989 0 net=1739
rlabel metal2 583 -1989 583 -1989 0 net=9551
rlabel metal2 1255 -1989 1255 -1989 0 net=7505
rlabel metal2 1283 -1989 1283 -1989 0 net=7915
rlabel metal2 1710 -1989 1710 -1989 0 net=10709
rlabel metal2 366 -1991 366 -1991 0 net=2433
rlabel metal2 1171 -1991 1171 -1991 0 net=7819
rlabel metal2 1374 -1991 1374 -1991 0 net=8563
rlabel metal2 1640 -1991 1640 -1991 0 net=10119
rlabel metal2 408 -1993 408 -1993 0 net=3039
rlabel metal2 765 -1993 765 -1993 0 net=4673
rlabel metal2 1192 -1993 1192 -1993 0 net=7529
rlabel metal2 1388 -1993 1388 -1993 0 net=7617
rlabel metal2 1556 -1993 1556 -1993 0 net=10087
rlabel metal2 471 -1995 471 -1995 0 net=4527
rlabel metal2 765 -1995 765 -1995 0 net=6477
rlabel metal2 1157 -1995 1157 -1995 0 net=7703
rlabel metal2 1514 -1995 1514 -1995 0 net=9313
rlabel metal2 520 -1997 520 -1997 0 net=4045
rlabel metal2 989 -1997 989 -1997 0 net=7039
rlabel metal2 1143 -1997 1143 -1997 0 net=7049
rlabel metal2 1514 -1997 1514 -1997 0 net=9773
rlabel metal2 635 -1999 635 -1999 0 net=2193
rlabel metal2 779 -1999 779 -1999 0 net=7003
rlabel metal2 1493 -1999 1493 -1999 0 net=10025
rlabel metal2 968 -2001 968 -2001 0 net=6149
rlabel metal2 1493 -2001 1493 -2001 0 net=11764
rlabel metal2 884 -2003 884 -2003 0 net=3927
rlabel metal2 2214 -2003 2214 -2003 0 net=13643
rlabel metal2 884 -2005 884 -2005 0 net=10171
rlabel metal2 2039 -2005 2039 -2005 0 net=13985
rlabel metal2 1668 -2007 1668 -2007 0 net=11079
rlabel metal2 2039 -2007 2039 -2007 0 net=12527
rlabel metal2 1794 -2009 1794 -2009 0 net=12203
rlabel metal2 2095 -2009 2095 -2009 0 net=14231
rlabel metal2 1808 -2011 1808 -2011 0 net=12397
rlabel metal2 2354 -2011 2354 -2011 0 net=14529
rlabel metal2 1808 -2013 1808 -2013 0 net=11301
rlabel metal2 1871 -2015 1871 -2015 0 net=11477
rlabel metal2 1906 -2017 1906 -2017 0 net=11707
rlabel metal2 1920 -2019 1920 -2019 0 net=12253
rlabel metal2 1717 -2021 1717 -2021 0 net=12645
rlabel metal2 779 -2023 779 -2023 0 net=10723
rlabel metal2 9 -2034 9 -2034 0 net=12432
rlabel metal2 800 -2034 800 -2034 0 net=3880
rlabel metal2 898 -2034 898 -2034 0 net=5654
rlabel metal2 1111 -2034 1111 -2034 0 net=7582
rlabel metal2 1230 -2034 1230 -2034 0 net=847
rlabel metal2 1335 -2034 1335 -2034 0 net=11192
rlabel metal2 2368 -2034 2368 -2034 0 net=14469
rlabel metal2 2368 -2034 2368 -2034 0 net=14469
rlabel metal2 2403 -2034 2403 -2034 0 net=14745
rlabel metal2 9 -2036 9 -2036 0 net=5011
rlabel metal2 51 -2036 51 -2036 0 net=8440
rlabel metal2 86 -2036 86 -2036 0 net=4677
rlabel metal2 138 -2036 138 -2036 0 net=4482
rlabel metal2 1024 -2036 1024 -2036 0 net=6273
rlabel metal2 1115 -2036 1115 -2036 0 net=6623
rlabel metal2 1115 -2036 1115 -2036 0 net=6623
rlabel metal2 1122 -2036 1122 -2036 0 net=8390
rlabel metal2 1437 -2036 1437 -2036 0 net=2040
rlabel metal2 37 -2038 37 -2038 0 net=4020
rlabel metal2 898 -2038 898 -2038 0 net=7961
rlabel metal2 1360 -2038 1360 -2038 0 net=10088
rlabel metal2 1713 -2038 1713 -2038 0 net=12130
rlabel metal2 37 -2040 37 -2040 0 net=5840
rlabel metal2 296 -2040 296 -2040 0 net=2094
rlabel metal2 1073 -2040 1073 -2040 0 net=6517
rlabel metal2 1297 -2040 1297 -2040 0 net=10472
rlabel metal2 1934 -2040 1934 -2040 0 net=11879
rlabel metal2 30 -2042 30 -2042 0 net=2652
rlabel metal2 296 -2042 296 -2042 0 net=4529
rlabel metal2 492 -2042 492 -2042 0 net=5731
rlabel metal2 1024 -2042 1024 -2042 0 net=9025
rlabel metal2 1437 -2042 1437 -2042 0 net=9251
rlabel metal2 1472 -2042 1472 -2042 0 net=11489
rlabel metal2 1969 -2042 1969 -2042 0 net=14509
rlabel metal2 16 -2044 16 -2044 0 net=2553
rlabel metal2 499 -2044 499 -2044 0 net=1871
rlabel metal2 569 -2044 569 -2044 0 net=6333
rlabel metal2 1150 -2044 1150 -2044 0 net=14070
rlabel metal2 2340 -2044 2340 -2044 0 net=14335
rlabel metal2 16 -2046 16 -2046 0 net=6453
rlabel metal2 828 -2046 828 -2046 0 net=8170
rlabel metal2 1430 -2046 1430 -2046 0 net=12233
rlabel metal2 2249 -2046 2249 -2046 0 net=13807
rlabel metal2 2298 -2046 2298 -2046 0 net=14085
rlabel metal2 30 -2048 30 -2048 0 net=4219
rlabel metal2 89 -2048 89 -2048 0 net=10172
rlabel metal2 919 -2048 919 -2048 0 net=6814
rlabel metal2 954 -2048 954 -2048 0 net=14530
rlabel metal2 44 -2050 44 -2050 0 net=4275
rlabel metal2 751 -2050 751 -2050 0 net=4949
rlabel metal2 922 -2050 922 -2050 0 net=7040
rlabel metal2 1087 -2050 1087 -2050 0 net=6705
rlabel metal2 1087 -2050 1087 -2050 0 net=6705
rlabel metal2 1153 -2050 1153 -2050 0 net=9020
rlabel metal2 1402 -2050 1402 -2050 0 net=8597
rlabel metal2 1440 -2050 1440 -2050 0 net=12922
rlabel metal2 2214 -2050 2214 -2050 0 net=13645
rlabel metal2 2 -2052 2 -2052 0 net=2192
rlabel metal2 1171 -2052 1171 -2052 0 net=4674
rlabel metal2 1363 -2052 1363 -2052 0 net=13774
rlabel metal2 51 -2054 51 -2054 0 net=10430
rlabel metal2 1766 -2054 1766 -2054 0 net=11119
rlabel metal2 58 -2056 58 -2056 0 net=6427
rlabel metal2 1384 -2056 1384 -2056 0 net=9742
rlabel metal2 1605 -2056 1605 -2056 0 net=9969
rlabel metal2 1808 -2056 1808 -2056 0 net=11303
rlabel metal2 2095 -2056 2095 -2056 0 net=14233
rlabel metal2 58 -2058 58 -2058 0 net=4647
rlabel metal2 100 -2058 100 -2058 0 net=3486
rlabel metal2 156 -2058 156 -2058 0 net=14358
rlabel metal2 65 -2060 65 -2060 0 net=6253
rlabel metal2 758 -2060 758 -2060 0 net=4824
rlabel metal2 807 -2060 807 -2060 0 net=8003
rlabel metal2 1402 -2060 1402 -2060 0 net=11506
rlabel metal2 2095 -2060 2095 -2060 0 net=13935
rlabel metal2 2228 -2060 2228 -2060 0 net=13447
rlabel metal2 2305 -2060 2305 -2060 0 net=14149
rlabel metal2 72 -2062 72 -2062 0 net=6079
rlabel metal2 1031 -2062 1031 -2062 0 net=5549
rlabel metal2 1178 -2062 1178 -2062 0 net=9557
rlabel metal2 1654 -2062 1654 -2062 0 net=10833
rlabel metal2 1815 -2062 1815 -2062 0 net=11291
rlabel metal2 2046 -2062 2046 -2062 0 net=12647
rlabel metal2 100 -2064 100 -2064 0 net=2205
rlabel metal2 1409 -2064 1409 -2064 0 net=11527
rlabel metal2 1920 -2064 1920 -2064 0 net=12255
rlabel metal2 2116 -2064 2116 -2064 0 net=13173
rlabel metal2 2172 -2064 2172 -2064 0 net=13393
rlabel metal2 2256 -2064 2256 -2064 0 net=13855
rlabel metal2 107 -2066 107 -2066 0 net=6819
rlabel metal2 1178 -2066 1178 -2066 0 net=7705
rlabel metal2 1220 -2066 1220 -2066 0 net=7435
rlabel metal2 1486 -2066 1486 -2066 0 net=11750
rlabel metal2 2074 -2066 2074 -2066 0 net=12835
rlabel metal2 2137 -2066 2137 -2066 0 net=13215
rlabel metal2 2186 -2066 2186 -2066 0 net=14381
rlabel metal2 156 -2068 156 -2068 0 net=7061
rlabel metal2 516 -2068 516 -2068 0 net=4576
rlabel metal2 1038 -2068 1038 -2068 0 net=6375
rlabel metal2 1192 -2068 1192 -2068 0 net=7973
rlabel metal2 1297 -2068 1297 -2068 0 net=7321
rlabel metal2 1486 -2068 1486 -2068 0 net=10102
rlabel metal2 1745 -2068 1745 -2068 0 net=10889
rlabel metal2 1871 -2068 1871 -2068 0 net=11479
rlabel metal2 1948 -2068 1948 -2068 0 net=12017
rlabel metal2 2018 -2068 2018 -2068 0 net=12399
rlabel metal2 2081 -2068 2081 -2068 0 net=12857
rlabel metal2 2207 -2068 2207 -2068 0 net=13547
rlabel metal2 2333 -2068 2333 -2068 0 net=14289
rlabel metal2 159 -2070 159 -2070 0 net=10080
rlabel metal2 1003 -2070 1003 -2070 0 net=7821
rlabel metal2 1269 -2070 1269 -2070 0 net=7233
rlabel metal2 173 -2072 173 -2072 0 net=8132
rlabel metal2 1276 -2072 1276 -2072 0 net=7849
rlabel metal2 1489 -2072 1489 -2072 0 net=13907
rlabel metal2 191 -2074 191 -2074 0 net=5760
rlabel metal2 569 -2074 569 -2074 0 net=5111
rlabel metal2 1038 -2074 1038 -2074 0 net=5869
rlabel metal2 1080 -2074 1080 -2074 0 net=6557
rlabel metal2 1234 -2074 1234 -2074 0 net=8047
rlabel metal2 1521 -2074 1521 -2074 0 net=10310
rlabel metal2 1843 -2074 1843 -2074 0 net=12483
rlabel metal2 191 -2076 191 -2076 0 net=1789
rlabel metal2 590 -2076 590 -2076 0 net=3674
rlabel metal2 670 -2076 670 -2076 0 net=5180
rlabel metal2 758 -2076 758 -2076 0 net=3461
rlabel metal2 891 -2076 891 -2076 0 net=5615
rlabel metal2 978 -2076 978 -2076 0 net=11240
rlabel metal2 1871 -2076 1871 -2076 0 net=11937
rlabel metal2 1955 -2076 1955 -2076 0 net=12155
rlabel metal2 170 -2078 170 -2078 0 net=3235
rlabel metal2 604 -2078 604 -2078 0 net=4842
rlabel metal2 786 -2078 786 -2078 0 net=9553
rlabel metal2 828 -2078 828 -2078 0 net=3929
rlabel metal2 989 -2078 989 -2078 0 net=6151
rlabel metal2 1283 -2078 1283 -2078 0 net=7531
rlabel metal2 1304 -2078 1304 -2078 0 net=9512
rlabel metal2 1521 -2078 1521 -2078 0 net=10045
rlabel metal2 1622 -2078 1622 -2078 0 net=13022
rlabel metal2 170 -2080 170 -2080 0 net=4819
rlabel metal2 740 -2080 740 -2080 0 net=12177
rlabel metal2 194 -2082 194 -2082 0 net=10187
rlabel metal2 1752 -2082 1752 -2082 0 net=11045
rlabel metal2 1899 -2082 1899 -2082 0 net=11539
rlabel metal2 1955 -2082 1955 -2082 0 net=14666
rlabel metal2 212 -2084 212 -2084 0 net=4798
rlabel metal2 331 -2084 331 -2084 0 net=7893
rlabel metal2 1059 -2084 1059 -2084 0 net=13991
rlabel metal2 2361 -2084 2361 -2084 0 net=14407
rlabel metal2 93 -2086 93 -2086 0 net=2165
rlabel metal2 338 -2086 338 -2086 0 net=2385
rlabel metal2 464 -2086 464 -2086 0 net=3545
rlabel metal2 618 -2086 618 -2086 0 net=5847
rlabel metal2 793 -2086 793 -2086 0 net=5483
rlabel metal2 940 -2086 940 -2086 0 net=5189
rlabel metal2 1066 -2086 1066 -2086 0 net=4385
rlabel metal2 1689 -2086 1689 -2086 0 net=10501
rlabel metal2 1773 -2086 1773 -2086 0 net=11147
rlabel metal2 1850 -2086 1850 -2086 0 net=11397
rlabel metal2 1906 -2086 1906 -2086 0 net=11709
rlabel metal2 2326 -2086 2326 -2086 0 net=14249
rlabel metal2 93 -2088 93 -2088 0 net=9392
rlabel metal2 1479 -2088 1479 -2088 0 net=9377
rlabel metal2 1780 -2088 1780 -2088 0 net=11179
rlabel metal2 2004 -2088 2004 -2088 0 net=12333
rlabel metal2 103 -2090 103 -2090 0 net=10617
rlabel metal2 1780 -2090 1780 -2090 0 net=11787
rlabel metal2 114 -2092 114 -2092 0 net=6775
rlabel metal2 835 -2092 835 -2092 0 net=5389
rlabel metal2 940 -2092 940 -2092 0 net=6109
rlabel metal2 1080 -2092 1080 -2092 0 net=6843
rlabel metal2 1143 -2092 1143 -2092 0 net=7005
rlabel metal2 1311 -2092 1311 -2092 0 net=7947
rlabel metal2 1451 -2092 1451 -2092 0 net=9875
rlabel metal2 1703 -2092 1703 -2092 0 net=11425
rlabel metal2 114 -2094 114 -2094 0 net=1723
rlabel metal2 366 -2094 366 -2094 0 net=2435
rlabel metal2 562 -2094 562 -2094 0 net=4463
rlabel metal2 653 -2094 653 -2094 0 net=5507
rlabel metal2 1094 -2094 1094 -2094 0 net=6699
rlabel metal2 1136 -2094 1136 -2094 0 net=7419
rlabel metal2 1332 -2094 1332 -2094 0 net=8209
rlabel metal2 1500 -2094 1500 -2094 0 net=9425
rlabel metal2 1626 -2094 1626 -2094 0 net=10333
rlabel metal2 1794 -2094 1794 -2094 0 net=12205
rlabel metal2 205 -2096 205 -2096 0 net=1579
rlabel metal2 404 -2096 404 -2096 0 net=2081
rlabel metal2 1010 -2096 1010 -2096 0 net=6257
rlabel metal2 1136 -2096 1136 -2096 0 net=7833
rlabel metal2 1325 -2096 1325 -2096 0 net=8525
rlabel metal2 1528 -2096 1528 -2096 0 net=9651
rlabel metal2 1703 -2096 1703 -2096 0 net=11459
rlabel metal2 177 -2098 177 -2098 0 net=5355
rlabel metal2 215 -2098 215 -2098 0 net=10205
rlabel metal2 1801 -2098 1801 -2098 0 net=11269
rlabel metal2 163 -2100 163 -2100 0 net=2053
rlabel metal2 219 -2100 219 -2100 0 net=9623
rlabel metal2 1143 -2100 1143 -2100 0 net=7665
rlabel metal2 1262 -2100 1262 -2100 0 net=7507
rlabel metal2 1332 -2100 1332 -2100 0 net=13930
rlabel metal2 124 -2102 124 -2102 0 net=1607
rlabel metal2 219 -2102 219 -2102 0 net=4895
rlabel metal2 2221 -2102 2221 -2102 0 net=13665
rlabel metal2 236 -2104 236 -2104 0 net=6948
rlabel metal2 688 -2104 688 -2104 0 net=7175
rlabel metal2 1353 -2104 1353 -2104 0 net=8619
rlabel metal2 1535 -2104 1535 -2104 0 net=12050
rlabel metal2 2179 -2104 2179 -2104 0 net=13417
rlabel metal2 247 -2106 247 -2106 0 net=9363
rlabel metal2 1927 -2106 1927 -2106 0 net=11841
rlabel metal2 2165 -2106 2165 -2106 0 net=13383
rlabel metal2 247 -2108 247 -2108 0 net=1591
rlabel metal2 303 -2108 303 -2108 0 net=3719
rlabel metal2 583 -2108 583 -2108 0 net=4309
rlabel metal2 625 -2108 625 -2108 0 net=2735
rlabel metal2 695 -2108 695 -2108 0 net=3549
rlabel metal2 1010 -2108 1010 -2108 0 net=6593
rlabel metal2 1164 -2108 1164 -2108 0 net=12071
rlabel metal2 2123 -2108 2123 -2108 0 net=13129
rlabel metal2 261 -2110 261 -2110 0 net=1567
rlabel metal2 338 -2110 338 -2110 0 net=1775
rlabel metal2 1563 -2110 1563 -2110 0 net=7917
rlabel metal2 2067 -2110 2067 -2110 0 net=12775
rlabel metal2 142 -2112 142 -2112 0 net=2251
rlabel metal2 275 -2112 275 -2112 0 net=3611
rlabel metal2 702 -2112 702 -2112 0 net=3617
rlabel metal2 1262 -2112 1262 -2112 0 net=7099
rlabel metal2 1538 -2112 1538 -2112 0 net=8231
rlabel metal2 2011 -2112 2011 -2112 0 net=12371
rlabel metal2 142 -2114 142 -2114 0 net=2573
rlabel metal2 1584 -2114 1584 -2114 0 net=10773
rlabel metal2 275 -2116 275 -2116 0 net=3335
rlabel metal2 597 -2116 597 -2116 0 net=6741
rlabel metal2 625 -2116 625 -2116 0 net=5535
rlabel metal2 863 -2116 863 -2116 0 net=7115
rlabel metal2 1367 -2116 1367 -2116 0 net=8645
rlabel metal2 1542 -2116 1542 -2116 0 net=10027
rlabel metal2 289 -2118 289 -2118 0 net=3143
rlabel metal2 422 -2118 422 -2118 0 net=6693
rlabel metal2 1164 -2118 1164 -2118 0 net=7291
rlabel metal2 1213 -2118 1213 -2118 0 net=3283
rlabel metal2 1549 -2118 1549 -2118 0 net=13654
rlabel metal2 226 -2120 226 -2120 0 net=2103
rlabel metal2 436 -2120 436 -2120 0 net=3257
rlabel metal2 653 -2120 653 -2120 0 net=13497
rlabel metal2 226 -2122 226 -2122 0 net=5627
rlabel metal2 660 -2122 660 -2122 0 net=9521
rlabel metal2 1636 -2122 1636 -2122 0 net=12101
rlabel metal2 2060 -2122 2060 -2122 0 net=12735
rlabel metal2 233 -2124 233 -2124 0 net=3405
rlabel metal2 443 -2124 443 -2124 0 net=3467
rlabel metal2 660 -2124 660 -2124 0 net=3951
rlabel metal2 1188 -2124 1188 -2124 0 net=11947
rlabel metal2 1339 -2124 1339 -2124 0 net=8407
rlabel metal2 1549 -2124 1549 -2124 0 net=8875
rlabel metal2 2060 -2124 2060 -2124 0 net=13987
rlabel metal2 303 -2126 303 -2126 0 net=1771
rlabel metal2 576 -2126 576 -2126 0 net=5063
rlabel metal2 891 -2126 891 -2126 0 net=4849
rlabel metal2 1633 -2126 1633 -2126 0 net=10711
rlabel metal2 2235 -2126 2235 -2126 0 net=13777
rlabel metal2 23 -2128 23 -2128 0 net=9497
rlabel metal2 2193 -2128 2193 -2128 0 net=13451
rlabel metal2 23 -2130 23 -2130 0 net=5541
rlabel metal2 310 -2130 310 -2130 0 net=1633
rlabel metal2 310 -2130 310 -2130 0 net=1633
rlabel metal2 345 -2130 345 -2130 0 net=1741
rlabel metal2 373 -2130 373 -2130 0 net=2913
rlabel metal2 555 -2130 555 -2130 0 net=5727
rlabel metal2 933 -2130 933 -2130 0 net=5919
rlabel metal2 1188 -2130 1188 -2130 0 net=11348
rlabel metal2 2151 -2130 2151 -2130 0 net=13343
rlabel metal2 131 -2132 131 -2132 0 net=1601
rlabel metal2 345 -2132 345 -2132 0 net=2143
rlabel metal2 443 -2132 443 -2132 0 net=6225
rlabel metal2 1199 -2132 1199 -2132 0 net=14522
rlabel metal2 149 -2134 149 -2134 0 net=3173
rlabel metal2 947 -2134 947 -2134 0 net=5965
rlabel metal2 1248 -2134 1248 -2134 0 net=7643
rlabel metal2 1381 -2134 1381 -2134 0 net=8843
rlabel metal2 1563 -2134 1563 -2134 0 net=11231
rlabel metal2 2151 -2134 2151 -2134 0 net=14545
rlabel metal2 54 -2136 54 -2136 0 net=1897
rlabel metal2 373 -2136 373 -2136 0 net=1939
rlabel metal2 1381 -2136 1381 -2136 0 net=12059
rlabel metal2 2144 -2136 2144 -2136 0 net=13327
rlabel metal2 394 -2138 394 -2138 0 net=2615
rlabel metal2 450 -2138 450 -2138 0 net=4094
rlabel metal2 639 -2138 639 -2138 0 net=5669
rlabel metal2 1157 -2138 1157 -2138 0 net=7051
rlabel metal2 1570 -2138 1570 -2138 0 net=10787
rlabel metal2 2088 -2138 2088 -2138 0 net=12999
rlabel metal2 79 -2140 79 -2140 0 net=4751
rlabel metal2 401 -2140 401 -2140 0 net=3040
rlabel metal2 492 -2140 492 -2140 0 net=8321
rlabel metal2 632 -2140 632 -2140 0 net=2701
rlabel metal2 1125 -2140 1125 -2140 0 net=8289
rlabel metal2 1458 -2140 1458 -2140 0 net=9195
rlabel metal2 1577 -2140 1577 -2140 0 net=9863
rlabel metal2 2039 -2140 2039 -2140 0 net=12529
rlabel metal2 79 -2142 79 -2142 0 net=2669
rlabel metal2 674 -2142 674 -2142 0 net=5479
rlabel metal2 1052 -2142 1052 -2142 0 net=8147
rlabel metal2 1584 -2142 1584 -2142 0 net=9287
rlabel metal2 1598 -2142 1598 -2142 0 net=10385
rlabel metal2 1787 -2142 1787 -2142 0 net=8919
rlabel metal2 121 -2144 121 -2144 0 net=2345
rlabel metal2 527 -2144 527 -2144 0 net=3279
rlabel metal2 709 -2144 709 -2144 0 net=4605
rlabel metal2 821 -2144 821 -2144 0 net=8093
rlabel metal2 1556 -2144 1556 -2144 0 net=9315
rlabel metal2 1605 -2144 1605 -2144 0 net=10363
rlabel metal2 1682 -2144 1682 -2144 0 net=11331
rlabel metal2 2396 -2144 2396 -2144 0 net=14775
rlabel metal2 135 -2146 135 -2146 0 net=2855
rlabel metal2 534 -2146 534 -2146 0 net=2903
rlabel metal2 1507 -2146 1507 -2146 0 net=9825
rlabel metal2 2102 -2146 2102 -2146 0 net=13027
rlabel metal2 254 -2148 254 -2148 0 net=5763
rlabel metal2 716 -2148 716 -2148 0 net=3876
rlabel metal2 842 -2148 842 -2148 0 net=5413
rlabel metal2 1052 -2148 1052 -2148 0 net=10120
rlabel metal2 2053 -2148 2053 -2148 0 net=12681
rlabel metal2 257 -2150 257 -2150 0 net=5261
rlabel metal2 1185 -2150 1185 -2150 0 net=12753
rlabel metal2 268 -2152 268 -2152 0 net=5239
rlabel metal2 723 -2152 723 -2152 0 net=4729
rlabel metal2 1185 -2152 1185 -2152 0 net=13866
rlabel metal2 268 -2154 268 -2154 0 net=3175
rlabel metal2 1374 -2154 1374 -2154 0 net=8565
rlabel metal2 1556 -2154 1556 -2154 0 net=10725
rlabel metal2 2200 -2154 2200 -2154 0 net=13475
rlabel metal2 408 -2156 408 -2156 0 net=2011
rlabel metal2 478 -2156 478 -2156 0 net=4025
rlabel metal2 730 -2156 730 -2156 0 net=6057
rlabel metal2 1230 -2156 1230 -2156 0 net=10259
rlabel metal2 2158 -2156 2158 -2156 0 net=13355
rlabel metal2 233 -2158 233 -2158 0 net=4543
rlabel metal2 513 -2158 513 -2158 0 net=4129
rlabel metal2 747 -2158 747 -2158 0 net=5451
rlabel metal2 1255 -2158 1255 -2158 0 net=7791
rlabel metal2 1647 -2158 1647 -2158 0 net=12317
rlabel metal2 282 -2160 282 -2160 0 net=3058
rlabel metal2 520 -2160 520 -2160 0 net=4047
rlabel metal2 765 -2160 765 -2160 0 net=6479
rlabel metal2 1647 -2160 1647 -2160 0 net=13978
rlabel metal2 282 -2162 282 -2162 0 net=1809
rlabel metal2 359 -2162 359 -2162 0 net=2831
rlabel metal2 765 -2162 765 -2162 0 net=5117
rlabel metal2 814 -2162 814 -2162 0 net=5345
rlabel metal2 877 -2162 877 -2162 0 net=1989
rlabel metal2 1668 -2162 1668 -2162 0 net=11081
rlabel metal2 1892 -2162 1892 -2162 0 net=13119
rlabel metal2 324 -2164 324 -2164 0 net=3211
rlabel metal2 667 -2164 667 -2164 0 net=2195
rlabel metal2 1346 -2164 1346 -2164 0 net=9813
rlabel metal2 1717 -2164 1717 -2164 0 net=10155
rlabel metal2 359 -2166 359 -2166 0 net=2945
rlabel metal2 499 -2166 499 -2166 0 net=3419
rlabel metal2 772 -2166 772 -2166 0 net=7603
rlabel metal2 1346 -2166 1346 -2166 0 net=7619
rlabel metal2 1496 -2166 1496 -2166 0 net=13719
rlabel metal2 198 -2168 198 -2168 0 net=6309
rlabel metal2 737 -2168 737 -2168 0 net=6393
rlabel metal2 1514 -2168 1514 -2168 0 net=9775
rlabel metal2 1836 -2168 1836 -2168 0 net=11373
rlabel metal2 184 -2170 184 -2170 0 net=3047
rlabel metal2 380 -2170 380 -2170 0 net=2791
rlabel metal2 429 -2170 429 -2170 0 net=4661
rlabel metal2 912 -2170 912 -2170 0 net=5703
rlabel metal2 1836 -2170 1836 -2170 0 net=13939
rlabel metal2 121 -2172 121 -2172 0 net=4735
rlabel metal2 737 -2172 737 -2172 0 net=3997
rlabel metal2 184 -2174 184 -2174 0 net=7399
rlabel metal2 1220 -2174 1220 -2174 0 net=8569
rlabel metal2 2 -2185 2 -2185 0 net=5765
rlabel metal2 744 -2185 744 -2185 0 net=6152
rlabel metal2 1258 -2185 1258 -2185 0 net=12648
rlabel metal2 2343 -2185 2343 -2185 0 net=14776
rlabel metal2 9 -2187 9 -2187 0 net=5012
rlabel metal2 54 -2187 54 -2187 0 net=6394
rlabel metal2 1398 -2187 1398 -2187 0 net=9864
rlabel metal2 1937 -2187 1937 -2187 0 net=13908
rlabel metal2 37 -2189 37 -2189 0 net=5671
rlabel metal2 1038 -2189 1038 -2189 0 net=5870
rlabel metal2 1227 -2189 1227 -2189 0 net=14150
rlabel metal2 51 -2191 51 -2191 0 net=5551
rlabel metal2 1080 -2191 1080 -2191 0 net=6845
rlabel metal2 1157 -2191 1157 -2191 0 net=8291
rlabel metal2 1405 -2191 1405 -2191 0 net=9252
rlabel metal2 1489 -2191 1489 -2191 0 net=11880
rlabel metal2 65 -2193 65 -2193 0 net=6254
rlabel metal2 1080 -2193 1080 -2193 0 net=6259
rlabel metal2 1115 -2193 1115 -2193 0 net=6624
rlabel metal2 1143 -2193 1143 -2193 0 net=7667
rlabel metal2 1293 -2193 1293 -2193 0 net=7234
rlabel metal2 2151 -2193 2151 -2193 0 net=14547
rlabel metal2 65 -2195 65 -2195 0 net=7177
rlabel metal2 1304 -2195 1304 -2195 0 net=8232
rlabel metal2 1969 -2195 1969 -2195 0 net=14511
rlabel metal2 93 -2197 93 -2197 0 net=6480
rlabel metal2 1496 -2197 1496 -2197 0 net=9378
rlabel metal2 1780 -2197 1780 -2197 0 net=11789
rlabel metal2 1836 -2197 1836 -2197 0 net=11939
rlabel metal2 1885 -2197 1885 -2197 0 net=11843
rlabel metal2 1969 -2197 1969 -2197 0 net=12207
rlabel metal2 2151 -2197 2151 -2197 0 net=13667
rlabel metal2 93 -2199 93 -2199 0 net=6428
rlabel metal2 1367 -2199 1367 -2199 0 net=13216
rlabel metal2 2228 -2199 2228 -2199 0 net=13448
rlabel metal2 96 -2201 96 -2201 0 net=5484
rlabel metal2 936 -2201 936 -2201 0 net=6594
rlabel metal2 1031 -2201 1031 -2201 0 net=5921
rlabel metal2 1094 -2201 1094 -2201 0 net=6701
rlabel metal2 1192 -2201 1192 -2201 0 net=7974
rlabel metal2 1304 -2201 1304 -2201 0 net=7949
rlabel metal2 1437 -2201 1437 -2201 0 net=8571
rlabel metal2 1521 -2201 1521 -2201 0 net=10047
rlabel metal2 1780 -2201 1780 -2201 0 net=11149
rlabel metal2 1860 -2201 1860 -2201 0 net=14470
rlabel metal2 107 -2203 107 -2203 0 net=6820
rlabel metal2 131 -2203 131 -2203 0 net=1455
rlabel metal2 296 -2203 296 -2203 0 net=4530
rlabel metal2 674 -2203 674 -2203 0 net=4503
rlabel metal2 1927 -2203 1927 -2203 0 net=12019
rlabel metal2 2032 -2203 2032 -2203 0 net=12683
rlabel metal2 107 -2205 107 -2205 0 net=3721
rlabel metal2 527 -2205 527 -2205 0 net=2856
rlabel metal2 1416 -2205 1416 -2205 0 net=8409
rlabel metal2 1521 -2205 1521 -2205 0 net=9523
rlabel metal2 1629 -2205 1629 -2205 0 net=13646
rlabel metal2 121 -2207 121 -2207 0 net=10561
rlabel metal2 1843 -2207 1843 -2207 0 net=11427
rlabel metal2 1962 -2207 1962 -2207 0 net=12179
rlabel metal2 2060 -2207 2060 -2207 0 net=13989
rlabel metal2 16 -2209 16 -2209 0 net=6455
rlabel metal2 124 -2209 124 -2209 0 net=2104
rlabel metal2 450 -2209 450 -2209 0 net=2346
rlabel metal2 506 -2209 506 -2209 0 net=4607
rlabel metal2 782 -2209 782 -2209 0 net=532
rlabel metal2 996 -2209 996 -2209 0 net=11541
rlabel metal2 1983 -2209 1983 -2209 0 net=12257
rlabel metal2 2060 -2209 2060 -2209 0 net=12837
rlabel metal2 16 -2211 16 -2211 0 net=4679
rlabel metal2 128 -2211 128 -2211 0 net=3281
rlabel metal2 1192 -2211 1192 -2211 0 net=7117
rlabel metal2 1332 -2211 1332 -2211 0 net=7620
rlabel metal2 1367 -2211 1367 -2211 0 net=8647
rlabel metal2 1545 -2211 1545 -2211 0 net=14290
rlabel metal2 86 -2213 86 -2213 0 net=5537
rlabel metal2 681 -2213 681 -2213 0 net=2737
rlabel metal2 800 -2213 800 -2213 0 net=9554
rlabel metal2 1202 -2213 1202 -2213 0 net=5181
rlabel metal2 1283 -2213 1283 -2213 0 net=11949
rlabel metal2 1381 -2213 1381 -2213 0 net=8876
rlabel metal2 1580 -2213 1580 -2213 0 net=13174
rlabel metal2 2130 -2213 2130 -2213 0 net=13549
rlabel metal2 138 -2215 138 -2215 0 net=13778
rlabel metal2 145 -2217 145 -2217 0 net=5480
rlabel metal2 877 -2217 877 -2217 0 net=1990
rlabel metal2 1517 -2217 1517 -2217 0 net=4531
rlabel metal2 166 -2219 166 -2219 0 net=13498
rlabel metal2 2256 -2219 2256 -2219 0 net=14235
rlabel metal2 236 -2221 236 -2221 0 net=6110
rlabel metal2 947 -2221 947 -2221 0 net=5415
rlabel metal2 947 -2221 947 -2221 0 net=5415
rlabel metal2 975 -2221 975 -2221 0 net=9364
rlabel metal2 1941 -2221 1941 -2221 0 net=12061
rlabel metal2 2025 -2221 2025 -2221 0 net=12531
rlabel metal2 2102 -2221 2102 -2221 0 net=13357
rlabel metal2 2207 -2221 2207 -2221 0 net=14087
rlabel metal2 243 -2223 243 -2223 0 net=3462
rlabel metal2 912 -2223 912 -2223 0 net=5705
rlabel metal2 1094 -2223 1094 -2223 0 net=6559
rlabel metal2 1185 -2223 1185 -2223 0 net=7101
rlabel metal2 1269 -2223 1269 -2223 0 net=7533
rlabel metal2 1342 -2223 1342 -2223 0 net=12234
rlabel metal2 1479 -2223 1479 -2223 0 net=8921
rlabel metal2 1871 -2223 1871 -2223 0 net=11711
rlabel metal2 1990 -2223 1990 -2223 0 net=12319
rlabel metal2 2088 -2223 2088 -2223 0 net=13131
rlabel metal2 2200 -2223 2200 -2223 0 net=13993
rlabel metal2 156 -2225 156 -2225 0 net=7063
rlabel metal2 1220 -2225 1220 -2225 0 net=13856
rlabel metal2 40 -2227 40 -2227 0 net=3911
rlabel metal2 250 -2227 250 -2227 0 net=7357
rlabel metal2 1227 -2227 1227 -2227 0 net=8095
rlabel metal2 1535 -2227 1535 -2227 0 net=9815
rlabel metal2 1759 -2227 1759 -2227 0 net=10891
rlabel metal2 1934 -2227 1934 -2227 0 net=7919
rlabel metal2 2186 -2227 2186 -2227 0 net=14383
rlabel metal2 289 -2229 289 -2229 0 net=3144
rlabel metal2 821 -2229 821 -2229 0 net=5263
rlabel metal2 940 -2229 940 -2229 0 net=5509
rlabel metal2 975 -2229 975 -2229 0 net=1115
rlabel metal2 1997 -2229 1997 -2229 0 net=12373
rlabel metal2 2116 -2229 2116 -2229 0 net=13419
rlabel metal2 289 -2231 289 -2231 0 net=1581
rlabel metal2 359 -2231 359 -2231 0 net=2946
rlabel metal2 1101 -2231 1101 -2231 0 net=6377
rlabel metal2 1136 -2231 1136 -2231 0 net=7835
rlabel metal2 1381 -2231 1381 -2231 0 net=8211
rlabel metal2 1549 -2231 1549 -2231 0 net=9317
rlabel metal2 1647 -2231 1647 -2231 0 net=14385
rlabel metal2 261 -2233 261 -2233 0 net=2253
rlabel metal2 457 -2233 457 -2233 0 net=2386
rlabel metal2 527 -2233 527 -2233 0 net=4311
rlabel metal2 590 -2233 590 -2233 0 net=3237
rlabel metal2 978 -2233 978 -2233 0 net=14553
rlabel metal2 100 -2235 100 -2235 0 net=2207
rlabel metal2 296 -2235 296 -2235 0 net=3547
rlabel metal2 618 -2235 618 -2235 0 net=4464
rlabel metal2 681 -2235 681 -2235 0 net=4027
rlabel metal2 726 -2235 726 -2235 0 net=13727
rlabel metal2 2186 -2235 2186 -2235 0 net=14747
rlabel metal2 100 -2237 100 -2237 0 net=5733
rlabel metal2 1115 -2237 1115 -2237 0 net=9971
rlabel metal2 1787 -2237 1787 -2237 0 net=11181
rlabel metal2 1934 -2237 1934 -2237 0 net=13384
rlabel metal2 2221 -2237 2221 -2237 0 net=13941
rlabel metal2 170 -2239 170 -2239 0 net=4821
rlabel metal2 492 -2239 492 -2239 0 net=6694
rlabel metal2 1129 -2239 1129 -2239 0 net=7293
rlabel metal2 1248 -2239 1248 -2239 0 net=7053
rlabel metal2 1423 -2239 1423 -2239 0 net=8599
rlabel metal2 1465 -2239 1465 -2239 0 net=9197
rlabel metal2 1591 -2239 1591 -2239 0 net=9877
rlabel metal2 1703 -2239 1703 -2239 0 net=11461
rlabel metal2 1948 -2239 1948 -2239 0 net=12073
rlabel metal2 2046 -2239 2046 -2239 0 net=14697
rlabel metal2 79 -2241 79 -2241 0 net=2671
rlabel metal2 555 -2241 555 -2241 0 net=5728
rlabel metal2 1248 -2241 1248 -2241 0 net=14273
rlabel metal2 79 -2243 79 -2243 0 net=5241
rlabel metal2 653 -2243 653 -2243 0 net=3687
rlabel metal2 1143 -2243 1143 -2243 0 net=6519
rlabel metal2 1255 -2243 1255 -2243 0 net=7793
rlabel metal2 1423 -2243 1423 -2243 0 net=8441
rlabel metal2 1570 -2243 1570 -2243 0 net=9777
rlabel metal2 1682 -2243 1682 -2243 0 net=11333
rlabel metal2 1857 -2243 1857 -2243 0 net=12403
rlabel metal2 2053 -2243 2053 -2243 0 net=12777
rlabel metal2 2179 -2243 2179 -2243 0 net=13809
rlabel metal2 170 -2245 170 -2245 0 net=2055
rlabel metal2 338 -2245 338 -2245 0 net=1777
rlabel metal2 576 -2245 576 -2245 0 net=3280
rlabel metal2 621 -2245 621 -2245 0 net=9795
rlabel metal2 1605 -2245 1605 -2245 0 net=10365
rlabel metal2 1703 -2245 1703 -2245 0 net=10503
rlabel metal2 1857 -2245 1857 -2245 0 net=11481
rlabel metal2 2067 -2245 2067 -2245 0 net=12859
rlabel metal2 177 -2247 177 -2247 0 net=2105
rlabel metal2 1766 -2247 1766 -2247 0 net=11047
rlabel metal2 2123 -2247 2123 -2247 0 net=13453
rlabel metal2 317 -2249 317 -2249 0 net=1569
rlabel metal2 352 -2249 352 -2249 0 net=1743
rlabel metal2 394 -2249 394 -2249 0 net=4753
rlabel metal2 583 -2249 583 -2249 0 net=3259
rlabel metal2 604 -2249 604 -2249 0 net=3551
rlabel metal2 709 -2249 709 -2249 0 net=5391
rlabel metal2 978 -2249 978 -2249 0 net=14421
rlabel metal2 275 -2251 275 -2251 0 net=3337
rlabel metal2 639 -2251 639 -2251 0 net=4851
rlabel metal2 912 -2251 912 -2251 0 net=5191
rlabel metal2 1073 -2251 1073 -2251 0 net=6335
rlabel metal2 1164 -2251 1164 -2251 0 net=7007
rlabel metal2 1262 -2251 1262 -2251 0 net=7851
rlabel metal2 1430 -2251 1430 -2251 0 net=8527
rlabel metal2 1605 -2251 1605 -2251 0 net=9559
rlabel metal2 1647 -2251 1647 -2251 0 net=10835
rlabel metal2 2074 -2251 2074 -2251 0 net=12401
rlabel metal2 275 -2253 275 -2253 0 net=1523
rlabel metal2 688 -2253 688 -2253 0 net=3613
rlabel metal2 828 -2253 828 -2253 0 net=3931
rlabel metal2 982 -2253 982 -2253 0 net=5967
rlabel metal2 1087 -2253 1087 -2253 0 net=6707
rlabel metal2 1178 -2253 1178 -2253 0 net=7707
rlabel metal2 1283 -2253 1283 -2253 0 net=7437
rlabel metal2 1339 -2253 1339 -2253 0 net=11377
rlabel metal2 2018 -2253 2018 -2253 0 net=12157
rlabel metal2 310 -2255 310 -2255 0 net=1635
rlabel metal2 324 -2255 324 -2255 0 net=3213
rlabel metal2 443 -2255 443 -2255 0 net=6227
rlabel metal2 961 -2255 961 -2255 0 net=7895
rlabel metal2 1178 -2255 1178 -2255 0 net=8049
rlabel metal2 1486 -2255 1486 -2255 0 net=11969
rlabel metal2 2018 -2255 2018 -2255 0 net=14251
rlabel metal2 114 -2257 114 -2257 0 net=1725
rlabel metal2 366 -2257 366 -2257 0 net=5269
rlabel metal2 695 -2257 695 -2257 0 net=4693
rlabel metal2 1318 -2257 1318 -2257 0 net=13028
rlabel metal2 114 -2259 114 -2259 0 net=5629
rlabel metal2 310 -2259 310 -2259 0 net=1873
rlabel metal2 590 -2259 590 -2259 0 net=3174
rlabel metal2 933 -2259 933 -2259 0 net=5453
rlabel metal2 989 -2259 989 -2259 0 net=11120
rlabel metal2 163 -2261 163 -2261 0 net=1609
rlabel metal2 380 -2261 380 -2261 0 net=4737
rlabel metal2 751 -2261 751 -2261 0 net=5849
rlabel metal2 1206 -2261 1206 -2261 0 net=7323
rlabel metal2 1339 -2261 1339 -2261 0 net=8149
rlabel metal2 1472 -2261 1472 -2261 0 net=11491
rlabel metal2 1500 -2261 1500 -2261 0 net=13328
rlabel metal2 163 -2263 163 -2263 0 net=14175
rlabel metal2 380 -2265 380 -2265 0 net=4731
rlabel metal2 856 -2265 856 -2265 0 net=11292
rlabel metal2 443 -2267 443 -2267 0 net=2555
rlabel metal2 478 -2267 478 -2267 0 net=4545
rlabel metal2 593 -2267 593 -2267 0 net=12754
rlabel metal2 142 -2269 142 -2269 0 net=2575
rlabel metal2 478 -2269 478 -2269 0 net=2591
rlabel metal2 1290 -2269 1290 -2269 0 net=10028
rlabel metal2 2039 -2269 2039 -2269 0 net=12737
rlabel metal2 142 -2271 142 -2271 0 net=2125
rlabel metal2 513 -2271 513 -2271 0 net=5029
rlabel metal2 1297 -2271 1297 -2271 0 net=7645
rlabel metal2 1370 -2271 1370 -2271 0 net=9987
rlabel metal2 1472 -2271 1472 -2271 0 net=9121
rlabel metal2 2109 -2271 2109 -2271 0 net=13395
rlabel metal2 513 -2273 513 -2273 0 net=2905
rlabel metal2 541 -2273 541 -2273 0 net=2915
rlabel metal2 737 -2273 737 -2273 0 net=3999
rlabel metal2 758 -2273 758 -2273 0 net=10193
rlabel metal2 1808 -2273 1808 -2273 0 net=12103
rlabel metal2 2095 -2273 2095 -2273 0 net=13937
rlabel metal2 422 -2275 422 -2275 0 net=3407
rlabel metal2 548 -2275 548 -2275 0 net=4049
rlabel metal2 758 -2275 758 -2275 0 net=5065
rlabel metal2 1353 -2275 1353 -2275 0 net=8621
rlabel metal2 1563 -2275 1563 -2275 0 net=11233
rlabel metal2 2011 -2275 2011 -2275 0 net=12485
rlabel metal2 2095 -2275 2095 -2275 0 net=13345
rlabel metal2 184 -2277 184 -2277 0 net=7401
rlabel metal2 765 -2277 765 -2277 0 net=5119
rlabel metal2 1059 -2277 1059 -2277 0 net=9625
rlabel metal2 1563 -2277 1563 -2277 0 net=9653
rlabel metal2 1661 -2277 1661 -2277 0 net=10261
rlabel metal2 1892 -2277 1892 -2277 0 net=11375
rlabel metal2 2081 -2277 2081 -2277 0 net=13121
rlabel metal2 149 -2279 149 -2279 0 net=1899
rlabel metal2 219 -2279 219 -2279 0 net=4897
rlabel metal2 485 -2279 485 -2279 0 net=6311
rlabel metal2 772 -2279 772 -2279 0 net=7605
rlabel metal2 814 -2279 814 -2279 0 net=2197
rlabel metal2 1059 -2279 1059 -2279 0 net=6083
rlabel metal2 1374 -2279 1374 -2279 0 net=8845
rlabel metal2 1619 -2279 1619 -2279 0 net=9499
rlabel metal2 1738 -2279 1738 -2279 0 net=10775
rlabel metal2 135 -2281 135 -2281 0 net=4715
rlabel metal2 191 -2281 191 -2281 0 net=1791
rlabel metal2 373 -2281 373 -2281 0 net=1940
rlabel metal2 786 -2281 786 -2281 0 net=14677
rlabel metal2 135 -2283 135 -2283 0 net=5113
rlabel metal2 611 -2283 611 -2283 0 net=6743
rlabel metal2 828 -2283 828 -2283 0 net=5347
rlabel metal2 859 -2283 859 -2283 0 net=13585
rlabel metal2 191 -2285 191 -2285 0 net=4387
rlabel metal2 1321 -2285 1321 -2285 0 net=13829
rlabel metal2 373 -2287 373 -2287 0 net=2833
rlabel metal2 569 -2287 569 -2287 0 net=4131
rlabel metal2 786 -2287 786 -2287 0 net=7823
rlabel metal2 1066 -2287 1066 -2287 0 net=6275
rlabel metal2 1395 -2287 1395 -2287 0 net=1485
rlabel metal2 415 -2289 415 -2289 0 net=2793
rlabel metal2 646 -2289 646 -2289 0 net=3469
rlabel metal2 807 -2289 807 -2289 0 net=8005
rlabel metal2 968 -2289 968 -2289 0 net=2082
rlabel metal2 1619 -2289 1619 -2289 0 net=10157
rlabel metal2 1794 -2289 1794 -2289 0 net=11271
rlabel metal2 331 -2291 331 -2291 0 net=2167
rlabel metal2 436 -2291 436 -2291 0 net=2617
rlabel metal2 499 -2291 499 -2291 0 net=3421
rlabel metal2 646 -2291 646 -2291 0 net=3953
rlabel metal2 723 -2291 723 -2291 0 net=9075
rlabel metal2 1052 -2291 1052 -2291 0 net=12657
rlabel metal2 1402 -2291 1402 -2291 0 net=13563
rlabel metal2 233 -2293 233 -2293 0 net=4353
rlabel metal2 562 -2293 562 -2293 0 net=8323
rlabel metal2 1409 -2293 1409 -2293 0 net=11529
rlabel metal2 233 -2295 233 -2295 0 net=4181
rlabel metal2 730 -2295 730 -2295 0 net=6059
rlabel metal2 1409 -2295 1409 -2295 0 net=8191
rlabel metal2 1633 -2295 1633 -2295 0 net=10713
rlabel metal2 268 -2297 268 -2297 0 net=3177
rlabel metal2 730 -2297 730 -2297 0 net=7963
rlabel metal2 905 -2297 905 -2297 0 net=5617
rlabel metal2 1444 -2297 1444 -2297 0 net=9289
rlabel metal2 1633 -2297 1633 -2297 0 net=10189
rlabel metal2 205 -2299 205 -2299 0 net=5357
rlabel metal2 905 -2299 905 -2299 0 net=7509
rlabel metal2 1584 -2299 1584 -2299 0 net=9827
rlabel metal2 44 -2301 44 -2301 0 net=4277
rlabel metal2 212 -2301 212 -2301 0 net=1603
rlabel metal2 331 -2301 331 -2301 0 net=2145
rlabel metal2 429 -2301 429 -2301 0 net=4663
rlabel metal2 747 -2301 747 -2301 0 net=5633
rlabel metal2 1024 -2301 1024 -2301 0 net=9027
rlabel metal2 44 -2303 44 -2303 0 net=4649
rlabel metal2 72 -2303 72 -2303 0 net=6081
rlabel metal2 1325 -2303 1325 -2303 0 net=9427
rlabel metal2 1640 -2303 1640 -2303 0 net=10207
rlabel metal2 23 -2305 23 -2305 0 net=5543
rlabel metal2 72 -2305 72 -2305 0 net=2303
rlabel metal2 807 -2305 807 -2305 0 net=4951
rlabel metal2 1507 -2305 1507 -2305 0 net=8567
rlabel metal2 1650 -2305 1650 -2305 0 net=12334
rlabel metal2 23 -2307 23 -2307 0 net=3049
rlabel metal2 212 -2307 212 -2307 0 net=1593
rlabel metal2 282 -2307 282 -2307 0 net=1811
rlabel metal2 401 -2307 401 -2307 0 net=2437
rlabel metal2 835 -2307 835 -2307 0 net=3285
rlabel metal2 1507 -2307 1507 -2307 0 net=10727
rlabel metal2 1675 -2307 1675 -2307 0 net=10335
rlabel metal2 2277 -2307 2277 -2307 0 net=13721
rlabel metal2 198 -2309 198 -2309 0 net=1849
rlabel metal2 793 -2309 793 -2309 0 net=6777
rlabel metal2 1556 -2309 1556 -2309 0 net=10387
rlabel metal2 1731 -2309 1731 -2309 0 net=13001
rlabel metal2 2277 -2309 2277 -2309 0 net=14409
rlabel metal2 247 -2311 247 -2311 0 net=468
rlabel metal2 464 -2311 464 -2311 0 net=2703
rlabel metal2 789 -2311 789 -2311 0 net=9999
rlabel metal2 1745 -2311 1745 -2311 0 net=10789
rlabel metal2 2144 -2311 2144 -2311 0 net=13477
rlabel metal2 282 -2313 282 -2313 0 net=1773
rlabel metal2 387 -2313 387 -2313 0 net=1931
rlabel metal2 793 -2313 793 -2313 0 net=4655
rlabel metal2 1801 -2313 1801 -2313 0 net=11305
rlabel metal2 2242 -2313 2242 -2313 0 net=14337
rlabel metal2 303 -2315 303 -2315 0 net=2013
rlabel metal2 632 -2315 632 -2315 0 net=3619
rlabel metal2 849 -2315 849 -2315 0 net=7421
rlabel metal2 1773 -2315 1773 -2315 0 net=10619
rlabel metal2 30 -2317 30 -2317 0 net=4221
rlabel metal2 660 -2317 660 -2317 0 net=8013
rlabel metal2 1773 -2317 1773 -2317 0 net=11083
rlabel metal2 702 -2319 702 -2319 0 net=10247
rlabel metal2 1829 -2319 1829 -2319 0 net=11399
rlabel metal2 1199 -2321 1199 -2321 0 net=11861
rlabel metal2 33 -2323 33 -2323 0 net=13709
rlabel metal2 5 -2334 5 -2334 0 net=7178
rlabel metal2 163 -2334 163 -2334 0 net=6082
rlabel metal2 1038 -2334 1038 -2334 0 net=7054
rlabel metal2 1363 -2334 1363 -2334 0 net=13942
rlabel metal2 2326 -2334 2326 -2334 0 net=13722
rlabel metal2 9 -2336 9 -2336 0 net=967
rlabel metal2 905 -2336 905 -2336 0 net=7510
rlabel metal2 1272 -2336 1272 -2336 0 net=12158
rlabel metal2 2165 -2336 2165 -2336 0 net=7920
rlabel metal2 23 -2338 23 -2338 0 net=3050
rlabel metal2 170 -2338 170 -2338 0 net=2057
rlabel metal2 226 -2338 226 -2338 0 net=1610
rlabel metal2 597 -2338 597 -2338 0 net=3338
rlabel metal2 782 -2338 782 -2338 0 net=9816
rlabel metal2 1542 -2338 1542 -2338 0 net=10620
rlabel metal2 1892 -2338 1892 -2338 0 net=12075
rlabel metal2 1976 -2338 1976 -2338 0 net=12739
rlabel metal2 2165 -2338 2165 -2338 0 net=13831
rlabel metal2 2221 -2338 2221 -2338 0 net=14339
rlabel metal2 16 -2340 16 -2340 0 net=4681
rlabel metal2 240 -2340 240 -2340 0 net=7805
rlabel metal2 618 -2340 618 -2340 0 net=65
rlabel metal2 1374 -2340 1374 -2340 0 net=8847
rlabel metal2 1398 -2340 1398 -2340 0 net=8192
rlabel metal2 1493 -2340 1493 -2340 0 net=12402
rlabel metal2 2242 -2340 2242 -2340 0 net=14423
rlabel metal2 16 -2342 16 -2342 0 net=5672
rlabel metal2 51 -2342 51 -2342 0 net=5553
rlabel metal2 1041 -2342 1041 -2342 0 net=9745
rlabel metal2 1517 -2342 1517 -2342 0 net=11790
rlabel metal2 1934 -2342 1934 -2342 0 net=14384
rlabel metal2 30 -2344 30 -2344 0 net=6260
rlabel metal2 1108 -2344 1108 -2344 0 net=12658
rlabel metal2 2039 -2344 2039 -2344 0 net=13133
rlabel metal2 2186 -2344 2186 -2344 0 net=14749
rlabel metal2 33 -2346 33 -2346 0 net=4650
rlabel metal2 51 -2346 51 -2346 0 net=9797
rlabel metal2 1580 -2346 1580 -2346 0 net=14236
rlabel metal2 44 -2348 44 -2348 0 net=5631
rlabel metal2 170 -2348 170 -2348 0 net=2107
rlabel metal2 243 -2348 243 -2348 0 net=4608
rlabel metal2 569 -2348 569 -2348 0 net=4133
rlabel metal2 625 -2348 625 -2348 0 net=6229
rlabel metal2 905 -2348 905 -2348 0 net=5511
rlabel metal2 954 -2348 954 -2348 0 net=3238
rlabel metal2 1377 -2348 1377 -2348 0 net=8600
rlabel metal2 1542 -2348 1542 -2348 0 net=10001
rlabel metal2 1682 -2348 1682 -2348 0 net=13990
rlabel metal2 2235 -2348 2235 -2348 0 net=14411
rlabel metal2 65 -2350 65 -2350 0 net=1525
rlabel metal2 282 -2350 282 -2350 0 net=1774
rlabel metal2 1080 -2350 1080 -2350 0 net=8568
rlabel metal2 1682 -2350 1682 -2350 0 net=10791
rlabel metal2 1850 -2350 1850 -2350 0 net=11463
rlabel metal2 1878 -2350 1878 -2350 0 net=13359
rlabel metal2 2179 -2350 2179 -2350 0 net=13811
rlabel metal2 2193 -2350 2193 -2350 0 net=14089
rlabel metal2 2228 -2350 2228 -2350 0 net=14387
rlabel metal2 114 -2352 114 -2352 0 net=2209
rlabel metal2 275 -2352 275 -2352 0 net=1933
rlabel metal2 408 -2352 408 -2352 0 net=4223
rlabel metal2 775 -2352 775 -2352 0 net=8249
rlabel metal2 978 -2352 978 -2352 0 net=6778
rlabel metal2 1248 -2352 1248 -2352 0 net=7853
rlabel metal2 1276 -2352 1276 -2352 0 net=5182
rlabel metal2 1451 -2352 1451 -2352 0 net=9627
rlabel metal2 1685 -2352 1685 -2352 0 net=13564
rlabel metal2 2207 -2352 2207 -2352 0 net=14127
rlabel metal2 166 -2354 166 -2354 0 net=14007
rlabel metal2 2256 -2354 2256 -2354 0 net=14555
rlabel metal2 247 -2356 247 -2356 0 net=8006
rlabel metal2 859 -2356 859 -2356 0 net=10313
rlabel metal2 1745 -2356 1745 -2356 0 net=11085
rlabel metal2 1850 -2356 1850 -2356 0 net=11845
rlabel metal2 1895 -2356 1895 -2356 0 net=13938
rlabel metal2 2263 -2356 2263 -2356 0 net=14679
rlabel metal2 247 -2358 247 -2358 0 net=2593
rlabel metal2 481 -2358 481 -2358 0 net=865
rlabel metal2 1773 -2358 1773 -2358 0 net=11183
rlabel metal2 1885 -2358 1885 -2358 0 net=12063
rlabel metal2 1948 -2358 1948 -2358 0 net=13421
rlabel metal2 254 -2360 254 -2360 0 net=2127
rlabel metal2 254 -2360 254 -2360 0 net=2127
rlabel metal2 261 -2360 261 -2360 0 net=2439
rlabel metal2 408 -2360 408 -2360 0 net=2619
rlabel metal2 492 -2360 492 -2360 0 net=2673
rlabel metal2 527 -2360 527 -2360 0 net=4313
rlabel metal2 576 -2360 576 -2360 0 net=4547
rlabel metal2 786 -2360 786 -2360 0 net=7824
rlabel metal2 982 -2360 982 -2360 0 net=9077
rlabel metal2 1055 -2360 1055 -2360 0 net=11492
rlabel metal2 1528 -2360 1528 -2360 0 net=9879
rlabel metal2 1787 -2360 1787 -2360 0 net=11429
rlabel metal2 1853 -2360 1853 -2360 0 net=1
rlabel metal2 2011 -2360 2011 -2360 0 net=12487
rlabel metal2 282 -2362 282 -2362 0 net=3287
rlabel metal2 842 -2362 842 -2362 0 net=5193
rlabel metal2 919 -2362 919 -2362 0 net=9500
rlabel metal2 1843 -2362 1843 -2362 0 net=11483
rlabel metal2 1906 -2362 1906 -2362 0 net=12021
rlabel metal2 1934 -2362 1934 -2362 0 net=12375
rlabel metal2 2011 -2362 2011 -2362 0 net=12861
rlabel metal2 2088 -2362 2088 -2362 0 net=14549
rlabel metal2 296 -2364 296 -2364 0 net=3548
rlabel metal2 730 -2364 730 -2364 0 net=7965
rlabel metal2 1486 -2364 1486 -2364 0 net=9779
rlabel metal2 1591 -2364 1591 -2364 0 net=11379
rlabel metal2 1836 -2364 1836 -2364 0 net=11941
rlabel metal2 1927 -2364 1927 -2364 0 net=12321
rlabel metal2 1997 -2364 1997 -2364 0 net=12839
rlabel metal2 2102 -2364 2102 -2364 0 net=13551
rlabel metal2 2305 -2364 2305 -2364 0 net=4533
rlabel metal2 191 -2366 191 -2366 0 net=4389
rlabel metal2 730 -2366 730 -2366 0 net=4657
rlabel metal2 796 -2366 796 -2366 0 net=10194
rlabel metal2 1678 -2366 1678 -2366 0 net=10693
rlabel metal2 1836 -2366 1836 -2366 0 net=12259
rlabel metal2 1990 -2366 1990 -2366 0 net=13455
rlabel metal2 72 -2368 72 -2368 0 net=2305
rlabel metal2 296 -2368 296 -2368 0 net=6061
rlabel metal2 1108 -2368 1108 -2368 0 net=6847
rlabel metal2 1262 -2368 1262 -2368 0 net=7951
rlabel metal2 1318 -2368 1318 -2368 0 net=8213
rlabel metal2 1668 -2368 1668 -2368 0 net=10777
rlabel metal2 1983 -2368 1983 -2368 0 net=12779
rlabel metal2 2060 -2368 2060 -2368 0 net=13397
rlabel metal2 2123 -2368 2123 -2368 0 net=13587
rlabel metal2 310 -2370 310 -2370 0 net=1875
rlabel metal2 457 -2370 457 -2370 0 net=4822
rlabel metal2 859 -2370 859 -2370 0 net=7836
rlabel metal2 1381 -2370 1381 -2370 0 net=8573
rlabel metal2 1738 -2370 1738 -2370 0 net=11049
rlabel metal2 1969 -2370 1969 -2370 0 net=12209
rlabel metal2 2137 -2370 2137 -2370 0 net=13669
rlabel metal2 268 -2372 268 -2372 0 net=1605
rlabel metal2 317 -2372 317 -2372 0 net=1637
rlabel metal2 317 -2372 317 -2372 0 net=1637
rlabel metal2 387 -2372 387 -2372 0 net=6531
rlabel metal2 863 -2372 863 -2372 0 net=2199
rlabel metal2 1052 -2372 1052 -2372 0 net=13537
rlabel metal2 2151 -2372 2151 -2372 0 net=13729
rlabel metal2 401 -2374 401 -2374 0 net=4029
rlabel metal2 716 -2374 716 -2374 0 net=7403
rlabel metal2 2172 -2374 2172 -2374 0 net=13995
rlabel metal2 37 -2376 37 -2376 0 net=14107
rlabel metal2 100 -2378 100 -2378 0 net=5735
rlabel metal2 786 -2378 786 -2378 0 net=7009
rlabel metal2 1227 -2378 1227 -2378 0 net=8097
rlabel metal2 1437 -2378 1437 -2378 0 net=9291
rlabel metal2 1766 -2378 1766 -2378 0 net=11401
rlabel metal2 2018 -2378 2018 -2378 0 net=14253
rlabel metal2 100 -2380 100 -2380 0 net=5455
rlabel metal2 1087 -2380 1087 -2380 0 net=7897
rlabel metal2 1227 -2380 1227 -2380 0 net=7795
rlabel metal2 1276 -2380 1276 -2380 0 net=8787
rlabel metal2 1647 -2380 1647 -2380 0 net=10837
rlabel metal2 2046 -2380 2046 -2380 0 net=14699
rlabel metal2 422 -2382 422 -2382 0 net=4898
rlabel metal2 821 -2382 821 -2382 0 net=3614
rlabel metal2 1087 -2382 1087 -2382 0 net=7295
rlabel metal2 1136 -2382 1136 -2382 0 net=7646
rlabel metal2 1444 -2382 1444 -2382 0 net=8923
rlabel metal2 1549 -2382 1549 -2382 0 net=9319
rlabel metal2 1801 -2382 1801 -2382 0 net=11307
rlabel metal2 2053 -2382 2053 -2382 0 net=13347
rlabel metal2 110 -2384 110 -2384 0 net=7611
rlabel metal2 1150 -2384 1150 -2384 0 net=7103
rlabel metal2 1293 -2384 1293 -2384 0 net=10048
rlabel metal2 1899 -2384 1899 -2384 0 net=11863
rlabel metal2 324 -2386 324 -2386 0 net=1727
rlabel metal2 457 -2386 457 -2386 0 net=3955
rlabel metal2 660 -2386 660 -2386 0 net=5066
rlabel metal2 821 -2386 821 -2386 0 net=5121
rlabel metal2 884 -2386 884 -2386 0 net=3933
rlabel metal2 912 -2386 912 -2386 0 net=5485
rlabel metal2 1479 -2386 1479 -2386 0 net=10505
rlabel metal2 1752 -2386 1752 -2386 0 net=11151
rlabel metal2 1801 -2386 1801 -2386 0 net=12079
rlabel metal2 324 -2388 324 -2388 0 net=3215
rlabel metal2 464 -2388 464 -2388 0 net=2705
rlabel metal2 492 -2388 492 -2388 0 net=8015
rlabel metal2 1465 -2388 1465 -2388 0 net=9199
rlabel metal2 303 -2390 303 -2390 0 net=2015
rlabel metal2 464 -2390 464 -2390 0 net=5851
rlabel metal2 1115 -2390 1115 -2390 0 net=9973
rlabel metal2 1703 -2390 1703 -2390 0 net=10715
rlabel metal2 303 -2392 303 -2392 0 net=2147
rlabel metal2 520 -2392 520 -2392 0 net=2795
rlabel metal2 702 -2392 702 -2392 0 net=13199
rlabel metal2 1311 -2392 1311 -2392 0 net=8151
rlabel metal2 1710 -2392 1710 -2392 0 net=10563
rlabel metal2 331 -2394 331 -2394 0 net=1745
rlabel metal2 380 -2394 380 -2394 0 net=4733
rlabel metal2 527 -2394 527 -2394 0 net=10485
rlabel metal2 1339 -2394 1339 -2394 0 net=8293
rlabel metal2 1598 -2394 1598 -2394 0 net=10935
rlabel metal2 345 -2396 345 -2396 0 net=1813
rlabel metal2 380 -2396 380 -2396 0 net=3179
rlabel metal2 499 -2396 499 -2396 0 net=4355
rlabel metal2 758 -2396 758 -2396 0 net=6085
rlabel metal2 1115 -2396 1115 -2396 0 net=7119
rlabel metal2 1367 -2396 1367 -2396 0 net=8649
rlabel metal2 219 -2398 219 -2398 0 net=1793
rlabel metal2 436 -2398 436 -2398 0 net=2577
rlabel metal2 499 -2398 499 -2398 0 net=3409
rlabel metal2 576 -2398 576 -2398 0 net=4053
rlabel metal2 814 -2398 814 -2398 0 net=6745
rlabel metal2 1129 -2398 1129 -2398 0 net=8325
rlabel metal2 149 -2400 149 -2400 0 net=4717
rlabel metal2 233 -2400 233 -2400 0 net=4183
rlabel metal2 590 -2400 590 -2400 0 net=3423
rlabel metal2 621 -2400 621 -2400 0 net=13595
rlabel metal2 149 -2402 149 -2402 0 net=7013
rlabel metal2 233 -2402 233 -2402 0 net=1779
rlabel metal2 597 -2402 597 -2402 0 net=5923
rlabel metal2 1171 -2402 1171 -2402 0 net=7065
rlabel metal2 359 -2404 359 -2404 0 net=2255
rlabel metal2 611 -2404 611 -2404 0 net=3621
rlabel metal2 646 -2404 646 -2404 0 net=6313
rlabel metal2 814 -2404 814 -2404 0 net=5031
rlabel metal2 884 -2404 884 -2404 0 net=5517
rlabel metal2 198 -2406 198 -2406 0 net=1851
rlabel metal2 443 -2406 443 -2406 0 net=2557
rlabel metal2 478 -2406 478 -2406 0 net=301
rlabel metal2 919 -2406 919 -2406 0 net=14176
rlabel metal2 184 -2408 184 -2408 0 net=1901
rlabel metal2 443 -2408 443 -2408 0 net=3553
rlabel metal2 628 -2408 628 -2408 0 net=7606
rlabel metal2 828 -2408 828 -2408 0 net=5349
rlabel metal2 922 -2408 922 -2408 0 net=6319
rlabel metal2 135 -2410 135 -2410 0 net=5114
rlabel metal2 632 -2410 632 -2410 0 net=5393
rlabel metal2 737 -2410 737 -2410 0 net=9865
rlabel metal2 135 -2412 135 -2412 0 net=2169
rlabel metal2 660 -2412 660 -2412 0 net=2063
rlabel metal2 1013 -2412 1013 -2412 0 net=9029
rlabel metal2 184 -2414 184 -2414 0 net=4853
rlabel metal2 670 -2414 670 -2414 0 net=14274
rlabel metal2 268 -2416 268 -2416 0 net=8109
rlabel metal2 800 -2416 800 -2416 0 net=4953
rlabel metal2 828 -2416 828 -2416 0 net=5359
rlabel metal2 922 -2416 922 -2416 0 net=9028
rlabel metal2 2270 -2416 2270 -2416 0 net=14513
rlabel metal2 366 -2418 366 -2418 0 net=5271
rlabel metal2 835 -2418 835 -2418 0 net=5635
rlabel metal2 1017 -2418 1017 -2418 0 net=6702
rlabel metal2 1171 -2418 1171 -2418 0 net=11376
rlabel metal2 121 -2420 121 -2420 0 net=6457
rlabel metal2 1031 -2420 1031 -2420 0 net=13003
rlabel metal2 1808 -2420 1808 -2420 0 net=12105
rlabel metal2 121 -2422 121 -2422 0 net=6867
rlabel metal2 863 -2422 863 -2422 0 net=5417
rlabel metal2 957 -2422 957 -2422 0 net=6669
rlabel metal2 1174 -2422 1174 -2422 0 net=12383
rlabel metal2 1332 -2422 1332 -2422 0 net=8011
rlabel metal2 107 -2424 107 -2424 0 net=3722
rlabel metal2 898 -2424 898 -2424 0 net=5619
rlabel metal2 975 -2424 975 -2424 0 net=10051
rlabel metal2 1633 -2424 1633 -2424 0 net=10191
rlabel metal2 107 -2426 107 -2426 0 net=3282
rlabel metal2 156 -2426 156 -2426 0 net=3913
rlabel metal2 415 -2426 415 -2426 0 net=2907
rlabel metal2 555 -2426 555 -2426 0 net=4755
rlabel metal2 933 -2426 933 -2426 0 net=13779
rlabel metal2 79 -2428 79 -2428 0 net=5243
rlabel metal2 639 -2428 639 -2428 0 net=2739
rlabel metal2 936 -2428 936 -2428 0 net=183
rlabel metal2 1724 -2428 1724 -2428 0 net=10955
rlabel metal2 2 -2430 2 -2430 0 net=5767
rlabel metal2 86 -2430 86 -2430 0 net=5539
rlabel metal2 947 -2430 947 -2430 0 net=6277
rlabel metal2 1139 -2430 1139 -2430 0 net=14441
rlabel metal2 2 -2432 2 -2432 0 net=8041
rlabel metal2 86 -2432 86 -2432 0 net=3979
rlabel metal2 1507 -2432 1507 -2432 0 net=10729
rlabel metal2 1731 -2432 1731 -2432 0 net=11531
rlabel metal2 128 -2434 128 -2434 0 net=4051
rlabel metal2 695 -2434 695 -2434 0 net=4695
rlabel metal2 961 -2434 961 -2434 0 net=6709
rlabel metal2 1178 -2434 1178 -2434 0 net=8051
rlabel metal2 1346 -2434 1346 -2434 0 net=11951
rlabel metal2 96 -2436 96 -2436 0 net=13349
rlabel metal2 1192 -2436 1192 -2436 0 net=9429
rlabel metal2 1346 -2436 1346 -2436 0 net=8443
rlabel metal2 1500 -2436 1500 -2436 0 net=9829
rlabel metal2 1605 -2436 1605 -2436 0 net=9561
rlabel metal2 58 -2438 58 -2438 0 net=5544
rlabel metal2 156 -2438 156 -2438 0 net=1595
rlabel metal2 513 -2438 513 -2438 0 net=4665
rlabel metal2 688 -2438 688 -2438 0 net=4739
rlabel metal2 968 -2438 968 -2438 0 net=5707
rlabel metal2 1066 -2438 1066 -2438 0 net=6521
rlabel metal2 1213 -2438 1213 -2438 0 net=10581
rlabel metal2 58 -2440 58 -2440 0 net=11542
rlabel metal2 1010 -2440 1010 -2440 0 net=6378
rlabel metal2 1122 -2440 1122 -2440 0 net=7325
rlabel metal2 1325 -2440 1325 -2440 0 net=8267
rlabel metal2 1507 -2440 1507 -2440 0 net=10389
rlabel metal2 1584 -2440 1584 -2440 0 net=10249
rlabel metal2 142 -2442 142 -2442 0 net=10243
rlabel metal2 793 -2442 793 -2442 0 net=6783
rlabel metal2 1143 -2442 1143 -2442 0 net=9525
rlabel metal2 1556 -2442 1556 -2442 0 net=10159
rlabel metal2 93 -2444 93 -2444 0 net=8335
rlabel metal2 205 -2444 205 -2444 0 net=4279
rlabel metal2 975 -2444 975 -2444 0 net=12881
rlabel metal2 93 -2446 93 -2446 0 net=11765
rlabel metal2 205 -2448 205 -2448 0 net=4505
rlabel metal2 996 -2448 996 -2448 0 net=5969
rlabel metal2 1206 -2448 1206 -2448 0 net=7669
rlabel metal2 1353 -2448 1353 -2448 0 net=8623
rlabel metal2 1458 -2448 1458 -2448 0 net=9989
rlabel metal2 212 -2450 212 -2450 0 net=1583
rlabel metal2 548 -2450 548 -2450 0 net=3001
rlabel metal2 289 -2452 289 -2452 0 net=1571
rlabel metal2 674 -2452 674 -2452 0 net=1535
rlabel metal2 1045 -2452 1045 -2452 0 net=6561
rlabel metal2 1234 -2452 1234 -2452 0 net=7953
rlabel metal2 338 -2454 338 -2454 0 net=2917
rlabel metal2 926 -2454 926 -2454 0 net=5265
rlabel metal2 1353 -2454 1353 -2454 0 net=13478
rlabel metal2 541 -2456 541 -2456 0 net=7423
rlabel metal2 992 -2456 992 -2456 0 net=13221
rlabel metal2 772 -2458 772 -2458 0 net=3471
rlabel metal2 1199 -2458 1199 -2458 0 net=13711
rlabel metal2 23 -2460 23 -2460 0 net=4297
rlabel metal2 849 -2460 849 -2460 0 net=5221
rlabel metal2 1367 -2460 1367 -2460 0 net=8529
rlabel metal2 1458 -2460 1458 -2460 0 net=11187
rlabel metal2 1199 -2462 1199 -2462 0 net=7439
rlabel metal2 1430 -2462 1430 -2462 0 net=10209
rlabel metal2 1283 -2464 1283 -2464 0 net=8411
rlabel metal2 1521 -2464 1521 -2464 0 net=10263
rlabel metal2 373 -2466 373 -2466 0 net=2835
rlabel metal2 373 -2468 373 -2468 0 net=3261
rlabel metal2 1416 -2468 1416 -2468 0 net=9123
rlabel metal2 1563 -2468 1563 -2468 0 net=9655
rlabel metal2 583 -2470 583 -2470 0 net=3689
rlabel metal2 1472 -2470 1472 -2470 0 net=10373
rlabel metal2 1640 -2470 1640 -2470 0 net=11335
rlabel metal2 653 -2472 653 -2472 0 net=4001
rlabel metal2 1563 -2472 1563 -2472 0 net=10367
rlabel metal2 1815 -2472 1815 -2472 0 net=11713
rlabel metal2 751 -2474 751 -2474 0 net=6337
rlabel metal2 1689 -2474 1689 -2474 0 net=10893
rlabel metal2 1871 -2474 1871 -2474 0 net=11971
rlabel metal2 1073 -2476 1073 -2476 0 net=11234
rlabel metal2 1759 -2478 1759 -2478 0 net=11273
rlabel metal2 1920 -2478 1920 -2478 0 net=12181
rlabel metal2 1675 -2480 1675 -2480 0 net=10337
rlabel metal2 1955 -2480 1955 -2480 0 net=12405
rlabel metal2 1962 -2482 1962 -2482 0 net=12533
rlabel metal2 1083 -2484 1083 -2484 0 net=12969
rlabel metal2 2004 -2486 2004 -2486 0 net=12685
rlabel metal2 2032 -2488 2032 -2488 0 net=13123
rlabel metal2 1220 -2490 1220 -2490 0 net=7359
rlabel metal2 1220 -2492 1220 -2492 0 net=7709
rlabel metal2 1241 -2494 1241 -2494 0 net=7535
rlabel metal2 1269 -2496 1269 -2496 0 net=10229
rlabel metal2 5 -2507 5 -2507 0 net=2908
rlabel metal2 464 -2507 464 -2507 0 net=5852
rlabel metal2 992 -2507 992 -2507 0 net=1292
rlabel metal2 1080 -2507 1080 -2507 0 net=10338
rlabel metal2 1801 -2507 1801 -2507 0 net=12377
rlabel metal2 2088 -2507 2088 -2507 0 net=14551
rlabel metal2 9 -2509 9 -2509 0 net=7966
rlabel metal2 1510 -2509 1510 -2509 0 net=13348
rlabel metal2 2088 -2509 2088 -2509 0 net=13781
rlabel metal2 9 -2511 9 -2511 0 net=9799
rlabel metal2 54 -2511 54 -2511 0 net=4224
rlabel metal2 775 -2511 775 -2511 0 net=5350
rlabel metal2 926 -2511 926 -2511 0 net=3472
rlabel metal2 1188 -2511 1188 -2511 0 net=10694
rlabel metal2 1717 -2511 1717 -2511 0 net=10565
rlabel metal2 1717 -2511 1717 -2511 0 net=10565
rlabel metal2 1794 -2511 1794 -2511 0 net=12065
rlabel metal2 1934 -2511 1934 -2511 0 net=12971
rlabel metal2 2053 -2511 2053 -2511 0 net=13597
rlabel metal2 16 -2513 16 -2513 0 net=2767
rlabel metal2 40 -2513 40 -2513 0 net=7854
rlabel metal2 1290 -2513 1290 -2513 0 net=10192
rlabel metal2 1885 -2513 1885 -2513 0 net=12841
rlabel metal2 2025 -2513 2025 -2513 0 net=13553
rlabel metal2 2130 -2513 2130 -2513 0 net=14091
rlabel metal2 33 -2515 33 -2515 0 net=5540
rlabel metal2 950 -2515 950 -2515 0 net=8807
rlabel metal2 1335 -2515 1335 -2515 0 net=12210
rlabel metal2 37 -2517 37 -2517 0 net=9695
rlabel metal2 58 -2517 58 -2517 0 net=7066
rlabel metal2 1521 -2517 1521 -2517 0 net=10265
rlabel metal2 1521 -2517 1521 -2517 0 net=10265
rlabel metal2 1580 -2517 1580 -2517 0 net=9320
rlabel metal2 1678 -2517 1678 -2517 0 net=11308
rlabel metal2 1997 -2517 1997 -2517 0 net=13399
rlabel metal2 2102 -2517 2102 -2517 0 net=14425
rlabel metal2 44 -2519 44 -2519 0 net=5632
rlabel metal2 93 -2519 93 -2519 0 net=7104
rlabel metal2 1195 -2519 1195 -2519 0 net=12022
rlabel metal2 1969 -2519 1969 -2519 0 net=13125
rlabel metal2 2109 -2519 2109 -2519 0 net=13997
rlabel metal2 2242 -2519 2242 -2519 0 net=14751
rlabel metal2 44 -2521 44 -2521 0 net=10487
rlabel metal2 541 -2521 541 -2521 0 net=7424
rlabel metal2 989 -2521 989 -2521 0 net=9983
rlabel metal2 1199 -2521 1199 -2521 0 net=7440
rlabel metal2 1356 -2521 1356 -2521 0 net=11349
rlabel metal2 1804 -2521 1804 -2521 0 net=13812
rlabel metal2 58 -2523 58 -2523 0 net=1941
rlabel metal2 72 -2523 72 -2523 0 net=8042
rlabel metal2 1332 -2523 1332 -2523 0 net=9125
rlabel metal2 1458 -2523 1458 -2523 0 net=11189
rlabel metal2 2172 -2523 2172 -2523 0 net=14413
rlabel metal2 72 -2525 72 -2525 0 net=3914
rlabel metal2 373 -2525 373 -2525 0 net=3262
rlabel metal2 817 -2525 817 -2525 0 net=13889
rlabel metal2 2186 -2525 2186 -2525 0 net=14557
rlabel metal2 93 -2527 93 -2527 0 net=2211
rlabel metal2 128 -2527 128 -2527 0 net=4052
rlabel metal2 859 -2527 859 -2527 0 net=11159
rlabel metal2 1808 -2527 1808 -2527 0 net=11973
rlabel metal2 2235 -2527 2235 -2527 0 net=14701
rlabel metal2 107 -2529 107 -2529 0 net=2441
rlabel metal2 268 -2529 268 -2529 0 net=8111
rlabel metal2 877 -2529 877 -2529 0 net=8153
rlabel metal2 1360 -2529 1360 -2529 0 net=12488
rlabel metal2 110 -2531 110 -2531 0 net=10681
rlabel metal2 1374 -2531 1374 -2531 0 net=11464
rlabel metal2 2116 -2531 2116 -2531 0 net=13589
rlabel metal2 131 -2533 131 -2533 0 net=5708
rlabel metal2 1006 -2533 1006 -2533 0 net=13004
rlabel metal2 1038 -2533 1038 -2533 0 net=9079
rlabel metal2 1216 -2533 1216 -2533 0 net=14514
rlabel metal2 19 -2535 19 -2535 0 net=8877
rlabel metal2 1038 -2535 1038 -2535 0 net=6670
rlabel metal2 1311 -2535 1311 -2535 0 net=11484
rlabel metal2 1871 -2535 1871 -2535 0 net=12323
rlabel metal2 1941 -2535 1941 -2535 0 net=13833
rlabel metal2 2270 -2535 2270 -2535 0 net=6321
rlabel metal2 149 -2537 149 -2537 0 net=7015
rlabel metal2 275 -2537 275 -2537 0 net=1934
rlabel metal2 898 -2537 898 -2537 0 net=5621
rlabel metal2 940 -2537 940 -2537 0 net=8251
rlabel metal2 1377 -2537 1377 -2537 0 net=9656
rlabel metal2 1843 -2537 1843 -2537 0 net=12081
rlabel metal2 2123 -2537 2123 -2537 0 net=14009
rlabel metal2 103 -2539 103 -2539 0 net=5901
rlabel metal2 919 -2539 919 -2539 0 net=9513
rlabel metal2 1010 -2539 1010 -2539 0 net=7326
rlabel metal2 1402 -2539 1402 -2539 0 net=9031
rlabel metal2 1416 -2539 1416 -2539 0 net=9293
rlabel metal2 1458 -2539 1458 -2539 0 net=9867
rlabel metal2 1580 -2539 1580 -2539 0 net=12686
rlabel metal2 2165 -2539 2165 -2539 0 net=14389
rlabel metal2 128 -2541 128 -2541 0 net=6403
rlabel metal2 1013 -2541 1013 -2541 0 net=9303
rlabel metal2 1402 -2541 1402 -2541 0 net=8925
rlabel metal2 1465 -2541 1465 -2541 0 net=10003
rlabel metal2 1601 -2541 1601 -2541 0 net=11864
rlabel metal2 2179 -2541 2179 -2541 0 net=14443
rlabel metal2 149 -2543 149 -2543 0 net=1877
rlabel metal2 478 -2543 478 -2543 0 net=2836
rlabel metal2 1766 -2543 1766 -2543 0 net=11403
rlabel metal2 163 -2545 163 -2545 0 net=2058
rlabel metal2 191 -2545 191 -2545 0 net=2307
rlabel metal2 303 -2545 303 -2545 0 net=2148
rlabel metal2 429 -2545 429 -2545 0 net=4615
rlabel metal2 1444 -2545 1444 -2545 0 net=9990
rlabel metal2 1647 -2545 1647 -2545 0 net=10937
rlabel metal2 1899 -2545 1899 -2545 0 net=12535
rlabel metal2 163 -2547 163 -2547 0 net=3339
rlabel metal2 1437 -2547 1437 -2547 0 net=10716
rlabel metal2 1710 -2547 1710 -2547 0 net=12183
rlabel metal2 96 -2549 96 -2549 0 net=9201
rlabel metal2 1500 -2549 1500 -2549 0 net=9831
rlabel metal2 1542 -2549 1542 -2549 0 net=10369
rlabel metal2 1612 -2549 1612 -2549 0 net=10315
rlabel metal2 177 -2551 177 -2551 0 net=3691
rlabel metal2 604 -2551 604 -2551 0 net=3935
rlabel metal2 894 -2551 894 -2551 0 net=11725
rlabel metal2 1920 -2551 1920 -2551 0 net=12863
rlabel metal2 191 -2553 191 -2553 0 net=7447
rlabel metal2 1619 -2553 1619 -2553 0 net=12741
rlabel metal2 201 -2555 201 -2555 0 net=1399
rlabel metal2 632 -2555 632 -2555 0 net=5394
rlabel metal2 1272 -2555 1272 -2555 0 net=14619
rlabel metal2 1948 -2555 1948 -2555 0 net=13423
rlabel metal2 205 -2557 205 -2557 0 net=4507
rlabel metal2 310 -2557 310 -2557 0 net=1606
rlabel metal2 1314 -2557 1314 -2557 0 net=13913
rlabel metal2 198 -2559 198 -2559 0 net=1903
rlabel metal2 240 -2559 240 -2559 0 net=7807
rlabel metal2 555 -2559 555 -2559 0 net=5244
rlabel metal2 751 -2559 751 -2559 0 net=6339
rlabel metal2 926 -2559 926 -2559 0 net=12385
rlabel metal2 1451 -2559 1451 -2559 0 net=9629
rlabel metal2 1654 -2559 1654 -2559 0 net=11021
rlabel metal2 1948 -2559 1948 -2559 0 net=13135
rlabel metal2 198 -2561 198 -2561 0 net=3622
rlabel metal2 709 -2561 709 -2561 0 net=5272
rlabel metal2 1066 -2561 1066 -2561 0 net=6522
rlabel metal2 1451 -2561 1451 -2561 0 net=10231
rlabel metal2 1661 -2561 1661 -2561 0 net=11051
rlabel metal2 1976 -2561 1976 -2561 0 net=13223
rlabel metal2 240 -2563 240 -2563 0 net=10431
rlabel metal2 457 -2563 457 -2563 0 net=3957
rlabel metal2 709 -2563 709 -2563 0 net=4659
rlabel metal2 737 -2563 737 -2563 0 net=13495
rlabel metal2 2046 -2563 2046 -2563 0 net=14129
rlabel metal2 254 -2565 254 -2565 0 net=2129
rlabel metal2 310 -2565 310 -2565 0 net=1729
rlabel metal2 457 -2565 457 -2565 0 net=1949
rlabel metal2 562 -2565 562 -2565 0 net=10245
rlabel metal2 873 -2565 873 -2565 0 net=13535
rlabel metal2 135 -2567 135 -2567 0 net=2171
rlabel metal2 352 -2567 352 -2567 0 net=1814
rlabel metal2 1017 -2567 1017 -2567 0 net=14607
rlabel metal2 135 -2569 135 -2569 0 net=2595
rlabel metal2 352 -2569 352 -2569 0 net=2257
rlabel metal2 492 -2569 492 -2569 0 net=8017
rlabel metal2 1185 -2569 1185 -2569 0 net=13201
rlabel metal2 184 -2571 184 -2571 0 net=4855
rlabel metal2 562 -2571 562 -2571 0 net=5419
rlabel metal2 1017 -2571 1017 -2571 0 net=6849
rlabel metal2 1122 -2571 1122 -2571 0 net=8624
rlabel metal2 1479 -2571 1479 -2571 0 net=10507
rlabel metal2 1570 -2571 1570 -2571 0 net=10583
rlabel metal2 1738 -2571 1738 -2571 0 net=11431
rlabel metal2 142 -2573 142 -2573 0 net=8337
rlabel metal2 1024 -2573 1024 -2573 0 net=5555
rlabel metal2 1024 -2573 1024 -2573 0 net=5555
rlabel metal2 1052 -2573 1052 -2573 0 net=7121
rlabel metal2 1213 -2573 1213 -2573 0 net=8269
rlabel metal2 1423 -2573 1423 -2573 0 net=9881
rlabel metal2 1605 -2573 1605 -2573 0 net=10793
rlabel metal2 1787 -2573 1787 -2573 0 net=11953
rlabel metal2 142 -2575 142 -2575 0 net=6183
rlabel metal2 1066 -2575 1066 -2575 0 net=8215
rlabel metal2 1479 -2575 1479 -2575 0 net=9781
rlabel metal2 1500 -2575 1500 -2575 0 net=10251
rlabel metal2 1682 -2575 1682 -2575 0 net=11275
rlabel metal2 1850 -2575 1850 -2575 0 net=11847
rlabel metal2 184 -2577 184 -2577 0 net=3305
rlabel metal2 1073 -2577 1073 -2577 0 net=5267
rlabel metal2 1269 -2577 1269 -2577 0 net=8651
rlabel metal2 1486 -2577 1486 -2577 0 net=10053
rlabel metal2 1584 -2577 1584 -2577 0 net=9563
rlabel metal2 1731 -2577 1731 -2577 0 net=11533
rlabel metal2 1850 -2577 1850 -2577 0 net=12407
rlabel metal2 219 -2579 219 -2579 0 net=4719
rlabel metal2 450 -2579 450 -2579 0 net=5361
rlabel metal2 842 -2579 842 -2579 0 net=5195
rlabel metal2 1080 -2579 1080 -2579 0 net=7297
rlabel metal2 1094 -2579 1094 -2579 0 net=9527
rlabel metal2 1297 -2579 1297 -2579 0 net=8849
rlabel metal2 1528 -2579 1528 -2579 0 net=10731
rlabel metal2 1955 -2579 1955 -2579 0 net=12883
rlabel metal2 86 -2581 86 -2581 0 net=3981
rlabel metal2 1087 -2581 1087 -2581 0 net=8575
rlabel metal2 1388 -2581 1388 -2581 0 net=9747
rlabel metal2 1549 -2581 1549 -2581 0 net=11087
rlabel metal2 1990 -2581 1990 -2581 0 net=13457
rlabel metal2 86 -2583 86 -2583 0 net=7487
rlabel metal2 1143 -2583 1143 -2583 0 net=7711
rlabel metal2 1234 -2583 1234 -2583 0 net=7955
rlabel metal2 1395 -2583 1395 -2583 0 net=10838
rlabel metal2 1878 -2583 1878 -2583 0 net=13361
rlabel metal2 26 -2585 26 -2585 0 net=12461
rlabel metal2 219 -2587 219 -2587 0 net=1639
rlabel metal2 359 -2587 359 -2587 0 net=1852
rlabel metal2 1430 -2587 1430 -2587 0 net=10211
rlabel metal2 1591 -2587 1591 -2587 0 net=11381
rlabel metal2 1745 -2587 1745 -2587 0 net=11715
rlabel metal2 1829 -2587 1829 -2587 0 net=12261
rlabel metal2 212 -2589 212 -2589 0 net=1585
rlabel metal2 331 -2589 331 -2589 0 net=1747
rlabel metal2 366 -2589 366 -2589 0 net=2675
rlabel metal2 569 -2589 569 -2589 0 net=4315
rlabel metal2 646 -2589 646 -2589 0 net=6314
rlabel metal2 1220 -2589 1220 -2589 0 net=8295
rlabel metal2 1430 -2589 1430 -2589 0 net=534
rlabel metal2 1626 -2589 1626 -2589 0 net=10895
rlabel metal2 1815 -2589 1815 -2589 0 net=11943
rlabel metal2 212 -2591 212 -2591 0 net=5925
rlabel metal2 646 -2591 646 -2591 0 net=4281
rlabel metal2 716 -2591 716 -2591 0 net=5737
rlabel metal2 828 -2591 828 -2591 0 net=8099
rlabel metal2 1318 -2591 1318 -2591 0 net=9975
rlabel metal2 1591 -2591 1591 -2591 0 net=11185
rlabel metal2 1836 -2591 1836 -2591 0 net=12077
rlabel metal2 68 -2593 68 -2593 0 net=12449
rlabel metal2 716 -2593 716 -2593 0 net=7671
rlabel metal2 1234 -2593 1234 -2593 0 net=7952
rlabel metal2 1339 -2593 1339 -2593 0 net=7905
rlabel metal2 1472 -2593 1472 -2593 0 net=10375
rlabel metal2 1598 -2593 1598 -2593 0 net=10779
rlabel metal2 1773 -2593 1773 -2593 0 net=11767
rlabel metal2 1857 -2593 1857 -2593 0 net=13539
rlabel metal2 226 -2595 226 -2595 0 net=4683
rlabel metal2 282 -2595 282 -2595 0 net=3289
rlabel metal2 1171 -2595 1171 -2595 0 net=4713
rlabel metal2 2074 -2595 2074 -2595 0 net=13713
rlabel metal2 170 -2597 170 -2597 0 net=2109
rlabel metal2 282 -2597 282 -2597 0 net=13149
rlabel metal2 723 -2597 723 -2597 0 net=4391
rlabel metal2 751 -2597 751 -2597 0 net=2991
rlabel metal2 1171 -2597 1171 -2597 0 net=8053
rlabel metal2 1262 -2597 1262 -2597 0 net=8445
rlabel metal2 1412 -2597 1412 -2597 0 net=9885
rlabel metal2 1633 -2597 1633 -2597 0 net=10939
rlabel metal2 166 -2599 166 -2599 0 net=8303
rlabel metal2 331 -2599 331 -2599 0 net=1795
rlabel metal2 373 -2599 373 -2599 0 net=2017
rlabel metal2 401 -2599 401 -2599 0 net=4030
rlabel metal2 954 -2599 954 -2599 0 net=9149
rlabel metal2 1640 -2599 1640 -2599 0 net=11337
rlabel metal2 1822 -2599 1822 -2599 0 net=12107
rlabel metal2 2144 -2599 2144 -2599 0 net=14255
rlabel metal2 30 -2601 30 -2601 0 net=1891
rlabel metal2 380 -2601 380 -2601 0 net=3181
rlabel metal2 569 -2601 569 -2601 0 net=5033
rlabel metal2 824 -2601 824 -2601 0 net=9051
rlabel metal2 1640 -2601 1640 -2601 0 net=10957
rlabel metal2 1913 -2601 1913 -2601 0 net=12781
rlabel metal2 2214 -2601 2214 -2601 0 net=14681
rlabel metal2 30 -2603 30 -2603 0 net=2707
rlabel metal2 506 -2603 506 -2603 0 net=5223
rlabel metal2 1178 -2603 1178 -2603 0 net=13351
rlabel metal2 2263 -2603 2263 -2603 0 net=4535
rlabel metal2 79 -2605 79 -2605 0 net=5769
rlabel metal2 1003 -2605 1003 -2605 0 net=6459
rlabel metal2 1206 -2605 1206 -2605 0 net=8413
rlabel metal2 1447 -2605 1447 -2605 0 net=11361
rlabel metal2 79 -2607 79 -2607 0 net=3003
rlabel metal2 583 -2607 583 -2607 0 net=4955
rlabel metal2 807 -2607 807 -2607 0 net=4756
rlabel metal2 1255 -2607 1255 -2607 0 net=5745
rlabel metal2 1668 -2607 1668 -2607 0 net=11153
rlabel metal2 156 -2609 156 -2609 0 net=1597
rlabel metal2 408 -2609 408 -2609 0 net=2621
rlabel metal2 485 -2609 485 -2609 0 net=2741
rlabel metal2 726 -2609 726 -2609 0 net=7360
rlabel metal2 156 -2611 156 -2611 0 net=5109
rlabel metal2 597 -2611 597 -2611 0 net=3775
rlabel metal2 1752 -2611 1752 -2611 0 net=8012
rlabel metal2 289 -2613 289 -2613 0 net=1572
rlabel metal2 520 -2613 520 -2613 0 net=4734
rlabel metal2 2081 -2613 2081 -2613 0 net=13731
rlabel metal2 65 -2615 65 -2615 0 net=1527
rlabel metal2 380 -2615 380 -2615 0 net=2065
rlabel metal2 730 -2615 730 -2615 0 net=2201
rlabel metal2 2151 -2615 2151 -2615 0 net=14341
rlabel metal2 65 -2617 65 -2617 0 net=7404
rlabel metal2 387 -2619 387 -2619 0 net=6533
rlabel metal2 513 -2619 513 -2619 0 net=4667
rlabel metal2 758 -2619 758 -2619 0 net=6087
rlabel metal2 2067 -2619 2067 -2619 0 net=13671
rlabel metal2 338 -2621 338 -2621 0 net=2919
rlabel metal2 394 -2621 394 -2621 0 net=6017
rlabel metal2 2137 -2621 2137 -2621 0 net=14109
rlabel metal2 338 -2623 338 -2623 0 net=3411
rlabel metal2 513 -2623 513 -2623 0 net=4741
rlabel metal2 786 -2623 786 -2623 0 net=7011
rlabel metal2 443 -2625 443 -2625 0 net=3555
rlabel metal2 520 -2625 520 -2625 0 net=4055
rlabel metal2 590 -2625 590 -2625 0 net=3425
rlabel metal2 800 -2625 800 -2625 0 net=10161
rlabel metal2 233 -2627 233 -2627 0 net=1781
rlabel metal2 534 -2627 534 -2627 0 net=4185
rlabel metal2 618 -2627 618 -2627 0 net=4134
rlabel metal2 849 -2627 849 -2627 0 net=6785
rlabel metal2 1507 -2627 1507 -2627 0 net=10391
rlabel metal2 233 -2629 233 -2629 0 net=1537
rlabel metal2 695 -2629 695 -2629 0 net=5971
rlabel metal2 1101 -2629 1101 -2629 0 net=7613
rlabel metal2 1248 -2629 1248 -2629 0 net=7541
rlabel metal2 324 -2631 324 -2631 0 net=3217
rlabel metal2 548 -2631 548 -2631 0 net=5637
rlabel metal2 982 -2631 982 -2631 0 net=6747
rlabel metal2 1136 -2631 1136 -2631 0 net=9537
rlabel metal2 324 -2633 324 -2633 0 net=2559
rlabel metal2 576 -2633 576 -2633 0 net=3447
rlabel metal2 796 -2633 796 -2633 0 net=7469
rlabel metal2 23 -2635 23 -2635 0 net=4299
rlabel metal2 618 -2635 618 -2635 0 net=5519
rlabel metal2 996 -2635 996 -2635 0 net=6563
rlabel metal2 639 -2637 639 -2637 0 net=2797
rlabel metal2 779 -2637 779 -2637 0 net=4549
rlabel metal2 884 -2637 884 -2637 0 net=5513
rlabel metal2 1045 -2637 1045 -2637 0 net=8789
rlabel metal2 121 -2639 121 -2639 0 net=6869
rlabel metal2 1241 -2639 1241 -2639 0 net=7537
rlabel metal2 481 -2641 481 -2641 0 net=6021
rlabel metal2 1241 -2641 1241 -2641 0 net=9200
rlabel metal2 625 -2643 625 -2643 0 net=6231
rlabel metal2 1013 -2643 1013 -2643 0 net=11805
rlabel metal2 625 -2645 625 -2645 0 net=5487
rlabel metal2 667 -2647 667 -2647 0 net=14609
rlabel metal2 667 -2649 667 -2649 0 net=4357
rlabel metal2 912 -2649 912 -2649 0 net=8327
rlabel metal2 674 -2651 674 -2651 0 net=5123
rlabel metal2 1129 -2651 1129 -2651 0 net=7899
rlabel metal2 114 -2653 114 -2653 0 net=7133
rlabel metal2 1164 -2653 1164 -2653 0 net=7797
rlabel metal2 702 -2655 702 -2655 0 net=4697
rlabel metal2 1227 -2655 1227 -2655 0 net=8531
rlabel metal2 744 -2657 744 -2657 0 net=6711
rlabel metal2 1192 -2657 1192 -2657 0 net=9431
rlabel metal2 947 -2659 947 -2659 0 net=6279
rlabel metal2 1192 -2659 1192 -2659 0 net=12705
rlabel metal2 296 -2661 296 -2661 0 net=6062
rlabel metal2 296 -2663 296 -2663 0 net=2579
rlabel metal2 436 -2665 436 -2665 0 net=4003
rlabel metal2 100 -2667 100 -2667 0 net=5457
rlabel metal2 100 -2669 100 -2669 0 net=5693
rlabel metal2 2 -2680 2 -2680 0 net=8391
rlabel metal2 103 -2680 103 -2680 0 net=3412
rlabel metal2 373 -2680 373 -2680 0 net=2019
rlabel metal2 373 -2680 373 -2680 0 net=2019
rlabel metal2 432 -2680 432 -2680 0 net=2622
rlabel metal2 506 -2680 506 -2680 0 net=5224
rlabel metal2 758 -2680 758 -2680 0 net=3426
rlabel metal2 915 -2680 915 -2680 0 net=14130
rlabel metal2 2200 -2680 2200 -2680 0 net=14611
rlabel metal2 2200 -2680 2200 -2680 0 net=14611
rlabel metal2 2224 -2680 2224 -2680 0 net=6322
rlabel metal2 16 -2682 16 -2682 0 net=2768
rlabel metal2 338 -2682 338 -2682 0 net=1893
rlabel metal2 506 -2682 506 -2682 0 net=6871
rlabel metal2 786 -2682 786 -2682 0 net=9080
rlabel metal2 1185 -2682 1185 -2682 0 net=12842
rlabel metal2 1927 -2682 1927 -2682 0 net=10316
rlabel metal2 16 -2684 16 -2684 0 net=5973
rlabel metal2 709 -2684 709 -2684 0 net=4660
rlabel metal2 978 -2684 978 -2684 0 net=7012
rlabel metal2 1286 -2684 1286 -2684 0 net=9868
rlabel metal2 1489 -2684 1489 -2684 0 net=11186
rlabel metal2 1605 -2684 1605 -2684 0 net=10795
rlabel metal2 1605 -2684 1605 -2684 0 net=10795
rlabel metal2 1619 -2684 1619 -2684 0 net=12743
rlabel metal2 1934 -2684 1934 -2684 0 net=12973
rlabel metal2 1934 -2684 1934 -2684 0 net=12973
rlabel metal2 1948 -2684 1948 -2684 0 net=13137
rlabel metal2 1948 -2684 1948 -2684 0 net=13137
rlabel metal2 2235 -2684 2235 -2684 0 net=14703
rlabel metal2 2235 -2684 2235 -2684 0 net=14703
rlabel metal2 2242 -2684 2242 -2684 0 net=14753
rlabel metal2 2242 -2684 2242 -2684 0 net=14753
rlabel metal2 23 -2686 23 -2686 0 net=2596
rlabel metal2 156 -2686 156 -2686 0 net=5110
rlabel metal2 1062 -2686 1062 -2686 0 net=11585
rlabel metal2 1139 -2686 1139 -2686 0 net=9782
rlabel metal2 1577 -2686 1577 -2686 0 net=7513
rlabel metal2 23 -2688 23 -2688 0 net=4057
rlabel metal2 548 -2688 548 -2688 0 net=5638
rlabel metal2 821 -2688 821 -2688 0 net=5622
rlabel metal2 954 -2688 954 -2688 0 net=7712
rlabel metal2 1185 -2688 1185 -2688 0 net=8415
rlabel metal2 1234 -2688 1234 -2688 0 net=13496
rlabel metal2 26 -2690 26 -2690 0 net=3982
rlabel metal2 919 -2690 919 -2690 0 net=12884
rlabel metal2 58 -2692 58 -2692 0 net=1943
rlabel metal2 58 -2692 58 -2692 0 net=1943
rlabel metal2 65 -2692 65 -2692 0 net=7488
rlabel metal2 110 -2692 110 -2692 0 net=13150
rlabel metal2 345 -2692 345 -2692 0 net=1749
rlabel metal2 387 -2692 387 -2692 0 net=2921
rlabel metal2 555 -2692 555 -2692 0 net=4316
rlabel metal2 653 -2692 653 -2692 0 net=5459
rlabel metal2 653 -2692 653 -2692 0 net=5459
rlabel metal2 681 -2692 681 -2692 0 net=6233
rlabel metal2 765 -2692 765 -2692 0 net=10246
rlabel metal2 954 -2692 954 -2692 0 net=5197
rlabel metal2 1013 -2692 1013 -2692 0 net=14426
rlabel metal2 65 -2694 65 -2694 0 net=6565
rlabel metal2 1041 -2694 1041 -2694 0 net=12324
rlabel metal2 1955 -2694 1955 -2694 0 net=13225
rlabel metal2 2102 -2694 2102 -2694 0 net=14111
rlabel metal2 82 -2696 82 -2696 0 net=4147
rlabel metal2 681 -2696 681 -2696 0 net=7673
rlabel metal2 765 -2696 765 -2696 0 net=8297
rlabel metal2 1234 -2696 1234 -2696 0 net=9365
rlabel metal2 1423 -2696 1423 -2696 0 net=9883
rlabel metal2 1479 -2696 1479 -2696 0 net=10393
rlabel metal2 1584 -2696 1584 -2696 0 net=9564
rlabel metal2 1755 -2696 1755 -2696 0 net=14552
rlabel metal2 86 -2698 86 -2698 0 net=9991
rlabel metal2 1318 -2698 1318 -2698 0 net=9977
rlabel metal2 107 -2700 107 -2700 0 net=2443
rlabel metal2 558 -2700 558 -2700 0 net=4668
rlabel metal2 695 -2700 695 -2700 0 net=4393
rlabel metal2 772 -2700 772 -2700 0 net=6341
rlabel metal2 919 -2700 919 -2700 0 net=6281
rlabel metal2 975 -2700 975 -2700 0 net=12929
rlabel metal2 1976 -2700 1976 -2700 0 net=13459
rlabel metal2 2130 -2700 2130 -2700 0 net=14093
rlabel metal2 2158 -2700 2158 -2700 0 net=14415
rlabel metal2 121 -2702 121 -2702 0 net=5694
rlabel metal2 163 -2702 163 -2702 0 net=3341
rlabel metal2 562 -2702 562 -2702 0 net=5420
rlabel metal2 1066 -2702 1066 -2702 0 net=8217
rlabel metal2 1195 -2702 1195 -2702 0 net=1037
rlabel metal2 1556 -2702 1556 -2702 0 net=11955
rlabel metal2 1871 -2702 1871 -2702 0 net=12707
rlabel metal2 2011 -2702 2011 -2702 0 net=13425
rlabel metal2 2130 -2702 2130 -2702 0 net=14257
rlabel metal2 51 -2704 51 -2704 0 net=11029
rlabel metal2 1584 -2704 1584 -2704 0 net=11351
rlabel metal2 1759 -2704 1759 -2704 0 net=11535
rlabel metal2 2144 -2704 2144 -2704 0 net=14343
rlabel metal2 51 -2706 51 -2706 0 net=6748
rlabel metal2 996 -2706 996 -2706 0 net=8271
rlabel metal2 1220 -2706 1220 -2706 0 net=8447
rlabel metal2 1360 -2706 1360 -2706 0 net=10683
rlabel metal2 1619 -2706 1619 -2706 0 net=10941
rlabel metal2 1647 -2706 1647 -2706 0 net=10938
rlabel metal2 1759 -2706 1759 -2706 0 net=11727
rlabel metal2 1773 -2706 1773 -2706 0 net=11769
rlabel metal2 1773 -2706 1773 -2706 0 net=11769
rlabel metal2 1899 -2706 1899 -2706 0 net=12537
rlabel metal2 2151 -2706 2151 -2706 0 net=14391
rlabel metal2 121 -2708 121 -2708 0 net=4359
rlabel metal2 730 -2708 730 -2708 0 net=2203
rlabel metal2 1066 -2708 1066 -2708 0 net=7901
rlabel metal2 1206 -2708 1206 -2708 0 net=8533
rlabel metal2 1241 -2708 1241 -2708 0 net=4714
rlabel metal2 1899 -2708 1899 -2708 0 net=12783
rlabel metal2 2165 -2708 2165 -2708 0 net=14445
rlabel metal2 128 -2710 128 -2710 0 net=4005
rlabel metal2 457 -2710 457 -2710 0 net=1951
rlabel metal2 576 -2710 576 -2710 0 net=3449
rlabel metal2 730 -2710 730 -2710 0 net=14577
rlabel metal2 93 -2712 93 -2712 0 net=2213
rlabel metal2 513 -2712 513 -2712 0 net=4743
rlabel metal2 772 -2712 772 -2712 0 net=8055
rlabel metal2 1213 -2712 1213 -2712 0 net=8653
rlabel metal2 1276 -2712 1276 -2712 0 net=7539
rlabel metal2 1374 -2712 1374 -2712 0 net=9304
rlabel metal2 1598 -2712 1598 -2712 0 net=10781
rlabel metal2 1647 -2712 1647 -2712 0 net=11023
rlabel metal2 1668 -2712 1668 -2712 0 net=11155
rlabel metal2 1766 -2712 1766 -2712 0 net=13599
rlabel metal2 93 -2714 93 -2714 0 net=7135
rlabel metal2 163 -2714 163 -2714 0 net=2259
rlabel metal2 366 -2714 366 -2714 0 net=2676
rlabel metal2 663 -2714 663 -2714 0 net=8999
rlabel metal2 1388 -2714 1388 -2714 0 net=9749
rlabel metal2 1430 -2714 1430 -2714 0 net=13352
rlabel metal2 2053 -2714 2053 -2714 0 net=13733
rlabel metal2 114 -2716 114 -2716 0 net=6535
rlabel metal2 513 -2716 513 -2716 0 net=8879
rlabel metal2 1073 -2716 1073 -2716 0 net=5268
rlabel metal2 1395 -2716 1395 -2716 0 net=9539
rlabel metal2 184 -2718 184 -2718 0 net=3306
rlabel metal2 1398 -2718 1398 -2718 0 net=13609
rlabel metal2 2060 -2718 2060 -2718 0 net=13891
rlabel metal2 2221 -2718 2221 -2718 0 net=4536
rlabel metal2 75 -2720 75 -2720 0 net=3755
rlabel metal2 226 -2720 226 -2720 0 net=2111
rlabel metal2 478 -2720 478 -2720 0 net=5771
rlabel metal2 877 -2720 877 -2720 0 net=8155
rlabel metal2 1227 -2720 1227 -2720 0 net=8717
rlabel metal2 1433 -2720 1433 -2720 0 net=11404
rlabel metal2 44 -2722 44 -2722 0 net=10489
rlabel metal2 877 -2722 877 -2722 0 net=8577
rlabel metal2 1097 -2722 1097 -2722 0 net=11190
rlabel metal2 2060 -2722 2060 -2722 0 net=13783
rlabel metal2 2214 -2722 2214 -2722 0 net=14683
rlabel metal2 44 -2724 44 -2724 0 net=4301
rlabel metal2 576 -2724 576 -2724 0 net=4283
rlabel metal2 667 -2724 667 -2724 0 net=4699
rlabel metal2 779 -2724 779 -2724 0 net=6787
rlabel metal2 912 -2724 912 -2724 0 net=8329
rlabel metal2 1262 -2724 1262 -2724 0 net=8809
rlabel metal2 1437 -2724 1437 -2724 0 net=11848
rlabel metal2 1962 -2724 1962 -2724 0 net=13203
rlabel metal2 2088 -2724 2088 -2724 0 net=13915
rlabel metal2 135 -2726 135 -2726 0 net=7493
rlabel metal2 933 -2726 933 -2726 0 net=7659
rlabel metal2 1010 -2726 1010 -2726 0 net=8767
rlabel metal2 1244 -2726 1244 -2726 0 net=12573
rlabel metal2 2095 -2726 2095 -2726 0 net=13999
rlabel metal2 142 -2728 142 -2728 0 net=6185
rlabel metal2 688 -2728 688 -2728 0 net=12451
rlabel metal2 142 -2730 142 -2730 0 net=8305
rlabel metal2 226 -2730 226 -2730 0 net=1797
rlabel metal2 352 -2730 352 -2730 0 net=7809
rlabel metal2 583 -2730 583 -2730 0 net=4957
rlabel metal2 583 -2730 583 -2730 0 net=4957
rlabel metal2 604 -2730 604 -2730 0 net=3936
rlabel metal2 1269 -2730 1269 -2730 0 net=8851
rlabel metal2 1437 -2730 1437 -2730 0 net=10055
rlabel metal2 1500 -2730 1500 -2730 0 net=10253
rlabel metal2 1528 -2730 1528 -2730 0 net=10733
rlabel metal2 1626 -2730 1626 -2730 0 net=10897
rlabel metal2 1668 -2730 1668 -2730 0 net=11277
rlabel metal2 1780 -2730 1780 -2730 0 net=11807
rlabel metal2 79 -2732 79 -2732 0 net=3005
rlabel metal2 625 -2732 625 -2732 0 net=5489
rlabel metal2 786 -2732 786 -2732 0 net=14573
rlabel metal2 9 -2734 9 -2734 0 net=9800
rlabel metal2 149 -2734 149 -2734 0 net=1879
rlabel metal2 415 -2734 415 -2734 0 net=10433
rlabel metal2 1073 -2734 1073 -2734 0 net=8019
rlabel metal2 1192 -2734 1192 -2734 0 net=9203
rlabel metal2 1440 -2734 1440 -2734 0 net=14671
rlabel metal2 9 -2736 9 -2736 0 net=8339
rlabel metal2 870 -2736 870 -2736 0 net=8113
rlabel metal2 1290 -2736 1290 -2736 0 net=9127
rlabel metal2 1353 -2736 1353 -2736 0 net=9433
rlabel metal2 1472 -2736 1472 -2736 0 net=9887
rlabel metal2 30 -2738 30 -2738 0 net=2709
rlabel metal2 471 -2738 471 -2738 0 net=4857
rlabel metal2 527 -2738 527 -2738 0 net=3182
rlabel metal2 870 -2738 870 -2738 0 net=8791
rlabel metal2 1087 -2738 1087 -2738 0 net=7615
rlabel metal2 1108 -2738 1108 -2738 0 net=6089
rlabel metal2 1332 -2738 1332 -2738 0 net=9033
rlabel metal2 30 -2740 30 -2740 0 net=2173
rlabel metal2 261 -2740 261 -2740 0 net=2309
rlabel metal2 408 -2740 408 -2740 0 net=8027
rlabel metal2 1115 -2740 1115 -2740 0 net=3290
rlabel metal2 1314 -2740 1314 -2740 0 net=14667
rlabel metal2 54 -2742 54 -2742 0 net=9379
rlabel metal2 1101 -2742 1101 -2742 0 net=5395
rlabel metal2 1367 -2742 1367 -2742 0 net=8927
rlabel metal2 1451 -2742 1451 -2742 0 net=10233
rlabel metal2 1521 -2742 1521 -2742 0 net=10267
rlabel metal2 1580 -2742 1580 -2742 0 net=13253
rlabel metal2 37 -2744 37 -2744 0 net=9697
rlabel metal2 1521 -2744 1521 -2744 0 net=11089
rlabel metal2 1626 -2744 1626 -2744 0 net=10959
rlabel metal2 1850 -2744 1850 -2744 0 net=12409
rlabel metal2 37 -2746 37 -2746 0 net=5363
rlabel metal2 492 -2746 492 -2746 0 net=4371
rlabel metal2 793 -2746 793 -2746 0 net=5739
rlabel metal2 849 -2746 849 -2746 0 net=5747
rlabel metal2 1549 -2746 1549 -2746 0 net=10585
rlabel metal2 1689 -2746 1689 -2746 0 net=11339
rlabel metal2 54 -2748 54 -2748 0 net=12875
rlabel metal2 131 -2750 131 -2750 0 net=2369
rlabel metal2 156 -2750 156 -2750 0 net=2755
rlabel metal2 1570 -2750 1570 -2750 0 net=11053
rlabel metal2 1689 -2750 1689 -2750 0 net=10567
rlabel metal2 170 -2752 170 -2752 0 net=1587
rlabel metal2 408 -2752 408 -2752 0 net=4721
rlabel metal2 450 -2752 450 -2752 0 net=3777
rlabel metal2 625 -2752 625 -2752 0 net=4139
rlabel metal2 968 -2752 968 -2752 0 net=9515
rlabel metal2 1542 -2752 1542 -2752 0 net=10371
rlabel metal2 205 -2754 205 -2754 0 net=1905
rlabel metal2 282 -2754 282 -2754 0 net=1731
rlabel metal2 317 -2754 317 -2754 0 net=1783
rlabel metal2 527 -2754 527 -2754 0 net=2993
rlabel metal2 793 -2754 793 -2754 0 net=1909
rlabel metal2 1542 -2754 1542 -2754 0 net=10509
rlabel metal2 1661 -2754 1661 -2754 0 net=11161
rlabel metal2 205 -2756 205 -2756 0 net=4317
rlabel metal2 233 -2758 233 -2758 0 net=1539
rlabel metal2 289 -2758 289 -2758 0 net=1529
rlabel metal2 411 -2758 411 -2758 0 net=9143
rlabel metal2 1675 -2758 1675 -2758 0 net=11383
rlabel metal2 240 -2760 240 -2760 0 net=6460
rlabel metal2 1255 -2760 1255 -2760 0 net=9832
rlabel metal2 1731 -2760 1731 -2760 0 net=13541
rlabel metal2 243 -2762 243 -2762 0 net=1598
rlabel metal2 443 -2762 443 -2762 0 net=2605
rlabel metal2 744 -2762 744 -2762 0 net=6713
rlabel metal2 982 -2762 982 -2762 0 net=6851
rlabel metal2 1059 -2762 1059 -2762 0 net=7471
rlabel metal2 1514 -2762 1514 -2762 0 net=11363
rlabel metal2 1857 -2762 1857 -2762 0 net=12463
rlabel metal2 212 -2764 212 -2764 0 net=5927
rlabel metal2 464 -2764 464 -2764 0 net=2465
rlabel metal2 1115 -2764 1115 -2764 0 net=7799
rlabel metal2 1724 -2764 1724 -2764 0 net=11433
rlabel metal2 1878 -2764 1878 -2764 0 net=14011
rlabel metal2 212 -2766 212 -2766 0 net=2131
rlabel metal2 310 -2766 310 -2766 0 net=4187
rlabel metal2 597 -2766 597 -2766 0 net=10005
rlabel metal2 1738 -2766 1738 -2766 0 net=11717
rlabel metal2 177 -2768 177 -2768 0 net=3693
rlabel metal2 621 -2768 621 -2768 0 net=4873
rlabel metal2 789 -2768 789 -2768 0 net=14201
rlabel metal2 177 -2770 177 -2770 0 net=5903
rlabel metal2 943 -2770 943 -2770 0 net=11915
rlabel metal2 247 -2772 247 -2772 0 net=4685
rlabel metal2 324 -2772 324 -2772 0 net=2561
rlabel metal2 541 -2772 541 -2772 0 net=9081
rlabel metal2 1465 -2772 1465 -2772 0 net=10213
rlabel metal2 1496 -2772 1496 -2772 0 net=11721
rlabel metal2 289 -2774 289 -2774 0 net=5035
rlabel metal2 639 -2774 639 -2774 0 net=2799
rlabel metal2 744 -2774 744 -2774 0 net=10599
rlabel metal2 296 -2776 296 -2776 0 net=2581
rlabel metal2 569 -2776 569 -2776 0 net=5125
rlabel metal2 688 -2776 688 -2776 0 net=6405
rlabel metal2 947 -2776 947 -2776 0 net=8343
rlabel metal2 1122 -2776 1122 -2776 0 net=9039
rlabel metal2 1493 -2776 1493 -2776 0 net=12184
rlabel metal2 72 -2778 72 -2778 0 net=5695
rlabel metal2 460 -2778 460 -2778 0 net=8085
rlabel metal2 1125 -2778 1125 -2778 0 net=12082
rlabel metal2 72 -2780 72 -2780 0 net=4373
rlabel metal2 268 -2780 268 -2780 0 net=7017
rlabel metal2 702 -2780 702 -2780 0 net=4149
rlabel metal2 1710 -2780 1710 -2780 0 net=12379
rlabel metal2 198 -2782 198 -2782 0 net=6509
rlabel metal2 961 -2782 961 -2782 0 net=13536
rlabel metal2 198 -2784 198 -2784 0 net=2295
rlabel metal2 1794 -2784 1794 -2784 0 net=12067
rlabel metal2 2039 -2784 2039 -2784 0 net=13715
rlabel metal2 219 -2786 219 -2786 0 net=1641
rlabel metal2 611 -2786 611 -2786 0 net=3959
rlabel metal2 789 -2786 789 -2786 0 net=11009
rlabel metal2 1794 -2786 1794 -2786 0 net=11975
rlabel metal2 2074 -2786 2074 -2786 0 net=13591
rlabel metal2 100 -2788 100 -2788 0 net=3983
rlabel metal2 800 -2788 800 -2788 0 net=10162
rlabel metal2 1703 -2788 1703 -2788 0 net=14621
rlabel metal2 100 -2790 100 -2790 0 net=9591
rlabel metal2 380 -2790 380 -2790 0 net=2067
rlabel metal2 807 -2790 807 -2790 0 net=13575
rlabel metal2 219 -2792 219 -2792 0 net=6359
rlabel metal2 940 -2792 940 -2792 0 net=12439
rlabel metal2 380 -2794 380 -2794 0 net=5521
rlabel metal2 807 -2794 807 -2794 0 net=8101
rlabel metal2 835 -2794 835 -2794 0 net=4550
rlabel metal2 1003 -2794 1003 -2794 0 net=5557
rlabel metal2 1164 -2794 1164 -2794 0 net=8253
rlabel metal2 810 -2796 810 -2796 0 net=14608
rlabel metal2 814 -2798 814 -2798 0 net=7956
rlabel metal2 2186 -2798 2186 -2798 0 net=14559
rlabel metal2 544 -2800 544 -2800 0 net=14631
rlabel metal2 814 -2802 814 -2802 0 net=5515
rlabel metal2 1017 -2802 1017 -2802 0 net=7299
rlabel metal2 1199 -2802 1199 -2802 0 net=7907
rlabel metal2 1381 -2802 1381 -2802 0 net=9631
rlabel metal2 394 -2804 394 -2804 0 net=6019
rlabel metal2 1024 -2804 1024 -2804 0 net=7769
rlabel metal2 394 -2806 394 -2806 0 net=3603
rlabel metal2 821 -2806 821 -2806 0 net=6023
rlabel metal2 1080 -2806 1080 -2806 0 net=7543
rlabel metal2 1339 -2806 1339 -2806 0 net=9151
rlabel metal2 1409 -2806 1409 -2806 0 net=10841
rlabel metal2 618 -2808 618 -2808 0 net=8801
rlabel metal2 1346 -2808 1346 -2808 0 net=13126
rlabel metal2 824 -2810 824 -2810 0 net=11903
rlabel metal2 1969 -2810 1969 -2810 0 net=13363
rlabel metal2 828 -2812 828 -2812 0 net=7123
rlabel metal2 1409 -2812 1409 -2812 0 net=9295
rlabel metal2 1815 -2812 1815 -2812 0 net=11945
rlabel metal2 835 -2814 835 -2814 0 net=12386
rlabel metal2 1052 -2814 1052 -2814 0 net=12078
rlabel metal2 191 -2816 191 -2816 0 net=7449
rlabel metal2 1815 -2816 1815 -2816 0 net=12109
rlabel metal2 1836 -2816 1836 -2816 0 net=12865
rlabel metal2 191 -2818 191 -2818 0 net=3219
rlabel metal2 866 -2818 866 -2818 0 net=14165
rlabel metal2 275 -2820 275 -2820 0 net=4509
rlabel metal2 894 -2820 894 -2820 0 net=9715
rlabel metal2 1535 -2820 1535 -2820 0 net=10377
rlabel metal2 275 -2822 275 -2822 0 net=3557
rlabel metal2 905 -2822 905 -2822 0 net=9053
rlabel metal2 1822 -2822 1822 -2822 0 net=12263
rlabel metal2 485 -2824 485 -2824 0 net=2743
rlabel metal2 989 -2824 989 -2824 0 net=9985
rlabel metal2 1829 -2824 1829 -2824 0 net=13401
rlabel metal2 429 -2826 429 -2826 0 net=4617
rlabel metal2 989 -2826 989 -2826 0 net=9529
rlabel metal2 1304 -2826 1304 -2826 0 net=9059
rlabel metal2 1997 -2826 1997 -2826 0 net=13555
rlabel metal2 240 -2828 240 -2828 0 net=2235
rlabel metal2 2025 -2828 2025 -2828 0 net=13673
rlabel metal2 1941 -2830 1941 -2830 0 net=13835
rlabel metal2 222 -2832 222 -2832 0 net=13041
rlabel metal2 23 -2843 23 -2843 0 net=4058
rlabel metal2 541 -2843 541 -2843 0 net=320
rlabel metal2 1500 -2843 1500 -2843 0 net=4150
rlabel metal2 23 -2845 23 -2845 0 net=3757
rlabel metal2 219 -2845 219 -2845 0 net=5522
rlabel metal2 429 -2845 429 -2845 0 net=4372
rlabel metal2 548 -2845 548 -2845 0 net=3343
rlabel metal2 814 -2845 814 -2845 0 net=5516
rlabel metal2 943 -2845 943 -2845 0 net=9034
rlabel metal2 1346 -2845 1346 -2845 0 net=10782
rlabel metal2 1682 -2845 1682 -2845 0 net=14094
rlabel metal2 2144 -2845 2144 -2845 0 net=14345
rlabel metal2 2144 -2845 2144 -2845 0 net=14345
rlabel metal2 2221 -2845 2221 -2845 0 net=7514
rlabel metal2 30 -2847 30 -2847 0 net=2174
rlabel metal2 548 -2847 548 -2847 0 net=6343
rlabel metal2 919 -2847 919 -2847 0 net=6282
rlabel metal2 1202 -2847 1202 -2847 0 net=1088
rlabel metal2 1255 -2847 1255 -2847 0 net=9145
rlabel metal2 1332 -2847 1332 -2847 0 net=10943
rlabel metal2 1682 -2847 1682 -2847 0 net=13785
rlabel metal2 2074 -2847 2074 -2847 0 net=13593
rlabel metal2 30 -2849 30 -2849 0 net=9305
rlabel metal2 317 -2849 317 -2849 0 net=1784
rlabel metal2 828 -2849 828 -2849 0 net=7125
rlabel metal2 922 -2849 922 -2849 0 net=10641
rlabel metal2 1566 -2849 1566 -2849 0 net=11536
rlabel metal2 2060 -2849 2060 -2849 0 net=14669
rlabel metal2 51 -2851 51 -2851 0 net=5772
rlabel metal2 492 -2851 492 -2851 0 net=2995
rlabel metal2 544 -2851 544 -2851 0 net=776
rlabel metal2 964 -2851 964 -2851 0 net=9366
rlabel metal2 1258 -2851 1258 -2851 0 net=10378
rlabel metal2 2004 -2851 2004 -2851 0 net=14113
rlabel metal2 82 -2853 82 -2853 0 net=4722
rlabel metal2 436 -2853 436 -2853 0 net=2215
rlabel metal2 436 -2853 436 -2853 0 net=2215
rlabel metal2 457 -2853 457 -2853 0 net=2745
rlabel metal2 527 -2853 527 -2853 0 net=4745
rlabel metal2 744 -2853 744 -2853 0 net=5740
rlabel metal2 863 -2853 863 -2853 0 net=13204
rlabel metal2 2074 -2853 2074 -2853 0 net=14673
rlabel metal2 103 -2855 103 -2855 0 net=7810
rlabel metal2 373 -2855 373 -2855 0 net=2021
rlabel metal2 460 -2855 460 -2855 0 net=2444
rlabel metal2 565 -2855 565 -2855 0 net=7725
rlabel metal2 968 -2855 968 -2855 0 net=6714
rlabel metal2 975 -2855 975 -2855 0 net=9517
rlabel metal2 1391 -2855 1391 -2855 0 net=11340
rlabel metal2 1983 -2855 1983 -2855 0 net=13917
rlabel metal2 2098 -2855 2098 -2855 0 net=1853
rlabel metal2 107 -2857 107 -2857 0 net=2112
rlabel metal2 401 -2857 401 -2857 0 net=5929
rlabel metal2 835 -2857 835 -2857 0 net=7451
rlabel metal2 968 -2857 968 -2857 0 net=6853
rlabel metal2 1017 -2857 1017 -2857 0 net=7300
rlabel metal2 1062 -2857 1062 -2857 0 net=7616
rlabel metal2 1136 -2857 1136 -2857 0 net=11587
rlabel metal2 1703 -2857 1703 -2857 0 net=11808
rlabel metal2 2088 -2857 2088 -2857 0 net=14705
rlabel metal2 117 -2859 117 -2859 0 net=12452
rlabel metal2 2032 -2859 2032 -2859 0 net=14393
rlabel metal2 124 -2861 124 -2861 0 net=10490
rlabel metal2 866 -2861 866 -2861 0 net=1275
rlabel metal2 1234 -2861 1234 -2861 0 net=9129
rlabel metal2 1314 -2861 1314 -2861 0 net=11956
rlabel metal2 1703 -2861 1703 -2861 0 net=11771
rlabel metal2 1850 -2861 1850 -2861 0 net=13557
rlabel metal2 191 -2863 191 -2863 0 net=3221
rlabel metal2 485 -2863 485 -2863 0 net=4619
rlabel metal2 597 -2863 597 -2863 0 net=10006
rlabel metal2 674 -2863 674 -2863 0 net=7019
rlabel metal2 1017 -2863 1017 -2863 0 net=13267
rlabel metal2 1283 -2863 1283 -2863 0 net=9633
rlabel metal2 1433 -2863 1433 -2863 0 net=10372
rlabel metal2 1731 -2863 1731 -2863 0 net=13543
rlabel metal2 128 -2865 128 -2865 0 net=4007
rlabel metal2 611 -2865 611 -2865 0 net=3984
rlabel metal2 1286 -2865 1286 -2865 0 net=11156
rlabel metal2 1706 -2865 1706 -2865 0 net=13426
rlabel metal2 86 -2867 86 -2867 0 net=9993
rlabel metal2 191 -2867 191 -2867 0 net=2133
rlabel metal2 219 -2867 219 -2867 0 net=2607
rlabel metal2 485 -2867 485 -2867 0 net=2923
rlabel metal2 583 -2867 583 -2867 0 net=4959
rlabel metal2 621 -2867 621 -2867 0 net=2068
rlabel metal2 856 -2867 856 -2867 0 net=8769
rlabel metal2 1290 -2867 1290 -2867 0 net=9153
rlabel metal2 1346 -2867 1346 -2867 0 net=10235
rlabel metal2 1486 -2867 1486 -2867 0 net=12410
rlabel metal2 86 -2869 86 -2869 0 net=5445
rlabel metal2 250 -2869 250 -2869 0 net=9698
rlabel metal2 1419 -2869 1419 -2869 0 net=10607
rlabel metal2 1489 -2869 1489 -2869 0 net=11575
rlabel metal2 1696 -2869 1696 -2869 0 net=12111
rlabel metal2 1878 -2869 1878 -2869 0 net=14013
rlabel metal2 2018 -2869 2018 -2869 0 net=14203
rlabel metal2 72 -2871 72 -2871 0 net=4375
rlabel metal2 289 -2871 289 -2871 0 net=5037
rlabel metal2 324 -2871 324 -2871 0 net=2583
rlabel metal2 443 -2871 443 -2871 0 net=4859
rlabel metal2 499 -2871 499 -2871 0 net=3007
rlabel metal2 674 -2871 674 -2871 0 net=4497
rlabel metal2 1314 -2871 1314 -2871 0 net=14612
rlabel metal2 58 -2873 58 -2873 0 net=1945
rlabel metal2 135 -2873 135 -2873 0 net=7495
rlabel metal2 681 -2873 681 -2873 0 net=7674
rlabel metal2 1038 -2873 1038 -2873 0 net=2204
rlabel metal2 1360 -2873 1360 -2873 0 net=7540
rlabel metal2 1374 -2873 1374 -2873 0 net=9751
rlabel metal2 1451 -2873 1451 -2873 0 net=14560
rlabel metal2 58 -2875 58 -2875 0 net=8803
rlabel metal2 1339 -2875 1339 -2875 0 net=8929
rlabel metal2 1381 -2875 1381 -2875 0 net=10057
rlabel metal2 1493 -2875 1493 -2875 0 net=1179
rlabel metal2 1717 -2875 1717 -2875 0 net=12465
rlabel metal2 1892 -2875 1892 -2875 0 net=13461
rlabel metal2 2109 -2875 2109 -2875 0 net=14755
rlabel metal2 100 -2877 100 -2877 0 net=9593
rlabel metal2 1402 -2877 1402 -2877 0 net=9297
rlabel metal2 1437 -2877 1437 -2877 0 net=9979
rlabel metal2 100 -2879 100 -2879 0 net=13511
rlabel metal2 1752 -2879 1752 -2879 0 net=12538
rlabel metal2 1976 -2879 1976 -2879 0 net=14579
rlabel metal2 110 -2881 110 -2881 0 net=10281
rlabel metal2 1493 -2881 1493 -2881 0 net=10511
rlabel metal2 1556 -2881 1556 -2881 0 net=11011
rlabel metal2 1752 -2881 1752 -2881 0 net=12709
rlabel metal2 1906 -2881 1906 -2881 0 net=13611
rlabel metal2 2123 -2881 2123 -2881 0 net=14353
rlabel metal2 135 -2883 135 -2883 0 net=4285
rlabel metal2 583 -2883 583 -2883 0 net=5749
rlabel metal2 880 -2883 880 -2883 0 net=5396
rlabel metal2 1115 -2883 1115 -2883 0 net=7801
rlabel metal2 1444 -2883 1444 -2883 0 net=11031
rlabel metal2 1640 -2883 1640 -2883 0 net=11729
rlabel metal2 1773 -2883 1773 -2883 0 net=12745
rlabel metal2 2011 -2883 2011 -2883 0 net=14167
rlabel metal2 65 -2885 65 -2885 0 net=6567
rlabel metal2 961 -2885 961 -2885 0 net=3623
rlabel metal2 205 -2887 205 -2887 0 net=4319
rlabel metal2 520 -2887 520 -2887 0 net=6399
rlabel metal2 1059 -2887 1059 -2887 0 net=9884
rlabel metal2 1755 -2887 1755 -2887 0 net=11946
rlabel metal2 2 -2889 2 -2889 0 net=8393
rlabel metal2 212 -2889 212 -2889 0 net=4148
rlabel metal2 642 -2889 642 -2889 0 net=10411
rlabel metal2 1759 -2889 1759 -2889 0 net=13403
rlabel metal2 1871 -2889 1871 -2889 0 net=13037
rlabel metal2 222 -2891 222 -2891 0 net=13576
rlabel metal2 233 -2893 233 -2893 0 net=4686
rlabel metal2 310 -2893 310 -2893 0 net=4189
rlabel metal2 373 -2893 373 -2893 0 net=2711
rlabel metal2 576 -2893 576 -2893 0 net=9717
rlabel metal2 1444 -2893 1444 -2893 0 net=10395
rlabel metal2 1801 -2893 1801 -2893 0 net=12069
rlabel metal2 1990 -2893 1990 -2893 0 net=14001
rlabel metal2 233 -2895 233 -2895 0 net=1643
rlabel metal2 289 -2895 289 -2895 0 net=4511
rlabel metal2 590 -2895 590 -2895 0 net=3695
rlabel metal2 688 -2895 688 -2895 0 net=6407
rlabel metal2 961 -2895 961 -2895 0 net=3375
rlabel metal2 163 -2897 163 -2897 0 net=2261
rlabel metal2 275 -2897 275 -2897 0 net=3559
rlabel metal2 590 -2897 590 -2897 0 net=8103
rlabel metal2 978 -2897 978 -2897 0 net=13313
rlabel metal2 2046 -2897 2046 -2897 0 net=14447
rlabel metal2 163 -2899 163 -2899 0 net=7661
rlabel metal2 1010 -2899 1010 -2899 0 net=10435
rlabel metal2 1479 -2899 1479 -2899 0 net=10735
rlabel metal2 1801 -2899 1801 -2899 0 net=13043
rlabel metal2 236 -2901 236 -2901 0 net=3939
rlabel metal2 310 -2901 310 -2901 0 net=2563
rlabel metal2 632 -2901 632 -2901 0 net=6235
rlabel metal2 730 -2901 730 -2901 0 net=688
rlabel metal2 1598 -2901 1598 -2901 0 net=10843
rlabel metal2 1815 -2901 1815 -2901 0 net=12867
rlabel metal2 1941 -2901 1941 -2901 0 net=13717
rlabel metal2 16 -2903 16 -2903 0 net=5975
rlabel metal2 744 -2903 744 -2903 0 net=8021
rlabel metal2 1087 -2903 1087 -2903 0 net=8087
rlabel metal2 1199 -2903 1199 -2903 0 net=7909
rlabel metal2 2039 -2903 2039 -2903 0 net=14417
rlabel metal2 37 -2905 37 -2905 0 net=5365
rlabel metal2 747 -2905 747 -2905 0 net=6510
rlabel metal2 954 -2905 954 -2905 0 net=5198
rlabel metal2 1241 -2905 1241 -2905 0 net=9041
rlabel metal2 1360 -2905 1360 -2905 0 net=11090
rlabel metal2 1612 -2905 1612 -2905 0 net=11385
rlabel metal2 1829 -2905 1829 -2905 0 net=13139
rlabel metal2 37 -2907 37 -2907 0 net=8307
rlabel metal2 275 -2907 275 -2907 0 net=1531
rlabel metal2 380 -2907 380 -2907 0 net=2851
rlabel metal2 737 -2907 737 -2907 0 net=12289
rlabel metal2 1836 -2907 1836 -2907 0 net=12877
rlabel metal2 142 -2909 142 -2909 0 net=8299
rlabel metal2 772 -2909 772 -2909 0 net=8057
rlabel metal2 933 -2909 933 -2909 0 net=8747
rlabel metal2 1101 -2909 1101 -2909 0 net=8219
rlabel metal2 1248 -2909 1248 -2909 0 net=9001
rlabel metal2 1297 -2909 1297 -2909 0 net=9541
rlabel metal2 1521 -2909 1521 -2909 0 net=10961
rlabel metal2 1913 -2909 1913 -2909 0 net=13675
rlabel metal2 324 -2911 324 -2911 0 net=3605
rlabel metal2 415 -2911 415 -2911 0 net=5253
rlabel metal2 1066 -2911 1066 -2911 0 net=7903
rlabel metal2 1388 -2911 1388 -2911 0 net=10215
rlabel metal2 2025 -2911 2025 -2911 0 net=14259
rlabel metal2 44 -2913 44 -2913 0 net=4302
rlabel metal2 1069 -2913 1069 -2913 0 net=10898
rlabel metal2 2130 -2913 2130 -2913 0 net=9889
rlabel metal2 44 -2915 44 -2915 0 net=1549
rlabel metal2 646 -2915 646 -2915 0 net=6187
rlabel metal2 842 -2915 842 -2915 0 net=10757
rlabel metal2 1276 -2915 1276 -2915 0 net=9435
rlabel metal2 1395 -2915 1395 -2915 0 net=10255
rlabel metal2 1654 -2915 1654 -2915 0 net=10569
rlabel metal2 9 -2917 9 -2917 0 net=8341
rlabel metal2 660 -2917 660 -2917 0 net=11633
rlabel metal2 1689 -2917 1689 -2917 0 net=11723
rlabel metal2 198 -2919 198 -2919 0 net=2297
rlabel metal2 422 -2919 422 -2919 0 net=2467
rlabel metal2 562 -2919 562 -2919 0 net=1953
rlabel metal2 663 -2919 663 -2919 0 net=7775
rlabel metal2 954 -2919 954 -2919 0 net=9759
rlabel metal2 1045 -2919 1045 -2919 0 net=9381
rlabel metal2 1507 -2919 1507 -2919 0 net=10685
rlabel metal2 1745 -2919 1745 -2919 0 net=12575
rlabel metal2 65 -2921 65 -2921 0 net=5639
rlabel metal2 506 -2921 506 -2921 0 net=6872
rlabel metal2 663 -2921 663 -2921 0 net=7472
rlabel metal2 1465 -2921 1465 -2921 0 net=10601
rlabel metal2 1710 -2921 1710 -2921 0 net=12381
rlabel metal2 121 -2923 121 -2923 0 net=4361
rlabel metal2 688 -2923 688 -2923 0 net=8331
rlabel metal2 1178 -2923 1178 -2923 0 net=9061
rlabel metal2 1430 -2923 1430 -2923 0 net=11241
rlabel metal2 1710 -2923 1710 -2923 0 net=11977
rlabel metal2 121 -2925 121 -2925 0 net=3523
rlabel metal2 331 -2925 331 -2925 0 net=1881
rlabel metal2 702 -2925 702 -2925 0 net=8114
rlabel metal2 1171 -2925 1171 -2925 0 net=8655
rlabel metal2 1304 -2925 1304 -2925 0 net=12441
rlabel metal2 149 -2927 149 -2927 0 net=2371
rlabel metal2 240 -2927 240 -2927 0 net=2237
rlabel metal2 345 -2927 345 -2927 0 net=1751
rlabel metal2 387 -2927 387 -2927 0 net=6395
rlabel metal2 1073 -2927 1073 -2927 0 net=8157
rlabel metal2 1213 -2927 1213 -2927 0 net=8811
rlabel metal2 1430 -2927 1430 -2927 0 net=10269
rlabel metal2 1570 -2927 1570 -2927 0 net=11055
rlabel metal2 1794 -2927 1794 -2927 0 net=13227
rlabel metal2 149 -2929 149 -2929 0 net=7771
rlabel metal2 1031 -2929 1031 -2929 0 net=8345
rlabel metal2 1080 -2929 1080 -2929 0 net=7545
rlabel metal2 1528 -2929 1528 -2929 0 net=11353
rlabel metal2 1843 -2929 1843 -2929 0 net=13255
rlabel metal2 156 -2931 156 -2931 0 net=2757
rlabel metal2 345 -2931 345 -2931 0 net=1911
rlabel metal2 989 -2931 989 -2931 0 net=9531
rlabel metal2 1080 -2931 1080 -2931 0 net=11163
rlabel metal2 1955 -2931 1955 -2931 0 net=13837
rlabel metal2 513 -2933 513 -2933 0 net=8881
rlabel metal2 1192 -2933 1192 -2933 0 net=9205
rlabel metal2 1514 -2933 1514 -2933 0 net=11365
rlabel metal2 1661 -2933 1661 -2933 0 net=11719
rlabel metal2 1962 -2933 1962 -2933 0 net=13893
rlabel metal2 296 -2935 296 -2935 0 net=5697
rlabel metal2 569 -2935 569 -2935 0 net=5127
rlabel metal2 705 -2935 705 -2935 0 net=6020
rlabel metal2 989 -2935 989 -2935 0 net=7743
rlabel metal2 1094 -2935 1094 -2935 0 net=7157
rlabel metal2 1192 -2935 1192 -2935 0 net=8853
rlabel metal2 1514 -2935 1514 -2935 0 net=10797
rlabel metal2 1738 -2935 1738 -2935 0 net=12489
rlabel metal2 54 -2937 54 -2937 0 net=9383
rlabel metal2 1605 -2937 1605 -2937 0 net=11279
rlabel metal2 2067 -2937 2067 -2937 0 net=14633
rlabel metal2 170 -2939 170 -2939 0 net=1588
rlabel metal2 709 -2939 709 -2939 0 net=3451
rlabel metal2 1010 -2939 1010 -2939 0 net=8535
rlabel metal2 1668 -2939 1668 -2939 0 net=11917
rlabel metal2 2081 -2939 2081 -2939 0 net=14685
rlabel metal2 170 -2941 170 -2941 0 net=1541
rlabel metal2 296 -2941 296 -2941 0 net=1895
rlabel metal2 695 -2941 695 -2941 0 net=4395
rlabel metal2 740 -2941 740 -2941 0 net=13751
rlabel metal2 254 -2943 254 -2943 0 net=1907
rlabel metal2 667 -2943 667 -2943 0 net=4701
rlabel metal2 751 -2943 751 -2943 0 net=4874
rlabel metal2 1787 -2943 1787 -2943 0 net=12975
rlabel metal2 16 -2945 16 -2945 0 net=3703
rlabel metal2 261 -2945 261 -2945 0 net=2311
rlabel metal2 667 -2945 667 -2945 0 net=6111
rlabel metal2 177 -2947 177 -2947 0 net=5905
rlabel metal2 765 -2947 765 -2947 0 net=6091
rlabel metal2 1157 -2947 1157 -2947 0 net=13573
rlabel metal2 177 -2949 177 -2949 0 net=4171
rlabel metal2 226 -2949 226 -2949 0 net=1799
rlabel metal2 772 -2949 772 -2949 0 net=5559
rlabel metal2 1115 -2949 1115 -2949 0 net=8255
rlabel metal2 1206 -2949 1206 -2949 0 net=9986
rlabel metal2 1563 -2949 1563 -2949 0 net=11025
rlabel metal2 159 -2951 159 -2951 0 net=3837
rlabel metal2 779 -2951 779 -2951 0 net=6789
rlabel metal2 870 -2951 870 -2951 0 net=8793
rlabel metal2 1150 -2951 1150 -2951 0 net=8417
rlabel metal2 1535 -2951 1535 -2951 0 net=11435
rlabel metal2 779 -2953 779 -2953 0 net=8579
rlabel metal2 905 -2953 905 -2953 0 net=9055
rlabel metal2 1185 -2953 1185 -2953 0 net=8449
rlabel metal2 1647 -2953 1647 -2953 0 net=11905
rlabel metal2 93 -2955 93 -2955 0 net=7137
rlabel metal2 1097 -2955 1097 -2955 0 net=9445
rlabel metal2 1724 -2955 1724 -2955 0 net=12265
rlabel metal2 79 -2957 79 -2957 0 net=4121
rlabel metal2 793 -2957 793 -2957 0 net=6025
rlabel metal2 870 -2957 870 -2957 0 net=6361
rlabel metal2 1780 -2957 1780 -2957 0 net=12931
rlabel metal2 79 -2959 79 -2959 0 net=8273
rlabel metal2 1822 -2959 1822 -2959 0 net=13365
rlabel metal2 114 -2961 114 -2961 0 net=6537
rlabel metal2 996 -2961 996 -2961 0 net=8029
rlabel metal2 1927 -2961 1927 -2961 0 net=13735
rlabel metal2 114 -2963 114 -2963 0 net=3778
rlabel metal2 758 -2963 758 -2963 0 net=5491
rlabel metal2 1108 -2963 1108 -2963 0 net=8719
rlabel metal2 1808 -2963 1808 -2963 0 net=14623
rlabel metal2 450 -2965 450 -2965 0 net=7201
rlabel metal2 1227 -2965 1227 -2965 0 net=9083
rlabel metal2 1808 -2965 1808 -2965 0 net=12785
rlabel metal2 1969 -2965 1969 -2965 0 net=14575
rlabel metal2 653 -2967 653 -2967 0 net=5461
rlabel metal2 1318 -2967 1318 -2967 0 net=10587
rlabel metal2 1766 -2967 1766 -2967 0 net=13601
rlabel metal2 639 -2969 639 -2969 0 net=3961
rlabel metal2 1160 -2969 1160 -2969 0 net=10399
rlabel metal2 282 -2971 282 -2971 0 net=1732
rlabel metal2 282 -2973 282 -2973 0 net=4141
rlabel metal2 625 -2975 625 -2975 0 net=2801
rlabel metal2 716 -2977 716 -2977 0 net=5685
rlabel metal2 16 -2988 16 -2988 0 net=3704
rlabel metal2 114 -2988 114 -2988 0 net=6397
rlabel metal2 422 -2988 422 -2988 0 net=2468
rlabel metal2 471 -2988 471 -2988 0 net=1883
rlabel metal2 569 -2988 569 -2988 0 net=9518
rlabel metal2 1041 -2988 1041 -2988 0 net=14670
rlabel metal2 2095 -2988 2095 -2988 0 net=13594
rlabel metal2 51 -2990 51 -2990 0 net=1946
rlabel metal2 100 -2990 100 -2990 0 net=8748
rlabel metal2 961 -2990 961 -2990 0 net=6854
rlabel metal2 1052 -2990 1052 -2990 0 net=7904
rlabel metal2 1346 -2990 1346 -2990 0 net=10237
rlabel metal2 1346 -2990 1346 -2990 0 net=10237
rlabel metal2 1360 -2990 1360 -2990 0 net=10283
rlabel metal2 1416 -2990 1416 -2990 0 net=7910
rlabel metal2 1871 -2990 1871 -2990 0 net=13039
rlabel metal2 2098 -2990 2098 -2990 0 net=3624
rlabel metal2 37 -2992 37 -2992 0 net=8309
rlabel metal2 93 -2992 93 -2992 0 net=4123
rlabel metal2 107 -2992 107 -2992 0 net=8581
rlabel metal2 880 -2992 880 -2992 0 net=11724
rlabel metal2 1769 -2992 1769 -2992 0 net=12868
rlabel metal2 1836 -2992 1836 -2992 0 net=12879
rlabel metal2 1871 -2992 1871 -2992 0 net=14003
rlabel metal2 30 -2994 30 -2994 0 net=9306
rlabel metal2 142 -2994 142 -2994 0 net=8300
rlabel metal2 964 -2994 964 -2994 0 net=736
rlabel metal2 1055 -2994 1055 -2994 0 net=14065
rlabel metal2 1892 -2994 1892 -2994 0 net=13463
rlabel metal2 30 -2996 30 -2996 0 net=8805
rlabel metal2 65 -2996 65 -2996 0 net=5640
rlabel metal2 572 -2996 572 -2996 0 net=6951
rlabel metal2 968 -2996 968 -2996 0 net=8089
rlabel metal2 1125 -2996 1125 -2996 0 net=10512
rlabel metal2 1566 -2996 1566 -2996 0 net=13314
rlabel metal2 37 -2998 37 -2998 0 net=6401
rlabel metal2 541 -2998 541 -2998 0 net=5930
rlabel metal2 884 -2998 884 -2998 0 net=3453
rlabel metal2 1031 -2998 1031 -2998 0 net=8451
rlabel metal2 1199 -2998 1199 -2998 0 net=14580
rlabel metal2 44 -3000 44 -3000 0 net=1551
rlabel metal2 135 -3000 135 -3000 0 net=4287
rlabel metal2 590 -3000 590 -3000 0 net=8104
rlabel metal2 954 -3000 954 -3000 0 net=9761
rlabel metal2 1199 -3000 1199 -3000 0 net=9003
rlabel metal2 1318 -3000 1318 -3000 0 net=10589
rlabel metal2 1419 -3000 1419 -3000 0 net=13544
rlabel metal2 1976 -3000 1976 -3000 0 net=1855
rlabel metal2 58 -3002 58 -3002 0 net=2373
rlabel metal2 208 -3002 208 -3002 0 net=4860
rlabel metal2 471 -3002 471 -3002 0 net=4899
rlabel metal2 894 -3002 894 -3002 0 net=12070
rlabel metal2 1885 -3002 1885 -3002 0 net=13919
rlabel metal2 142 -3004 142 -3004 0 net=8395
rlabel metal2 212 -3004 212 -3004 0 net=1908
rlabel metal2 422 -3004 422 -3004 0 net=2585
rlabel metal2 436 -3004 436 -3004 0 net=2217
rlabel metal2 436 -3004 436 -3004 0 net=2217
rlabel metal2 443 -3004 443 -3004 0 net=9437
rlabel metal2 1318 -3004 1318 -3004 0 net=8931
rlabel metal2 1398 -3004 1398 -3004 0 net=13718
rlabel metal2 86 -3006 86 -3006 0 net=5447
rlabel metal2 236 -3006 236 -3006 0 net=8342
rlabel metal2 642 -3006 642 -3006 0 net=5462
rlabel metal2 786 -3006 786 -3006 0 net=3345
rlabel metal2 1055 -3006 1055 -3006 0 net=11772
rlabel metal2 1808 -3006 1808 -3006 0 net=12786
rlabel metal2 1920 -3006 1920 -3006 0 net=14261
rlabel metal2 86 -3008 86 -3008 0 net=2609
rlabel metal2 240 -3008 240 -3008 0 net=2759
rlabel metal2 478 -3008 478 -3008 0 net=4321
rlabel metal2 688 -3008 688 -3008 0 net=8332
rlabel metal2 1066 -3008 1066 -3008 0 net=11019
rlabel metal2 1139 -3008 1139 -3008 0 net=11576
rlabel metal2 1654 -3008 1654 -3008 0 net=10571
rlabel metal2 131 -3010 131 -3010 0 net=6967
rlabel metal2 905 -3010 905 -3010 0 net=7139
rlabel metal2 1038 -3010 1038 -3010 0 net=9447
rlabel metal2 1325 -3010 1325 -3010 0 net=6897
rlabel metal2 1570 -3010 1570 -3010 0 net=12382
rlabel metal2 149 -3012 149 -3012 0 net=7773
rlabel metal2 478 -3012 478 -3012 0 net=6113
rlabel metal2 688 -3012 688 -3012 0 net=9147
rlabel metal2 1339 -3012 1339 -3012 0 net=10271
rlabel metal2 1486 -3012 1486 -3012 0 net=9382
rlabel metal2 1808 -3012 1808 -3012 0 net=14625
rlabel metal2 138 -3014 138 -3014 0 net=2499
rlabel metal2 156 -3014 156 -3014 0 net=1157
rlabel metal2 667 -3014 667 -3014 0 net=4703
rlabel metal2 716 -3014 716 -3014 0 net=5687
rlabel metal2 730 -3014 730 -3014 0 net=5976
rlabel metal2 1045 -3014 1045 -3014 0 net=8347
rlabel metal2 1069 -3014 1069 -3014 0 net=8812
rlabel metal2 1220 -3014 1220 -3014 0 net=9085
rlabel metal2 1255 -3014 1255 -3014 0 net=9385
rlabel metal2 1402 -3014 1402 -3014 0 net=9298
rlabel metal2 1430 -3014 1430 -3014 0 net=10643
rlabel metal2 1570 -3014 1570 -3014 0 net=11281
rlabel metal2 1633 -3014 1633 -3014 0 net=12291
rlabel metal2 1689 -3014 1689 -3014 0 net=12747
rlabel metal2 1815 -3014 1815 -3014 0 net=13753
rlabel metal2 156 -3016 156 -3016 0 net=2135
rlabel metal2 198 -3016 198 -3016 0 net=2313
rlabel metal2 282 -3016 282 -3016 0 net=4143
rlabel metal2 590 -3016 590 -3016 0 net=5129
rlabel metal2 716 -3016 716 -3016 0 net=6791
rlabel metal2 849 -3016 849 -3016 0 net=6569
rlabel metal2 1045 -3016 1045 -3016 0 net=7159
rlabel metal2 1160 -3016 1160 -3016 0 net=7546
rlabel metal2 1402 -3016 1402 -3016 0 net=11354
rlabel metal2 1549 -3016 1549 -3016 0 net=10401
rlabel metal2 1703 -3016 1703 -3016 0 net=12933
rlabel metal2 1864 -3016 1864 -3016 0 net=14419
rlabel metal2 128 -3018 128 -3018 0 net=9994
rlabel metal2 1178 -3018 1178 -3018 0 net=9063
rlabel metal2 1213 -3018 1213 -3018 0 net=7802
rlabel metal2 1486 -3018 1486 -3018 0 net=11027
rlabel metal2 1573 -3018 1573 -3018 0 net=9890
rlabel metal2 159 -3020 159 -3020 0 net=8158
rlabel metal2 1076 -3020 1076 -3020 0 net=9980
rlabel metal2 1493 -3020 1493 -3020 0 net=10963
rlabel metal2 1528 -3020 1528 -3020 0 net=13787
rlabel metal2 1759 -3020 1759 -3020 0 net=13405
rlabel metal2 1874 -3020 1874 -3020 0 net=1
rlabel metal2 1948 -3020 1948 -3020 0 net=14707
rlabel metal2 163 -3022 163 -3022 0 net=7663
rlabel metal2 597 -3022 597 -3022 0 net=4009
rlabel metal2 695 -3022 695 -3022 0 net=4397
rlabel metal2 730 -3022 730 -3022 0 net=11165
rlabel metal2 1083 -3022 1083 -3022 0 net=13574
rlabel metal2 166 -3024 166 -3024 0 net=7020
rlabel metal2 1087 -3024 1087 -3024 0 net=8257
rlabel metal2 1143 -3024 1143 -3024 0 net=12443
rlabel metal2 1353 -3024 1353 -3024 0 net=10257
rlabel metal2 1423 -3024 1423 -3024 0 net=10737
rlabel metal2 1500 -3024 1500 -3024 0 net=11013
rlabel metal2 1654 -3024 1654 -3024 0 net=12577
rlabel metal2 1759 -3024 1759 -3024 0 net=13559
rlabel metal2 1934 -3024 1934 -3024 0 net=14169
rlabel metal2 79 -3026 79 -3026 0 net=8275
rlabel metal2 985 -3026 985 -3026 0 net=14151
rlabel metal2 170 -3028 170 -3028 0 net=1543
rlabel metal2 282 -3028 282 -3028 0 net=2853
rlabel metal2 457 -3028 457 -3028 0 net=2747
rlabel metal2 614 -3028 614 -3028 0 net=6538
rlabel metal2 1178 -3028 1178 -3028 0 net=9043
rlabel metal2 1269 -3028 1269 -3028 0 net=9155
rlabel metal2 1304 -3028 1304 -3028 0 net=10609
rlabel metal2 1549 -3028 1549 -3028 0 net=11387
rlabel metal2 1661 -3028 1661 -3028 0 net=11720
rlabel metal2 1745 -3028 1745 -3028 0 net=13839
rlabel metal2 173 -3030 173 -3030 0 net=7496
rlabel metal2 625 -3030 625 -3030 0 net=2803
rlabel metal2 1192 -3030 1192 -3030 0 net=8855
rlabel metal2 1612 -3030 1612 -3030 0 net=11731
rlabel metal2 1661 -3030 1661 -3030 0 net=12267
rlabel metal2 1766 -3030 1766 -3030 0 net=13257
rlabel metal2 184 -3032 184 -3032 0 net=3525
rlabel metal2 219 -3032 219 -3032 0 net=2713
rlabel metal2 457 -3032 457 -3032 0 net=7547
rlabel metal2 1164 -3032 1164 -3032 0 net=9057
rlabel metal2 1202 -3032 1202 -3032 0 net=10483
rlabel metal2 1437 -3032 1437 -3032 0 net=10799
rlabel metal2 1598 -3032 1598 -3032 0 net=10845
rlabel metal2 1682 -3032 1682 -3032 0 net=6037
rlabel metal2 184 -3034 184 -3034 0 net=11091
rlabel metal2 215 -3034 215 -3034 0 net=4799
rlabel metal2 485 -3034 485 -3034 0 net=2924
rlabel metal2 740 -3034 740 -3034 0 net=6362
rlabel metal2 1136 -3034 1136 -3034 0 net=11675
rlabel metal2 1724 -3034 1724 -3034 0 net=14675
rlabel metal2 240 -3036 240 -3036 0 net=2263
rlabel metal2 296 -3036 296 -3036 0 net=1896
rlabel metal2 702 -3036 702 -3036 0 net=5367
rlabel metal2 737 -3036 737 -3036 0 net=4011
rlabel metal2 1136 -3036 1136 -3036 0 net=9131
rlabel metal2 1241 -3036 1241 -3036 0 net=10217
rlabel metal2 1451 -3036 1451 -3036 0 net=10413
rlabel metal2 1773 -3036 1773 -3036 0 net=13367
rlabel metal2 1843 -3036 1843 -3036 0 net=14115
rlabel metal2 2074 -3036 2074 -3036 0 net=3377
rlabel metal2 254 -3038 254 -3038 0 net=9594
rlabel metal2 1388 -3038 1388 -3038 0 net=12467
rlabel metal2 1822 -3038 1822 -3038 0 net=14205
rlabel metal2 247 -3040 247 -3040 0 net=4377
rlabel metal2 268 -3040 268 -3040 0 net=2077
rlabel metal2 1157 -3040 1157 -3040 0 net=10325
rlabel metal2 1451 -3040 1451 -3040 0 net=13513
rlabel metal2 2004 -3040 2004 -3040 0 net=14687
rlabel metal2 103 -3042 103 -3042 0 net=11193
rlabel metal2 296 -3042 296 -3042 0 net=3223
rlabel metal2 415 -3042 415 -3042 0 net=5255
rlabel metal2 758 -3042 758 -3042 0 net=3417
rlabel metal2 870 -3042 870 -3042 0 net=7777
rlabel metal2 1017 -3042 1017 -3042 0 net=13269
rlabel metal2 275 -3044 275 -3044 0 net=1533
rlabel metal2 415 -3044 415 -3044 0 net=4363
rlabel metal2 513 -3044 513 -3044 0 net=5699
rlabel metal2 835 -3044 835 -3044 0 net=7453
rlabel metal2 1003 -3044 1003 -3044 0 net=8795
rlabel metal2 1059 -3044 1059 -3044 0 net=8221
rlabel metal2 1164 -3044 1164 -3044 0 net=11611
rlabel metal2 1283 -3044 1283 -3044 0 net=9635
rlabel metal2 1332 -3044 1332 -3044 0 net=10945
rlabel metal2 1514 -3044 1514 -3044 0 net=11033
rlabel metal2 1717 -3044 1717 -3044 0 net=13229
rlabel metal2 275 -3046 275 -3046 0 net=3607
rlabel metal2 338 -3046 338 -3046 0 net=1753
rlabel metal2 485 -3046 485 -3046 0 net=4621
rlabel metal2 625 -3046 625 -3046 0 net=4499
rlabel metal2 709 -3046 709 -3046 0 net=5013
rlabel metal2 1097 -3046 1097 -3046 0 net=10239
rlabel metal2 1465 -3046 1465 -3046 0 net=10603
rlabel metal2 289 -3048 289 -3048 0 net=4513
rlabel metal2 660 -3048 660 -3048 0 net=3697
rlabel metal2 765 -3048 765 -3048 0 net=6093
rlabel metal2 884 -3048 884 -3048 0 net=13571
rlabel metal2 1283 -3048 1283 -3048 0 net=9543
rlabel metal2 1465 -3048 1465 -3048 0 net=12491
rlabel metal2 1794 -3048 1794 -3048 0 net=13737
rlabel metal2 289 -3050 289 -3050 0 net=6237
rlabel metal2 674 -3050 674 -3050 0 net=8883
rlabel metal2 1227 -3050 1227 -3050 0 net=9207
rlabel metal2 1297 -3050 1297 -3050 0 net=7237
rlabel metal2 1472 -3050 1472 -3050 0 net=5027
rlabel metal2 310 -3052 310 -3052 0 net=2565
rlabel metal2 506 -3052 506 -3052 0 net=8031
rlabel metal2 1024 -3052 1024 -3052 0 net=9533
rlabel metal2 1311 -3052 1311 -3052 0 net=11436
rlabel metal2 1542 -3052 1542 -3052 0 net=11367
rlabel metal2 1738 -3052 1738 -3052 0 net=13045
rlabel metal2 1927 -3052 1927 -3052 0 net=14635
rlabel metal2 310 -3054 310 -3054 0 net=6047
rlabel metal2 1101 -3054 1101 -3054 0 net=8419
rlabel metal2 1535 -3054 1535 -3054 0 net=11057
rlabel metal2 1801 -3054 1801 -3054 0 net=13613
rlabel metal2 324 -3056 324 -3056 0 net=3009
rlabel metal2 513 -3056 513 -3056 0 net=3561
rlabel metal2 548 -3056 548 -3056 0 net=6344
rlabel metal2 1584 -3056 1584 -3056 0 net=11589
rlabel metal2 1906 -3056 1906 -3056 0 net=14395
rlabel metal2 226 -3058 226 -3058 0 net=3839
rlabel metal2 632 -3058 632 -3058 0 net=6409
rlabel metal2 835 -3058 835 -3058 0 net=10059
rlabel metal2 1591 -3058 1591 -3058 0 net=11635
rlabel metal2 2032 -3058 2032 -3058 0 net=14757
rlabel metal2 121 -3060 121 -3060 0 net=6505
rlabel metal2 352 -3060 352 -3060 0 net=4191
rlabel metal2 681 -3060 681 -3060 0 net=10759
rlabel metal2 940 -3060 940 -3060 0 net=7727
rlabel metal2 1024 -3060 1024 -3060 0 net=8721
rlabel metal2 1122 -3060 1122 -3060 0 net=8857
rlabel metal2 1381 -3060 1381 -3060 0 net=10397
rlabel metal2 1619 -3060 1619 -3060 0 net=11907
rlabel metal2 121 -3062 121 -3062 0 net=9719
rlabel metal2 765 -3062 765 -3062 0 net=8771
rlabel metal2 940 -3062 940 -3062 0 net=9753
rlabel metal2 1626 -3062 1626 -3062 0 net=12113
rlabel metal2 124 -3064 124 -3064 0 net=10949
rlabel metal2 359 -3064 359 -3064 0 net=1801
rlabel metal2 450 -3064 450 -3064 0 net=7203
rlabel metal2 856 -3064 856 -3064 0 net=8059
rlabel metal2 996 -3064 996 -3064 0 net=7675
rlabel metal2 1556 -3064 1556 -3064 0 net=14023
rlabel metal2 359 -3066 359 -3066 0 net=2677
rlabel metal2 576 -3066 576 -3066 0 net=3963
rlabel metal2 772 -3066 772 -3066 0 net=5561
rlabel metal2 1010 -3066 1010 -3066 0 net=8537
rlabel metal2 1129 -3066 1129 -3066 0 net=8657
rlabel metal2 1647 -3066 1647 -3066 0 net=11979
rlabel metal2 366 -3068 366 -3068 0 net=2299
rlabel metal2 450 -3068 450 -3068 0 net=2997
rlabel metal2 499 -3068 499 -3068 0 net=3291
rlabel metal2 1710 -3068 1710 -3068 0 net=12977
rlabel metal2 317 -3070 317 -3070 0 net=5039
rlabel metal2 492 -3070 492 -3070 0 net=1955
rlabel metal2 653 -3070 653 -3070 0 net=7127
rlabel metal2 1034 -3070 1034 -3070 0 net=10551
rlabel metal2 1787 -3070 1787 -3070 0 net=13603
rlabel metal2 177 -3072 177 -3072 0 net=4173
rlabel metal2 527 -3072 527 -3072 0 net=4747
rlabel metal2 611 -3072 611 -3072 0 net=4961
rlabel metal2 744 -3072 744 -3072 0 net=8023
rlabel metal2 1171 -3072 1171 -3072 0 net=8939
rlabel metal2 1899 -3072 1899 -3072 0 net=14015
rlabel metal2 23 -3074 23 -3074 0 net=3758
rlabel metal2 772 -3074 772 -3074 0 net=5493
rlabel metal2 863 -3074 863 -3074 0 net=14576
rlabel metal2 23 -3076 23 -3076 0 net=13845
rlabel metal2 1507 -3076 1507 -3076 0 net=10687
rlabel metal2 177 -3078 177 -3078 0 net=3941
rlabel metal2 331 -3078 331 -3078 0 net=2239
rlabel metal2 982 -3078 982 -3078 0 net=7745
rlabel metal2 1507 -3078 1507 -3078 0 net=11243
rlabel metal2 1913 -3078 1913 -3078 0 net=13677
rlabel metal2 233 -3080 233 -3080 0 net=1645
rlabel metal2 331 -3080 331 -3080 0 net=1913
rlabel metal2 583 -3080 583 -3080 0 net=5751
rlabel metal2 807 -3080 807 -3080 0 net=6189
rlabel metal2 877 -3080 877 -3080 0 net=11447
rlabel metal2 1913 -3080 1913 -3080 0 net=14449
rlabel metal2 345 -3082 345 -3082 0 net=2023
rlabel metal2 583 -3082 583 -3082 0 net=5907
rlabel metal2 793 -3082 793 -3082 0 net=6027
rlabel metal2 989 -3082 989 -3082 0 net=10437
rlabel metal2 2046 -3082 2046 -3082 0 net=14355
rlabel metal2 117 -3084 117 -3084 0 net=4977
rlabel metal2 751 -3084 751 -3084 0 net=5245
rlabel metal2 1458 -3084 1458 -3084 0 net=11919
rlabel metal2 793 -3086 793 -3086 0 net=5655
rlabel metal2 1668 -3086 1668 -3086 0 net=12711
rlabel metal2 1752 -3088 1752 -3088 0 net=13141
rlabel metal2 1829 -3090 1829 -3090 0 net=13895
rlabel metal2 1962 -3092 1962 -3092 0 net=14346
rlabel metal2 23 -3103 23 -3103 0 net=13846
rlabel metal2 212 -3103 212 -3103 0 net=5449
rlabel metal2 303 -3103 303 -3103 0 net=1647
rlabel metal2 303 -3103 303 -3103 0 net=1647
rlabel metal2 380 -3103 380 -3103 0 net=1802
rlabel metal2 520 -3103 520 -3103 0 net=7664
rlabel metal2 821 -3103 821 -3103 0 net=2240
rlabel metal2 1381 -3103 1381 -3103 0 net=10398
rlabel metal2 1461 -3103 1461 -3103 0 net=14420
rlabel metal2 1962 -3103 1962 -3103 0 net=14356
rlabel metal2 30 -3105 30 -3105 0 net=8806
rlabel metal2 212 -3105 212 -3105 0 net=9455
rlabel metal2 1199 -3105 1199 -3105 0 net=9004
rlabel metal2 1276 -3105 1276 -3105 0 net=13514
rlabel metal2 1465 -3105 1465 -3105 0 net=12492
rlabel metal2 1566 -3105 1566 -3105 0 net=757
rlabel metal2 1853 -3105 1853 -3105 0 net=13040
rlabel metal2 1997 -3105 1997 -3105 0 net=13679
rlabel metal2 2046 -3105 2046 -3105 0 net=3379
rlabel metal2 58 -3107 58 -3107 0 net=2374
rlabel metal2 187 -3107 187 -3107 0 net=9148
rlabel metal2 737 -3107 737 -3107 0 net=4012
rlabel metal2 1451 -3107 1451 -3107 0 net=11059
rlabel metal2 1640 -3107 1640 -3107 0 net=10846
rlabel metal2 1892 -3107 1892 -3107 0 net=14709
rlabel metal2 65 -3109 65 -3109 0 net=1552
rlabel metal2 1129 -3109 1129 -3109 0 net=8659
rlabel metal2 1129 -3109 1129 -3109 0 net=8659
rlabel metal2 1199 -3109 1199 -3109 0 net=10611
rlabel metal2 1311 -3109 1311 -3109 0 net=12935
rlabel metal2 1864 -3109 1864 -3109 0 net=14005
rlabel metal2 1878 -3109 1878 -3109 0 net=14017
rlabel metal2 72 -3111 72 -3111 0 net=8310
rlabel metal2 289 -3111 289 -3111 0 net=6239
rlabel metal2 835 -3111 835 -3111 0 net=10060
rlabel metal2 1216 -3111 1216 -3111 0 net=8856
rlabel metal2 1671 -3111 1671 -3111 0 net=12880
rlabel metal2 79 -3113 79 -3113 0 net=8884
rlabel metal2 681 -3113 681 -3113 0 net=10760
rlabel metal2 1234 -3113 1234 -3113 0 net=10238
rlabel metal2 1381 -3113 1381 -3113 0 net=12293
rlabel metal2 1675 -3113 1675 -3113 0 net=10402
rlabel metal2 86 -3115 86 -3115 0 net=2610
rlabel metal2 194 -3115 194 -3115 0 net=2854
rlabel metal2 289 -3115 289 -3115 0 net=1965
rlabel metal2 436 -3115 436 -3115 0 net=2219
rlabel metal2 436 -3115 436 -3115 0 net=2219
rlabel metal2 506 -3115 506 -3115 0 net=8033
rlabel metal2 758 -3115 758 -3115 0 net=3418
rlabel metal2 1857 -3115 1857 -3115 0 net=13921
rlabel metal2 93 -3117 93 -3117 0 net=8397
rlabel metal2 198 -3117 198 -3117 0 net=2315
rlabel metal2 198 -3117 198 -3117 0 net=2315
rlabel metal2 254 -3117 254 -3117 0 net=4379
rlabel metal2 352 -3117 352 -3117 0 net=10951
rlabel metal2 1388 -3117 1388 -3117 0 net=12469
rlabel metal2 1388 -3117 1388 -3117 0 net=12469
rlabel metal2 1395 -3117 1395 -3117 0 net=5028
rlabel metal2 1486 -3117 1486 -3117 0 net=11028
rlabel metal2 1605 -3117 1605 -3117 0 net=14153
rlabel metal2 1885 -3117 1885 -3117 0 net=14263
rlabel metal2 107 -3119 107 -3119 0 net=8582
rlabel metal2 891 -3119 891 -3119 0 net=2804
rlabel metal2 1122 -3119 1122 -3119 0 net=6899
rlabel metal2 1395 -3119 1395 -3119 0 net=12979
rlabel metal2 1920 -3119 1920 -3119 0 net=1857
rlabel metal2 107 -3121 107 -3121 0 net=3943
rlabel metal2 226 -3121 226 -3121 0 net=6507
rlabel metal2 380 -3121 380 -3121 0 net=6511
rlabel metal2 604 -3121 604 -3121 0 net=4748
rlabel metal2 898 -3121 898 -3121 0 net=5563
rlabel metal2 1237 -3121 1237 -3121 0 net=10484
rlabel metal2 1437 -3121 1437 -3121 0 net=10801
rlabel metal2 1633 -3121 1633 -3121 0 net=13605
rlabel metal2 1976 -3121 1976 -3121 0 net=14689
rlabel metal2 114 -3123 114 -3123 0 net=6398
rlabel metal2 177 -3123 177 -3123 0 net=6029
rlabel metal2 828 -3123 828 -3123 0 net=7205
rlabel metal2 926 -3123 926 -3123 0 net=8277
rlabel metal2 926 -3123 926 -3123 0 net=8277
rlabel metal2 943 -3123 943 -3123 0 net=14676
rlabel metal2 100 -3125 100 -3125 0 net=4124
rlabel metal2 121 -3125 121 -3125 0 net=9720
rlabel metal2 254 -3125 254 -3125 0 net=2679
rlabel metal2 401 -3125 401 -3125 0 net=1534
rlabel metal2 555 -3125 555 -3125 0 net=4514
rlabel metal2 877 -3125 877 -3125 0 net=7197
rlabel metal2 1465 -3125 1465 -3125 0 net=11733
rlabel metal2 1647 -3125 1647 -3125 0 net=11981
rlabel metal2 100 -3127 100 -3127 0 net=6049
rlabel metal2 359 -3127 359 -3127 0 net=2301
rlabel metal2 373 -3127 373 -3127 0 net=4801
rlabel metal2 569 -3127 569 -3127 0 net=4144
rlabel metal2 828 -3127 828 -3127 0 net=9065
rlabel metal2 1248 -3127 1248 -3127 0 net=9156
rlabel metal2 1276 -3127 1276 -3127 0 net=5991
rlabel metal2 121 -3129 121 -3129 0 net=2137
rlabel metal2 191 -3129 191 -3129 0 net=3527
rlabel metal2 275 -3129 275 -3129 0 net=3608
rlabel metal2 404 -3129 404 -3129 0 net=3107
rlabel metal2 471 -3129 471 -3129 0 net=4901
rlabel metal2 625 -3129 625 -3129 0 net=4500
rlabel metal2 1094 -3129 1094 -3129 0 net=11020
rlabel metal2 1185 -3129 1185 -3129 0 net=9763
rlabel metal2 1297 -3129 1297 -3129 0 net=7238
rlabel metal2 1318 -3129 1318 -3129 0 net=8932
rlabel metal2 1647 -3129 1647 -3129 0 net=10604
rlabel metal2 135 -3131 135 -3131 0 net=10543
rlabel metal2 296 -3131 296 -3131 0 net=3225
rlabel metal2 471 -3131 471 -3131 0 net=3841
rlabel metal2 541 -3131 541 -3131 0 net=4289
rlabel metal2 625 -3131 625 -3131 0 net=5015
rlabel metal2 716 -3131 716 -3131 0 net=6793
rlabel metal2 863 -3131 863 -3131 0 net=7141
rlabel metal2 961 -3131 961 -3131 0 net=6953
rlabel metal2 135 -3133 135 -3133 0 net=2079
rlabel metal2 310 -3133 310 -3133 0 net=4175
rlabel metal2 366 -3133 366 -3133 0 net=2761
rlabel metal2 443 -3133 443 -3133 0 net=9439
rlabel metal2 758 -3133 758 -3133 0 net=3347
rlabel metal2 961 -3133 961 -3133 0 net=8453
rlabel metal2 1045 -3133 1045 -3133 0 net=7161
rlabel metal2 142 -3135 142 -3135 0 net=13175
rlabel metal2 968 -3135 968 -3135 0 net=8090
rlabel metal2 1612 -3135 1612 -3135 0 net=14207
rlabel metal2 156 -3137 156 -3137 0 net=7465
rlabel metal2 219 -3137 219 -3137 0 net=2715
rlabel metal2 317 -3137 317 -3137 0 net=1915
rlabel metal2 429 -3137 429 -3137 0 net=2749
rlabel metal2 632 -3137 632 -3137 0 net=6411
rlabel metal2 856 -3137 856 -3137 0 net=8061
rlabel metal2 968 -3137 968 -3137 0 net=9209
rlabel metal2 1248 -3137 1248 -3137 0 net=10327
rlabel metal2 1402 -3137 1402 -3137 0 net=11389
rlabel metal2 1556 -3137 1556 -3137 0 net=14397
rlabel metal2 173 -3139 173 -3139 0 net=11735
rlabel metal2 1073 -3139 1073 -3139 0 net=10847
rlabel metal2 1318 -3139 1318 -3139 0 net=13231
rlabel metal2 1766 -3139 1766 -3139 0 net=13259
rlabel metal2 1906 -3139 1906 -3139 0 net=14171
rlabel metal2 205 -3141 205 -3141 0 net=13029
rlabel metal2 639 -3141 639 -3141 0 net=4010
rlabel metal2 912 -3141 912 -3141 0 net=10553
rlabel metal2 1409 -3141 1409 -3141 0 net=11369
rlabel metal2 1549 -3141 1549 -3141 0 net=12115
rlabel metal2 1661 -3141 1661 -3141 0 net=12269
rlabel metal2 219 -3143 219 -3143 0 net=1545
rlabel metal2 268 -3143 268 -3143 0 net=2025
rlabel metal2 394 -3143 394 -3143 0 net=5041
rlabel metal2 681 -3143 681 -3143 0 net=5369
rlabel metal2 765 -3143 765 -3143 0 net=8773
rlabel metal2 1073 -3143 1073 -3143 0 net=8941
rlabel metal2 1185 -3143 1185 -3143 0 net=10285
rlabel metal2 1367 -3143 1367 -3143 0 net=11449
rlabel metal2 1626 -3143 1626 -3143 0 net=14637
rlabel metal2 261 -3145 261 -3145 0 net=2031
rlabel metal2 1171 -3145 1171 -3145 0 net=11921
rlabel metal2 1472 -3145 1472 -3145 0 net=12713
rlabel metal2 1675 -3145 1675 -3145 0 net=14581
rlabel metal2 331 -3147 331 -3147 0 net=5909
rlabel metal2 597 -3147 597 -3147 0 net=4323
rlabel metal2 688 -3147 688 -3147 0 net=5657
rlabel metal2 800 -3147 800 -3147 0 net=5689
rlabel metal2 1017 -3147 1017 -3147 0 net=8797
rlabel metal2 1076 -3147 1076 -3147 0 net=445
rlabel metal2 1661 -3147 1661 -3147 0 net=14117
rlabel metal2 338 -3149 338 -3149 0 net=1755
rlabel metal2 394 -3149 394 -3149 0 net=3699
rlabel metal2 702 -3149 702 -3149 0 net=8723
rlabel metal2 1094 -3149 1094 -3149 0 net=9087
rlabel metal2 1227 -3149 1227 -3149 0 net=10241
rlabel metal2 1360 -3149 1360 -3149 0 net=11245
rlabel metal2 1535 -3149 1535 -3149 0 net=11637
rlabel metal2 338 -3151 338 -3151 0 net=2999
rlabel metal2 485 -3151 485 -3151 0 net=4623
rlabel metal2 576 -3151 576 -3151 0 net=3964
rlabel metal2 768 -3151 768 -3151 0 net=9058
rlabel metal2 1206 -3151 1206 -3151 0 net=10473
rlabel metal2 1220 -3151 1220 -3151 0 net=10219
rlabel metal2 1262 -3151 1262 -3151 0 net=9535
rlabel metal2 1486 -3151 1486 -3151 0 net=12579
rlabel metal2 37 -3153 37 -3153 0 net=6402
rlabel metal2 583 -3153 583 -3153 0 net=4465
rlabel metal2 1101 -3153 1101 -3153 0 net=8420
rlabel metal2 1241 -3153 1241 -3153 0 net=10591
rlabel metal2 1437 -3153 1437 -3153 0 net=12305
rlabel metal2 418 -3155 418 -3155 0 net=10339
rlabel metal2 485 -3155 485 -3155 0 net=5257
rlabel metal2 793 -3155 793 -3155 0 net=6191
rlabel metal2 985 -3155 985 -3155 0 net=13479
rlabel metal2 1542 -3155 1542 -3155 0 net=13755
rlabel metal2 443 -3157 443 -3157 0 net=2847
rlabel metal2 1262 -3157 1262 -3157 0 net=10965
rlabel metal2 1570 -3157 1570 -3157 0 net=11283
rlabel metal2 1738 -3157 1738 -3157 0 net=13047
rlabel metal2 506 -3159 506 -3159 0 net=3455
rlabel metal2 989 -3159 989 -3159 0 net=10439
rlabel metal2 1297 -3159 1297 -3159 0 net=10699
rlabel metal2 520 -3161 520 -3161 0 net=3529
rlabel metal2 1416 -3161 1416 -3161 0 net=11591
rlabel metal2 1591 -3161 1591 -3161 0 net=13615
rlabel metal2 1965 -3161 1965 -3161 0 net=14758
rlabel metal2 527 -3163 527 -3163 0 net=13572
rlabel metal2 905 -3163 905 -3163 0 net=6571
rlabel metal2 1003 -3163 1003 -3163 0 net=7729
rlabel metal2 1024 -3163 1024 -3163 0 net=8223
rlabel metal2 1101 -3163 1101 -3163 0 net=9133
rlabel metal2 1157 -3163 1157 -3163 0 net=9637
rlabel metal2 1325 -3163 1325 -3163 0 net=11035
rlabel metal2 1521 -3163 1521 -3163 0 net=10415
rlabel metal2 324 -3165 324 -3165 0 net=3011
rlabel metal2 1332 -3165 1332 -3165 0 net=10947
rlabel metal2 1493 -3165 1493 -3165 0 net=12749
rlabel metal2 324 -3167 324 -3167 0 net=2567
rlabel metal2 527 -3167 527 -3167 0 net=5753
rlabel metal2 786 -3167 786 -3167 0 net=6969
rlabel metal2 905 -3167 905 -3167 0 net=7549
rlabel metal2 1003 -3167 1003 -3167 0 net=8349
rlabel metal2 1143 -3167 1143 -3167 0 net=12445
rlabel metal2 1500 -3167 1500 -3167 0 net=11015
rlabel metal2 1577 -3167 1577 -3167 0 net=10572
rlabel metal2 387 -3169 387 -3169 0 net=3563
rlabel metal2 534 -3169 534 -3169 0 net=5495
rlabel metal2 800 -3169 800 -3169 0 net=1501
rlabel metal2 464 -3171 464 -3171 0 net=7774
rlabel metal2 814 -3171 814 -3171 0 net=11549
rlabel metal2 1500 -3171 1500 -3171 0 net=11677
rlabel metal2 1650 -3171 1650 -3171 0 net=922
rlabel metal2 163 -3173 163 -3173 0 net=6965
rlabel metal2 492 -3173 492 -3173 0 net=1957
rlabel metal2 1059 -3173 1059 -3173 0 net=8859
rlabel metal2 1356 -3173 1356 -3173 0 net=14327
rlabel metal2 1584 -3173 1584 -3173 0 net=13271
rlabel metal2 163 -3175 163 -3175 0 net=5021
rlabel metal2 933 -3175 933 -3175 0 net=7747
rlabel metal2 1066 -3175 1066 -3175 0 net=8539
rlabel metal2 1143 -3175 1143 -3175 0 net=9045
rlabel metal2 1514 -3175 1514 -3175 0 net=14025
rlabel metal2 1731 -3175 1731 -3175 0 net=13841
rlabel metal2 415 -3177 415 -3177 0 net=4364
rlabel metal2 513 -3177 513 -3177 0 net=5131
rlabel metal2 611 -3177 611 -3177 0 net=6779
rlabel metal2 940 -3177 940 -3177 0 net=9755
rlabel metal2 1150 -3177 1150 -3177 0 net=9545
rlabel metal2 1598 -3177 1598 -3177 0 net=14067
rlabel metal2 415 -3179 415 -3179 0 net=7473
rlabel metal2 954 -3179 954 -3179 0 net=9949
rlabel metal2 1283 -3179 1283 -3179 0 net=10273
rlabel metal2 1654 -3179 1654 -3179 0 net=10688
rlabel metal2 184 -3181 184 -3181 0 net=11093
rlabel metal2 1696 -3181 1696 -3181 0 net=14627
rlabel metal2 1969 -3181 1969 -3181 0 net=6039
rlabel metal2 590 -3183 590 -3183 0 net=4399
rlabel metal2 730 -3183 730 -3183 0 net=11166
rlabel metal2 1108 -3183 1108 -3183 0 net=10258
rlabel metal2 1745 -3183 1745 -3183 0 net=13561
rlabel metal2 1780 -3183 1780 -3183 0 net=13407
rlabel metal2 1983 -3183 1983 -3183 0 net=13465
rlabel metal2 82 -3185 82 -3185 0 net=10667
rlabel metal2 772 -3185 772 -3185 0 net=7235
rlabel metal2 1752 -3185 1752 -3185 0 net=13143
rlabel metal2 1773 -3185 1773 -3185 0 net=13369
rlabel metal2 562 -3187 562 -3187 0 net=1885
rlabel metal2 1752 -3187 1752 -3187 0 net=13739
rlabel metal2 499 -3189 499 -3189 0 net=3293
rlabel metal2 611 -3189 611 -3189 0 net=4704
rlabel metal2 674 -3189 674 -3189 0 net=3413
rlabel metal2 1773 -3189 1773 -3189 0 net=13897
rlabel metal2 499 -3191 499 -3191 0 net=5701
rlabel metal2 614 -3193 614 -3193 0 net=730
rlabel metal2 247 -3195 247 -3195 0 net=11194
rlabel metal2 618 -3195 618 -3195 0 net=4963
rlabel metal2 653 -3195 653 -3195 0 net=7129
rlabel metal2 240 -3197 240 -3197 0 net=2265
rlabel metal2 478 -3197 478 -3197 0 net=6115
rlabel metal2 660 -3197 660 -3197 0 net=8245
rlabel metal2 170 -3199 170 -3199 0 net=5463
rlabel metal2 408 -3199 408 -3199 0 net=4979
rlabel metal2 548 -3199 548 -3199 0 net=4193
rlabel metal2 667 -3199 667 -3199 0 net=7779
rlabel metal2 170 -3201 170 -3201 0 net=5246
rlabel metal2 779 -3201 779 -3201 0 net=7455
rlabel metal2 128 -3203 128 -3203 0 net=8107
rlabel metal2 849 -3203 849 -3203 0 net=6095
rlabel metal2 128 -3205 128 -3205 0 net=2501
rlabel metal2 408 -3205 408 -3205 0 net=2587
rlabel metal2 548 -3205 548 -3205 0 net=10121
rlabel metal2 849 -3205 849 -3205 0 net=9449
rlabel metal2 149 -3207 149 -3207 0 net=9215
rlabel metal2 947 -3207 947 -3207 0 net=7677
rlabel metal2 1038 -3207 1038 -3207 0 net=8259
rlabel metal2 996 -3209 996 -3209 0 net=8025
rlabel metal2 1087 -3209 1087 -3209 0 net=9387
rlabel metal2 1010 -3211 1010 -3211 0 net=5089
rlabel metal2 1255 -3213 1255 -3213 0 net=10738
rlabel metal2 1164 -3215 1164 -3215 0 net=11613
rlabel metal2 1164 -3217 1164 -3217 0 net=13788
rlabel metal2 1430 -3219 1430 -3219 0 net=10645
rlabel metal2 1430 -3221 1430 -3221 0 net=11909
rlabel metal2 1619 -3223 1619 -3223 0 net=14451
rlabel metal2 93 -3234 93 -3234 0 net=8398
rlabel metal2 184 -3234 184 -3234 0 net=11209
rlabel metal2 541 -3234 541 -3234 0 net=4625
rlabel metal2 541 -3234 541 -3234 0 net=4625
rlabel metal2 548 -3234 548 -3234 0 net=10122
rlabel metal2 642 -3234 642 -3234 0 net=7236
rlabel metal2 800 -3234 800 -3234 0 net=9536
rlabel metal2 1563 -3234 1563 -3234 0 net=10802
rlabel metal2 1668 -3234 1668 -3234 0 net=13147
rlabel metal2 1738 -3234 1738 -3234 0 net=10416
rlabel metal2 1969 -3234 1969 -3234 0 net=6041
rlabel metal2 1969 -3234 1969 -3234 0 net=6041
rlabel metal2 2018 -3234 2018 -3234 0 net=13681
rlabel metal2 2032 -3234 2032 -3234 0 net=3381
rlabel metal2 107 -3236 107 -3236 0 net=3944
rlabel metal2 688 -3236 688 -3236 0 net=5658
rlabel metal2 1213 -3236 1213 -3236 0 net=14068
rlabel metal2 1640 -3236 1640 -3236 0 net=13562
rlabel metal2 1766 -3236 1766 -3236 0 net=12271
rlabel metal2 1808 -3236 1808 -3236 0 net=13408
rlabel metal2 1857 -3236 1857 -3236 0 net=13923
rlabel metal2 1857 -3236 1857 -3236 0 net=13923
rlabel metal2 1871 -3236 1871 -3236 0 net=14265
rlabel metal2 1962 -3236 1962 -3236 0 net=13466
rlabel metal2 121 -3238 121 -3238 0 net=2138
rlabel metal2 208 -3238 208 -3238 0 net=3528
rlabel metal2 233 -3238 233 -3238 0 net=5450
rlabel metal2 275 -3238 275 -3238 0 net=10544
rlabel metal2 800 -3238 800 -3238 0 net=7475
rlabel metal2 929 -3238 929 -3238 0 net=14154
rlabel metal2 1689 -3238 1689 -3238 0 net=1503
rlabel metal2 1815 -3238 1815 -3238 0 net=13049
rlabel metal2 1878 -3238 1878 -3238 0 net=14019
rlabel metal2 1878 -3238 1878 -3238 0 net=14019
rlabel metal2 1962 -3238 1962 -3238 0 net=14691
rlabel metal2 100 -3240 100 -3240 0 net=6050
rlabel metal2 247 -3240 247 -3240 0 net=2267
rlabel metal2 282 -3240 282 -3240 0 net=4380
rlabel metal2 464 -3240 464 -3240 0 net=6966
rlabel metal2 873 -3240 873 -3240 0 net=11734
rlabel metal2 1528 -3240 1528 -3240 0 net=10646
rlabel metal2 1703 -3240 1703 -3240 0 net=6955
rlabel metal2 1815 -3240 1815 -3240 0 net=13565
rlabel metal2 128 -3242 128 -3242 0 net=2502
rlabel metal2 191 -3242 191 -3242 0 net=13272
rlabel metal2 1598 -3242 1598 -3242 0 net=13607
rlabel metal2 1717 -3242 1717 -3242 0 net=11285
rlabel metal2 1745 -3242 1745 -3242 0 net=13899
rlabel metal2 1780 -3242 1780 -3242 0 net=13371
rlabel metal2 1780 -3242 1780 -3242 0 net=13371
rlabel metal2 1822 -3242 1822 -3242 0 net=13261
rlabel metal2 135 -3244 135 -3244 0 net=2080
rlabel metal2 751 -3244 751 -3244 0 net=8108
rlabel metal2 957 -3244 957 -3244 0 net=8026
rlabel metal2 1104 -3244 1104 -3244 0 net=10220
rlabel metal2 1237 -3244 1237 -3244 0 net=14452
rlabel metal2 1717 -3244 1717 -3244 0 net=13843
rlabel metal2 1759 -3244 1759 -3244 0 net=13145
rlabel metal2 156 -3246 156 -3246 0 net=7467
rlabel metal2 191 -3246 191 -3246 0 net=6013
rlabel metal2 1731 -3246 1731 -3246 0 net=13741
rlabel metal2 205 -3248 205 -3248 0 net=9457
rlabel metal2 215 -3248 215 -3248 0 net=277
rlabel metal2 1108 -3248 1108 -3248 0 net=1
rlabel metal2 1724 -3248 1724 -3248 0 net=11983
rlabel metal2 219 -3250 219 -3250 0 net=1546
rlabel metal2 814 -3250 814 -3250 0 net=5091
rlabel metal2 1108 -3250 1108 -3250 0 net=8661
rlabel metal2 1216 -3250 1216 -3250 0 net=11370
rlabel metal2 1465 -3250 1465 -3250 0 net=2469
rlabel metal2 219 -3252 219 -3252 0 net=2155
rlabel metal2 464 -3252 464 -3252 0 net=3457
rlabel metal2 513 -3252 513 -3252 0 net=5132
rlabel metal2 632 -3252 632 -3252 0 net=13031
rlabel metal2 1216 -3252 1216 -3252 0 net=10952
rlabel metal2 1353 -3252 1353 -3252 0 net=13616
rlabel metal2 1654 -3252 1654 -3252 0 net=14629
rlabel metal2 240 -3254 240 -3254 0 net=5465
rlabel metal2 569 -3254 569 -3254 0 net=4291
rlabel metal2 569 -3254 569 -3254 0 net=4291
rlabel metal2 576 -3254 576 -3254 0 net=1318
rlabel metal2 240 -3256 240 -3256 0 net=5043
rlabel metal2 653 -3256 653 -3256 0 net=6117
rlabel metal2 716 -3256 716 -3256 0 net=10948
rlabel metal2 1346 -3256 1346 -3256 0 net=12581
rlabel metal2 1549 -3256 1549 -3256 0 net=12117
rlabel metal2 247 -3258 247 -3258 0 net=2033
rlabel metal2 282 -3258 282 -3258 0 net=8247
rlabel metal2 674 -3258 674 -3258 0 net=8725
rlabel metal2 716 -3258 716 -3258 0 net=7587
rlabel metal2 1080 -3258 1080 -3258 0 net=6097
rlabel metal2 1374 -3258 1374 -3258 0 net=11551
rlabel metal2 1472 -3258 1472 -3258 0 net=12715
rlabel metal2 1563 -3258 1563 -3258 0 net=14119
rlabel metal2 254 -3260 254 -3260 0 net=2681
rlabel metal2 303 -3260 303 -3260 0 net=1649
rlabel metal2 303 -3260 303 -3260 0 net=1649
rlabel metal2 331 -3260 331 -3260 0 net=5911
rlabel metal2 751 -3260 751 -3260 0 net=6413
rlabel metal2 856 -3260 856 -3260 0 net=5691
rlabel metal2 985 -3260 985 -3260 0 net=9764
rlabel metal2 1290 -3260 1290 -3260 0 net=3012
rlabel metal2 1486 -3260 1486 -3260 0 net=3679
rlabel metal2 1661 -3260 1661 -3260 0 net=14583
rlabel metal2 268 -3262 268 -3262 0 net=2027
rlabel metal2 338 -3262 338 -3262 0 net=3000
rlabel metal2 772 -3262 772 -3262 0 net=6193
rlabel metal2 807 -3262 807 -3262 0 net=7679
rlabel metal2 957 -3262 957 -3262 0 net=10803
rlabel metal2 1167 -3262 1167 -3262 0 net=4843
rlabel metal2 268 -3264 268 -3264 0 net=1967
rlabel metal2 338 -3264 338 -3264 0 net=4903
rlabel metal2 653 -3264 653 -3264 0 net=1887
rlabel metal2 702 -3264 702 -3264 0 net=4409
rlabel metal2 1269 -3264 1269 -3264 0 net=14208
rlabel metal2 289 -3266 289 -3266 0 net=1757
rlabel metal2 352 -3266 352 -3266 0 net=6508
rlabel metal2 485 -3266 485 -3266 0 net=5259
rlabel metal2 562 -3266 562 -3266 0 net=3295
rlabel metal2 863 -3266 863 -3266 0 net=7143
rlabel metal2 898 -3266 898 -3266 0 net=9089
rlabel metal2 1115 -3266 1115 -3266 0 net=5564
rlabel metal2 1237 -3266 1237 -3266 0 net=1127
rlabel metal2 345 -3268 345 -3268 0 net=4195
rlabel metal2 660 -3268 660 -3268 0 net=7781
rlabel metal2 695 -3268 695 -3268 0 net=10669
rlabel metal2 793 -3268 793 -3268 0 net=8775
rlabel metal2 1115 -3268 1115 -3268 0 net=10441
rlabel metal2 1220 -3268 1220 -3268 0 net=12751
rlabel metal2 352 -3270 352 -3270 0 net=2849
rlabel metal2 485 -3270 485 -3270 0 net=6781
rlabel metal2 912 -3270 912 -3270 0 net=10555
rlabel metal2 1031 -3270 1031 -3270 0 net=9547
rlabel metal2 1171 -3270 1171 -3270 0 net=11923
rlabel metal2 1290 -3270 1290 -3270 0 net=12937
rlabel metal2 1332 -3270 1332 -3270 0 net=11095
rlabel metal2 1374 -3270 1374 -3270 0 net=14027
rlabel metal2 229 -3272 229 -3272 0 net=3855
rlabel metal2 495 -3272 495 -3272 0 net=37
rlabel metal2 583 -3272 583 -3272 0 net=4466
rlabel metal2 646 -3272 646 -3272 0 net=5371
rlabel metal2 786 -3272 786 -3272 0 net=8861
rlabel metal2 1066 -3272 1066 -3272 0 net=8541
rlabel metal2 1500 -3272 1500 -3272 0 net=11679
rlabel metal2 359 -3274 359 -3274 0 net=2302
rlabel metal2 499 -3274 499 -3274 0 net=5702
rlabel metal2 912 -3274 912 -3274 0 net=7749
rlabel metal2 947 -3274 947 -3274 0 net=8351
rlabel metal2 1059 -3274 1059 -3274 0 net=9951
rlabel metal2 1192 -3274 1192 -3274 0 net=10967
rlabel metal2 1283 -3274 1283 -3274 0 net=10275
rlabel metal2 177 -3276 177 -3276 0 net=6031
rlabel metal2 527 -3276 527 -3276 0 net=5755
rlabel metal2 709 -3276 709 -3276 0 net=9441
rlabel metal2 1066 -3276 1066 -3276 0 net=10242
rlabel metal2 1262 -3276 1262 -3276 0 net=14399
rlabel metal2 177 -3278 177 -3278 0 net=2317
rlabel metal2 359 -3278 359 -3278 0 net=2221
rlabel metal2 527 -3278 527 -3278 0 net=2059
rlabel metal2 919 -3278 919 -3278 0 net=8063
rlabel metal2 968 -3278 968 -3278 0 net=9211
rlabel metal2 1150 -3278 1150 -3278 0 net=10701
rlabel metal2 1311 -3278 1311 -3278 0 net=13233
rlabel metal2 1409 -3278 1409 -3278 0 net=2775
rlabel metal2 163 -3280 163 -3280 0 net=5023
rlabel metal2 366 -3280 366 -3280 0 net=2763
rlabel metal2 555 -3280 555 -3280 0 net=4802
rlabel metal2 1458 -3280 1458 -3280 0 net=13757
rlabel metal2 1853 -3280 1853 -3280 0 net=14006
rlabel metal2 142 -3282 142 -3282 0 net=13177
rlabel metal2 324 -3282 324 -3282 0 net=2569
rlabel metal2 373 -3282 373 -3282 0 net=3227
rlabel metal2 478 -3282 478 -3282 0 net=4981
rlabel metal2 562 -3282 562 -3282 0 net=4325
rlabel metal2 604 -3282 604 -3282 0 net=8035
rlabel metal2 919 -3282 919 -3282 0 net=9299
rlabel metal2 968 -3282 968 -3282 0 net=6900
rlabel metal2 1157 -3282 1157 -3282 0 net=9639
rlabel metal2 1283 -3282 1283 -3282 0 net=12295
rlabel metal2 1535 -3282 1535 -3282 0 net=11639
rlabel metal2 1864 -3282 1864 -3282 0 net=14711
rlabel metal2 117 -3284 117 -3284 0 net=8301
rlabel metal2 310 -3284 310 -3284 0 net=4176
rlabel metal2 667 -3284 667 -3284 0 net=7457
rlabel metal2 1122 -3284 1122 -3284 0 net=10475
rlabel metal2 1297 -3284 1297 -3284 0 net=11451
rlabel metal2 1892 -3284 1892 -3284 0 net=14173
rlabel metal2 310 -3286 310 -3286 0 net=1917
rlabel metal2 324 -3286 324 -3286 0 net=2751
rlabel metal2 576 -3286 576 -3286 0 net=5795
rlabel metal2 1143 -3286 1143 -3286 0 net=9047
rlabel metal2 1171 -3286 1171 -3286 0 net=12471
rlabel metal2 1906 -3286 1906 -3286 0 net=1859
rlabel metal2 317 -3288 317 -3288 0 net=5017
rlabel metal2 709 -3288 709 -3288 0 net=6795
rlabel metal2 940 -3288 940 -3288 0 net=8225
rlabel metal2 1178 -3288 1178 -3288 0 net=11593
rlabel metal2 373 -3290 373 -3290 0 net=10341
rlabel metal2 583 -3290 583 -3290 0 net=8457
rlabel metal2 625 -3290 625 -3290 0 net=3583
rlabel metal2 1206 -3290 1206 -3290 0 net=12307
rlabel metal2 149 -3292 149 -3292 0 net=9217
rlabel metal2 737 -3292 737 -3292 0 net=7731
rlabel metal2 1024 -3292 1024 -3292 0 net=8799
rlabel metal2 1318 -3292 1318 -3292 0 net=11911
rlabel metal2 383 -3294 383 -3294 0 net=12509
rlabel metal2 961 -3294 961 -3294 0 net=8455
rlabel metal2 1402 -3294 1402 -3294 0 net=11391
rlabel metal2 387 -3296 387 -3296 0 net=3565
rlabel metal2 590 -3296 590 -3296 0 net=4401
rlabel metal2 765 -3296 765 -3296 0 net=4063
rlabel metal2 1038 -3296 1038 -3296 0 net=8261
rlabel metal2 1136 -3296 1136 -3296 0 net=9757
rlabel metal2 387 -3298 387 -3298 0 net=3843
rlabel metal2 590 -3298 590 -3298 0 net=9389
rlabel metal2 1136 -3298 1136 -3298 0 net=10613
rlabel metal2 1325 -3298 1325 -3298 0 net=11037
rlabel metal2 394 -3300 394 -3300 0 net=3701
rlabel metal2 765 -3300 765 -3300 0 net=7551
rlabel metal2 961 -3300 961 -3300 0 net=6573
rlabel metal2 1038 -3300 1038 -3300 0 net=3985
rlabel metal2 1087 -3300 1087 -3300 0 net=10287
rlabel metal2 1199 -3300 1199 -3300 0 net=11247
rlabel metal2 1367 -3300 1367 -3300 0 net=11016
rlabel metal2 394 -3302 394 -3302 0 net=2589
rlabel metal2 429 -3302 429 -3302 0 net=5497
rlabel metal2 723 -3302 723 -3302 0 net=3415
rlabel metal2 1325 -3302 1325 -3302 0 net=14329
rlabel metal2 380 -3304 380 -3304 0 net=6513
rlabel metal2 450 -3304 450 -3304 0 net=4965
rlabel metal2 779 -3304 779 -3304 0 net=5992
rlabel metal2 1451 -3304 1451 -3304 0 net=11061
rlabel metal2 380 -3306 380 -3306 0 net=7563
rlabel metal2 534 -3306 534 -3306 0 net=1293
rlabel metal2 401 -3308 401 -3308 0 net=9803
rlabel metal2 821 -3308 821 -3308 0 net=6241
rlabel metal2 884 -3308 884 -3308 0 net=6971
rlabel metal2 1451 -3308 1451 -3308 0 net=13481
rlabel metal2 296 -3310 296 -3310 0 net=2717
rlabel metal2 404 -3310 404 -3310 0 net=3108
rlabel metal2 471 -3310 471 -3310 0 net=1959
rlabel metal2 978 -3310 978 -3310 0 net=10513
rlabel metal2 1248 -3310 1248 -3310 0 net=10329
rlabel metal2 1423 -3310 1423 -3310 0 net=11615
rlabel metal2 296 -3312 296 -3312 0 net=12099
rlabel metal2 821 -3312 821 -3312 0 net=7131
rlabel metal2 849 -3312 849 -3312 0 net=9451
rlabel metal2 905 -3312 905 -3312 0 net=6901
rlabel metal2 1248 -3312 1248 -3312 0 net=12447
rlabel metal2 457 -3314 457 -3314 0 net=3531
rlabel metal2 842 -3314 842 -3314 0 net=7199
rlabel metal2 989 -3314 989 -3314 0 net=14638
rlabel metal2 520 -3316 520 -3316 0 net=3349
rlabel metal2 877 -3316 877 -3316 0 net=7207
rlabel metal2 1304 -3316 1304 -3316 0 net=10849
rlabel metal2 1479 -3316 1479 -3316 0 net=6625
rlabel metal2 758 -3318 758 -3318 0 net=6873
rlabel metal2 1304 -3318 1304 -3318 0 net=12981
rlabel metal2 1626 -3318 1626 -3318 0 net=7163
rlabel metal2 828 -3320 828 -3320 0 net=9067
rlabel metal2 1073 -3320 1073 -3320 0 net=8943
rlabel metal2 828 -3322 828 -3322 0 net=8279
rlabel metal2 1073 -3322 1073 -3322 0 net=10593
rlabel metal2 254 -3324 254 -3324 0 net=319
rlabel metal2 1045 -3324 1045 -3324 0 net=11737
rlabel metal2 1045 -3326 1045 -3326 0 net=9135
rlabel metal2 142 -3337 142 -3337 0 net=8302
rlabel metal2 177 -3337 177 -3337 0 net=2318
rlabel metal2 257 -3337 257 -3337 0 net=10342
rlabel metal2 394 -3337 394 -3337 0 net=2590
rlabel metal2 541 -3337 541 -3337 0 net=4627
rlabel metal2 590 -3337 590 -3337 0 net=9390
rlabel metal2 814 -3337 814 -3337 0 net=5092
rlabel metal2 1160 -3337 1160 -3337 0 net=9640
rlabel metal2 1234 -3337 1234 -3337 0 net=13482
rlabel metal2 1500 -3337 1500 -3337 0 net=10277
rlabel metal2 1500 -3337 1500 -3337 0 net=10277
rlabel metal2 1521 -3337 1521 -3337 0 net=11062
rlabel metal2 1591 -3337 1591 -3337 0 net=12119
rlabel metal2 1647 -3337 1647 -3337 0 net=14585
rlabel metal2 1717 -3337 1717 -3337 0 net=13844
rlabel metal2 1731 -3337 1731 -3337 0 net=13743
rlabel metal2 1731 -3337 1731 -3337 0 net=13743
rlabel metal2 1738 -3337 1738 -3337 0 net=11287
rlabel metal2 1738 -3337 1738 -3337 0 net=11287
rlabel metal2 1752 -3337 1752 -3337 0 net=11985
rlabel metal2 1766 -3337 1766 -3337 0 net=13146
rlabel metal2 1780 -3337 1780 -3337 0 net=13373
rlabel metal2 1780 -3337 1780 -3337 0 net=13373
rlabel metal2 1787 -3337 1787 -3337 0 net=12272
rlabel metal2 1829 -3337 1829 -3337 0 net=13051
rlabel metal2 1885 -3337 1885 -3337 0 net=1860
rlabel metal2 1955 -3337 1955 -3337 0 net=14693
rlabel metal2 2025 -3337 2025 -3337 0 net=13683
rlabel metal2 163 -3339 163 -3339 0 net=13178
rlabel metal2 415 -3339 415 -3339 0 net=6782
rlabel metal2 488 -3339 488 -3339 0 net=5466
rlabel metal2 513 -3339 513 -3339 0 net=5260
rlabel metal2 1034 -3339 1034 -3339 0 net=12752
rlabel metal2 1234 -3339 1234 -3339 0 net=12297
rlabel metal2 1339 -3339 1339 -3339 0 net=13758
rlabel metal2 1521 -3339 1521 -3339 0 net=12717
rlabel metal2 1549 -3339 1549 -3339 0 net=7164
rlabel metal2 1724 -3339 1724 -3339 0 net=13901
rlabel metal2 1787 -3339 1787 -3339 0 net=6315
rlabel metal2 1888 -3339 1888 -3339 0 net=14174
rlabel metal2 1962 -3339 1962 -3339 0 net=6043
rlabel metal2 2025 -3339 2025 -3339 0 net=3383
rlabel metal2 170 -3341 170 -3341 0 net=7468
rlabel metal2 212 -3341 212 -3341 0 net=6514
rlabel metal2 429 -3341 429 -3341 0 net=5498
rlabel metal2 968 -3341 968 -3341 0 net=11096
rlabel metal2 1367 -3341 1367 -3341 0 net=8543
rlabel metal2 1528 -3341 1528 -3341 0 net=14121
rlabel metal2 1605 -3341 1605 -3341 0 net=14630
rlabel metal2 1794 -3341 1794 -3341 0 net=1505
rlabel metal2 1836 -3341 1836 -3341 0 net=13263
rlabel metal2 1850 -3341 1850 -3341 0 net=13925
rlabel metal2 215 -3343 215 -3343 0 net=1459
rlabel metal2 821 -3343 821 -3343 0 net=7132
rlabel metal2 968 -3343 968 -3343 0 net=9443
rlabel metal2 1031 -3343 1031 -3343 0 net=9549
rlabel metal2 1237 -3343 1237 -3343 0 net=11452
rlabel metal2 1332 -3343 1332 -3343 0 net=14029
rlabel metal2 1381 -3343 1381 -3343 0 net=11552
rlabel metal2 1451 -3343 1451 -3343 0 net=3681
rlabel metal2 1552 -3343 1552 -3343 0 net=13608
rlabel metal2 1608 -3343 1608 -3343 0 net=13148
rlabel metal2 1801 -3343 1801 -3343 0 net=6957
rlabel metal2 1857 -3343 1857 -3343 0 net=14267
rlabel metal2 240 -3345 240 -3345 0 net=5045
rlabel metal2 541 -3345 541 -3345 0 net=5797
rlabel metal2 597 -3345 597 -3345 0 net=375
rlabel metal2 1097 -3345 1097 -3345 0 net=13234
rlabel metal2 1374 -3345 1374 -3345 0 net=10621
rlabel metal2 1556 -3345 1556 -3345 0 net=11640
rlabel metal2 1654 -3345 1654 -3345 0 net=10739
rlabel metal2 1864 -3345 1864 -3345 0 net=14713
rlabel metal2 275 -3347 275 -3347 0 net=2269
rlabel metal2 422 -3347 422 -3347 0 net=2765
rlabel metal2 474 -3347 474 -3347 0 net=66
rlabel metal2 1384 -3347 1384 -3347 0 net=10850
rlabel metal2 1801 -3347 1801 -3347 0 net=13567
rlabel metal2 1864 -3347 1864 -3347 0 net=14021
rlabel metal2 2028 -3347 2028 -3347 0 net=1
rlabel metal2 205 -3349 205 -3349 0 net=9459
rlabel metal2 548 -3349 548 -3349 0 net=3702
rlabel metal2 1066 -3349 1066 -3349 0 net=11038
rlabel metal2 282 -3351 282 -3351 0 net=8248
rlabel metal2 877 -3351 877 -3351 0 net=7209
rlabel metal2 1080 -3351 1080 -3351 0 net=10614
rlabel metal2 1199 -3351 1199 -3351 0 net=11249
rlabel metal2 1269 -3351 1269 -3351 0 net=6098
rlabel metal2 1388 -3351 1388 -3351 0 net=8456
rlabel metal2 296 -3353 296 -3353 0 net=12100
rlabel metal2 492 -3353 492 -3353 0 net=3567
rlabel metal2 555 -3353 555 -3353 0 net=4983
rlabel metal2 597 -3353 597 -3353 0 net=5373
rlabel metal2 653 -3353 653 -3353 0 net=1889
rlabel metal2 891 -3353 891 -3353 0 net=9068
rlabel metal2 961 -3353 961 -3353 0 net=6575
rlabel metal2 1101 -3353 1101 -3353 0 net=11595
rlabel metal2 1199 -3353 1199 -3353 0 net=14331
rlabel metal2 1416 -3353 1416 -3353 0 net=11392
rlabel metal2 268 -3355 268 -3355 0 net=1969
rlabel metal2 317 -3355 317 -3355 0 net=5019
rlabel metal2 450 -3355 450 -3355 0 net=4967
rlabel metal2 534 -3355 534 -3355 0 net=11625
rlabel metal2 674 -3355 674 -3355 0 net=8726
rlabel metal2 1045 -3355 1045 -3355 0 net=9137
rlabel metal2 1213 -3355 1213 -3355 0 net=9758
rlabel metal2 359 -3357 359 -3357 0 net=2223
rlabel metal2 534 -3357 534 -3357 0 net=8459
rlabel metal2 618 -3357 618 -3357 0 net=9805
rlabel metal2 660 -3357 660 -3357 0 net=7783
rlabel metal2 681 -3357 681 -3357 0 net=5756
rlabel metal2 1157 -3357 1157 -3357 0 net=9049
rlabel metal2 1269 -3357 1269 -3357 0 net=4845
rlabel metal2 303 -3359 303 -3359 0 net=1651
rlabel metal2 366 -3359 366 -3359 0 net=2571
rlabel metal2 478 -3359 478 -3359 0 net=7564
rlabel metal2 562 -3359 562 -3359 0 net=4327
rlabel metal2 716 -3359 716 -3359 0 net=7589
rlabel metal2 716 -3359 716 -3359 0 net=7589
rlabel metal2 723 -3359 723 -3359 0 net=8944
rlabel metal2 1472 -3359 1472 -3359 0 net=11681
rlabel metal2 331 -3361 331 -3361 0 net=2029
rlabel metal2 562 -3361 562 -3361 0 net=5157
rlabel metal2 730 -3361 730 -3361 0 net=1345
rlabel metal2 198 -3363 198 -3363 0 net=5025
rlabel metal2 345 -3363 345 -3363 0 net=4197
rlabel metal2 723 -3363 723 -3363 0 net=6874
rlabel metal2 772 -3363 772 -3363 0 net=6195
rlabel metal2 821 -3363 821 -3363 0 net=9953
rlabel metal2 1272 -3363 1272 -3363 0 net=14057
rlabel metal2 1290 -3363 1290 -3363 0 net=12939
rlabel metal2 289 -3365 289 -3365 0 net=1759
rlabel metal2 387 -3365 387 -3365 0 net=3845
rlabel metal2 583 -3365 583 -3365 0 net=7459
rlabel metal2 737 -3365 737 -3365 0 net=7733
rlabel metal2 978 -3365 978 -3365 0 net=8800
rlabel metal2 1045 -3365 1045 -3365 0 net=10515
rlabel metal2 1255 -3365 1255 -3365 0 net=11925
rlabel metal2 219 -3367 219 -3367 0 net=2156
rlabel metal2 443 -3367 443 -3367 0 net=3857
rlabel metal2 751 -3367 751 -3367 0 net=6414
rlabel metal2 1192 -3367 1192 -3367 0 net=10969
rlabel metal2 352 -3369 352 -3369 0 net=2850
rlabel metal2 772 -3369 772 -3369 0 net=7477
rlabel metal2 835 -3369 835 -3369 0 net=6242
rlabel metal2 852 -3369 852 -3369 0 net=10556
rlabel metal2 1024 -3369 1024 -3369 0 net=3986
rlabel metal2 1059 -3369 1059 -3369 0 net=10595
rlabel metal2 1094 -3369 1094 -3369 0 net=11739
rlabel metal2 401 -3371 401 -3371 0 net=2719
rlabel metal2 471 -3371 471 -3371 0 net=1961
rlabel metal2 779 -3371 779 -3371 0 net=8663
rlabel metal2 982 -3371 982 -3371 0 net=5692
rlabel metal2 1192 -3371 1192 -3371 0 net=2471
rlabel metal2 401 -3373 401 -3373 0 net=10311
rlabel metal2 793 -3373 793 -3373 0 net=8777
rlabel metal2 842 -3373 842 -3373 0 net=7200
rlabel metal2 989 -3373 989 -3373 0 net=6972
rlabel metal2 1465 -3373 1465 -3373 0 net=11617
rlabel metal2 600 -3375 600 -3375 0 net=7041
rlabel metal2 1241 -3375 1241 -3375 0 net=12983
rlabel metal2 1346 -3375 1346 -3375 0 net=12583
rlabel metal2 604 -3377 604 -3377 0 net=8037
rlabel metal2 800 -3377 800 -3377 0 net=1215
rlabel metal2 604 -3379 604 -3379 0 net=9219
rlabel metal2 618 -3379 618 -3379 0 net=6797
rlabel metal2 842 -3379 842 -3379 0 net=12308
rlabel metal2 1318 -3379 1318 -3379 0 net=11913
rlabel metal2 520 -3381 520 -3381 0 net=3351
rlabel metal2 849 -3381 849 -3381 0 net=10703
rlabel metal2 1185 -3381 1185 -3381 0 net=3416
rlabel metal2 418 -3383 418 -3383 0 net=13505
rlabel metal2 527 -3383 527 -3383 0 net=2061
rlabel metal2 625 -3383 625 -3383 0 net=3585
rlabel metal2 688 -3383 688 -3383 0 net=6119
rlabel metal2 856 -3383 856 -3383 0 net=3297
rlabel metal2 989 -3383 989 -3383 0 net=12448
rlabel metal2 457 -3385 457 -3385 0 net=3533
rlabel metal2 688 -3385 688 -3385 0 net=8863
rlabel metal2 870 -3385 870 -3385 0 net=7145
rlabel metal2 1108 -3385 1108 -3385 0 net=8662
rlabel metal2 1209 -3385 1209 -3385 0 net=10605
rlabel metal2 310 -3387 310 -3387 0 net=1919
rlabel metal2 527 -3387 527 -3387 0 net=4293
rlabel metal2 786 -3387 786 -3387 0 net=9453
rlabel metal2 891 -3387 891 -3387 0 net=10477
rlabel metal2 1185 -3387 1185 -3387 0 net=6627
rlabel metal2 184 -3389 184 -3389 0 net=11211
rlabel metal2 807 -3389 807 -3389 0 net=7681
rlabel metal2 1122 -3389 1122 -3389 0 net=12605
rlabel metal2 261 -3391 261 -3391 0 net=2683
rlabel metal2 695 -3391 695 -3391 0 net=10671
rlabel metal2 863 -3391 863 -3391 0 net=12511
rlabel metal2 898 -3391 898 -3391 0 net=9091
rlabel metal2 324 -3393 324 -3393 0 net=2753
rlabel metal2 744 -3393 744 -3393 0 net=5913
rlabel metal2 870 -3393 870 -3393 0 net=6903
rlabel metal2 919 -3393 919 -3393 0 net=9301
rlabel metal2 702 -3395 702 -3395 0 net=4411
rlabel metal2 901 -3395 901 -3395 0 net=10330
rlabel metal2 464 -3397 464 -3397 0 net=3459
rlabel metal2 905 -3397 905 -3397 0 net=10443
rlabel metal2 436 -3399 436 -3399 0 net=3229
rlabel metal2 912 -3399 912 -3399 0 net=7750
rlabel metal2 926 -3399 926 -3399 0 net=13033
rlabel metal2 380 -3401 380 -3401 0 net=666
rlabel metal2 765 -3401 765 -3401 0 net=7553
rlabel metal2 940 -3401 940 -3401 0 net=8227
rlabel metal2 247 -3403 247 -3403 0 net=2035
rlabel metal2 632 -3403 632 -3403 0 net=4403
rlabel metal2 940 -3403 940 -3403 0 net=3041
rlabel metal2 499 -3405 499 -3405 0 net=6033
rlabel metal2 947 -3405 947 -3405 0 net=8353
rlabel metal2 338 -3407 338 -3407 0 net=4905
rlabel metal2 828 -3407 828 -3407 0 net=8281
rlabel metal2 954 -3407 954 -3407 0 net=9213
rlabel metal2 1052 -3407 1052 -3407 0 net=8263
rlabel metal2 191 -3409 191 -3409 0 net=6015
rlabel metal2 828 -3409 828 -3409 0 net=8065
rlabel metal2 996 -3409 996 -3409 0 net=12473
rlabel metal2 933 -3411 933 -3411 0 net=4064
rlabel metal2 1052 -3411 1052 -3411 0 net=10289
rlabel metal2 1171 -3411 1171 -3411 0 net=14401
rlabel metal2 971 -3413 971 -3413 0 net=7341
rlabel metal2 1087 -3413 1087 -3413 0 net=10805
rlabel metal2 1262 -3413 1262 -3413 0 net=2777
rlabel metal2 173 -3424 173 -3424 0 net=612
rlabel metal2 296 -3424 296 -3424 0 net=1970
rlabel metal2 338 -3424 338 -3424 0 net=6016
rlabel metal2 478 -3424 478 -3424 0 net=2030
rlabel metal2 621 -3424 621 -3424 0 net=6034
rlabel metal2 639 -3424 639 -3424 0 net=9806
rlabel metal2 726 -3424 726 -3424 0 net=3042
rlabel metal2 961 -3424 961 -3424 0 net=7734
rlabel metal2 1213 -3424 1213 -3424 0 net=9050
rlabel metal2 1290 -3424 1290 -3424 0 net=11927
rlabel metal2 1290 -3424 1290 -3424 0 net=11927
rlabel metal2 1297 -3424 1297 -3424 0 net=12940
rlabel metal2 1311 -3424 1311 -3424 0 net=14031
rlabel metal2 1346 -3424 1346 -3424 0 net=11914
rlabel metal2 1437 -3424 1437 -3424 0 net=3683
rlabel metal2 1458 -3424 1458 -3424 0 net=10623
rlabel metal2 1500 -3424 1500 -3424 0 net=10279
rlabel metal2 1500 -3424 1500 -3424 0 net=10279
rlabel metal2 1514 -3424 1514 -3424 0 net=14123
rlabel metal2 1584 -3424 1584 -3424 0 net=326
rlabel metal2 1822 -3424 1822 -3424 0 net=1506
rlabel metal2 1955 -3424 1955 -3424 0 net=14695
rlabel metal2 1955 -3424 1955 -3424 0 net=14695
rlabel metal2 1962 -3424 1962 -3424 0 net=6045
rlabel metal2 1962 -3424 1962 -3424 0 net=6045
rlabel metal2 2025 -3424 2025 -3424 0 net=3385
rlabel metal2 2025 -3424 2025 -3424 0 net=3385
rlabel metal2 2032 -3424 2032 -3424 0 net=13685
rlabel metal2 2032 -3424 2032 -3424 0 net=13685
rlabel metal2 170 -3426 170 -3426 0 net=1383
rlabel metal2 310 -3426 310 -3426 0 net=2685
rlabel metal2 345 -3426 345 -3426 0 net=1760
rlabel metal2 394 -3426 394 -3426 0 net=2572
rlabel metal2 404 -3426 404 -3426 0 net=4239
rlabel metal2 429 -3426 429 -3426 0 net=2766
rlabel metal2 492 -3426 492 -3426 0 net=4968
rlabel metal2 646 -3426 646 -3426 0 net=11627
rlabel metal2 758 -3426 758 -3426 0 net=8039
rlabel metal2 807 -3426 807 -3426 0 net=10672
rlabel metal2 884 -3426 884 -3426 0 net=12512
rlabel metal2 975 -3426 975 -3426 0 net=7147
rlabel metal2 1038 -3426 1038 -3426 0 net=9093
rlabel metal2 1038 -3426 1038 -3426 0 net=9093
rlabel metal2 1066 -3426 1066 -3426 0 net=14332
rlabel metal2 1206 -3426 1206 -3426 0 net=12299
rlabel metal2 1248 -3426 1248 -3426 0 net=10606
rlabel metal2 1321 -3426 1321 -3426 0 net=12961
rlabel metal2 1360 -3426 1360 -3426 0 net=12585
rlabel metal2 1360 -3426 1360 -3426 0 net=12585
rlabel metal2 1444 -3426 1444 -3426 0 net=11619
rlabel metal2 1521 -3426 1521 -3426 0 net=12719
rlabel metal2 1521 -3426 1521 -3426 0 net=12719
rlabel metal2 1612 -3426 1612 -3426 0 net=12120
rlabel metal2 1640 -3426 1640 -3426 0 net=14587
rlabel metal2 1724 -3426 1724 -3426 0 net=13903
rlabel metal2 1738 -3426 1738 -3426 0 net=11288
rlabel metal2 1759 -3426 1759 -3426 0 net=11986
rlabel metal2 1780 -3426 1780 -3426 0 net=13375
rlabel metal2 1780 -3426 1780 -3426 0 net=13375
rlabel metal2 1794 -3426 1794 -3426 0 net=13569
rlabel metal2 1822 -3426 1822 -3426 0 net=13053
rlabel metal2 1850 -3426 1850 -3426 0 net=13927
rlabel metal2 1850 -3426 1850 -3426 0 net=13927
rlabel metal2 1857 -3426 1857 -3426 0 net=14269
rlabel metal2 373 -3428 373 -3428 0 net=2270
rlabel metal2 492 -3428 492 -3428 0 net=5159
rlabel metal2 576 -3428 576 -3428 0 net=4628
rlabel metal2 576 -3428 576 -3428 0 net=4628
rlabel metal2 611 -3428 611 -3428 0 net=2062
rlabel metal2 653 -3428 653 -3428 0 net=3587
rlabel metal2 684 -3428 684 -3428 0 net=7590
rlabel metal2 744 -3428 744 -3428 0 net=4413
rlabel metal2 793 -3428 793 -3428 0 net=6121
rlabel metal2 793 -3428 793 -3428 0 net=6121
rlabel metal2 807 -3428 807 -3428 0 net=6749
rlabel metal2 992 -3428 992 -3428 0 net=10290
rlabel metal2 1066 -3428 1066 -3428 0 net=11597
rlabel metal2 1108 -3428 1108 -3428 0 net=7683
rlabel metal2 1220 -3428 1220 -3428 0 net=9550
rlabel metal2 1461 -3428 1461 -3428 0 net=10740
rlabel metal2 1724 -3428 1724 -3428 0 net=13745
rlabel metal2 1766 -3428 1766 -3428 0 net=6317
rlabel metal2 1829 -3428 1829 -3428 0 net=13265
rlabel metal2 1857 -3428 1857 -3428 0 net=14022
rlabel metal2 408 -3430 408 -3430 0 net=5020
rlabel metal2 499 -3430 499 -3430 0 net=4907
rlabel metal2 625 -3430 625 -3430 0 net=3535
rlabel metal2 695 -3430 695 -3430 0 net=2754
rlabel metal2 1052 -3430 1052 -3430 0 net=10807
rlabel metal2 1101 -3430 1101 -3430 0 net=6629
rlabel metal2 1255 -3430 1255 -3430 0 net=10970
rlabel metal2 1325 -3430 1325 -3430 0 net=8545
rlabel metal2 1381 -3430 1381 -3430 0 net=12607
rlabel metal2 1836 -3430 1836 -3430 0 net=6959
rlabel metal2 1864 -3430 1864 -3430 0 net=14715
rlabel metal2 450 -3432 450 -3432 0 net=3847
rlabel metal2 506 -3432 506 -3432 0 net=5047
rlabel metal2 653 -3432 653 -3432 0 net=8865
rlabel metal2 702 -3432 702 -3432 0 net=3460
rlabel metal2 1003 -3432 1003 -3432 0 net=7211
rlabel metal2 1069 -3432 1069 -3432 0 net=397
rlabel metal2 1136 -3432 1136 -3432 0 net=8355
rlabel metal2 1276 -3432 1276 -3432 0 net=14058
rlabel metal2 1451 -3432 1451 -3432 0 net=11683
rlabel metal2 422 -3434 422 -3434 0 net=9461
rlabel metal2 534 -3434 534 -3434 0 net=8461
rlabel metal2 534 -3434 534 -3434 0 net=8461
rlabel metal2 548 -3434 548 -3434 0 net=3568
rlabel metal2 660 -3434 660 -3434 0 net=4199
rlabel metal2 702 -3434 702 -3434 0 net=9454
rlabel metal2 814 -3434 814 -3434 0 net=6196
rlabel metal2 863 -3434 863 -3434 0 net=5915
rlabel metal2 901 -3434 901 -3434 0 net=11740
rlabel metal2 1108 -3434 1108 -3434 0 net=2473
rlabel metal2 1867 -3434 1867 -3434 0 net=1
rlabel metal2 380 -3436 380 -3436 0 net=2037
rlabel metal2 464 -3436 464 -3436 0 net=3231
rlabel metal2 555 -3436 555 -3436 0 net=9220
rlabel metal2 660 -3436 660 -3436 0 net=12803
rlabel metal2 709 -3436 709 -3436 0 net=3352
rlabel metal2 912 -3436 912 -3436 0 net=7555
rlabel metal2 1010 -3436 1010 -3436 0 net=9302
rlabel metal2 1143 -3436 1143 -3436 0 net=8229
rlabel metal2 331 -3438 331 -3438 0 net=5026
rlabel metal2 541 -3438 541 -3438 0 net=5799
rlabel metal2 558 -3438 558 -3438 0 net=8664
rlabel metal2 814 -3438 814 -3438 0 net=8067
rlabel metal2 835 -3438 835 -3438 0 net=8778
rlabel metal2 915 -3438 915 -3438 0 net=9444
rlabel metal2 982 -3438 982 -3438 0 net=3299
rlabel metal2 1017 -3438 1017 -3438 0 net=7343
rlabel metal2 1017 -3438 1017 -3438 0 net=7343
rlabel metal2 1034 -3438 1034 -3438 0 net=6011
rlabel metal2 1115 -3438 1115 -3438 0 net=8264
rlabel metal2 1185 -3438 1185 -3438 0 net=2779
rlabel metal2 359 -3440 359 -3440 0 net=1653
rlabel metal2 541 -3440 541 -3440 0 net=6799
rlabel metal2 674 -3440 674 -3440 0 net=7785
rlabel metal2 737 -3440 737 -3440 0 net=1963
rlabel metal2 835 -3440 835 -3440 0 net=6905
rlabel metal2 919 -3440 919 -3440 0 net=9214
rlabel metal2 1073 -3440 1073 -3440 0 net=7043
rlabel metal2 562 -3442 562 -3442 0 net=5375
rlabel metal2 604 -3442 604 -3442 0 net=2335
rlabel metal2 681 -3442 681 -3442 0 net=4329
rlabel metal2 744 -3442 744 -3442 0 net=9955
rlabel metal2 842 -3442 842 -3442 0 net=10479
rlabel metal2 947 -3442 947 -3442 0 net=8283
rlabel metal2 1059 -3442 1059 -3442 0 net=10597
rlabel metal2 1080 -3442 1080 -3442 0 net=6577
rlabel metal2 1157 -3442 1157 -3442 0 net=14155
rlabel metal2 1157 -3442 1157 -3442 0 net=14155
rlabel metal2 1164 -3442 1164 -3442 0 net=13877
rlabel metal2 520 -3444 520 -3444 0 net=13506
rlabel metal2 751 -3444 751 -3444 0 net=10312
rlabel metal2 1192 -3444 1192 -3444 0 net=12985
rlabel metal2 436 -3446 436 -3446 0 net=661
rlabel metal2 569 -3446 569 -3446 0 net=11213
rlabel metal2 751 -3446 751 -3446 0 net=10705
rlabel metal2 877 -3446 877 -3446 0 net=1890
rlabel metal2 1083 -3446 1083 -3446 0 net=14402
rlabel metal2 1227 -3446 1227 -3446 0 net=11251
rlabel metal2 527 -3448 527 -3448 0 net=4295
rlabel metal2 583 -3448 583 -3448 0 net=7461
rlabel metal2 632 -3448 632 -3448 0 net=13943
rlabel metal2 1087 -3448 1087 -3448 0 net=5649
rlabel metal2 513 -3450 513 -3450 0 net=2225
rlabel metal2 590 -3450 590 -3450 0 net=4985
rlabel metal2 730 -3450 730 -3450 0 net=3859
rlabel metal2 877 -3450 877 -3450 0 net=10445
rlabel metal2 954 -3450 954 -3450 0 net=12475
rlabel metal2 1171 -3450 1171 -3450 0 net=4847
rlabel metal2 457 -3452 457 -3452 0 net=1921
rlabel metal2 730 -3452 730 -3452 0 net=13034
rlabel metal2 996 -3452 996 -3452 0 net=10517
rlabel metal2 1178 -3452 1178 -3452 0 net=9139
rlabel metal2 443 -3454 443 -3454 0 net=2721
rlabel metal2 590 -3454 590 -3454 0 net=13707
rlabel metal2 1178 -3454 1178 -3454 0 net=13439
rlabel metal2 439 -3456 439 -3456 0 net=5827
rlabel metal2 765 -3456 765 -3456 0 net=4405
rlabel metal2 772 -3458 772 -3458 0 net=7479
rlabel metal2 271 -3469 271 -3469 0 net=353
rlabel metal2 369 -3469 369 -3469 0 net=7803
rlabel metal2 415 -3469 415 -3469 0 net=4240
rlabel metal2 439 -3469 439 -3469 0 net=5828
rlabel metal2 457 -3469 457 -3469 0 net=2723
rlabel metal2 478 -3469 478 -3469 0 net=5161
rlabel metal2 499 -3469 499 -3469 0 net=3232
rlabel metal2 569 -3469 569 -3469 0 net=4296
rlabel metal2 642 -3469 642 -3469 0 net=10706
rlabel metal2 765 -3469 765 -3469 0 net=6751
rlabel metal2 828 -3469 828 -3469 0 net=1964
rlabel metal2 919 -3469 919 -3469 0 net=12476
rlabel metal2 975 -3469 975 -3469 0 net=7557
rlabel metal2 1031 -3469 1031 -3469 0 net=7212
rlabel metal2 1066 -3469 1066 -3469 0 net=11599
rlabel metal2 1066 -3469 1066 -3469 0 net=11599
rlabel metal2 1080 -3469 1080 -3469 0 net=2475
rlabel metal2 1122 -3469 1122 -3469 0 net=2780
rlabel metal2 1199 -3469 1199 -3469 0 net=7684
rlabel metal2 1360 -3469 1360 -3469 0 net=12587
rlabel metal2 1360 -3469 1360 -3469 0 net=12587
rlabel metal2 1430 -3469 1430 -3469 0 net=11620
rlabel metal2 1458 -3469 1458 -3469 0 net=5429
rlabel metal2 1640 -3469 1640 -3469 0 net=14589
rlabel metal2 1640 -3469 1640 -3469 0 net=14589
rlabel metal2 1724 -3469 1724 -3469 0 net=13746
rlabel metal2 1724 -3469 1724 -3469 0 net=13746
rlabel metal2 1731 -3469 1731 -3469 0 net=13905
rlabel metal2 1731 -3469 1731 -3469 0 net=13905
rlabel metal2 1745 -3469 1745 -3469 0 net=6318
rlabel metal2 1780 -3469 1780 -3469 0 net=13377
rlabel metal2 1780 -3469 1780 -3469 0 net=13377
rlabel metal2 1790 -3469 1790 -3469 0 net=13570
rlabel metal2 1829 -3469 1829 -3469 0 net=13266
rlabel metal2 1839 -3469 1839 -3469 0 net=13928
rlabel metal2 1860 -3469 1860 -3469 0 net=14716
rlabel metal2 1955 -3469 1955 -3469 0 net=14696
rlabel metal2 1955 -3469 1955 -3469 0 net=14696
rlabel metal2 1958 -3469 1958 -3469 0 net=6046
rlabel metal2 2025 -3469 2025 -3469 0 net=3387
rlabel metal2 324 -3471 324 -3471 0 net=2687
rlabel metal2 380 -3471 380 -3471 0 net=1655
rlabel metal2 422 -3471 422 -3471 0 net=2038
rlabel metal2 485 -3471 485 -3471 0 net=3848
rlabel metal2 541 -3471 541 -3471 0 net=6801
rlabel metal2 579 -3471 579 -3471 0 net=2336
rlabel metal2 618 -3471 618 -3471 0 net=5225
rlabel metal2 639 -3471 639 -3471 0 net=8867
rlabel metal2 667 -3471 667 -3471 0 net=3536
rlabel metal2 730 -3471 730 -3471 0 net=4330
rlabel metal2 772 -3471 772 -3471 0 net=7481
rlabel metal2 789 -3471 789 -3471 0 net=8068
rlabel metal2 828 -3471 828 -3471 0 net=10481
rlabel metal2 849 -3471 849 -3471 0 net=3860
rlabel metal2 975 -3471 975 -3471 0 net=10519
rlabel metal2 1017 -3471 1017 -3471 0 net=7345
rlabel metal2 1052 -3471 1052 -3471 0 net=10809
rlabel metal2 1052 -3471 1052 -3471 0 net=10809
rlabel metal2 1059 -3471 1059 -3471 0 net=10598
rlabel metal2 1083 -3471 1083 -3471 0 net=4848
rlabel metal2 1178 -3471 1178 -3471 0 net=12300
rlabel metal2 1213 -3471 1213 -3471 0 net=13440
rlabel metal2 1276 -3471 1276 -3471 0 net=10913
rlabel metal2 1307 -3471 1307 -3471 0 net=14032
rlabel metal2 1433 -3471 1433 -3471 0 net=11684
rlabel metal2 1500 -3471 1500 -3471 0 net=10280
rlabel metal2 1507 -3471 1507 -3471 0 net=14125
rlabel metal2 1521 -3471 1521 -3471 0 net=12721
rlabel metal2 1521 -3471 1521 -3471 0 net=12721
rlabel metal2 1843 -3471 1843 -3471 0 net=6961
rlabel metal2 1864 -3471 1864 -3471 0 net=14271
rlabel metal2 2025 -3471 2025 -3471 0 net=13687
rlabel metal2 471 -3473 471 -3473 0 net=6551
rlabel metal2 562 -3473 562 -3473 0 net=5377
rlabel metal2 646 -3473 646 -3473 0 net=5049
rlabel metal2 646 -3473 646 -3473 0 net=5049
rlabel metal2 653 -3473 653 -3473 0 net=9956
rlabel metal2 793 -3473 793 -3473 0 net=6123
rlabel metal2 793 -3473 793 -3473 0 net=6123
rlabel metal2 800 -3473 800 -3473 0 net=8040
rlabel metal2 1010 -3473 1010 -3473 0 net=3301
rlabel metal2 1045 -3473 1045 -3473 0 net=13708
rlabel metal2 1822 -3473 1822 -3473 0 net=13055
rlabel metal2 2028 -3473 2028 -3473 0 net=1
rlabel metal2 485 -3475 485 -3475 0 net=13945
rlabel metal2 674 -3475 674 -3475 0 net=4986
rlabel metal2 709 -3475 709 -3475 0 net=7787
rlabel metal2 814 -3475 814 -3475 0 net=6907
rlabel metal2 866 -3475 866 -3475 0 net=5650
rlabel metal2 1094 -3475 1094 -3475 0 net=6012
rlabel metal2 1129 -3475 1129 -3475 0 net=6579
rlabel metal2 1178 -3475 1178 -3475 0 net=12987
rlabel metal2 1234 -3475 1234 -3475 0 net=8230
rlabel metal2 1269 -3475 1269 -3475 0 net=8546
rlabel metal2 1437 -3475 1437 -3475 0 net=3685
rlabel metal2 1437 -3475 1437 -3475 0 net=3685
rlabel metal2 1493 -3475 1493 -3475 0 net=10625
rlabel metal2 506 -3477 506 -3477 0 net=9463
rlabel metal2 583 -3477 583 -3477 0 net=2227
rlabel metal2 583 -3477 583 -3477 0 net=2227
rlabel metal2 590 -3477 590 -3477 0 net=7462
rlabel metal2 632 -3477 632 -3477 0 net=12805
rlabel metal2 681 -3477 681 -3477 0 net=7855
rlabel metal2 821 -3477 821 -3477 0 net=4407
rlabel metal2 870 -3477 870 -3477 0 net=10447
rlabel metal2 884 -3477 884 -3477 0 net=5916
rlabel metal2 1003 -3477 1003 -3477 0 net=8285
rlabel metal2 1038 -3477 1038 -3477 0 net=9095
rlabel metal2 1059 -3477 1059 -3477 0 net=6631
rlabel metal2 1157 -3477 1157 -3477 0 net=14157
rlabel metal2 1220 -3477 1220 -3477 0 net=8357
rlabel metal2 1255 -3477 1255 -3477 0 net=2805
rlabel metal2 1311 -3477 1311 -3477 0 net=12962
rlabel metal2 1465 -3477 1465 -3477 0 net=12609
rlabel metal2 520 -3479 520 -3479 0 net=1785
rlabel metal2 1024 -3479 1024 -3479 0 net=7149
rlabel metal2 1248 -3479 1248 -3479 0 net=7045
rlabel metal2 534 -3481 534 -3481 0 net=8463
rlabel metal2 611 -3481 611 -3481 0 net=4909
rlabel metal2 695 -3481 695 -3481 0 net=4200
rlabel metal2 1024 -3481 1024 -3481 0 net=13879
rlabel metal2 1241 -3481 1241 -3481 0 net=11252
rlabel metal2 1283 -3481 1283 -3481 0 net=11928
rlabel metal2 513 -3483 513 -3483 0 net=1923
rlabel metal2 555 -3483 555 -3483 0 net=5801
rlabel metal2 716 -3483 716 -3483 0 net=11215
rlabel metal2 1227 -3483 1227 -3483 0 net=9141
rlabel metal2 1290 -3483 1290 -3483 0 net=3965
rlabel metal2 688 -3485 688 -3485 0 net=3589
rlabel metal2 737 -3485 737 -3485 0 net=4415
rlabel metal2 723 -3487 723 -3487 0 net=11629
rlabel metal2 331 -3498 331 -3498 0 net=2688
rlabel metal2 394 -3498 394 -3498 0 net=7804
rlabel metal2 432 -3498 432 -3498 0 net=6552
rlabel metal2 478 -3498 478 -3498 0 net=5163
rlabel metal2 478 -3498 478 -3498 0 net=5163
rlabel metal2 523 -3498 523 -3498 0 net=1274
rlabel metal2 681 -3498 681 -3498 0 net=4911
rlabel metal2 716 -3498 716 -3498 0 net=3591
rlabel metal2 737 -3498 737 -3498 0 net=4417
rlabel metal2 737 -3498 737 -3498 0 net=4417
rlabel metal2 775 -3498 775 -3498 0 net=11965
rlabel metal2 968 -3498 968 -3498 0 net=10521
rlabel metal2 996 -3498 996 -3498 0 net=7559
rlabel metal2 1010 -3498 1010 -3498 0 net=8287
rlabel metal2 1010 -3498 1010 -3498 0 net=8287
rlabel metal2 1017 -3498 1017 -3498 0 net=3303
rlabel metal2 1017 -3498 1017 -3498 0 net=3303
rlabel metal2 1038 -3498 1038 -3498 0 net=7150
rlabel metal2 1122 -3498 1122 -3498 0 net=3967
rlabel metal2 1304 -3498 1304 -3498 0 net=7046
rlabel metal2 1430 -3498 1430 -3498 0 net=3686
rlabel metal2 1500 -3498 1500 -3498 0 net=14126
rlabel metal2 1514 -3498 1514 -3498 0 net=10627
rlabel metal2 1514 -3498 1514 -3498 0 net=10627
rlabel metal2 1521 -3498 1521 -3498 0 net=12723
rlabel metal2 1521 -3498 1521 -3498 0 net=12723
rlabel metal2 1570 -3498 1570 -3498 0 net=5431
rlabel metal2 1640 -3498 1640 -3498 0 net=14591
rlabel metal2 1640 -3498 1640 -3498 0 net=14591
rlabel metal2 1724 -3498 1724 -3498 0 net=13906
rlabel metal2 1780 -3498 1780 -3498 0 net=13378
rlabel metal2 1850 -3498 1850 -3498 0 net=6962
rlabel metal2 2025 -3498 2025 -3498 0 net=13689
rlabel metal2 2025 -3498 2025 -3498 0 net=13689
rlabel metal2 2032 -3498 2032 -3498 0 net=3389
rlabel metal2 2032 -3498 2032 -3498 0 net=3389
rlabel metal2 387 -3500 387 -3500 0 net=1657
rlabel metal2 429 -3500 429 -3500 0 net=13947
rlabel metal2 534 -3500 534 -3500 0 net=1925
rlabel metal2 569 -3500 569 -3500 0 net=6803
rlabel metal2 583 -3500 583 -3500 0 net=2229
rlabel metal2 583 -3500 583 -3500 0 net=2229
rlabel metal2 625 -3500 625 -3500 0 net=12807
rlabel metal2 639 -3500 639 -3500 0 net=8869
rlabel metal2 639 -3500 639 -3500 0 net=8869
rlabel metal2 646 -3500 646 -3500 0 net=5050
rlabel metal2 779 -3500 779 -3500 0 net=11217
rlabel metal2 810 -3500 810 -3500 0 net=10482
rlabel metal2 842 -3500 842 -3500 0 net=4408
rlabel metal2 884 -3500 884 -3500 0 net=13880
rlabel metal2 1038 -3500 1038 -3500 0 net=9097
rlabel metal2 1052 -3500 1052 -3500 0 net=10811
rlabel metal2 1052 -3500 1052 -3500 0 net=10811
rlabel metal2 1143 -3500 1143 -3500 0 net=6581
rlabel metal2 1160 -3500 1160 -3500 0 net=12988
rlabel metal2 1192 -3500 1192 -3500 0 net=14159
rlabel metal2 1234 -3500 1234 -3500 0 net=8358
rlabel metal2 1262 -3500 1262 -3500 0 net=10914
rlabel metal2 1283 -3500 1283 -3500 0 net=1042
rlabel metal2 1360 -3500 1360 -3500 0 net=12589
rlabel metal2 1360 -3500 1360 -3500 0 net=12589
rlabel metal2 1493 -3500 1493 -3500 0 net=12611
rlabel metal2 1843 -3500 1843 -3500 0 net=13057
rlabel metal2 1857 -3500 1857 -3500 0 net=14272
rlabel metal2 464 -3502 464 -3502 0 net=2725
rlabel metal2 464 -3502 464 -3502 0 net=2725
rlabel metal2 541 -3502 541 -3502 0 net=9465
rlabel metal2 541 -3502 541 -3502 0 net=9465
rlabel metal2 611 -3502 611 -3502 0 net=5803
rlabel metal2 751 -3502 751 -3502 0 net=7857
rlabel metal2 789 -3502 789 -3502 0 net=6908
rlabel metal2 863 -3502 863 -3502 0 net=10448
rlabel metal2 898 -3502 898 -3502 0 net=1787
rlabel metal2 1031 -3502 1031 -3502 0 net=7347
rlabel metal2 1234 -3502 1234 -3502 0 net=2807
rlabel metal2 611 -3504 611 -3504 0 net=5227
rlabel metal2 751 -3504 751 -3504 0 net=11631
rlabel metal2 793 -3504 793 -3504 0 net=6125
rlabel metal2 793 -3504 793 -3504 0 net=6125
rlabel metal2 1031 -3504 1031 -3504 0 net=6633
rlabel metal2 1241 -3504 1241 -3504 0 net=9142
rlabel metal2 604 -3506 604 -3506 0 net=5379
rlabel metal2 744 -3506 744 -3506 0 net=7789
rlabel metal2 1059 -3506 1059 -3506 0 net=11600
rlabel metal2 590 -3508 590 -3508 0 net=8465
rlabel metal2 744 -3508 744 -3508 0 net=6753
rlabel metal2 1066 -3508 1066 -3508 0 net=2477
rlabel metal2 765 -3510 765 -3510 0 net=7483
rlabel metal2 394 -3521 394 -3521 0 net=1659
rlabel metal2 394 -3521 394 -3521 0 net=1659
rlabel metal2 408 -3521 408 -3521 0 net=13949
rlabel metal2 464 -3521 464 -3521 0 net=2727
rlabel metal2 464 -3521 464 -3521 0 net=2727
rlabel metal2 478 -3521 478 -3521 0 net=5165
rlabel metal2 478 -3521 478 -3521 0 net=5165
rlabel metal2 541 -3521 541 -3521 0 net=9467
rlabel metal2 541 -3521 541 -3521 0 net=9467
rlabel metal2 548 -3521 548 -3521 0 net=1927
rlabel metal2 548 -3521 548 -3521 0 net=1927
rlabel metal2 576 -3521 576 -3521 0 net=6805
rlabel metal2 576 -3521 576 -3521 0 net=6805
rlabel metal2 583 -3521 583 -3521 0 net=2231
rlabel metal2 583 -3521 583 -3521 0 net=2231
rlabel metal2 618 -3521 618 -3521 0 net=5380
rlabel metal2 639 -3521 639 -3521 0 net=8871
rlabel metal2 639 -3521 639 -3521 0 net=8871
rlabel metal2 709 -3521 709 -3521 0 net=4913
rlabel metal2 723 -3521 723 -3521 0 net=4419
rlabel metal2 744 -3521 744 -3521 0 net=6755
rlabel metal2 744 -3521 744 -3521 0 net=6755
rlabel metal2 751 -3521 751 -3521 0 net=11632
rlabel metal2 793 -3521 793 -3521 0 net=6127
rlabel metal2 793 -3521 793 -3521 0 net=6127
rlabel metal2 800 -3521 800 -3521 0 net=11218
rlabel metal2 891 -3521 891 -3521 0 net=11967
rlabel metal2 968 -3521 968 -3521 0 net=10522
rlabel metal2 1017 -3521 1017 -3521 0 net=3304
rlabel metal2 1031 -3521 1031 -3521 0 net=6635
rlabel metal2 1031 -3521 1031 -3521 0 net=6635
rlabel metal2 1038 -3521 1038 -3521 0 net=9099
rlabel metal2 1059 -3521 1059 -3521 0 net=2478
rlabel metal2 1150 -3521 1150 -3521 0 net=6582
rlabel metal2 1206 -3521 1206 -3521 0 net=14161
rlabel metal2 1223 -3521 1223 -3521 0 net=2808
rlabel metal2 1360 -3521 1360 -3521 0 net=12590
rlabel metal2 1507 -3521 1507 -3521 0 net=12613
rlabel metal2 1521 -3521 1521 -3521 0 net=12725
rlabel metal2 1521 -3521 1521 -3521 0 net=12725
rlabel metal2 1612 -3521 1612 -3521 0 net=5433
rlabel metal2 1640 -3521 1640 -3521 0 net=14593
rlabel metal2 1640 -3521 1640 -3521 0 net=14593
rlabel metal2 1850 -3521 1850 -3521 0 net=13058
rlabel metal2 2025 -3521 2025 -3521 0 net=13691
rlabel metal2 2025 -3521 2025 -3521 0 net=13691
rlabel metal2 2032 -3521 2032 -3521 0 net=3391
rlabel metal2 2032 -3521 2032 -3521 0 net=3391
rlabel metal2 611 -3523 611 -3523 0 net=5229
rlabel metal2 632 -3523 632 -3523 0 net=5805
rlabel metal2 709 -3523 709 -3523 0 net=8707
rlabel metal2 758 -3523 758 -3523 0 net=7790
rlabel metal2 779 -3523 779 -3523 0 net=7859
rlabel metal2 1024 -3523 1024 -3523 0 net=1788
rlabel metal2 1507 -3523 1507 -3523 0 net=10629
rlabel metal2 604 -3525 604 -3525 0 net=8467
rlabel metal2 730 -3525 730 -3525 0 net=3593
rlabel metal2 730 -3525 730 -3525 0 net=3593
rlabel metal2 765 -3525 765 -3525 0 net=7484
rlabel metal2 1010 -3525 1010 -3525 0 net=8288
rlabel metal2 1038 -3525 1038 -3525 0 net=7348
rlabel metal2 1052 -3525 1052 -3525 0 net=10813
rlabel metal2 1066 -3525 1066 -3525 0 net=3969
rlabel metal2 604 -3527 604 -3527 0 net=12809
rlabel metal2 765 -3527 765 -3527 0 net=11097
rlabel metal2 1003 -3527 1003 -3527 0 net=7561
rlabel metal2 1510 -3527 1510 -3527 0 net=1
rlabel metal2 625 -3529 625 -3529 0 net=104
rlabel metal2 394 -3540 394 -3540 0 net=1661
rlabel metal2 408 -3540 408 -3540 0 net=13951
rlabel metal2 408 -3540 408 -3540 0 net=13951
rlabel metal2 464 -3540 464 -3540 0 net=2728
rlabel metal2 541 -3540 541 -3540 0 net=9469
rlabel metal2 541 -3540 541 -3540 0 net=9469
rlabel metal2 548 -3540 548 -3540 0 net=1929
rlabel metal2 583 -3540 583 -3540 0 net=2233
rlabel metal2 604 -3540 604 -3540 0 net=12811
rlabel metal2 604 -3540 604 -3540 0 net=12811
rlabel metal2 611 -3540 611 -3540 0 net=8469
rlabel metal2 611 -3540 611 -3540 0 net=8469
rlabel metal2 618 -3540 618 -3540 0 net=5231
rlabel metal2 618 -3540 618 -3540 0 net=5231
rlabel metal2 635 -3540 635 -3540 0 net=8872
rlabel metal2 646 -3540 646 -3540 0 net=5807
rlabel metal2 646 -3540 646 -3540 0 net=5807
rlabel metal2 702 -3540 702 -3540 0 net=8709
rlabel metal2 716 -3540 716 -3540 0 net=4915
rlabel metal2 716 -3540 716 -3540 0 net=4915
rlabel metal2 723 -3540 723 -3540 0 net=4421
rlabel metal2 723 -3540 723 -3540 0 net=4421
rlabel metal2 730 -3540 730 -3540 0 net=3594
rlabel metal2 758 -3540 758 -3540 0 net=11099
rlabel metal2 786 -3540 786 -3540 0 net=7860
rlabel metal2 793 -3540 793 -3540 0 net=6129
rlabel metal2 793 -3540 793 -3540 0 net=6129
rlabel metal2 926 -3540 926 -3540 0 net=11968
rlabel metal2 1010 -3540 1010 -3540 0 net=7562
rlabel metal2 1027 -3540 1027 -3540 0 net=6636
rlabel metal2 1038 -3540 1038 -3540 0 net=9100
rlabel metal2 1059 -3540 1059 -3540 0 net=10815
rlabel metal2 1059 -3540 1059 -3540 0 net=10815
rlabel metal2 1213 -3540 1213 -3540 0 net=14162
rlabel metal2 1507 -3540 1507 -3540 0 net=10631
rlabel metal2 1514 -3540 1514 -3540 0 net=12615
rlabel metal2 1514 -3540 1514 -3540 0 net=12615
rlabel metal2 1640 -3540 1640 -3540 0 net=14595
rlabel metal2 2025 -3540 2025 -3540 0 net=13693
rlabel metal2 2025 -3540 2025 -3540 0 net=13693
rlabel metal2 2032 -3540 2032 -3540 0 net=3393
rlabel metal2 2032 -3540 2032 -3540 0 net=3393
rlabel metal2 471 -3542 471 -3542 0 net=5166
rlabel metal2 576 -3542 576 -3542 0 net=6806
rlabel metal2 730 -3542 730 -3542 0 net=6757
rlabel metal2 1038 -3542 1038 -3542 0 net=3971
rlabel metal2 1507 -3542 1507 -3542 0 net=12727
rlabel metal2 1633 -3542 1633 -3542 0 net=5435
rlabel metal2 401 -3555 401 -3555 0 net=1663
rlabel metal2 541 -3555 541 -3555 0 net=9470
rlabel metal2 551 -3555 551 -3555 0 net=1930
rlabel metal2 586 -3555 586 -3555 0 net=2234
rlabel metal2 604 -3555 604 -3555 0 net=12813
rlabel metal2 618 -3555 618 -3555 0 net=5233
rlabel metal2 618 -3555 618 -3555 0 net=5233
rlabel metal2 646 -3555 646 -3555 0 net=5808
rlabel metal2 702 -3555 702 -3555 0 net=8711
rlabel metal2 702 -3555 702 -3555 0 net=8711
rlabel metal2 716 -3555 716 -3555 0 net=4917
rlabel metal2 716 -3555 716 -3555 0 net=4917
rlabel metal2 723 -3555 723 -3555 0 net=4423
rlabel metal2 723 -3555 723 -3555 0 net=4423
rlabel metal2 730 -3555 730 -3555 0 net=6759
rlabel metal2 730 -3555 730 -3555 0 net=6759
rlabel metal2 758 -3555 758 -3555 0 net=11101
rlabel metal2 758 -3555 758 -3555 0 net=11101
rlabel metal2 789 -3555 789 -3555 0 net=6130
rlabel metal2 1017 -3555 1017 -3555 0 net=3972
rlabel metal2 1059 -3555 1059 -3555 0 net=10817
rlabel metal2 1517 -3555 1517 -3555 0 net=10632
rlabel metal2 1640 -3555 1640 -3555 0 net=5437
rlabel metal2 1640 -3555 1640 -3555 0 net=5437
rlabel metal2 1647 -3555 1647 -3555 0 net=14597
rlabel metal2 1647 -3555 1647 -3555 0 net=14597
rlabel metal2 2025 -3555 2025 -3555 0 net=13694
rlabel metal2 2025 -3555 2025 -3555 0 net=13694
rlabel metal2 2028 -3555 2028 -3555 0 net=3394
rlabel metal2 401 -3557 401 -3557 0 net=13953
rlabel metal2 604 -3557 604 -3557 0 net=8471
rlabel metal2 1514 -3557 1514 -3557 0 net=12617
rlabel metal2 607 -3559 607 -3559 0 net=1
rlabel metal2 1507 -3559 1507 -3559 0 net=12728
rlabel metal2 401 -3570 401 -3570 0 net=13955
rlabel metal2 604 -3570 604 -3570 0 net=8473
rlabel metal2 604 -3570 604 -3570 0 net=8473
rlabel metal2 611 -3570 611 -3570 0 net=12815
rlabel metal2 611 -3570 611 -3570 0 net=12815
rlabel metal2 618 -3570 618 -3570 0 net=5235
rlabel metal2 618 -3570 618 -3570 0 net=5235
rlabel metal2 702 -3570 702 -3570 0 net=8713
rlabel metal2 702 -3570 702 -3570 0 net=8713
rlabel metal2 716 -3570 716 -3570 0 net=4919
rlabel metal2 716 -3570 716 -3570 0 net=4919
rlabel metal2 723 -3570 723 -3570 0 net=4425
rlabel metal2 723 -3570 723 -3570 0 net=4425
rlabel metal2 730 -3570 730 -3570 0 net=6761
rlabel metal2 730 -3570 730 -3570 0 net=6761
rlabel metal2 758 -3570 758 -3570 0 net=11103
rlabel metal2 758 -3570 758 -3570 0 net=11103
rlabel metal2 1062 -3570 1062 -3570 0 net=10818
rlabel metal2 1514 -3570 1514 -3570 0 net=12618
rlabel metal2 1640 -3570 1640 -3570 0 net=5439
rlabel metal2 1640 -3570 1640 -3570 0 net=5439
rlabel metal2 1647 -3570 1647 -3570 0 net=14599
rlabel metal2 1647 -3570 1647 -3570 0 net=14599
rlabel metal2 401 -3572 401 -3572 0 net=1665
rlabel metal2 394 -3585 394 -3585 0 net=1667
rlabel metal2 604 -3585 604 -3585 0 net=8475
rlabel metal2 604 -3585 604 -3585 0 net=8475
rlabel metal2 611 -3585 611 -3585 0 net=12817
rlabel metal2 611 -3585 611 -3585 0 net=12817
rlabel metal2 618 -3585 618 -3585 0 net=5236
rlabel metal2 702 -3585 702 -3585 0 net=8715
rlabel metal2 702 -3585 702 -3585 0 net=8715
rlabel metal2 723 -3585 723 -3585 0 net=4426
rlabel metal2 730 -3585 730 -3585 0 net=6763
rlabel metal2 730 -3585 730 -3585 0 net=6763
rlabel metal2 758 -3585 758 -3585 0 net=11105
rlabel metal2 758 -3585 758 -3585 0 net=11105
rlabel metal2 1640 -3585 1640 -3585 0 net=5441
rlabel metal2 1640 -3585 1640 -3585 0 net=5441
rlabel metal2 1647 -3585 1647 -3585 0 net=14601
rlabel metal2 1647 -3585 1647 -3585 0 net=14601
rlabel metal2 401 -3587 401 -3587 0 net=13957
rlabel metal2 716 -3587 716 -3587 0 net=4920
rlabel metal2 394 -3598 394 -3598 0 net=1669
rlabel metal2 394 -3598 394 -3598 0 net=1669
rlabel metal2 401 -3598 401 -3598 0 net=13959
rlabel metal2 401 -3598 401 -3598 0 net=13959
rlabel metal2 604 -3598 604 -3598 0 net=8477
rlabel metal2 604 -3598 604 -3598 0 net=8477
rlabel metal2 611 -3598 611 -3598 0 net=12819
rlabel metal2 611 -3598 611 -3598 0 net=12819
rlabel metal2 702 -3598 702 -3598 0 net=8716
rlabel metal2 702 -3598 702 -3598 0 net=8716
rlabel metal2 723 -3598 723 -3598 0 net=6764
rlabel metal2 758 -3598 758 -3598 0 net=11107
rlabel metal2 758 -3598 758 -3598 0 net=11107
rlabel metal2 1640 -3598 1640 -3598 0 net=5443
rlabel metal2 1640 -3598 1640 -3598 0 net=5443
rlabel metal2 1647 -3598 1647 -3598 0 net=14603
rlabel metal2 1647 -3598 1647 -3598 0 net=14603
rlabel metal2 394 -3609 394 -3609 0 net=1671
rlabel metal2 394 -3609 394 -3609 0 net=1671
rlabel metal2 401 -3609 401 -3609 0 net=13961
rlabel metal2 401 -3609 401 -3609 0 net=13961
rlabel metal2 604 -3609 604 -3609 0 net=8479
rlabel metal2 604 -3609 604 -3609 0 net=8479
rlabel metal2 611 -3609 611 -3609 0 net=12821
rlabel metal2 611 -3609 611 -3609 0 net=12821
rlabel metal2 695 -3609 695 -3609 0 net=2809
rlabel metal2 758 -3609 758 -3609 0 net=11109
rlabel metal2 758 -3609 758 -3609 0 net=11109
rlabel metal2 1640 -3609 1640 -3609 0 net=5444
rlabel metal2 1647 -3609 1647 -3609 0 net=14605
rlabel metal2 1647 -3609 1647 -3609 0 net=14605
rlabel metal2 394 -3620 394 -3620 0 net=1673
rlabel metal2 394 -3620 394 -3620 0 net=1673
rlabel metal2 401 -3620 401 -3620 0 net=13963
rlabel metal2 401 -3620 401 -3620 0 net=13963
rlabel metal2 604 -3620 604 -3620 0 net=8481
rlabel metal2 604 -3620 604 -3620 0 net=8481
rlabel metal2 611 -3620 611 -3620 0 net=12823
rlabel metal2 611 -3620 611 -3620 0 net=12823
rlabel metal2 695 -3620 695 -3620 0 net=2811
rlabel metal2 695 -3620 695 -3620 0 net=2811
rlabel metal2 758 -3620 758 -3620 0 net=11111
rlabel metal2 1640 -3620 1640 -3620 0 net=14606
rlabel metal2 394 -3631 394 -3631 0 net=1675
rlabel metal2 394 -3631 394 -3631 0 net=1675
rlabel metal2 401 -3631 401 -3631 0 net=13965
rlabel metal2 401 -3631 401 -3631 0 net=13965
rlabel metal2 604 -3631 604 -3631 0 net=8483
rlabel metal2 604 -3631 604 -3631 0 net=8483
rlabel metal2 611 -3631 611 -3631 0 net=12825
rlabel metal2 611 -3631 611 -3631 0 net=12825
rlabel metal2 695 -3631 695 -3631 0 net=2813
rlabel metal2 695 -3631 695 -3631 0 net=2813
rlabel metal2 761 -3631 761 -3631 0 net=11112
rlabel metal2 394 -3642 394 -3642 0 net=1677
rlabel metal2 394 -3642 394 -3642 0 net=1677
rlabel metal2 401 -3642 401 -3642 0 net=13967
rlabel metal2 401 -3642 401 -3642 0 net=13967
rlabel metal2 604 -3642 604 -3642 0 net=8485
rlabel metal2 604 -3642 604 -3642 0 net=8485
rlabel metal2 611 -3642 611 -3642 0 net=12827
rlabel metal2 611 -3642 611 -3642 0 net=12827
rlabel metal2 695 -3642 695 -3642 0 net=2815
rlabel metal2 695 -3642 695 -3642 0 net=2815
rlabel metal2 394 -3653 394 -3653 0 net=1679
rlabel metal2 604 -3653 604 -3653 0 net=8487
rlabel metal2 604 -3653 604 -3653 0 net=8487
rlabel metal2 611 -3653 611 -3653 0 net=12828
rlabel metal2 611 -3653 611 -3653 0 net=12828
rlabel metal2 695 -3653 695 -3653 0 net=2816
rlabel metal2 394 -3655 394 -3655 0 net=13968
rlabel metal2 397 -3668 397 -3668 0 net=1680
rlabel metal2 604 -3668 604 -3668 0 net=8488
<< end >>
