magic
tech scmos
timestamp 1555016836 
<< pdiffusion >>
rect 1 -12 7 -6
rect 8 -12 14 -6
rect 15 -12 21 -6
rect 22 -12 28 -6
rect 29 -12 35 -6
rect 36 -12 42 -6
rect 43 -12 49 -6
rect 50 -12 56 -6
rect 57 -12 63 -6
rect 64 -12 70 -6
rect 71 -12 77 -6
rect 106 -12 112 -6
rect 113 -12 119 -6
rect 127 -12 133 -6
rect 134 -12 140 -6
rect 141 -12 147 -6
rect 155 -12 158 -6
rect 162 -12 165 -6
rect 169 -12 175 -6
rect 176 -12 179 -6
rect 183 -12 189 -6
rect 190 -12 193 -6
rect 197 -12 203 -6
rect 204 -12 210 -6
rect 211 -12 217 -6
rect 218 -12 224 -6
rect 225 -12 228 -6
rect 232 -12 238 -6
rect 239 -12 245 -6
rect 246 -12 249 -6
rect 253 -12 259 -6
rect 260 -12 263 -6
rect 267 -12 270 -6
rect 274 -12 280 -6
rect 281 -12 287 -6
rect 323 -12 329 -6
rect 1 -39 7 -33
rect 8 -39 14 -33
rect 15 -39 21 -33
rect 22 -39 28 -33
rect 29 -39 35 -33
rect 36 -39 42 -33
rect 43 -39 49 -33
rect 71 -39 77 -33
rect 78 -39 84 -33
rect 85 -39 88 -33
rect 92 -39 95 -33
rect 99 -39 105 -33
rect 106 -39 112 -33
rect 113 -39 119 -33
rect 120 -39 126 -33
rect 127 -39 133 -33
rect 134 -39 140 -33
rect 141 -39 144 -33
rect 148 -39 151 -33
rect 155 -39 158 -33
rect 162 -39 168 -33
rect 169 -39 172 -33
rect 176 -39 182 -33
rect 183 -39 186 -33
rect 190 -39 193 -33
rect 197 -39 200 -33
rect 204 -39 210 -33
rect 211 -39 217 -33
rect 218 -39 221 -33
rect 225 -39 231 -33
rect 232 -39 235 -33
rect 239 -39 242 -33
rect 246 -39 249 -33
rect 253 -39 256 -33
rect 260 -39 263 -33
rect 267 -39 270 -33
rect 274 -39 277 -33
rect 281 -39 287 -33
rect 288 -39 291 -33
rect 295 -39 298 -33
rect 302 -39 305 -33
rect 309 -39 315 -33
rect 316 -39 319 -33
rect 323 -39 329 -33
rect 330 -39 333 -33
rect 337 -39 343 -33
rect 344 -39 347 -33
rect 351 -39 354 -33
rect 358 -39 361 -33
rect 365 -39 371 -33
rect 372 -39 378 -33
rect 379 -39 382 -33
rect 386 -39 389 -33
rect 393 -39 399 -33
rect 400 -39 403 -33
rect 414 -39 420 -33
rect 1 -82 7 -76
rect 8 -82 14 -76
rect 15 -82 21 -76
rect 22 -82 28 -76
rect 29 -82 35 -76
rect 36 -82 42 -76
rect 43 -82 46 -76
rect 50 -82 53 -76
rect 57 -82 63 -76
rect 64 -82 67 -76
rect 71 -82 77 -76
rect 78 -82 81 -76
rect 85 -82 91 -76
rect 92 -82 98 -76
rect 99 -82 105 -76
rect 106 -82 109 -76
rect 113 -82 119 -76
rect 120 -82 126 -76
rect 127 -82 133 -76
rect 134 -82 137 -76
rect 141 -82 147 -76
rect 148 -82 151 -76
rect 155 -82 161 -76
rect 162 -82 165 -76
rect 169 -82 175 -76
rect 176 -82 182 -76
rect 183 -82 186 -76
rect 190 -82 196 -76
rect 197 -82 203 -76
rect 204 -82 210 -76
rect 211 -82 217 -76
rect 218 -82 224 -76
rect 225 -82 231 -76
rect 232 -82 235 -76
rect 239 -82 242 -76
rect 246 -82 249 -76
rect 253 -82 259 -76
rect 260 -82 263 -76
rect 267 -82 273 -76
rect 274 -82 280 -76
rect 281 -82 287 -76
rect 288 -82 291 -76
rect 295 -82 298 -76
rect 302 -82 305 -76
rect 309 -82 312 -76
rect 316 -82 319 -76
rect 323 -82 326 -76
rect 330 -82 333 -76
rect 337 -82 340 -76
rect 344 -82 347 -76
rect 351 -82 357 -76
rect 358 -82 361 -76
rect 365 -82 368 -76
rect 372 -82 375 -76
rect 379 -82 382 -76
rect 386 -82 389 -76
rect 393 -82 396 -76
rect 400 -82 403 -76
rect 407 -82 410 -76
rect 428 -82 434 -76
rect 1 -127 7 -121
rect 8 -127 14 -121
rect 15 -127 21 -121
rect 22 -127 28 -121
rect 29 -127 35 -121
rect 36 -127 42 -121
rect 43 -127 49 -121
rect 50 -127 56 -121
rect 57 -127 60 -121
rect 64 -127 70 -121
rect 78 -127 81 -121
rect 85 -127 88 -121
rect 92 -127 95 -121
rect 99 -127 105 -121
rect 106 -127 109 -121
rect 113 -127 119 -121
rect 120 -127 123 -121
rect 127 -127 133 -121
rect 134 -127 140 -121
rect 141 -127 147 -121
rect 148 -127 151 -121
rect 155 -127 161 -121
rect 162 -127 168 -121
rect 169 -127 172 -121
rect 176 -127 179 -121
rect 183 -127 189 -121
rect 190 -127 193 -121
rect 197 -127 203 -121
rect 204 -127 207 -121
rect 211 -127 217 -121
rect 218 -127 224 -121
rect 225 -127 228 -121
rect 232 -127 238 -121
rect 239 -127 245 -121
rect 246 -127 252 -121
rect 253 -127 256 -121
rect 260 -127 266 -121
rect 267 -127 273 -121
rect 274 -127 280 -121
rect 281 -127 284 -121
rect 288 -127 291 -121
rect 295 -127 298 -121
rect 302 -127 305 -121
rect 309 -127 315 -121
rect 316 -127 319 -121
rect 323 -127 326 -121
rect 330 -127 333 -121
rect 337 -127 340 -121
rect 344 -127 347 -121
rect 351 -127 354 -121
rect 358 -127 361 -121
rect 365 -127 371 -121
rect 372 -127 375 -121
rect 379 -127 385 -121
rect 386 -127 389 -121
rect 393 -127 396 -121
rect 400 -127 403 -121
rect 407 -127 410 -121
rect 414 -127 417 -121
rect 421 -127 424 -121
rect 428 -127 431 -121
rect 435 -127 441 -121
rect 442 -127 445 -121
rect 449 -127 455 -121
rect 1 -180 7 -174
rect 8 -180 14 -174
rect 15 -180 21 -174
rect 22 -180 28 -174
rect 29 -180 35 -174
rect 36 -180 39 -174
rect 43 -180 46 -174
rect 50 -180 53 -174
rect 57 -180 60 -174
rect 64 -180 70 -174
rect 71 -180 74 -174
rect 78 -180 81 -174
rect 85 -180 91 -174
rect 92 -180 98 -174
rect 99 -180 102 -174
rect 106 -180 112 -174
rect 113 -180 116 -174
rect 120 -180 126 -174
rect 127 -180 130 -174
rect 134 -180 140 -174
rect 141 -180 147 -174
rect 148 -180 154 -174
rect 155 -180 158 -174
rect 162 -180 168 -174
rect 169 -180 172 -174
rect 176 -180 182 -174
rect 183 -180 189 -174
rect 190 -180 193 -174
rect 197 -180 200 -174
rect 204 -180 210 -174
rect 211 -180 217 -174
rect 218 -180 221 -174
rect 225 -180 228 -174
rect 232 -180 238 -174
rect 239 -180 245 -174
rect 246 -180 249 -174
rect 253 -180 259 -174
rect 260 -180 263 -174
rect 267 -180 270 -174
rect 274 -180 280 -174
rect 281 -180 287 -174
rect 288 -180 294 -174
rect 295 -180 301 -174
rect 302 -180 308 -174
rect 309 -180 315 -174
rect 316 -180 322 -174
rect 323 -180 326 -174
rect 330 -180 336 -174
rect 337 -180 340 -174
rect 344 -180 347 -174
rect 351 -180 354 -174
rect 358 -180 361 -174
rect 365 -180 368 -174
rect 372 -180 375 -174
rect 379 -180 382 -174
rect 386 -180 389 -174
rect 393 -180 396 -174
rect 400 -180 403 -174
rect 407 -180 410 -174
rect 414 -180 417 -174
rect 428 -180 431 -174
rect 435 -180 438 -174
rect 442 -180 445 -174
rect 449 -180 452 -174
rect 456 -180 459 -174
rect 463 -180 466 -174
rect 470 -180 473 -174
rect 477 -180 483 -174
rect 484 -180 487 -174
rect 491 -180 494 -174
rect 547 -180 553 -174
rect 1 -237 7 -231
rect 15 -237 18 -231
rect 22 -237 28 -231
rect 29 -237 32 -231
rect 36 -237 42 -231
rect 43 -237 49 -231
rect 57 -237 63 -231
rect 64 -237 70 -231
rect 78 -237 84 -231
rect 85 -237 91 -231
rect 92 -237 95 -231
rect 99 -237 105 -231
rect 106 -237 109 -231
rect 113 -237 116 -231
rect 120 -237 126 -231
rect 127 -237 130 -231
rect 134 -237 137 -231
rect 141 -237 147 -231
rect 148 -237 154 -231
rect 155 -237 161 -231
rect 162 -237 168 -231
rect 169 -237 172 -231
rect 176 -237 179 -231
rect 183 -237 186 -231
rect 190 -237 193 -231
rect 197 -237 200 -231
rect 204 -237 207 -231
rect 211 -237 217 -231
rect 218 -237 224 -231
rect 225 -237 228 -231
rect 232 -237 235 -231
rect 239 -237 245 -231
rect 246 -237 249 -231
rect 253 -237 259 -231
rect 260 -237 263 -231
rect 267 -237 270 -231
rect 274 -237 277 -231
rect 281 -237 287 -231
rect 288 -237 291 -231
rect 302 -237 305 -231
rect 309 -237 315 -231
rect 316 -237 319 -231
rect 323 -237 329 -231
rect 330 -237 333 -231
rect 337 -237 343 -231
rect 344 -237 347 -231
rect 351 -237 357 -231
rect 358 -237 364 -231
rect 365 -237 368 -231
rect 372 -237 375 -231
rect 379 -237 382 -231
rect 386 -237 389 -231
rect 393 -237 396 -231
rect 400 -237 403 -231
rect 407 -237 410 -231
rect 414 -237 417 -231
rect 421 -237 424 -231
rect 428 -237 431 -231
rect 435 -237 438 -231
rect 442 -237 445 -231
rect 449 -237 452 -231
rect 456 -237 459 -231
rect 463 -237 466 -231
rect 470 -237 473 -231
rect 477 -237 480 -231
rect 484 -237 487 -231
rect 491 -237 494 -231
rect 498 -237 501 -231
rect 505 -237 508 -231
rect 512 -237 515 -231
rect 519 -237 525 -231
rect 526 -237 529 -231
rect 533 -237 536 -231
rect 540 -237 546 -231
rect 547 -237 553 -231
rect 554 -237 560 -231
rect 561 -237 567 -231
rect 582 -237 588 -231
rect 638 -237 641 -231
rect 652 -237 658 -231
rect 1 -294 7 -288
rect 8 -294 14 -288
rect 15 -294 21 -288
rect 22 -294 28 -288
rect 29 -294 32 -288
rect 36 -294 42 -288
rect 43 -294 46 -288
rect 50 -294 56 -288
rect 57 -294 60 -288
rect 64 -294 70 -288
rect 71 -294 74 -288
rect 78 -294 84 -288
rect 85 -294 88 -288
rect 92 -294 95 -288
rect 99 -294 102 -288
rect 106 -294 109 -288
rect 113 -294 116 -288
rect 120 -294 126 -288
rect 127 -294 130 -288
rect 134 -294 137 -288
rect 141 -294 147 -288
rect 148 -294 154 -288
rect 155 -294 158 -288
rect 162 -294 168 -288
rect 169 -294 172 -288
rect 176 -294 182 -288
rect 183 -294 186 -288
rect 190 -294 196 -288
rect 197 -294 200 -288
rect 204 -294 210 -288
rect 211 -294 217 -288
rect 218 -294 224 -288
rect 225 -294 228 -288
rect 232 -294 235 -288
rect 239 -294 242 -288
rect 246 -294 252 -288
rect 253 -294 259 -288
rect 260 -294 263 -288
rect 267 -294 270 -288
rect 274 -294 280 -288
rect 281 -294 287 -288
rect 288 -294 291 -288
rect 295 -294 301 -288
rect 302 -294 305 -288
rect 309 -294 315 -288
rect 316 -294 322 -288
rect 323 -294 326 -288
rect 330 -294 336 -288
rect 337 -294 343 -288
rect 344 -294 347 -288
rect 351 -294 354 -288
rect 358 -294 364 -288
rect 365 -294 368 -288
rect 372 -294 375 -288
rect 379 -294 382 -288
rect 386 -294 392 -288
rect 393 -294 396 -288
rect 400 -294 403 -288
rect 407 -294 410 -288
rect 414 -294 417 -288
rect 421 -294 424 -288
rect 428 -294 431 -288
rect 435 -294 441 -288
rect 442 -294 445 -288
rect 449 -294 452 -288
rect 456 -294 459 -288
rect 463 -294 466 -288
rect 470 -294 473 -288
rect 477 -294 483 -288
rect 484 -294 487 -288
rect 491 -294 494 -288
rect 498 -294 501 -288
rect 505 -294 508 -288
rect 512 -294 515 -288
rect 519 -294 522 -288
rect 526 -294 529 -288
rect 533 -294 536 -288
rect 540 -294 543 -288
rect 547 -294 550 -288
rect 554 -294 557 -288
rect 561 -294 564 -288
rect 568 -294 571 -288
rect 575 -294 578 -288
rect 582 -294 585 -288
rect 589 -294 592 -288
rect 596 -294 599 -288
rect 603 -294 606 -288
rect 610 -294 613 -288
rect 617 -294 620 -288
rect 624 -294 627 -288
rect 631 -294 634 -288
rect 652 -294 655 -288
rect 659 -294 662 -288
rect 1 -363 7 -357
rect 8 -363 11 -357
rect 15 -363 21 -357
rect 22 -363 25 -357
rect 29 -363 32 -357
rect 43 -363 49 -357
rect 50 -363 56 -357
rect 57 -363 60 -357
rect 71 -363 74 -357
rect 78 -363 81 -357
rect 85 -363 88 -357
rect 92 -363 95 -357
rect 99 -363 105 -357
rect 106 -363 112 -357
rect 113 -363 119 -357
rect 120 -363 126 -357
rect 127 -363 130 -357
rect 134 -363 137 -357
rect 141 -363 144 -357
rect 148 -363 154 -357
rect 155 -363 161 -357
rect 162 -363 168 -357
rect 169 -363 175 -357
rect 176 -363 182 -357
rect 183 -363 189 -357
rect 190 -363 196 -357
rect 197 -363 200 -357
rect 204 -363 210 -357
rect 211 -363 214 -357
rect 218 -363 224 -357
rect 225 -363 228 -357
rect 232 -363 235 -357
rect 239 -363 242 -357
rect 246 -363 249 -357
rect 253 -363 256 -357
rect 260 -363 263 -357
rect 267 -363 270 -357
rect 274 -363 280 -357
rect 281 -363 287 -357
rect 288 -363 291 -357
rect 295 -363 301 -357
rect 302 -363 305 -357
rect 309 -363 312 -357
rect 316 -363 319 -357
rect 323 -363 329 -357
rect 330 -363 333 -357
rect 337 -363 340 -357
rect 344 -363 347 -357
rect 351 -363 357 -357
rect 358 -363 364 -357
rect 365 -363 371 -357
rect 372 -363 375 -357
rect 379 -363 385 -357
rect 386 -363 392 -357
rect 393 -363 396 -357
rect 400 -363 403 -357
rect 407 -363 410 -357
rect 414 -363 417 -357
rect 421 -363 424 -357
rect 428 -363 434 -357
rect 435 -363 438 -357
rect 442 -363 445 -357
rect 449 -363 455 -357
rect 456 -363 459 -357
rect 463 -363 466 -357
rect 470 -363 473 -357
rect 477 -363 480 -357
rect 484 -363 487 -357
rect 491 -363 494 -357
rect 505 -363 508 -357
rect 512 -363 515 -357
rect 519 -363 522 -357
rect 526 -363 529 -357
rect 533 -363 536 -357
rect 540 -363 543 -357
rect 547 -363 550 -357
rect 554 -363 557 -357
rect 561 -363 564 -357
rect 568 -363 571 -357
rect 575 -363 578 -357
rect 582 -363 585 -357
rect 589 -363 592 -357
rect 596 -363 599 -357
rect 603 -363 606 -357
rect 610 -363 613 -357
rect 617 -363 623 -357
rect 652 -363 658 -357
rect 659 -363 662 -357
rect 666 -363 672 -357
rect 673 -363 676 -357
rect 1 -430 7 -424
rect 8 -430 14 -424
rect 15 -430 18 -424
rect 29 -430 35 -424
rect 36 -430 42 -424
rect 43 -430 46 -424
rect 50 -430 53 -424
rect 57 -430 63 -424
rect 64 -430 67 -424
rect 71 -430 74 -424
rect 78 -430 84 -424
rect 85 -430 88 -424
rect 92 -430 95 -424
rect 99 -430 102 -424
rect 106 -430 109 -424
rect 113 -430 119 -424
rect 120 -430 123 -424
rect 127 -430 130 -424
rect 134 -430 140 -424
rect 141 -430 144 -424
rect 148 -430 151 -424
rect 155 -430 158 -424
rect 162 -430 168 -424
rect 169 -430 175 -424
rect 176 -430 182 -424
rect 183 -430 186 -424
rect 190 -430 196 -424
rect 197 -430 203 -424
rect 204 -430 210 -424
rect 211 -430 217 -424
rect 218 -430 224 -424
rect 225 -430 231 -424
rect 232 -430 238 -424
rect 239 -430 242 -424
rect 246 -430 252 -424
rect 253 -430 259 -424
rect 260 -430 266 -424
rect 267 -430 270 -424
rect 274 -430 277 -424
rect 281 -430 287 -424
rect 288 -430 291 -424
rect 295 -430 298 -424
rect 302 -430 305 -424
rect 309 -430 315 -424
rect 316 -430 322 -424
rect 323 -430 329 -424
rect 330 -430 333 -424
rect 337 -430 343 -424
rect 344 -430 347 -424
rect 351 -430 354 -424
rect 358 -430 364 -424
rect 365 -430 368 -424
rect 372 -430 375 -424
rect 379 -430 385 -424
rect 386 -430 392 -424
rect 393 -430 396 -424
rect 400 -430 403 -424
rect 407 -430 410 -424
rect 414 -430 417 -424
rect 421 -430 424 -424
rect 428 -430 431 -424
rect 435 -430 438 -424
rect 442 -430 445 -424
rect 449 -430 452 -424
rect 456 -430 459 -424
rect 463 -430 466 -424
rect 470 -430 476 -424
rect 477 -430 483 -424
rect 484 -430 487 -424
rect 491 -430 494 -424
rect 498 -430 501 -424
rect 505 -430 508 -424
rect 512 -430 515 -424
rect 519 -430 522 -424
rect 526 -430 529 -424
rect 533 -430 536 -424
rect 540 -430 543 -424
rect 547 -430 550 -424
rect 554 -430 557 -424
rect 561 -430 564 -424
rect 568 -430 571 -424
rect 575 -430 578 -424
rect 582 -430 585 -424
rect 589 -430 592 -424
rect 596 -430 599 -424
rect 603 -430 606 -424
rect 610 -430 613 -424
rect 617 -430 620 -424
rect 624 -430 627 -424
rect 631 -430 634 -424
rect 638 -430 641 -424
rect 645 -430 648 -424
rect 652 -430 655 -424
rect 659 -430 662 -424
rect 666 -430 669 -424
rect 673 -430 679 -424
rect 680 -430 683 -424
rect 1 -517 7 -511
rect 8 -517 14 -511
rect 15 -517 21 -511
rect 22 -517 28 -511
rect 29 -517 35 -511
rect 36 -517 42 -511
rect 43 -517 46 -511
rect 50 -517 56 -511
rect 57 -517 60 -511
rect 64 -517 67 -511
rect 71 -517 74 -511
rect 78 -517 81 -511
rect 85 -517 91 -511
rect 92 -517 95 -511
rect 99 -517 102 -511
rect 106 -517 112 -511
rect 113 -517 116 -511
rect 120 -517 126 -511
rect 127 -517 130 -511
rect 134 -517 137 -511
rect 141 -517 147 -511
rect 148 -517 151 -511
rect 155 -517 158 -511
rect 162 -517 165 -511
rect 169 -517 175 -511
rect 176 -517 179 -511
rect 183 -517 186 -511
rect 190 -517 193 -511
rect 197 -517 203 -511
rect 204 -517 207 -511
rect 211 -517 217 -511
rect 218 -517 224 -511
rect 225 -517 231 -511
rect 232 -517 235 -511
rect 239 -517 245 -511
rect 246 -517 249 -511
rect 253 -517 259 -511
rect 260 -517 263 -511
rect 267 -517 273 -511
rect 274 -517 280 -511
rect 281 -517 287 -511
rect 288 -517 291 -511
rect 295 -517 301 -511
rect 302 -517 305 -511
rect 309 -517 312 -511
rect 316 -517 322 -511
rect 323 -517 329 -511
rect 330 -517 333 -511
rect 337 -517 340 -511
rect 344 -517 350 -511
rect 351 -517 357 -511
rect 358 -517 364 -511
rect 365 -517 368 -511
rect 372 -517 375 -511
rect 379 -517 382 -511
rect 386 -517 392 -511
rect 393 -517 396 -511
rect 400 -517 406 -511
rect 407 -517 410 -511
rect 414 -517 417 -511
rect 421 -517 427 -511
rect 428 -517 431 -511
rect 435 -517 441 -511
rect 442 -517 445 -511
rect 449 -517 455 -511
rect 456 -517 459 -511
rect 463 -517 466 -511
rect 470 -517 473 -511
rect 477 -517 480 -511
rect 484 -517 487 -511
rect 491 -517 494 -511
rect 498 -517 501 -511
rect 505 -517 508 -511
rect 512 -517 515 -511
rect 519 -517 522 -511
rect 526 -517 529 -511
rect 533 -517 536 -511
rect 540 -517 543 -511
rect 547 -517 550 -511
rect 554 -517 557 -511
rect 561 -517 564 -511
rect 568 -517 571 -511
rect 575 -517 578 -511
rect 582 -517 585 -511
rect 589 -517 592 -511
rect 596 -517 599 -511
rect 603 -517 606 -511
rect 610 -517 613 -511
rect 617 -517 620 -511
rect 624 -517 627 -511
rect 631 -517 634 -511
rect 638 -517 641 -511
rect 645 -517 648 -511
rect 652 -517 655 -511
rect 659 -517 662 -511
rect 666 -517 669 -511
rect 673 -517 676 -511
rect 680 -517 683 -511
rect 687 -517 690 -511
rect 694 -517 697 -511
rect 701 -517 704 -511
rect 708 -517 711 -511
rect 1 -604 7 -598
rect 8 -604 14 -598
rect 15 -604 21 -598
rect 22 -604 25 -598
rect 29 -604 32 -598
rect 36 -604 39 -598
rect 43 -604 46 -598
rect 50 -604 56 -598
rect 57 -604 60 -598
rect 64 -604 70 -598
rect 71 -604 77 -598
rect 78 -604 81 -598
rect 85 -604 88 -598
rect 92 -604 95 -598
rect 99 -604 105 -598
rect 106 -604 112 -598
rect 113 -604 119 -598
rect 120 -604 123 -598
rect 127 -604 133 -598
rect 134 -604 140 -598
rect 141 -604 144 -598
rect 148 -604 151 -598
rect 155 -604 161 -598
rect 162 -604 165 -598
rect 169 -604 172 -598
rect 176 -604 179 -598
rect 183 -604 186 -598
rect 190 -604 196 -598
rect 197 -604 203 -598
rect 204 -604 207 -598
rect 211 -604 217 -598
rect 218 -604 224 -598
rect 225 -604 228 -598
rect 232 -604 235 -598
rect 239 -604 242 -598
rect 246 -604 249 -598
rect 253 -604 256 -598
rect 260 -604 263 -598
rect 267 -604 270 -598
rect 274 -604 280 -598
rect 281 -604 287 -598
rect 288 -604 291 -598
rect 295 -604 298 -598
rect 302 -604 308 -598
rect 309 -604 312 -598
rect 316 -604 322 -598
rect 323 -604 326 -598
rect 330 -604 333 -598
rect 337 -604 343 -598
rect 344 -604 350 -598
rect 351 -604 354 -598
rect 358 -604 361 -598
rect 365 -604 368 -598
rect 372 -604 378 -598
rect 379 -604 382 -598
rect 386 -604 389 -598
rect 393 -604 396 -598
rect 400 -604 403 -598
rect 407 -604 413 -598
rect 414 -604 420 -598
rect 421 -604 424 -598
rect 428 -604 431 -598
rect 435 -604 441 -598
rect 442 -604 448 -598
rect 449 -604 452 -598
rect 456 -604 462 -598
rect 463 -604 466 -598
rect 470 -604 476 -598
rect 477 -604 480 -598
rect 484 -604 487 -598
rect 491 -604 497 -598
rect 498 -604 504 -598
rect 505 -604 508 -598
rect 512 -604 515 -598
rect 519 -604 522 -598
rect 526 -604 529 -598
rect 533 -604 536 -598
rect 540 -604 543 -598
rect 547 -604 550 -598
rect 554 -604 560 -598
rect 561 -604 564 -598
rect 568 -604 571 -598
rect 575 -604 578 -598
rect 582 -604 585 -598
rect 589 -604 592 -598
rect 596 -604 599 -598
rect 603 -604 606 -598
rect 610 -604 613 -598
rect 617 -604 620 -598
rect 624 -604 627 -598
rect 631 -604 634 -598
rect 638 -604 641 -598
rect 645 -604 648 -598
rect 652 -604 655 -598
rect 659 -604 662 -598
rect 666 -604 669 -598
rect 673 -604 676 -598
rect 680 -604 683 -598
rect 708 -604 711 -598
rect 1 -683 7 -677
rect 8 -683 14 -677
rect 15 -683 21 -677
rect 22 -683 28 -677
rect 29 -683 35 -677
rect 36 -683 39 -677
rect 43 -683 46 -677
rect 50 -683 53 -677
rect 57 -683 63 -677
rect 64 -683 67 -677
rect 71 -683 77 -677
rect 78 -683 81 -677
rect 85 -683 88 -677
rect 92 -683 95 -677
rect 99 -683 102 -677
rect 106 -683 109 -677
rect 113 -683 116 -677
rect 120 -683 126 -677
rect 127 -683 133 -677
rect 134 -683 140 -677
rect 141 -683 147 -677
rect 148 -683 151 -677
rect 155 -683 161 -677
rect 162 -683 165 -677
rect 169 -683 172 -677
rect 176 -683 179 -677
rect 183 -683 189 -677
rect 190 -683 193 -677
rect 197 -683 203 -677
rect 204 -683 207 -677
rect 211 -683 214 -677
rect 218 -683 224 -677
rect 225 -683 228 -677
rect 232 -683 235 -677
rect 239 -683 242 -677
rect 246 -683 249 -677
rect 253 -683 256 -677
rect 260 -683 263 -677
rect 267 -683 270 -677
rect 274 -683 280 -677
rect 281 -683 287 -677
rect 288 -683 291 -677
rect 295 -683 298 -677
rect 302 -683 305 -677
rect 309 -683 312 -677
rect 316 -683 322 -677
rect 323 -683 329 -677
rect 330 -683 333 -677
rect 337 -683 340 -677
rect 344 -683 350 -677
rect 351 -683 357 -677
rect 358 -683 361 -677
rect 365 -683 368 -677
rect 372 -683 375 -677
rect 379 -683 382 -677
rect 386 -683 389 -677
rect 393 -683 399 -677
rect 400 -683 406 -677
rect 407 -683 410 -677
rect 414 -683 417 -677
rect 421 -683 427 -677
rect 428 -683 431 -677
rect 435 -683 441 -677
rect 442 -683 445 -677
rect 449 -683 455 -677
rect 456 -683 462 -677
rect 463 -683 469 -677
rect 477 -683 483 -677
rect 484 -683 487 -677
rect 491 -683 497 -677
rect 498 -683 501 -677
rect 505 -683 511 -677
rect 512 -683 515 -677
rect 519 -683 522 -677
rect 526 -683 529 -677
rect 533 -683 536 -677
rect 540 -683 543 -677
rect 547 -683 550 -677
rect 554 -683 557 -677
rect 561 -683 564 -677
rect 568 -683 571 -677
rect 575 -683 578 -677
rect 582 -683 588 -677
rect 589 -683 592 -677
rect 596 -683 599 -677
rect 603 -683 606 -677
rect 610 -683 613 -677
rect 617 -683 620 -677
rect 624 -683 627 -677
rect 631 -683 634 -677
rect 638 -683 641 -677
rect 645 -683 648 -677
rect 652 -683 655 -677
rect 659 -683 662 -677
rect 666 -683 669 -677
rect 673 -683 676 -677
rect 680 -683 683 -677
rect 687 -683 690 -677
rect 694 -683 697 -677
rect 701 -683 704 -677
rect 708 -683 711 -677
rect 715 -683 718 -677
rect 722 -683 725 -677
rect 729 -683 732 -677
rect 736 -683 739 -677
rect 743 -683 746 -677
rect 750 -683 753 -677
rect 757 -683 760 -677
rect 764 -683 767 -677
rect 771 -683 774 -677
rect 1 -768 7 -762
rect 15 -768 21 -762
rect 22 -768 28 -762
rect 29 -768 35 -762
rect 36 -768 39 -762
rect 43 -768 46 -762
rect 50 -768 56 -762
rect 57 -768 60 -762
rect 64 -768 67 -762
rect 71 -768 74 -762
rect 78 -768 84 -762
rect 85 -768 91 -762
rect 92 -768 98 -762
rect 99 -768 102 -762
rect 106 -768 109 -762
rect 113 -768 119 -762
rect 120 -768 126 -762
rect 127 -768 133 -762
rect 134 -768 137 -762
rect 141 -768 144 -762
rect 148 -768 154 -762
rect 155 -768 158 -762
rect 162 -768 165 -762
rect 169 -768 172 -762
rect 176 -768 179 -762
rect 183 -768 186 -762
rect 190 -768 193 -762
rect 197 -768 203 -762
rect 204 -768 207 -762
rect 211 -768 214 -762
rect 218 -768 224 -762
rect 225 -768 228 -762
rect 232 -768 235 -762
rect 239 -768 242 -762
rect 246 -768 249 -762
rect 253 -768 256 -762
rect 260 -768 263 -762
rect 267 -768 270 -762
rect 274 -768 277 -762
rect 281 -768 287 -762
rect 288 -768 294 -762
rect 295 -768 298 -762
rect 302 -768 308 -762
rect 309 -768 315 -762
rect 316 -768 322 -762
rect 323 -768 326 -762
rect 330 -768 333 -762
rect 337 -768 340 -762
rect 344 -768 350 -762
rect 351 -768 357 -762
rect 358 -768 364 -762
rect 365 -768 368 -762
rect 372 -768 375 -762
rect 379 -768 385 -762
rect 386 -768 389 -762
rect 393 -768 399 -762
rect 400 -768 403 -762
rect 407 -768 410 -762
rect 414 -768 417 -762
rect 421 -768 424 -762
rect 428 -768 434 -762
rect 435 -768 441 -762
rect 442 -768 448 -762
rect 449 -768 452 -762
rect 456 -768 459 -762
rect 463 -768 466 -762
rect 470 -768 473 -762
rect 477 -768 483 -762
rect 484 -768 490 -762
rect 491 -768 494 -762
rect 498 -768 501 -762
rect 505 -768 508 -762
rect 512 -768 515 -762
rect 519 -768 522 -762
rect 526 -768 529 -762
rect 533 -768 539 -762
rect 540 -768 543 -762
rect 547 -768 550 -762
rect 554 -768 557 -762
rect 561 -768 564 -762
rect 568 -768 571 -762
rect 575 -768 578 -762
rect 582 -768 585 -762
rect 589 -768 592 -762
rect 596 -768 599 -762
rect 603 -768 606 -762
rect 610 -768 613 -762
rect 617 -768 623 -762
rect 624 -768 627 -762
rect 631 -768 634 -762
rect 638 -768 641 -762
rect 645 -768 648 -762
rect 652 -768 655 -762
rect 659 -768 662 -762
rect 666 -768 669 -762
rect 673 -768 676 -762
rect 680 -768 683 -762
rect 687 -768 690 -762
rect 694 -768 697 -762
rect 701 -768 704 -762
rect 708 -768 711 -762
rect 715 -768 718 -762
rect 722 -768 725 -762
rect 729 -768 735 -762
rect 736 -768 739 -762
rect 743 -768 746 -762
rect 750 -768 753 -762
rect 757 -768 760 -762
rect 764 -768 767 -762
rect 771 -768 774 -762
rect 778 -768 781 -762
rect 785 -768 788 -762
rect 792 -768 795 -762
rect 848 -768 851 -762
rect 1 -857 7 -851
rect 8 -857 14 -851
rect 15 -857 21 -851
rect 22 -857 25 -851
rect 29 -857 32 -851
rect 36 -857 42 -851
rect 43 -857 46 -851
rect 50 -857 56 -851
rect 57 -857 60 -851
rect 64 -857 67 -851
rect 71 -857 77 -851
rect 78 -857 81 -851
rect 85 -857 91 -851
rect 92 -857 95 -851
rect 99 -857 105 -851
rect 106 -857 109 -851
rect 113 -857 116 -851
rect 120 -857 123 -851
rect 127 -857 130 -851
rect 134 -857 137 -851
rect 141 -857 147 -851
rect 148 -857 154 -851
rect 155 -857 161 -851
rect 162 -857 168 -851
rect 169 -857 172 -851
rect 176 -857 179 -851
rect 183 -857 186 -851
rect 190 -857 193 -851
rect 197 -857 200 -851
rect 204 -857 207 -851
rect 211 -857 214 -851
rect 218 -857 221 -851
rect 225 -857 228 -851
rect 232 -857 235 -851
rect 239 -857 242 -851
rect 246 -857 252 -851
rect 253 -857 256 -851
rect 260 -857 266 -851
rect 267 -857 270 -851
rect 274 -857 277 -851
rect 281 -857 284 -851
rect 288 -857 291 -851
rect 295 -857 301 -851
rect 302 -857 308 -851
rect 309 -857 312 -851
rect 316 -857 319 -851
rect 323 -857 329 -851
rect 330 -857 336 -851
rect 337 -857 343 -851
rect 344 -857 347 -851
rect 351 -857 354 -851
rect 358 -857 364 -851
rect 365 -857 368 -851
rect 372 -857 375 -851
rect 379 -857 385 -851
rect 386 -857 389 -851
rect 393 -857 399 -851
rect 400 -857 403 -851
rect 407 -857 413 -851
rect 414 -857 417 -851
rect 421 -857 424 -851
rect 428 -857 434 -851
rect 435 -857 441 -851
rect 442 -857 448 -851
rect 449 -857 455 -851
rect 456 -857 462 -851
rect 463 -857 469 -851
rect 470 -857 473 -851
rect 477 -857 480 -851
rect 484 -857 487 -851
rect 491 -857 494 -851
rect 498 -857 501 -851
rect 505 -857 511 -851
rect 512 -857 518 -851
rect 519 -857 522 -851
rect 526 -857 529 -851
rect 533 -857 536 -851
rect 540 -857 543 -851
rect 547 -857 550 -851
rect 554 -857 557 -851
rect 561 -857 564 -851
rect 568 -857 571 -851
rect 575 -857 578 -851
rect 582 -857 585 -851
rect 589 -857 592 -851
rect 596 -857 599 -851
rect 603 -857 606 -851
rect 610 -857 613 -851
rect 617 -857 620 -851
rect 624 -857 627 -851
rect 631 -857 634 -851
rect 638 -857 641 -851
rect 645 -857 648 -851
rect 652 -857 655 -851
rect 659 -857 662 -851
rect 666 -857 669 -851
rect 673 -857 679 -851
rect 680 -857 683 -851
rect 687 -857 690 -851
rect 694 -857 697 -851
rect 701 -857 704 -851
rect 708 -857 711 -851
rect 715 -857 718 -851
rect 722 -857 725 -851
rect 729 -857 732 -851
rect 736 -857 739 -851
rect 743 -857 746 -851
rect 750 -857 753 -851
rect 757 -857 760 -851
rect 764 -857 767 -851
rect 771 -857 774 -851
rect 778 -857 781 -851
rect 785 -857 788 -851
rect 799 -857 802 -851
rect 806 -857 809 -851
rect 813 -857 816 -851
rect 820 -857 823 -851
rect 827 -857 830 -851
rect 834 -857 837 -851
rect 841 -857 844 -851
rect 848 -857 851 -851
rect 855 -857 858 -851
rect 862 -857 865 -851
rect 869 -857 872 -851
rect 939 -857 942 -851
rect 1 -934 7 -928
rect 8 -934 11 -928
rect 15 -934 18 -928
rect 22 -934 25 -928
rect 29 -934 32 -928
rect 36 -934 42 -928
rect 43 -934 46 -928
rect 50 -934 56 -928
rect 57 -934 60 -928
rect 64 -934 70 -928
rect 71 -934 74 -928
rect 78 -934 84 -928
rect 85 -934 88 -928
rect 92 -934 95 -928
rect 99 -934 102 -928
rect 106 -934 109 -928
rect 113 -934 116 -928
rect 120 -934 126 -928
rect 127 -934 130 -928
rect 134 -934 137 -928
rect 141 -934 144 -928
rect 148 -934 154 -928
rect 155 -934 158 -928
rect 162 -934 168 -928
rect 169 -934 172 -928
rect 176 -934 179 -928
rect 183 -934 189 -928
rect 190 -934 193 -928
rect 197 -934 203 -928
rect 204 -934 210 -928
rect 211 -934 217 -928
rect 218 -934 224 -928
rect 225 -934 228 -928
rect 232 -934 235 -928
rect 239 -934 242 -928
rect 246 -934 252 -928
rect 253 -934 256 -928
rect 260 -934 263 -928
rect 267 -934 270 -928
rect 274 -934 280 -928
rect 281 -934 287 -928
rect 288 -934 291 -928
rect 295 -934 301 -928
rect 302 -934 305 -928
rect 309 -934 312 -928
rect 316 -934 319 -928
rect 323 -934 326 -928
rect 330 -934 333 -928
rect 337 -934 343 -928
rect 344 -934 350 -928
rect 351 -934 357 -928
rect 358 -934 361 -928
rect 365 -934 368 -928
rect 372 -934 375 -928
rect 379 -934 382 -928
rect 386 -934 389 -928
rect 393 -934 399 -928
rect 400 -934 406 -928
rect 407 -934 410 -928
rect 414 -934 417 -928
rect 421 -934 424 -928
rect 428 -934 431 -928
rect 435 -934 438 -928
rect 442 -934 448 -928
rect 449 -934 455 -928
rect 456 -934 459 -928
rect 463 -934 469 -928
rect 470 -934 473 -928
rect 477 -934 480 -928
rect 484 -934 487 -928
rect 491 -934 494 -928
rect 498 -934 501 -928
rect 505 -934 511 -928
rect 512 -934 518 -928
rect 519 -934 522 -928
rect 526 -934 529 -928
rect 533 -934 536 -928
rect 540 -934 546 -928
rect 547 -934 553 -928
rect 554 -934 557 -928
rect 561 -934 564 -928
rect 568 -934 571 -928
rect 575 -934 578 -928
rect 582 -934 585 -928
rect 589 -934 595 -928
rect 596 -934 599 -928
rect 603 -934 606 -928
rect 610 -934 613 -928
rect 617 -934 620 -928
rect 624 -934 627 -928
rect 631 -934 634 -928
rect 638 -934 641 -928
rect 645 -934 648 -928
rect 652 -934 655 -928
rect 659 -934 662 -928
rect 666 -934 669 -928
rect 673 -934 676 -928
rect 680 -934 683 -928
rect 687 -934 690 -928
rect 694 -934 697 -928
rect 701 -934 704 -928
rect 708 -934 711 -928
rect 715 -934 718 -928
rect 722 -934 725 -928
rect 729 -934 732 -928
rect 736 -934 739 -928
rect 743 -934 746 -928
rect 750 -934 753 -928
rect 757 -934 760 -928
rect 764 -934 767 -928
rect 771 -934 774 -928
rect 778 -934 781 -928
rect 785 -934 788 -928
rect 792 -934 795 -928
rect 799 -934 802 -928
rect 806 -934 809 -928
rect 813 -934 816 -928
rect 820 -934 823 -928
rect 827 -934 833 -928
rect 834 -934 837 -928
rect 841 -934 844 -928
rect 848 -934 854 -928
rect 1 -1013 4 -1007
rect 8 -1013 11 -1007
rect 15 -1013 21 -1007
rect 22 -1013 25 -1007
rect 29 -1013 35 -1007
rect 36 -1013 39 -1007
rect 43 -1013 46 -1007
rect 50 -1013 53 -1007
rect 57 -1013 63 -1007
rect 64 -1013 67 -1007
rect 71 -1013 74 -1007
rect 78 -1013 81 -1007
rect 85 -1013 88 -1007
rect 92 -1013 95 -1007
rect 99 -1013 105 -1007
rect 106 -1013 109 -1007
rect 113 -1013 119 -1007
rect 120 -1013 126 -1007
rect 127 -1013 133 -1007
rect 134 -1013 137 -1007
rect 141 -1013 144 -1007
rect 148 -1013 151 -1007
rect 155 -1013 158 -1007
rect 162 -1013 165 -1007
rect 169 -1013 175 -1007
rect 176 -1013 179 -1007
rect 183 -1013 186 -1007
rect 190 -1013 196 -1007
rect 197 -1013 203 -1007
rect 204 -1013 207 -1007
rect 211 -1013 214 -1007
rect 218 -1013 224 -1007
rect 225 -1013 228 -1007
rect 232 -1013 235 -1007
rect 239 -1013 242 -1007
rect 246 -1013 249 -1007
rect 253 -1013 256 -1007
rect 260 -1013 263 -1007
rect 267 -1013 273 -1007
rect 274 -1013 277 -1007
rect 281 -1013 284 -1007
rect 288 -1013 291 -1007
rect 295 -1013 298 -1007
rect 302 -1013 305 -1007
rect 309 -1013 315 -1007
rect 316 -1013 319 -1007
rect 323 -1013 326 -1007
rect 330 -1013 336 -1007
rect 337 -1013 343 -1007
rect 344 -1013 347 -1007
rect 351 -1013 354 -1007
rect 358 -1013 361 -1007
rect 365 -1013 371 -1007
rect 372 -1013 378 -1007
rect 379 -1013 382 -1007
rect 386 -1013 392 -1007
rect 393 -1013 399 -1007
rect 400 -1013 406 -1007
rect 407 -1013 413 -1007
rect 414 -1013 417 -1007
rect 421 -1013 427 -1007
rect 428 -1013 434 -1007
rect 435 -1013 441 -1007
rect 442 -1013 445 -1007
rect 449 -1013 452 -1007
rect 456 -1013 459 -1007
rect 463 -1013 466 -1007
rect 470 -1013 476 -1007
rect 477 -1013 483 -1007
rect 484 -1013 487 -1007
rect 491 -1013 494 -1007
rect 498 -1013 504 -1007
rect 505 -1013 511 -1007
rect 512 -1013 518 -1007
rect 519 -1013 522 -1007
rect 526 -1013 529 -1007
rect 533 -1013 536 -1007
rect 540 -1013 543 -1007
rect 547 -1013 550 -1007
rect 554 -1013 560 -1007
rect 561 -1013 564 -1007
rect 568 -1013 571 -1007
rect 575 -1013 578 -1007
rect 589 -1013 592 -1007
rect 596 -1013 599 -1007
rect 603 -1013 606 -1007
rect 610 -1013 613 -1007
rect 617 -1013 620 -1007
rect 624 -1013 627 -1007
rect 631 -1013 634 -1007
rect 638 -1013 641 -1007
rect 645 -1013 648 -1007
rect 652 -1013 655 -1007
rect 659 -1013 662 -1007
rect 666 -1013 669 -1007
rect 673 -1013 676 -1007
rect 680 -1013 683 -1007
rect 687 -1013 690 -1007
rect 694 -1013 697 -1007
rect 701 -1013 704 -1007
rect 708 -1013 711 -1007
rect 715 -1013 718 -1007
rect 722 -1013 725 -1007
rect 729 -1013 732 -1007
rect 736 -1013 739 -1007
rect 743 -1013 746 -1007
rect 750 -1013 753 -1007
rect 757 -1013 760 -1007
rect 764 -1013 767 -1007
rect 771 -1013 774 -1007
rect 778 -1013 781 -1007
rect 785 -1013 788 -1007
rect 792 -1013 795 -1007
rect 799 -1013 802 -1007
rect 806 -1013 809 -1007
rect 813 -1013 816 -1007
rect 820 -1013 823 -1007
rect 827 -1013 830 -1007
rect 834 -1013 837 -1007
rect 841 -1013 844 -1007
rect 848 -1013 851 -1007
rect 855 -1013 861 -1007
rect 862 -1013 865 -1007
rect 869 -1013 875 -1007
rect 897 -1013 900 -1007
rect 1 -1090 7 -1084
rect 8 -1090 14 -1084
rect 15 -1090 18 -1084
rect 22 -1090 25 -1084
rect 29 -1090 32 -1084
rect 36 -1090 39 -1084
rect 43 -1090 46 -1084
rect 50 -1090 56 -1084
rect 57 -1090 60 -1084
rect 64 -1090 70 -1084
rect 71 -1090 74 -1084
rect 78 -1090 84 -1084
rect 85 -1090 88 -1084
rect 92 -1090 98 -1084
rect 99 -1090 105 -1084
rect 106 -1090 109 -1084
rect 113 -1090 116 -1084
rect 120 -1090 123 -1084
rect 127 -1090 130 -1084
rect 134 -1090 140 -1084
rect 141 -1090 144 -1084
rect 148 -1090 154 -1084
rect 155 -1090 161 -1084
rect 162 -1090 168 -1084
rect 169 -1090 172 -1084
rect 176 -1090 179 -1084
rect 183 -1090 186 -1084
rect 190 -1090 193 -1084
rect 197 -1090 203 -1084
rect 204 -1090 207 -1084
rect 211 -1090 214 -1084
rect 218 -1090 224 -1084
rect 225 -1090 228 -1084
rect 232 -1090 235 -1084
rect 239 -1090 245 -1084
rect 246 -1090 252 -1084
rect 253 -1090 256 -1084
rect 260 -1090 263 -1084
rect 267 -1090 270 -1084
rect 274 -1090 280 -1084
rect 281 -1090 284 -1084
rect 288 -1090 291 -1084
rect 295 -1090 298 -1084
rect 302 -1090 305 -1084
rect 309 -1090 312 -1084
rect 316 -1090 319 -1084
rect 323 -1090 326 -1084
rect 330 -1090 333 -1084
rect 337 -1090 340 -1084
rect 344 -1090 350 -1084
rect 351 -1090 357 -1084
rect 358 -1090 361 -1084
rect 365 -1090 368 -1084
rect 372 -1090 375 -1084
rect 379 -1090 382 -1084
rect 386 -1090 392 -1084
rect 393 -1090 396 -1084
rect 400 -1090 403 -1084
rect 407 -1090 410 -1084
rect 414 -1090 417 -1084
rect 421 -1090 424 -1084
rect 428 -1090 431 -1084
rect 435 -1090 438 -1084
rect 442 -1090 448 -1084
rect 449 -1090 455 -1084
rect 456 -1090 459 -1084
rect 463 -1090 469 -1084
rect 470 -1090 473 -1084
rect 477 -1090 480 -1084
rect 484 -1090 487 -1084
rect 491 -1090 497 -1084
rect 498 -1090 501 -1084
rect 505 -1090 508 -1084
rect 512 -1090 515 -1084
rect 519 -1090 522 -1084
rect 526 -1090 532 -1084
rect 533 -1090 539 -1084
rect 540 -1090 543 -1084
rect 547 -1090 553 -1084
rect 554 -1090 560 -1084
rect 561 -1090 567 -1084
rect 568 -1090 574 -1084
rect 575 -1090 578 -1084
rect 582 -1090 585 -1084
rect 589 -1090 592 -1084
rect 596 -1090 599 -1084
rect 603 -1090 609 -1084
rect 610 -1090 613 -1084
rect 617 -1090 620 -1084
rect 624 -1090 627 -1084
rect 631 -1090 634 -1084
rect 638 -1090 644 -1084
rect 645 -1090 648 -1084
rect 652 -1090 655 -1084
rect 659 -1090 662 -1084
rect 666 -1090 669 -1084
rect 673 -1090 676 -1084
rect 680 -1090 683 -1084
rect 687 -1090 690 -1084
rect 694 -1090 697 -1084
rect 701 -1090 704 -1084
rect 708 -1090 711 -1084
rect 715 -1090 718 -1084
rect 722 -1090 725 -1084
rect 729 -1090 732 -1084
rect 736 -1090 739 -1084
rect 743 -1090 746 -1084
rect 750 -1090 753 -1084
rect 757 -1090 760 -1084
rect 764 -1090 767 -1084
rect 771 -1090 774 -1084
rect 778 -1090 781 -1084
rect 785 -1090 788 -1084
rect 792 -1090 795 -1084
rect 799 -1090 802 -1084
rect 806 -1090 809 -1084
rect 813 -1090 816 -1084
rect 820 -1090 823 -1084
rect 827 -1090 830 -1084
rect 834 -1090 837 -1084
rect 841 -1090 844 -1084
rect 848 -1090 851 -1084
rect 855 -1090 858 -1084
rect 862 -1090 865 -1084
rect 869 -1090 872 -1084
rect 876 -1090 879 -1084
rect 883 -1090 886 -1084
rect 890 -1090 893 -1084
rect 897 -1090 900 -1084
rect 904 -1090 907 -1084
rect 911 -1090 914 -1084
rect 918 -1090 921 -1084
rect 925 -1090 931 -1084
rect 939 -1090 942 -1084
rect 1 -1187 7 -1181
rect 8 -1187 11 -1181
rect 15 -1187 18 -1181
rect 22 -1187 28 -1181
rect 29 -1187 32 -1181
rect 36 -1187 39 -1181
rect 43 -1187 46 -1181
rect 50 -1187 53 -1181
rect 57 -1187 60 -1181
rect 64 -1187 67 -1181
rect 71 -1187 77 -1181
rect 78 -1187 81 -1181
rect 85 -1187 88 -1181
rect 92 -1187 98 -1181
rect 99 -1187 105 -1181
rect 106 -1187 109 -1181
rect 113 -1187 116 -1181
rect 120 -1187 126 -1181
rect 127 -1187 130 -1181
rect 134 -1187 140 -1181
rect 141 -1187 144 -1181
rect 148 -1187 154 -1181
rect 155 -1187 158 -1181
rect 162 -1187 165 -1181
rect 169 -1187 175 -1181
rect 176 -1187 179 -1181
rect 183 -1187 186 -1181
rect 190 -1187 193 -1181
rect 197 -1187 203 -1181
rect 204 -1187 207 -1181
rect 211 -1187 217 -1181
rect 218 -1187 224 -1181
rect 225 -1187 228 -1181
rect 232 -1187 235 -1181
rect 239 -1187 242 -1181
rect 246 -1187 249 -1181
rect 253 -1187 256 -1181
rect 260 -1187 263 -1181
rect 267 -1187 270 -1181
rect 274 -1187 277 -1181
rect 281 -1187 287 -1181
rect 288 -1187 291 -1181
rect 295 -1187 298 -1181
rect 302 -1187 305 -1181
rect 309 -1187 312 -1181
rect 316 -1187 322 -1181
rect 323 -1187 326 -1181
rect 330 -1187 333 -1181
rect 337 -1187 340 -1181
rect 344 -1187 347 -1181
rect 351 -1187 357 -1181
rect 358 -1187 364 -1181
rect 365 -1187 368 -1181
rect 372 -1187 375 -1181
rect 379 -1187 382 -1181
rect 386 -1187 389 -1181
rect 393 -1187 396 -1181
rect 400 -1187 403 -1181
rect 407 -1187 413 -1181
rect 414 -1187 417 -1181
rect 421 -1187 427 -1181
rect 428 -1187 431 -1181
rect 435 -1187 438 -1181
rect 442 -1187 445 -1181
rect 449 -1187 455 -1181
rect 456 -1187 459 -1181
rect 463 -1187 469 -1181
rect 470 -1187 473 -1181
rect 477 -1187 483 -1181
rect 484 -1187 487 -1181
rect 491 -1187 494 -1181
rect 498 -1187 501 -1181
rect 505 -1187 511 -1181
rect 512 -1187 515 -1181
rect 519 -1187 522 -1181
rect 526 -1187 529 -1181
rect 533 -1187 536 -1181
rect 540 -1187 546 -1181
rect 547 -1187 550 -1181
rect 554 -1187 557 -1181
rect 561 -1187 564 -1181
rect 568 -1187 571 -1181
rect 575 -1187 581 -1181
rect 582 -1187 585 -1181
rect 589 -1187 592 -1181
rect 596 -1187 599 -1181
rect 603 -1187 606 -1181
rect 610 -1187 613 -1181
rect 617 -1187 623 -1181
rect 624 -1187 627 -1181
rect 631 -1187 634 -1181
rect 638 -1187 641 -1181
rect 645 -1187 648 -1181
rect 652 -1187 658 -1181
rect 659 -1187 662 -1181
rect 666 -1187 669 -1181
rect 673 -1187 676 -1181
rect 680 -1187 686 -1181
rect 687 -1187 690 -1181
rect 694 -1187 697 -1181
rect 701 -1187 704 -1181
rect 708 -1187 711 -1181
rect 715 -1187 721 -1181
rect 722 -1187 725 -1181
rect 729 -1187 732 -1181
rect 736 -1187 739 -1181
rect 743 -1187 746 -1181
rect 750 -1187 753 -1181
rect 757 -1187 760 -1181
rect 764 -1187 767 -1181
rect 771 -1187 774 -1181
rect 778 -1187 781 -1181
rect 785 -1187 788 -1181
rect 792 -1187 795 -1181
rect 799 -1187 802 -1181
rect 806 -1187 809 -1181
rect 813 -1187 816 -1181
rect 820 -1187 823 -1181
rect 827 -1187 830 -1181
rect 834 -1187 837 -1181
rect 841 -1187 844 -1181
rect 848 -1187 851 -1181
rect 855 -1187 858 -1181
rect 862 -1187 865 -1181
rect 869 -1187 872 -1181
rect 876 -1187 879 -1181
rect 883 -1187 886 -1181
rect 890 -1187 893 -1181
rect 897 -1187 900 -1181
rect 904 -1187 907 -1181
rect 911 -1187 914 -1181
rect 918 -1187 921 -1181
rect 925 -1187 928 -1181
rect 932 -1187 935 -1181
rect 939 -1187 942 -1181
rect 946 -1187 949 -1181
rect 953 -1187 959 -1181
rect 960 -1187 966 -1181
rect 967 -1187 973 -1181
rect 974 -1187 977 -1181
rect 981 -1187 987 -1181
rect 988 -1187 991 -1181
rect 1 -1282 7 -1276
rect 8 -1282 14 -1276
rect 15 -1282 18 -1276
rect 22 -1282 28 -1276
rect 29 -1282 32 -1276
rect 36 -1282 42 -1276
rect 43 -1282 46 -1276
rect 50 -1282 53 -1276
rect 57 -1282 60 -1276
rect 64 -1282 67 -1276
rect 71 -1282 74 -1276
rect 78 -1282 81 -1276
rect 85 -1282 88 -1276
rect 92 -1282 98 -1276
rect 99 -1282 102 -1276
rect 106 -1282 112 -1276
rect 113 -1282 116 -1276
rect 120 -1282 123 -1276
rect 127 -1282 133 -1276
rect 134 -1282 137 -1276
rect 141 -1282 144 -1276
rect 148 -1282 151 -1276
rect 155 -1282 158 -1276
rect 162 -1282 165 -1276
rect 169 -1282 175 -1276
rect 176 -1282 179 -1276
rect 183 -1282 189 -1276
rect 190 -1282 193 -1276
rect 197 -1282 200 -1276
rect 204 -1282 207 -1276
rect 211 -1282 217 -1276
rect 218 -1282 224 -1276
rect 225 -1282 228 -1276
rect 232 -1282 235 -1276
rect 239 -1282 242 -1276
rect 246 -1282 249 -1276
rect 253 -1282 256 -1276
rect 260 -1282 263 -1276
rect 267 -1282 270 -1276
rect 274 -1282 277 -1276
rect 281 -1282 284 -1276
rect 288 -1282 291 -1276
rect 295 -1282 298 -1276
rect 302 -1282 308 -1276
rect 309 -1282 315 -1276
rect 316 -1282 319 -1276
rect 323 -1282 326 -1276
rect 330 -1282 333 -1276
rect 337 -1282 343 -1276
rect 344 -1282 347 -1276
rect 351 -1282 354 -1276
rect 358 -1282 364 -1276
rect 365 -1282 368 -1276
rect 372 -1282 375 -1276
rect 379 -1282 385 -1276
rect 386 -1282 389 -1276
rect 393 -1282 396 -1276
rect 400 -1282 403 -1276
rect 407 -1282 413 -1276
rect 414 -1282 417 -1276
rect 421 -1282 424 -1276
rect 428 -1282 431 -1276
rect 435 -1282 438 -1276
rect 442 -1282 448 -1276
rect 449 -1282 452 -1276
rect 456 -1282 462 -1276
rect 463 -1282 469 -1276
rect 470 -1282 476 -1276
rect 477 -1282 480 -1276
rect 484 -1282 487 -1276
rect 491 -1282 497 -1276
rect 498 -1282 504 -1276
rect 505 -1282 511 -1276
rect 512 -1282 515 -1276
rect 519 -1282 522 -1276
rect 526 -1282 529 -1276
rect 533 -1282 536 -1276
rect 540 -1282 543 -1276
rect 547 -1282 550 -1276
rect 554 -1282 557 -1276
rect 561 -1282 564 -1276
rect 568 -1282 574 -1276
rect 575 -1282 578 -1276
rect 582 -1282 585 -1276
rect 589 -1282 592 -1276
rect 596 -1282 602 -1276
rect 603 -1282 609 -1276
rect 610 -1282 613 -1276
rect 617 -1282 623 -1276
rect 624 -1282 627 -1276
rect 631 -1282 637 -1276
rect 638 -1282 641 -1276
rect 645 -1282 648 -1276
rect 652 -1282 658 -1276
rect 659 -1282 662 -1276
rect 666 -1282 672 -1276
rect 673 -1282 676 -1276
rect 680 -1282 683 -1276
rect 687 -1282 690 -1276
rect 694 -1282 697 -1276
rect 701 -1282 704 -1276
rect 708 -1282 711 -1276
rect 715 -1282 718 -1276
rect 722 -1282 725 -1276
rect 729 -1282 732 -1276
rect 736 -1282 739 -1276
rect 743 -1282 746 -1276
rect 750 -1282 753 -1276
rect 757 -1282 760 -1276
rect 764 -1282 767 -1276
rect 771 -1282 774 -1276
rect 778 -1282 781 -1276
rect 785 -1282 788 -1276
rect 792 -1282 795 -1276
rect 799 -1282 802 -1276
rect 806 -1282 809 -1276
rect 813 -1282 816 -1276
rect 820 -1282 823 -1276
rect 827 -1282 830 -1276
rect 834 -1282 837 -1276
rect 841 -1282 844 -1276
rect 848 -1282 851 -1276
rect 855 -1282 858 -1276
rect 862 -1282 865 -1276
rect 869 -1282 872 -1276
rect 876 -1282 879 -1276
rect 883 -1282 886 -1276
rect 890 -1282 893 -1276
rect 897 -1282 900 -1276
rect 904 -1282 907 -1276
rect 911 -1282 914 -1276
rect 918 -1282 921 -1276
rect 925 -1282 928 -1276
rect 932 -1282 935 -1276
rect 939 -1282 945 -1276
rect 946 -1282 949 -1276
rect 953 -1282 956 -1276
rect 960 -1282 963 -1276
rect 967 -1282 970 -1276
rect 974 -1282 977 -1276
rect 981 -1282 984 -1276
rect 988 -1282 991 -1276
rect 995 -1282 998 -1276
rect 1002 -1282 1005 -1276
rect 1009 -1282 1012 -1276
rect 8 -1367 14 -1361
rect 15 -1367 18 -1361
rect 22 -1367 28 -1361
rect 29 -1367 35 -1361
rect 36 -1367 39 -1361
rect 43 -1367 46 -1361
rect 50 -1367 53 -1361
rect 57 -1367 63 -1361
rect 64 -1367 70 -1361
rect 71 -1367 77 -1361
rect 78 -1367 81 -1361
rect 85 -1367 91 -1361
rect 92 -1367 95 -1361
rect 99 -1367 102 -1361
rect 106 -1367 109 -1361
rect 113 -1367 116 -1361
rect 120 -1367 126 -1361
rect 127 -1367 130 -1361
rect 134 -1367 137 -1361
rect 141 -1367 144 -1361
rect 148 -1367 151 -1361
rect 155 -1367 161 -1361
rect 162 -1367 165 -1361
rect 169 -1367 172 -1361
rect 176 -1367 179 -1361
rect 183 -1367 186 -1361
rect 190 -1367 196 -1361
rect 197 -1367 200 -1361
rect 204 -1367 210 -1361
rect 211 -1367 217 -1361
rect 218 -1367 224 -1361
rect 225 -1367 231 -1361
rect 232 -1367 235 -1361
rect 239 -1367 242 -1361
rect 246 -1367 249 -1361
rect 253 -1367 256 -1361
rect 260 -1367 263 -1361
rect 267 -1367 270 -1361
rect 274 -1367 277 -1361
rect 281 -1367 284 -1361
rect 288 -1367 291 -1361
rect 295 -1367 298 -1361
rect 302 -1367 305 -1361
rect 309 -1367 312 -1361
rect 316 -1367 319 -1361
rect 323 -1367 326 -1361
rect 330 -1367 336 -1361
rect 337 -1367 340 -1361
rect 344 -1367 350 -1361
rect 351 -1367 354 -1361
rect 358 -1367 361 -1361
rect 365 -1367 368 -1361
rect 372 -1367 378 -1361
rect 379 -1367 385 -1361
rect 386 -1367 389 -1361
rect 393 -1367 399 -1361
rect 400 -1367 403 -1361
rect 407 -1367 410 -1361
rect 414 -1367 417 -1361
rect 421 -1367 424 -1361
rect 428 -1367 434 -1361
rect 435 -1367 438 -1361
rect 442 -1367 445 -1361
rect 449 -1367 455 -1361
rect 456 -1367 459 -1361
rect 463 -1367 469 -1361
rect 470 -1367 473 -1361
rect 477 -1367 483 -1361
rect 484 -1367 490 -1361
rect 491 -1367 494 -1361
rect 498 -1367 501 -1361
rect 505 -1367 508 -1361
rect 512 -1367 518 -1361
rect 519 -1367 522 -1361
rect 526 -1367 532 -1361
rect 533 -1367 536 -1361
rect 540 -1367 543 -1361
rect 547 -1367 550 -1361
rect 554 -1367 557 -1361
rect 561 -1367 564 -1361
rect 568 -1367 571 -1361
rect 575 -1367 581 -1361
rect 582 -1367 585 -1361
rect 589 -1367 592 -1361
rect 596 -1367 599 -1361
rect 603 -1367 609 -1361
rect 610 -1367 613 -1361
rect 617 -1367 620 -1361
rect 624 -1367 627 -1361
rect 631 -1367 634 -1361
rect 638 -1367 641 -1361
rect 645 -1367 648 -1361
rect 652 -1367 655 -1361
rect 659 -1367 662 -1361
rect 666 -1367 669 -1361
rect 673 -1367 676 -1361
rect 680 -1367 683 -1361
rect 687 -1367 690 -1361
rect 694 -1367 697 -1361
rect 701 -1367 704 -1361
rect 708 -1367 711 -1361
rect 715 -1367 718 -1361
rect 722 -1367 725 -1361
rect 729 -1367 732 -1361
rect 736 -1367 739 -1361
rect 743 -1367 746 -1361
rect 750 -1367 753 -1361
rect 757 -1367 760 -1361
rect 764 -1367 767 -1361
rect 771 -1367 774 -1361
rect 778 -1367 781 -1361
rect 785 -1367 788 -1361
rect 792 -1367 795 -1361
rect 799 -1367 802 -1361
rect 806 -1367 809 -1361
rect 813 -1367 816 -1361
rect 820 -1367 823 -1361
rect 827 -1367 830 -1361
rect 834 -1367 837 -1361
rect 841 -1367 844 -1361
rect 848 -1367 851 -1361
rect 855 -1367 858 -1361
rect 862 -1367 865 -1361
rect 869 -1367 872 -1361
rect 876 -1367 879 -1361
rect 883 -1367 886 -1361
rect 890 -1367 893 -1361
rect 897 -1367 900 -1361
rect 904 -1367 910 -1361
rect 911 -1367 914 -1361
rect 918 -1367 924 -1361
rect 939 -1367 945 -1361
rect 953 -1367 956 -1361
rect 967 -1367 973 -1361
rect 988 -1367 991 -1361
rect 1 -1446 4 -1440
rect 8 -1446 14 -1440
rect 15 -1446 18 -1440
rect 22 -1446 25 -1440
rect 29 -1446 32 -1440
rect 36 -1446 39 -1440
rect 50 -1446 53 -1440
rect 57 -1446 60 -1440
rect 64 -1446 67 -1440
rect 71 -1446 74 -1440
rect 78 -1446 81 -1440
rect 85 -1446 88 -1440
rect 92 -1446 95 -1440
rect 99 -1446 102 -1440
rect 106 -1446 109 -1440
rect 113 -1446 119 -1440
rect 120 -1446 126 -1440
rect 127 -1446 133 -1440
rect 134 -1446 137 -1440
rect 141 -1446 147 -1440
rect 148 -1446 151 -1440
rect 155 -1446 161 -1440
rect 162 -1446 168 -1440
rect 169 -1446 172 -1440
rect 176 -1446 179 -1440
rect 183 -1446 189 -1440
rect 190 -1446 193 -1440
rect 197 -1446 200 -1440
rect 204 -1446 207 -1440
rect 211 -1446 217 -1440
rect 218 -1446 221 -1440
rect 225 -1446 228 -1440
rect 232 -1446 235 -1440
rect 239 -1446 242 -1440
rect 246 -1446 249 -1440
rect 253 -1446 256 -1440
rect 260 -1446 263 -1440
rect 267 -1446 270 -1440
rect 274 -1446 277 -1440
rect 281 -1446 284 -1440
rect 288 -1446 291 -1440
rect 295 -1446 298 -1440
rect 302 -1446 305 -1440
rect 309 -1446 312 -1440
rect 316 -1446 319 -1440
rect 323 -1446 329 -1440
rect 330 -1446 333 -1440
rect 337 -1446 343 -1440
rect 344 -1446 347 -1440
rect 351 -1446 357 -1440
rect 358 -1446 361 -1440
rect 365 -1446 368 -1440
rect 372 -1446 378 -1440
rect 379 -1446 382 -1440
rect 386 -1446 392 -1440
rect 393 -1446 399 -1440
rect 400 -1446 403 -1440
rect 407 -1446 410 -1440
rect 414 -1446 417 -1440
rect 421 -1446 424 -1440
rect 428 -1446 434 -1440
rect 435 -1446 438 -1440
rect 442 -1446 445 -1440
rect 449 -1446 455 -1440
rect 456 -1446 462 -1440
rect 463 -1446 469 -1440
rect 470 -1446 473 -1440
rect 477 -1446 480 -1440
rect 484 -1446 490 -1440
rect 491 -1446 494 -1440
rect 498 -1446 501 -1440
rect 505 -1446 511 -1440
rect 512 -1446 515 -1440
rect 519 -1446 522 -1440
rect 526 -1446 529 -1440
rect 533 -1446 539 -1440
rect 540 -1446 543 -1440
rect 547 -1446 553 -1440
rect 554 -1446 560 -1440
rect 561 -1446 564 -1440
rect 568 -1446 571 -1440
rect 575 -1446 581 -1440
rect 582 -1446 585 -1440
rect 589 -1446 595 -1440
rect 596 -1446 599 -1440
rect 603 -1446 609 -1440
rect 610 -1446 613 -1440
rect 617 -1446 620 -1440
rect 624 -1446 627 -1440
rect 631 -1446 637 -1440
rect 638 -1446 641 -1440
rect 645 -1446 648 -1440
rect 652 -1446 658 -1440
rect 659 -1446 662 -1440
rect 666 -1446 669 -1440
rect 673 -1446 676 -1440
rect 680 -1446 683 -1440
rect 687 -1446 690 -1440
rect 694 -1446 697 -1440
rect 701 -1446 704 -1440
rect 708 -1446 714 -1440
rect 715 -1446 718 -1440
rect 722 -1446 725 -1440
rect 729 -1446 732 -1440
rect 736 -1446 739 -1440
rect 743 -1446 746 -1440
rect 750 -1446 753 -1440
rect 757 -1446 760 -1440
rect 764 -1446 767 -1440
rect 771 -1446 774 -1440
rect 778 -1446 781 -1440
rect 785 -1446 788 -1440
rect 792 -1446 795 -1440
rect 799 -1446 802 -1440
rect 806 -1446 809 -1440
rect 813 -1446 816 -1440
rect 820 -1446 823 -1440
rect 834 -1446 837 -1440
rect 841 -1446 844 -1440
rect 848 -1446 851 -1440
rect 855 -1446 858 -1440
rect 862 -1446 865 -1440
rect 869 -1446 872 -1440
rect 876 -1446 879 -1440
rect 883 -1446 886 -1440
rect 890 -1446 893 -1440
rect 897 -1446 900 -1440
rect 904 -1446 907 -1440
rect 911 -1446 914 -1440
rect 918 -1446 921 -1440
rect 925 -1446 928 -1440
rect 932 -1446 935 -1440
rect 939 -1446 945 -1440
rect 946 -1446 952 -1440
rect 953 -1446 956 -1440
rect 967 -1446 970 -1440
rect 981 -1446 984 -1440
rect 8 -1535 11 -1529
rect 15 -1535 18 -1529
rect 22 -1535 28 -1529
rect 29 -1535 32 -1529
rect 36 -1535 42 -1529
rect 43 -1535 46 -1529
rect 50 -1535 53 -1529
rect 57 -1535 60 -1529
rect 64 -1535 67 -1529
rect 71 -1535 77 -1529
rect 78 -1535 81 -1529
rect 85 -1535 88 -1529
rect 92 -1535 95 -1529
rect 99 -1535 102 -1529
rect 106 -1535 109 -1529
rect 113 -1535 116 -1529
rect 120 -1535 123 -1529
rect 127 -1535 130 -1529
rect 134 -1535 140 -1529
rect 141 -1535 144 -1529
rect 148 -1535 154 -1529
rect 155 -1535 161 -1529
rect 162 -1535 168 -1529
rect 169 -1535 175 -1529
rect 176 -1535 182 -1529
rect 183 -1535 189 -1529
rect 190 -1535 196 -1529
rect 197 -1535 203 -1529
rect 204 -1535 207 -1529
rect 211 -1535 217 -1529
rect 218 -1535 224 -1529
rect 225 -1535 228 -1529
rect 232 -1535 235 -1529
rect 239 -1535 242 -1529
rect 246 -1535 249 -1529
rect 253 -1535 256 -1529
rect 260 -1535 263 -1529
rect 267 -1535 270 -1529
rect 274 -1535 277 -1529
rect 281 -1535 287 -1529
rect 288 -1535 291 -1529
rect 295 -1535 298 -1529
rect 302 -1535 308 -1529
rect 309 -1535 312 -1529
rect 316 -1535 319 -1529
rect 323 -1535 326 -1529
rect 330 -1535 333 -1529
rect 337 -1535 340 -1529
rect 344 -1535 347 -1529
rect 351 -1535 354 -1529
rect 358 -1535 364 -1529
rect 365 -1535 371 -1529
rect 372 -1535 375 -1529
rect 379 -1535 382 -1529
rect 386 -1535 389 -1529
rect 393 -1535 396 -1529
rect 400 -1535 403 -1529
rect 407 -1535 413 -1529
rect 414 -1535 417 -1529
rect 421 -1535 424 -1529
rect 428 -1535 434 -1529
rect 435 -1535 438 -1529
rect 442 -1535 448 -1529
rect 449 -1535 455 -1529
rect 456 -1535 459 -1529
rect 463 -1535 469 -1529
rect 470 -1535 473 -1529
rect 477 -1535 483 -1529
rect 484 -1535 487 -1529
rect 491 -1535 494 -1529
rect 498 -1535 504 -1529
rect 505 -1535 511 -1529
rect 512 -1535 515 -1529
rect 519 -1535 522 -1529
rect 526 -1535 529 -1529
rect 533 -1535 539 -1529
rect 540 -1535 543 -1529
rect 547 -1535 550 -1529
rect 554 -1535 560 -1529
rect 561 -1535 564 -1529
rect 568 -1535 571 -1529
rect 575 -1535 578 -1529
rect 582 -1535 585 -1529
rect 589 -1535 592 -1529
rect 596 -1535 599 -1529
rect 603 -1535 606 -1529
rect 610 -1535 613 -1529
rect 617 -1535 620 -1529
rect 624 -1535 627 -1529
rect 631 -1535 634 -1529
rect 638 -1535 641 -1529
rect 645 -1535 648 -1529
rect 652 -1535 655 -1529
rect 659 -1535 662 -1529
rect 666 -1535 669 -1529
rect 673 -1535 676 -1529
rect 680 -1535 683 -1529
rect 687 -1535 690 -1529
rect 694 -1535 697 -1529
rect 701 -1535 704 -1529
rect 708 -1535 711 -1529
rect 715 -1535 718 -1529
rect 722 -1535 725 -1529
rect 729 -1535 732 -1529
rect 736 -1535 739 -1529
rect 743 -1535 746 -1529
rect 750 -1535 753 -1529
rect 764 -1535 767 -1529
rect 771 -1535 774 -1529
rect 778 -1535 781 -1529
rect 785 -1535 788 -1529
rect 792 -1535 795 -1529
rect 799 -1535 802 -1529
rect 806 -1535 809 -1529
rect 813 -1535 816 -1529
rect 820 -1535 823 -1529
rect 827 -1535 830 -1529
rect 834 -1535 837 -1529
rect 841 -1535 844 -1529
rect 848 -1535 851 -1529
rect 855 -1535 858 -1529
rect 883 -1535 889 -1529
rect 890 -1535 893 -1529
rect 897 -1535 900 -1529
rect 904 -1535 907 -1529
rect 911 -1535 914 -1529
rect 918 -1535 921 -1529
rect 932 -1535 938 -1529
rect 939 -1535 942 -1529
rect 953 -1535 956 -1529
rect 960 -1535 966 -1529
rect 981 -1535 987 -1529
rect 988 -1535 991 -1529
rect 8 -1620 14 -1614
rect 15 -1620 18 -1614
rect 22 -1620 25 -1614
rect 29 -1620 32 -1614
rect 36 -1620 39 -1614
rect 43 -1620 46 -1614
rect 50 -1620 53 -1614
rect 57 -1620 63 -1614
rect 64 -1620 67 -1614
rect 71 -1620 74 -1614
rect 78 -1620 81 -1614
rect 85 -1620 88 -1614
rect 92 -1620 98 -1614
rect 99 -1620 102 -1614
rect 106 -1620 112 -1614
rect 120 -1620 126 -1614
rect 127 -1620 130 -1614
rect 134 -1620 137 -1614
rect 141 -1620 144 -1614
rect 148 -1620 151 -1614
rect 155 -1620 161 -1614
rect 162 -1620 168 -1614
rect 169 -1620 175 -1614
rect 176 -1620 179 -1614
rect 183 -1620 189 -1614
rect 190 -1620 196 -1614
rect 197 -1620 200 -1614
rect 204 -1620 210 -1614
rect 211 -1620 214 -1614
rect 218 -1620 221 -1614
rect 225 -1620 228 -1614
rect 232 -1620 235 -1614
rect 239 -1620 242 -1614
rect 246 -1620 249 -1614
rect 253 -1620 256 -1614
rect 260 -1620 263 -1614
rect 267 -1620 270 -1614
rect 274 -1620 277 -1614
rect 281 -1620 284 -1614
rect 288 -1620 294 -1614
rect 295 -1620 298 -1614
rect 302 -1620 305 -1614
rect 309 -1620 312 -1614
rect 316 -1620 319 -1614
rect 323 -1620 326 -1614
rect 330 -1620 333 -1614
rect 337 -1620 343 -1614
rect 344 -1620 350 -1614
rect 351 -1620 354 -1614
rect 358 -1620 364 -1614
rect 365 -1620 368 -1614
rect 372 -1620 375 -1614
rect 379 -1620 385 -1614
rect 386 -1620 389 -1614
rect 393 -1620 396 -1614
rect 400 -1620 403 -1614
rect 407 -1620 410 -1614
rect 414 -1620 417 -1614
rect 421 -1620 427 -1614
rect 428 -1620 431 -1614
rect 435 -1620 438 -1614
rect 442 -1620 445 -1614
rect 449 -1620 455 -1614
rect 456 -1620 459 -1614
rect 463 -1620 466 -1614
rect 470 -1620 473 -1614
rect 477 -1620 483 -1614
rect 484 -1620 487 -1614
rect 491 -1620 497 -1614
rect 498 -1620 501 -1614
rect 505 -1620 508 -1614
rect 512 -1620 515 -1614
rect 519 -1620 522 -1614
rect 526 -1620 532 -1614
rect 533 -1620 539 -1614
rect 540 -1620 543 -1614
rect 547 -1620 550 -1614
rect 554 -1620 557 -1614
rect 561 -1620 567 -1614
rect 568 -1620 571 -1614
rect 575 -1620 578 -1614
rect 582 -1620 588 -1614
rect 589 -1620 592 -1614
rect 596 -1620 599 -1614
rect 603 -1620 606 -1614
rect 610 -1620 613 -1614
rect 624 -1620 627 -1614
rect 631 -1620 634 -1614
rect 638 -1620 641 -1614
rect 645 -1620 648 -1614
rect 652 -1620 655 -1614
rect 659 -1620 662 -1614
rect 666 -1620 672 -1614
rect 673 -1620 676 -1614
rect 680 -1620 683 -1614
rect 687 -1620 690 -1614
rect 694 -1620 697 -1614
rect 701 -1620 707 -1614
rect 708 -1620 711 -1614
rect 715 -1620 718 -1614
rect 722 -1620 725 -1614
rect 729 -1620 735 -1614
rect 743 -1620 746 -1614
rect 750 -1620 753 -1614
rect 757 -1620 760 -1614
rect 764 -1620 767 -1614
rect 785 -1620 788 -1614
rect 792 -1620 795 -1614
rect 799 -1620 802 -1614
rect 813 -1620 816 -1614
rect 827 -1620 830 -1614
rect 841 -1620 844 -1614
rect 848 -1620 854 -1614
rect 855 -1620 858 -1614
rect 869 -1620 872 -1614
rect 876 -1620 882 -1614
rect 897 -1620 900 -1614
rect 911 -1620 917 -1614
rect 918 -1620 921 -1614
rect 925 -1620 928 -1614
rect 939 -1620 945 -1614
rect 946 -1620 949 -1614
rect 953 -1620 956 -1614
rect 967 -1620 973 -1614
rect 974 -1620 977 -1614
rect 981 -1620 984 -1614
rect 8 -1713 11 -1707
rect 15 -1713 21 -1707
rect 22 -1713 25 -1707
rect 29 -1713 32 -1707
rect 36 -1713 39 -1707
rect 43 -1713 46 -1707
rect 50 -1713 53 -1707
rect 57 -1713 63 -1707
rect 64 -1713 67 -1707
rect 71 -1713 77 -1707
rect 78 -1713 81 -1707
rect 85 -1713 88 -1707
rect 92 -1713 95 -1707
rect 99 -1713 105 -1707
rect 106 -1713 109 -1707
rect 113 -1713 119 -1707
rect 120 -1713 123 -1707
rect 127 -1713 130 -1707
rect 134 -1713 137 -1707
rect 141 -1713 147 -1707
rect 148 -1713 154 -1707
rect 155 -1713 158 -1707
rect 162 -1713 165 -1707
rect 169 -1713 175 -1707
rect 176 -1713 182 -1707
rect 183 -1713 186 -1707
rect 190 -1713 193 -1707
rect 197 -1713 200 -1707
rect 204 -1713 210 -1707
rect 211 -1713 214 -1707
rect 218 -1713 221 -1707
rect 225 -1713 228 -1707
rect 232 -1713 238 -1707
rect 239 -1713 242 -1707
rect 246 -1713 249 -1707
rect 253 -1713 256 -1707
rect 260 -1713 263 -1707
rect 267 -1713 270 -1707
rect 274 -1713 277 -1707
rect 281 -1713 284 -1707
rect 288 -1713 291 -1707
rect 295 -1713 301 -1707
rect 302 -1713 305 -1707
rect 309 -1713 312 -1707
rect 316 -1713 319 -1707
rect 323 -1713 326 -1707
rect 330 -1713 336 -1707
rect 337 -1713 343 -1707
rect 344 -1713 347 -1707
rect 351 -1713 354 -1707
rect 358 -1713 361 -1707
rect 365 -1713 368 -1707
rect 372 -1713 378 -1707
rect 379 -1713 382 -1707
rect 386 -1713 392 -1707
rect 393 -1713 399 -1707
rect 400 -1713 406 -1707
rect 407 -1713 410 -1707
rect 414 -1713 417 -1707
rect 421 -1713 424 -1707
rect 428 -1713 431 -1707
rect 435 -1713 441 -1707
rect 442 -1713 445 -1707
rect 449 -1713 455 -1707
rect 456 -1713 459 -1707
rect 463 -1713 469 -1707
rect 470 -1713 473 -1707
rect 477 -1713 480 -1707
rect 484 -1713 490 -1707
rect 491 -1713 494 -1707
rect 498 -1713 501 -1707
rect 505 -1713 511 -1707
rect 512 -1713 515 -1707
rect 519 -1713 522 -1707
rect 526 -1713 529 -1707
rect 533 -1713 536 -1707
rect 540 -1713 546 -1707
rect 547 -1713 550 -1707
rect 554 -1713 557 -1707
rect 561 -1713 564 -1707
rect 568 -1713 574 -1707
rect 575 -1713 578 -1707
rect 582 -1713 585 -1707
rect 589 -1713 592 -1707
rect 596 -1713 599 -1707
rect 603 -1713 606 -1707
rect 610 -1713 613 -1707
rect 617 -1713 620 -1707
rect 624 -1713 627 -1707
rect 631 -1713 634 -1707
rect 638 -1713 641 -1707
rect 645 -1713 648 -1707
rect 652 -1713 655 -1707
rect 659 -1713 665 -1707
rect 666 -1713 669 -1707
rect 673 -1713 676 -1707
rect 680 -1713 683 -1707
rect 687 -1713 690 -1707
rect 694 -1713 697 -1707
rect 701 -1713 704 -1707
rect 708 -1713 714 -1707
rect 715 -1713 718 -1707
rect 722 -1713 725 -1707
rect 729 -1713 732 -1707
rect 736 -1713 739 -1707
rect 743 -1713 746 -1707
rect 750 -1713 753 -1707
rect 757 -1713 760 -1707
rect 764 -1713 767 -1707
rect 771 -1713 774 -1707
rect 778 -1713 781 -1707
rect 785 -1713 788 -1707
rect 799 -1713 802 -1707
rect 813 -1713 816 -1707
rect 820 -1713 823 -1707
rect 827 -1713 830 -1707
rect 834 -1713 837 -1707
rect 841 -1713 844 -1707
rect 862 -1713 865 -1707
rect 869 -1713 872 -1707
rect 883 -1713 889 -1707
rect 890 -1713 896 -1707
rect 911 -1713 914 -1707
rect 925 -1713 928 -1707
rect 939 -1713 945 -1707
rect 960 -1713 963 -1707
rect 967 -1713 973 -1707
rect 974 -1713 980 -1707
rect 8 -1808 14 -1802
rect 15 -1808 18 -1802
rect 22 -1808 25 -1802
rect 29 -1808 32 -1802
rect 36 -1808 42 -1802
rect 43 -1808 46 -1802
rect 50 -1808 56 -1802
rect 57 -1808 60 -1802
rect 64 -1808 67 -1802
rect 71 -1808 74 -1802
rect 78 -1808 84 -1802
rect 85 -1808 91 -1802
rect 92 -1808 95 -1802
rect 99 -1808 105 -1802
rect 106 -1808 109 -1802
rect 113 -1808 119 -1802
rect 120 -1808 126 -1802
rect 127 -1808 133 -1802
rect 134 -1808 140 -1802
rect 141 -1808 144 -1802
rect 148 -1808 151 -1802
rect 155 -1808 161 -1802
rect 162 -1808 168 -1802
rect 169 -1808 175 -1802
rect 176 -1808 182 -1802
rect 183 -1808 189 -1802
rect 190 -1808 193 -1802
rect 197 -1808 200 -1802
rect 204 -1808 207 -1802
rect 211 -1808 217 -1802
rect 218 -1808 224 -1802
rect 225 -1808 228 -1802
rect 232 -1808 235 -1802
rect 239 -1808 242 -1802
rect 246 -1808 249 -1802
rect 253 -1808 256 -1802
rect 260 -1808 263 -1802
rect 267 -1808 273 -1802
rect 274 -1808 277 -1802
rect 281 -1808 284 -1802
rect 288 -1808 291 -1802
rect 295 -1808 298 -1802
rect 302 -1808 305 -1802
rect 309 -1808 312 -1802
rect 316 -1808 322 -1802
rect 323 -1808 326 -1802
rect 330 -1808 333 -1802
rect 337 -1808 340 -1802
rect 344 -1808 347 -1802
rect 351 -1808 357 -1802
rect 358 -1808 361 -1802
rect 365 -1808 371 -1802
rect 372 -1808 378 -1802
rect 379 -1808 385 -1802
rect 386 -1808 389 -1802
rect 393 -1808 399 -1802
rect 400 -1808 403 -1802
rect 407 -1808 410 -1802
rect 414 -1808 417 -1802
rect 421 -1808 424 -1802
rect 428 -1808 431 -1802
rect 435 -1808 438 -1802
rect 442 -1808 445 -1802
rect 449 -1808 452 -1802
rect 456 -1808 459 -1802
rect 463 -1808 466 -1802
rect 470 -1808 476 -1802
rect 477 -1808 480 -1802
rect 484 -1808 487 -1802
rect 491 -1808 497 -1802
rect 498 -1808 504 -1802
rect 505 -1808 511 -1802
rect 512 -1808 518 -1802
rect 519 -1808 525 -1802
rect 526 -1808 529 -1802
rect 533 -1808 536 -1802
rect 540 -1808 543 -1802
rect 547 -1808 550 -1802
rect 554 -1808 557 -1802
rect 561 -1808 564 -1802
rect 568 -1808 571 -1802
rect 575 -1808 578 -1802
rect 582 -1808 585 -1802
rect 589 -1808 592 -1802
rect 596 -1808 599 -1802
rect 603 -1808 606 -1802
rect 610 -1808 613 -1802
rect 617 -1808 620 -1802
rect 624 -1808 627 -1802
rect 631 -1808 634 -1802
rect 638 -1808 644 -1802
rect 645 -1808 648 -1802
rect 652 -1808 655 -1802
rect 659 -1808 662 -1802
rect 666 -1808 669 -1802
rect 673 -1808 676 -1802
rect 680 -1808 683 -1802
rect 687 -1808 690 -1802
rect 694 -1808 697 -1802
rect 701 -1808 704 -1802
rect 708 -1808 711 -1802
rect 715 -1808 718 -1802
rect 722 -1808 725 -1802
rect 729 -1808 732 -1802
rect 736 -1808 739 -1802
rect 743 -1808 746 -1802
rect 750 -1808 753 -1802
rect 757 -1808 760 -1802
rect 904 -1808 910 -1802
rect 1 -1889 7 -1883
rect 8 -1889 14 -1883
rect 15 -1889 18 -1883
rect 22 -1889 28 -1883
rect 29 -1889 35 -1883
rect 36 -1889 39 -1883
rect 43 -1889 49 -1883
rect 50 -1889 53 -1883
rect 57 -1889 60 -1883
rect 64 -1889 67 -1883
rect 71 -1889 74 -1883
rect 78 -1889 81 -1883
rect 85 -1889 88 -1883
rect 92 -1889 95 -1883
rect 99 -1889 102 -1883
rect 106 -1889 109 -1883
rect 113 -1889 116 -1883
rect 120 -1889 123 -1883
rect 127 -1889 133 -1883
rect 134 -1889 137 -1883
rect 141 -1889 147 -1883
rect 148 -1889 154 -1883
rect 155 -1889 158 -1883
rect 162 -1889 168 -1883
rect 169 -1889 175 -1883
rect 176 -1889 179 -1883
rect 183 -1889 186 -1883
rect 190 -1889 196 -1883
rect 197 -1889 203 -1883
rect 204 -1889 207 -1883
rect 211 -1889 214 -1883
rect 218 -1889 221 -1883
rect 225 -1889 231 -1883
rect 232 -1889 235 -1883
rect 239 -1889 242 -1883
rect 246 -1889 249 -1883
rect 253 -1889 256 -1883
rect 260 -1889 263 -1883
rect 267 -1889 270 -1883
rect 274 -1889 277 -1883
rect 281 -1889 284 -1883
rect 288 -1889 294 -1883
rect 295 -1889 298 -1883
rect 302 -1889 308 -1883
rect 309 -1889 312 -1883
rect 316 -1889 319 -1883
rect 323 -1889 329 -1883
rect 330 -1889 333 -1883
rect 337 -1889 343 -1883
rect 344 -1889 350 -1883
rect 351 -1889 357 -1883
rect 358 -1889 364 -1883
rect 365 -1889 368 -1883
rect 372 -1889 378 -1883
rect 379 -1889 382 -1883
rect 386 -1889 392 -1883
rect 393 -1889 396 -1883
rect 400 -1889 403 -1883
rect 407 -1889 410 -1883
rect 414 -1889 417 -1883
rect 421 -1889 424 -1883
rect 428 -1889 431 -1883
rect 435 -1889 441 -1883
rect 442 -1889 448 -1883
rect 449 -1889 455 -1883
rect 456 -1889 459 -1883
rect 463 -1889 469 -1883
rect 470 -1889 473 -1883
rect 477 -1889 480 -1883
rect 484 -1889 487 -1883
rect 491 -1889 494 -1883
rect 498 -1889 504 -1883
rect 505 -1889 508 -1883
rect 512 -1889 515 -1883
rect 519 -1889 522 -1883
rect 526 -1889 529 -1883
rect 533 -1889 536 -1883
rect 540 -1889 543 -1883
rect 547 -1889 553 -1883
rect 554 -1889 557 -1883
rect 561 -1889 564 -1883
rect 568 -1889 571 -1883
rect 575 -1889 581 -1883
rect 582 -1889 585 -1883
rect 589 -1889 592 -1883
rect 596 -1889 599 -1883
rect 603 -1889 606 -1883
rect 610 -1889 613 -1883
rect 617 -1889 620 -1883
rect 624 -1889 627 -1883
rect 631 -1889 634 -1883
rect 638 -1889 644 -1883
rect 645 -1889 648 -1883
rect 652 -1889 655 -1883
rect 659 -1889 662 -1883
rect 666 -1889 669 -1883
rect 673 -1889 676 -1883
rect 680 -1889 683 -1883
rect 687 -1889 690 -1883
rect 694 -1889 697 -1883
rect 701 -1889 704 -1883
rect 708 -1889 711 -1883
rect 715 -1889 718 -1883
rect 722 -1889 725 -1883
rect 729 -1889 732 -1883
rect 736 -1889 739 -1883
rect 743 -1889 749 -1883
rect 750 -1889 753 -1883
rect 1 -1972 4 -1966
rect 8 -1972 11 -1966
rect 15 -1972 21 -1966
rect 22 -1972 25 -1966
rect 29 -1972 35 -1966
rect 36 -1972 42 -1966
rect 43 -1972 46 -1966
rect 50 -1972 56 -1966
rect 57 -1972 63 -1966
rect 64 -1972 67 -1966
rect 71 -1972 77 -1966
rect 78 -1972 84 -1966
rect 85 -1972 88 -1966
rect 92 -1972 95 -1966
rect 99 -1972 105 -1966
rect 106 -1972 112 -1966
rect 113 -1972 119 -1966
rect 120 -1972 123 -1966
rect 127 -1972 130 -1966
rect 134 -1972 137 -1966
rect 141 -1972 144 -1966
rect 148 -1972 151 -1966
rect 155 -1972 161 -1966
rect 162 -1972 165 -1966
rect 169 -1972 175 -1966
rect 176 -1972 182 -1966
rect 183 -1972 186 -1966
rect 190 -1972 193 -1966
rect 197 -1972 203 -1966
rect 204 -1972 210 -1966
rect 211 -1972 217 -1966
rect 218 -1972 224 -1966
rect 225 -1972 228 -1966
rect 232 -1972 235 -1966
rect 239 -1972 242 -1966
rect 246 -1972 249 -1966
rect 253 -1972 256 -1966
rect 260 -1972 263 -1966
rect 267 -1972 273 -1966
rect 274 -1972 277 -1966
rect 281 -1972 284 -1966
rect 288 -1972 291 -1966
rect 295 -1972 298 -1966
rect 302 -1972 305 -1966
rect 309 -1972 315 -1966
rect 316 -1972 319 -1966
rect 323 -1972 326 -1966
rect 330 -1972 333 -1966
rect 337 -1972 340 -1966
rect 344 -1972 350 -1966
rect 351 -1972 357 -1966
rect 358 -1972 361 -1966
rect 365 -1972 371 -1966
rect 372 -1972 375 -1966
rect 379 -1972 382 -1966
rect 386 -1972 392 -1966
rect 393 -1972 399 -1966
rect 400 -1972 403 -1966
rect 407 -1972 410 -1966
rect 414 -1972 420 -1966
rect 421 -1972 427 -1966
rect 428 -1972 434 -1966
rect 435 -1972 438 -1966
rect 442 -1972 445 -1966
rect 449 -1972 452 -1966
rect 456 -1972 462 -1966
rect 463 -1972 469 -1966
rect 470 -1972 473 -1966
rect 477 -1972 483 -1966
rect 484 -1972 487 -1966
rect 491 -1972 494 -1966
rect 498 -1972 501 -1966
rect 505 -1972 508 -1966
rect 512 -1972 515 -1966
rect 519 -1972 522 -1966
rect 526 -1972 529 -1966
rect 533 -1972 536 -1966
rect 540 -1972 543 -1966
rect 547 -1972 553 -1966
rect 554 -1972 557 -1966
rect 561 -1972 564 -1966
rect 568 -1972 571 -1966
rect 575 -1972 578 -1966
rect 582 -1972 585 -1966
rect 589 -1972 592 -1966
rect 596 -1972 599 -1966
rect 603 -1972 606 -1966
rect 610 -1972 613 -1966
rect 617 -1972 620 -1966
rect 624 -1972 627 -1966
rect 631 -1972 634 -1966
rect 638 -1972 644 -1966
rect 645 -1972 648 -1966
rect 652 -1972 655 -1966
rect 659 -1972 662 -1966
rect 666 -1972 669 -1966
rect 673 -1972 676 -1966
rect 680 -1972 683 -1966
rect 687 -1972 690 -1966
rect 694 -1972 697 -1966
rect 701 -1972 704 -1966
rect 708 -1972 711 -1966
rect 715 -1972 718 -1966
rect 722 -1972 725 -1966
rect 729 -1972 732 -1966
rect 8 -2033 11 -2027
rect 15 -2033 18 -2027
rect 22 -2033 28 -2027
rect 29 -2033 32 -2027
rect 36 -2033 39 -2027
rect 43 -2033 46 -2027
rect 50 -2033 56 -2027
rect 57 -2033 60 -2027
rect 64 -2033 70 -2027
rect 71 -2033 74 -2027
rect 78 -2033 81 -2027
rect 85 -2033 91 -2027
rect 92 -2033 98 -2027
rect 99 -2033 105 -2027
rect 106 -2033 112 -2027
rect 113 -2033 119 -2027
rect 120 -2033 123 -2027
rect 127 -2033 133 -2027
rect 134 -2033 137 -2027
rect 141 -2033 144 -2027
rect 148 -2033 151 -2027
rect 155 -2033 158 -2027
rect 162 -2033 165 -2027
rect 169 -2033 172 -2027
rect 176 -2033 179 -2027
rect 183 -2033 189 -2027
rect 190 -2033 196 -2027
rect 197 -2033 203 -2027
rect 204 -2033 207 -2027
rect 211 -2033 217 -2027
rect 218 -2033 224 -2027
rect 225 -2033 228 -2027
rect 232 -2033 235 -2027
rect 239 -2033 242 -2027
rect 246 -2033 252 -2027
rect 253 -2033 259 -2027
rect 260 -2033 263 -2027
rect 267 -2033 270 -2027
rect 274 -2033 277 -2027
rect 281 -2033 287 -2027
rect 288 -2033 291 -2027
rect 295 -2033 298 -2027
rect 302 -2033 308 -2027
rect 309 -2033 312 -2027
rect 316 -2033 319 -2027
rect 323 -2033 326 -2027
rect 330 -2033 333 -2027
rect 337 -2033 340 -2027
rect 344 -2033 347 -2027
rect 351 -2033 354 -2027
rect 358 -2033 361 -2027
rect 365 -2033 368 -2027
rect 372 -2033 375 -2027
rect 379 -2033 385 -2027
rect 386 -2033 389 -2027
rect 393 -2033 396 -2027
rect 400 -2033 406 -2027
rect 407 -2033 410 -2027
rect 414 -2033 420 -2027
rect 421 -2033 424 -2027
rect 428 -2033 431 -2027
rect 435 -2033 441 -2027
rect 442 -2033 445 -2027
rect 449 -2033 452 -2027
rect 456 -2033 459 -2027
rect 463 -2033 466 -2027
rect 470 -2033 476 -2027
rect 477 -2033 480 -2027
rect 484 -2033 490 -2027
rect 491 -2033 494 -2027
rect 498 -2033 501 -2027
rect 505 -2033 508 -2027
rect 512 -2033 515 -2027
rect 519 -2033 525 -2027
rect 526 -2033 529 -2027
rect 533 -2033 536 -2027
rect 540 -2033 543 -2027
rect 547 -2033 553 -2027
rect 554 -2033 557 -2027
rect 561 -2033 564 -2027
rect 568 -2033 571 -2027
rect 575 -2033 578 -2027
rect 582 -2033 585 -2027
rect 589 -2033 592 -2027
rect 596 -2033 599 -2027
rect 603 -2033 606 -2027
rect 610 -2033 613 -2027
rect 617 -2033 620 -2027
rect 624 -2033 627 -2027
rect 631 -2033 637 -2027
rect 638 -2033 644 -2027
rect 645 -2033 651 -2027
rect 652 -2033 658 -2027
rect 659 -2033 662 -2027
rect 666 -2033 672 -2027
rect 694 -2033 697 -2027
rect 15 -2098 18 -2092
rect 22 -2098 28 -2092
rect 29 -2098 35 -2092
rect 36 -2098 39 -2092
rect 43 -2098 46 -2092
rect 50 -2098 53 -2092
rect 57 -2098 63 -2092
rect 64 -2098 67 -2092
rect 71 -2098 77 -2092
rect 78 -2098 81 -2092
rect 85 -2098 88 -2092
rect 92 -2098 98 -2092
rect 99 -2098 102 -2092
rect 106 -2098 109 -2092
rect 113 -2098 119 -2092
rect 120 -2098 123 -2092
rect 127 -2098 130 -2092
rect 134 -2098 137 -2092
rect 141 -2098 144 -2092
rect 148 -2098 151 -2092
rect 155 -2098 161 -2092
rect 162 -2098 165 -2092
rect 169 -2098 172 -2092
rect 176 -2098 179 -2092
rect 183 -2098 189 -2092
rect 190 -2098 196 -2092
rect 197 -2098 200 -2092
rect 204 -2098 210 -2092
rect 211 -2098 214 -2092
rect 218 -2098 224 -2092
rect 225 -2098 228 -2092
rect 232 -2098 238 -2092
rect 239 -2098 242 -2092
rect 246 -2098 249 -2092
rect 253 -2098 256 -2092
rect 260 -2098 263 -2092
rect 267 -2098 270 -2092
rect 274 -2098 277 -2092
rect 281 -2098 284 -2092
rect 288 -2098 291 -2092
rect 295 -2098 298 -2092
rect 302 -2098 308 -2092
rect 309 -2098 315 -2092
rect 316 -2098 322 -2092
rect 323 -2098 329 -2092
rect 330 -2098 333 -2092
rect 337 -2098 340 -2092
rect 344 -2098 347 -2092
rect 351 -2098 357 -2092
rect 358 -2098 361 -2092
rect 365 -2098 371 -2092
rect 372 -2098 375 -2092
rect 379 -2098 385 -2092
rect 386 -2098 389 -2092
rect 393 -2098 396 -2092
rect 400 -2098 406 -2092
rect 407 -2098 413 -2092
rect 414 -2098 420 -2092
rect 421 -2098 427 -2092
rect 428 -2098 431 -2092
rect 435 -2098 438 -2092
rect 442 -2098 445 -2092
rect 449 -2098 452 -2092
rect 456 -2098 459 -2092
rect 463 -2098 466 -2092
rect 470 -2098 473 -2092
rect 477 -2098 483 -2092
rect 484 -2098 487 -2092
rect 491 -2098 494 -2092
rect 498 -2098 504 -2092
rect 505 -2098 508 -2092
rect 512 -2098 515 -2092
rect 519 -2098 522 -2092
rect 526 -2098 529 -2092
rect 533 -2098 536 -2092
rect 540 -2098 543 -2092
rect 547 -2098 550 -2092
rect 554 -2098 560 -2092
rect 561 -2098 564 -2092
rect 568 -2098 571 -2092
rect 575 -2098 578 -2092
rect 582 -2098 585 -2092
rect 589 -2098 595 -2092
rect 603 -2098 606 -2092
rect 610 -2098 613 -2092
rect 617 -2098 623 -2092
rect 638 -2098 644 -2092
rect 645 -2098 648 -2092
rect 673 -2098 679 -2092
rect 687 -2098 690 -2092
rect 22 -2155 28 -2149
rect 29 -2155 35 -2149
rect 36 -2155 39 -2149
rect 43 -2155 46 -2149
rect 50 -2155 53 -2149
rect 57 -2155 60 -2149
rect 64 -2155 67 -2149
rect 71 -2155 77 -2149
rect 78 -2155 84 -2149
rect 85 -2155 88 -2149
rect 92 -2155 98 -2149
rect 99 -2155 102 -2149
rect 106 -2155 109 -2149
rect 113 -2155 119 -2149
rect 120 -2155 126 -2149
rect 127 -2155 133 -2149
rect 134 -2155 137 -2149
rect 141 -2155 144 -2149
rect 148 -2155 154 -2149
rect 155 -2155 158 -2149
rect 162 -2155 165 -2149
rect 169 -2155 172 -2149
rect 176 -2155 182 -2149
rect 183 -2155 189 -2149
rect 190 -2155 193 -2149
rect 197 -2155 200 -2149
rect 204 -2155 207 -2149
rect 211 -2155 217 -2149
rect 218 -2155 224 -2149
rect 225 -2155 228 -2149
rect 232 -2155 235 -2149
rect 239 -2155 242 -2149
rect 246 -2155 249 -2149
rect 253 -2155 259 -2149
rect 260 -2155 266 -2149
rect 267 -2155 270 -2149
rect 274 -2155 277 -2149
rect 281 -2155 287 -2149
rect 288 -2155 294 -2149
rect 295 -2155 298 -2149
rect 302 -2155 308 -2149
rect 309 -2155 312 -2149
rect 316 -2155 322 -2149
rect 323 -2155 326 -2149
rect 330 -2155 336 -2149
rect 337 -2155 343 -2149
rect 344 -2155 347 -2149
rect 351 -2155 354 -2149
rect 358 -2155 364 -2149
rect 365 -2155 371 -2149
rect 372 -2155 378 -2149
rect 379 -2155 382 -2149
rect 386 -2155 389 -2149
rect 393 -2155 396 -2149
rect 400 -2155 403 -2149
rect 407 -2155 410 -2149
rect 414 -2155 420 -2149
rect 421 -2155 424 -2149
rect 428 -2155 431 -2149
rect 435 -2155 438 -2149
rect 442 -2155 445 -2149
rect 449 -2155 452 -2149
rect 456 -2155 459 -2149
rect 463 -2155 469 -2149
rect 470 -2155 473 -2149
rect 477 -2155 480 -2149
rect 484 -2155 487 -2149
rect 491 -2155 494 -2149
rect 498 -2155 504 -2149
rect 505 -2155 511 -2149
rect 512 -2155 515 -2149
rect 519 -2155 525 -2149
rect 526 -2155 532 -2149
rect 533 -2155 536 -2149
rect 540 -2155 543 -2149
rect 547 -2155 550 -2149
rect 554 -2155 557 -2149
rect 561 -2155 564 -2149
rect 568 -2155 571 -2149
rect 589 -2155 592 -2149
rect 596 -2155 599 -2149
rect 610 -2155 613 -2149
rect 8 -2202 11 -2196
rect 15 -2202 21 -2196
rect 22 -2202 28 -2196
rect 36 -2202 42 -2196
rect 43 -2202 49 -2196
rect 50 -2202 53 -2196
rect 57 -2202 60 -2196
rect 64 -2202 67 -2196
rect 71 -2202 74 -2196
rect 78 -2202 81 -2196
rect 85 -2202 88 -2196
rect 92 -2202 95 -2196
rect 99 -2202 102 -2196
rect 106 -2202 109 -2196
rect 113 -2202 119 -2196
rect 120 -2202 123 -2196
rect 127 -2202 133 -2196
rect 134 -2202 140 -2196
rect 141 -2202 147 -2196
rect 148 -2202 154 -2196
rect 155 -2202 158 -2196
rect 162 -2202 165 -2196
rect 169 -2202 172 -2196
rect 176 -2202 179 -2196
rect 183 -2202 189 -2196
rect 190 -2202 193 -2196
rect 197 -2202 203 -2196
rect 204 -2202 210 -2196
rect 211 -2202 217 -2196
rect 218 -2202 221 -2196
rect 225 -2202 228 -2196
rect 232 -2202 238 -2196
rect 246 -2202 249 -2196
rect 253 -2202 259 -2196
rect 260 -2202 263 -2196
rect 267 -2202 270 -2196
rect 274 -2202 280 -2196
rect 281 -2202 287 -2196
rect 288 -2202 291 -2196
rect 295 -2202 301 -2196
rect 302 -2202 305 -2196
rect 316 -2202 319 -2196
rect 323 -2202 329 -2196
rect 330 -2202 333 -2196
rect 344 -2202 350 -2196
rect 351 -2202 354 -2196
rect 358 -2202 364 -2196
rect 365 -2202 371 -2196
rect 372 -2202 378 -2196
rect 379 -2202 382 -2196
rect 386 -2202 389 -2196
rect 393 -2202 396 -2196
rect 400 -2202 403 -2196
rect 407 -2202 410 -2196
rect 414 -2202 420 -2196
rect 421 -2202 427 -2196
rect 428 -2202 431 -2196
rect 435 -2202 438 -2196
rect 442 -2202 445 -2196
rect 449 -2202 455 -2196
rect 456 -2202 459 -2196
rect 463 -2202 466 -2196
rect 477 -2202 483 -2196
rect 491 -2202 497 -2196
rect 498 -2202 504 -2196
rect 519 -2202 522 -2196
rect 533 -2202 536 -2196
rect 547 -2202 553 -2196
rect 554 -2202 557 -2196
rect 596 -2202 602 -2196
rect 603 -2202 606 -2196
rect 610 -2202 613 -2196
rect 15 -2231 21 -2225
rect 22 -2231 28 -2225
rect 43 -2231 49 -2225
rect 50 -2231 56 -2225
rect 57 -2231 60 -2225
rect 71 -2231 77 -2225
rect 78 -2231 84 -2225
rect 92 -2231 98 -2225
rect 99 -2231 105 -2225
rect 106 -2231 109 -2225
rect 113 -2231 116 -2225
rect 127 -2231 133 -2225
rect 148 -2231 151 -2225
rect 162 -2231 168 -2225
rect 169 -2231 175 -2225
rect 176 -2231 182 -2225
rect 183 -2231 189 -2225
rect 190 -2231 196 -2225
rect 197 -2231 203 -2225
rect 204 -2231 210 -2225
rect 211 -2231 217 -2225
rect 218 -2231 224 -2225
rect 225 -2231 228 -2225
rect 239 -2231 242 -2225
rect 246 -2231 249 -2225
rect 253 -2231 256 -2225
rect 267 -2231 270 -2225
rect 274 -2231 277 -2225
rect 281 -2231 284 -2225
rect 288 -2231 291 -2225
rect 302 -2231 308 -2225
rect 309 -2231 315 -2225
rect 323 -2231 329 -2225
rect 330 -2231 333 -2225
rect 337 -2231 343 -2225
rect 344 -2231 350 -2225
rect 351 -2231 357 -2225
rect 372 -2231 375 -2225
rect 379 -2231 385 -2225
rect 386 -2231 392 -2225
rect 407 -2231 410 -2225
rect 428 -2231 434 -2225
rect 449 -2231 452 -2225
rect 470 -2231 476 -2225
rect 484 -2231 490 -2225
rect 505 -2231 508 -2225
rect 533 -2231 539 -2225
rect 610 -2231 616 -2225
<< polysilicon >>
rect 26 -13 27 -11
rect 107 -13 108 -11
rect 110 -13 111 -11
rect 117 -13 118 -11
rect 131 -7 132 -5
rect 138 -13 139 -11
rect 142 -13 143 -11
rect 156 -7 157 -5
rect 156 -13 157 -11
rect 163 -7 164 -5
rect 163 -13 164 -11
rect 170 -13 171 -11
rect 177 -7 178 -5
rect 177 -13 178 -11
rect 187 -7 188 -5
rect 191 -7 192 -5
rect 191 -13 192 -11
rect 198 -13 199 -11
rect 205 -13 206 -11
rect 212 -7 213 -5
rect 215 -7 216 -5
rect 222 -13 223 -11
rect 226 -7 227 -5
rect 226 -13 227 -11
rect 233 -7 234 -5
rect 243 -13 244 -11
rect 247 -7 248 -5
rect 247 -13 248 -11
rect 257 -7 258 -5
rect 257 -13 258 -11
rect 261 -7 262 -5
rect 261 -13 262 -11
rect 268 -7 269 -5
rect 268 -13 269 -11
rect 278 -7 279 -5
rect 282 -7 283 -5
rect 282 -13 283 -11
rect 327 -13 328 -11
rect 26 -34 27 -32
rect 72 -40 73 -38
rect 86 -34 87 -32
rect 86 -40 87 -38
rect 93 -34 94 -32
rect 93 -40 94 -38
rect 100 -34 101 -32
rect 110 -34 111 -32
rect 114 -40 115 -38
rect 121 -40 122 -38
rect 128 -34 129 -32
rect 135 -40 136 -38
rect 142 -34 143 -32
rect 142 -40 143 -38
rect 149 -34 150 -32
rect 149 -40 150 -38
rect 156 -34 157 -32
rect 156 -40 157 -38
rect 166 -34 167 -32
rect 170 -34 171 -32
rect 170 -40 171 -38
rect 177 -34 178 -32
rect 180 -34 181 -32
rect 177 -40 178 -38
rect 180 -40 181 -38
rect 184 -34 185 -32
rect 184 -40 185 -38
rect 191 -34 192 -32
rect 191 -40 192 -38
rect 198 -34 199 -32
rect 198 -40 199 -38
rect 208 -34 209 -32
rect 212 -34 213 -32
rect 215 -34 216 -32
rect 212 -40 213 -38
rect 219 -34 220 -32
rect 219 -40 220 -38
rect 229 -40 230 -38
rect 233 -34 234 -32
rect 233 -40 234 -38
rect 240 -34 241 -32
rect 240 -40 241 -38
rect 247 -34 248 -32
rect 247 -40 248 -38
rect 254 -34 255 -32
rect 254 -40 255 -38
rect 261 -34 262 -32
rect 261 -40 262 -38
rect 268 -34 269 -32
rect 268 -40 269 -38
rect 275 -34 276 -32
rect 275 -40 276 -38
rect 282 -34 283 -32
rect 282 -40 283 -38
rect 285 -40 286 -38
rect 289 -34 290 -32
rect 289 -40 290 -38
rect 296 -34 297 -32
rect 296 -40 297 -38
rect 303 -34 304 -32
rect 303 -40 304 -38
rect 313 -40 314 -38
rect 317 -34 318 -32
rect 317 -40 318 -38
rect 324 -40 325 -38
rect 331 -34 332 -32
rect 331 -40 332 -38
rect 338 -40 339 -38
rect 345 -34 346 -32
rect 345 -40 346 -38
rect 352 -34 353 -32
rect 352 -40 353 -38
rect 359 -34 360 -32
rect 359 -40 360 -38
rect 369 -34 370 -32
rect 376 -34 377 -32
rect 380 -34 381 -32
rect 380 -40 381 -38
rect 387 -34 388 -32
rect 387 -40 388 -38
rect 394 -40 395 -38
rect 401 -34 402 -32
rect 401 -40 402 -38
rect 418 -34 419 -32
rect 44 -77 45 -75
rect 44 -83 45 -81
rect 51 -77 52 -75
rect 51 -83 52 -81
rect 65 -77 66 -75
rect 65 -83 66 -81
rect 75 -77 76 -75
rect 79 -77 80 -75
rect 79 -83 80 -81
rect 86 -77 87 -75
rect 96 -83 97 -81
rect 100 -77 101 -75
rect 107 -77 108 -75
rect 107 -83 108 -81
rect 114 -77 115 -75
rect 117 -77 118 -75
rect 114 -83 115 -81
rect 121 -77 122 -75
rect 124 -83 125 -81
rect 128 -77 129 -75
rect 131 -77 132 -75
rect 135 -77 136 -75
rect 135 -83 136 -81
rect 142 -83 143 -81
rect 145 -83 146 -81
rect 149 -77 150 -75
rect 149 -83 150 -81
rect 156 -77 157 -75
rect 159 -83 160 -81
rect 163 -77 164 -75
rect 163 -83 164 -81
rect 170 -77 171 -75
rect 173 -77 174 -75
rect 184 -77 185 -75
rect 184 -83 185 -81
rect 191 -83 192 -81
rect 194 -83 195 -81
rect 198 -77 199 -75
rect 198 -83 199 -81
rect 205 -77 206 -75
rect 212 -77 213 -75
rect 215 -77 216 -75
rect 212 -83 213 -81
rect 215 -83 216 -81
rect 219 -77 220 -75
rect 222 -77 223 -75
rect 219 -83 220 -81
rect 222 -83 223 -81
rect 226 -77 227 -75
rect 233 -77 234 -75
rect 233 -83 234 -81
rect 240 -77 241 -75
rect 240 -83 241 -81
rect 247 -77 248 -75
rect 247 -83 248 -81
rect 254 -77 255 -75
rect 257 -77 258 -75
rect 254 -83 255 -81
rect 257 -83 258 -81
rect 261 -77 262 -75
rect 261 -83 262 -81
rect 271 -83 272 -81
rect 275 -77 276 -75
rect 278 -83 279 -81
rect 282 -77 283 -75
rect 289 -77 290 -75
rect 289 -83 290 -81
rect 296 -77 297 -75
rect 296 -83 297 -81
rect 303 -77 304 -75
rect 303 -83 304 -81
rect 310 -77 311 -75
rect 310 -83 311 -81
rect 317 -77 318 -75
rect 317 -83 318 -81
rect 324 -77 325 -75
rect 324 -83 325 -81
rect 331 -77 332 -75
rect 331 -83 332 -81
rect 338 -77 339 -75
rect 338 -83 339 -81
rect 345 -77 346 -75
rect 345 -83 346 -81
rect 352 -83 353 -81
rect 359 -77 360 -75
rect 359 -83 360 -81
rect 366 -77 367 -75
rect 366 -83 367 -81
rect 373 -77 374 -75
rect 373 -83 374 -81
rect 380 -77 381 -75
rect 380 -83 381 -81
rect 387 -77 388 -75
rect 387 -83 388 -81
rect 394 -77 395 -75
rect 394 -83 395 -81
rect 401 -77 402 -75
rect 401 -83 402 -81
rect 408 -77 409 -75
rect 408 -83 409 -81
rect 432 -83 433 -81
rect 58 -122 59 -120
rect 58 -128 59 -126
rect 65 -122 66 -120
rect 79 -122 80 -120
rect 79 -128 80 -126
rect 86 -122 87 -120
rect 86 -128 87 -126
rect 93 -122 94 -120
rect 93 -128 94 -126
rect 100 -122 101 -120
rect 100 -128 101 -126
rect 103 -128 104 -126
rect 107 -122 108 -120
rect 107 -128 108 -126
rect 117 -128 118 -126
rect 121 -122 122 -120
rect 121 -128 122 -126
rect 128 -122 129 -120
rect 131 -122 132 -120
rect 131 -128 132 -126
rect 138 -128 139 -126
rect 142 -128 143 -126
rect 145 -128 146 -126
rect 149 -122 150 -120
rect 149 -128 150 -126
rect 156 -122 157 -120
rect 163 -122 164 -120
rect 166 -128 167 -126
rect 170 -122 171 -120
rect 170 -128 171 -126
rect 177 -122 178 -120
rect 177 -128 178 -126
rect 184 -122 185 -120
rect 184 -128 185 -126
rect 191 -122 192 -120
rect 191 -128 192 -126
rect 201 -122 202 -120
rect 198 -128 199 -126
rect 205 -122 206 -120
rect 205 -128 206 -126
rect 212 -122 213 -120
rect 215 -122 216 -120
rect 215 -128 216 -126
rect 222 -128 223 -126
rect 226 -122 227 -120
rect 226 -128 227 -126
rect 236 -128 237 -126
rect 240 -122 241 -120
rect 247 -122 248 -120
rect 250 -122 251 -120
rect 247 -128 248 -126
rect 250 -128 251 -126
rect 254 -122 255 -120
rect 254 -128 255 -126
rect 261 -122 262 -120
rect 271 -122 272 -120
rect 275 -122 276 -120
rect 278 -122 279 -120
rect 282 -122 283 -120
rect 282 -128 283 -126
rect 289 -122 290 -120
rect 289 -128 290 -126
rect 296 -122 297 -120
rect 296 -128 297 -126
rect 303 -122 304 -120
rect 303 -128 304 -126
rect 310 -128 311 -126
rect 317 -122 318 -120
rect 317 -128 318 -126
rect 324 -122 325 -120
rect 324 -128 325 -126
rect 331 -122 332 -120
rect 331 -128 332 -126
rect 338 -122 339 -120
rect 338 -128 339 -126
rect 345 -122 346 -120
rect 345 -128 346 -126
rect 352 -122 353 -120
rect 352 -128 353 -126
rect 359 -122 360 -120
rect 359 -128 360 -126
rect 366 -122 367 -120
rect 373 -122 374 -120
rect 373 -128 374 -126
rect 383 -122 384 -120
rect 380 -128 381 -126
rect 387 -122 388 -120
rect 387 -128 388 -126
rect 394 -122 395 -120
rect 394 -128 395 -126
rect 401 -122 402 -120
rect 401 -128 402 -126
rect 408 -122 409 -120
rect 408 -128 409 -126
rect 415 -122 416 -120
rect 415 -128 416 -126
rect 422 -122 423 -120
rect 422 -128 423 -126
rect 429 -122 430 -120
rect 429 -128 430 -126
rect 439 -128 440 -126
rect 443 -122 444 -120
rect 443 -128 444 -126
rect 453 -122 454 -120
rect 37 -175 38 -173
rect 37 -181 38 -179
rect 44 -175 45 -173
rect 44 -181 45 -179
rect 51 -175 52 -173
rect 51 -181 52 -179
rect 58 -175 59 -173
rect 58 -181 59 -179
rect 68 -181 69 -179
rect 72 -175 73 -173
rect 72 -181 73 -179
rect 79 -175 80 -173
rect 79 -181 80 -179
rect 89 -175 90 -173
rect 89 -181 90 -179
rect 93 -175 94 -173
rect 96 -181 97 -179
rect 100 -175 101 -173
rect 100 -181 101 -179
rect 110 -175 111 -173
rect 114 -175 115 -173
rect 114 -181 115 -179
rect 121 -175 122 -173
rect 121 -181 122 -179
rect 128 -175 129 -173
rect 128 -181 129 -179
rect 138 -175 139 -173
rect 135 -181 136 -179
rect 142 -181 143 -179
rect 145 -181 146 -179
rect 149 -181 150 -179
rect 152 -181 153 -179
rect 156 -175 157 -173
rect 156 -181 157 -179
rect 166 -175 167 -173
rect 170 -175 171 -173
rect 170 -181 171 -179
rect 177 -175 178 -173
rect 177 -181 178 -179
rect 184 -175 185 -173
rect 187 -181 188 -179
rect 191 -175 192 -173
rect 191 -181 192 -179
rect 198 -175 199 -173
rect 198 -181 199 -179
rect 208 -175 209 -173
rect 208 -181 209 -179
rect 212 -181 213 -179
rect 215 -181 216 -179
rect 219 -175 220 -173
rect 219 -181 220 -179
rect 226 -175 227 -173
rect 226 -181 227 -179
rect 233 -175 234 -173
rect 236 -175 237 -173
rect 233 -181 234 -179
rect 243 -181 244 -179
rect 247 -175 248 -173
rect 247 -181 248 -179
rect 254 -175 255 -173
rect 257 -181 258 -179
rect 261 -175 262 -173
rect 261 -181 262 -179
rect 268 -175 269 -173
rect 268 -181 269 -179
rect 275 -175 276 -173
rect 278 -181 279 -179
rect 285 -175 286 -173
rect 289 -181 290 -179
rect 292 -181 293 -179
rect 296 -175 297 -173
rect 296 -181 297 -179
rect 306 -175 307 -173
rect 306 -181 307 -179
rect 313 -175 314 -173
rect 317 -175 318 -173
rect 320 -175 321 -173
rect 324 -175 325 -173
rect 324 -181 325 -179
rect 331 -175 332 -173
rect 331 -181 332 -179
rect 334 -181 335 -179
rect 338 -175 339 -173
rect 338 -181 339 -179
rect 345 -175 346 -173
rect 345 -181 346 -179
rect 352 -175 353 -173
rect 352 -181 353 -179
rect 359 -175 360 -173
rect 359 -181 360 -179
rect 366 -175 367 -173
rect 366 -181 367 -179
rect 373 -175 374 -173
rect 373 -181 374 -179
rect 380 -175 381 -173
rect 380 -181 381 -179
rect 387 -175 388 -173
rect 387 -181 388 -179
rect 394 -175 395 -173
rect 394 -181 395 -179
rect 401 -175 402 -173
rect 401 -181 402 -179
rect 408 -175 409 -173
rect 408 -181 409 -179
rect 415 -175 416 -173
rect 415 -181 416 -179
rect 429 -175 430 -173
rect 429 -181 430 -179
rect 436 -175 437 -173
rect 436 -181 437 -179
rect 443 -175 444 -173
rect 443 -181 444 -179
rect 450 -175 451 -173
rect 450 -181 451 -179
rect 457 -175 458 -173
rect 457 -181 458 -179
rect 464 -175 465 -173
rect 464 -181 465 -179
rect 471 -175 472 -173
rect 471 -181 472 -179
rect 481 -175 482 -173
rect 485 -175 486 -173
rect 485 -181 486 -179
rect 492 -175 493 -173
rect 492 -181 493 -179
rect 548 -181 549 -179
rect 16 -232 17 -230
rect 16 -238 17 -236
rect 30 -232 31 -230
rect 30 -238 31 -236
rect 37 -232 38 -230
rect 58 -232 59 -230
rect 65 -232 66 -230
rect 79 -232 80 -230
rect 82 -232 83 -230
rect 82 -238 83 -236
rect 86 -232 87 -230
rect 89 -232 90 -230
rect 93 -232 94 -230
rect 93 -238 94 -236
rect 100 -232 101 -230
rect 103 -232 104 -230
rect 100 -238 101 -236
rect 103 -238 104 -236
rect 107 -232 108 -230
rect 107 -238 108 -236
rect 114 -232 115 -230
rect 114 -238 115 -236
rect 121 -232 122 -230
rect 124 -232 125 -230
rect 128 -232 129 -230
rect 128 -238 129 -236
rect 135 -232 136 -230
rect 135 -238 136 -236
rect 142 -232 143 -230
rect 152 -232 153 -230
rect 149 -238 150 -236
rect 152 -238 153 -236
rect 156 -232 157 -230
rect 156 -238 157 -236
rect 163 -232 164 -230
rect 163 -238 164 -236
rect 166 -238 167 -236
rect 170 -232 171 -230
rect 170 -238 171 -236
rect 177 -232 178 -230
rect 177 -238 178 -236
rect 184 -232 185 -230
rect 184 -238 185 -236
rect 191 -232 192 -230
rect 191 -238 192 -236
rect 198 -232 199 -230
rect 198 -238 199 -236
rect 205 -232 206 -230
rect 205 -238 206 -236
rect 212 -232 213 -230
rect 215 -238 216 -236
rect 219 -232 220 -230
rect 222 -232 223 -230
rect 222 -238 223 -236
rect 226 -232 227 -230
rect 226 -238 227 -236
rect 233 -232 234 -230
rect 233 -238 234 -236
rect 240 -232 241 -230
rect 243 -232 244 -230
rect 240 -238 241 -236
rect 243 -238 244 -236
rect 247 -232 248 -230
rect 247 -238 248 -236
rect 254 -232 255 -230
rect 257 -238 258 -236
rect 261 -232 262 -230
rect 261 -238 262 -236
rect 268 -232 269 -230
rect 268 -238 269 -236
rect 275 -232 276 -230
rect 275 -238 276 -236
rect 282 -232 283 -230
rect 285 -232 286 -230
rect 282 -238 283 -236
rect 285 -238 286 -236
rect 289 -232 290 -230
rect 289 -238 290 -236
rect 303 -232 304 -230
rect 303 -238 304 -236
rect 310 -232 311 -230
rect 317 -232 318 -230
rect 317 -238 318 -236
rect 324 -232 325 -230
rect 324 -238 325 -236
rect 331 -232 332 -230
rect 331 -238 332 -236
rect 341 -232 342 -230
rect 345 -232 346 -230
rect 345 -238 346 -236
rect 352 -238 353 -236
rect 359 -232 360 -230
rect 362 -238 363 -236
rect 366 -232 367 -230
rect 366 -238 367 -236
rect 373 -232 374 -230
rect 373 -238 374 -236
rect 380 -232 381 -230
rect 380 -238 381 -236
rect 387 -232 388 -230
rect 387 -238 388 -236
rect 394 -232 395 -230
rect 394 -238 395 -236
rect 401 -232 402 -230
rect 401 -238 402 -236
rect 408 -232 409 -230
rect 408 -238 409 -236
rect 415 -232 416 -230
rect 415 -238 416 -236
rect 422 -232 423 -230
rect 422 -238 423 -236
rect 429 -232 430 -230
rect 429 -238 430 -236
rect 436 -232 437 -230
rect 436 -238 437 -236
rect 443 -232 444 -230
rect 443 -238 444 -236
rect 450 -232 451 -230
rect 450 -238 451 -236
rect 457 -232 458 -230
rect 457 -238 458 -236
rect 464 -232 465 -230
rect 464 -238 465 -236
rect 471 -232 472 -230
rect 471 -238 472 -236
rect 478 -232 479 -230
rect 478 -238 479 -236
rect 485 -232 486 -230
rect 485 -238 486 -236
rect 492 -232 493 -230
rect 492 -238 493 -236
rect 499 -232 500 -230
rect 499 -238 500 -236
rect 506 -232 507 -230
rect 506 -238 507 -236
rect 513 -232 514 -230
rect 513 -238 514 -236
rect 520 -232 521 -230
rect 527 -232 528 -230
rect 527 -238 528 -236
rect 534 -232 535 -230
rect 534 -238 535 -236
rect 541 -238 542 -236
rect 548 -232 549 -230
rect 555 -232 556 -230
rect 555 -238 556 -236
rect 558 -238 559 -236
rect 565 -232 566 -230
rect 565 -238 566 -236
rect 583 -232 584 -230
rect 586 -238 587 -236
rect 639 -232 640 -230
rect 639 -238 640 -236
rect 653 -238 654 -236
rect 26 -295 27 -293
rect 30 -289 31 -287
rect 30 -295 31 -293
rect 40 -289 41 -287
rect 44 -289 45 -287
rect 44 -295 45 -293
rect 51 -289 52 -287
rect 51 -295 52 -293
rect 58 -289 59 -287
rect 58 -295 59 -293
rect 65 -295 66 -293
rect 72 -289 73 -287
rect 72 -295 73 -293
rect 79 -289 80 -287
rect 79 -295 80 -293
rect 86 -289 87 -287
rect 86 -295 87 -293
rect 93 -289 94 -287
rect 93 -295 94 -293
rect 100 -289 101 -287
rect 100 -295 101 -293
rect 107 -289 108 -287
rect 107 -295 108 -293
rect 114 -289 115 -287
rect 114 -295 115 -293
rect 124 -289 125 -287
rect 128 -289 129 -287
rect 128 -295 129 -293
rect 135 -289 136 -287
rect 135 -295 136 -293
rect 145 -289 146 -287
rect 142 -295 143 -293
rect 152 -289 153 -287
rect 149 -295 150 -293
rect 156 -289 157 -287
rect 156 -295 157 -293
rect 163 -289 164 -287
rect 163 -295 164 -293
rect 166 -295 167 -293
rect 170 -289 171 -287
rect 170 -295 171 -293
rect 180 -289 181 -287
rect 177 -295 178 -293
rect 184 -289 185 -287
rect 184 -295 185 -293
rect 194 -289 195 -287
rect 191 -295 192 -293
rect 198 -289 199 -287
rect 198 -295 199 -293
rect 205 -289 206 -287
rect 205 -295 206 -293
rect 212 -289 213 -287
rect 215 -289 216 -287
rect 215 -295 216 -293
rect 219 -289 220 -287
rect 219 -295 220 -293
rect 222 -295 223 -293
rect 226 -289 227 -287
rect 226 -295 227 -293
rect 233 -289 234 -287
rect 233 -295 234 -293
rect 240 -289 241 -287
rect 240 -295 241 -293
rect 247 -289 248 -287
rect 247 -295 248 -293
rect 250 -295 251 -293
rect 254 -289 255 -287
rect 254 -295 255 -293
rect 257 -295 258 -293
rect 261 -289 262 -287
rect 261 -295 262 -293
rect 268 -289 269 -287
rect 268 -295 269 -293
rect 275 -289 276 -287
rect 278 -289 279 -287
rect 278 -295 279 -293
rect 285 -289 286 -287
rect 282 -295 283 -293
rect 289 -289 290 -287
rect 289 -295 290 -293
rect 296 -289 297 -287
rect 299 -289 300 -287
rect 299 -295 300 -293
rect 303 -289 304 -287
rect 303 -295 304 -293
rect 310 -289 311 -287
rect 313 -289 314 -287
rect 310 -295 311 -293
rect 313 -295 314 -293
rect 317 -295 318 -293
rect 320 -295 321 -293
rect 324 -289 325 -287
rect 324 -295 325 -293
rect 331 -289 332 -287
rect 331 -295 332 -293
rect 338 -289 339 -287
rect 338 -295 339 -293
rect 341 -295 342 -293
rect 345 -289 346 -287
rect 345 -295 346 -293
rect 352 -289 353 -287
rect 352 -295 353 -293
rect 359 -289 360 -287
rect 359 -295 360 -293
rect 362 -295 363 -293
rect 366 -289 367 -287
rect 366 -295 367 -293
rect 373 -289 374 -287
rect 373 -295 374 -293
rect 380 -289 381 -287
rect 380 -295 381 -293
rect 387 -289 388 -287
rect 387 -295 388 -293
rect 394 -289 395 -287
rect 394 -295 395 -293
rect 401 -289 402 -287
rect 401 -295 402 -293
rect 408 -289 409 -287
rect 408 -295 409 -293
rect 415 -289 416 -287
rect 415 -295 416 -293
rect 422 -289 423 -287
rect 422 -295 423 -293
rect 429 -289 430 -287
rect 429 -295 430 -293
rect 439 -289 440 -287
rect 436 -295 437 -293
rect 443 -289 444 -287
rect 443 -295 444 -293
rect 450 -289 451 -287
rect 450 -295 451 -293
rect 457 -289 458 -287
rect 457 -295 458 -293
rect 464 -289 465 -287
rect 464 -295 465 -293
rect 471 -289 472 -287
rect 471 -295 472 -293
rect 481 -289 482 -287
rect 485 -289 486 -287
rect 485 -295 486 -293
rect 492 -289 493 -287
rect 492 -295 493 -293
rect 499 -289 500 -287
rect 499 -295 500 -293
rect 506 -289 507 -287
rect 506 -295 507 -293
rect 513 -289 514 -287
rect 513 -295 514 -293
rect 520 -289 521 -287
rect 520 -295 521 -293
rect 527 -289 528 -287
rect 527 -295 528 -293
rect 534 -289 535 -287
rect 534 -295 535 -293
rect 541 -289 542 -287
rect 541 -295 542 -293
rect 548 -289 549 -287
rect 548 -295 549 -293
rect 555 -289 556 -287
rect 555 -295 556 -293
rect 562 -289 563 -287
rect 562 -295 563 -293
rect 569 -289 570 -287
rect 569 -295 570 -293
rect 576 -289 577 -287
rect 576 -295 577 -293
rect 583 -289 584 -287
rect 583 -295 584 -293
rect 590 -289 591 -287
rect 590 -295 591 -293
rect 597 -289 598 -287
rect 597 -295 598 -293
rect 604 -289 605 -287
rect 604 -295 605 -293
rect 611 -289 612 -287
rect 611 -295 612 -293
rect 618 -289 619 -287
rect 618 -295 619 -293
rect 625 -289 626 -287
rect 625 -295 626 -293
rect 632 -289 633 -287
rect 632 -295 633 -293
rect 653 -289 654 -287
rect 653 -295 654 -293
rect 660 -289 661 -287
rect 660 -295 661 -293
rect 9 -358 10 -356
rect 9 -364 10 -362
rect 23 -358 24 -356
rect 23 -364 24 -362
rect 30 -358 31 -356
rect 30 -364 31 -362
rect 58 -358 59 -356
rect 58 -364 59 -362
rect 72 -358 73 -356
rect 72 -364 73 -362
rect 79 -358 80 -356
rect 79 -364 80 -362
rect 86 -358 87 -356
rect 86 -364 87 -362
rect 93 -358 94 -356
rect 93 -364 94 -362
rect 100 -358 101 -356
rect 107 -358 108 -356
rect 110 -358 111 -356
rect 107 -364 108 -362
rect 114 -358 115 -356
rect 117 -364 118 -362
rect 121 -358 122 -356
rect 121 -364 122 -362
rect 128 -358 129 -356
rect 128 -364 129 -362
rect 135 -358 136 -356
rect 135 -364 136 -362
rect 142 -358 143 -356
rect 142 -364 143 -362
rect 152 -358 153 -356
rect 149 -364 150 -362
rect 152 -364 153 -362
rect 159 -364 160 -362
rect 163 -358 164 -356
rect 163 -364 164 -362
rect 170 -358 171 -356
rect 170 -364 171 -362
rect 177 -358 178 -356
rect 177 -364 178 -362
rect 180 -364 181 -362
rect 184 -358 185 -356
rect 187 -358 188 -356
rect 191 -358 192 -356
rect 191 -364 192 -362
rect 194 -364 195 -362
rect 198 -358 199 -356
rect 198 -364 199 -362
rect 208 -364 209 -362
rect 212 -358 213 -356
rect 212 -364 213 -362
rect 219 -358 220 -356
rect 222 -358 223 -356
rect 219 -364 220 -362
rect 222 -364 223 -362
rect 226 -358 227 -356
rect 226 -364 227 -362
rect 233 -358 234 -356
rect 233 -364 234 -362
rect 240 -358 241 -356
rect 240 -364 241 -362
rect 247 -358 248 -356
rect 247 -364 248 -362
rect 254 -358 255 -356
rect 254 -364 255 -362
rect 261 -358 262 -356
rect 261 -364 262 -362
rect 268 -358 269 -356
rect 268 -364 269 -362
rect 275 -358 276 -356
rect 278 -358 279 -356
rect 275 -364 276 -362
rect 282 -364 283 -362
rect 289 -358 290 -356
rect 289 -364 290 -362
rect 296 -358 297 -356
rect 299 -358 300 -356
rect 296 -364 297 -362
rect 303 -358 304 -356
rect 303 -364 304 -362
rect 310 -358 311 -356
rect 310 -364 311 -362
rect 317 -358 318 -356
rect 317 -364 318 -362
rect 324 -364 325 -362
rect 327 -364 328 -362
rect 331 -358 332 -356
rect 331 -364 332 -362
rect 338 -358 339 -356
rect 338 -364 339 -362
rect 345 -358 346 -356
rect 345 -364 346 -362
rect 352 -358 353 -356
rect 352 -364 353 -362
rect 355 -364 356 -362
rect 362 -358 363 -356
rect 362 -364 363 -362
rect 366 -364 367 -362
rect 373 -358 374 -356
rect 373 -364 374 -362
rect 383 -358 384 -356
rect 383 -364 384 -362
rect 390 -358 391 -356
rect 387 -364 388 -362
rect 390 -364 391 -362
rect 394 -358 395 -356
rect 394 -364 395 -362
rect 401 -358 402 -356
rect 401 -364 402 -362
rect 408 -358 409 -356
rect 408 -364 409 -362
rect 415 -358 416 -356
rect 415 -364 416 -362
rect 422 -358 423 -356
rect 422 -364 423 -362
rect 429 -358 430 -356
rect 432 -358 433 -356
rect 429 -364 430 -362
rect 436 -358 437 -356
rect 436 -364 437 -362
rect 443 -358 444 -356
rect 443 -364 444 -362
rect 453 -358 454 -356
rect 453 -364 454 -362
rect 457 -358 458 -356
rect 457 -364 458 -362
rect 464 -358 465 -356
rect 464 -364 465 -362
rect 471 -358 472 -356
rect 471 -364 472 -362
rect 478 -358 479 -356
rect 478 -364 479 -362
rect 485 -358 486 -356
rect 485 -364 486 -362
rect 492 -358 493 -356
rect 492 -364 493 -362
rect 506 -358 507 -356
rect 506 -364 507 -362
rect 513 -358 514 -356
rect 513 -364 514 -362
rect 520 -358 521 -356
rect 520 -364 521 -362
rect 527 -358 528 -356
rect 527 -364 528 -362
rect 534 -358 535 -356
rect 534 -364 535 -362
rect 541 -358 542 -356
rect 541 -364 542 -362
rect 548 -358 549 -356
rect 548 -364 549 -362
rect 555 -358 556 -356
rect 555 -364 556 -362
rect 562 -358 563 -356
rect 562 -364 563 -362
rect 569 -358 570 -356
rect 569 -364 570 -362
rect 576 -358 577 -356
rect 576 -364 577 -362
rect 583 -358 584 -356
rect 583 -364 584 -362
rect 590 -358 591 -356
rect 590 -364 591 -362
rect 597 -358 598 -356
rect 597 -364 598 -362
rect 604 -358 605 -356
rect 604 -364 605 -362
rect 611 -358 612 -356
rect 611 -364 612 -362
rect 621 -358 622 -356
rect 653 -358 654 -356
rect 656 -358 657 -356
rect 653 -364 654 -362
rect 660 -358 661 -356
rect 660 -364 661 -362
rect 670 -364 671 -362
rect 674 -358 675 -356
rect 674 -364 675 -362
rect 16 -425 17 -423
rect 16 -431 17 -429
rect 33 -425 34 -423
rect 40 -431 41 -429
rect 44 -425 45 -423
rect 44 -431 45 -429
rect 51 -425 52 -423
rect 51 -431 52 -429
rect 61 -431 62 -429
rect 65 -425 66 -423
rect 65 -431 66 -429
rect 72 -425 73 -423
rect 72 -431 73 -429
rect 82 -431 83 -429
rect 86 -425 87 -423
rect 86 -431 87 -429
rect 93 -425 94 -423
rect 93 -431 94 -429
rect 100 -425 101 -423
rect 100 -431 101 -429
rect 107 -425 108 -423
rect 107 -431 108 -429
rect 114 -425 115 -423
rect 117 -425 118 -423
rect 114 -431 115 -429
rect 117 -431 118 -429
rect 121 -425 122 -423
rect 121 -431 122 -429
rect 128 -425 129 -423
rect 128 -431 129 -429
rect 135 -425 136 -423
rect 138 -425 139 -423
rect 142 -425 143 -423
rect 142 -431 143 -429
rect 149 -425 150 -423
rect 149 -431 150 -429
rect 156 -425 157 -423
rect 156 -431 157 -429
rect 163 -425 164 -423
rect 166 -425 167 -423
rect 166 -431 167 -429
rect 170 -425 171 -423
rect 173 -431 174 -429
rect 177 -425 178 -423
rect 177 -431 178 -429
rect 184 -425 185 -423
rect 184 -431 185 -429
rect 191 -425 192 -423
rect 194 -431 195 -429
rect 198 -425 199 -423
rect 198 -431 199 -429
rect 201 -431 202 -429
rect 205 -431 206 -429
rect 215 -425 216 -423
rect 215 -431 216 -429
rect 222 -425 223 -423
rect 222 -431 223 -429
rect 226 -425 227 -423
rect 229 -425 230 -423
rect 226 -431 227 -429
rect 229 -431 230 -429
rect 233 -425 234 -423
rect 233 -431 234 -429
rect 240 -425 241 -423
rect 240 -431 241 -429
rect 247 -425 248 -423
rect 250 -425 251 -423
rect 247 -431 248 -429
rect 254 -425 255 -423
rect 257 -431 258 -429
rect 261 -425 262 -423
rect 264 -425 265 -423
rect 261 -431 262 -429
rect 264 -431 265 -429
rect 268 -425 269 -423
rect 268 -431 269 -429
rect 275 -425 276 -423
rect 275 -431 276 -429
rect 282 -425 283 -423
rect 285 -425 286 -423
rect 282 -431 283 -429
rect 289 -425 290 -423
rect 296 -425 297 -423
rect 296 -431 297 -429
rect 303 -425 304 -423
rect 303 -431 304 -429
rect 310 -431 311 -429
rect 317 -425 318 -423
rect 317 -431 318 -429
rect 320 -431 321 -429
rect 324 -425 325 -423
rect 327 -431 328 -429
rect 331 -425 332 -423
rect 331 -431 332 -429
rect 341 -425 342 -423
rect 338 -431 339 -429
rect 345 -425 346 -423
rect 345 -431 346 -429
rect 352 -425 353 -423
rect 352 -431 353 -429
rect 359 -425 360 -423
rect 362 -425 363 -423
rect 359 -431 360 -429
rect 362 -431 363 -429
rect 366 -425 367 -423
rect 366 -431 367 -429
rect 373 -425 374 -423
rect 373 -431 374 -429
rect 383 -425 384 -423
rect 380 -431 381 -429
rect 383 -431 384 -429
rect 387 -425 388 -423
rect 387 -431 388 -429
rect 390 -431 391 -429
rect 394 -425 395 -423
rect 394 -431 395 -429
rect 401 -425 402 -423
rect 401 -431 402 -429
rect 408 -425 409 -423
rect 408 -431 409 -429
rect 415 -425 416 -423
rect 415 -431 416 -429
rect 422 -425 423 -423
rect 422 -431 423 -429
rect 429 -425 430 -423
rect 429 -431 430 -429
rect 436 -425 437 -423
rect 436 -431 437 -429
rect 443 -425 444 -423
rect 443 -431 444 -429
rect 450 -425 451 -423
rect 450 -431 451 -429
rect 457 -425 458 -423
rect 457 -431 458 -429
rect 464 -425 465 -423
rect 464 -431 465 -429
rect 474 -425 475 -423
rect 471 -431 472 -429
rect 481 -425 482 -423
rect 478 -431 479 -429
rect 485 -425 486 -423
rect 485 -431 486 -429
rect 492 -425 493 -423
rect 492 -431 493 -429
rect 499 -425 500 -423
rect 499 -431 500 -429
rect 506 -425 507 -423
rect 506 -431 507 -429
rect 513 -425 514 -423
rect 513 -431 514 -429
rect 520 -425 521 -423
rect 520 -431 521 -429
rect 527 -425 528 -423
rect 527 -431 528 -429
rect 534 -425 535 -423
rect 534 -431 535 -429
rect 541 -425 542 -423
rect 541 -431 542 -429
rect 544 -431 545 -429
rect 548 -425 549 -423
rect 548 -431 549 -429
rect 555 -425 556 -423
rect 555 -431 556 -429
rect 562 -425 563 -423
rect 562 -431 563 -429
rect 569 -425 570 -423
rect 569 -431 570 -429
rect 576 -425 577 -423
rect 576 -431 577 -429
rect 583 -425 584 -423
rect 583 -431 584 -429
rect 590 -425 591 -423
rect 590 -431 591 -429
rect 597 -425 598 -423
rect 597 -431 598 -429
rect 604 -425 605 -423
rect 604 -431 605 -429
rect 611 -425 612 -423
rect 611 -431 612 -429
rect 618 -425 619 -423
rect 618 -431 619 -429
rect 625 -425 626 -423
rect 625 -431 626 -429
rect 632 -425 633 -423
rect 632 -431 633 -429
rect 639 -425 640 -423
rect 639 -431 640 -429
rect 646 -425 647 -423
rect 646 -431 647 -429
rect 653 -425 654 -423
rect 653 -431 654 -429
rect 660 -425 661 -423
rect 660 -431 661 -429
rect 667 -425 668 -423
rect 667 -431 668 -429
rect 674 -425 675 -423
rect 681 -425 682 -423
rect 681 -431 682 -429
rect 26 -518 27 -516
rect 33 -512 34 -510
rect 30 -518 31 -516
rect 37 -512 38 -510
rect 44 -512 45 -510
rect 44 -518 45 -516
rect 51 -518 52 -516
rect 58 -512 59 -510
rect 58 -518 59 -516
rect 65 -512 66 -510
rect 65 -518 66 -516
rect 72 -512 73 -510
rect 72 -518 73 -516
rect 79 -512 80 -510
rect 79 -518 80 -516
rect 86 -512 87 -510
rect 93 -512 94 -510
rect 93 -518 94 -516
rect 100 -512 101 -510
rect 100 -518 101 -516
rect 110 -512 111 -510
rect 107 -518 108 -516
rect 114 -512 115 -510
rect 114 -518 115 -516
rect 121 -518 122 -516
rect 124 -518 125 -516
rect 128 -512 129 -510
rect 128 -518 129 -516
rect 135 -512 136 -510
rect 135 -518 136 -516
rect 142 -518 143 -516
rect 145 -518 146 -516
rect 149 -512 150 -510
rect 149 -518 150 -516
rect 156 -512 157 -510
rect 156 -518 157 -516
rect 163 -512 164 -510
rect 163 -518 164 -516
rect 173 -518 174 -516
rect 177 -512 178 -510
rect 177 -518 178 -516
rect 184 -512 185 -510
rect 184 -518 185 -516
rect 191 -512 192 -510
rect 191 -518 192 -516
rect 198 -512 199 -510
rect 201 -518 202 -516
rect 205 -512 206 -510
rect 205 -518 206 -516
rect 212 -512 213 -510
rect 215 -512 216 -510
rect 215 -518 216 -516
rect 219 -512 220 -510
rect 219 -518 220 -516
rect 226 -512 227 -510
rect 229 -512 230 -510
rect 233 -512 234 -510
rect 233 -518 234 -516
rect 240 -512 241 -510
rect 243 -512 244 -510
rect 240 -518 241 -516
rect 243 -518 244 -516
rect 247 -512 248 -510
rect 247 -518 248 -516
rect 254 -512 255 -510
rect 257 -512 258 -510
rect 254 -518 255 -516
rect 257 -518 258 -516
rect 261 -512 262 -510
rect 261 -518 262 -516
rect 268 -512 269 -510
rect 271 -512 272 -510
rect 275 -512 276 -510
rect 275 -518 276 -516
rect 282 -512 283 -510
rect 282 -518 283 -516
rect 285 -518 286 -516
rect 289 -518 290 -516
rect 296 -518 297 -516
rect 299 -518 300 -516
rect 303 -512 304 -510
rect 303 -518 304 -516
rect 310 -512 311 -510
rect 310 -518 311 -516
rect 317 -512 318 -510
rect 320 -512 321 -510
rect 317 -518 318 -516
rect 320 -518 321 -516
rect 327 -512 328 -510
rect 324 -518 325 -516
rect 327 -518 328 -516
rect 331 -512 332 -510
rect 331 -518 332 -516
rect 338 -512 339 -510
rect 338 -518 339 -516
rect 348 -512 349 -510
rect 348 -518 349 -516
rect 352 -512 353 -510
rect 355 -512 356 -510
rect 355 -518 356 -516
rect 359 -512 360 -510
rect 362 -518 363 -516
rect 366 -512 367 -510
rect 366 -518 367 -516
rect 373 -512 374 -510
rect 373 -518 374 -516
rect 380 -512 381 -510
rect 380 -518 381 -516
rect 390 -512 391 -510
rect 387 -518 388 -516
rect 390 -518 391 -516
rect 394 -512 395 -510
rect 394 -518 395 -516
rect 401 -518 402 -516
rect 404 -518 405 -516
rect 408 -512 409 -510
rect 408 -518 409 -516
rect 415 -512 416 -510
rect 415 -518 416 -516
rect 422 -512 423 -510
rect 425 -512 426 -510
rect 425 -518 426 -516
rect 429 -512 430 -510
rect 429 -518 430 -516
rect 439 -512 440 -510
rect 439 -518 440 -516
rect 443 -512 444 -510
rect 443 -518 444 -516
rect 450 -512 451 -510
rect 450 -518 451 -516
rect 457 -512 458 -510
rect 457 -518 458 -516
rect 464 -512 465 -510
rect 464 -518 465 -516
rect 471 -512 472 -510
rect 471 -518 472 -516
rect 478 -512 479 -510
rect 478 -518 479 -516
rect 485 -512 486 -510
rect 485 -518 486 -516
rect 492 -512 493 -510
rect 492 -518 493 -516
rect 499 -512 500 -510
rect 499 -518 500 -516
rect 506 -512 507 -510
rect 506 -518 507 -516
rect 513 -512 514 -510
rect 513 -518 514 -516
rect 520 -512 521 -510
rect 520 -518 521 -516
rect 527 -512 528 -510
rect 527 -518 528 -516
rect 534 -512 535 -510
rect 534 -518 535 -516
rect 541 -512 542 -510
rect 544 -512 545 -510
rect 541 -518 542 -516
rect 548 -512 549 -510
rect 548 -518 549 -516
rect 555 -512 556 -510
rect 555 -518 556 -516
rect 562 -512 563 -510
rect 562 -518 563 -516
rect 569 -512 570 -510
rect 569 -518 570 -516
rect 576 -512 577 -510
rect 576 -518 577 -516
rect 583 -512 584 -510
rect 583 -518 584 -516
rect 590 -512 591 -510
rect 590 -518 591 -516
rect 597 -512 598 -510
rect 597 -518 598 -516
rect 604 -512 605 -510
rect 604 -518 605 -516
rect 611 -512 612 -510
rect 611 -518 612 -516
rect 618 -512 619 -510
rect 618 -518 619 -516
rect 625 -512 626 -510
rect 625 -518 626 -516
rect 632 -512 633 -510
rect 632 -518 633 -516
rect 639 -512 640 -510
rect 639 -518 640 -516
rect 646 -512 647 -510
rect 646 -518 647 -516
rect 653 -512 654 -510
rect 653 -518 654 -516
rect 660 -512 661 -510
rect 660 -518 661 -516
rect 667 -512 668 -510
rect 667 -518 668 -516
rect 674 -512 675 -510
rect 674 -518 675 -516
rect 681 -512 682 -510
rect 681 -518 682 -516
rect 688 -512 689 -510
rect 688 -518 689 -516
rect 695 -512 696 -510
rect 695 -518 696 -516
rect 702 -512 703 -510
rect 702 -518 703 -516
rect 709 -512 710 -510
rect 709 -518 710 -516
rect 16 -599 17 -597
rect 23 -599 24 -597
rect 23 -605 24 -603
rect 30 -599 31 -597
rect 30 -605 31 -603
rect 37 -599 38 -597
rect 37 -605 38 -603
rect 44 -599 45 -597
rect 44 -605 45 -603
rect 54 -599 55 -597
rect 54 -605 55 -603
rect 58 -599 59 -597
rect 58 -605 59 -603
rect 65 -599 66 -597
rect 68 -599 69 -597
rect 65 -605 66 -603
rect 72 -599 73 -597
rect 79 -599 80 -597
rect 79 -605 80 -603
rect 86 -599 87 -597
rect 86 -605 87 -603
rect 93 -599 94 -597
rect 93 -605 94 -603
rect 100 -605 101 -603
rect 103 -605 104 -603
rect 107 -599 108 -597
rect 107 -605 108 -603
rect 114 -599 115 -597
rect 117 -599 118 -597
rect 117 -605 118 -603
rect 121 -599 122 -597
rect 121 -605 122 -603
rect 131 -599 132 -597
rect 128 -605 129 -603
rect 135 -599 136 -597
rect 135 -605 136 -603
rect 142 -599 143 -597
rect 142 -605 143 -603
rect 149 -599 150 -597
rect 149 -605 150 -603
rect 159 -599 160 -597
rect 163 -599 164 -597
rect 163 -605 164 -603
rect 170 -599 171 -597
rect 170 -605 171 -603
rect 177 -599 178 -597
rect 177 -605 178 -603
rect 184 -599 185 -597
rect 184 -605 185 -603
rect 194 -599 195 -597
rect 194 -605 195 -603
rect 198 -599 199 -597
rect 201 -599 202 -597
rect 198 -605 199 -603
rect 201 -605 202 -603
rect 205 -599 206 -597
rect 205 -605 206 -603
rect 212 -599 213 -597
rect 215 -599 216 -597
rect 215 -605 216 -603
rect 219 -599 220 -597
rect 222 -605 223 -603
rect 226 -599 227 -597
rect 226 -605 227 -603
rect 233 -599 234 -597
rect 233 -605 234 -603
rect 240 -599 241 -597
rect 240 -605 241 -603
rect 247 -599 248 -597
rect 247 -605 248 -603
rect 254 -599 255 -597
rect 254 -605 255 -603
rect 261 -599 262 -597
rect 261 -605 262 -603
rect 268 -599 269 -597
rect 268 -605 269 -603
rect 275 -599 276 -597
rect 285 -599 286 -597
rect 285 -605 286 -603
rect 289 -599 290 -597
rect 289 -605 290 -603
rect 296 -599 297 -597
rect 296 -605 297 -603
rect 306 -599 307 -597
rect 303 -605 304 -603
rect 310 -599 311 -597
rect 310 -605 311 -603
rect 317 -599 318 -597
rect 320 -599 321 -597
rect 317 -605 318 -603
rect 320 -605 321 -603
rect 324 -599 325 -597
rect 324 -605 325 -603
rect 331 -599 332 -597
rect 331 -605 332 -603
rect 338 -599 339 -597
rect 345 -599 346 -597
rect 348 -605 349 -603
rect 352 -599 353 -597
rect 352 -605 353 -603
rect 359 -599 360 -597
rect 359 -605 360 -603
rect 366 -599 367 -597
rect 366 -605 367 -603
rect 373 -605 374 -603
rect 376 -605 377 -603
rect 380 -599 381 -597
rect 380 -605 381 -603
rect 387 -599 388 -597
rect 387 -605 388 -603
rect 394 -599 395 -597
rect 394 -605 395 -603
rect 401 -599 402 -597
rect 401 -605 402 -603
rect 408 -599 409 -597
rect 411 -599 412 -597
rect 408 -605 409 -603
rect 411 -605 412 -603
rect 418 -599 419 -597
rect 418 -605 419 -603
rect 422 -599 423 -597
rect 422 -605 423 -603
rect 429 -599 430 -597
rect 429 -605 430 -603
rect 436 -599 437 -597
rect 439 -599 440 -597
rect 439 -605 440 -603
rect 443 -599 444 -597
rect 446 -605 447 -603
rect 450 -599 451 -597
rect 450 -605 451 -603
rect 457 -599 458 -597
rect 460 -599 461 -597
rect 457 -605 458 -603
rect 464 -599 465 -597
rect 464 -605 465 -603
rect 471 -605 472 -603
rect 478 -599 479 -597
rect 478 -605 479 -603
rect 485 -599 486 -597
rect 485 -605 486 -603
rect 492 -599 493 -597
rect 495 -599 496 -597
rect 492 -605 493 -603
rect 502 -599 503 -597
rect 499 -605 500 -603
rect 506 -599 507 -597
rect 506 -605 507 -603
rect 513 -599 514 -597
rect 513 -605 514 -603
rect 520 -599 521 -597
rect 520 -605 521 -603
rect 527 -599 528 -597
rect 527 -605 528 -603
rect 534 -599 535 -597
rect 534 -605 535 -603
rect 541 -599 542 -597
rect 541 -605 542 -603
rect 548 -599 549 -597
rect 548 -605 549 -603
rect 558 -599 559 -597
rect 555 -605 556 -603
rect 562 -599 563 -597
rect 562 -605 563 -603
rect 569 -599 570 -597
rect 569 -605 570 -603
rect 576 -599 577 -597
rect 576 -605 577 -603
rect 583 -599 584 -597
rect 583 -605 584 -603
rect 590 -599 591 -597
rect 590 -605 591 -603
rect 597 -599 598 -597
rect 597 -605 598 -603
rect 604 -599 605 -597
rect 604 -605 605 -603
rect 611 -599 612 -597
rect 611 -605 612 -603
rect 618 -599 619 -597
rect 618 -605 619 -603
rect 625 -599 626 -597
rect 625 -605 626 -603
rect 632 -599 633 -597
rect 632 -605 633 -603
rect 639 -599 640 -597
rect 639 -605 640 -603
rect 646 -599 647 -597
rect 646 -605 647 -603
rect 653 -599 654 -597
rect 653 -605 654 -603
rect 660 -599 661 -597
rect 660 -605 661 -603
rect 667 -599 668 -597
rect 667 -605 668 -603
rect 674 -599 675 -597
rect 674 -605 675 -603
rect 681 -599 682 -597
rect 681 -605 682 -603
rect 709 -599 710 -597
rect 709 -605 710 -603
rect 19 -678 20 -676
rect 23 -678 24 -676
rect 30 -684 31 -682
rect 37 -678 38 -676
rect 37 -684 38 -682
rect 44 -678 45 -676
rect 44 -684 45 -682
rect 51 -678 52 -676
rect 51 -684 52 -682
rect 58 -678 59 -676
rect 61 -684 62 -682
rect 65 -678 66 -676
rect 65 -684 66 -682
rect 72 -678 73 -676
rect 75 -678 76 -676
rect 72 -684 73 -682
rect 79 -678 80 -676
rect 79 -684 80 -682
rect 86 -678 87 -676
rect 86 -684 87 -682
rect 93 -678 94 -676
rect 93 -684 94 -682
rect 100 -678 101 -676
rect 100 -684 101 -682
rect 107 -678 108 -676
rect 107 -684 108 -682
rect 114 -678 115 -676
rect 114 -684 115 -682
rect 124 -678 125 -676
rect 121 -684 122 -682
rect 124 -684 125 -682
rect 128 -684 129 -682
rect 135 -678 136 -676
rect 135 -684 136 -682
rect 142 -678 143 -676
rect 142 -684 143 -682
rect 145 -684 146 -682
rect 149 -678 150 -676
rect 149 -684 150 -682
rect 159 -678 160 -676
rect 156 -684 157 -682
rect 159 -684 160 -682
rect 163 -678 164 -676
rect 163 -684 164 -682
rect 170 -678 171 -676
rect 170 -684 171 -682
rect 177 -678 178 -676
rect 177 -684 178 -682
rect 187 -678 188 -676
rect 184 -684 185 -682
rect 187 -684 188 -682
rect 191 -678 192 -676
rect 191 -684 192 -682
rect 198 -678 199 -676
rect 201 -678 202 -676
rect 201 -684 202 -682
rect 205 -678 206 -676
rect 205 -684 206 -682
rect 212 -678 213 -676
rect 212 -684 213 -682
rect 219 -678 220 -676
rect 222 -678 223 -676
rect 222 -684 223 -682
rect 226 -678 227 -676
rect 226 -684 227 -682
rect 233 -678 234 -676
rect 233 -684 234 -682
rect 240 -678 241 -676
rect 240 -684 241 -682
rect 247 -678 248 -676
rect 247 -684 248 -682
rect 254 -678 255 -676
rect 254 -684 255 -682
rect 261 -678 262 -676
rect 261 -684 262 -682
rect 268 -678 269 -676
rect 268 -684 269 -682
rect 275 -678 276 -676
rect 275 -684 276 -682
rect 278 -684 279 -682
rect 282 -678 283 -676
rect 285 -678 286 -676
rect 282 -684 283 -682
rect 289 -678 290 -676
rect 289 -684 290 -682
rect 296 -678 297 -676
rect 296 -684 297 -682
rect 303 -678 304 -676
rect 303 -684 304 -682
rect 310 -678 311 -676
rect 310 -684 311 -682
rect 317 -678 318 -676
rect 320 -684 321 -682
rect 324 -678 325 -676
rect 327 -684 328 -682
rect 331 -678 332 -676
rect 331 -684 332 -682
rect 338 -678 339 -676
rect 338 -684 339 -682
rect 345 -684 346 -682
rect 348 -684 349 -682
rect 355 -678 356 -676
rect 355 -684 356 -682
rect 359 -678 360 -676
rect 359 -684 360 -682
rect 366 -678 367 -676
rect 366 -684 367 -682
rect 373 -678 374 -676
rect 373 -684 374 -682
rect 380 -678 381 -676
rect 380 -684 381 -682
rect 387 -678 388 -676
rect 387 -684 388 -682
rect 394 -678 395 -676
rect 394 -684 395 -682
rect 397 -684 398 -682
rect 401 -678 402 -676
rect 404 -678 405 -676
rect 401 -684 402 -682
rect 404 -684 405 -682
rect 408 -678 409 -676
rect 408 -684 409 -682
rect 415 -678 416 -676
rect 415 -684 416 -682
rect 422 -678 423 -676
rect 425 -678 426 -676
rect 429 -678 430 -676
rect 429 -684 430 -682
rect 439 -678 440 -676
rect 436 -684 437 -682
rect 439 -684 440 -682
rect 443 -678 444 -676
rect 443 -684 444 -682
rect 453 -678 454 -676
rect 453 -684 454 -682
rect 457 -678 458 -676
rect 460 -678 461 -676
rect 457 -684 458 -682
rect 464 -678 465 -676
rect 467 -678 468 -676
rect 467 -684 468 -682
rect 478 -678 479 -676
rect 481 -684 482 -682
rect 485 -678 486 -676
rect 485 -684 486 -682
rect 495 -684 496 -682
rect 499 -678 500 -676
rect 499 -684 500 -682
rect 506 -684 507 -682
rect 509 -684 510 -682
rect 513 -678 514 -676
rect 513 -684 514 -682
rect 520 -678 521 -676
rect 520 -684 521 -682
rect 527 -678 528 -676
rect 527 -684 528 -682
rect 534 -678 535 -676
rect 534 -684 535 -682
rect 541 -678 542 -676
rect 541 -684 542 -682
rect 548 -678 549 -676
rect 548 -684 549 -682
rect 555 -678 556 -676
rect 555 -684 556 -682
rect 562 -678 563 -676
rect 562 -684 563 -682
rect 569 -678 570 -676
rect 569 -684 570 -682
rect 576 -678 577 -676
rect 576 -684 577 -682
rect 583 -678 584 -676
rect 586 -684 587 -682
rect 590 -678 591 -676
rect 590 -684 591 -682
rect 597 -678 598 -676
rect 597 -684 598 -682
rect 604 -678 605 -676
rect 604 -684 605 -682
rect 611 -678 612 -676
rect 611 -684 612 -682
rect 618 -678 619 -676
rect 618 -684 619 -682
rect 625 -678 626 -676
rect 625 -684 626 -682
rect 632 -678 633 -676
rect 632 -684 633 -682
rect 639 -678 640 -676
rect 639 -684 640 -682
rect 646 -678 647 -676
rect 646 -684 647 -682
rect 653 -678 654 -676
rect 653 -684 654 -682
rect 660 -678 661 -676
rect 660 -684 661 -682
rect 667 -678 668 -676
rect 667 -684 668 -682
rect 674 -678 675 -676
rect 674 -684 675 -682
rect 681 -678 682 -676
rect 681 -684 682 -682
rect 688 -678 689 -676
rect 688 -684 689 -682
rect 695 -678 696 -676
rect 695 -684 696 -682
rect 702 -678 703 -676
rect 702 -684 703 -682
rect 709 -678 710 -676
rect 709 -684 710 -682
rect 716 -678 717 -676
rect 716 -684 717 -682
rect 723 -678 724 -676
rect 723 -684 724 -682
rect 730 -678 731 -676
rect 730 -684 731 -682
rect 737 -678 738 -676
rect 737 -684 738 -682
rect 744 -678 745 -676
rect 744 -684 745 -682
rect 751 -678 752 -676
rect 751 -684 752 -682
rect 758 -678 759 -676
rect 758 -684 759 -682
rect 765 -678 766 -676
rect 765 -684 766 -682
rect 772 -678 773 -676
rect 772 -684 773 -682
rect 16 -763 17 -761
rect 19 -769 20 -767
rect 23 -769 24 -767
rect 30 -763 31 -761
rect 37 -763 38 -761
rect 37 -769 38 -767
rect 44 -763 45 -761
rect 44 -769 45 -767
rect 54 -763 55 -761
rect 58 -763 59 -761
rect 58 -769 59 -767
rect 65 -763 66 -761
rect 65 -769 66 -767
rect 72 -763 73 -761
rect 72 -769 73 -767
rect 79 -763 80 -761
rect 79 -769 80 -767
rect 86 -763 87 -761
rect 89 -763 90 -761
rect 86 -769 87 -767
rect 89 -769 90 -767
rect 93 -763 94 -761
rect 96 -763 97 -761
rect 96 -769 97 -767
rect 100 -763 101 -761
rect 100 -769 101 -767
rect 107 -763 108 -761
rect 107 -769 108 -767
rect 114 -763 115 -761
rect 117 -769 118 -767
rect 124 -763 125 -761
rect 121 -769 122 -767
rect 131 -763 132 -761
rect 128 -769 129 -767
rect 135 -763 136 -761
rect 135 -769 136 -767
rect 142 -763 143 -761
rect 142 -769 143 -767
rect 149 -763 150 -761
rect 149 -769 150 -767
rect 152 -769 153 -767
rect 156 -763 157 -761
rect 156 -769 157 -767
rect 163 -763 164 -761
rect 163 -769 164 -767
rect 170 -763 171 -761
rect 170 -769 171 -767
rect 177 -763 178 -761
rect 177 -769 178 -767
rect 184 -763 185 -761
rect 184 -769 185 -767
rect 191 -763 192 -761
rect 191 -769 192 -767
rect 201 -763 202 -761
rect 198 -769 199 -767
rect 201 -769 202 -767
rect 205 -763 206 -761
rect 212 -763 213 -761
rect 212 -769 213 -767
rect 222 -763 223 -761
rect 219 -769 220 -767
rect 222 -769 223 -767
rect 226 -763 227 -761
rect 226 -769 227 -767
rect 233 -763 234 -761
rect 233 -769 234 -767
rect 240 -763 241 -761
rect 240 -769 241 -767
rect 243 -769 244 -767
rect 247 -763 248 -761
rect 247 -769 248 -767
rect 254 -763 255 -761
rect 254 -769 255 -767
rect 261 -763 262 -761
rect 261 -769 262 -767
rect 268 -763 269 -761
rect 268 -769 269 -767
rect 275 -763 276 -761
rect 275 -769 276 -767
rect 282 -763 283 -761
rect 282 -769 283 -767
rect 289 -763 290 -761
rect 292 -763 293 -761
rect 289 -769 290 -767
rect 292 -769 293 -767
rect 296 -763 297 -761
rect 296 -769 297 -767
rect 303 -763 304 -761
rect 306 -763 307 -761
rect 306 -769 307 -767
rect 313 -763 314 -761
rect 310 -769 311 -767
rect 320 -763 321 -761
rect 317 -769 318 -767
rect 320 -769 321 -767
rect 324 -763 325 -761
rect 324 -769 325 -767
rect 331 -763 332 -761
rect 331 -769 332 -767
rect 338 -763 339 -761
rect 338 -769 339 -767
rect 345 -763 346 -761
rect 348 -763 349 -761
rect 352 -763 353 -761
rect 355 -763 356 -761
rect 352 -769 353 -767
rect 355 -769 356 -767
rect 362 -763 363 -761
rect 359 -769 360 -767
rect 366 -763 367 -761
rect 366 -769 367 -767
rect 373 -763 374 -761
rect 373 -769 374 -767
rect 383 -763 384 -761
rect 380 -769 381 -767
rect 387 -763 388 -761
rect 387 -769 388 -767
rect 394 -763 395 -761
rect 397 -763 398 -761
rect 397 -769 398 -767
rect 401 -763 402 -761
rect 401 -769 402 -767
rect 408 -763 409 -761
rect 408 -769 409 -767
rect 415 -763 416 -761
rect 415 -769 416 -767
rect 422 -763 423 -761
rect 422 -769 423 -767
rect 429 -763 430 -761
rect 429 -769 430 -767
rect 432 -769 433 -767
rect 436 -763 437 -761
rect 439 -763 440 -761
rect 446 -763 447 -761
rect 443 -769 444 -767
rect 446 -769 447 -767
rect 450 -763 451 -761
rect 450 -769 451 -767
rect 457 -763 458 -761
rect 457 -769 458 -767
rect 464 -763 465 -761
rect 464 -769 465 -767
rect 471 -763 472 -761
rect 471 -769 472 -767
rect 478 -763 479 -761
rect 481 -763 482 -761
rect 488 -763 489 -761
rect 488 -769 489 -767
rect 492 -763 493 -761
rect 492 -769 493 -767
rect 499 -763 500 -761
rect 499 -769 500 -767
rect 506 -763 507 -761
rect 506 -769 507 -767
rect 513 -763 514 -761
rect 513 -769 514 -767
rect 520 -763 521 -761
rect 520 -769 521 -767
rect 527 -763 528 -761
rect 527 -769 528 -767
rect 534 -763 535 -761
rect 534 -769 535 -767
rect 537 -769 538 -767
rect 541 -763 542 -761
rect 541 -769 542 -767
rect 548 -763 549 -761
rect 548 -769 549 -767
rect 555 -763 556 -761
rect 555 -769 556 -767
rect 562 -763 563 -761
rect 562 -769 563 -767
rect 569 -763 570 -761
rect 569 -769 570 -767
rect 576 -763 577 -761
rect 576 -769 577 -767
rect 583 -763 584 -761
rect 583 -769 584 -767
rect 590 -763 591 -761
rect 590 -769 591 -767
rect 597 -763 598 -761
rect 597 -769 598 -767
rect 604 -763 605 -761
rect 604 -769 605 -767
rect 611 -763 612 -761
rect 611 -769 612 -767
rect 621 -763 622 -761
rect 621 -769 622 -767
rect 625 -763 626 -761
rect 625 -769 626 -767
rect 632 -763 633 -761
rect 632 -769 633 -767
rect 639 -763 640 -761
rect 639 -769 640 -767
rect 646 -763 647 -761
rect 646 -769 647 -767
rect 653 -763 654 -761
rect 653 -769 654 -767
rect 660 -763 661 -761
rect 660 -769 661 -767
rect 667 -763 668 -761
rect 667 -769 668 -767
rect 674 -763 675 -761
rect 674 -769 675 -767
rect 681 -763 682 -761
rect 681 -769 682 -767
rect 688 -763 689 -761
rect 688 -769 689 -767
rect 695 -763 696 -761
rect 695 -769 696 -767
rect 702 -763 703 -761
rect 702 -769 703 -767
rect 709 -763 710 -761
rect 709 -769 710 -767
rect 716 -763 717 -761
rect 716 -769 717 -767
rect 723 -763 724 -761
rect 723 -769 724 -767
rect 733 -763 734 -761
rect 737 -763 738 -761
rect 737 -769 738 -767
rect 744 -763 745 -761
rect 744 -769 745 -767
rect 751 -763 752 -761
rect 751 -769 752 -767
rect 758 -763 759 -761
rect 758 -769 759 -767
rect 765 -763 766 -761
rect 765 -769 766 -767
rect 772 -763 773 -761
rect 772 -769 773 -767
rect 779 -763 780 -761
rect 779 -769 780 -767
rect 786 -763 787 -761
rect 786 -769 787 -767
rect 793 -763 794 -761
rect 793 -769 794 -767
rect 849 -763 850 -761
rect 849 -769 850 -767
rect 19 -858 20 -856
rect 23 -852 24 -850
rect 23 -858 24 -856
rect 30 -852 31 -850
rect 30 -858 31 -856
rect 37 -852 38 -850
rect 40 -852 41 -850
rect 44 -852 45 -850
rect 44 -858 45 -856
rect 54 -852 55 -850
rect 51 -858 52 -856
rect 58 -852 59 -850
rect 58 -858 59 -856
rect 65 -852 66 -850
rect 65 -858 66 -856
rect 72 -852 73 -850
rect 72 -858 73 -856
rect 75 -858 76 -856
rect 79 -852 80 -850
rect 79 -858 80 -856
rect 86 -852 87 -850
rect 89 -852 90 -850
rect 86 -858 87 -856
rect 93 -852 94 -850
rect 93 -858 94 -856
rect 100 -852 101 -850
rect 100 -858 101 -856
rect 103 -858 104 -856
rect 107 -852 108 -850
rect 107 -858 108 -856
rect 114 -852 115 -850
rect 114 -858 115 -856
rect 121 -852 122 -850
rect 121 -858 122 -856
rect 128 -852 129 -850
rect 128 -858 129 -856
rect 135 -852 136 -850
rect 135 -858 136 -856
rect 142 -852 143 -850
rect 142 -858 143 -856
rect 145 -858 146 -856
rect 149 -852 150 -850
rect 152 -852 153 -850
rect 156 -852 157 -850
rect 159 -852 160 -850
rect 156 -858 157 -856
rect 159 -858 160 -856
rect 163 -852 164 -850
rect 166 -852 167 -850
rect 163 -858 164 -856
rect 170 -852 171 -850
rect 170 -858 171 -856
rect 177 -852 178 -850
rect 177 -858 178 -856
rect 184 -852 185 -850
rect 184 -858 185 -856
rect 191 -852 192 -850
rect 191 -858 192 -856
rect 198 -852 199 -850
rect 198 -858 199 -856
rect 205 -858 206 -856
rect 212 -852 213 -850
rect 212 -858 213 -856
rect 219 -852 220 -850
rect 219 -858 220 -856
rect 226 -852 227 -850
rect 226 -858 227 -856
rect 233 -852 234 -850
rect 233 -858 234 -856
rect 240 -852 241 -850
rect 243 -852 244 -850
rect 240 -858 241 -856
rect 250 -852 251 -850
rect 254 -852 255 -850
rect 254 -858 255 -856
rect 261 -858 262 -856
rect 264 -858 265 -856
rect 268 -852 269 -850
rect 268 -858 269 -856
rect 275 -852 276 -850
rect 275 -858 276 -856
rect 282 -852 283 -850
rect 282 -858 283 -856
rect 289 -852 290 -850
rect 289 -858 290 -856
rect 296 -852 297 -850
rect 299 -852 300 -850
rect 296 -858 297 -856
rect 306 -852 307 -850
rect 303 -858 304 -856
rect 306 -858 307 -856
rect 310 -852 311 -850
rect 310 -858 311 -856
rect 317 -852 318 -850
rect 317 -858 318 -856
rect 324 -852 325 -850
rect 327 -852 328 -850
rect 327 -858 328 -856
rect 331 -852 332 -850
rect 331 -858 332 -856
rect 334 -858 335 -856
rect 338 -852 339 -850
rect 338 -858 339 -856
rect 345 -852 346 -850
rect 345 -858 346 -856
rect 352 -852 353 -850
rect 352 -858 353 -856
rect 359 -852 360 -850
rect 362 -852 363 -850
rect 359 -858 360 -856
rect 362 -858 363 -856
rect 366 -852 367 -850
rect 366 -858 367 -856
rect 373 -852 374 -850
rect 373 -858 374 -856
rect 383 -852 384 -850
rect 380 -858 381 -856
rect 387 -852 388 -850
rect 387 -858 388 -856
rect 394 -852 395 -850
rect 397 -852 398 -850
rect 401 -852 402 -850
rect 401 -858 402 -856
rect 408 -852 409 -850
rect 411 -852 412 -850
rect 411 -858 412 -856
rect 415 -852 416 -850
rect 415 -858 416 -856
rect 422 -852 423 -850
rect 422 -858 423 -856
rect 429 -852 430 -850
rect 432 -852 433 -850
rect 429 -858 430 -856
rect 436 -852 437 -850
rect 439 -858 440 -856
rect 446 -852 447 -850
rect 446 -858 447 -856
rect 450 -852 451 -850
rect 457 -852 458 -850
rect 460 -852 461 -850
rect 460 -858 461 -856
rect 464 -852 465 -850
rect 467 -852 468 -850
rect 471 -852 472 -850
rect 471 -858 472 -856
rect 478 -852 479 -850
rect 478 -858 479 -856
rect 485 -852 486 -850
rect 485 -858 486 -856
rect 492 -852 493 -850
rect 492 -858 493 -856
rect 499 -852 500 -850
rect 499 -858 500 -856
rect 506 -852 507 -850
rect 506 -858 507 -856
rect 513 -852 514 -850
rect 516 -852 517 -850
rect 516 -858 517 -856
rect 520 -852 521 -850
rect 520 -858 521 -856
rect 527 -852 528 -850
rect 527 -858 528 -856
rect 534 -852 535 -850
rect 534 -858 535 -856
rect 541 -852 542 -850
rect 541 -858 542 -856
rect 548 -852 549 -850
rect 548 -858 549 -856
rect 555 -852 556 -850
rect 555 -858 556 -856
rect 562 -852 563 -850
rect 562 -858 563 -856
rect 569 -852 570 -850
rect 569 -858 570 -856
rect 576 -852 577 -850
rect 576 -858 577 -856
rect 583 -852 584 -850
rect 583 -858 584 -856
rect 590 -852 591 -850
rect 590 -858 591 -856
rect 597 -852 598 -850
rect 597 -858 598 -856
rect 604 -852 605 -850
rect 604 -858 605 -856
rect 611 -852 612 -850
rect 611 -858 612 -856
rect 618 -852 619 -850
rect 618 -858 619 -856
rect 625 -852 626 -850
rect 625 -858 626 -856
rect 632 -852 633 -850
rect 632 -858 633 -856
rect 639 -852 640 -850
rect 639 -858 640 -856
rect 646 -852 647 -850
rect 646 -858 647 -856
rect 653 -852 654 -850
rect 653 -858 654 -856
rect 660 -852 661 -850
rect 660 -858 661 -856
rect 667 -852 668 -850
rect 667 -858 668 -856
rect 674 -852 675 -850
rect 674 -858 675 -856
rect 681 -852 682 -850
rect 681 -858 682 -856
rect 688 -852 689 -850
rect 688 -858 689 -856
rect 695 -852 696 -850
rect 695 -858 696 -856
rect 702 -852 703 -850
rect 702 -858 703 -856
rect 709 -852 710 -850
rect 709 -858 710 -856
rect 716 -852 717 -850
rect 716 -858 717 -856
rect 723 -852 724 -850
rect 723 -858 724 -856
rect 730 -852 731 -850
rect 730 -858 731 -856
rect 737 -852 738 -850
rect 737 -858 738 -856
rect 744 -852 745 -850
rect 744 -858 745 -856
rect 751 -852 752 -850
rect 751 -858 752 -856
rect 758 -852 759 -850
rect 758 -858 759 -856
rect 765 -852 766 -850
rect 765 -858 766 -856
rect 772 -852 773 -850
rect 772 -858 773 -856
rect 779 -852 780 -850
rect 779 -858 780 -856
rect 786 -852 787 -850
rect 786 -858 787 -856
rect 800 -852 801 -850
rect 800 -858 801 -856
rect 807 -852 808 -850
rect 807 -858 808 -856
rect 814 -852 815 -850
rect 814 -858 815 -856
rect 821 -852 822 -850
rect 821 -858 822 -856
rect 828 -852 829 -850
rect 828 -858 829 -856
rect 835 -852 836 -850
rect 835 -858 836 -856
rect 842 -852 843 -850
rect 842 -858 843 -856
rect 849 -852 850 -850
rect 849 -858 850 -856
rect 856 -852 857 -850
rect 856 -858 857 -856
rect 863 -852 864 -850
rect 863 -858 864 -856
rect 870 -852 871 -850
rect 870 -858 871 -856
rect 940 -852 941 -850
rect 940 -858 941 -856
rect 9 -929 10 -927
rect 9 -935 10 -933
rect 16 -929 17 -927
rect 16 -935 17 -933
rect 23 -929 24 -927
rect 23 -935 24 -933
rect 30 -929 31 -927
rect 30 -935 31 -933
rect 40 -929 41 -927
rect 40 -935 41 -933
rect 44 -929 45 -927
rect 44 -935 45 -933
rect 51 -929 52 -927
rect 54 -929 55 -927
rect 58 -929 59 -927
rect 58 -935 59 -933
rect 65 -935 66 -933
rect 72 -929 73 -927
rect 72 -935 73 -933
rect 79 -929 80 -927
rect 82 -929 83 -927
rect 82 -935 83 -933
rect 86 -929 87 -927
rect 86 -935 87 -933
rect 93 -929 94 -927
rect 93 -935 94 -933
rect 100 -929 101 -927
rect 100 -935 101 -933
rect 107 -929 108 -927
rect 107 -935 108 -933
rect 114 -929 115 -927
rect 114 -935 115 -933
rect 124 -929 125 -927
rect 121 -935 122 -933
rect 124 -935 125 -933
rect 128 -929 129 -927
rect 128 -935 129 -933
rect 135 -929 136 -927
rect 135 -935 136 -933
rect 142 -929 143 -927
rect 142 -935 143 -933
rect 149 -929 150 -927
rect 152 -935 153 -933
rect 156 -929 157 -927
rect 156 -935 157 -933
rect 163 -929 164 -927
rect 166 -929 167 -927
rect 170 -929 171 -927
rect 170 -935 171 -933
rect 177 -929 178 -927
rect 177 -935 178 -933
rect 184 -929 185 -927
rect 184 -935 185 -933
rect 191 -929 192 -927
rect 191 -935 192 -933
rect 198 -929 199 -927
rect 201 -929 202 -927
rect 201 -935 202 -933
rect 205 -929 206 -927
rect 208 -935 209 -933
rect 215 -929 216 -927
rect 215 -935 216 -933
rect 219 -929 220 -927
rect 222 -929 223 -927
rect 226 -929 227 -927
rect 226 -935 227 -933
rect 233 -929 234 -927
rect 233 -935 234 -933
rect 240 -929 241 -927
rect 240 -935 241 -933
rect 250 -929 251 -927
rect 247 -935 248 -933
rect 254 -929 255 -927
rect 254 -935 255 -933
rect 261 -929 262 -927
rect 261 -935 262 -933
rect 268 -929 269 -927
rect 268 -935 269 -933
rect 278 -929 279 -927
rect 278 -935 279 -933
rect 282 -929 283 -927
rect 285 -935 286 -933
rect 289 -929 290 -927
rect 289 -935 290 -933
rect 299 -929 300 -927
rect 296 -935 297 -933
rect 299 -935 300 -933
rect 303 -929 304 -927
rect 303 -935 304 -933
rect 310 -929 311 -927
rect 310 -935 311 -933
rect 317 -929 318 -927
rect 317 -935 318 -933
rect 324 -929 325 -927
rect 324 -935 325 -933
rect 331 -929 332 -927
rect 331 -935 332 -933
rect 338 -929 339 -927
rect 341 -929 342 -927
rect 338 -935 339 -933
rect 345 -929 346 -927
rect 348 -929 349 -927
rect 345 -935 346 -933
rect 348 -935 349 -933
rect 352 -935 353 -933
rect 359 -929 360 -927
rect 359 -935 360 -933
rect 366 -929 367 -927
rect 366 -935 367 -933
rect 373 -929 374 -927
rect 373 -935 374 -933
rect 380 -929 381 -927
rect 380 -935 381 -933
rect 387 -929 388 -927
rect 387 -935 388 -933
rect 394 -935 395 -933
rect 401 -929 402 -927
rect 404 -929 405 -927
rect 401 -935 402 -933
rect 404 -935 405 -933
rect 408 -929 409 -927
rect 408 -935 409 -933
rect 415 -929 416 -927
rect 415 -935 416 -933
rect 422 -929 423 -927
rect 422 -935 423 -933
rect 429 -929 430 -927
rect 429 -935 430 -933
rect 436 -929 437 -927
rect 436 -935 437 -933
rect 443 -929 444 -927
rect 446 -929 447 -927
rect 443 -935 444 -933
rect 446 -935 447 -933
rect 453 -929 454 -927
rect 450 -935 451 -933
rect 453 -935 454 -933
rect 457 -929 458 -927
rect 457 -935 458 -933
rect 464 -929 465 -927
rect 467 -929 468 -927
rect 471 -929 472 -927
rect 471 -935 472 -933
rect 478 -929 479 -927
rect 478 -935 479 -933
rect 485 -929 486 -927
rect 485 -935 486 -933
rect 492 -929 493 -927
rect 492 -935 493 -933
rect 499 -929 500 -927
rect 499 -935 500 -933
rect 506 -929 507 -927
rect 506 -935 507 -933
rect 509 -935 510 -933
rect 516 -929 517 -927
rect 513 -935 514 -933
rect 516 -935 517 -933
rect 520 -929 521 -927
rect 520 -935 521 -933
rect 527 -929 528 -927
rect 527 -935 528 -933
rect 534 -929 535 -927
rect 534 -935 535 -933
rect 541 -935 542 -933
rect 548 -929 549 -927
rect 548 -935 549 -933
rect 555 -929 556 -927
rect 555 -935 556 -933
rect 562 -929 563 -927
rect 562 -935 563 -933
rect 569 -929 570 -927
rect 569 -935 570 -933
rect 576 -929 577 -927
rect 576 -935 577 -933
rect 583 -929 584 -927
rect 583 -935 584 -933
rect 590 -929 591 -927
rect 593 -929 594 -927
rect 590 -935 591 -933
rect 597 -929 598 -927
rect 597 -935 598 -933
rect 604 -929 605 -927
rect 604 -935 605 -933
rect 611 -929 612 -927
rect 611 -935 612 -933
rect 618 -929 619 -927
rect 618 -935 619 -933
rect 625 -929 626 -927
rect 625 -935 626 -933
rect 632 -929 633 -927
rect 632 -935 633 -933
rect 639 -929 640 -927
rect 639 -935 640 -933
rect 646 -929 647 -927
rect 646 -935 647 -933
rect 653 -929 654 -927
rect 653 -935 654 -933
rect 660 -929 661 -927
rect 660 -935 661 -933
rect 667 -929 668 -927
rect 667 -935 668 -933
rect 674 -929 675 -927
rect 674 -935 675 -933
rect 681 -929 682 -927
rect 681 -935 682 -933
rect 688 -929 689 -927
rect 688 -935 689 -933
rect 695 -929 696 -927
rect 695 -935 696 -933
rect 702 -929 703 -927
rect 702 -935 703 -933
rect 709 -929 710 -927
rect 709 -935 710 -933
rect 716 -929 717 -927
rect 716 -935 717 -933
rect 723 -929 724 -927
rect 723 -935 724 -933
rect 730 -929 731 -927
rect 730 -935 731 -933
rect 737 -929 738 -927
rect 737 -935 738 -933
rect 744 -929 745 -927
rect 744 -935 745 -933
rect 751 -929 752 -927
rect 751 -935 752 -933
rect 758 -929 759 -927
rect 758 -935 759 -933
rect 765 -929 766 -927
rect 765 -935 766 -933
rect 772 -929 773 -927
rect 772 -935 773 -933
rect 779 -929 780 -927
rect 779 -935 780 -933
rect 786 -929 787 -927
rect 786 -935 787 -933
rect 793 -929 794 -927
rect 793 -935 794 -933
rect 800 -929 801 -927
rect 800 -935 801 -933
rect 807 -929 808 -927
rect 807 -935 808 -933
rect 814 -929 815 -927
rect 814 -935 815 -933
rect 821 -929 822 -927
rect 821 -935 822 -933
rect 828 -929 829 -927
rect 831 -929 832 -927
rect 828 -935 829 -933
rect 835 -929 836 -927
rect 835 -935 836 -933
rect 842 -929 843 -927
rect 842 -935 843 -933
rect 849 -929 850 -927
rect 2 -1008 3 -1006
rect 2 -1014 3 -1012
rect 9 -1008 10 -1006
rect 9 -1014 10 -1012
rect 19 -1014 20 -1012
rect 23 -1008 24 -1006
rect 23 -1014 24 -1012
rect 33 -1014 34 -1012
rect 37 -1008 38 -1006
rect 37 -1014 38 -1012
rect 44 -1008 45 -1006
rect 44 -1014 45 -1012
rect 51 -1008 52 -1006
rect 51 -1014 52 -1012
rect 58 -1008 59 -1006
rect 61 -1008 62 -1006
rect 65 -1008 66 -1006
rect 65 -1014 66 -1012
rect 72 -1008 73 -1006
rect 72 -1014 73 -1012
rect 79 -1008 80 -1006
rect 79 -1014 80 -1012
rect 86 -1008 87 -1006
rect 86 -1014 87 -1012
rect 93 -1008 94 -1006
rect 93 -1014 94 -1012
rect 100 -1014 101 -1012
rect 107 -1008 108 -1006
rect 107 -1014 108 -1012
rect 114 -1008 115 -1006
rect 117 -1008 118 -1006
rect 114 -1014 115 -1012
rect 117 -1014 118 -1012
rect 121 -1008 122 -1006
rect 128 -1008 129 -1006
rect 131 -1008 132 -1006
rect 128 -1014 129 -1012
rect 135 -1008 136 -1006
rect 135 -1014 136 -1012
rect 142 -1008 143 -1006
rect 142 -1014 143 -1012
rect 149 -1008 150 -1006
rect 149 -1014 150 -1012
rect 156 -1008 157 -1006
rect 163 -1008 164 -1006
rect 163 -1014 164 -1012
rect 170 -1008 171 -1006
rect 173 -1008 174 -1006
rect 170 -1014 171 -1012
rect 177 -1008 178 -1006
rect 177 -1014 178 -1012
rect 184 -1008 185 -1006
rect 184 -1014 185 -1012
rect 194 -1008 195 -1006
rect 191 -1014 192 -1012
rect 194 -1014 195 -1012
rect 201 -1008 202 -1006
rect 201 -1014 202 -1012
rect 205 -1008 206 -1006
rect 205 -1014 206 -1012
rect 212 -1008 213 -1006
rect 212 -1014 213 -1012
rect 219 -1008 220 -1006
rect 222 -1008 223 -1006
rect 219 -1014 220 -1012
rect 222 -1014 223 -1012
rect 226 -1008 227 -1006
rect 226 -1014 227 -1012
rect 233 -1008 234 -1006
rect 233 -1014 234 -1012
rect 240 -1008 241 -1006
rect 240 -1014 241 -1012
rect 247 -1008 248 -1006
rect 247 -1014 248 -1012
rect 254 -1008 255 -1006
rect 254 -1014 255 -1012
rect 261 -1008 262 -1006
rect 261 -1014 262 -1012
rect 268 -1008 269 -1006
rect 268 -1014 269 -1012
rect 275 -1008 276 -1006
rect 275 -1014 276 -1012
rect 282 -1008 283 -1006
rect 282 -1014 283 -1012
rect 289 -1008 290 -1006
rect 289 -1014 290 -1012
rect 296 -1008 297 -1006
rect 296 -1014 297 -1012
rect 303 -1008 304 -1006
rect 303 -1014 304 -1012
rect 313 -1008 314 -1006
rect 317 -1008 318 -1006
rect 317 -1014 318 -1012
rect 324 -1008 325 -1006
rect 324 -1014 325 -1012
rect 331 -1008 332 -1006
rect 334 -1008 335 -1006
rect 331 -1014 332 -1012
rect 334 -1014 335 -1012
rect 338 -1008 339 -1006
rect 341 -1014 342 -1012
rect 345 -1008 346 -1006
rect 345 -1014 346 -1012
rect 352 -1008 353 -1006
rect 352 -1014 353 -1012
rect 359 -1008 360 -1006
rect 359 -1014 360 -1012
rect 366 -1008 367 -1006
rect 366 -1014 367 -1012
rect 373 -1008 374 -1006
rect 376 -1008 377 -1006
rect 376 -1014 377 -1012
rect 380 -1008 381 -1006
rect 380 -1014 381 -1012
rect 387 -1008 388 -1006
rect 390 -1008 391 -1006
rect 390 -1014 391 -1012
rect 394 -1008 395 -1006
rect 397 -1008 398 -1006
rect 404 -1008 405 -1006
rect 401 -1014 402 -1012
rect 404 -1014 405 -1012
rect 408 -1008 409 -1006
rect 411 -1008 412 -1006
rect 411 -1014 412 -1012
rect 415 -1008 416 -1006
rect 415 -1014 416 -1012
rect 425 -1008 426 -1006
rect 429 -1008 430 -1006
rect 429 -1014 430 -1012
rect 432 -1014 433 -1012
rect 436 -1008 437 -1006
rect 439 -1014 440 -1012
rect 443 -1008 444 -1006
rect 443 -1014 444 -1012
rect 450 -1008 451 -1006
rect 450 -1014 451 -1012
rect 457 -1008 458 -1006
rect 457 -1014 458 -1012
rect 464 -1008 465 -1006
rect 464 -1014 465 -1012
rect 474 -1008 475 -1006
rect 478 -1008 479 -1006
rect 481 -1008 482 -1006
rect 478 -1014 479 -1012
rect 485 -1008 486 -1006
rect 485 -1014 486 -1012
rect 492 -1008 493 -1006
rect 492 -1014 493 -1012
rect 499 -1008 500 -1006
rect 499 -1014 500 -1012
rect 502 -1014 503 -1012
rect 506 -1008 507 -1006
rect 506 -1014 507 -1012
rect 513 -1014 514 -1012
rect 516 -1014 517 -1012
rect 520 -1008 521 -1006
rect 520 -1014 521 -1012
rect 527 -1008 528 -1006
rect 527 -1014 528 -1012
rect 534 -1008 535 -1006
rect 534 -1014 535 -1012
rect 541 -1008 542 -1006
rect 541 -1014 542 -1012
rect 548 -1008 549 -1006
rect 548 -1014 549 -1012
rect 555 -1008 556 -1006
rect 558 -1008 559 -1006
rect 562 -1008 563 -1006
rect 562 -1014 563 -1012
rect 569 -1008 570 -1006
rect 569 -1014 570 -1012
rect 576 -1008 577 -1006
rect 576 -1014 577 -1012
rect 590 -1008 591 -1006
rect 590 -1014 591 -1012
rect 597 -1008 598 -1006
rect 597 -1014 598 -1012
rect 604 -1008 605 -1006
rect 604 -1014 605 -1012
rect 611 -1008 612 -1006
rect 611 -1014 612 -1012
rect 614 -1014 615 -1012
rect 618 -1008 619 -1006
rect 618 -1014 619 -1012
rect 625 -1008 626 -1006
rect 625 -1014 626 -1012
rect 632 -1008 633 -1006
rect 632 -1014 633 -1012
rect 639 -1008 640 -1006
rect 639 -1014 640 -1012
rect 646 -1008 647 -1006
rect 646 -1014 647 -1012
rect 653 -1008 654 -1006
rect 653 -1014 654 -1012
rect 660 -1008 661 -1006
rect 660 -1014 661 -1012
rect 667 -1008 668 -1006
rect 667 -1014 668 -1012
rect 674 -1008 675 -1006
rect 674 -1014 675 -1012
rect 681 -1008 682 -1006
rect 681 -1014 682 -1012
rect 688 -1008 689 -1006
rect 688 -1014 689 -1012
rect 695 -1008 696 -1006
rect 695 -1014 696 -1012
rect 702 -1008 703 -1006
rect 702 -1014 703 -1012
rect 709 -1008 710 -1006
rect 709 -1014 710 -1012
rect 716 -1008 717 -1006
rect 716 -1014 717 -1012
rect 723 -1008 724 -1006
rect 723 -1014 724 -1012
rect 730 -1008 731 -1006
rect 730 -1014 731 -1012
rect 737 -1008 738 -1006
rect 737 -1014 738 -1012
rect 744 -1008 745 -1006
rect 744 -1014 745 -1012
rect 751 -1008 752 -1006
rect 751 -1014 752 -1012
rect 758 -1008 759 -1006
rect 758 -1014 759 -1012
rect 765 -1008 766 -1006
rect 765 -1014 766 -1012
rect 772 -1008 773 -1006
rect 772 -1014 773 -1012
rect 779 -1008 780 -1006
rect 779 -1014 780 -1012
rect 786 -1008 787 -1006
rect 786 -1014 787 -1012
rect 793 -1008 794 -1006
rect 793 -1014 794 -1012
rect 800 -1008 801 -1006
rect 800 -1014 801 -1012
rect 807 -1008 808 -1006
rect 807 -1014 808 -1012
rect 814 -1008 815 -1006
rect 814 -1014 815 -1012
rect 821 -1008 822 -1006
rect 821 -1014 822 -1012
rect 828 -1008 829 -1006
rect 828 -1014 829 -1012
rect 835 -1008 836 -1006
rect 835 -1014 836 -1012
rect 842 -1008 843 -1006
rect 842 -1014 843 -1012
rect 849 -1008 850 -1006
rect 849 -1014 850 -1012
rect 856 -1008 857 -1006
rect 859 -1008 860 -1006
rect 859 -1014 860 -1012
rect 863 -1008 864 -1006
rect 863 -1014 864 -1012
rect 873 -1008 874 -1006
rect 898 -1008 899 -1006
rect 898 -1014 899 -1012
rect 9 -1091 10 -1089
rect 16 -1085 17 -1083
rect 16 -1091 17 -1089
rect 23 -1085 24 -1083
rect 23 -1091 24 -1089
rect 30 -1085 31 -1083
rect 30 -1091 31 -1089
rect 37 -1085 38 -1083
rect 37 -1091 38 -1089
rect 44 -1085 45 -1083
rect 44 -1091 45 -1089
rect 54 -1085 55 -1083
rect 58 -1085 59 -1083
rect 58 -1091 59 -1089
rect 65 -1085 66 -1083
rect 72 -1085 73 -1083
rect 72 -1091 73 -1089
rect 79 -1085 80 -1083
rect 79 -1091 80 -1089
rect 82 -1091 83 -1089
rect 86 -1085 87 -1083
rect 86 -1091 87 -1089
rect 93 -1091 94 -1089
rect 96 -1091 97 -1089
rect 103 -1085 104 -1083
rect 103 -1091 104 -1089
rect 107 -1085 108 -1083
rect 107 -1091 108 -1089
rect 114 -1085 115 -1083
rect 114 -1091 115 -1089
rect 121 -1085 122 -1083
rect 121 -1091 122 -1089
rect 128 -1085 129 -1083
rect 128 -1091 129 -1089
rect 135 -1091 136 -1089
rect 138 -1091 139 -1089
rect 142 -1085 143 -1083
rect 142 -1091 143 -1089
rect 152 -1085 153 -1083
rect 152 -1091 153 -1089
rect 159 -1085 160 -1083
rect 163 -1085 164 -1083
rect 166 -1085 167 -1083
rect 166 -1091 167 -1089
rect 170 -1085 171 -1083
rect 170 -1091 171 -1089
rect 177 -1085 178 -1083
rect 177 -1091 178 -1089
rect 184 -1085 185 -1083
rect 184 -1091 185 -1089
rect 191 -1085 192 -1083
rect 191 -1091 192 -1089
rect 198 -1085 199 -1083
rect 198 -1091 199 -1089
rect 205 -1085 206 -1083
rect 205 -1091 206 -1089
rect 212 -1085 213 -1083
rect 212 -1091 213 -1089
rect 222 -1085 223 -1083
rect 219 -1091 220 -1089
rect 222 -1091 223 -1089
rect 226 -1085 227 -1083
rect 226 -1091 227 -1089
rect 233 -1085 234 -1083
rect 233 -1091 234 -1089
rect 243 -1085 244 -1083
rect 250 -1091 251 -1089
rect 254 -1085 255 -1083
rect 254 -1091 255 -1089
rect 261 -1085 262 -1083
rect 261 -1091 262 -1089
rect 268 -1085 269 -1083
rect 268 -1091 269 -1089
rect 275 -1085 276 -1083
rect 278 -1085 279 -1083
rect 278 -1091 279 -1089
rect 282 -1085 283 -1083
rect 282 -1091 283 -1089
rect 289 -1085 290 -1083
rect 289 -1091 290 -1089
rect 296 -1085 297 -1083
rect 296 -1091 297 -1089
rect 303 -1085 304 -1083
rect 303 -1091 304 -1089
rect 310 -1085 311 -1083
rect 310 -1091 311 -1089
rect 317 -1085 318 -1083
rect 317 -1091 318 -1089
rect 324 -1085 325 -1083
rect 324 -1091 325 -1089
rect 331 -1085 332 -1083
rect 331 -1091 332 -1089
rect 338 -1085 339 -1083
rect 338 -1091 339 -1089
rect 345 -1085 346 -1083
rect 348 -1085 349 -1083
rect 348 -1091 349 -1089
rect 352 -1085 353 -1083
rect 355 -1091 356 -1089
rect 359 -1085 360 -1083
rect 359 -1091 360 -1089
rect 366 -1085 367 -1083
rect 366 -1091 367 -1089
rect 373 -1085 374 -1083
rect 373 -1091 374 -1089
rect 380 -1085 381 -1083
rect 380 -1091 381 -1089
rect 387 -1085 388 -1083
rect 390 -1085 391 -1083
rect 390 -1091 391 -1089
rect 394 -1085 395 -1083
rect 394 -1091 395 -1089
rect 401 -1085 402 -1083
rect 401 -1091 402 -1089
rect 408 -1085 409 -1083
rect 408 -1091 409 -1089
rect 415 -1085 416 -1083
rect 415 -1091 416 -1089
rect 422 -1085 423 -1083
rect 422 -1091 423 -1089
rect 429 -1085 430 -1083
rect 429 -1091 430 -1089
rect 436 -1085 437 -1083
rect 436 -1091 437 -1089
rect 446 -1085 447 -1083
rect 446 -1091 447 -1089
rect 450 -1085 451 -1083
rect 453 -1085 454 -1083
rect 450 -1091 451 -1089
rect 453 -1091 454 -1089
rect 457 -1085 458 -1083
rect 457 -1091 458 -1089
rect 467 -1085 468 -1083
rect 464 -1091 465 -1089
rect 471 -1085 472 -1083
rect 471 -1091 472 -1089
rect 478 -1085 479 -1083
rect 478 -1091 479 -1089
rect 485 -1085 486 -1083
rect 485 -1091 486 -1089
rect 492 -1085 493 -1083
rect 495 -1085 496 -1083
rect 492 -1091 493 -1089
rect 499 -1085 500 -1083
rect 499 -1091 500 -1089
rect 506 -1085 507 -1083
rect 506 -1091 507 -1089
rect 513 -1085 514 -1083
rect 513 -1091 514 -1089
rect 520 -1085 521 -1083
rect 520 -1091 521 -1089
rect 527 -1085 528 -1083
rect 530 -1085 531 -1083
rect 527 -1091 528 -1089
rect 530 -1091 531 -1089
rect 534 -1085 535 -1083
rect 537 -1085 538 -1083
rect 541 -1085 542 -1083
rect 541 -1091 542 -1089
rect 548 -1085 549 -1083
rect 551 -1085 552 -1083
rect 558 -1085 559 -1083
rect 558 -1091 559 -1089
rect 562 -1085 563 -1083
rect 565 -1085 566 -1083
rect 562 -1091 563 -1089
rect 572 -1085 573 -1083
rect 569 -1091 570 -1089
rect 572 -1091 573 -1089
rect 576 -1085 577 -1083
rect 576 -1091 577 -1089
rect 583 -1085 584 -1083
rect 583 -1091 584 -1089
rect 590 -1085 591 -1083
rect 590 -1091 591 -1089
rect 597 -1085 598 -1083
rect 597 -1091 598 -1089
rect 604 -1085 605 -1083
rect 607 -1085 608 -1083
rect 604 -1091 605 -1089
rect 607 -1091 608 -1089
rect 611 -1085 612 -1083
rect 614 -1085 615 -1083
rect 611 -1091 612 -1089
rect 618 -1085 619 -1083
rect 618 -1091 619 -1089
rect 625 -1085 626 -1083
rect 625 -1091 626 -1089
rect 632 -1085 633 -1083
rect 632 -1091 633 -1089
rect 642 -1085 643 -1083
rect 639 -1091 640 -1089
rect 642 -1091 643 -1089
rect 646 -1085 647 -1083
rect 646 -1091 647 -1089
rect 653 -1085 654 -1083
rect 653 -1091 654 -1089
rect 660 -1085 661 -1083
rect 660 -1091 661 -1089
rect 667 -1085 668 -1083
rect 667 -1091 668 -1089
rect 674 -1085 675 -1083
rect 674 -1091 675 -1089
rect 681 -1085 682 -1083
rect 681 -1091 682 -1089
rect 688 -1085 689 -1083
rect 688 -1091 689 -1089
rect 695 -1085 696 -1083
rect 695 -1091 696 -1089
rect 702 -1085 703 -1083
rect 702 -1091 703 -1089
rect 709 -1085 710 -1083
rect 709 -1091 710 -1089
rect 716 -1085 717 -1083
rect 716 -1091 717 -1089
rect 723 -1085 724 -1083
rect 723 -1091 724 -1089
rect 730 -1085 731 -1083
rect 730 -1091 731 -1089
rect 737 -1085 738 -1083
rect 737 -1091 738 -1089
rect 744 -1085 745 -1083
rect 744 -1091 745 -1089
rect 751 -1085 752 -1083
rect 751 -1091 752 -1089
rect 758 -1085 759 -1083
rect 758 -1091 759 -1089
rect 765 -1085 766 -1083
rect 765 -1091 766 -1089
rect 772 -1085 773 -1083
rect 772 -1091 773 -1089
rect 779 -1085 780 -1083
rect 779 -1091 780 -1089
rect 786 -1085 787 -1083
rect 786 -1091 787 -1089
rect 793 -1085 794 -1083
rect 793 -1091 794 -1089
rect 800 -1085 801 -1083
rect 800 -1091 801 -1089
rect 807 -1085 808 -1083
rect 807 -1091 808 -1089
rect 814 -1085 815 -1083
rect 814 -1091 815 -1089
rect 821 -1085 822 -1083
rect 821 -1091 822 -1089
rect 828 -1085 829 -1083
rect 828 -1091 829 -1089
rect 835 -1085 836 -1083
rect 835 -1091 836 -1089
rect 842 -1085 843 -1083
rect 842 -1091 843 -1089
rect 849 -1085 850 -1083
rect 849 -1091 850 -1089
rect 856 -1085 857 -1083
rect 856 -1091 857 -1089
rect 863 -1085 864 -1083
rect 863 -1091 864 -1089
rect 870 -1085 871 -1083
rect 870 -1091 871 -1089
rect 877 -1085 878 -1083
rect 877 -1091 878 -1089
rect 884 -1085 885 -1083
rect 884 -1091 885 -1089
rect 891 -1085 892 -1083
rect 891 -1091 892 -1089
rect 898 -1085 899 -1083
rect 898 -1091 899 -1089
rect 905 -1085 906 -1083
rect 905 -1091 906 -1089
rect 912 -1085 913 -1083
rect 912 -1091 913 -1089
rect 919 -1085 920 -1083
rect 919 -1091 920 -1089
rect 926 -1085 927 -1083
rect 926 -1091 927 -1089
rect 929 -1091 930 -1089
rect 940 -1085 941 -1083
rect 940 -1091 941 -1089
rect 5 -1188 6 -1186
rect 9 -1182 10 -1180
rect 9 -1188 10 -1186
rect 16 -1182 17 -1180
rect 16 -1188 17 -1186
rect 26 -1188 27 -1186
rect 30 -1182 31 -1180
rect 30 -1188 31 -1186
rect 37 -1182 38 -1180
rect 37 -1188 38 -1186
rect 44 -1182 45 -1180
rect 44 -1188 45 -1186
rect 51 -1182 52 -1180
rect 51 -1188 52 -1186
rect 58 -1182 59 -1180
rect 58 -1188 59 -1186
rect 65 -1182 66 -1180
rect 65 -1188 66 -1186
rect 72 -1182 73 -1180
rect 79 -1182 80 -1180
rect 79 -1188 80 -1186
rect 86 -1182 87 -1180
rect 86 -1188 87 -1186
rect 93 -1182 94 -1180
rect 93 -1188 94 -1186
rect 96 -1188 97 -1186
rect 103 -1182 104 -1180
rect 103 -1188 104 -1186
rect 107 -1182 108 -1180
rect 107 -1188 108 -1186
rect 114 -1182 115 -1180
rect 114 -1188 115 -1186
rect 121 -1188 122 -1186
rect 124 -1188 125 -1186
rect 128 -1182 129 -1180
rect 128 -1188 129 -1186
rect 135 -1182 136 -1180
rect 135 -1188 136 -1186
rect 142 -1182 143 -1180
rect 142 -1188 143 -1186
rect 152 -1182 153 -1180
rect 149 -1188 150 -1186
rect 152 -1188 153 -1186
rect 156 -1182 157 -1180
rect 156 -1188 157 -1186
rect 163 -1182 164 -1180
rect 163 -1188 164 -1186
rect 170 -1182 171 -1180
rect 173 -1188 174 -1186
rect 177 -1182 178 -1180
rect 177 -1188 178 -1186
rect 184 -1182 185 -1180
rect 184 -1188 185 -1186
rect 191 -1182 192 -1180
rect 191 -1188 192 -1186
rect 198 -1182 199 -1180
rect 201 -1182 202 -1180
rect 198 -1188 199 -1186
rect 201 -1188 202 -1186
rect 205 -1182 206 -1180
rect 205 -1188 206 -1186
rect 212 -1182 213 -1180
rect 212 -1188 213 -1186
rect 215 -1188 216 -1186
rect 222 -1182 223 -1180
rect 219 -1188 220 -1186
rect 222 -1188 223 -1186
rect 226 -1182 227 -1180
rect 226 -1188 227 -1186
rect 233 -1182 234 -1180
rect 233 -1188 234 -1186
rect 240 -1182 241 -1180
rect 240 -1188 241 -1186
rect 247 -1182 248 -1180
rect 247 -1188 248 -1186
rect 254 -1182 255 -1180
rect 254 -1188 255 -1186
rect 261 -1182 262 -1180
rect 261 -1188 262 -1186
rect 268 -1182 269 -1180
rect 268 -1188 269 -1186
rect 275 -1182 276 -1180
rect 275 -1188 276 -1186
rect 282 -1182 283 -1180
rect 282 -1188 283 -1186
rect 285 -1188 286 -1186
rect 289 -1182 290 -1180
rect 289 -1188 290 -1186
rect 296 -1182 297 -1180
rect 296 -1188 297 -1186
rect 303 -1182 304 -1180
rect 303 -1188 304 -1186
rect 310 -1182 311 -1180
rect 310 -1188 311 -1186
rect 320 -1182 321 -1180
rect 320 -1188 321 -1186
rect 324 -1182 325 -1180
rect 324 -1188 325 -1186
rect 331 -1182 332 -1180
rect 331 -1188 332 -1186
rect 338 -1182 339 -1180
rect 338 -1188 339 -1186
rect 345 -1182 346 -1180
rect 345 -1188 346 -1186
rect 355 -1182 356 -1180
rect 355 -1188 356 -1186
rect 359 -1182 360 -1180
rect 362 -1182 363 -1180
rect 366 -1182 367 -1180
rect 366 -1188 367 -1186
rect 373 -1182 374 -1180
rect 373 -1188 374 -1186
rect 380 -1182 381 -1180
rect 380 -1188 381 -1186
rect 387 -1182 388 -1180
rect 387 -1188 388 -1186
rect 394 -1182 395 -1180
rect 394 -1188 395 -1186
rect 401 -1182 402 -1180
rect 401 -1188 402 -1186
rect 408 -1188 409 -1186
rect 411 -1188 412 -1186
rect 415 -1182 416 -1180
rect 415 -1188 416 -1186
rect 422 -1182 423 -1180
rect 425 -1182 426 -1180
rect 425 -1188 426 -1186
rect 429 -1182 430 -1180
rect 429 -1188 430 -1186
rect 436 -1182 437 -1180
rect 436 -1188 437 -1186
rect 443 -1182 444 -1180
rect 443 -1188 444 -1186
rect 450 -1182 451 -1180
rect 453 -1182 454 -1180
rect 450 -1188 451 -1186
rect 453 -1188 454 -1186
rect 457 -1182 458 -1180
rect 457 -1188 458 -1186
rect 464 -1188 465 -1186
rect 467 -1188 468 -1186
rect 471 -1182 472 -1180
rect 471 -1188 472 -1186
rect 478 -1182 479 -1180
rect 478 -1188 479 -1186
rect 485 -1182 486 -1180
rect 485 -1188 486 -1186
rect 492 -1182 493 -1180
rect 492 -1188 493 -1186
rect 499 -1182 500 -1180
rect 499 -1188 500 -1186
rect 506 -1182 507 -1180
rect 509 -1182 510 -1180
rect 506 -1188 507 -1186
rect 513 -1182 514 -1180
rect 513 -1188 514 -1186
rect 520 -1182 521 -1180
rect 520 -1188 521 -1186
rect 527 -1182 528 -1180
rect 527 -1188 528 -1186
rect 534 -1182 535 -1180
rect 534 -1188 535 -1186
rect 541 -1182 542 -1180
rect 544 -1182 545 -1180
rect 541 -1188 542 -1186
rect 544 -1188 545 -1186
rect 548 -1182 549 -1180
rect 548 -1188 549 -1186
rect 555 -1182 556 -1180
rect 555 -1188 556 -1186
rect 562 -1182 563 -1180
rect 562 -1188 563 -1186
rect 569 -1182 570 -1180
rect 569 -1188 570 -1186
rect 579 -1182 580 -1180
rect 579 -1188 580 -1186
rect 583 -1182 584 -1180
rect 583 -1188 584 -1186
rect 590 -1182 591 -1180
rect 590 -1188 591 -1186
rect 597 -1182 598 -1180
rect 597 -1188 598 -1186
rect 604 -1182 605 -1180
rect 604 -1188 605 -1186
rect 611 -1182 612 -1180
rect 611 -1188 612 -1186
rect 618 -1182 619 -1180
rect 625 -1182 626 -1180
rect 625 -1188 626 -1186
rect 632 -1182 633 -1180
rect 632 -1188 633 -1186
rect 639 -1182 640 -1180
rect 639 -1188 640 -1186
rect 646 -1182 647 -1180
rect 646 -1188 647 -1186
rect 656 -1182 657 -1180
rect 656 -1188 657 -1186
rect 660 -1182 661 -1180
rect 660 -1188 661 -1186
rect 667 -1182 668 -1180
rect 667 -1188 668 -1186
rect 674 -1182 675 -1180
rect 674 -1188 675 -1186
rect 681 -1182 682 -1180
rect 684 -1182 685 -1180
rect 688 -1182 689 -1180
rect 688 -1188 689 -1186
rect 695 -1182 696 -1180
rect 695 -1188 696 -1186
rect 702 -1182 703 -1180
rect 702 -1188 703 -1186
rect 709 -1182 710 -1180
rect 709 -1188 710 -1186
rect 716 -1182 717 -1180
rect 719 -1188 720 -1186
rect 723 -1182 724 -1180
rect 723 -1188 724 -1186
rect 730 -1182 731 -1180
rect 730 -1188 731 -1186
rect 737 -1182 738 -1180
rect 737 -1188 738 -1186
rect 744 -1182 745 -1180
rect 744 -1188 745 -1186
rect 751 -1182 752 -1180
rect 751 -1188 752 -1186
rect 758 -1182 759 -1180
rect 758 -1188 759 -1186
rect 765 -1182 766 -1180
rect 765 -1188 766 -1186
rect 772 -1182 773 -1180
rect 772 -1188 773 -1186
rect 779 -1182 780 -1180
rect 779 -1188 780 -1186
rect 786 -1182 787 -1180
rect 786 -1188 787 -1186
rect 793 -1182 794 -1180
rect 793 -1188 794 -1186
rect 800 -1182 801 -1180
rect 800 -1188 801 -1186
rect 807 -1182 808 -1180
rect 807 -1188 808 -1186
rect 814 -1182 815 -1180
rect 814 -1188 815 -1186
rect 821 -1182 822 -1180
rect 821 -1188 822 -1186
rect 828 -1182 829 -1180
rect 828 -1188 829 -1186
rect 835 -1182 836 -1180
rect 835 -1188 836 -1186
rect 842 -1182 843 -1180
rect 842 -1188 843 -1186
rect 849 -1182 850 -1180
rect 849 -1188 850 -1186
rect 856 -1182 857 -1180
rect 856 -1188 857 -1186
rect 863 -1182 864 -1180
rect 863 -1188 864 -1186
rect 870 -1182 871 -1180
rect 870 -1188 871 -1186
rect 877 -1182 878 -1180
rect 877 -1188 878 -1186
rect 884 -1182 885 -1180
rect 884 -1188 885 -1186
rect 891 -1182 892 -1180
rect 891 -1188 892 -1186
rect 898 -1182 899 -1180
rect 898 -1188 899 -1186
rect 905 -1182 906 -1180
rect 905 -1188 906 -1186
rect 912 -1182 913 -1180
rect 912 -1188 913 -1186
rect 919 -1182 920 -1180
rect 919 -1188 920 -1186
rect 926 -1182 927 -1180
rect 926 -1188 927 -1186
rect 933 -1182 934 -1180
rect 933 -1188 934 -1186
rect 940 -1182 941 -1180
rect 940 -1188 941 -1186
rect 947 -1182 948 -1180
rect 947 -1188 948 -1186
rect 957 -1188 958 -1186
rect 961 -1182 962 -1180
rect 961 -1188 962 -1186
rect 964 -1188 965 -1186
rect 968 -1182 969 -1180
rect 968 -1188 969 -1186
rect 975 -1182 976 -1180
rect 975 -1188 976 -1186
rect 982 -1182 983 -1180
rect 985 -1188 986 -1186
rect 989 -1182 990 -1180
rect 989 -1188 990 -1186
rect 12 -1277 13 -1275
rect 16 -1277 17 -1275
rect 16 -1283 17 -1281
rect 26 -1277 27 -1275
rect 30 -1277 31 -1275
rect 30 -1283 31 -1281
rect 40 -1277 41 -1275
rect 44 -1277 45 -1275
rect 44 -1283 45 -1281
rect 51 -1277 52 -1275
rect 51 -1283 52 -1281
rect 58 -1277 59 -1275
rect 58 -1283 59 -1281
rect 65 -1277 66 -1275
rect 65 -1283 66 -1281
rect 72 -1277 73 -1275
rect 72 -1283 73 -1281
rect 79 -1277 80 -1275
rect 79 -1283 80 -1281
rect 86 -1277 87 -1275
rect 86 -1283 87 -1281
rect 93 -1277 94 -1275
rect 96 -1277 97 -1275
rect 96 -1283 97 -1281
rect 100 -1277 101 -1275
rect 100 -1283 101 -1281
rect 110 -1277 111 -1275
rect 110 -1283 111 -1281
rect 114 -1277 115 -1275
rect 114 -1283 115 -1281
rect 121 -1277 122 -1275
rect 121 -1283 122 -1281
rect 128 -1277 129 -1275
rect 128 -1283 129 -1281
rect 135 -1277 136 -1275
rect 135 -1283 136 -1281
rect 142 -1277 143 -1275
rect 142 -1283 143 -1281
rect 149 -1277 150 -1275
rect 149 -1283 150 -1281
rect 156 -1277 157 -1275
rect 156 -1283 157 -1281
rect 163 -1277 164 -1275
rect 163 -1283 164 -1281
rect 170 -1277 171 -1275
rect 173 -1283 174 -1281
rect 177 -1277 178 -1275
rect 177 -1283 178 -1281
rect 184 -1277 185 -1275
rect 184 -1283 185 -1281
rect 191 -1277 192 -1275
rect 191 -1283 192 -1281
rect 198 -1277 199 -1275
rect 198 -1283 199 -1281
rect 205 -1277 206 -1275
rect 205 -1283 206 -1281
rect 212 -1277 213 -1275
rect 215 -1277 216 -1275
rect 222 -1277 223 -1275
rect 219 -1283 220 -1281
rect 222 -1283 223 -1281
rect 226 -1277 227 -1275
rect 226 -1283 227 -1281
rect 233 -1277 234 -1275
rect 233 -1283 234 -1281
rect 240 -1277 241 -1275
rect 240 -1283 241 -1281
rect 247 -1277 248 -1275
rect 247 -1283 248 -1281
rect 254 -1277 255 -1275
rect 254 -1283 255 -1281
rect 261 -1277 262 -1275
rect 261 -1283 262 -1281
rect 268 -1277 269 -1275
rect 268 -1283 269 -1281
rect 275 -1277 276 -1275
rect 275 -1283 276 -1281
rect 282 -1277 283 -1275
rect 282 -1283 283 -1281
rect 289 -1277 290 -1275
rect 289 -1283 290 -1281
rect 296 -1277 297 -1275
rect 296 -1283 297 -1281
rect 303 -1277 304 -1275
rect 306 -1277 307 -1275
rect 303 -1283 304 -1281
rect 310 -1277 311 -1275
rect 313 -1277 314 -1275
rect 310 -1283 311 -1281
rect 313 -1283 314 -1281
rect 317 -1277 318 -1275
rect 317 -1283 318 -1281
rect 324 -1277 325 -1275
rect 324 -1283 325 -1281
rect 331 -1277 332 -1275
rect 331 -1283 332 -1281
rect 341 -1277 342 -1275
rect 338 -1283 339 -1281
rect 341 -1283 342 -1281
rect 345 -1277 346 -1275
rect 345 -1283 346 -1281
rect 352 -1277 353 -1275
rect 352 -1283 353 -1281
rect 359 -1277 360 -1275
rect 362 -1277 363 -1275
rect 359 -1283 360 -1281
rect 366 -1277 367 -1275
rect 366 -1283 367 -1281
rect 373 -1277 374 -1275
rect 373 -1283 374 -1281
rect 380 -1277 381 -1275
rect 380 -1283 381 -1281
rect 383 -1283 384 -1281
rect 387 -1277 388 -1275
rect 387 -1283 388 -1281
rect 394 -1277 395 -1275
rect 394 -1283 395 -1281
rect 401 -1277 402 -1275
rect 401 -1283 402 -1281
rect 408 -1277 409 -1275
rect 411 -1277 412 -1275
rect 408 -1283 409 -1281
rect 411 -1283 412 -1281
rect 415 -1277 416 -1275
rect 415 -1283 416 -1281
rect 422 -1277 423 -1275
rect 422 -1283 423 -1281
rect 429 -1277 430 -1275
rect 429 -1283 430 -1281
rect 436 -1277 437 -1275
rect 436 -1283 437 -1281
rect 443 -1277 444 -1275
rect 446 -1277 447 -1275
rect 443 -1283 444 -1281
rect 446 -1283 447 -1281
rect 450 -1277 451 -1275
rect 450 -1283 451 -1281
rect 457 -1277 458 -1275
rect 460 -1277 461 -1275
rect 460 -1283 461 -1281
rect 464 -1277 465 -1275
rect 467 -1277 468 -1275
rect 464 -1283 465 -1281
rect 471 -1277 472 -1275
rect 474 -1277 475 -1275
rect 471 -1283 472 -1281
rect 474 -1283 475 -1281
rect 478 -1277 479 -1275
rect 478 -1283 479 -1281
rect 485 -1277 486 -1275
rect 485 -1283 486 -1281
rect 492 -1277 493 -1275
rect 495 -1277 496 -1275
rect 499 -1283 500 -1281
rect 502 -1283 503 -1281
rect 506 -1283 507 -1281
rect 509 -1283 510 -1281
rect 513 -1277 514 -1275
rect 513 -1283 514 -1281
rect 520 -1277 521 -1275
rect 520 -1283 521 -1281
rect 527 -1277 528 -1275
rect 527 -1283 528 -1281
rect 534 -1277 535 -1275
rect 534 -1283 535 -1281
rect 541 -1277 542 -1275
rect 541 -1283 542 -1281
rect 548 -1277 549 -1275
rect 548 -1283 549 -1281
rect 555 -1277 556 -1275
rect 555 -1283 556 -1281
rect 562 -1277 563 -1275
rect 562 -1283 563 -1281
rect 569 -1277 570 -1275
rect 569 -1283 570 -1281
rect 576 -1277 577 -1275
rect 576 -1283 577 -1281
rect 583 -1277 584 -1275
rect 583 -1283 584 -1281
rect 590 -1277 591 -1275
rect 590 -1283 591 -1281
rect 597 -1277 598 -1275
rect 600 -1277 601 -1275
rect 604 -1277 605 -1275
rect 607 -1277 608 -1275
rect 604 -1283 605 -1281
rect 611 -1277 612 -1275
rect 611 -1283 612 -1281
rect 618 -1277 619 -1275
rect 618 -1283 619 -1281
rect 625 -1277 626 -1275
rect 625 -1283 626 -1281
rect 635 -1277 636 -1275
rect 639 -1277 640 -1275
rect 639 -1283 640 -1281
rect 646 -1277 647 -1275
rect 646 -1283 647 -1281
rect 653 -1277 654 -1275
rect 656 -1277 657 -1275
rect 653 -1283 654 -1281
rect 656 -1283 657 -1281
rect 660 -1277 661 -1275
rect 660 -1283 661 -1281
rect 670 -1277 671 -1275
rect 667 -1283 668 -1281
rect 674 -1277 675 -1275
rect 674 -1283 675 -1281
rect 681 -1277 682 -1275
rect 681 -1283 682 -1281
rect 688 -1277 689 -1275
rect 688 -1283 689 -1281
rect 695 -1277 696 -1275
rect 695 -1283 696 -1281
rect 702 -1277 703 -1275
rect 702 -1283 703 -1281
rect 709 -1277 710 -1275
rect 709 -1283 710 -1281
rect 716 -1277 717 -1275
rect 716 -1283 717 -1281
rect 723 -1277 724 -1275
rect 723 -1283 724 -1281
rect 730 -1277 731 -1275
rect 730 -1283 731 -1281
rect 737 -1277 738 -1275
rect 737 -1283 738 -1281
rect 744 -1277 745 -1275
rect 744 -1283 745 -1281
rect 751 -1277 752 -1275
rect 751 -1283 752 -1281
rect 758 -1277 759 -1275
rect 758 -1283 759 -1281
rect 765 -1277 766 -1275
rect 765 -1283 766 -1281
rect 772 -1277 773 -1275
rect 772 -1283 773 -1281
rect 779 -1277 780 -1275
rect 779 -1283 780 -1281
rect 786 -1277 787 -1275
rect 786 -1283 787 -1281
rect 793 -1277 794 -1275
rect 793 -1283 794 -1281
rect 800 -1277 801 -1275
rect 800 -1283 801 -1281
rect 807 -1277 808 -1275
rect 807 -1283 808 -1281
rect 814 -1277 815 -1275
rect 814 -1283 815 -1281
rect 821 -1277 822 -1275
rect 821 -1283 822 -1281
rect 828 -1277 829 -1275
rect 828 -1283 829 -1281
rect 835 -1277 836 -1275
rect 835 -1283 836 -1281
rect 842 -1277 843 -1275
rect 842 -1283 843 -1281
rect 849 -1277 850 -1275
rect 849 -1283 850 -1281
rect 856 -1277 857 -1275
rect 856 -1283 857 -1281
rect 863 -1277 864 -1275
rect 863 -1283 864 -1281
rect 870 -1277 871 -1275
rect 870 -1283 871 -1281
rect 877 -1277 878 -1275
rect 877 -1283 878 -1281
rect 884 -1277 885 -1275
rect 884 -1283 885 -1281
rect 891 -1277 892 -1275
rect 891 -1283 892 -1281
rect 898 -1277 899 -1275
rect 898 -1283 899 -1281
rect 905 -1277 906 -1275
rect 905 -1283 906 -1281
rect 912 -1277 913 -1275
rect 912 -1283 913 -1281
rect 919 -1277 920 -1275
rect 919 -1283 920 -1281
rect 926 -1277 927 -1275
rect 926 -1283 927 -1281
rect 933 -1277 934 -1275
rect 933 -1283 934 -1281
rect 943 -1277 944 -1275
rect 943 -1283 944 -1281
rect 947 -1277 948 -1275
rect 947 -1283 948 -1281
rect 954 -1277 955 -1275
rect 954 -1283 955 -1281
rect 961 -1277 962 -1275
rect 961 -1283 962 -1281
rect 968 -1277 969 -1275
rect 968 -1283 969 -1281
rect 975 -1277 976 -1275
rect 975 -1283 976 -1281
rect 982 -1277 983 -1275
rect 982 -1283 983 -1281
rect 989 -1277 990 -1275
rect 989 -1283 990 -1281
rect 996 -1277 997 -1275
rect 996 -1283 997 -1281
rect 1003 -1277 1004 -1275
rect 1003 -1283 1004 -1281
rect 1010 -1277 1011 -1275
rect 1010 -1283 1011 -1281
rect 9 -1362 10 -1360
rect 12 -1362 13 -1360
rect 9 -1368 10 -1366
rect 16 -1362 17 -1360
rect 16 -1368 17 -1366
rect 23 -1368 24 -1366
rect 30 -1362 31 -1360
rect 33 -1368 34 -1366
rect 37 -1362 38 -1360
rect 37 -1368 38 -1366
rect 44 -1362 45 -1360
rect 44 -1368 45 -1366
rect 51 -1362 52 -1360
rect 51 -1368 52 -1366
rect 61 -1362 62 -1360
rect 65 -1362 66 -1360
rect 65 -1368 66 -1366
rect 72 -1362 73 -1360
rect 72 -1368 73 -1366
rect 79 -1362 80 -1360
rect 79 -1368 80 -1366
rect 89 -1362 90 -1360
rect 89 -1368 90 -1366
rect 93 -1362 94 -1360
rect 93 -1368 94 -1366
rect 100 -1362 101 -1360
rect 100 -1368 101 -1366
rect 107 -1362 108 -1360
rect 107 -1368 108 -1366
rect 114 -1362 115 -1360
rect 114 -1368 115 -1366
rect 121 -1362 122 -1360
rect 124 -1362 125 -1360
rect 121 -1368 122 -1366
rect 128 -1362 129 -1360
rect 128 -1368 129 -1366
rect 135 -1362 136 -1360
rect 135 -1368 136 -1366
rect 142 -1362 143 -1360
rect 142 -1368 143 -1366
rect 149 -1362 150 -1360
rect 149 -1368 150 -1366
rect 156 -1362 157 -1360
rect 156 -1368 157 -1366
rect 159 -1368 160 -1366
rect 163 -1362 164 -1360
rect 163 -1368 164 -1366
rect 170 -1362 171 -1360
rect 170 -1368 171 -1366
rect 177 -1362 178 -1360
rect 177 -1368 178 -1366
rect 184 -1362 185 -1360
rect 184 -1368 185 -1366
rect 191 -1362 192 -1360
rect 191 -1368 192 -1366
rect 194 -1368 195 -1366
rect 198 -1362 199 -1360
rect 198 -1368 199 -1366
rect 208 -1362 209 -1360
rect 205 -1368 206 -1366
rect 212 -1362 213 -1360
rect 215 -1362 216 -1360
rect 219 -1362 220 -1360
rect 219 -1368 220 -1366
rect 222 -1368 223 -1366
rect 226 -1362 227 -1360
rect 229 -1362 230 -1360
rect 229 -1368 230 -1366
rect 233 -1362 234 -1360
rect 233 -1368 234 -1366
rect 240 -1362 241 -1360
rect 240 -1368 241 -1366
rect 247 -1362 248 -1360
rect 247 -1368 248 -1366
rect 254 -1362 255 -1360
rect 254 -1368 255 -1366
rect 261 -1362 262 -1360
rect 261 -1368 262 -1366
rect 268 -1362 269 -1360
rect 268 -1368 269 -1366
rect 275 -1362 276 -1360
rect 275 -1368 276 -1366
rect 282 -1362 283 -1360
rect 282 -1368 283 -1366
rect 289 -1362 290 -1360
rect 289 -1368 290 -1366
rect 296 -1362 297 -1360
rect 296 -1368 297 -1366
rect 303 -1362 304 -1360
rect 303 -1368 304 -1366
rect 310 -1362 311 -1360
rect 310 -1368 311 -1366
rect 317 -1362 318 -1360
rect 317 -1368 318 -1366
rect 324 -1362 325 -1360
rect 324 -1368 325 -1366
rect 331 -1362 332 -1360
rect 331 -1368 332 -1366
rect 334 -1368 335 -1366
rect 338 -1362 339 -1360
rect 338 -1368 339 -1366
rect 345 -1368 346 -1366
rect 348 -1368 349 -1366
rect 352 -1362 353 -1360
rect 352 -1368 353 -1366
rect 359 -1362 360 -1360
rect 359 -1368 360 -1366
rect 366 -1362 367 -1360
rect 366 -1368 367 -1366
rect 373 -1362 374 -1360
rect 373 -1368 374 -1366
rect 376 -1368 377 -1366
rect 383 -1362 384 -1360
rect 380 -1368 381 -1366
rect 387 -1362 388 -1360
rect 387 -1368 388 -1366
rect 394 -1362 395 -1360
rect 394 -1368 395 -1366
rect 397 -1368 398 -1366
rect 401 -1362 402 -1360
rect 401 -1368 402 -1366
rect 408 -1362 409 -1360
rect 408 -1368 409 -1366
rect 415 -1362 416 -1360
rect 415 -1368 416 -1366
rect 422 -1362 423 -1360
rect 422 -1368 423 -1366
rect 429 -1362 430 -1360
rect 432 -1362 433 -1360
rect 432 -1368 433 -1366
rect 436 -1362 437 -1360
rect 436 -1368 437 -1366
rect 443 -1362 444 -1360
rect 443 -1368 444 -1366
rect 450 -1362 451 -1360
rect 453 -1362 454 -1360
rect 457 -1362 458 -1360
rect 457 -1368 458 -1366
rect 464 -1362 465 -1360
rect 467 -1362 468 -1360
rect 464 -1368 465 -1366
rect 467 -1368 468 -1366
rect 471 -1362 472 -1360
rect 471 -1368 472 -1366
rect 478 -1362 479 -1360
rect 481 -1362 482 -1360
rect 478 -1368 479 -1366
rect 481 -1368 482 -1366
rect 485 -1362 486 -1360
rect 488 -1362 489 -1360
rect 485 -1368 486 -1366
rect 492 -1362 493 -1360
rect 492 -1368 493 -1366
rect 499 -1362 500 -1360
rect 499 -1368 500 -1366
rect 506 -1362 507 -1360
rect 506 -1368 507 -1366
rect 513 -1362 514 -1360
rect 513 -1368 514 -1366
rect 516 -1368 517 -1366
rect 520 -1362 521 -1360
rect 520 -1368 521 -1366
rect 527 -1362 528 -1360
rect 530 -1362 531 -1360
rect 527 -1368 528 -1366
rect 530 -1368 531 -1366
rect 534 -1362 535 -1360
rect 534 -1368 535 -1366
rect 541 -1362 542 -1360
rect 541 -1368 542 -1366
rect 548 -1362 549 -1360
rect 548 -1368 549 -1366
rect 555 -1362 556 -1360
rect 555 -1368 556 -1366
rect 562 -1362 563 -1360
rect 562 -1368 563 -1366
rect 569 -1362 570 -1360
rect 569 -1368 570 -1366
rect 576 -1362 577 -1360
rect 579 -1362 580 -1360
rect 579 -1368 580 -1366
rect 583 -1362 584 -1360
rect 583 -1368 584 -1366
rect 590 -1362 591 -1360
rect 590 -1368 591 -1366
rect 597 -1362 598 -1360
rect 597 -1368 598 -1366
rect 604 -1362 605 -1360
rect 604 -1368 605 -1366
rect 611 -1362 612 -1360
rect 611 -1368 612 -1366
rect 618 -1362 619 -1360
rect 618 -1368 619 -1366
rect 625 -1362 626 -1360
rect 625 -1368 626 -1366
rect 632 -1362 633 -1360
rect 632 -1368 633 -1366
rect 639 -1362 640 -1360
rect 639 -1368 640 -1366
rect 646 -1362 647 -1360
rect 646 -1368 647 -1366
rect 653 -1362 654 -1360
rect 653 -1368 654 -1366
rect 660 -1362 661 -1360
rect 660 -1368 661 -1366
rect 667 -1362 668 -1360
rect 667 -1368 668 -1366
rect 674 -1362 675 -1360
rect 674 -1368 675 -1366
rect 681 -1362 682 -1360
rect 681 -1368 682 -1366
rect 688 -1362 689 -1360
rect 688 -1368 689 -1366
rect 695 -1362 696 -1360
rect 695 -1368 696 -1366
rect 702 -1362 703 -1360
rect 702 -1368 703 -1366
rect 709 -1362 710 -1360
rect 709 -1368 710 -1366
rect 716 -1362 717 -1360
rect 716 -1368 717 -1366
rect 723 -1362 724 -1360
rect 723 -1368 724 -1366
rect 730 -1362 731 -1360
rect 730 -1368 731 -1366
rect 737 -1362 738 -1360
rect 737 -1368 738 -1366
rect 744 -1362 745 -1360
rect 744 -1368 745 -1366
rect 751 -1362 752 -1360
rect 751 -1368 752 -1366
rect 758 -1362 759 -1360
rect 758 -1368 759 -1366
rect 765 -1362 766 -1360
rect 765 -1368 766 -1366
rect 772 -1362 773 -1360
rect 772 -1368 773 -1366
rect 779 -1362 780 -1360
rect 779 -1368 780 -1366
rect 786 -1362 787 -1360
rect 786 -1368 787 -1366
rect 793 -1362 794 -1360
rect 793 -1368 794 -1366
rect 800 -1362 801 -1360
rect 800 -1368 801 -1366
rect 807 -1362 808 -1360
rect 807 -1368 808 -1366
rect 814 -1362 815 -1360
rect 814 -1368 815 -1366
rect 821 -1362 822 -1360
rect 821 -1368 822 -1366
rect 828 -1362 829 -1360
rect 828 -1368 829 -1366
rect 835 -1362 836 -1360
rect 835 -1368 836 -1366
rect 842 -1362 843 -1360
rect 842 -1368 843 -1366
rect 849 -1362 850 -1360
rect 849 -1368 850 -1366
rect 856 -1362 857 -1360
rect 856 -1368 857 -1366
rect 863 -1362 864 -1360
rect 863 -1368 864 -1366
rect 870 -1362 871 -1360
rect 870 -1368 871 -1366
rect 877 -1362 878 -1360
rect 877 -1368 878 -1366
rect 884 -1362 885 -1360
rect 884 -1368 885 -1366
rect 891 -1362 892 -1360
rect 891 -1368 892 -1366
rect 898 -1362 899 -1360
rect 898 -1368 899 -1366
rect 905 -1362 906 -1360
rect 908 -1368 909 -1366
rect 912 -1362 913 -1360
rect 912 -1368 913 -1366
rect 919 -1362 920 -1360
rect 940 -1362 941 -1360
rect 943 -1362 944 -1360
rect 943 -1368 944 -1366
rect 954 -1362 955 -1360
rect 954 -1368 955 -1366
rect 971 -1362 972 -1360
rect 971 -1368 972 -1366
rect 989 -1362 990 -1360
rect 989 -1368 990 -1366
rect 2 -1441 3 -1439
rect 2 -1447 3 -1445
rect 9 -1441 10 -1439
rect 16 -1441 17 -1439
rect 16 -1447 17 -1445
rect 23 -1441 24 -1439
rect 23 -1447 24 -1445
rect 30 -1441 31 -1439
rect 30 -1447 31 -1445
rect 37 -1441 38 -1439
rect 37 -1447 38 -1445
rect 51 -1441 52 -1439
rect 51 -1447 52 -1445
rect 58 -1441 59 -1439
rect 58 -1447 59 -1445
rect 65 -1441 66 -1439
rect 65 -1447 66 -1445
rect 72 -1441 73 -1439
rect 72 -1447 73 -1445
rect 79 -1441 80 -1439
rect 79 -1447 80 -1445
rect 86 -1441 87 -1439
rect 86 -1447 87 -1445
rect 93 -1441 94 -1439
rect 93 -1447 94 -1445
rect 100 -1441 101 -1439
rect 100 -1447 101 -1445
rect 107 -1441 108 -1439
rect 107 -1447 108 -1445
rect 117 -1441 118 -1439
rect 117 -1447 118 -1445
rect 121 -1441 122 -1439
rect 124 -1441 125 -1439
rect 128 -1441 129 -1439
rect 131 -1447 132 -1445
rect 135 -1441 136 -1439
rect 135 -1447 136 -1445
rect 142 -1447 143 -1445
rect 149 -1441 150 -1439
rect 149 -1447 150 -1445
rect 159 -1441 160 -1439
rect 156 -1447 157 -1445
rect 166 -1441 167 -1439
rect 163 -1447 164 -1445
rect 170 -1441 171 -1439
rect 170 -1447 171 -1445
rect 177 -1441 178 -1439
rect 177 -1447 178 -1445
rect 187 -1441 188 -1439
rect 184 -1447 185 -1445
rect 187 -1447 188 -1445
rect 191 -1441 192 -1439
rect 191 -1447 192 -1445
rect 198 -1441 199 -1439
rect 198 -1447 199 -1445
rect 205 -1441 206 -1439
rect 205 -1447 206 -1445
rect 212 -1441 213 -1439
rect 219 -1441 220 -1439
rect 219 -1447 220 -1445
rect 226 -1441 227 -1439
rect 226 -1447 227 -1445
rect 233 -1441 234 -1439
rect 233 -1447 234 -1445
rect 240 -1441 241 -1439
rect 240 -1447 241 -1445
rect 247 -1441 248 -1439
rect 247 -1447 248 -1445
rect 254 -1441 255 -1439
rect 254 -1447 255 -1445
rect 261 -1441 262 -1439
rect 261 -1447 262 -1445
rect 268 -1441 269 -1439
rect 268 -1447 269 -1445
rect 275 -1441 276 -1439
rect 275 -1447 276 -1445
rect 282 -1441 283 -1439
rect 282 -1447 283 -1445
rect 289 -1441 290 -1439
rect 289 -1447 290 -1445
rect 296 -1441 297 -1439
rect 296 -1447 297 -1445
rect 303 -1441 304 -1439
rect 303 -1447 304 -1445
rect 310 -1441 311 -1439
rect 310 -1447 311 -1445
rect 317 -1441 318 -1439
rect 317 -1447 318 -1445
rect 324 -1447 325 -1445
rect 331 -1441 332 -1439
rect 331 -1447 332 -1445
rect 338 -1441 339 -1439
rect 345 -1441 346 -1439
rect 345 -1447 346 -1445
rect 352 -1441 353 -1439
rect 352 -1447 353 -1445
rect 355 -1447 356 -1445
rect 359 -1441 360 -1439
rect 359 -1447 360 -1445
rect 366 -1441 367 -1439
rect 366 -1447 367 -1445
rect 373 -1441 374 -1439
rect 376 -1441 377 -1439
rect 376 -1447 377 -1445
rect 380 -1441 381 -1439
rect 380 -1447 381 -1445
rect 390 -1441 391 -1439
rect 390 -1447 391 -1445
rect 394 -1447 395 -1445
rect 397 -1447 398 -1445
rect 401 -1441 402 -1439
rect 401 -1447 402 -1445
rect 408 -1441 409 -1439
rect 408 -1447 409 -1445
rect 415 -1441 416 -1439
rect 415 -1447 416 -1445
rect 422 -1441 423 -1439
rect 422 -1447 423 -1445
rect 429 -1447 430 -1445
rect 432 -1447 433 -1445
rect 436 -1441 437 -1439
rect 436 -1447 437 -1445
rect 443 -1441 444 -1439
rect 443 -1447 444 -1445
rect 450 -1441 451 -1439
rect 453 -1441 454 -1439
rect 460 -1441 461 -1439
rect 460 -1447 461 -1445
rect 464 -1441 465 -1439
rect 467 -1441 468 -1439
rect 464 -1447 465 -1445
rect 467 -1447 468 -1445
rect 471 -1441 472 -1439
rect 471 -1447 472 -1445
rect 478 -1441 479 -1439
rect 478 -1447 479 -1445
rect 488 -1441 489 -1439
rect 485 -1447 486 -1445
rect 492 -1441 493 -1439
rect 492 -1447 493 -1445
rect 499 -1441 500 -1439
rect 499 -1447 500 -1445
rect 506 -1441 507 -1439
rect 509 -1441 510 -1439
rect 506 -1447 507 -1445
rect 509 -1447 510 -1445
rect 513 -1441 514 -1439
rect 513 -1447 514 -1445
rect 520 -1441 521 -1439
rect 520 -1447 521 -1445
rect 527 -1441 528 -1439
rect 527 -1447 528 -1445
rect 537 -1441 538 -1439
rect 537 -1447 538 -1445
rect 541 -1441 542 -1439
rect 541 -1447 542 -1445
rect 551 -1441 552 -1439
rect 548 -1447 549 -1445
rect 551 -1447 552 -1445
rect 555 -1441 556 -1439
rect 558 -1441 559 -1439
rect 555 -1447 556 -1445
rect 562 -1441 563 -1439
rect 562 -1447 563 -1445
rect 569 -1441 570 -1439
rect 569 -1447 570 -1445
rect 576 -1441 577 -1439
rect 579 -1441 580 -1439
rect 583 -1441 584 -1439
rect 583 -1447 584 -1445
rect 593 -1441 594 -1439
rect 590 -1447 591 -1445
rect 593 -1447 594 -1445
rect 597 -1441 598 -1439
rect 597 -1447 598 -1445
rect 604 -1441 605 -1439
rect 604 -1447 605 -1445
rect 607 -1447 608 -1445
rect 611 -1441 612 -1439
rect 611 -1447 612 -1445
rect 618 -1441 619 -1439
rect 618 -1447 619 -1445
rect 625 -1441 626 -1439
rect 625 -1447 626 -1445
rect 632 -1441 633 -1439
rect 632 -1447 633 -1445
rect 635 -1447 636 -1445
rect 639 -1441 640 -1439
rect 639 -1447 640 -1445
rect 646 -1441 647 -1439
rect 646 -1447 647 -1445
rect 653 -1447 654 -1445
rect 656 -1447 657 -1445
rect 660 -1441 661 -1439
rect 660 -1447 661 -1445
rect 667 -1441 668 -1439
rect 667 -1447 668 -1445
rect 674 -1441 675 -1439
rect 674 -1447 675 -1445
rect 681 -1441 682 -1439
rect 681 -1447 682 -1445
rect 688 -1441 689 -1439
rect 688 -1447 689 -1445
rect 695 -1441 696 -1439
rect 695 -1447 696 -1445
rect 702 -1441 703 -1439
rect 702 -1447 703 -1445
rect 712 -1441 713 -1439
rect 712 -1447 713 -1445
rect 716 -1441 717 -1439
rect 716 -1447 717 -1445
rect 723 -1441 724 -1439
rect 723 -1447 724 -1445
rect 730 -1441 731 -1439
rect 730 -1447 731 -1445
rect 737 -1441 738 -1439
rect 737 -1447 738 -1445
rect 744 -1441 745 -1439
rect 744 -1447 745 -1445
rect 751 -1441 752 -1439
rect 751 -1447 752 -1445
rect 758 -1441 759 -1439
rect 758 -1447 759 -1445
rect 765 -1441 766 -1439
rect 765 -1447 766 -1445
rect 772 -1441 773 -1439
rect 772 -1447 773 -1445
rect 779 -1441 780 -1439
rect 779 -1447 780 -1445
rect 786 -1441 787 -1439
rect 786 -1447 787 -1445
rect 793 -1441 794 -1439
rect 793 -1447 794 -1445
rect 800 -1441 801 -1439
rect 800 -1447 801 -1445
rect 807 -1441 808 -1439
rect 807 -1447 808 -1445
rect 814 -1441 815 -1439
rect 814 -1447 815 -1445
rect 821 -1441 822 -1439
rect 821 -1447 822 -1445
rect 835 -1441 836 -1439
rect 835 -1447 836 -1445
rect 842 -1441 843 -1439
rect 842 -1447 843 -1445
rect 849 -1441 850 -1439
rect 849 -1447 850 -1445
rect 856 -1441 857 -1439
rect 856 -1447 857 -1445
rect 863 -1441 864 -1439
rect 863 -1447 864 -1445
rect 870 -1441 871 -1439
rect 870 -1447 871 -1445
rect 877 -1441 878 -1439
rect 877 -1447 878 -1445
rect 884 -1441 885 -1439
rect 884 -1447 885 -1445
rect 891 -1441 892 -1439
rect 891 -1447 892 -1445
rect 898 -1441 899 -1439
rect 898 -1447 899 -1445
rect 905 -1441 906 -1439
rect 905 -1447 906 -1445
rect 912 -1441 913 -1439
rect 912 -1447 913 -1445
rect 919 -1441 920 -1439
rect 919 -1447 920 -1445
rect 926 -1441 927 -1439
rect 926 -1447 927 -1445
rect 933 -1441 934 -1439
rect 933 -1447 934 -1445
rect 940 -1441 941 -1439
rect 943 -1441 944 -1439
rect 947 -1441 948 -1439
rect 950 -1447 951 -1445
rect 954 -1441 955 -1439
rect 954 -1447 955 -1445
rect 968 -1441 969 -1439
rect 968 -1447 969 -1445
rect 982 -1441 983 -1439
rect 982 -1447 983 -1445
rect 9 -1530 10 -1528
rect 9 -1536 10 -1534
rect 16 -1530 17 -1528
rect 16 -1536 17 -1534
rect 23 -1530 24 -1528
rect 26 -1536 27 -1534
rect 30 -1530 31 -1528
rect 30 -1536 31 -1534
rect 40 -1530 41 -1528
rect 37 -1536 38 -1534
rect 40 -1536 41 -1534
rect 44 -1530 45 -1528
rect 44 -1536 45 -1534
rect 51 -1530 52 -1528
rect 51 -1536 52 -1534
rect 58 -1530 59 -1528
rect 58 -1536 59 -1534
rect 65 -1530 66 -1528
rect 65 -1536 66 -1534
rect 72 -1536 73 -1534
rect 75 -1536 76 -1534
rect 79 -1530 80 -1528
rect 79 -1536 80 -1534
rect 86 -1530 87 -1528
rect 86 -1536 87 -1534
rect 93 -1530 94 -1528
rect 93 -1536 94 -1534
rect 100 -1530 101 -1528
rect 100 -1536 101 -1534
rect 107 -1530 108 -1528
rect 107 -1536 108 -1534
rect 114 -1530 115 -1528
rect 114 -1536 115 -1534
rect 121 -1530 122 -1528
rect 121 -1536 122 -1534
rect 128 -1530 129 -1528
rect 128 -1536 129 -1534
rect 135 -1536 136 -1534
rect 138 -1536 139 -1534
rect 142 -1530 143 -1528
rect 142 -1536 143 -1534
rect 149 -1530 150 -1528
rect 152 -1530 153 -1528
rect 149 -1536 150 -1534
rect 156 -1530 157 -1528
rect 159 -1530 160 -1528
rect 156 -1536 157 -1534
rect 163 -1530 164 -1528
rect 166 -1530 167 -1528
rect 163 -1536 164 -1534
rect 173 -1530 174 -1528
rect 177 -1530 178 -1528
rect 180 -1530 181 -1528
rect 177 -1536 178 -1534
rect 184 -1530 185 -1528
rect 187 -1530 188 -1528
rect 184 -1536 185 -1534
rect 191 -1530 192 -1528
rect 194 -1530 195 -1528
rect 198 -1530 199 -1528
rect 201 -1530 202 -1528
rect 201 -1536 202 -1534
rect 205 -1530 206 -1528
rect 205 -1536 206 -1534
rect 215 -1536 216 -1534
rect 219 -1530 220 -1528
rect 222 -1530 223 -1528
rect 226 -1530 227 -1528
rect 226 -1536 227 -1534
rect 233 -1530 234 -1528
rect 233 -1536 234 -1534
rect 240 -1530 241 -1528
rect 240 -1536 241 -1534
rect 247 -1530 248 -1528
rect 247 -1536 248 -1534
rect 254 -1530 255 -1528
rect 254 -1536 255 -1534
rect 261 -1530 262 -1528
rect 261 -1536 262 -1534
rect 268 -1530 269 -1528
rect 268 -1536 269 -1534
rect 275 -1530 276 -1528
rect 275 -1536 276 -1534
rect 282 -1530 283 -1528
rect 285 -1530 286 -1528
rect 282 -1536 283 -1534
rect 289 -1530 290 -1528
rect 289 -1536 290 -1534
rect 296 -1530 297 -1528
rect 296 -1536 297 -1534
rect 303 -1530 304 -1528
rect 306 -1530 307 -1528
rect 303 -1536 304 -1534
rect 306 -1536 307 -1534
rect 310 -1530 311 -1528
rect 310 -1536 311 -1534
rect 317 -1530 318 -1528
rect 317 -1536 318 -1534
rect 324 -1530 325 -1528
rect 324 -1536 325 -1534
rect 331 -1530 332 -1528
rect 331 -1536 332 -1534
rect 338 -1530 339 -1528
rect 338 -1536 339 -1534
rect 345 -1530 346 -1528
rect 345 -1536 346 -1534
rect 352 -1530 353 -1528
rect 352 -1536 353 -1534
rect 359 -1530 360 -1528
rect 362 -1530 363 -1528
rect 359 -1536 360 -1534
rect 362 -1536 363 -1534
rect 366 -1530 367 -1528
rect 369 -1530 370 -1528
rect 366 -1536 367 -1534
rect 369 -1536 370 -1534
rect 373 -1530 374 -1528
rect 373 -1536 374 -1534
rect 380 -1530 381 -1528
rect 380 -1536 381 -1534
rect 387 -1530 388 -1528
rect 394 -1530 395 -1528
rect 394 -1536 395 -1534
rect 401 -1530 402 -1528
rect 401 -1536 402 -1534
rect 411 -1530 412 -1528
rect 408 -1536 409 -1534
rect 411 -1536 412 -1534
rect 415 -1530 416 -1528
rect 415 -1536 416 -1534
rect 422 -1530 423 -1528
rect 422 -1536 423 -1534
rect 429 -1530 430 -1528
rect 432 -1530 433 -1528
rect 429 -1536 430 -1534
rect 432 -1536 433 -1534
rect 436 -1530 437 -1528
rect 436 -1536 437 -1534
rect 443 -1530 444 -1528
rect 446 -1530 447 -1528
rect 443 -1536 444 -1534
rect 446 -1536 447 -1534
rect 450 -1530 451 -1528
rect 453 -1530 454 -1528
rect 450 -1536 451 -1534
rect 453 -1536 454 -1534
rect 457 -1530 458 -1528
rect 457 -1536 458 -1534
rect 464 -1530 465 -1528
rect 467 -1530 468 -1528
rect 467 -1536 468 -1534
rect 471 -1530 472 -1528
rect 471 -1536 472 -1534
rect 478 -1530 479 -1528
rect 478 -1536 479 -1534
rect 481 -1536 482 -1534
rect 485 -1530 486 -1528
rect 485 -1536 486 -1534
rect 492 -1530 493 -1528
rect 492 -1536 493 -1534
rect 499 -1530 500 -1528
rect 502 -1530 503 -1528
rect 499 -1536 500 -1534
rect 506 -1530 507 -1528
rect 506 -1536 507 -1534
rect 509 -1536 510 -1534
rect 513 -1530 514 -1528
rect 513 -1536 514 -1534
rect 520 -1530 521 -1528
rect 520 -1536 521 -1534
rect 523 -1536 524 -1534
rect 527 -1530 528 -1528
rect 527 -1536 528 -1534
rect 537 -1530 538 -1528
rect 534 -1536 535 -1534
rect 537 -1536 538 -1534
rect 541 -1530 542 -1528
rect 541 -1536 542 -1534
rect 548 -1530 549 -1528
rect 548 -1536 549 -1534
rect 555 -1530 556 -1528
rect 558 -1530 559 -1528
rect 555 -1536 556 -1534
rect 562 -1530 563 -1528
rect 562 -1536 563 -1534
rect 569 -1530 570 -1528
rect 569 -1536 570 -1534
rect 576 -1530 577 -1528
rect 576 -1536 577 -1534
rect 583 -1530 584 -1528
rect 583 -1536 584 -1534
rect 590 -1530 591 -1528
rect 590 -1536 591 -1534
rect 597 -1530 598 -1528
rect 597 -1536 598 -1534
rect 604 -1530 605 -1528
rect 604 -1536 605 -1534
rect 611 -1530 612 -1528
rect 611 -1536 612 -1534
rect 618 -1530 619 -1528
rect 618 -1536 619 -1534
rect 625 -1530 626 -1528
rect 625 -1536 626 -1534
rect 632 -1530 633 -1528
rect 632 -1536 633 -1534
rect 639 -1530 640 -1528
rect 639 -1536 640 -1534
rect 646 -1530 647 -1528
rect 646 -1536 647 -1534
rect 653 -1530 654 -1528
rect 653 -1536 654 -1534
rect 660 -1530 661 -1528
rect 660 -1536 661 -1534
rect 667 -1530 668 -1528
rect 667 -1536 668 -1534
rect 674 -1530 675 -1528
rect 674 -1536 675 -1534
rect 681 -1530 682 -1528
rect 681 -1536 682 -1534
rect 688 -1530 689 -1528
rect 688 -1536 689 -1534
rect 695 -1530 696 -1528
rect 695 -1536 696 -1534
rect 702 -1530 703 -1528
rect 702 -1536 703 -1534
rect 709 -1530 710 -1528
rect 709 -1536 710 -1534
rect 716 -1530 717 -1528
rect 716 -1536 717 -1534
rect 723 -1530 724 -1528
rect 723 -1536 724 -1534
rect 730 -1530 731 -1528
rect 730 -1536 731 -1534
rect 737 -1530 738 -1528
rect 737 -1536 738 -1534
rect 744 -1530 745 -1528
rect 744 -1536 745 -1534
rect 751 -1530 752 -1528
rect 751 -1536 752 -1534
rect 765 -1530 766 -1528
rect 765 -1536 766 -1534
rect 772 -1530 773 -1528
rect 772 -1536 773 -1534
rect 779 -1530 780 -1528
rect 779 -1536 780 -1534
rect 786 -1530 787 -1528
rect 786 -1536 787 -1534
rect 793 -1530 794 -1528
rect 793 -1536 794 -1534
rect 800 -1530 801 -1528
rect 800 -1536 801 -1534
rect 807 -1530 808 -1528
rect 807 -1536 808 -1534
rect 814 -1530 815 -1528
rect 814 -1536 815 -1534
rect 821 -1530 822 -1528
rect 821 -1536 822 -1534
rect 828 -1530 829 -1528
rect 828 -1536 829 -1534
rect 835 -1530 836 -1528
rect 835 -1536 836 -1534
rect 842 -1530 843 -1528
rect 842 -1536 843 -1534
rect 849 -1530 850 -1528
rect 849 -1536 850 -1534
rect 856 -1530 857 -1528
rect 856 -1536 857 -1534
rect 884 -1530 885 -1528
rect 887 -1530 888 -1528
rect 884 -1536 885 -1534
rect 891 -1530 892 -1528
rect 891 -1536 892 -1534
rect 898 -1530 899 -1528
rect 898 -1536 899 -1534
rect 905 -1530 906 -1528
rect 905 -1536 906 -1534
rect 912 -1530 913 -1528
rect 912 -1536 913 -1534
rect 919 -1530 920 -1528
rect 919 -1536 920 -1534
rect 933 -1530 934 -1528
rect 940 -1530 941 -1528
rect 940 -1536 941 -1534
rect 954 -1530 955 -1528
rect 954 -1536 955 -1534
rect 961 -1530 962 -1528
rect 982 -1530 983 -1528
rect 989 -1530 990 -1528
rect 989 -1536 990 -1534
rect 9 -1621 10 -1619
rect 16 -1615 17 -1613
rect 16 -1621 17 -1619
rect 23 -1615 24 -1613
rect 23 -1621 24 -1619
rect 30 -1615 31 -1613
rect 30 -1621 31 -1619
rect 37 -1615 38 -1613
rect 37 -1621 38 -1619
rect 44 -1615 45 -1613
rect 44 -1621 45 -1619
rect 51 -1615 52 -1613
rect 51 -1621 52 -1619
rect 58 -1615 59 -1613
rect 58 -1621 59 -1619
rect 65 -1615 66 -1613
rect 65 -1621 66 -1619
rect 72 -1615 73 -1613
rect 72 -1621 73 -1619
rect 79 -1615 80 -1613
rect 79 -1621 80 -1619
rect 86 -1615 87 -1613
rect 86 -1621 87 -1619
rect 96 -1615 97 -1613
rect 93 -1621 94 -1619
rect 96 -1621 97 -1619
rect 100 -1615 101 -1613
rect 100 -1621 101 -1619
rect 110 -1615 111 -1613
rect 110 -1621 111 -1619
rect 121 -1615 122 -1613
rect 124 -1621 125 -1619
rect 128 -1615 129 -1613
rect 128 -1621 129 -1619
rect 135 -1615 136 -1613
rect 135 -1621 136 -1619
rect 142 -1615 143 -1613
rect 142 -1621 143 -1619
rect 149 -1615 150 -1613
rect 149 -1621 150 -1619
rect 156 -1615 157 -1613
rect 159 -1615 160 -1613
rect 156 -1621 157 -1619
rect 166 -1615 167 -1613
rect 163 -1621 164 -1619
rect 166 -1621 167 -1619
rect 173 -1615 174 -1613
rect 170 -1621 171 -1619
rect 173 -1621 174 -1619
rect 177 -1615 178 -1613
rect 177 -1621 178 -1619
rect 184 -1621 185 -1619
rect 187 -1621 188 -1619
rect 194 -1615 195 -1613
rect 191 -1621 192 -1619
rect 198 -1615 199 -1613
rect 198 -1621 199 -1619
rect 205 -1621 206 -1619
rect 208 -1621 209 -1619
rect 212 -1615 213 -1613
rect 212 -1621 213 -1619
rect 219 -1615 220 -1613
rect 219 -1621 220 -1619
rect 226 -1615 227 -1613
rect 226 -1621 227 -1619
rect 233 -1615 234 -1613
rect 233 -1621 234 -1619
rect 240 -1615 241 -1613
rect 240 -1621 241 -1619
rect 247 -1615 248 -1613
rect 247 -1621 248 -1619
rect 254 -1615 255 -1613
rect 254 -1621 255 -1619
rect 261 -1615 262 -1613
rect 261 -1621 262 -1619
rect 268 -1615 269 -1613
rect 268 -1621 269 -1619
rect 275 -1615 276 -1613
rect 275 -1621 276 -1619
rect 282 -1615 283 -1613
rect 282 -1621 283 -1619
rect 289 -1615 290 -1613
rect 292 -1615 293 -1613
rect 296 -1615 297 -1613
rect 296 -1621 297 -1619
rect 303 -1615 304 -1613
rect 303 -1621 304 -1619
rect 310 -1615 311 -1613
rect 310 -1621 311 -1619
rect 317 -1615 318 -1613
rect 317 -1621 318 -1619
rect 324 -1615 325 -1613
rect 324 -1621 325 -1619
rect 331 -1615 332 -1613
rect 331 -1621 332 -1619
rect 338 -1615 339 -1613
rect 341 -1615 342 -1613
rect 338 -1621 339 -1619
rect 341 -1621 342 -1619
rect 345 -1615 346 -1613
rect 348 -1615 349 -1613
rect 345 -1621 346 -1619
rect 348 -1621 349 -1619
rect 352 -1615 353 -1613
rect 352 -1621 353 -1619
rect 359 -1615 360 -1613
rect 362 -1615 363 -1613
rect 366 -1615 367 -1613
rect 366 -1621 367 -1619
rect 373 -1615 374 -1613
rect 373 -1621 374 -1619
rect 383 -1621 384 -1619
rect 387 -1621 388 -1619
rect 394 -1615 395 -1613
rect 394 -1621 395 -1619
rect 401 -1615 402 -1613
rect 401 -1621 402 -1619
rect 408 -1615 409 -1613
rect 408 -1621 409 -1619
rect 415 -1615 416 -1613
rect 415 -1621 416 -1619
rect 422 -1621 423 -1619
rect 425 -1621 426 -1619
rect 429 -1615 430 -1613
rect 429 -1621 430 -1619
rect 436 -1615 437 -1613
rect 436 -1621 437 -1619
rect 443 -1615 444 -1613
rect 443 -1621 444 -1619
rect 453 -1615 454 -1613
rect 450 -1621 451 -1619
rect 453 -1621 454 -1619
rect 457 -1615 458 -1613
rect 457 -1621 458 -1619
rect 464 -1615 465 -1613
rect 464 -1621 465 -1619
rect 471 -1615 472 -1613
rect 471 -1621 472 -1619
rect 478 -1615 479 -1613
rect 481 -1615 482 -1613
rect 481 -1621 482 -1619
rect 485 -1615 486 -1613
rect 485 -1621 486 -1619
rect 492 -1615 493 -1613
rect 492 -1621 493 -1619
rect 495 -1621 496 -1619
rect 499 -1615 500 -1613
rect 499 -1621 500 -1619
rect 506 -1615 507 -1613
rect 506 -1621 507 -1619
rect 513 -1615 514 -1613
rect 513 -1621 514 -1619
rect 520 -1615 521 -1613
rect 523 -1615 524 -1613
rect 520 -1621 521 -1619
rect 530 -1615 531 -1613
rect 527 -1621 528 -1619
rect 534 -1615 535 -1613
rect 537 -1615 538 -1613
rect 534 -1621 535 -1619
rect 537 -1621 538 -1619
rect 541 -1615 542 -1613
rect 541 -1621 542 -1619
rect 548 -1615 549 -1613
rect 548 -1621 549 -1619
rect 555 -1615 556 -1613
rect 555 -1621 556 -1619
rect 562 -1615 563 -1613
rect 565 -1615 566 -1613
rect 562 -1621 563 -1619
rect 565 -1621 566 -1619
rect 569 -1615 570 -1613
rect 569 -1621 570 -1619
rect 576 -1615 577 -1613
rect 576 -1621 577 -1619
rect 586 -1615 587 -1613
rect 583 -1621 584 -1619
rect 586 -1621 587 -1619
rect 590 -1615 591 -1613
rect 590 -1621 591 -1619
rect 597 -1615 598 -1613
rect 597 -1621 598 -1619
rect 604 -1615 605 -1613
rect 604 -1621 605 -1619
rect 611 -1615 612 -1613
rect 611 -1621 612 -1619
rect 625 -1615 626 -1613
rect 625 -1621 626 -1619
rect 632 -1615 633 -1613
rect 632 -1621 633 -1619
rect 639 -1615 640 -1613
rect 639 -1621 640 -1619
rect 646 -1615 647 -1613
rect 646 -1621 647 -1619
rect 653 -1615 654 -1613
rect 653 -1621 654 -1619
rect 660 -1615 661 -1613
rect 660 -1621 661 -1619
rect 667 -1615 668 -1613
rect 667 -1621 668 -1619
rect 674 -1615 675 -1613
rect 674 -1621 675 -1619
rect 681 -1615 682 -1613
rect 681 -1621 682 -1619
rect 688 -1615 689 -1613
rect 688 -1621 689 -1619
rect 695 -1615 696 -1613
rect 695 -1621 696 -1619
rect 702 -1615 703 -1613
rect 705 -1615 706 -1613
rect 702 -1621 703 -1619
rect 705 -1621 706 -1619
rect 709 -1615 710 -1613
rect 709 -1621 710 -1619
rect 716 -1615 717 -1613
rect 716 -1621 717 -1619
rect 723 -1615 724 -1613
rect 723 -1621 724 -1619
rect 733 -1615 734 -1613
rect 730 -1621 731 -1619
rect 733 -1621 734 -1619
rect 744 -1615 745 -1613
rect 744 -1621 745 -1619
rect 751 -1615 752 -1613
rect 751 -1621 752 -1619
rect 758 -1615 759 -1613
rect 758 -1621 759 -1619
rect 765 -1615 766 -1613
rect 765 -1621 766 -1619
rect 786 -1615 787 -1613
rect 786 -1621 787 -1619
rect 793 -1615 794 -1613
rect 793 -1621 794 -1619
rect 800 -1615 801 -1613
rect 800 -1621 801 -1619
rect 814 -1615 815 -1613
rect 814 -1621 815 -1619
rect 828 -1615 829 -1613
rect 828 -1621 829 -1619
rect 842 -1615 843 -1613
rect 842 -1621 843 -1619
rect 849 -1615 850 -1613
rect 852 -1615 853 -1613
rect 849 -1621 850 -1619
rect 856 -1615 857 -1613
rect 856 -1621 857 -1619
rect 870 -1615 871 -1613
rect 870 -1621 871 -1619
rect 880 -1615 881 -1613
rect 877 -1621 878 -1619
rect 898 -1615 899 -1613
rect 898 -1621 899 -1619
rect 915 -1615 916 -1613
rect 919 -1615 920 -1613
rect 919 -1621 920 -1619
rect 926 -1615 927 -1613
rect 926 -1621 927 -1619
rect 940 -1615 941 -1613
rect 940 -1621 941 -1619
rect 943 -1621 944 -1619
rect 947 -1615 948 -1613
rect 947 -1621 948 -1619
rect 954 -1615 955 -1613
rect 954 -1621 955 -1619
rect 968 -1615 969 -1613
rect 971 -1615 972 -1613
rect 975 -1615 976 -1613
rect 975 -1621 976 -1619
rect 982 -1615 983 -1613
rect 982 -1621 983 -1619
rect 9 -1708 10 -1706
rect 9 -1714 10 -1712
rect 16 -1708 17 -1706
rect 16 -1714 17 -1712
rect 23 -1708 24 -1706
rect 23 -1714 24 -1712
rect 30 -1708 31 -1706
rect 30 -1714 31 -1712
rect 37 -1708 38 -1706
rect 37 -1714 38 -1712
rect 44 -1708 45 -1706
rect 44 -1714 45 -1712
rect 51 -1708 52 -1706
rect 51 -1714 52 -1712
rect 58 -1708 59 -1706
rect 61 -1708 62 -1706
rect 58 -1714 59 -1712
rect 65 -1708 66 -1706
rect 65 -1714 66 -1712
rect 75 -1714 76 -1712
rect 79 -1708 80 -1706
rect 79 -1714 80 -1712
rect 86 -1708 87 -1706
rect 86 -1714 87 -1712
rect 93 -1708 94 -1706
rect 93 -1714 94 -1712
rect 103 -1708 104 -1706
rect 103 -1714 104 -1712
rect 107 -1708 108 -1706
rect 107 -1714 108 -1712
rect 117 -1708 118 -1706
rect 117 -1714 118 -1712
rect 121 -1708 122 -1706
rect 121 -1714 122 -1712
rect 128 -1708 129 -1706
rect 128 -1714 129 -1712
rect 135 -1708 136 -1706
rect 135 -1714 136 -1712
rect 142 -1708 143 -1706
rect 145 -1708 146 -1706
rect 149 -1708 150 -1706
rect 152 -1708 153 -1706
rect 156 -1708 157 -1706
rect 156 -1714 157 -1712
rect 163 -1708 164 -1706
rect 163 -1714 164 -1712
rect 173 -1708 174 -1706
rect 170 -1714 171 -1712
rect 180 -1708 181 -1706
rect 184 -1708 185 -1706
rect 184 -1714 185 -1712
rect 191 -1708 192 -1706
rect 191 -1714 192 -1712
rect 198 -1708 199 -1706
rect 198 -1714 199 -1712
rect 205 -1708 206 -1706
rect 208 -1708 209 -1706
rect 212 -1708 213 -1706
rect 212 -1714 213 -1712
rect 219 -1708 220 -1706
rect 219 -1714 220 -1712
rect 226 -1708 227 -1706
rect 226 -1714 227 -1712
rect 233 -1714 234 -1712
rect 236 -1714 237 -1712
rect 240 -1708 241 -1706
rect 240 -1714 241 -1712
rect 247 -1708 248 -1706
rect 247 -1714 248 -1712
rect 254 -1708 255 -1706
rect 254 -1714 255 -1712
rect 261 -1708 262 -1706
rect 261 -1714 262 -1712
rect 268 -1708 269 -1706
rect 268 -1714 269 -1712
rect 275 -1708 276 -1706
rect 275 -1714 276 -1712
rect 282 -1708 283 -1706
rect 282 -1714 283 -1712
rect 289 -1708 290 -1706
rect 289 -1714 290 -1712
rect 296 -1708 297 -1706
rect 299 -1708 300 -1706
rect 296 -1714 297 -1712
rect 299 -1714 300 -1712
rect 303 -1708 304 -1706
rect 303 -1714 304 -1712
rect 310 -1708 311 -1706
rect 310 -1714 311 -1712
rect 317 -1708 318 -1706
rect 317 -1714 318 -1712
rect 324 -1708 325 -1706
rect 324 -1714 325 -1712
rect 331 -1708 332 -1706
rect 331 -1714 332 -1712
rect 334 -1714 335 -1712
rect 341 -1708 342 -1706
rect 338 -1714 339 -1712
rect 341 -1714 342 -1712
rect 345 -1708 346 -1706
rect 345 -1714 346 -1712
rect 352 -1708 353 -1706
rect 352 -1714 353 -1712
rect 359 -1708 360 -1706
rect 359 -1714 360 -1712
rect 366 -1708 367 -1706
rect 366 -1714 367 -1712
rect 373 -1714 374 -1712
rect 376 -1714 377 -1712
rect 380 -1708 381 -1706
rect 380 -1714 381 -1712
rect 387 -1708 388 -1706
rect 390 -1708 391 -1706
rect 387 -1714 388 -1712
rect 397 -1708 398 -1706
rect 394 -1714 395 -1712
rect 397 -1714 398 -1712
rect 401 -1708 402 -1706
rect 404 -1708 405 -1706
rect 401 -1714 402 -1712
rect 408 -1708 409 -1706
rect 408 -1714 409 -1712
rect 415 -1708 416 -1706
rect 415 -1714 416 -1712
rect 422 -1708 423 -1706
rect 422 -1714 423 -1712
rect 429 -1708 430 -1706
rect 429 -1714 430 -1712
rect 436 -1708 437 -1706
rect 439 -1708 440 -1706
rect 439 -1714 440 -1712
rect 443 -1708 444 -1706
rect 443 -1714 444 -1712
rect 450 -1708 451 -1706
rect 450 -1714 451 -1712
rect 453 -1714 454 -1712
rect 457 -1708 458 -1706
rect 457 -1714 458 -1712
rect 464 -1708 465 -1706
rect 464 -1714 465 -1712
rect 467 -1714 468 -1712
rect 471 -1708 472 -1706
rect 471 -1714 472 -1712
rect 478 -1708 479 -1706
rect 478 -1714 479 -1712
rect 488 -1708 489 -1706
rect 485 -1714 486 -1712
rect 488 -1714 489 -1712
rect 492 -1708 493 -1706
rect 492 -1714 493 -1712
rect 499 -1708 500 -1706
rect 499 -1714 500 -1712
rect 509 -1708 510 -1706
rect 509 -1714 510 -1712
rect 513 -1708 514 -1706
rect 513 -1714 514 -1712
rect 520 -1708 521 -1706
rect 520 -1714 521 -1712
rect 527 -1708 528 -1706
rect 527 -1714 528 -1712
rect 534 -1708 535 -1706
rect 534 -1714 535 -1712
rect 541 -1708 542 -1706
rect 544 -1708 545 -1706
rect 541 -1714 542 -1712
rect 548 -1708 549 -1706
rect 548 -1714 549 -1712
rect 555 -1708 556 -1706
rect 555 -1714 556 -1712
rect 562 -1708 563 -1706
rect 562 -1714 563 -1712
rect 569 -1708 570 -1706
rect 572 -1708 573 -1706
rect 572 -1714 573 -1712
rect 576 -1708 577 -1706
rect 576 -1714 577 -1712
rect 583 -1708 584 -1706
rect 583 -1714 584 -1712
rect 590 -1708 591 -1706
rect 590 -1714 591 -1712
rect 597 -1708 598 -1706
rect 597 -1714 598 -1712
rect 604 -1708 605 -1706
rect 604 -1714 605 -1712
rect 611 -1708 612 -1706
rect 611 -1714 612 -1712
rect 618 -1708 619 -1706
rect 618 -1714 619 -1712
rect 625 -1708 626 -1706
rect 625 -1714 626 -1712
rect 632 -1708 633 -1706
rect 632 -1714 633 -1712
rect 639 -1708 640 -1706
rect 639 -1714 640 -1712
rect 646 -1708 647 -1706
rect 646 -1714 647 -1712
rect 653 -1708 654 -1706
rect 653 -1714 654 -1712
rect 660 -1708 661 -1706
rect 660 -1714 661 -1712
rect 667 -1708 668 -1706
rect 667 -1714 668 -1712
rect 674 -1708 675 -1706
rect 674 -1714 675 -1712
rect 681 -1708 682 -1706
rect 681 -1714 682 -1712
rect 688 -1708 689 -1706
rect 688 -1714 689 -1712
rect 695 -1708 696 -1706
rect 695 -1714 696 -1712
rect 702 -1708 703 -1706
rect 702 -1714 703 -1712
rect 712 -1708 713 -1706
rect 716 -1708 717 -1706
rect 716 -1714 717 -1712
rect 723 -1708 724 -1706
rect 723 -1714 724 -1712
rect 730 -1708 731 -1706
rect 730 -1714 731 -1712
rect 737 -1708 738 -1706
rect 737 -1714 738 -1712
rect 744 -1708 745 -1706
rect 744 -1714 745 -1712
rect 751 -1708 752 -1706
rect 751 -1714 752 -1712
rect 758 -1708 759 -1706
rect 758 -1714 759 -1712
rect 765 -1708 766 -1706
rect 765 -1714 766 -1712
rect 772 -1708 773 -1706
rect 772 -1714 773 -1712
rect 779 -1708 780 -1706
rect 779 -1714 780 -1712
rect 786 -1708 787 -1706
rect 786 -1714 787 -1712
rect 800 -1708 801 -1706
rect 800 -1714 801 -1712
rect 814 -1708 815 -1706
rect 814 -1714 815 -1712
rect 821 -1708 822 -1706
rect 821 -1714 822 -1712
rect 828 -1708 829 -1706
rect 828 -1714 829 -1712
rect 835 -1708 836 -1706
rect 835 -1714 836 -1712
rect 842 -1708 843 -1706
rect 842 -1714 843 -1712
rect 863 -1708 864 -1706
rect 863 -1714 864 -1712
rect 870 -1708 871 -1706
rect 870 -1714 871 -1712
rect 887 -1708 888 -1706
rect 887 -1714 888 -1712
rect 894 -1708 895 -1706
rect 912 -1708 913 -1706
rect 912 -1714 913 -1712
rect 926 -1708 927 -1706
rect 926 -1714 927 -1712
rect 940 -1714 941 -1712
rect 961 -1708 962 -1706
rect 961 -1714 962 -1712
rect 971 -1708 972 -1706
rect 975 -1708 976 -1706
rect 978 -1714 979 -1712
rect 9 -1803 10 -1801
rect 9 -1809 10 -1807
rect 12 -1809 13 -1807
rect 16 -1803 17 -1801
rect 16 -1809 17 -1807
rect 23 -1803 24 -1801
rect 23 -1809 24 -1807
rect 30 -1803 31 -1801
rect 30 -1809 31 -1807
rect 37 -1803 38 -1801
rect 40 -1809 41 -1807
rect 44 -1803 45 -1801
rect 44 -1809 45 -1807
rect 51 -1803 52 -1801
rect 58 -1803 59 -1801
rect 58 -1809 59 -1807
rect 65 -1803 66 -1801
rect 65 -1809 66 -1807
rect 72 -1803 73 -1801
rect 72 -1809 73 -1807
rect 82 -1803 83 -1801
rect 82 -1809 83 -1807
rect 86 -1803 87 -1801
rect 89 -1809 90 -1807
rect 93 -1803 94 -1801
rect 93 -1809 94 -1807
rect 103 -1803 104 -1801
rect 103 -1809 104 -1807
rect 107 -1803 108 -1801
rect 107 -1809 108 -1807
rect 114 -1803 115 -1801
rect 117 -1803 118 -1801
rect 114 -1809 115 -1807
rect 124 -1803 125 -1801
rect 121 -1809 122 -1807
rect 124 -1809 125 -1807
rect 128 -1809 129 -1807
rect 135 -1809 136 -1807
rect 138 -1809 139 -1807
rect 142 -1803 143 -1801
rect 142 -1809 143 -1807
rect 149 -1803 150 -1801
rect 149 -1809 150 -1807
rect 156 -1803 157 -1801
rect 159 -1803 160 -1801
rect 166 -1803 167 -1801
rect 163 -1809 164 -1807
rect 166 -1809 167 -1807
rect 170 -1803 171 -1801
rect 173 -1803 174 -1801
rect 170 -1809 171 -1807
rect 173 -1809 174 -1807
rect 180 -1803 181 -1801
rect 180 -1809 181 -1807
rect 184 -1803 185 -1801
rect 187 -1803 188 -1801
rect 187 -1809 188 -1807
rect 191 -1803 192 -1801
rect 191 -1809 192 -1807
rect 198 -1803 199 -1801
rect 198 -1809 199 -1807
rect 205 -1803 206 -1801
rect 205 -1809 206 -1807
rect 212 -1803 213 -1801
rect 215 -1809 216 -1807
rect 219 -1803 220 -1801
rect 222 -1803 223 -1801
rect 219 -1809 220 -1807
rect 222 -1809 223 -1807
rect 226 -1803 227 -1801
rect 226 -1809 227 -1807
rect 233 -1803 234 -1801
rect 233 -1809 234 -1807
rect 240 -1803 241 -1801
rect 240 -1809 241 -1807
rect 247 -1803 248 -1801
rect 247 -1809 248 -1807
rect 254 -1803 255 -1801
rect 254 -1809 255 -1807
rect 261 -1803 262 -1801
rect 261 -1809 262 -1807
rect 271 -1803 272 -1801
rect 268 -1809 269 -1807
rect 275 -1803 276 -1801
rect 275 -1809 276 -1807
rect 282 -1803 283 -1801
rect 282 -1809 283 -1807
rect 289 -1803 290 -1801
rect 289 -1809 290 -1807
rect 296 -1803 297 -1801
rect 296 -1809 297 -1807
rect 303 -1803 304 -1801
rect 303 -1809 304 -1807
rect 310 -1803 311 -1801
rect 310 -1809 311 -1807
rect 320 -1803 321 -1801
rect 317 -1809 318 -1807
rect 324 -1803 325 -1801
rect 324 -1809 325 -1807
rect 331 -1803 332 -1801
rect 331 -1809 332 -1807
rect 338 -1803 339 -1801
rect 338 -1809 339 -1807
rect 345 -1803 346 -1801
rect 345 -1809 346 -1807
rect 352 -1803 353 -1801
rect 355 -1803 356 -1801
rect 352 -1809 353 -1807
rect 355 -1809 356 -1807
rect 359 -1803 360 -1801
rect 359 -1809 360 -1807
rect 369 -1803 370 -1801
rect 369 -1809 370 -1807
rect 376 -1803 377 -1801
rect 373 -1809 374 -1807
rect 383 -1803 384 -1801
rect 380 -1809 381 -1807
rect 387 -1803 388 -1801
rect 387 -1809 388 -1807
rect 394 -1809 395 -1807
rect 401 -1803 402 -1801
rect 401 -1809 402 -1807
rect 408 -1803 409 -1801
rect 408 -1809 409 -1807
rect 415 -1803 416 -1801
rect 415 -1809 416 -1807
rect 422 -1803 423 -1801
rect 422 -1809 423 -1807
rect 429 -1803 430 -1801
rect 429 -1809 430 -1807
rect 436 -1803 437 -1801
rect 436 -1809 437 -1807
rect 443 -1803 444 -1801
rect 443 -1809 444 -1807
rect 450 -1803 451 -1801
rect 450 -1809 451 -1807
rect 457 -1803 458 -1801
rect 457 -1809 458 -1807
rect 464 -1803 465 -1801
rect 464 -1809 465 -1807
rect 471 -1803 472 -1801
rect 474 -1803 475 -1801
rect 478 -1803 479 -1801
rect 478 -1809 479 -1807
rect 485 -1803 486 -1801
rect 485 -1809 486 -1807
rect 495 -1803 496 -1801
rect 492 -1809 493 -1807
rect 495 -1809 496 -1807
rect 499 -1803 500 -1801
rect 499 -1809 500 -1807
rect 506 -1803 507 -1801
rect 506 -1809 507 -1807
rect 509 -1809 510 -1807
rect 513 -1803 514 -1801
rect 516 -1809 517 -1807
rect 523 -1803 524 -1801
rect 527 -1803 528 -1801
rect 527 -1809 528 -1807
rect 534 -1803 535 -1801
rect 534 -1809 535 -1807
rect 541 -1803 542 -1801
rect 541 -1809 542 -1807
rect 548 -1803 549 -1801
rect 548 -1809 549 -1807
rect 555 -1803 556 -1801
rect 555 -1809 556 -1807
rect 562 -1803 563 -1801
rect 562 -1809 563 -1807
rect 569 -1803 570 -1801
rect 569 -1809 570 -1807
rect 576 -1803 577 -1801
rect 576 -1809 577 -1807
rect 583 -1803 584 -1801
rect 583 -1809 584 -1807
rect 590 -1803 591 -1801
rect 590 -1809 591 -1807
rect 597 -1803 598 -1801
rect 597 -1809 598 -1807
rect 604 -1803 605 -1801
rect 604 -1809 605 -1807
rect 611 -1803 612 -1801
rect 611 -1809 612 -1807
rect 618 -1803 619 -1801
rect 618 -1809 619 -1807
rect 625 -1803 626 -1801
rect 625 -1809 626 -1807
rect 632 -1803 633 -1801
rect 632 -1809 633 -1807
rect 639 -1803 640 -1801
rect 642 -1803 643 -1801
rect 646 -1803 647 -1801
rect 646 -1809 647 -1807
rect 653 -1803 654 -1801
rect 653 -1809 654 -1807
rect 660 -1803 661 -1801
rect 660 -1809 661 -1807
rect 667 -1803 668 -1801
rect 667 -1809 668 -1807
rect 674 -1803 675 -1801
rect 674 -1809 675 -1807
rect 681 -1803 682 -1801
rect 681 -1809 682 -1807
rect 688 -1803 689 -1801
rect 688 -1809 689 -1807
rect 695 -1803 696 -1801
rect 695 -1809 696 -1807
rect 702 -1803 703 -1801
rect 702 -1809 703 -1807
rect 709 -1803 710 -1801
rect 709 -1809 710 -1807
rect 716 -1803 717 -1801
rect 716 -1809 717 -1807
rect 723 -1803 724 -1801
rect 723 -1809 724 -1807
rect 730 -1803 731 -1801
rect 730 -1809 731 -1807
rect 737 -1803 738 -1801
rect 737 -1809 738 -1807
rect 744 -1803 745 -1801
rect 744 -1809 745 -1807
rect 751 -1803 752 -1801
rect 751 -1809 752 -1807
rect 758 -1803 759 -1801
rect 758 -1809 759 -1807
rect 905 -1803 906 -1801
rect 5 -1890 6 -1888
rect 12 -1890 13 -1888
rect 16 -1884 17 -1882
rect 16 -1890 17 -1888
rect 23 -1890 24 -1888
rect 26 -1890 27 -1888
rect 33 -1884 34 -1882
rect 37 -1884 38 -1882
rect 37 -1890 38 -1888
rect 47 -1884 48 -1882
rect 51 -1884 52 -1882
rect 51 -1890 52 -1888
rect 58 -1884 59 -1882
rect 58 -1890 59 -1888
rect 65 -1884 66 -1882
rect 65 -1890 66 -1888
rect 72 -1884 73 -1882
rect 72 -1890 73 -1888
rect 79 -1884 80 -1882
rect 79 -1890 80 -1888
rect 86 -1884 87 -1882
rect 86 -1890 87 -1888
rect 93 -1884 94 -1882
rect 93 -1890 94 -1888
rect 100 -1884 101 -1882
rect 100 -1890 101 -1888
rect 107 -1884 108 -1882
rect 107 -1890 108 -1888
rect 114 -1884 115 -1882
rect 114 -1890 115 -1888
rect 121 -1884 122 -1882
rect 121 -1890 122 -1888
rect 131 -1884 132 -1882
rect 131 -1890 132 -1888
rect 135 -1884 136 -1882
rect 135 -1890 136 -1888
rect 142 -1884 143 -1882
rect 142 -1890 143 -1888
rect 145 -1890 146 -1888
rect 149 -1890 150 -1888
rect 156 -1884 157 -1882
rect 156 -1890 157 -1888
rect 163 -1884 164 -1882
rect 166 -1890 167 -1888
rect 170 -1884 171 -1882
rect 170 -1890 171 -1888
rect 177 -1884 178 -1882
rect 177 -1890 178 -1888
rect 184 -1884 185 -1882
rect 184 -1890 185 -1888
rect 191 -1884 192 -1882
rect 194 -1890 195 -1888
rect 198 -1884 199 -1882
rect 201 -1884 202 -1882
rect 198 -1890 199 -1888
rect 205 -1884 206 -1882
rect 205 -1890 206 -1888
rect 212 -1884 213 -1882
rect 212 -1890 213 -1888
rect 219 -1884 220 -1882
rect 219 -1890 220 -1888
rect 226 -1884 227 -1882
rect 233 -1884 234 -1882
rect 233 -1890 234 -1888
rect 240 -1884 241 -1882
rect 240 -1890 241 -1888
rect 247 -1884 248 -1882
rect 247 -1890 248 -1888
rect 254 -1884 255 -1882
rect 254 -1890 255 -1888
rect 261 -1884 262 -1882
rect 261 -1890 262 -1888
rect 268 -1884 269 -1882
rect 268 -1890 269 -1888
rect 275 -1884 276 -1882
rect 275 -1890 276 -1888
rect 282 -1884 283 -1882
rect 282 -1890 283 -1888
rect 292 -1884 293 -1882
rect 292 -1890 293 -1888
rect 296 -1884 297 -1882
rect 296 -1890 297 -1888
rect 303 -1884 304 -1882
rect 306 -1884 307 -1882
rect 303 -1890 304 -1888
rect 306 -1890 307 -1888
rect 310 -1884 311 -1882
rect 310 -1890 311 -1888
rect 317 -1884 318 -1882
rect 317 -1890 318 -1888
rect 324 -1884 325 -1882
rect 324 -1890 325 -1888
rect 327 -1890 328 -1888
rect 331 -1884 332 -1882
rect 331 -1890 332 -1888
rect 338 -1884 339 -1882
rect 348 -1884 349 -1882
rect 352 -1884 353 -1882
rect 355 -1884 356 -1882
rect 362 -1884 363 -1882
rect 359 -1890 360 -1888
rect 362 -1890 363 -1888
rect 366 -1884 367 -1882
rect 366 -1890 367 -1888
rect 373 -1884 374 -1882
rect 376 -1884 377 -1882
rect 376 -1890 377 -1888
rect 380 -1884 381 -1882
rect 380 -1890 381 -1888
rect 387 -1884 388 -1882
rect 390 -1884 391 -1882
rect 387 -1890 388 -1888
rect 394 -1884 395 -1882
rect 394 -1890 395 -1888
rect 401 -1884 402 -1882
rect 401 -1890 402 -1888
rect 408 -1884 409 -1882
rect 408 -1890 409 -1888
rect 415 -1884 416 -1882
rect 415 -1890 416 -1888
rect 422 -1884 423 -1882
rect 422 -1890 423 -1888
rect 429 -1884 430 -1882
rect 429 -1890 430 -1888
rect 436 -1890 437 -1888
rect 439 -1890 440 -1888
rect 443 -1884 444 -1882
rect 450 -1884 451 -1882
rect 453 -1884 454 -1882
rect 450 -1890 451 -1888
rect 457 -1884 458 -1882
rect 457 -1890 458 -1888
rect 464 -1884 465 -1882
rect 464 -1890 465 -1888
rect 467 -1890 468 -1888
rect 471 -1884 472 -1882
rect 471 -1890 472 -1888
rect 478 -1884 479 -1882
rect 478 -1890 479 -1888
rect 485 -1884 486 -1882
rect 485 -1890 486 -1888
rect 492 -1884 493 -1882
rect 492 -1890 493 -1888
rect 499 -1884 500 -1882
rect 502 -1884 503 -1882
rect 502 -1890 503 -1888
rect 506 -1884 507 -1882
rect 506 -1890 507 -1888
rect 513 -1884 514 -1882
rect 513 -1890 514 -1888
rect 520 -1884 521 -1882
rect 520 -1890 521 -1888
rect 527 -1884 528 -1882
rect 527 -1890 528 -1888
rect 534 -1884 535 -1882
rect 534 -1890 535 -1888
rect 541 -1884 542 -1882
rect 541 -1890 542 -1888
rect 548 -1890 549 -1888
rect 555 -1884 556 -1882
rect 555 -1890 556 -1888
rect 562 -1884 563 -1882
rect 562 -1890 563 -1888
rect 569 -1884 570 -1882
rect 569 -1890 570 -1888
rect 579 -1884 580 -1882
rect 579 -1890 580 -1888
rect 583 -1884 584 -1882
rect 583 -1890 584 -1888
rect 590 -1884 591 -1882
rect 590 -1890 591 -1888
rect 597 -1884 598 -1882
rect 597 -1890 598 -1888
rect 604 -1884 605 -1882
rect 604 -1890 605 -1888
rect 611 -1884 612 -1882
rect 611 -1890 612 -1888
rect 618 -1884 619 -1882
rect 618 -1890 619 -1888
rect 625 -1884 626 -1882
rect 625 -1890 626 -1888
rect 632 -1884 633 -1882
rect 632 -1890 633 -1888
rect 642 -1884 643 -1882
rect 639 -1890 640 -1888
rect 646 -1884 647 -1882
rect 646 -1890 647 -1888
rect 653 -1884 654 -1882
rect 653 -1890 654 -1888
rect 660 -1884 661 -1882
rect 660 -1890 661 -1888
rect 667 -1884 668 -1882
rect 667 -1890 668 -1888
rect 674 -1884 675 -1882
rect 674 -1890 675 -1888
rect 681 -1884 682 -1882
rect 681 -1890 682 -1888
rect 688 -1884 689 -1882
rect 688 -1890 689 -1888
rect 695 -1884 696 -1882
rect 695 -1890 696 -1888
rect 702 -1884 703 -1882
rect 702 -1890 703 -1888
rect 709 -1884 710 -1882
rect 709 -1890 710 -1888
rect 716 -1884 717 -1882
rect 716 -1890 717 -1888
rect 723 -1884 724 -1882
rect 723 -1890 724 -1888
rect 730 -1884 731 -1882
rect 730 -1890 731 -1888
rect 737 -1884 738 -1882
rect 737 -1890 738 -1888
rect 744 -1884 745 -1882
rect 747 -1884 748 -1882
rect 747 -1890 748 -1888
rect 751 -1884 752 -1882
rect 751 -1890 752 -1888
rect 2 -1967 3 -1965
rect 2 -1973 3 -1971
rect 9 -1967 10 -1965
rect 9 -1973 10 -1971
rect 19 -1967 20 -1965
rect 19 -1973 20 -1971
rect 23 -1967 24 -1965
rect 23 -1973 24 -1971
rect 33 -1967 34 -1965
rect 30 -1973 31 -1971
rect 37 -1967 38 -1965
rect 44 -1967 45 -1965
rect 44 -1973 45 -1971
rect 51 -1967 52 -1965
rect 54 -1967 55 -1965
rect 54 -1973 55 -1971
rect 61 -1967 62 -1965
rect 65 -1967 66 -1965
rect 65 -1973 66 -1971
rect 72 -1967 73 -1965
rect 75 -1973 76 -1971
rect 79 -1967 80 -1965
rect 86 -1967 87 -1965
rect 86 -1973 87 -1971
rect 93 -1967 94 -1965
rect 93 -1973 94 -1971
rect 100 -1967 101 -1965
rect 100 -1973 101 -1971
rect 107 -1973 108 -1971
rect 110 -1973 111 -1971
rect 117 -1967 118 -1965
rect 117 -1973 118 -1971
rect 121 -1967 122 -1965
rect 121 -1973 122 -1971
rect 128 -1967 129 -1965
rect 128 -1973 129 -1971
rect 135 -1967 136 -1965
rect 135 -1973 136 -1971
rect 142 -1967 143 -1965
rect 142 -1973 143 -1971
rect 149 -1967 150 -1965
rect 149 -1973 150 -1971
rect 156 -1967 157 -1965
rect 156 -1973 157 -1971
rect 159 -1973 160 -1971
rect 163 -1967 164 -1965
rect 163 -1973 164 -1971
rect 170 -1967 171 -1965
rect 170 -1973 171 -1971
rect 173 -1973 174 -1971
rect 177 -1967 178 -1965
rect 177 -1973 178 -1971
rect 184 -1967 185 -1965
rect 184 -1973 185 -1971
rect 191 -1967 192 -1965
rect 191 -1973 192 -1971
rect 201 -1967 202 -1965
rect 201 -1973 202 -1971
rect 205 -1967 206 -1965
rect 208 -1967 209 -1965
rect 208 -1973 209 -1971
rect 212 -1967 213 -1965
rect 212 -1973 213 -1971
rect 215 -1973 216 -1971
rect 219 -1967 220 -1965
rect 222 -1967 223 -1965
rect 219 -1973 220 -1971
rect 226 -1967 227 -1965
rect 226 -1973 227 -1971
rect 233 -1967 234 -1965
rect 233 -1973 234 -1971
rect 240 -1967 241 -1965
rect 240 -1973 241 -1971
rect 247 -1967 248 -1965
rect 247 -1973 248 -1971
rect 254 -1967 255 -1965
rect 254 -1973 255 -1971
rect 261 -1967 262 -1965
rect 261 -1973 262 -1971
rect 268 -1967 269 -1965
rect 271 -1967 272 -1965
rect 268 -1973 269 -1971
rect 275 -1967 276 -1965
rect 275 -1973 276 -1971
rect 282 -1967 283 -1965
rect 282 -1973 283 -1971
rect 289 -1967 290 -1965
rect 289 -1973 290 -1971
rect 296 -1967 297 -1965
rect 296 -1973 297 -1971
rect 303 -1967 304 -1965
rect 303 -1973 304 -1971
rect 310 -1967 311 -1965
rect 313 -1973 314 -1971
rect 317 -1967 318 -1965
rect 317 -1973 318 -1971
rect 324 -1967 325 -1965
rect 324 -1973 325 -1971
rect 331 -1967 332 -1965
rect 331 -1973 332 -1971
rect 338 -1967 339 -1965
rect 338 -1973 339 -1971
rect 345 -1967 346 -1965
rect 348 -1967 349 -1965
rect 345 -1973 346 -1971
rect 348 -1973 349 -1971
rect 352 -1967 353 -1965
rect 355 -1967 356 -1965
rect 359 -1967 360 -1965
rect 359 -1973 360 -1971
rect 366 -1967 367 -1965
rect 369 -1967 370 -1965
rect 366 -1973 367 -1971
rect 369 -1973 370 -1971
rect 373 -1967 374 -1965
rect 373 -1973 374 -1971
rect 380 -1967 381 -1965
rect 380 -1973 381 -1971
rect 387 -1973 388 -1971
rect 394 -1967 395 -1965
rect 397 -1967 398 -1965
rect 397 -1973 398 -1971
rect 401 -1967 402 -1965
rect 401 -1973 402 -1971
rect 408 -1967 409 -1965
rect 408 -1973 409 -1971
rect 418 -1967 419 -1965
rect 415 -1973 416 -1971
rect 418 -1973 419 -1971
rect 422 -1967 423 -1965
rect 429 -1967 430 -1965
rect 432 -1967 433 -1965
rect 429 -1973 430 -1971
rect 432 -1973 433 -1971
rect 436 -1967 437 -1965
rect 436 -1973 437 -1971
rect 443 -1967 444 -1965
rect 443 -1973 444 -1971
rect 450 -1967 451 -1965
rect 450 -1973 451 -1971
rect 460 -1967 461 -1965
rect 457 -1973 458 -1971
rect 464 -1973 465 -1971
rect 471 -1967 472 -1965
rect 471 -1973 472 -1971
rect 478 -1967 479 -1965
rect 481 -1967 482 -1965
rect 481 -1973 482 -1971
rect 485 -1967 486 -1965
rect 485 -1973 486 -1971
rect 492 -1967 493 -1965
rect 492 -1973 493 -1971
rect 499 -1967 500 -1965
rect 499 -1973 500 -1971
rect 506 -1967 507 -1965
rect 506 -1973 507 -1971
rect 513 -1967 514 -1965
rect 513 -1973 514 -1971
rect 520 -1967 521 -1965
rect 520 -1973 521 -1971
rect 527 -1967 528 -1965
rect 527 -1973 528 -1971
rect 534 -1967 535 -1965
rect 534 -1973 535 -1971
rect 541 -1967 542 -1965
rect 541 -1973 542 -1971
rect 548 -1973 549 -1971
rect 551 -1973 552 -1971
rect 555 -1967 556 -1965
rect 555 -1973 556 -1971
rect 562 -1967 563 -1965
rect 562 -1973 563 -1971
rect 569 -1967 570 -1965
rect 569 -1973 570 -1971
rect 576 -1967 577 -1965
rect 576 -1973 577 -1971
rect 583 -1967 584 -1965
rect 583 -1973 584 -1971
rect 590 -1967 591 -1965
rect 590 -1973 591 -1971
rect 597 -1967 598 -1965
rect 597 -1973 598 -1971
rect 604 -1967 605 -1965
rect 604 -1973 605 -1971
rect 611 -1967 612 -1965
rect 611 -1973 612 -1971
rect 618 -1967 619 -1965
rect 618 -1973 619 -1971
rect 625 -1967 626 -1965
rect 625 -1973 626 -1971
rect 632 -1967 633 -1965
rect 632 -1973 633 -1971
rect 639 -1973 640 -1971
rect 642 -1973 643 -1971
rect 646 -1967 647 -1965
rect 646 -1973 647 -1971
rect 653 -1967 654 -1965
rect 653 -1973 654 -1971
rect 660 -1967 661 -1965
rect 660 -1973 661 -1971
rect 667 -1967 668 -1965
rect 667 -1973 668 -1971
rect 674 -1967 675 -1965
rect 674 -1973 675 -1971
rect 681 -1967 682 -1965
rect 681 -1973 682 -1971
rect 688 -1967 689 -1965
rect 688 -1973 689 -1971
rect 695 -1967 696 -1965
rect 695 -1973 696 -1971
rect 702 -1967 703 -1965
rect 702 -1973 703 -1971
rect 709 -1967 710 -1965
rect 709 -1973 710 -1971
rect 716 -1967 717 -1965
rect 716 -1973 717 -1971
rect 723 -1967 724 -1965
rect 723 -1973 724 -1971
rect 730 -1967 731 -1965
rect 730 -1973 731 -1971
rect 9 -2028 10 -2026
rect 9 -2034 10 -2032
rect 16 -2028 17 -2026
rect 16 -2034 17 -2032
rect 23 -2028 24 -2026
rect 30 -2028 31 -2026
rect 30 -2034 31 -2032
rect 37 -2028 38 -2026
rect 37 -2034 38 -2032
rect 44 -2028 45 -2026
rect 44 -2034 45 -2032
rect 51 -2028 52 -2026
rect 54 -2028 55 -2026
rect 51 -2034 52 -2032
rect 58 -2028 59 -2026
rect 58 -2034 59 -2032
rect 65 -2028 66 -2026
rect 68 -2028 69 -2026
rect 65 -2034 66 -2032
rect 72 -2028 73 -2026
rect 72 -2034 73 -2032
rect 79 -2028 80 -2026
rect 79 -2034 80 -2032
rect 89 -2028 90 -2026
rect 86 -2034 87 -2032
rect 89 -2034 90 -2032
rect 96 -2034 97 -2032
rect 100 -2028 101 -2026
rect 103 -2028 104 -2026
rect 107 -2028 108 -2026
rect 107 -2034 108 -2032
rect 117 -2028 118 -2026
rect 114 -2034 115 -2032
rect 117 -2034 118 -2032
rect 121 -2028 122 -2026
rect 121 -2034 122 -2032
rect 128 -2028 129 -2026
rect 131 -2028 132 -2026
rect 128 -2034 129 -2032
rect 135 -2028 136 -2026
rect 135 -2034 136 -2032
rect 142 -2028 143 -2026
rect 142 -2034 143 -2032
rect 149 -2028 150 -2026
rect 149 -2034 150 -2032
rect 156 -2028 157 -2026
rect 156 -2034 157 -2032
rect 163 -2028 164 -2026
rect 163 -2034 164 -2032
rect 170 -2028 171 -2026
rect 170 -2034 171 -2032
rect 177 -2028 178 -2026
rect 177 -2034 178 -2032
rect 184 -2028 185 -2026
rect 184 -2034 185 -2032
rect 191 -2034 192 -2032
rect 198 -2034 199 -2032
rect 201 -2034 202 -2032
rect 205 -2028 206 -2026
rect 205 -2034 206 -2032
rect 212 -2034 213 -2032
rect 215 -2034 216 -2032
rect 219 -2028 220 -2026
rect 219 -2034 220 -2032
rect 222 -2034 223 -2032
rect 226 -2028 227 -2026
rect 226 -2034 227 -2032
rect 233 -2028 234 -2026
rect 233 -2034 234 -2032
rect 240 -2028 241 -2026
rect 240 -2034 241 -2032
rect 247 -2028 248 -2026
rect 254 -2034 255 -2032
rect 257 -2034 258 -2032
rect 261 -2028 262 -2026
rect 261 -2034 262 -2032
rect 268 -2028 269 -2026
rect 268 -2034 269 -2032
rect 275 -2028 276 -2026
rect 275 -2034 276 -2032
rect 282 -2028 283 -2026
rect 285 -2028 286 -2026
rect 282 -2034 283 -2032
rect 289 -2028 290 -2026
rect 289 -2034 290 -2032
rect 296 -2028 297 -2026
rect 296 -2034 297 -2032
rect 303 -2028 304 -2026
rect 306 -2028 307 -2026
rect 303 -2034 304 -2032
rect 310 -2028 311 -2026
rect 310 -2034 311 -2032
rect 317 -2028 318 -2026
rect 317 -2034 318 -2032
rect 324 -2028 325 -2026
rect 324 -2034 325 -2032
rect 331 -2028 332 -2026
rect 331 -2034 332 -2032
rect 338 -2028 339 -2026
rect 338 -2034 339 -2032
rect 345 -2028 346 -2026
rect 345 -2034 346 -2032
rect 352 -2028 353 -2026
rect 352 -2034 353 -2032
rect 359 -2028 360 -2026
rect 359 -2034 360 -2032
rect 366 -2028 367 -2026
rect 366 -2034 367 -2032
rect 373 -2028 374 -2026
rect 373 -2034 374 -2032
rect 380 -2034 381 -2032
rect 387 -2028 388 -2026
rect 387 -2034 388 -2032
rect 394 -2028 395 -2026
rect 394 -2034 395 -2032
rect 404 -2028 405 -2026
rect 401 -2034 402 -2032
rect 404 -2034 405 -2032
rect 408 -2028 409 -2026
rect 408 -2034 409 -2032
rect 415 -2028 416 -2026
rect 418 -2034 419 -2032
rect 422 -2028 423 -2026
rect 422 -2034 423 -2032
rect 429 -2028 430 -2026
rect 429 -2034 430 -2032
rect 436 -2028 437 -2026
rect 439 -2028 440 -2026
rect 436 -2034 437 -2032
rect 443 -2028 444 -2026
rect 443 -2034 444 -2032
rect 450 -2028 451 -2026
rect 450 -2034 451 -2032
rect 457 -2028 458 -2026
rect 457 -2034 458 -2032
rect 464 -2028 465 -2026
rect 464 -2034 465 -2032
rect 474 -2028 475 -2026
rect 471 -2034 472 -2032
rect 474 -2034 475 -2032
rect 478 -2028 479 -2026
rect 478 -2034 479 -2032
rect 488 -2028 489 -2026
rect 492 -2028 493 -2026
rect 492 -2034 493 -2032
rect 499 -2028 500 -2026
rect 499 -2034 500 -2032
rect 506 -2028 507 -2026
rect 506 -2034 507 -2032
rect 513 -2028 514 -2026
rect 513 -2034 514 -2032
rect 520 -2028 521 -2026
rect 527 -2028 528 -2026
rect 527 -2034 528 -2032
rect 534 -2028 535 -2026
rect 534 -2034 535 -2032
rect 541 -2028 542 -2026
rect 541 -2034 542 -2032
rect 551 -2028 552 -2026
rect 548 -2034 549 -2032
rect 555 -2028 556 -2026
rect 555 -2034 556 -2032
rect 562 -2028 563 -2026
rect 562 -2034 563 -2032
rect 569 -2028 570 -2026
rect 569 -2034 570 -2032
rect 576 -2028 577 -2026
rect 576 -2034 577 -2032
rect 583 -2028 584 -2026
rect 583 -2034 584 -2032
rect 590 -2028 591 -2026
rect 590 -2034 591 -2032
rect 597 -2028 598 -2026
rect 597 -2034 598 -2032
rect 604 -2028 605 -2026
rect 604 -2034 605 -2032
rect 611 -2028 612 -2026
rect 611 -2034 612 -2032
rect 618 -2028 619 -2026
rect 618 -2034 619 -2032
rect 625 -2028 626 -2026
rect 625 -2034 626 -2032
rect 632 -2028 633 -2026
rect 635 -2028 636 -2026
rect 632 -2034 633 -2032
rect 635 -2034 636 -2032
rect 642 -2028 643 -2026
rect 639 -2034 640 -2032
rect 642 -2034 643 -2032
rect 646 -2028 647 -2026
rect 649 -2028 650 -2026
rect 653 -2028 654 -2026
rect 653 -2034 654 -2032
rect 660 -2028 661 -2026
rect 660 -2034 661 -2032
rect 670 -2034 671 -2032
rect 695 -2028 696 -2026
rect 695 -2034 696 -2032
rect 16 -2093 17 -2091
rect 16 -2099 17 -2097
rect 23 -2099 24 -2097
rect 33 -2093 34 -2091
rect 37 -2093 38 -2091
rect 37 -2099 38 -2097
rect 44 -2093 45 -2091
rect 44 -2099 45 -2097
rect 51 -2093 52 -2091
rect 51 -2099 52 -2097
rect 58 -2093 59 -2091
rect 58 -2099 59 -2097
rect 65 -2093 66 -2091
rect 65 -2099 66 -2097
rect 75 -2093 76 -2091
rect 72 -2099 73 -2097
rect 75 -2099 76 -2097
rect 79 -2093 80 -2091
rect 79 -2099 80 -2097
rect 86 -2093 87 -2091
rect 86 -2099 87 -2097
rect 96 -2093 97 -2091
rect 100 -2093 101 -2091
rect 100 -2099 101 -2097
rect 107 -2093 108 -2091
rect 107 -2099 108 -2097
rect 114 -2093 115 -2091
rect 117 -2093 118 -2091
rect 117 -2099 118 -2097
rect 121 -2093 122 -2091
rect 121 -2099 122 -2097
rect 128 -2093 129 -2091
rect 128 -2099 129 -2097
rect 135 -2093 136 -2091
rect 135 -2099 136 -2097
rect 142 -2093 143 -2091
rect 142 -2099 143 -2097
rect 149 -2093 150 -2091
rect 149 -2099 150 -2097
rect 156 -2093 157 -2091
rect 159 -2093 160 -2091
rect 163 -2093 164 -2091
rect 163 -2099 164 -2097
rect 170 -2093 171 -2091
rect 170 -2099 171 -2097
rect 177 -2093 178 -2091
rect 177 -2099 178 -2097
rect 184 -2099 185 -2097
rect 187 -2099 188 -2097
rect 191 -2093 192 -2091
rect 194 -2093 195 -2091
rect 198 -2093 199 -2091
rect 198 -2099 199 -2097
rect 205 -2099 206 -2097
rect 208 -2099 209 -2097
rect 212 -2093 213 -2091
rect 212 -2099 213 -2097
rect 219 -2093 220 -2091
rect 222 -2093 223 -2091
rect 226 -2093 227 -2091
rect 226 -2099 227 -2097
rect 236 -2093 237 -2091
rect 233 -2099 234 -2097
rect 240 -2093 241 -2091
rect 240 -2099 241 -2097
rect 247 -2093 248 -2091
rect 247 -2099 248 -2097
rect 254 -2093 255 -2091
rect 254 -2099 255 -2097
rect 261 -2093 262 -2091
rect 261 -2099 262 -2097
rect 268 -2093 269 -2091
rect 268 -2099 269 -2097
rect 275 -2093 276 -2091
rect 275 -2099 276 -2097
rect 282 -2093 283 -2091
rect 282 -2099 283 -2097
rect 289 -2093 290 -2091
rect 289 -2099 290 -2097
rect 296 -2093 297 -2091
rect 296 -2099 297 -2097
rect 303 -2093 304 -2091
rect 306 -2093 307 -2091
rect 306 -2099 307 -2097
rect 313 -2093 314 -2091
rect 310 -2099 311 -2097
rect 317 -2093 318 -2091
rect 320 -2093 321 -2091
rect 317 -2099 318 -2097
rect 320 -2099 321 -2097
rect 324 -2093 325 -2091
rect 327 -2093 328 -2091
rect 331 -2093 332 -2091
rect 331 -2099 332 -2097
rect 338 -2093 339 -2091
rect 338 -2099 339 -2097
rect 345 -2093 346 -2091
rect 345 -2099 346 -2097
rect 352 -2093 353 -2091
rect 359 -2093 360 -2091
rect 359 -2099 360 -2097
rect 366 -2093 367 -2091
rect 369 -2093 370 -2091
rect 369 -2099 370 -2097
rect 373 -2093 374 -2091
rect 373 -2099 374 -2097
rect 380 -2093 381 -2091
rect 383 -2093 384 -2091
rect 383 -2099 384 -2097
rect 387 -2093 388 -2091
rect 387 -2099 388 -2097
rect 394 -2093 395 -2091
rect 394 -2099 395 -2097
rect 401 -2093 402 -2091
rect 404 -2093 405 -2091
rect 408 -2093 409 -2091
rect 415 -2093 416 -2091
rect 418 -2093 419 -2091
rect 425 -2093 426 -2091
rect 422 -2099 423 -2097
rect 429 -2093 430 -2091
rect 429 -2099 430 -2097
rect 436 -2093 437 -2091
rect 436 -2099 437 -2097
rect 443 -2093 444 -2091
rect 443 -2099 444 -2097
rect 450 -2093 451 -2091
rect 450 -2099 451 -2097
rect 457 -2093 458 -2091
rect 457 -2099 458 -2097
rect 464 -2093 465 -2091
rect 464 -2099 465 -2097
rect 471 -2093 472 -2091
rect 471 -2099 472 -2097
rect 478 -2093 479 -2091
rect 481 -2093 482 -2091
rect 485 -2093 486 -2091
rect 485 -2099 486 -2097
rect 492 -2093 493 -2091
rect 492 -2099 493 -2097
rect 499 -2093 500 -2091
rect 502 -2099 503 -2097
rect 506 -2093 507 -2091
rect 506 -2099 507 -2097
rect 513 -2093 514 -2091
rect 513 -2099 514 -2097
rect 520 -2093 521 -2091
rect 520 -2099 521 -2097
rect 527 -2093 528 -2091
rect 527 -2099 528 -2097
rect 534 -2093 535 -2091
rect 534 -2099 535 -2097
rect 541 -2093 542 -2091
rect 541 -2099 542 -2097
rect 548 -2093 549 -2091
rect 548 -2099 549 -2097
rect 555 -2093 556 -2091
rect 558 -2099 559 -2097
rect 562 -2093 563 -2091
rect 562 -2099 563 -2097
rect 569 -2093 570 -2091
rect 569 -2099 570 -2097
rect 576 -2093 577 -2091
rect 576 -2099 577 -2097
rect 583 -2093 584 -2091
rect 583 -2099 584 -2097
rect 590 -2093 591 -2091
rect 590 -2099 591 -2097
rect 604 -2093 605 -2091
rect 604 -2099 605 -2097
rect 611 -2093 612 -2091
rect 611 -2099 612 -2097
rect 618 -2099 619 -2097
rect 621 -2099 622 -2097
rect 642 -2093 643 -2091
rect 642 -2099 643 -2097
rect 646 -2093 647 -2091
rect 646 -2099 647 -2097
rect 674 -2093 675 -2091
rect 674 -2099 675 -2097
rect 688 -2093 689 -2091
rect 688 -2099 689 -2097
rect 26 -2150 27 -2148
rect 33 -2150 34 -2148
rect 37 -2150 38 -2148
rect 37 -2156 38 -2154
rect 44 -2150 45 -2148
rect 44 -2156 45 -2154
rect 51 -2150 52 -2148
rect 51 -2156 52 -2154
rect 58 -2150 59 -2148
rect 58 -2156 59 -2154
rect 65 -2150 66 -2148
rect 65 -2156 66 -2154
rect 72 -2156 73 -2154
rect 79 -2150 80 -2148
rect 86 -2150 87 -2148
rect 86 -2156 87 -2154
rect 93 -2156 94 -2154
rect 96 -2156 97 -2154
rect 100 -2150 101 -2148
rect 100 -2156 101 -2154
rect 107 -2150 108 -2148
rect 107 -2156 108 -2154
rect 117 -2150 118 -2148
rect 121 -2156 122 -2154
rect 128 -2156 129 -2154
rect 131 -2156 132 -2154
rect 135 -2150 136 -2148
rect 135 -2156 136 -2154
rect 142 -2150 143 -2148
rect 142 -2156 143 -2154
rect 152 -2150 153 -2148
rect 156 -2150 157 -2148
rect 156 -2156 157 -2154
rect 163 -2150 164 -2148
rect 163 -2156 164 -2154
rect 170 -2150 171 -2148
rect 170 -2156 171 -2154
rect 177 -2150 178 -2148
rect 177 -2156 178 -2154
rect 180 -2156 181 -2154
rect 184 -2156 185 -2154
rect 187 -2156 188 -2154
rect 191 -2150 192 -2148
rect 191 -2156 192 -2154
rect 198 -2150 199 -2148
rect 198 -2156 199 -2154
rect 205 -2150 206 -2148
rect 205 -2156 206 -2154
rect 215 -2150 216 -2148
rect 212 -2156 213 -2154
rect 222 -2150 223 -2148
rect 219 -2156 220 -2154
rect 226 -2150 227 -2148
rect 226 -2156 227 -2154
rect 233 -2150 234 -2148
rect 233 -2156 234 -2154
rect 240 -2150 241 -2148
rect 240 -2156 241 -2154
rect 247 -2150 248 -2148
rect 247 -2156 248 -2154
rect 254 -2150 255 -2148
rect 261 -2150 262 -2148
rect 264 -2150 265 -2148
rect 268 -2150 269 -2148
rect 268 -2156 269 -2154
rect 275 -2150 276 -2148
rect 275 -2156 276 -2154
rect 282 -2156 283 -2154
rect 289 -2150 290 -2148
rect 292 -2150 293 -2148
rect 292 -2156 293 -2154
rect 296 -2150 297 -2148
rect 296 -2156 297 -2154
rect 303 -2150 304 -2148
rect 306 -2150 307 -2148
rect 303 -2156 304 -2154
rect 310 -2150 311 -2148
rect 310 -2156 311 -2154
rect 317 -2156 318 -2154
rect 324 -2150 325 -2148
rect 324 -2156 325 -2154
rect 334 -2150 335 -2148
rect 334 -2156 335 -2154
rect 338 -2150 339 -2148
rect 338 -2156 339 -2154
rect 345 -2150 346 -2148
rect 345 -2156 346 -2154
rect 352 -2150 353 -2148
rect 352 -2156 353 -2154
rect 359 -2156 360 -2154
rect 362 -2156 363 -2154
rect 366 -2150 367 -2148
rect 366 -2156 367 -2154
rect 373 -2150 374 -2148
rect 380 -2150 381 -2148
rect 380 -2156 381 -2154
rect 387 -2150 388 -2148
rect 387 -2156 388 -2154
rect 394 -2150 395 -2148
rect 394 -2156 395 -2154
rect 401 -2150 402 -2148
rect 401 -2156 402 -2154
rect 408 -2150 409 -2148
rect 408 -2156 409 -2154
rect 415 -2156 416 -2154
rect 422 -2150 423 -2148
rect 422 -2156 423 -2154
rect 429 -2150 430 -2148
rect 429 -2156 430 -2154
rect 436 -2150 437 -2148
rect 436 -2156 437 -2154
rect 443 -2150 444 -2148
rect 443 -2156 444 -2154
rect 450 -2150 451 -2148
rect 450 -2156 451 -2154
rect 457 -2150 458 -2148
rect 457 -2156 458 -2154
rect 467 -2156 468 -2154
rect 471 -2150 472 -2148
rect 471 -2156 472 -2154
rect 478 -2150 479 -2148
rect 478 -2156 479 -2154
rect 485 -2150 486 -2148
rect 485 -2156 486 -2154
rect 492 -2150 493 -2148
rect 492 -2156 493 -2154
rect 499 -2156 500 -2154
rect 509 -2150 510 -2148
rect 509 -2156 510 -2154
rect 513 -2150 514 -2148
rect 513 -2156 514 -2154
rect 523 -2150 524 -2148
rect 530 -2150 531 -2148
rect 534 -2150 535 -2148
rect 534 -2156 535 -2154
rect 541 -2150 542 -2148
rect 541 -2156 542 -2154
rect 548 -2150 549 -2148
rect 548 -2156 549 -2154
rect 555 -2150 556 -2148
rect 555 -2156 556 -2154
rect 562 -2150 563 -2148
rect 562 -2156 563 -2154
rect 569 -2150 570 -2148
rect 569 -2156 570 -2154
rect 590 -2150 591 -2148
rect 590 -2156 591 -2154
rect 597 -2150 598 -2148
rect 597 -2156 598 -2154
rect 611 -2150 612 -2148
rect 611 -2156 612 -2154
rect 9 -2197 10 -2195
rect 9 -2203 10 -2201
rect 19 -2197 20 -2195
rect 23 -2203 24 -2201
rect 40 -2197 41 -2195
rect 44 -2203 45 -2201
rect 51 -2197 52 -2195
rect 51 -2203 52 -2201
rect 58 -2197 59 -2195
rect 58 -2203 59 -2201
rect 65 -2197 66 -2195
rect 65 -2203 66 -2201
rect 72 -2197 73 -2195
rect 72 -2203 73 -2201
rect 79 -2197 80 -2195
rect 79 -2203 80 -2201
rect 86 -2197 87 -2195
rect 86 -2203 87 -2201
rect 93 -2197 94 -2195
rect 93 -2203 94 -2201
rect 100 -2197 101 -2195
rect 100 -2203 101 -2201
rect 107 -2197 108 -2195
rect 107 -2203 108 -2201
rect 114 -2203 115 -2201
rect 121 -2197 122 -2195
rect 121 -2203 122 -2201
rect 128 -2197 129 -2195
rect 131 -2197 132 -2195
rect 128 -2203 129 -2201
rect 135 -2197 136 -2195
rect 138 -2197 139 -2195
rect 145 -2203 146 -2201
rect 149 -2197 150 -2195
rect 149 -2203 150 -2201
rect 156 -2197 157 -2195
rect 156 -2203 157 -2201
rect 163 -2197 164 -2195
rect 163 -2203 164 -2201
rect 170 -2197 171 -2195
rect 170 -2203 171 -2201
rect 177 -2197 178 -2195
rect 177 -2203 178 -2201
rect 187 -2197 188 -2195
rect 191 -2197 192 -2195
rect 191 -2203 192 -2201
rect 198 -2197 199 -2195
rect 201 -2203 202 -2201
rect 208 -2197 209 -2195
rect 205 -2203 206 -2201
rect 212 -2197 213 -2195
rect 215 -2197 216 -2195
rect 219 -2197 220 -2195
rect 219 -2203 220 -2201
rect 226 -2197 227 -2195
rect 226 -2203 227 -2201
rect 233 -2197 234 -2195
rect 247 -2197 248 -2195
rect 247 -2203 248 -2201
rect 257 -2197 258 -2195
rect 254 -2203 255 -2201
rect 261 -2197 262 -2195
rect 261 -2203 262 -2201
rect 268 -2197 269 -2195
rect 268 -2203 269 -2201
rect 278 -2197 279 -2195
rect 285 -2197 286 -2195
rect 289 -2197 290 -2195
rect 289 -2203 290 -2201
rect 296 -2197 297 -2195
rect 299 -2203 300 -2201
rect 303 -2197 304 -2195
rect 303 -2203 304 -2201
rect 317 -2197 318 -2195
rect 317 -2203 318 -2201
rect 324 -2197 325 -2195
rect 324 -2203 325 -2201
rect 331 -2197 332 -2195
rect 331 -2203 332 -2201
rect 345 -2197 346 -2195
rect 348 -2197 349 -2195
rect 345 -2203 346 -2201
rect 352 -2197 353 -2195
rect 352 -2203 353 -2201
rect 359 -2203 360 -2201
rect 362 -2203 363 -2201
rect 366 -2203 367 -2201
rect 373 -2197 374 -2195
rect 380 -2197 381 -2195
rect 380 -2203 381 -2201
rect 387 -2197 388 -2195
rect 387 -2203 388 -2201
rect 394 -2197 395 -2195
rect 394 -2203 395 -2201
rect 401 -2197 402 -2195
rect 401 -2203 402 -2201
rect 408 -2197 409 -2195
rect 408 -2203 409 -2201
rect 415 -2197 416 -2195
rect 418 -2203 419 -2201
rect 425 -2197 426 -2195
rect 422 -2203 423 -2201
rect 429 -2197 430 -2195
rect 429 -2203 430 -2201
rect 436 -2197 437 -2195
rect 436 -2203 437 -2201
rect 443 -2197 444 -2195
rect 443 -2203 444 -2201
rect 453 -2197 454 -2195
rect 457 -2197 458 -2195
rect 457 -2203 458 -2201
rect 464 -2197 465 -2195
rect 464 -2203 465 -2201
rect 481 -2197 482 -2195
rect 492 -2197 493 -2195
rect 492 -2203 493 -2201
rect 499 -2197 500 -2195
rect 520 -2197 521 -2195
rect 520 -2203 521 -2201
rect 534 -2197 535 -2195
rect 534 -2203 535 -2201
rect 548 -2203 549 -2201
rect 555 -2197 556 -2195
rect 555 -2203 556 -2201
rect 600 -2197 601 -2195
rect 600 -2203 601 -2201
rect 604 -2197 605 -2195
rect 604 -2203 605 -2201
rect 611 -2197 612 -2195
rect 611 -2203 612 -2201
rect 16 -2226 17 -2224
rect 26 -2226 27 -2224
rect 44 -2226 45 -2224
rect 51 -2226 52 -2224
rect 58 -2226 59 -2224
rect 58 -2232 59 -2230
rect 75 -2232 76 -2230
rect 82 -2226 83 -2224
rect 93 -2232 94 -2230
rect 103 -2226 104 -2224
rect 107 -2226 108 -2224
rect 107 -2232 108 -2230
rect 114 -2226 115 -2224
rect 114 -2232 115 -2230
rect 131 -2232 132 -2230
rect 149 -2226 150 -2224
rect 149 -2232 150 -2230
rect 163 -2232 164 -2230
rect 173 -2232 174 -2230
rect 177 -2226 178 -2224
rect 187 -2226 188 -2224
rect 191 -2226 192 -2224
rect 201 -2232 202 -2230
rect 205 -2226 206 -2224
rect 208 -2226 209 -2224
rect 212 -2226 213 -2224
rect 219 -2232 220 -2230
rect 226 -2226 227 -2224
rect 226 -2232 227 -2230
rect 240 -2226 241 -2224
rect 240 -2232 241 -2230
rect 247 -2226 248 -2224
rect 247 -2232 248 -2230
rect 254 -2226 255 -2224
rect 254 -2232 255 -2230
rect 268 -2226 269 -2224
rect 268 -2232 269 -2230
rect 275 -2226 276 -2224
rect 275 -2232 276 -2230
rect 282 -2226 283 -2224
rect 282 -2232 283 -2230
rect 289 -2226 290 -2224
rect 289 -2232 290 -2230
rect 303 -2232 304 -2230
rect 310 -2232 311 -2230
rect 313 -2232 314 -2230
rect 327 -2226 328 -2224
rect 327 -2232 328 -2230
rect 331 -2226 332 -2224
rect 331 -2232 332 -2230
rect 341 -2226 342 -2224
rect 348 -2226 349 -2224
rect 355 -2232 356 -2230
rect 373 -2226 374 -2224
rect 373 -2232 374 -2230
rect 383 -2232 384 -2230
rect 390 -2232 391 -2230
rect 408 -2226 409 -2224
rect 408 -2232 409 -2230
rect 429 -2232 430 -2230
rect 450 -2226 451 -2224
rect 450 -2232 451 -2230
rect 474 -2232 475 -2230
rect 485 -2232 486 -2230
rect 506 -2226 507 -2224
rect 506 -2232 507 -2230
rect 534 -2226 535 -2224
rect 537 -2226 538 -2224
rect 611 -2226 612 -2224
<< metal1 >>
rect 131 0 157 1
rect 163 0 188 1
rect 191 0 234 1
rect 261 0 283 1
rect 177 -2 213 -1
rect 215 -2 248 -1
rect 268 -2 279 -1
rect 226 -4 258 -3
rect 86 -15 164 -14
rect 170 -15 220 -14
rect 240 -15 262 -14
rect 268 -15 346 -14
rect 369 -15 402 -14
rect 93 -17 101 -16
rect 107 -17 111 -16
rect 142 -17 227 -16
rect 247 -17 290 -16
rect 327 -17 332 -16
rect 376 -17 381 -16
rect 110 -19 255 -18
rect 257 -19 388 -18
rect 138 -21 143 -20
rect 149 -21 167 -20
rect 170 -21 178 -20
rect 180 -21 234 -20
rect 243 -21 248 -20
rect 275 -21 419 -20
rect 156 -23 178 -22
rect 184 -23 213 -22
rect 215 -23 297 -22
rect 117 -25 157 -24
rect 191 -25 353 -24
rect 128 -27 192 -26
rect 198 -27 304 -26
rect 198 -29 209 -28
rect 222 -29 262 -28
rect 282 -29 360 -28
rect 205 -31 269 -30
rect 282 -31 318 -30
rect 65 -42 94 -41
rect 100 -42 185 -41
rect 212 -42 360 -41
rect 72 -44 129 -43
rect 149 -44 181 -43
rect 184 -44 199 -43
rect 226 -44 374 -43
rect 75 -46 150 -45
rect 156 -46 199 -45
rect 229 -46 262 -45
rect 275 -46 279 -45
rect 282 -46 409 -45
rect 79 -48 216 -47
rect 233 -48 314 -47
rect 324 -48 388 -47
rect 86 -50 223 -49
rect 233 -50 241 -49
rect 261 -50 269 -49
rect 275 -50 318 -49
rect 44 -52 87 -51
rect 114 -52 157 -51
rect 163 -52 213 -51
rect 240 -52 248 -51
rect 278 -52 318 -51
rect 107 -54 115 -53
rect 117 -54 174 -53
rect 191 -54 248 -53
rect 282 -54 381 -53
rect 121 -56 178 -55
rect 205 -56 381 -55
rect 121 -58 136 -57
rect 170 -58 360 -57
rect 131 -60 388 -59
rect 135 -62 143 -61
rect 170 -62 402 -61
rect 285 -64 346 -63
rect 289 -66 311 -65
rect 331 -66 402 -65
rect 219 -68 290 -67
rect 296 -68 325 -67
rect 338 -68 346 -67
rect 219 -70 367 -69
rect 254 -72 297 -71
rect 338 -72 395 -71
rect 51 -74 255 -73
rect 257 -74 332 -73
rect 352 -74 395 -73
rect 44 -85 101 -84
rect 121 -85 136 -84
rect 159 -85 192 -84
rect 194 -85 227 -84
rect 250 -85 402 -84
rect 51 -87 157 -86
rect 163 -87 171 -86
rect 201 -87 248 -86
rect 254 -87 304 -86
rect 331 -87 384 -86
rect 394 -87 444 -86
rect 58 -89 146 -88
rect 205 -89 241 -88
rect 257 -89 374 -88
rect 401 -89 454 -88
rect 65 -91 115 -90
rect 128 -91 395 -90
rect 65 -93 80 -92
rect 86 -93 108 -92
rect 131 -93 290 -92
rect 317 -93 332 -92
rect 352 -93 409 -92
rect 93 -95 125 -94
rect 142 -95 164 -94
rect 212 -95 262 -94
rect 271 -95 388 -94
rect 408 -95 433 -94
rect 107 -97 248 -96
rect 275 -97 283 -96
rect 289 -97 360 -96
rect 366 -97 416 -96
rect 96 -99 360 -98
rect 149 -101 374 -100
rect 149 -103 185 -102
rect 212 -103 220 -102
rect 222 -103 423 -102
rect 177 -105 262 -104
rect 278 -105 381 -104
rect 184 -107 192 -106
rect 215 -107 325 -106
rect 338 -107 388 -106
rect 79 -109 216 -108
rect 233 -109 255 -108
rect 271 -109 339 -108
rect 345 -109 353 -108
rect 198 -111 346 -110
rect 240 -113 430 -112
rect 278 -115 304 -114
rect 310 -115 325 -114
rect 296 -117 318 -116
rect 296 -119 367 -118
rect 37 -130 150 -129
rect 156 -130 199 -129
rect 215 -130 430 -129
rect 436 -130 482 -129
rect 44 -132 94 -131
rect 110 -132 115 -131
rect 128 -132 206 -131
rect 219 -132 223 -131
rect 226 -132 251 -131
rect 254 -132 269 -131
rect 275 -132 451 -131
rect 51 -134 167 -133
rect 170 -134 430 -133
rect 58 -136 143 -135
rect 145 -136 227 -135
rect 233 -136 237 -135
rect 247 -136 339 -135
rect 359 -136 367 -135
rect 380 -136 472 -135
rect 58 -138 167 -137
rect 170 -138 192 -137
rect 236 -138 416 -137
rect 72 -140 122 -139
rect 131 -140 423 -139
rect 79 -142 94 -141
rect 177 -142 199 -141
rect 254 -142 465 -141
rect 79 -144 122 -143
rect 184 -144 248 -143
rect 261 -144 286 -143
rect 289 -144 381 -143
rect 387 -144 486 -143
rect 89 -146 101 -145
rect 103 -146 178 -145
rect 191 -146 325 -145
rect 352 -146 360 -145
rect 401 -146 458 -145
rect 100 -148 108 -147
rect 117 -148 325 -147
rect 345 -148 353 -147
rect 415 -148 444 -147
rect 138 -150 185 -149
rect 208 -150 402 -149
rect 86 -152 139 -151
rect 282 -152 339 -151
rect 296 -154 314 -153
rect 317 -154 493 -153
rect 296 -156 388 -155
rect 303 -158 346 -157
rect 306 -160 444 -159
rect 310 -162 409 -161
rect 317 -164 409 -163
rect 320 -166 395 -165
rect 373 -168 395 -167
rect 331 -170 374 -169
rect 331 -172 440 -171
rect 16 -183 90 -182
rect 114 -183 153 -182
rect 191 -183 286 -182
rect 292 -183 374 -182
rect 380 -183 556 -182
rect 583 -183 640 -182
rect 30 -185 223 -184
rect 226 -185 479 -184
rect 534 -185 549 -184
rect 37 -187 209 -186
rect 254 -187 335 -186
rect 380 -187 566 -186
rect 37 -189 80 -188
rect 86 -189 108 -188
rect 114 -189 342 -188
rect 387 -189 549 -188
rect 44 -191 146 -190
rect 191 -191 234 -190
rect 257 -191 269 -190
rect 275 -191 339 -190
rect 366 -191 388 -190
rect 464 -191 500 -190
rect 51 -193 290 -192
rect 296 -193 325 -192
rect 450 -193 465 -192
rect 471 -193 507 -192
rect 58 -195 528 -194
rect 58 -197 94 -196
rect 121 -197 248 -196
rect 261 -197 290 -196
rect 306 -197 486 -196
rect 65 -199 69 -198
rect 72 -199 153 -198
rect 156 -199 262 -198
rect 278 -199 430 -198
rect 443 -199 451 -198
rect 457 -199 472 -198
rect 79 -201 423 -200
rect 436 -201 444 -200
rect 89 -203 416 -202
rect 103 -205 430 -204
rect 121 -207 374 -206
rect 408 -207 458 -206
rect 124 -209 241 -208
rect 243 -209 269 -208
rect 282 -209 416 -208
rect 128 -211 185 -210
rect 187 -211 367 -210
rect 408 -211 521 -210
rect 82 -213 129 -212
rect 135 -213 244 -212
rect 317 -213 493 -212
rect 135 -215 164 -214
rect 170 -215 248 -214
rect 324 -215 514 -214
rect 142 -217 227 -216
rect 233 -217 346 -216
rect 401 -217 493 -216
rect 96 -219 402 -218
rect 142 -221 304 -220
rect 331 -221 486 -220
rect 170 -223 178 -222
rect 198 -223 216 -222
rect 310 -223 332 -222
rect 345 -223 395 -222
rect 156 -225 178 -224
rect 198 -225 353 -224
rect 359 -225 395 -224
rect 205 -227 220 -226
rect 359 -227 437 -226
rect 149 -229 220 -228
rect 16 -240 150 -239
rect 180 -240 248 -239
rect 285 -240 493 -239
rect 499 -240 577 -239
rect 586 -240 626 -239
rect 639 -240 661 -239
rect 30 -242 146 -241
rect 205 -242 220 -241
rect 240 -242 605 -241
rect 30 -244 199 -243
rect 205 -244 241 -243
rect 243 -244 276 -243
rect 278 -244 493 -243
rect 506 -244 563 -243
rect 44 -246 80 -245
rect 82 -246 479 -245
rect 481 -246 591 -245
rect 51 -248 528 -247
rect 534 -248 566 -247
rect 58 -250 94 -249
rect 103 -250 346 -249
rect 352 -250 486 -249
rect 513 -250 584 -249
rect 72 -252 136 -251
rect 156 -252 353 -251
rect 362 -252 402 -251
rect 408 -252 507 -251
rect 555 -252 598 -251
rect 86 -254 195 -253
rect 198 -254 360 -253
rect 366 -254 486 -253
rect 558 -254 619 -253
rect 93 -256 101 -255
rect 124 -256 136 -255
rect 156 -256 178 -255
rect 212 -256 227 -255
rect 247 -256 409 -255
rect 422 -256 528 -255
rect 100 -258 167 -257
rect 226 -258 258 -257
rect 268 -258 276 -257
rect 285 -258 633 -257
rect 254 -260 423 -259
rect 429 -260 535 -259
rect 268 -262 325 -261
rect 331 -262 500 -261
rect 233 -264 332 -263
rect 338 -264 514 -263
rect 289 -266 297 -265
rect 303 -266 346 -265
rect 380 -266 440 -265
rect 443 -266 521 -265
rect 114 -268 290 -267
rect 310 -268 402 -267
rect 415 -268 430 -267
rect 457 -268 612 -267
rect 114 -270 262 -269
rect 282 -270 444 -269
rect 457 -270 465 -269
rect 471 -270 570 -269
rect 128 -272 381 -271
rect 387 -272 556 -271
rect 107 -274 129 -273
rect 152 -274 262 -273
rect 299 -274 416 -273
rect 107 -276 192 -275
rect 222 -276 465 -275
rect 152 -278 164 -277
rect 170 -278 304 -277
rect 313 -278 542 -277
rect 40 -280 171 -279
rect 317 -280 325 -279
rect 366 -280 388 -279
rect 394 -280 549 -279
rect 215 -282 395 -281
rect 450 -282 542 -281
rect 215 -284 234 -283
rect 373 -284 472 -283
rect 163 -286 374 -285
rect 436 -286 451 -285
rect 9 -297 318 -296
rect 320 -297 535 -296
rect 653 -297 657 -296
rect 660 -297 675 -296
rect 30 -299 164 -298
rect 191 -299 381 -298
rect 387 -299 570 -298
rect 653 -299 661 -298
rect 30 -301 220 -300
rect 247 -301 353 -300
rect 359 -301 612 -300
rect 44 -303 220 -302
rect 247 -303 297 -302
rect 310 -303 507 -302
rect 534 -303 563 -302
rect 569 -303 605 -302
rect 611 -303 633 -302
rect 51 -305 213 -304
rect 215 -305 486 -304
rect 506 -305 514 -304
rect 562 -305 598 -304
rect 604 -305 619 -304
rect 58 -307 153 -306
rect 156 -307 188 -306
rect 191 -307 227 -306
rect 254 -307 500 -306
rect 597 -307 626 -306
rect 65 -309 269 -308
rect 289 -309 514 -308
rect 79 -311 395 -310
rect 401 -311 405 -310
rect 429 -311 486 -310
rect 79 -313 136 -312
rect 170 -313 269 -312
rect 289 -313 391 -312
rect 401 -313 423 -312
rect 432 -313 577 -312
rect 23 -315 171 -314
rect 205 -315 234 -314
rect 240 -315 255 -314
rect 257 -315 304 -314
rect 310 -315 367 -314
rect 373 -315 384 -314
rect 408 -315 577 -314
rect 86 -317 150 -316
rect 313 -317 528 -316
rect 86 -319 276 -318
rect 317 -319 346 -318
rect 352 -319 556 -318
rect 26 -321 346 -320
rect 373 -321 472 -320
rect 478 -321 493 -320
rect 527 -321 591 -320
rect 93 -323 234 -322
rect 331 -323 556 -322
rect 93 -325 143 -324
rect 261 -325 332 -324
rect 338 -325 549 -324
rect 100 -327 251 -326
rect 324 -327 339 -326
rect 341 -327 395 -326
rect 408 -327 542 -326
rect 548 -327 622 -326
rect 100 -329 227 -328
rect 415 -329 423 -328
rect 436 -329 591 -328
rect 110 -331 178 -330
rect 222 -331 262 -330
rect 404 -331 416 -330
rect 457 -331 472 -330
rect 492 -331 521 -330
rect 541 -331 584 -330
rect 72 -333 178 -332
rect 222 -333 363 -332
rect 450 -333 521 -332
rect 72 -335 199 -334
rect 362 -335 430 -334
rect 457 -335 465 -334
rect 107 -337 199 -336
rect 299 -337 465 -336
rect 107 -339 437 -338
rect 114 -341 283 -340
rect 299 -341 444 -340
rect 114 -343 304 -342
rect 443 -343 454 -342
rect 121 -345 164 -344
rect 166 -345 584 -344
rect 128 -347 241 -346
rect 135 -349 279 -348
rect 58 -351 279 -350
rect 142 -353 185 -352
rect 128 -355 185 -354
rect 9 -366 118 -365
rect 128 -366 286 -365
rect 324 -366 640 -365
rect 653 -366 671 -365
rect 674 -366 682 -365
rect 16 -368 143 -367
rect 170 -368 437 -367
rect 453 -368 570 -367
rect 583 -368 654 -367
rect 660 -368 675 -367
rect 23 -370 122 -369
rect 128 -370 209 -369
rect 219 -370 500 -369
rect 520 -370 668 -369
rect 30 -372 325 -371
rect 341 -372 402 -371
rect 408 -372 570 -371
rect 583 -372 612 -371
rect 44 -374 195 -373
rect 212 -374 409 -373
rect 429 -374 619 -373
rect 51 -376 181 -375
rect 229 -376 633 -375
rect 58 -378 297 -377
rect 359 -378 493 -377
rect 506 -378 521 -377
rect 548 -378 612 -377
rect 33 -380 549 -379
rect 555 -380 647 -379
rect 72 -382 153 -381
rect 177 -382 251 -381
rect 254 -382 297 -381
rect 366 -382 458 -381
rect 464 -382 493 -381
rect 562 -382 626 -381
rect 72 -384 87 -383
rect 100 -384 164 -383
rect 275 -384 374 -383
rect 383 -384 577 -383
rect 604 -384 661 -383
rect 65 -386 164 -385
rect 275 -386 304 -385
rect 345 -386 465 -385
rect 471 -386 577 -385
rect 79 -388 223 -387
rect 240 -388 304 -387
rect 338 -388 346 -387
rect 352 -388 458 -387
rect 478 -388 507 -387
rect 527 -388 605 -387
rect 86 -390 265 -389
rect 282 -390 367 -389
rect 383 -390 528 -389
rect 93 -392 223 -391
rect 261 -392 283 -391
rect 289 -392 374 -391
rect 387 -392 451 -391
rect 481 -392 591 -391
rect 93 -394 160 -393
rect 198 -394 241 -393
rect 331 -394 353 -393
rect 355 -394 591 -393
rect 107 -396 167 -395
rect 233 -396 290 -395
rect 310 -396 332 -395
rect 362 -396 563 -395
rect 107 -398 262 -397
rect 317 -398 363 -397
rect 390 -398 598 -397
rect 114 -400 556 -399
rect 121 -402 328 -401
rect 401 -402 416 -401
rect 422 -402 430 -401
rect 436 -402 444 -401
rect 534 -402 598 -401
rect 135 -404 178 -403
rect 268 -404 423 -403
rect 135 -406 157 -405
rect 170 -406 234 -405
rect 317 -406 514 -405
rect 138 -408 255 -407
rect 387 -408 535 -407
rect 142 -410 216 -409
rect 226 -410 269 -409
rect 394 -410 416 -409
rect 485 -410 514 -409
rect 117 -412 486 -411
rect 149 -414 199 -413
rect 247 -414 395 -413
rect 149 -416 192 -415
rect 247 -416 444 -415
rect 184 -418 227 -417
rect 191 -420 542 -419
rect 474 -422 542 -421
rect 16 -433 244 -432
rect 257 -433 367 -432
rect 380 -433 514 -432
rect 541 -433 545 -432
rect 583 -433 703 -432
rect 33 -435 143 -434
rect 149 -435 167 -434
rect 201 -435 563 -434
rect 646 -435 675 -434
rect 40 -437 213 -436
rect 219 -437 549 -436
rect 653 -437 689 -436
rect 44 -439 514 -438
rect 527 -439 584 -438
rect 639 -439 654 -438
rect 44 -441 157 -440
rect 205 -441 465 -440
rect 471 -441 626 -440
rect 632 -441 640 -440
rect 51 -443 384 -442
rect 390 -443 577 -442
rect 611 -443 626 -442
rect 58 -445 297 -444
rect 320 -445 430 -444
rect 450 -445 612 -444
rect 618 -445 633 -444
rect 65 -447 206 -446
rect 222 -447 563 -446
rect 65 -449 349 -448
rect 352 -449 367 -448
rect 390 -449 668 -448
rect 72 -451 174 -450
rect 177 -451 668 -450
rect 72 -453 199 -452
rect 229 -453 241 -452
rect 257 -453 465 -452
rect 478 -453 647 -452
rect 79 -455 122 -454
rect 128 -455 132 -454
rect 135 -455 255 -454
rect 264 -455 416 -454
rect 425 -455 591 -454
rect 82 -457 150 -456
rect 156 -457 304 -456
rect 331 -457 430 -456
rect 439 -457 479 -456
rect 485 -457 528 -456
rect 534 -457 591 -456
rect 93 -459 164 -458
rect 177 -459 339 -458
rect 345 -459 381 -458
rect 401 -459 472 -458
rect 492 -459 535 -458
rect 541 -459 598 -458
rect 100 -461 332 -460
rect 338 -461 409 -460
rect 443 -461 486 -460
rect 499 -461 619 -460
rect 100 -463 199 -462
rect 215 -463 416 -462
rect 436 -463 500 -462
rect 520 -463 577 -462
rect 107 -465 248 -464
rect 275 -465 521 -464
rect 61 -467 276 -466
rect 310 -467 409 -466
rect 450 -467 710 -466
rect 110 -469 444 -468
rect 457 -469 493 -468
rect 114 -471 570 -470
rect 114 -473 363 -472
rect 117 -475 374 -474
rect 128 -477 290 -476
rect 327 -477 374 -476
rect 184 -479 311 -478
rect 355 -479 570 -478
rect 86 -481 185 -480
rect 191 -481 328 -480
rect 359 -481 507 -480
rect 544 -481 598 -480
rect 86 -483 94 -482
rect 194 -483 507 -482
rect 215 -485 423 -484
rect 226 -487 458 -486
rect 226 -489 269 -488
rect 359 -489 605 -488
rect 229 -491 262 -490
rect 268 -491 304 -490
rect 422 -491 549 -490
rect 555 -491 605 -490
rect 37 -493 556 -492
rect 233 -495 353 -494
rect 233 -497 272 -496
rect 240 -499 395 -498
rect 247 -501 321 -500
rect 387 -501 395 -500
rect 261 -503 318 -502
rect 317 -505 661 -504
rect 282 -507 661 -506
rect 282 -509 696 -508
rect 16 -520 346 -519
rect 348 -520 612 -519
rect 23 -522 500 -521
rect 558 -522 675 -521
rect 26 -524 311 -523
rect 324 -524 472 -523
rect 502 -524 675 -523
rect 30 -526 437 -525
rect 460 -526 619 -525
rect 30 -528 465 -527
rect 611 -528 696 -527
rect 37 -530 300 -529
rect 310 -530 419 -529
rect 464 -530 514 -529
rect 618 -530 640 -529
rect 44 -532 286 -531
rect 296 -532 430 -531
rect 513 -532 668 -531
rect 44 -534 101 -533
rect 107 -534 563 -533
rect 576 -534 668 -533
rect 58 -536 258 -535
rect 282 -536 290 -535
rect 327 -536 486 -535
rect 562 -536 584 -535
rect 639 -536 661 -535
rect 51 -538 661 -537
rect 58 -540 374 -539
rect 387 -540 496 -539
rect 65 -542 325 -541
rect 352 -542 391 -541
rect 401 -542 521 -541
rect 65 -544 297 -543
rect 306 -544 584 -543
rect 68 -546 577 -545
rect 72 -548 125 -547
rect 128 -548 321 -547
rect 355 -548 654 -547
rect 54 -550 73 -549
rect 79 -550 220 -549
rect 240 -550 251 -549
rect 254 -550 416 -549
rect 425 -550 430 -549
rect 520 -550 591 -549
rect 79 -552 118 -551
rect 131 -552 402 -551
rect 404 -552 689 -551
rect 86 -554 185 -553
rect 194 -554 556 -553
rect 114 -556 227 -555
rect 233 -556 255 -555
rect 285 -556 528 -555
rect 541 -556 591 -555
rect 107 -558 528 -557
rect 541 -558 598 -557
rect 114 -560 570 -559
rect 135 -562 360 -561
rect 387 -562 451 -561
rect 478 -562 598 -561
rect 135 -564 493 -563
rect 569 -564 626 -563
rect 145 -566 535 -565
rect 625 -566 647 -565
rect 170 -568 199 -567
rect 201 -568 339 -567
rect 408 -568 440 -567
rect 478 -568 507 -567
rect 534 -568 633 -567
rect 177 -570 202 -569
rect 205 -570 269 -569
rect 289 -570 318 -569
rect 320 -570 451 -569
rect 506 -570 605 -569
rect 163 -572 178 -571
rect 184 -572 363 -571
rect 394 -572 409 -571
rect 411 -572 654 -571
rect 159 -574 164 -573
rect 205 -574 213 -573
rect 215 -574 633 -573
rect 215 -576 458 -575
rect 492 -576 605 -575
rect 219 -578 332 -577
rect 422 -578 440 -577
rect 457 -578 710 -577
rect 233 -580 339 -579
rect 548 -580 647 -579
rect 681 -580 710 -579
rect 121 -582 549 -581
rect 121 -584 143 -583
rect 173 -584 682 -583
rect 142 -586 157 -585
rect 240 -586 262 -585
rect 275 -586 332 -585
rect 243 -588 486 -587
rect 247 -590 395 -589
rect 149 -592 248 -591
rect 250 -592 262 -591
rect 275 -592 444 -591
rect 149 -594 192 -593
rect 317 -594 381 -593
rect 443 -594 703 -593
rect 303 -596 381 -595
rect 23 -607 377 -606
rect 411 -607 584 -606
rect 611 -607 738 -606
rect 30 -609 703 -608
rect 709 -609 766 -608
rect 37 -611 73 -610
rect 93 -611 104 -610
rect 107 -611 563 -610
rect 632 -611 773 -610
rect 37 -613 185 -612
rect 187 -613 202 -612
rect 219 -613 661 -612
rect 674 -613 752 -612
rect 44 -615 66 -614
rect 93 -615 381 -614
rect 415 -615 528 -614
rect 541 -615 689 -614
rect 44 -617 216 -616
rect 222 -617 724 -616
rect 51 -619 353 -618
rect 355 -619 745 -618
rect 58 -621 66 -620
rect 100 -621 199 -620
rect 212 -621 223 -620
rect 233 -621 339 -620
rect 348 -621 563 -620
rect 569 -621 661 -620
rect 681 -621 759 -620
rect 23 -623 59 -622
rect 75 -623 234 -622
rect 275 -623 388 -622
rect 418 -623 507 -622
rect 513 -623 717 -622
rect 79 -625 101 -624
rect 107 -625 143 -624
rect 170 -625 192 -624
rect 282 -625 528 -624
rect 555 -625 696 -624
rect 79 -627 206 -626
rect 303 -627 332 -626
rect 380 -627 402 -626
rect 422 -627 444 -626
rect 450 -627 570 -626
rect 583 -627 633 -626
rect 639 -627 710 -626
rect 114 -629 262 -628
rect 296 -629 332 -628
rect 425 -629 654 -628
rect 117 -631 248 -630
rect 261 -631 409 -630
rect 439 -631 535 -630
rect 590 -631 654 -630
rect 54 -633 440 -632
rect 453 -633 640 -632
rect 121 -635 388 -634
rect 457 -635 612 -634
rect 618 -635 682 -634
rect 124 -637 675 -636
rect 128 -639 360 -638
rect 457 -639 521 -638
rect 135 -641 514 -640
rect 142 -643 402 -642
rect 464 -643 556 -642
rect 163 -645 171 -644
rect 198 -645 591 -644
rect 149 -647 164 -646
rect 247 -647 269 -646
rect 296 -647 423 -646
rect 429 -647 465 -646
rect 471 -647 535 -646
rect 19 -649 150 -648
rect 303 -649 405 -648
rect 478 -649 521 -648
rect 86 -651 269 -650
rect 310 -651 409 -650
rect 478 -651 668 -650
rect 86 -653 286 -652
rect 317 -653 731 -652
rect 177 -655 311 -654
rect 320 -655 577 -654
rect 604 -655 668 -654
rect 177 -657 241 -656
rect 359 -657 447 -656
rect 485 -657 542 -656
rect 548 -657 605 -656
rect 159 -659 241 -658
rect 373 -659 577 -658
rect 194 -661 286 -660
rect 324 -661 374 -660
rect 394 -661 430 -660
rect 467 -661 486 -660
rect 492 -661 647 -660
rect 201 -663 549 -662
rect 205 -665 395 -664
rect 460 -665 647 -664
rect 324 -667 619 -666
rect 499 -669 598 -668
rect 135 -671 598 -670
rect 289 -673 500 -672
rect 289 -675 318 -674
rect 30 -686 458 -685
rect 467 -686 759 -685
rect 765 -686 794 -685
rect 37 -688 325 -687
rect 345 -688 640 -687
rect 730 -688 780 -687
rect 37 -690 108 -689
rect 114 -690 423 -689
rect 443 -690 472 -689
rect 485 -690 493 -689
rect 506 -690 766 -689
rect 772 -690 850 -689
rect 44 -692 356 -691
rect 362 -692 367 -691
rect 380 -692 458 -691
rect 495 -692 773 -691
rect 44 -694 94 -693
rect 107 -694 304 -693
rect 320 -694 556 -693
rect 586 -694 752 -693
rect 51 -696 437 -695
rect 450 -696 591 -695
rect 604 -696 640 -695
rect 744 -696 787 -695
rect 54 -698 353 -697
rect 359 -698 367 -697
rect 383 -698 703 -697
rect 58 -700 62 -699
rect 65 -700 328 -699
rect 345 -700 356 -699
rect 397 -700 682 -699
rect 65 -702 500 -701
rect 506 -702 514 -701
rect 555 -702 563 -701
rect 597 -702 605 -701
rect 632 -702 759 -701
rect 72 -704 745 -703
rect 72 -706 94 -705
rect 124 -706 290 -705
rect 296 -706 465 -705
rect 478 -706 633 -705
rect 646 -706 682 -705
rect 86 -708 188 -707
rect 222 -708 311 -707
rect 320 -708 734 -707
rect 89 -710 405 -709
rect 415 -710 591 -709
rect 625 -710 647 -709
rect 653 -710 703 -709
rect 128 -712 262 -711
rect 268 -712 283 -711
rect 289 -712 510 -711
rect 562 -712 570 -711
rect 611 -712 654 -711
rect 79 -714 269 -713
rect 282 -714 752 -713
rect 79 -716 724 -715
rect 131 -718 388 -717
rect 397 -718 689 -717
rect 695 -718 724 -717
rect 16 -720 689 -719
rect 135 -722 584 -721
rect 618 -722 626 -721
rect 135 -724 206 -723
rect 233 -724 395 -723
rect 401 -724 738 -723
rect 114 -726 402 -725
rect 408 -726 416 -725
rect 429 -726 598 -725
rect 621 -726 696 -725
rect 121 -728 234 -727
rect 247 -728 307 -727
rect 348 -728 482 -727
rect 499 -728 535 -727
rect 142 -730 675 -729
rect 124 -732 143 -731
rect 145 -732 160 -731
rect 163 -732 409 -731
rect 429 -732 661 -731
rect 86 -734 661 -733
rect 156 -736 717 -735
rect 156 -738 223 -737
rect 247 -738 304 -737
rect 348 -738 717 -737
rect 163 -740 279 -739
rect 373 -740 388 -739
rect 394 -740 570 -739
rect 184 -742 738 -741
rect 170 -744 185 -743
rect 191 -744 206 -743
rect 254 -744 276 -743
rect 373 -744 489 -743
rect 149 -746 276 -745
rect 436 -746 675 -745
rect 149 -748 710 -747
rect 170 -750 227 -749
rect 254 -750 314 -749
rect 453 -750 514 -749
rect 576 -750 710 -749
rect 177 -752 192 -751
rect 201 -752 612 -751
rect 96 -754 178 -753
rect 201 -754 297 -753
rect 446 -754 577 -753
rect 226 -756 241 -755
rect 261 -756 332 -755
rect 481 -756 668 -755
rect 100 -758 332 -757
rect 439 -758 668 -757
rect 30 -760 101 -759
rect 240 -760 293 -759
rect 439 -760 535 -759
rect 19 -771 24 -770
rect 30 -771 395 -770
rect 408 -771 486 -770
rect 488 -771 836 -770
rect 849 -771 941 -770
rect 23 -773 150 -772
rect 159 -773 276 -772
rect 289 -773 297 -772
rect 310 -773 514 -772
rect 534 -773 710 -772
rect 751 -773 815 -772
rect 37 -775 153 -774
rect 177 -775 181 -774
rect 201 -775 262 -774
rect 268 -775 283 -774
rect 292 -775 458 -774
rect 460 -775 563 -774
rect 621 -775 773 -774
rect 779 -775 850 -774
rect 37 -777 433 -776
rect 446 -777 703 -776
rect 758 -777 829 -776
rect 40 -779 276 -778
rect 296 -779 619 -778
rect 646 -779 780 -778
rect 793 -779 864 -778
rect 54 -781 66 -780
rect 86 -781 220 -780
rect 222 -781 661 -780
rect 667 -781 710 -780
rect 765 -781 843 -780
rect 44 -783 220 -782
rect 226 -783 283 -782
rect 317 -783 346 -782
rect 352 -783 766 -782
rect 44 -785 157 -784
rect 166 -785 647 -784
rect 674 -785 808 -784
rect 58 -787 97 -786
rect 100 -787 311 -786
rect 320 -787 598 -786
rect 688 -787 857 -786
rect 65 -789 465 -788
rect 467 -789 738 -788
rect 72 -791 668 -790
rect 681 -791 738 -790
rect 79 -793 598 -792
rect 639 -793 682 -792
rect 695 -793 752 -792
rect 79 -795 108 -794
rect 114 -795 136 -794
rect 149 -795 290 -794
rect 327 -795 398 -794
rect 411 -795 717 -794
rect 86 -797 731 -796
rect 93 -799 363 -798
rect 397 -799 787 -798
rect 117 -801 584 -800
rect 604 -801 640 -800
rect 653 -801 689 -800
rect 702 -801 724 -800
rect 121 -803 402 -802
rect 408 -803 605 -802
rect 611 -803 654 -802
rect 723 -803 745 -802
rect 72 -805 122 -804
rect 135 -805 192 -804
rect 198 -805 433 -804
rect 436 -805 787 -804
rect 152 -807 318 -806
rect 338 -807 444 -806
rect 446 -807 773 -806
rect 58 -809 339 -808
rect 352 -809 374 -808
rect 429 -809 661 -808
rect 674 -809 745 -808
rect 156 -811 192 -810
rect 226 -811 381 -810
rect 401 -811 430 -810
rect 464 -811 584 -810
rect 625 -811 696 -810
rect 177 -813 185 -812
rect 233 -813 374 -812
rect 513 -813 871 -812
rect 170 -815 234 -814
rect 240 -815 244 -814
rect 247 -815 251 -814
rect 254 -815 517 -814
rect 520 -815 535 -814
rect 537 -815 717 -814
rect 142 -817 171 -816
rect 184 -817 206 -816
rect 240 -817 388 -816
rect 548 -817 563 -816
rect 569 -817 759 -816
rect 142 -819 591 -818
rect 163 -821 255 -820
rect 268 -821 458 -820
rect 499 -821 549 -820
rect 555 -821 570 -820
rect 576 -821 626 -820
rect 128 -823 577 -822
rect 128 -825 423 -824
rect 471 -825 500 -824
rect 541 -825 556 -824
rect 163 -827 325 -826
rect 331 -827 521 -826
rect 527 -827 542 -826
rect 107 -829 325 -828
rect 331 -829 801 -828
rect 243 -831 388 -830
rect 471 -831 493 -830
rect 506 -831 528 -830
rect 299 -833 423 -832
rect 506 -833 822 -832
rect 306 -835 591 -834
rect 100 -837 307 -836
rect 355 -837 416 -836
rect 359 -839 612 -838
rect 198 -841 360 -840
rect 366 -841 416 -840
rect 366 -843 633 -842
rect 383 -845 493 -844
rect 450 -847 633 -846
rect 450 -849 479 -848
rect 9 -860 594 -859
rect 674 -860 864 -859
rect 16 -862 192 -861
rect 201 -862 279 -861
rect 282 -862 335 -861
rect 338 -862 367 -861
rect 404 -862 563 -861
rect 660 -862 675 -861
rect 831 -862 941 -861
rect 30 -864 223 -863
rect 240 -864 307 -863
rect 317 -864 409 -863
rect 411 -864 787 -863
rect 44 -866 160 -865
rect 163 -866 794 -865
rect 44 -868 353 -867
rect 359 -868 535 -867
rect 562 -868 612 -867
rect 653 -868 661 -867
rect 58 -870 251 -869
rect 261 -870 367 -869
rect 429 -870 815 -869
rect 72 -872 640 -871
rect 653 -872 731 -871
rect 744 -872 815 -871
rect 72 -874 108 -873
rect 121 -874 125 -873
rect 135 -874 265 -873
rect 268 -874 325 -873
rect 327 -874 857 -873
rect 23 -876 136 -875
rect 142 -876 290 -875
rect 317 -876 381 -875
rect 387 -876 430 -875
rect 443 -876 836 -875
rect 23 -878 521 -877
rect 590 -878 787 -877
rect 75 -880 374 -879
rect 387 -880 423 -879
rect 453 -880 528 -879
rect 597 -880 640 -879
rect 730 -880 759 -879
rect 79 -882 297 -881
rect 310 -882 423 -881
rect 457 -882 500 -881
rect 506 -882 710 -881
rect 744 -882 766 -881
rect 79 -884 528 -883
rect 611 -884 626 -883
rect 702 -884 759 -883
rect 765 -884 801 -883
rect 82 -886 486 -885
rect 506 -886 689 -885
rect 709 -886 738 -885
rect 800 -886 829 -885
rect 86 -888 115 -887
rect 142 -888 164 -887
rect 166 -888 178 -887
rect 184 -888 311 -887
rect 345 -888 374 -887
rect 439 -888 500 -887
rect 534 -888 829 -887
rect 30 -890 346 -889
rect 362 -890 437 -889
rect 460 -890 843 -889
rect 51 -892 115 -891
rect 177 -892 227 -891
rect 233 -892 269 -891
rect 464 -892 598 -891
rect 625 -892 696 -891
rect 737 -892 752 -891
rect 842 -892 871 -891
rect 40 -894 234 -893
rect 254 -894 290 -893
rect 467 -894 570 -893
rect 583 -894 703 -893
rect 751 -894 773 -893
rect 51 -896 416 -895
rect 478 -896 517 -895
rect 555 -896 570 -895
rect 681 -896 689 -895
rect 695 -896 780 -895
rect 86 -898 157 -897
rect 170 -898 227 -897
rect 254 -898 300 -897
rect 471 -898 517 -897
rect 541 -898 556 -897
rect 667 -898 682 -897
rect 716 -898 780 -897
rect 93 -900 150 -899
rect 156 -900 283 -899
rect 446 -900 668 -899
rect 716 -900 724 -899
rect 772 -900 822 -899
rect 93 -902 402 -901
rect 471 -902 493 -901
rect 646 -902 724 -901
rect 821 -902 850 -901
rect 54 -904 493 -903
rect 632 -904 647 -903
rect 835 -904 850 -903
rect 100 -906 808 -905
rect 65 -908 101 -907
rect 103 -908 349 -907
rect 401 -908 584 -907
rect 618 -908 633 -907
rect 107 -910 146 -909
rect 191 -910 199 -909
rect 205 -910 360 -909
rect 485 -910 591 -909
rect 604 -910 619 -909
rect 58 -912 199 -911
rect 212 -912 241 -911
rect 261 -912 339 -911
rect 548 -912 605 -911
rect 128 -914 447 -913
rect 128 -916 185 -915
rect 215 -916 521 -915
rect 170 -918 206 -917
rect 219 -918 332 -917
rect 380 -918 549 -917
rect 219 -920 416 -919
rect 275 -922 479 -921
rect 303 -924 808 -923
rect 19 -926 304 -925
rect 331 -926 342 -925
rect 2 -937 234 -936
rect 247 -937 262 -936
rect 275 -937 360 -936
rect 390 -937 724 -936
rect 779 -937 899 -936
rect 9 -939 83 -938
rect 100 -939 339 -938
rect 348 -939 787 -938
rect 814 -939 850 -938
rect 9 -941 129 -940
rect 149 -941 171 -940
rect 173 -941 388 -940
rect 394 -941 437 -940
rect 450 -941 864 -940
rect 16 -943 335 -942
rect 352 -943 500 -942
rect 509 -943 738 -942
rect 786 -943 829 -942
rect 30 -945 297 -944
rect 331 -945 360 -944
rect 397 -945 675 -944
rect 716 -945 780 -944
rect 814 -945 836 -944
rect 37 -947 125 -946
rect 128 -947 223 -946
rect 247 -947 314 -946
rect 331 -947 703 -946
rect 737 -947 745 -946
rect 40 -949 73 -948
rect 79 -949 381 -948
rect 401 -949 668 -948
rect 744 -949 752 -948
rect 44 -951 286 -950
rect 404 -951 409 -950
rect 429 -951 500 -950
rect 513 -951 661 -950
rect 751 -951 808 -950
rect 51 -953 94 -952
rect 117 -953 577 -952
rect 590 -953 822 -952
rect 58 -955 395 -954
rect 408 -955 605 -954
rect 646 -955 668 -954
rect 793 -955 808 -954
rect 58 -957 94 -956
rect 121 -957 195 -956
rect 201 -957 283 -956
rect 303 -957 591 -956
rect 646 -957 689 -956
rect 44 -959 122 -958
rect 152 -959 836 -958
rect 61 -961 412 -960
rect 429 -961 829 -960
rect 65 -963 87 -962
rect 163 -963 486 -962
rect 516 -963 794 -962
rect 65 -965 374 -964
rect 436 -965 633 -964
rect 653 -965 703 -964
rect 72 -967 157 -966
rect 177 -967 304 -966
rect 373 -967 381 -966
rect 443 -967 822 -966
rect 86 -969 318 -968
rect 443 -969 458 -968
rect 464 -969 472 -968
rect 474 -969 724 -968
rect 135 -971 157 -970
rect 177 -971 227 -970
rect 254 -971 297 -970
rect 317 -971 346 -970
rect 446 -971 717 -970
rect 135 -973 202 -972
rect 205 -973 857 -972
rect 170 -975 227 -974
rect 254 -975 454 -974
rect 457 -975 493 -974
rect 541 -975 619 -974
rect 653 -975 682 -974
rect 688 -975 696 -974
rect 191 -977 234 -976
rect 261 -977 269 -976
rect 278 -977 423 -976
rect 450 -977 479 -976
rect 481 -977 542 -976
rect 548 -977 801 -976
rect 208 -979 640 -978
rect 695 -979 731 -978
rect 772 -979 801 -978
rect 212 -981 388 -980
rect 478 -981 661 -980
rect 765 -981 773 -980
rect 215 -983 311 -982
rect 338 -983 549 -982
rect 562 -983 619 -982
rect 639 -983 710 -982
rect 758 -983 766 -982
rect 184 -985 710 -984
rect 758 -985 874 -984
rect 142 -987 185 -986
rect 219 -987 241 -986
rect 268 -987 353 -986
rect 376 -987 731 -986
rect 114 -989 143 -988
rect 240 -989 416 -988
rect 485 -989 570 -988
rect 576 -989 598 -988
rect 114 -991 675 -990
rect 289 -993 633 -992
rect 289 -995 325 -994
rect 345 -995 367 -994
rect 404 -995 416 -994
rect 555 -995 563 -994
rect 583 -995 682 -994
rect 23 -997 367 -996
rect 555 -997 626 -996
rect 23 -999 108 -998
rect 299 -999 493 -998
rect 558 -999 570 -998
rect 597 -999 860 -998
rect 107 -1001 132 -1000
rect 324 -1001 507 -1000
rect 611 -1001 626 -1000
rect 425 -1003 612 -1002
rect 506 -1005 605 -1004
rect 2 -1016 412 -1015
rect 422 -1016 542 -1015
rect 551 -1016 724 -1015
rect 786 -1016 857 -1015
rect 863 -1016 920 -1015
rect 9 -1018 171 -1017
rect 212 -1018 339 -1017
rect 341 -1018 493 -1017
rect 502 -1018 843 -1017
rect 849 -1018 913 -1017
rect 16 -1020 206 -1019
rect 212 -1020 402 -1019
rect 404 -1020 486 -1019
rect 492 -1020 885 -1019
rect 898 -1020 927 -1019
rect 19 -1022 787 -1021
rect 800 -1022 878 -1021
rect 23 -1024 27 -1023
rect 30 -1024 199 -1023
rect 205 -1024 262 -1023
rect 303 -1024 468 -1023
rect 478 -1024 640 -1023
rect 642 -1024 843 -1023
rect 23 -1026 157 -1025
rect 166 -1026 234 -1025
rect 261 -1026 559 -1025
rect 590 -1026 892 -1025
rect 33 -1028 710 -1027
rect 772 -1028 801 -1027
rect 807 -1028 871 -1027
rect 37 -1030 192 -1029
rect 219 -1030 283 -1029
rect 303 -1030 325 -1029
rect 331 -1030 731 -1029
rect 772 -1030 860 -1029
rect 37 -1032 87 -1031
rect 93 -1032 437 -1031
rect 439 -1032 479 -1031
rect 506 -1032 612 -1031
rect 660 -1032 724 -1031
rect 779 -1032 850 -1031
rect 54 -1034 87 -1033
rect 107 -1034 409 -1033
rect 415 -1034 486 -1033
rect 513 -1034 752 -1033
rect 821 -1034 941 -1033
rect 58 -1036 160 -1035
rect 163 -1036 514 -1035
rect 516 -1036 598 -1035
rect 604 -1036 615 -1035
rect 681 -1036 731 -1035
rect 828 -1036 899 -1035
rect 65 -1038 416 -1037
rect 432 -1038 444 -1037
rect 446 -1038 808 -1037
rect 835 -1038 906 -1037
rect 65 -1040 255 -1039
rect 278 -1040 283 -1039
rect 289 -1040 507 -1039
rect 527 -1040 591 -1039
rect 604 -1040 745 -1039
rect 72 -1042 115 -1041
rect 121 -1042 143 -1041
rect 163 -1042 815 -1041
rect 72 -1044 150 -1043
rect 152 -1044 815 -1043
rect 79 -1046 311 -1045
rect 317 -1046 402 -1045
rect 453 -1046 573 -1045
rect 576 -1046 661 -1045
rect 674 -1046 745 -1045
rect 79 -1048 276 -1047
rect 296 -1048 325 -1047
rect 352 -1048 395 -1047
rect 499 -1048 829 -1047
rect 103 -1050 115 -1049
rect 128 -1050 668 -1049
rect 688 -1050 822 -1049
rect 107 -1052 118 -1051
rect 128 -1052 335 -1051
rect 352 -1052 584 -1051
rect 614 -1052 675 -1051
rect 695 -1052 864 -1051
rect 135 -1054 143 -1053
rect 170 -1054 269 -1053
rect 275 -1054 451 -1053
rect 464 -1054 500 -1053
rect 520 -1054 577 -1053
rect 716 -1054 780 -1053
rect 177 -1056 234 -1055
rect 243 -1056 290 -1055
rect 317 -1056 496 -1055
rect 527 -1056 682 -1055
rect 737 -1056 836 -1055
rect 100 -1058 178 -1057
rect 184 -1058 255 -1057
rect 268 -1058 349 -1057
rect 359 -1058 374 -1057
rect 380 -1058 391 -1057
rect 429 -1058 521 -1057
rect 534 -1058 696 -1057
rect 191 -1060 223 -1059
rect 226 -1060 542 -1059
rect 565 -1060 668 -1059
rect 44 -1062 223 -1061
rect 226 -1062 241 -1061
rect 247 -1062 297 -1061
rect 345 -1062 381 -1061
rect 387 -1062 633 -1061
rect 646 -1062 738 -1061
rect 44 -1064 52 -1063
rect 201 -1064 332 -1063
rect 345 -1064 759 -1063
rect 359 -1066 538 -1065
rect 548 -1066 633 -1065
rect 653 -1066 717 -1065
rect 758 -1066 766 -1065
rect 184 -1068 549 -1067
rect 562 -1068 647 -1067
rect 366 -1070 612 -1069
rect 625 -1070 766 -1069
rect 366 -1072 531 -1071
rect 534 -1072 752 -1071
rect 376 -1074 654 -1073
rect 390 -1076 472 -1075
rect 562 -1076 710 -1075
rect 429 -1078 458 -1077
rect 569 -1078 598 -1077
rect 607 -1078 626 -1077
rect 194 -1080 458 -1079
rect 450 -1082 689 -1081
rect 9 -1093 787 -1092
rect 884 -1093 976 -1092
rect 982 -1093 990 -1092
rect 9 -1095 171 -1094
rect 198 -1095 227 -1094
rect 240 -1095 283 -1094
rect 317 -1095 444 -1094
rect 446 -1095 892 -1094
rect 898 -1095 969 -1094
rect 16 -1097 580 -1096
rect 642 -1097 850 -1096
rect 856 -1097 899 -1096
rect 912 -1097 948 -1096
rect 16 -1099 31 -1098
rect 44 -1099 97 -1098
rect 103 -1099 717 -1098
rect 828 -1099 885 -1098
rect 30 -1101 38 -1100
rect 44 -1101 206 -1100
rect 226 -1101 311 -1100
rect 345 -1101 367 -1100
rect 387 -1101 409 -1100
rect 436 -1101 440 -1100
rect 450 -1101 640 -1100
rect 667 -1101 934 -1100
rect 37 -1103 269 -1102
rect 275 -1103 321 -1102
rect 348 -1103 416 -1102
rect 436 -1103 493 -1102
rect 506 -1103 535 -1102
rect 544 -1103 822 -1102
rect 842 -1103 892 -1102
rect 51 -1105 87 -1104
rect 93 -1105 913 -1104
rect 58 -1107 66 -1106
rect 72 -1107 153 -1106
rect 156 -1107 178 -1106
rect 198 -1107 556 -1106
rect 558 -1107 864 -1106
rect 58 -1109 255 -1108
rect 268 -1109 297 -1108
rect 303 -1109 311 -1108
rect 355 -1109 696 -1108
rect 702 -1109 857 -1108
rect 863 -1109 930 -1108
rect 72 -1111 202 -1110
rect 205 -1111 363 -1110
rect 366 -1111 633 -1110
rect 684 -1111 878 -1110
rect 82 -1113 220 -1112
rect 247 -1113 290 -1112
rect 303 -1113 325 -1112
rect 355 -1113 416 -1112
rect 439 -1113 493 -1112
rect 520 -1113 605 -1112
rect 607 -1113 668 -1112
rect 702 -1113 717 -1112
rect 751 -1113 843 -1112
rect 849 -1113 962 -1112
rect 86 -1115 108 -1114
rect 128 -1115 297 -1114
rect 331 -1115 605 -1114
rect 758 -1115 822 -1114
rect 103 -1117 255 -1116
rect 278 -1117 752 -1116
rect 800 -1117 829 -1116
rect 107 -1119 115 -1118
rect 128 -1119 143 -1118
rect 152 -1119 507 -1118
rect 527 -1119 738 -1118
rect 114 -1121 381 -1120
rect 390 -1121 920 -1120
rect 135 -1123 787 -1122
rect 870 -1123 920 -1122
rect 135 -1125 521 -1124
rect 530 -1125 906 -1124
rect 138 -1127 234 -1126
rect 250 -1127 696 -1126
rect 772 -1127 871 -1126
rect 23 -1129 234 -1128
rect 282 -1129 528 -1128
rect 562 -1129 815 -1128
rect 93 -1131 773 -1130
rect 793 -1131 906 -1130
rect 142 -1133 430 -1132
rect 453 -1133 689 -1132
rect 709 -1133 815 -1132
rect 163 -1135 262 -1134
rect 289 -1135 360 -1134
rect 380 -1135 395 -1134
rect 422 -1135 689 -1134
rect 166 -1137 878 -1136
rect 177 -1139 192 -1138
rect 261 -1139 486 -1138
rect 562 -1139 927 -1138
rect 184 -1141 430 -1140
rect 464 -1141 836 -1140
rect 170 -1143 185 -1142
rect 191 -1143 213 -1142
rect 324 -1143 454 -1142
rect 485 -1143 510 -1142
rect 569 -1143 801 -1142
rect 331 -1145 591 -1144
rect 618 -1145 759 -1144
rect 338 -1147 423 -1146
rect 513 -1147 570 -1146
rect 572 -1147 766 -1146
rect 222 -1149 766 -1148
rect 222 -1151 395 -1150
rect 401 -1151 514 -1150
rect 576 -1151 633 -1150
rect 646 -1151 710 -1150
rect 730 -1151 836 -1150
rect 338 -1153 374 -1152
rect 583 -1153 640 -1152
rect 646 -1153 682 -1152
rect 359 -1155 780 -1154
rect 373 -1157 451 -1156
rect 548 -1157 682 -1156
rect 744 -1157 780 -1156
rect 79 -1159 745 -1158
rect 79 -1161 122 -1160
rect 425 -1161 584 -1160
rect 618 -1161 724 -1160
rect 625 -1163 794 -1162
rect 611 -1165 626 -1164
rect 653 -1165 724 -1164
rect 597 -1167 612 -1166
rect 656 -1167 927 -1166
rect 499 -1169 598 -1168
rect 660 -1169 731 -1168
rect 478 -1171 500 -1170
rect 541 -1171 661 -1170
rect 674 -1171 738 -1170
rect 401 -1173 479 -1172
rect 541 -1173 591 -1172
rect 457 -1175 675 -1174
rect 457 -1177 472 -1176
rect 212 -1179 472 -1178
rect 5 -1190 220 -1189
rect 222 -1190 675 -1189
rect 719 -1190 829 -1189
rect 940 -1190 965 -1189
rect 975 -1190 983 -1189
rect 985 -1190 1011 -1189
rect 9 -1192 213 -1191
rect 215 -1192 724 -1191
rect 737 -1192 741 -1191
rect 751 -1192 955 -1191
rect 989 -1192 1004 -1191
rect 16 -1194 216 -1193
rect 254 -1194 307 -1193
rect 341 -1194 619 -1193
rect 625 -1194 717 -1193
rect 723 -1194 745 -1193
rect 800 -1194 829 -1193
rect 968 -1194 990 -1193
rect 16 -1196 178 -1195
rect 201 -1196 766 -1195
rect 800 -1196 885 -1195
rect 912 -1196 969 -1195
rect 44 -1198 314 -1197
rect 352 -1198 486 -1197
rect 506 -1198 899 -1197
rect 58 -1200 174 -1199
rect 254 -1200 363 -1199
rect 373 -1200 423 -1199
rect 429 -1200 766 -1199
rect 814 -1200 997 -1199
rect 58 -1202 461 -1201
rect 464 -1202 794 -1201
rect 814 -1202 927 -1201
rect 72 -1204 199 -1203
rect 268 -1204 318 -1203
rect 355 -1204 367 -1203
rect 411 -1204 689 -1203
rect 737 -1204 857 -1203
rect 65 -1206 367 -1205
rect 411 -1206 682 -1205
rect 842 -1206 857 -1205
rect 65 -1208 500 -1207
rect 534 -1208 689 -1207
rect 786 -1208 843 -1207
rect 849 -1208 913 -1207
rect 86 -1210 122 -1209
rect 135 -1210 227 -1209
rect 268 -1210 304 -1209
rect 310 -1210 374 -1209
rect 429 -1210 563 -1209
rect 579 -1210 976 -1209
rect 79 -1212 136 -1211
rect 142 -1212 321 -1211
rect 359 -1212 808 -1211
rect 30 -1214 143 -1213
rect 149 -1214 332 -1213
rect 446 -1214 710 -1213
rect 772 -1214 787 -1213
rect 30 -1216 409 -1215
rect 450 -1216 598 -1215
rect 604 -1216 675 -1215
rect 740 -1216 773 -1215
rect 779 -1216 850 -1215
rect 12 -1218 409 -1217
rect 436 -1218 451 -1217
rect 453 -1218 759 -1217
rect 79 -1220 325 -1219
rect 464 -1220 934 -1219
rect 86 -1222 153 -1221
rect 163 -1222 199 -1221
rect 226 -1222 496 -1221
rect 520 -1222 563 -1221
rect 583 -1222 927 -1221
rect 93 -1224 206 -1223
rect 233 -1224 325 -1223
rect 467 -1224 654 -1223
rect 656 -1224 906 -1223
rect 37 -1226 206 -1225
rect 233 -1226 402 -1225
rect 474 -1226 521 -1225
rect 527 -1226 535 -1225
rect 541 -1226 958 -1225
rect 93 -1228 633 -1227
rect 635 -1228 808 -1227
rect 877 -1228 934 -1227
rect 96 -1230 164 -1229
rect 170 -1230 178 -1229
rect 275 -1230 745 -1229
rect 758 -1230 871 -1229
rect 877 -1230 948 -1229
rect 96 -1232 332 -1231
rect 401 -1232 468 -1231
rect 471 -1232 542 -1231
rect 544 -1232 899 -1231
rect 100 -1234 157 -1233
rect 285 -1234 493 -1233
rect 555 -1234 626 -1233
rect 639 -1234 710 -1233
rect 863 -1234 871 -1233
rect 103 -1236 696 -1235
rect 107 -1238 122 -1237
rect 128 -1238 157 -1237
rect 296 -1238 437 -1237
rect 457 -1238 528 -1237
rect 583 -1238 591 -1237
rect 597 -1238 696 -1237
rect 44 -1240 129 -1239
rect 149 -1240 185 -1239
rect 296 -1240 346 -1239
rect 394 -1240 640 -1239
rect 646 -1240 794 -1239
rect 110 -1242 192 -1241
rect 303 -1242 426 -1241
rect 457 -1242 731 -1241
rect 114 -1244 577 -1243
rect 604 -1244 752 -1243
rect 51 -1246 115 -1245
rect 184 -1246 276 -1245
rect 338 -1246 395 -1245
rect 471 -1246 962 -1245
rect 51 -1248 262 -1247
rect 345 -1248 381 -1247
rect 478 -1248 906 -1247
rect 191 -1250 223 -1249
rect 261 -1250 290 -1249
rect 380 -1250 591 -1249
rect 607 -1250 822 -1249
rect 891 -1250 962 -1249
rect 212 -1252 731 -1251
rect 835 -1252 892 -1251
rect 289 -1254 388 -1253
rect 443 -1254 479 -1253
rect 492 -1254 780 -1253
rect 310 -1256 836 -1255
rect 387 -1258 416 -1257
rect 443 -1258 486 -1257
rect 513 -1258 556 -1257
rect 600 -1258 822 -1257
rect 282 -1260 416 -1259
rect 513 -1260 549 -1259
rect 646 -1260 944 -1259
rect 240 -1262 283 -1261
rect 548 -1262 570 -1261
rect 656 -1262 920 -1261
rect 40 -1264 241 -1263
rect 569 -1264 920 -1263
rect 660 -1266 864 -1265
rect 660 -1268 703 -1267
rect 124 -1270 703 -1269
rect 667 -1272 885 -1271
rect 670 -1274 948 -1273
rect 9 -1285 31 -1284
rect 37 -1285 150 -1284
rect 170 -1285 220 -1284
rect 222 -1285 290 -1284
rect 310 -1285 577 -1284
rect 579 -1285 927 -1284
rect 943 -1285 1011 -1284
rect 30 -1287 689 -1286
rect 971 -1287 990 -1286
rect 44 -1289 216 -1288
rect 226 -1289 507 -1288
rect 509 -1289 696 -1288
rect 940 -1289 990 -1288
rect 44 -1291 87 -1290
rect 89 -1291 454 -1290
rect 457 -1291 542 -1290
rect 569 -1291 955 -1290
rect 51 -1293 342 -1292
rect 408 -1293 437 -1292
rect 446 -1293 493 -1292
rect 499 -1293 710 -1292
rect 954 -1293 1004 -1292
rect 51 -1295 97 -1294
rect 124 -1295 227 -1294
rect 240 -1295 290 -1294
rect 310 -1295 318 -1294
rect 352 -1295 500 -1294
rect 569 -1295 584 -1294
rect 597 -1295 612 -1294
rect 618 -1295 920 -1294
rect 58 -1297 174 -1296
rect 184 -1297 864 -1296
rect 919 -1297 976 -1296
rect 61 -1299 108 -1298
rect 135 -1299 185 -1298
rect 198 -1299 220 -1298
rect 229 -1299 864 -1298
rect 65 -1301 353 -1300
rect 387 -1301 409 -1300
rect 411 -1301 899 -1300
rect 65 -1303 381 -1302
rect 387 -1303 556 -1302
rect 576 -1303 913 -1302
rect 72 -1305 129 -1304
rect 149 -1305 262 -1304
rect 282 -1305 360 -1304
rect 415 -1305 465 -1304
rect 467 -1305 489 -1304
rect 502 -1305 584 -1304
rect 632 -1305 661 -1304
rect 667 -1305 892 -1304
rect 898 -1305 983 -1304
rect 16 -1307 262 -1306
rect 296 -1307 360 -1306
rect 366 -1307 465 -1306
rect 471 -1307 794 -1306
rect 16 -1309 111 -1308
rect 114 -1309 136 -1308
rect 163 -1309 283 -1308
rect 303 -1309 472 -1308
rect 474 -1309 647 -1308
rect 653 -1309 892 -1308
rect 72 -1311 731 -1310
rect 793 -1311 850 -1310
rect 12 -1313 731 -1312
rect 93 -1315 531 -1314
rect 548 -1315 612 -1314
rect 646 -1315 717 -1314
rect 114 -1317 122 -1316
rect 128 -1317 255 -1316
rect 317 -1317 325 -1316
rect 331 -1317 619 -1316
rect 653 -1317 703 -1316
rect 709 -1317 836 -1316
rect 121 -1319 626 -1318
rect 656 -1319 997 -1318
rect 156 -1321 164 -1320
rect 177 -1321 325 -1320
rect 415 -1321 944 -1320
rect 142 -1323 178 -1322
rect 191 -1323 199 -1322
rect 208 -1323 507 -1322
rect 534 -1323 549 -1322
rect 590 -1323 661 -1322
rect 667 -1323 808 -1322
rect 835 -1323 934 -1322
rect 100 -1325 192 -1324
rect 212 -1325 297 -1324
rect 313 -1325 591 -1324
rect 625 -1325 682 -1324
rect 688 -1325 780 -1324
rect 100 -1327 157 -1326
rect 233 -1327 332 -1326
rect 429 -1327 556 -1326
rect 674 -1327 913 -1326
rect 142 -1329 528 -1328
rect 562 -1329 675 -1328
rect 702 -1329 787 -1328
rect 233 -1331 402 -1330
rect 432 -1331 766 -1330
rect 240 -1333 423 -1332
rect 436 -1333 451 -1332
rect 460 -1333 850 -1332
rect 247 -1335 384 -1334
rect 394 -1335 423 -1334
rect 443 -1335 808 -1334
rect 205 -1337 248 -1336
rect 254 -1337 346 -1336
rect 366 -1337 395 -1336
rect 443 -1337 479 -1336
rect 481 -1337 885 -1336
rect 303 -1339 430 -1338
rect 450 -1339 521 -1338
rect 527 -1339 542 -1338
rect 716 -1339 752 -1338
rect 765 -1339 829 -1338
rect 877 -1339 885 -1338
rect 338 -1341 402 -1340
rect 478 -1341 535 -1340
rect 639 -1341 752 -1340
rect 814 -1341 878 -1340
rect 338 -1343 374 -1342
rect 383 -1343 780 -1342
rect 814 -1343 857 -1342
rect 268 -1345 374 -1344
rect 485 -1345 682 -1344
rect 737 -1345 787 -1344
rect 800 -1345 857 -1344
rect 268 -1347 276 -1346
rect 513 -1347 563 -1346
rect 639 -1347 745 -1346
rect 758 -1347 801 -1346
rect 828 -1347 906 -1346
rect 79 -1349 276 -1348
rect 485 -1349 745 -1348
rect 758 -1349 969 -1348
rect 79 -1351 605 -1350
rect 695 -1351 906 -1350
rect 513 -1353 843 -1352
rect 520 -1355 605 -1354
rect 737 -1355 822 -1354
rect 842 -1355 948 -1354
rect 821 -1357 871 -1356
rect 870 -1359 962 -1358
rect 2 -1370 45 -1369
rect 58 -1370 80 -1369
rect 86 -1370 136 -1369
rect 156 -1370 353 -1369
rect 376 -1370 773 -1369
rect 856 -1370 906 -1369
rect 908 -1370 955 -1369
rect 971 -1370 990 -1369
rect 9 -1372 325 -1371
rect 394 -1372 682 -1371
rect 712 -1372 717 -1371
rect 765 -1372 927 -1371
rect 947 -1372 955 -1371
rect 9 -1374 731 -1373
rect 765 -1374 899 -1373
rect 912 -1374 969 -1373
rect 37 -1376 230 -1375
rect 240 -1376 381 -1375
rect 397 -1376 409 -1375
rect 450 -1376 461 -1375
rect 467 -1376 759 -1375
rect 856 -1376 871 -1375
rect 891 -1376 913 -1375
rect 37 -1378 195 -1377
rect 205 -1378 339 -1377
rect 348 -1378 717 -1377
rect 744 -1378 759 -1377
rect 800 -1378 871 -1377
rect 51 -1380 381 -1379
rect 401 -1380 468 -1379
rect 478 -1380 654 -1379
rect 681 -1380 696 -1379
rect 702 -1380 731 -1379
rect 800 -1380 822 -1379
rect 849 -1380 892 -1379
rect 51 -1382 269 -1381
rect 296 -1382 377 -1381
rect 401 -1382 563 -1381
rect 576 -1382 598 -1381
rect 604 -1382 829 -1381
rect 842 -1382 850 -1381
rect 863 -1382 934 -1381
rect 65 -1384 188 -1383
rect 191 -1384 773 -1383
rect 807 -1384 843 -1383
rect 863 -1384 941 -1383
rect 33 -1386 66 -1385
rect 72 -1386 552 -1385
rect 555 -1386 696 -1385
rect 702 -1386 738 -1385
rect 72 -1388 458 -1387
rect 464 -1388 563 -1387
rect 590 -1388 920 -1387
rect 79 -1390 335 -1389
rect 338 -1390 493 -1389
rect 516 -1390 689 -1389
rect 723 -1390 745 -1389
rect 89 -1392 584 -1391
rect 593 -1392 878 -1391
rect 93 -1394 206 -1393
rect 226 -1394 559 -1393
rect 569 -1394 584 -1393
rect 604 -1394 808 -1393
rect 877 -1394 885 -1393
rect 93 -1396 115 -1395
rect 124 -1396 752 -1395
rect 835 -1396 885 -1395
rect 100 -1398 556 -1397
rect 667 -1398 689 -1397
rect 709 -1398 724 -1397
rect 751 -1398 794 -1397
rect 835 -1398 944 -1397
rect 23 -1400 101 -1399
rect 128 -1400 297 -1399
rect 310 -1400 374 -1399
rect 453 -1400 738 -1399
rect 779 -1400 794 -1399
rect 943 -1400 983 -1399
rect 23 -1402 255 -1401
rect 261 -1402 346 -1401
rect 373 -1402 668 -1401
rect 121 -1404 346 -1403
rect 478 -1404 500 -1403
rect 527 -1404 787 -1403
rect 121 -1406 220 -1405
rect 233 -1406 409 -1405
rect 471 -1406 528 -1405
rect 530 -1406 675 -1405
rect 786 -1406 815 -1405
rect 135 -1408 290 -1407
rect 310 -1408 318 -1407
rect 331 -1408 570 -1407
rect 646 -1408 675 -1407
rect 149 -1410 262 -1409
rect 289 -1410 367 -1409
rect 390 -1410 472 -1409
rect 481 -1410 899 -1409
rect 107 -1412 150 -1411
rect 159 -1412 241 -1411
rect 247 -1412 353 -1411
rect 366 -1412 388 -1411
rect 485 -1412 549 -1411
rect 632 -1412 647 -1411
rect 660 -1412 780 -1411
rect 30 -1414 160 -1413
rect 166 -1414 192 -1413
rect 219 -1414 223 -1413
rect 233 -1414 514 -1413
rect 537 -1414 626 -1413
rect 632 -1414 815 -1413
rect 107 -1416 118 -1415
rect 170 -1416 269 -1415
rect 317 -1416 433 -1415
rect 492 -1416 507 -1415
rect 513 -1416 521 -1415
rect 534 -1416 626 -1415
rect 639 -1416 661 -1415
rect 16 -1418 507 -1417
rect 541 -1418 598 -1417
rect 16 -1420 304 -1419
rect 464 -1420 521 -1419
rect 541 -1420 612 -1419
rect 163 -1422 171 -1421
rect 177 -1422 248 -1421
rect 254 -1422 360 -1421
rect 488 -1422 640 -1421
rect 128 -1424 178 -1423
rect 184 -1424 332 -1423
rect 499 -1424 619 -1423
rect 212 -1426 304 -1425
rect 509 -1426 612 -1425
rect 282 -1428 360 -1427
rect 579 -1428 619 -1427
rect 282 -1430 416 -1429
rect 579 -1430 822 -1429
rect 415 -1432 423 -1431
rect 422 -1434 437 -1433
rect 436 -1436 444 -1435
rect 142 -1438 444 -1437
rect 9 -1449 17 -1448
rect 23 -1449 395 -1448
rect 432 -1449 521 -1448
rect 548 -1449 871 -1448
rect 940 -1449 969 -1448
rect 16 -1451 227 -1450
rect 282 -1451 395 -1450
rect 457 -1451 500 -1450
rect 502 -1451 731 -1450
rect 961 -1451 983 -1450
rect 23 -1453 38 -1452
rect 44 -1453 108 -1452
rect 114 -1453 283 -1452
rect 285 -1453 514 -1452
rect 555 -1453 885 -1452
rect 982 -1453 990 -1452
rect 51 -1455 363 -1454
rect 373 -1455 416 -1454
rect 432 -1455 500 -1454
rect 506 -1455 864 -1454
rect 51 -1457 552 -1456
rect 558 -1457 927 -1456
rect 79 -1459 591 -1458
rect 604 -1459 780 -1458
rect 79 -1461 223 -1460
rect 303 -1461 391 -1460
rect 397 -1461 780 -1460
rect 93 -1463 132 -1462
rect 142 -1463 332 -1462
rect 338 -1463 430 -1462
rect 460 -1463 899 -1462
rect 93 -1465 318 -1464
rect 345 -1465 549 -1464
rect 576 -1465 612 -1464
rect 632 -1465 906 -1464
rect 100 -1467 318 -1466
rect 352 -1467 367 -1466
rect 376 -1467 381 -1466
rect 415 -1467 423 -1466
rect 467 -1467 829 -1466
rect 887 -1467 899 -1466
rect 905 -1467 913 -1466
rect 100 -1469 412 -1468
rect 422 -1469 479 -1468
rect 485 -1469 608 -1468
rect 611 -1469 661 -1468
rect 688 -1469 710 -1468
rect 712 -1469 815 -1468
rect 912 -1469 934 -1468
rect 65 -1471 661 -1470
rect 688 -1471 794 -1470
rect 65 -1473 73 -1472
rect 117 -1473 150 -1472
rect 156 -1473 738 -1472
rect 793 -1473 843 -1472
rect 86 -1475 157 -1474
rect 159 -1475 626 -1474
rect 632 -1475 636 -1474
rect 653 -1475 892 -1474
rect 86 -1477 195 -1476
rect 201 -1477 269 -1476
rect 352 -1477 465 -1476
rect 467 -1477 696 -1476
rect 730 -1477 745 -1476
rect 821 -1477 892 -1476
rect 107 -1479 465 -1478
rect 471 -1479 556 -1478
rect 590 -1479 682 -1478
rect 695 -1479 724 -1478
rect 737 -1479 951 -1478
rect 58 -1481 472 -1480
rect 478 -1481 773 -1480
rect 842 -1481 920 -1480
rect 58 -1483 234 -1482
rect 240 -1483 346 -1482
rect 355 -1483 451 -1482
rect 485 -1483 542 -1482
rect 597 -1483 605 -1482
rect 625 -1483 657 -1482
rect 681 -1483 703 -1482
rect 723 -1483 752 -1482
rect 765 -1483 773 -1482
rect 919 -1483 955 -1482
rect 121 -1485 304 -1484
rect 324 -1485 542 -1484
rect 597 -1485 640 -1484
rect 653 -1485 717 -1484
rect 744 -1485 759 -1484
rect 933 -1485 955 -1484
rect 128 -1487 507 -1486
rect 509 -1487 675 -1486
rect 702 -1487 836 -1486
rect 135 -1489 381 -1488
rect 443 -1489 717 -1488
rect 751 -1489 787 -1488
rect 835 -1489 850 -1488
rect 40 -1491 850 -1490
rect 142 -1493 181 -1492
rect 184 -1493 332 -1492
rect 366 -1493 409 -1492
rect 443 -1493 521 -1492
rect 537 -1493 822 -1492
rect 149 -1495 255 -1494
rect 261 -1495 325 -1494
rect 369 -1495 766 -1494
rect 786 -1495 808 -1494
rect 163 -1497 171 -1496
rect 173 -1497 360 -1496
rect 492 -1497 514 -1496
rect 537 -1497 815 -1496
rect 30 -1499 164 -1498
rect 184 -1499 388 -1498
rect 492 -1499 528 -1498
rect 618 -1499 640 -1498
rect 667 -1499 675 -1498
rect 807 -1499 878 -1498
rect 30 -1501 290 -1500
rect 359 -1501 619 -1500
rect 646 -1501 668 -1500
rect 152 -1503 647 -1502
rect 187 -1505 248 -1504
rect 261 -1505 594 -1504
rect 187 -1507 570 -1506
rect 191 -1509 255 -1508
rect 289 -1509 447 -1508
rect 562 -1509 570 -1508
rect 191 -1511 307 -1510
rect 401 -1511 528 -1510
rect 562 -1511 584 -1510
rect 205 -1513 248 -1512
rect 401 -1513 437 -1512
rect 583 -1513 885 -1512
rect 166 -1515 437 -1514
rect 177 -1517 206 -1516
rect 219 -1517 227 -1516
rect 233 -1517 454 -1516
rect 177 -1519 269 -1518
rect 219 -1521 297 -1520
rect 240 -1523 430 -1522
rect 275 -1525 297 -1524
rect 2 -1527 276 -1526
rect 23 -1538 41 -1537
rect 44 -1538 164 -1537
rect 166 -1538 290 -1537
rect 306 -1538 374 -1537
rect 432 -1538 486 -1537
rect 509 -1538 843 -1537
rect 849 -1538 927 -1537
rect 947 -1538 969 -1537
rect 982 -1538 990 -1537
rect 30 -1540 293 -1539
rect 345 -1540 367 -1539
rect 373 -1540 402 -1539
rect 436 -1540 853 -1539
rect 884 -1540 941 -1539
rect 954 -1540 972 -1539
rect 16 -1542 31 -1541
rect 37 -1542 276 -1541
rect 282 -1542 286 -1541
rect 352 -1542 465 -1541
rect 478 -1542 591 -1541
rect 604 -1542 871 -1541
rect 898 -1542 916 -1541
rect 940 -1542 976 -1541
rect 16 -1544 349 -1543
rect 352 -1544 381 -1543
rect 401 -1544 647 -1543
rect 705 -1544 773 -1543
rect 800 -1544 850 -1543
rect 898 -1544 913 -1543
rect 37 -1546 97 -1545
rect 100 -1546 139 -1545
rect 149 -1546 458 -1545
rect 478 -1546 493 -1545
rect 520 -1546 524 -1545
rect 534 -1546 731 -1545
rect 733 -1546 808 -1545
rect 814 -1546 843 -1545
rect 44 -1548 129 -1547
rect 135 -1548 360 -1547
rect 436 -1548 482 -1547
rect 485 -1548 528 -1547
rect 586 -1548 717 -1547
rect 814 -1548 906 -1547
rect 9 -1550 482 -1549
rect 492 -1550 633 -1549
rect 646 -1550 696 -1549
rect 716 -1550 752 -1549
rect 65 -1552 409 -1551
rect 446 -1552 710 -1551
rect 751 -1552 892 -1551
rect 65 -1554 185 -1553
rect 194 -1554 598 -1553
rect 604 -1554 654 -1553
rect 709 -1554 829 -1553
rect 86 -1556 367 -1555
rect 408 -1556 472 -1555
rect 520 -1556 577 -1555
rect 590 -1556 689 -1555
rect 86 -1558 111 -1557
rect 114 -1558 500 -1557
rect 555 -1558 598 -1557
rect 618 -1558 955 -1557
rect 93 -1560 444 -1559
rect 450 -1560 738 -1559
rect 100 -1562 304 -1561
rect 341 -1562 829 -1561
rect 107 -1564 346 -1563
rect 369 -1564 444 -1563
rect 453 -1564 745 -1563
rect 58 -1566 454 -1565
rect 457 -1566 514 -1565
rect 530 -1566 556 -1565
rect 632 -1566 661 -1565
rect 688 -1566 703 -1565
rect 744 -1566 836 -1565
rect 58 -1568 696 -1567
rect 702 -1568 920 -1567
rect 128 -1570 332 -1569
rect 411 -1570 654 -1569
rect 660 -1570 682 -1569
rect 880 -1570 920 -1569
rect 135 -1572 206 -1571
rect 212 -1572 248 -1571
rect 261 -1572 276 -1571
rect 282 -1572 325 -1571
rect 331 -1572 468 -1571
rect 513 -1572 549 -1571
rect 75 -1574 262 -1573
rect 289 -1574 472 -1573
rect 534 -1574 682 -1573
rect 149 -1576 360 -1575
rect 429 -1576 500 -1575
rect 548 -1576 563 -1575
rect 156 -1578 255 -1577
rect 303 -1578 318 -1577
rect 324 -1578 542 -1577
rect 562 -1578 766 -1577
rect 156 -1580 794 -1579
rect 159 -1582 255 -1581
rect 317 -1582 395 -1581
rect 429 -1582 566 -1581
rect 765 -1582 822 -1581
rect 72 -1584 395 -1583
rect 793 -1584 857 -1583
rect 72 -1586 241 -1585
rect 247 -1586 297 -1585
rect 362 -1586 857 -1585
rect 177 -1588 612 -1587
rect 177 -1590 675 -1589
rect 198 -1592 269 -1591
rect 296 -1592 339 -1591
rect 362 -1592 423 -1591
rect 569 -1592 612 -1591
rect 674 -1592 780 -1591
rect 173 -1594 269 -1593
rect 338 -1594 626 -1593
rect 201 -1596 220 -1595
rect 240 -1596 538 -1595
rect 569 -1596 640 -1595
rect 215 -1598 227 -1597
rect 387 -1598 542 -1597
rect 639 -1598 668 -1597
rect 226 -1600 311 -1599
rect 506 -1600 626 -1599
rect 667 -1600 801 -1599
rect 233 -1602 311 -1601
rect 506 -1602 584 -1601
rect 51 -1604 234 -1603
rect 523 -1604 577 -1603
rect 51 -1606 80 -1605
rect 537 -1606 787 -1605
rect 26 -1608 787 -1607
rect 79 -1610 122 -1609
rect 121 -1612 759 -1611
rect 9 -1623 24 -1622
rect 30 -1623 122 -1622
rect 124 -1623 682 -1622
rect 695 -1623 941 -1622
rect 943 -1623 962 -1622
rect 971 -1623 976 -1622
rect 9 -1625 241 -1624
rect 247 -1625 251 -1624
rect 289 -1625 388 -1624
rect 390 -1625 738 -1624
rect 793 -1625 850 -1624
rect 877 -1625 899 -1624
rect 912 -1625 920 -1624
rect 975 -1625 983 -1624
rect 16 -1627 188 -1626
rect 240 -1627 297 -1626
rect 299 -1627 654 -1626
rect 660 -1627 668 -1626
rect 712 -1627 766 -1626
rect 835 -1627 857 -1626
rect 894 -1627 927 -1626
rect 16 -1629 62 -1628
rect 93 -1629 626 -1628
rect 639 -1629 864 -1628
rect 926 -1629 948 -1628
rect 23 -1631 97 -1630
rect 100 -1631 185 -1630
rect 247 -1631 311 -1630
rect 341 -1631 706 -1630
rect 723 -1631 731 -1630
rect 842 -1631 888 -1630
rect 30 -1633 297 -1632
rect 303 -1633 339 -1632
rect 341 -1633 633 -1632
rect 660 -1633 745 -1632
rect 828 -1633 843 -1632
rect 37 -1635 59 -1634
rect 93 -1635 118 -1634
rect 163 -1635 626 -1634
rect 667 -1635 752 -1634
rect 37 -1637 423 -1636
rect 439 -1637 619 -1636
rect 716 -1637 745 -1636
rect 44 -1639 206 -1638
rect 250 -1639 311 -1638
rect 331 -1639 633 -1638
rect 44 -1641 52 -1640
rect 58 -1641 87 -1640
rect 107 -1641 227 -1640
rect 303 -1641 398 -1640
rect 404 -1641 766 -1640
rect 51 -1643 213 -1642
rect 226 -1643 346 -1642
rect 348 -1643 374 -1642
rect 383 -1643 731 -1642
rect 86 -1645 104 -1644
rect 110 -1645 325 -1644
rect 359 -1645 367 -1644
rect 387 -1645 430 -1644
rect 450 -1645 724 -1644
rect 128 -1647 213 -1646
rect 282 -1647 325 -1646
rect 352 -1647 367 -1646
rect 429 -1647 458 -1646
rect 464 -1647 703 -1646
rect 65 -1649 353 -1648
rect 401 -1649 458 -1648
rect 464 -1649 682 -1648
rect 65 -1651 80 -1650
rect 128 -1651 181 -1650
rect 282 -1651 409 -1650
rect 450 -1651 780 -1650
rect 135 -1653 206 -1652
rect 317 -1653 346 -1652
rect 401 -1653 773 -1652
rect 135 -1655 150 -1654
rect 163 -1655 192 -1654
rect 219 -1655 318 -1654
rect 331 -1655 703 -1654
rect 72 -1657 192 -1656
rect 408 -1657 416 -1656
rect 453 -1657 710 -1656
rect 145 -1659 423 -1658
rect 471 -1659 654 -1658
rect 149 -1661 759 -1660
rect 166 -1663 269 -1662
rect 471 -1663 514 -1662
rect 527 -1663 675 -1662
rect 170 -1665 178 -1664
rect 198 -1665 416 -1664
rect 478 -1665 493 -1664
rect 495 -1665 689 -1664
rect 173 -1667 220 -1666
rect 254 -1667 514 -1666
rect 527 -1667 549 -1666
rect 555 -1667 717 -1666
rect 173 -1669 185 -1668
rect 198 -1669 209 -1668
rect 254 -1669 262 -1668
rect 268 -1669 426 -1668
rect 488 -1669 955 -1668
rect 79 -1671 209 -1670
rect 261 -1671 276 -1670
rect 492 -1671 500 -1670
rect 506 -1671 549 -1670
rect 555 -1671 577 -1670
rect 586 -1671 696 -1670
rect 233 -1673 276 -1672
rect 499 -1673 521 -1672
rect 534 -1673 801 -1672
rect 156 -1675 535 -1674
rect 537 -1675 829 -1674
rect 142 -1677 157 -1676
rect 509 -1677 871 -1676
rect 142 -1679 577 -1678
rect 590 -1679 759 -1678
rect 786 -1679 801 -1678
rect 814 -1679 871 -1678
rect 485 -1681 787 -1680
rect 541 -1683 815 -1682
rect 520 -1685 542 -1684
rect 544 -1685 647 -1684
rect 562 -1687 605 -1686
rect 611 -1687 675 -1686
rect 152 -1689 612 -1688
rect 443 -1691 605 -1690
rect 436 -1693 444 -1692
rect 481 -1693 563 -1692
rect 565 -1693 640 -1692
rect 380 -1695 437 -1694
rect 569 -1695 822 -1694
rect 569 -1697 689 -1696
rect 583 -1699 647 -1698
rect 572 -1701 584 -1700
rect 590 -1701 734 -1700
rect 597 -1703 752 -1702
rect 394 -1705 598 -1704
rect 16 -1716 59 -1715
rect 72 -1716 76 -1715
rect 79 -1716 496 -1715
rect 506 -1716 549 -1715
rect 572 -1716 864 -1715
rect 905 -1716 913 -1715
rect 926 -1716 941 -1715
rect 961 -1716 979 -1715
rect 16 -1718 346 -1717
rect 355 -1718 773 -1717
rect 37 -1720 395 -1719
rect 397 -1720 430 -1719
rect 436 -1720 689 -1719
rect 709 -1720 759 -1719
rect 37 -1722 510 -1721
rect 523 -1722 703 -1721
rect 51 -1724 342 -1723
rect 376 -1724 731 -1723
rect 58 -1726 66 -1725
rect 93 -1726 388 -1725
rect 439 -1726 787 -1725
rect 9 -1728 66 -1727
rect 103 -1728 458 -1727
rect 467 -1728 815 -1727
rect 9 -1730 374 -1729
rect 387 -1730 409 -1729
rect 450 -1730 822 -1729
rect 86 -1732 104 -1731
rect 117 -1732 535 -1731
rect 548 -1732 556 -1731
rect 642 -1732 871 -1731
rect 23 -1734 118 -1733
rect 121 -1734 150 -1733
rect 159 -1734 738 -1733
rect 23 -1736 188 -1735
rect 191 -1736 206 -1735
rect 222 -1736 384 -1735
rect 450 -1736 479 -1735
rect 485 -1736 493 -1735
rect 534 -1736 591 -1735
rect 667 -1736 759 -1735
rect 82 -1738 87 -1737
rect 124 -1738 570 -1737
rect 702 -1738 766 -1737
rect 128 -1740 591 -1739
rect 730 -1740 801 -1739
rect 142 -1742 661 -1741
rect 737 -1742 829 -1741
rect 163 -1744 171 -1743
rect 173 -1744 262 -1743
rect 268 -1744 335 -1743
rect 471 -1744 486 -1743
rect 488 -1744 668 -1743
rect 166 -1746 423 -1745
rect 474 -1746 717 -1745
rect 170 -1748 409 -1747
rect 422 -1748 888 -1747
rect 191 -1750 248 -1749
rect 261 -1750 304 -1749
rect 310 -1750 377 -1749
rect 478 -1750 528 -1749
rect 555 -1750 612 -1749
rect 660 -1750 724 -1749
rect 107 -1752 304 -1751
rect 324 -1752 346 -1751
rect 527 -1752 577 -1751
rect 716 -1752 843 -1751
rect 107 -1754 136 -1753
rect 156 -1754 248 -1753
rect 271 -1754 836 -1753
rect 30 -1756 157 -1755
rect 219 -1756 311 -1755
rect 324 -1756 339 -1755
rect 576 -1756 626 -1755
rect 723 -1756 780 -1755
rect 30 -1758 52 -1757
rect 219 -1758 430 -1757
rect 625 -1758 696 -1757
rect 226 -1760 542 -1759
rect 695 -1760 745 -1759
rect 114 -1762 227 -1761
rect 233 -1762 416 -1761
rect 541 -1762 598 -1761
rect 639 -1762 745 -1761
rect 198 -1764 234 -1763
rect 236 -1764 612 -1763
rect 198 -1766 321 -1765
rect 338 -1766 367 -1765
rect 415 -1766 521 -1765
rect 597 -1766 647 -1765
rect 240 -1768 402 -1767
rect 443 -1768 647 -1767
rect 44 -1770 444 -1769
rect 44 -1772 500 -1771
rect 240 -1774 370 -1773
rect 499 -1774 654 -1773
rect 254 -1776 640 -1775
rect 653 -1776 752 -1775
rect 184 -1778 255 -1777
rect 275 -1778 689 -1777
rect 184 -1780 360 -1779
rect 583 -1780 752 -1779
rect 212 -1782 276 -1781
rect 282 -1782 465 -1781
rect 583 -1782 619 -1781
rect 93 -1784 213 -1783
rect 282 -1784 454 -1783
rect 464 -1784 514 -1783
rect 618 -1784 682 -1783
rect 289 -1786 458 -1785
rect 562 -1786 682 -1785
rect 180 -1788 290 -1787
rect 296 -1788 332 -1787
rect 352 -1788 563 -1787
rect 296 -1790 381 -1789
rect 401 -1790 514 -1789
rect 299 -1792 472 -1791
rect 317 -1794 332 -1793
rect 359 -1794 605 -1793
rect 604 -1796 675 -1795
rect 632 -1798 675 -1797
rect 352 -1800 633 -1799
rect 9 -1811 31 -1810
rect 33 -1811 38 -1810
rect 40 -1811 83 -1810
rect 89 -1811 423 -1810
rect 471 -1811 479 -1810
rect 492 -1811 759 -1810
rect 23 -1813 87 -1812
rect 93 -1813 213 -1812
rect 219 -1813 276 -1812
rect 306 -1813 339 -1812
rect 345 -1813 356 -1812
rect 366 -1813 377 -1812
rect 380 -1813 556 -1812
rect 579 -1813 738 -1812
rect 44 -1815 479 -1814
rect 492 -1815 500 -1814
rect 506 -1815 605 -1814
rect 674 -1815 678 -1814
rect 737 -1815 752 -1814
rect 51 -1817 108 -1816
rect 121 -1817 332 -1816
rect 348 -1817 689 -1816
rect 65 -1819 216 -1818
rect 219 -1819 283 -1818
rect 331 -1819 465 -1818
rect 495 -1819 752 -1818
rect 65 -1821 234 -1820
rect 240 -1821 503 -1820
rect 513 -1821 528 -1820
rect 604 -1821 612 -1820
rect 653 -1821 689 -1820
rect 72 -1823 223 -1822
rect 240 -1823 297 -1822
rect 352 -1823 423 -1822
rect 464 -1823 535 -1822
rect 611 -1823 619 -1822
rect 674 -1823 682 -1822
rect 72 -1825 143 -1824
rect 149 -1825 178 -1824
rect 184 -1825 192 -1824
rect 201 -1825 395 -1824
rect 415 -1825 507 -1824
rect 516 -1825 731 -1824
rect 47 -1827 416 -1826
rect 453 -1827 535 -1826
rect 618 -1827 633 -1826
rect 681 -1827 710 -1826
rect 79 -1829 115 -1828
rect 121 -1829 192 -1828
rect 268 -1829 591 -1828
rect 695 -1829 710 -1828
rect 93 -1831 500 -1830
rect 509 -1831 633 -1830
rect 695 -1831 717 -1830
rect 103 -1833 290 -1832
rect 296 -1833 304 -1832
rect 338 -1833 731 -1832
rect 107 -1835 199 -1834
rect 275 -1835 444 -1834
rect 520 -1835 549 -1834
rect 590 -1835 626 -1834
rect 677 -1835 717 -1834
rect 100 -1837 199 -1836
rect 282 -1837 486 -1836
rect 625 -1837 661 -1836
rect 124 -1839 528 -1838
rect 642 -1839 661 -1838
rect 128 -1841 248 -1840
rect 352 -1841 654 -1840
rect 135 -1843 437 -1842
rect 443 -1843 542 -1842
rect 142 -1845 255 -1844
rect 355 -1845 570 -1844
rect 156 -1847 206 -1846
rect 247 -1847 262 -1846
rect 310 -1847 570 -1846
rect 16 -1849 206 -1848
rect 254 -1849 363 -1848
rect 369 -1849 598 -1848
rect 16 -1851 293 -1850
rect 310 -1851 325 -1850
rect 359 -1851 381 -1850
rect 387 -1851 395 -1850
rect 450 -1851 598 -1850
rect 163 -1853 563 -1852
rect 12 -1855 563 -1854
rect 131 -1857 164 -1856
rect 166 -1857 556 -1856
rect 170 -1859 234 -1858
rect 261 -1859 402 -1858
rect 485 -1859 748 -1858
rect 135 -1861 171 -1860
rect 173 -1861 402 -1860
rect 187 -1863 227 -1862
rect 268 -1863 451 -1862
rect 114 -1865 227 -1864
rect 324 -1865 542 -1864
rect 373 -1867 703 -1866
rect 303 -1869 374 -1868
rect 387 -1869 584 -1868
rect 390 -1871 647 -1870
rect 180 -1873 647 -1872
rect 408 -1875 703 -1874
rect 408 -1877 430 -1876
rect 576 -1877 584 -1876
rect 317 -1879 430 -1878
rect 138 -1881 318 -1880
rect 2 -1892 73 -1891
rect 107 -1892 171 -1891
rect 177 -1892 192 -1891
rect 194 -1892 416 -1891
rect 432 -1892 738 -1891
rect 5 -1894 199 -1893
rect 201 -1894 370 -1893
rect 376 -1894 647 -1893
rect 709 -1894 748 -1893
rect 9 -1896 388 -1895
rect 397 -1896 556 -1895
rect 12 -1898 171 -1897
rect 177 -1898 227 -1897
rect 240 -1898 328 -1897
rect 338 -1898 535 -1897
rect 541 -1898 556 -1897
rect 23 -1900 234 -1899
rect 292 -1900 570 -1899
rect 23 -1902 465 -1901
rect 471 -1902 549 -1901
rect 562 -1902 570 -1901
rect 33 -1904 38 -1903
rect 44 -1904 269 -1903
rect 296 -1904 307 -1903
rect 317 -1904 419 -1903
rect 436 -1904 598 -1903
rect 26 -1906 269 -1905
rect 296 -1906 325 -1905
rect 345 -1906 703 -1905
rect 51 -1908 150 -1907
rect 156 -1908 304 -1907
rect 324 -1908 507 -1907
rect 520 -1908 535 -1907
rect 541 -1908 591 -1907
rect 597 -1908 633 -1907
rect 674 -1908 703 -1907
rect 51 -1910 59 -1909
rect 61 -1910 80 -1909
rect 117 -1910 157 -1909
rect 184 -1910 223 -1909
rect 254 -1910 318 -1909
rect 359 -1910 563 -1909
rect 590 -1910 661 -1909
rect 667 -1910 675 -1909
rect 65 -1912 167 -1911
rect 184 -1912 220 -1911
rect 303 -1912 461 -1911
rect 471 -1912 482 -1911
rect 502 -1912 724 -1911
rect 65 -1914 283 -1913
rect 331 -1914 360 -1913
rect 362 -1914 367 -1913
rect 380 -1914 521 -1913
rect 625 -1914 661 -1913
rect 16 -1916 283 -1915
rect 366 -1916 647 -1915
rect 72 -1918 580 -1917
rect 618 -1918 626 -1917
rect 639 -1918 724 -1917
rect 79 -1920 500 -1919
rect 506 -1920 528 -1919
rect 618 -1920 752 -1919
rect 19 -1922 528 -1921
rect 114 -1924 255 -1923
rect 261 -1924 332 -1923
rect 380 -1924 395 -1923
rect 401 -1924 577 -1923
rect 100 -1926 262 -1925
rect 355 -1926 395 -1925
rect 401 -1926 423 -1925
rect 429 -1926 668 -1925
rect 100 -1928 633 -1927
rect 128 -1930 311 -1929
rect 429 -1930 468 -1929
rect 131 -1932 654 -1931
rect 145 -1934 374 -1933
rect 436 -1934 486 -1933
rect 205 -1936 290 -1935
rect 310 -1936 458 -1935
rect 485 -1936 514 -1935
rect 149 -1938 206 -1937
rect 208 -1938 731 -1937
rect 142 -1940 731 -1939
rect 86 -1942 143 -1941
rect 212 -1942 241 -1941
rect 271 -1942 654 -1941
rect 86 -1944 136 -1943
rect 163 -1944 213 -1943
rect 219 -1944 234 -1943
rect 352 -1944 514 -1943
rect 135 -1946 409 -1945
rect 439 -1946 710 -1945
rect 275 -1948 409 -1947
rect 443 -1948 493 -1947
rect 247 -1950 276 -1949
rect 422 -1950 493 -1949
rect 93 -1952 248 -1951
rect 450 -1952 689 -1951
rect 37 -1954 689 -1953
rect 93 -1956 349 -1955
rect 450 -1956 479 -1955
rect 478 -1958 717 -1957
rect 695 -1960 717 -1959
rect 681 -1962 696 -1961
rect 54 -1964 682 -1963
rect 16 -1975 143 -1974
rect 156 -1975 262 -1974
rect 285 -1975 633 -1974
rect 635 -1975 717 -1974
rect 19 -1977 332 -1976
rect 366 -1977 591 -1976
rect 642 -1977 696 -1976
rect 23 -1979 206 -1978
rect 240 -1979 314 -1978
rect 324 -1979 440 -1978
rect 450 -1979 489 -1978
rect 534 -1979 549 -1978
rect 551 -1979 661 -1978
rect 695 -1979 724 -1978
rect 23 -1981 31 -1980
rect 37 -1981 76 -1980
rect 100 -1981 360 -1980
rect 366 -1981 552 -1980
rect 562 -1981 640 -1980
rect 30 -1983 108 -1982
rect 110 -1983 160 -1982
rect 163 -1983 325 -1982
rect 331 -1983 398 -1982
rect 404 -1983 472 -1982
rect 478 -1983 633 -1982
rect 44 -1985 433 -1984
rect 443 -1985 451 -1984
rect 457 -1985 584 -1984
rect 618 -1985 661 -1984
rect 44 -1987 87 -1986
rect 93 -1987 164 -1986
rect 170 -1987 297 -1986
rect 303 -1987 311 -1986
rect 369 -1987 668 -1986
rect 51 -1989 689 -1988
rect 58 -1991 104 -1990
rect 107 -1991 136 -1990
rect 142 -1991 213 -1990
rect 219 -1991 297 -1990
rect 387 -1991 570 -1990
rect 583 -1991 647 -1990
rect 65 -1993 80 -1992
rect 100 -1993 710 -1992
rect 2 -1995 66 -1994
rect 68 -1995 157 -1994
rect 177 -1995 209 -1994
rect 215 -1995 647 -1994
rect 72 -1997 90 -1996
rect 117 -1997 500 -1996
rect 534 -1997 682 -1996
rect 117 -1999 136 -1998
rect 149 -1999 171 -1998
rect 177 -1999 185 -1998
rect 191 -1999 241 -1998
rect 254 -1999 269 -1998
rect 289 -1999 353 -1998
rect 387 -1999 409 -1998
rect 415 -1999 591 -1998
rect 604 -1999 619 -1998
rect 9 -2001 150 -2000
rect 184 -2001 556 -2000
rect 562 -2001 598 -2000
rect 604 -2001 675 -2000
rect 9 -2003 174 -2002
rect 219 -2003 234 -2002
rect 247 -2003 269 -2002
rect 289 -2003 339 -2002
rect 380 -2003 416 -2002
rect 418 -2003 507 -2002
rect 569 -2003 654 -2002
rect 54 -2005 339 -2004
rect 394 -2005 402 -2004
rect 408 -2005 437 -2004
rect 443 -2005 514 -2004
rect 597 -2005 731 -2004
rect 54 -2007 500 -2006
rect 506 -2007 577 -2006
rect 642 -2007 654 -2006
rect 121 -2009 202 -2008
rect 226 -2009 248 -2008
rect 261 -2009 276 -2008
rect 422 -2009 482 -2008
rect 513 -2009 542 -2008
rect 576 -2009 626 -2008
rect 128 -2011 360 -2010
rect 457 -2011 486 -2010
rect 541 -2011 612 -2010
rect 625 -2011 650 -2010
rect 121 -2013 129 -2012
rect 131 -2013 307 -2012
rect 464 -2013 521 -2012
rect 611 -2013 703 -2012
rect 226 -2015 374 -2014
rect 474 -2015 556 -2014
rect 233 -2017 346 -2016
rect 373 -2017 430 -2016
rect 492 -2017 521 -2016
rect 275 -2019 318 -2018
rect 429 -2019 528 -2018
rect 282 -2021 318 -2020
rect 348 -2021 528 -2020
rect 282 -2023 465 -2022
rect 303 -2025 346 -2024
rect 436 -2025 493 -2024
rect 9 -2036 202 -2035
rect 212 -2036 430 -2035
rect 436 -2036 626 -2035
rect 632 -2036 640 -2035
rect 646 -2036 661 -2035
rect 688 -2036 696 -2035
rect 16 -2038 97 -2037
rect 114 -2038 290 -2037
rect 303 -2038 353 -2037
rect 380 -2038 444 -2037
rect 474 -2038 514 -2037
rect 520 -2038 542 -2037
rect 548 -2038 584 -2037
rect 16 -2040 129 -2039
rect 191 -2040 388 -2039
rect 415 -2040 535 -2039
rect 541 -2040 563 -2039
rect 30 -2042 118 -2041
rect 128 -2042 136 -2041
rect 191 -2042 241 -2041
rect 257 -2042 262 -2041
rect 289 -2042 472 -2041
rect 481 -2042 570 -2041
rect 37 -2044 255 -2043
rect 303 -2044 437 -2043
rect 443 -2044 451 -2043
rect 471 -2044 507 -2043
rect 548 -2044 577 -2043
rect 33 -2046 38 -2045
rect 44 -2046 87 -2045
rect 100 -2046 115 -2045
rect 117 -2046 185 -2045
rect 198 -2046 405 -2045
rect 425 -2046 598 -2045
rect 44 -2048 143 -2047
rect 194 -2048 199 -2047
rect 205 -2048 262 -2047
rect 313 -2048 577 -2047
rect 51 -2050 73 -2049
rect 79 -2050 419 -2049
rect 429 -2050 479 -2049
rect 485 -2050 643 -2049
rect 51 -2052 97 -2051
rect 212 -2052 311 -2051
rect 320 -2052 514 -2051
rect 555 -2052 654 -2051
rect 65 -2054 500 -2053
rect 555 -2054 619 -2053
rect 642 -2054 675 -2053
rect 65 -2056 171 -2055
rect 215 -2056 671 -2055
rect 75 -2058 80 -2057
rect 86 -2058 108 -2057
rect 170 -2058 276 -2057
rect 327 -2058 346 -2057
rect 359 -2058 388 -2057
rect 418 -2058 584 -2057
rect 107 -2060 164 -2059
rect 219 -2060 528 -2059
rect 562 -2060 612 -2059
rect 58 -2062 220 -2061
rect 222 -2062 227 -2061
rect 236 -2062 570 -2061
rect 604 -2062 612 -2061
rect 58 -2064 90 -2063
rect 149 -2064 360 -2063
rect 383 -2064 409 -2063
rect 450 -2064 458 -2063
rect 492 -2064 507 -2063
rect 149 -2066 234 -2065
rect 240 -2066 325 -2065
rect 331 -2066 402 -2065
rect 408 -2066 528 -2065
rect 135 -2068 325 -2067
rect 338 -2068 493 -2067
rect 499 -2068 636 -2067
rect 156 -2070 458 -2069
rect 142 -2072 157 -2071
rect 159 -2072 164 -2071
rect 222 -2072 248 -2071
rect 254 -2072 374 -2071
rect 394 -2072 605 -2071
rect 226 -2074 370 -2073
rect 373 -2074 479 -2073
rect 268 -2076 339 -2075
rect 345 -2076 381 -2075
rect 394 -2076 423 -2075
rect 268 -2078 367 -2077
rect 401 -2078 465 -2077
rect 275 -2080 405 -2079
rect 317 -2082 332 -2081
rect 352 -2082 465 -2081
rect 317 -2084 535 -2083
rect 366 -2086 591 -2085
rect 282 -2088 591 -2087
rect 282 -2090 307 -2089
rect 23 -2101 59 -2100
rect 65 -2101 311 -2100
rect 324 -2101 346 -2100
rect 366 -2101 409 -2100
rect 509 -2101 521 -2100
rect 523 -2101 570 -2100
rect 590 -2101 598 -2100
rect 611 -2101 622 -2100
rect 642 -2101 647 -2100
rect 674 -2101 689 -2100
rect 26 -2103 76 -2102
rect 107 -2103 307 -2102
rect 310 -2103 339 -2102
rect 345 -2103 384 -2102
rect 394 -2103 402 -2102
rect 530 -2103 584 -2102
rect 611 -2103 619 -2102
rect 33 -2105 38 -2104
rect 44 -2105 318 -2104
rect 331 -2105 570 -2104
rect 37 -2107 129 -2106
rect 135 -2107 139 -2106
rect 156 -2107 178 -2106
rect 187 -2107 321 -2106
rect 338 -2107 381 -2106
rect 387 -2107 395 -2106
rect 534 -2107 556 -2106
rect 562 -2107 591 -2106
rect 44 -2109 185 -2108
rect 208 -2109 269 -2108
rect 282 -2109 353 -2108
rect 359 -2109 388 -2108
rect 464 -2109 535 -2108
rect 51 -2111 153 -2110
rect 163 -2111 206 -2110
rect 215 -2111 528 -2110
rect 51 -2113 199 -2112
rect 205 -2113 213 -2112
rect 222 -2113 503 -2112
rect 58 -2115 87 -2114
rect 107 -2115 122 -2114
rect 135 -2115 143 -2114
rect 149 -2115 164 -2114
rect 170 -2115 192 -2114
rect 198 -2115 290 -2114
rect 303 -2115 563 -2114
rect 65 -2117 80 -2116
rect 86 -2117 227 -2116
rect 233 -2117 241 -2116
rect 247 -2117 559 -2116
rect 16 -2119 80 -2118
rect 138 -2119 143 -2118
rect 170 -2119 265 -2118
rect 268 -2119 307 -2118
rect 369 -2119 605 -2118
rect 72 -2121 118 -2120
rect 177 -2121 479 -2120
rect 117 -2123 290 -2122
rect 233 -2125 276 -2124
rect 240 -2127 335 -2126
rect 247 -2129 444 -2128
rect 254 -2131 293 -2130
rect 443 -2131 451 -2130
rect 226 -2133 255 -2132
rect 261 -2133 276 -2132
rect 450 -2133 472 -2132
rect 261 -2135 514 -2134
rect 422 -2137 472 -2136
rect 513 -2137 549 -2136
rect 422 -2139 437 -2138
rect 492 -2139 549 -2138
rect 373 -2141 437 -2140
rect 492 -2141 507 -2140
rect 373 -2143 458 -2142
rect 457 -2145 486 -2144
rect 485 -2147 577 -2146
rect 9 -2158 20 -2157
rect 37 -2158 216 -2157
rect 240 -2158 283 -2157
rect 285 -2158 297 -2157
rect 317 -2158 409 -2157
rect 415 -2158 549 -2157
rect 590 -2158 605 -2157
rect 44 -2160 185 -2159
rect 208 -2160 290 -2159
rect 292 -2160 311 -2159
rect 317 -2160 388 -2159
rect 408 -2160 444 -2159
rect 450 -2160 468 -2159
rect 499 -2160 556 -2159
rect 597 -2160 601 -2159
rect 51 -2162 262 -2161
rect 275 -2162 304 -2161
rect 324 -2162 335 -2161
rect 352 -2162 360 -2161
rect 362 -2162 486 -2161
rect 541 -2162 556 -2161
rect 51 -2164 150 -2163
rect 163 -2164 188 -2163
rect 247 -2164 374 -2163
rect 387 -2164 423 -2163
rect 425 -2164 479 -2163
rect 58 -2166 97 -2165
rect 107 -2166 129 -2165
rect 131 -2166 136 -2165
rect 163 -2166 181 -2165
rect 268 -2166 304 -2165
rect 324 -2166 346 -2165
rect 352 -2166 570 -2165
rect 58 -2168 178 -2167
rect 278 -2168 349 -2167
rect 366 -2168 563 -2167
rect 65 -2170 73 -2169
rect 79 -2170 157 -2169
rect 177 -2170 339 -2169
rect 345 -2170 535 -2169
rect 40 -2172 73 -2171
rect 86 -2172 269 -2171
rect 296 -2172 465 -2171
rect 513 -2172 535 -2171
rect 65 -2174 220 -2173
rect 331 -2174 395 -2173
rect 415 -2174 521 -2173
rect 86 -2176 143 -2175
rect 156 -2176 171 -2175
rect 219 -2176 258 -2175
rect 394 -2176 482 -2175
rect 93 -2178 101 -2177
rect 107 -2178 129 -2177
rect 135 -2178 213 -2177
rect 429 -2178 444 -2177
rect 453 -2178 472 -2177
rect 93 -2180 139 -2179
rect 205 -2180 213 -2179
rect 429 -2180 493 -2179
rect 100 -2182 199 -2181
rect 380 -2182 493 -2181
rect 121 -2184 234 -2183
rect 380 -2184 402 -2183
rect 436 -2184 510 -2183
rect 121 -2186 132 -2185
rect 170 -2186 234 -2185
rect 436 -2186 458 -2185
rect 198 -2188 248 -2187
rect 457 -2188 500 -2187
rect 226 -2190 402 -2189
rect 191 -2192 227 -2191
rect 187 -2194 192 -2193
rect 9 -2205 17 -2204
rect 23 -2205 27 -2204
rect 51 -2205 104 -2204
rect 107 -2205 202 -2204
rect 240 -2205 381 -2204
rect 408 -2205 419 -2204
rect 429 -2205 451 -2204
rect 457 -2205 507 -2204
rect 534 -2205 549 -2204
rect 600 -2205 605 -2204
rect 51 -2207 83 -2206
rect 86 -2207 206 -2206
rect 254 -2207 465 -2206
rect 537 -2207 556 -2206
rect 58 -2209 129 -2208
rect 149 -2209 157 -2208
rect 177 -2209 206 -2208
rect 254 -2209 290 -2208
rect 299 -2209 363 -2208
rect 366 -2209 388 -2208
rect 394 -2209 409 -2208
rect 422 -2209 535 -2208
rect 58 -2211 94 -2210
rect 100 -2211 213 -2210
rect 247 -2211 290 -2210
rect 303 -2211 342 -2210
rect 359 -2211 521 -2210
rect 65 -2213 146 -2212
rect 149 -2213 164 -2212
rect 177 -2213 262 -2212
rect 268 -2213 349 -2212
rect 373 -2213 437 -2212
rect 443 -2213 493 -2212
rect 79 -2215 209 -2214
rect 247 -2215 318 -2214
rect 324 -2215 353 -2214
rect 107 -2217 171 -2216
rect 187 -2217 220 -2216
rect 268 -2217 346 -2216
rect 114 -2219 122 -2218
rect 191 -2219 283 -2218
rect 72 -2221 115 -2220
rect 191 -2221 227 -2220
rect 275 -2221 332 -2220
rect 226 -2223 328 -2222
rect 331 -2223 402 -2222
rect 58 -2234 94 -2233
rect 107 -2234 174 -2233
rect 201 -2234 269 -2233
rect 275 -2234 328 -2233
rect 331 -2234 384 -2233
rect 408 -2234 430 -2233
rect 450 -2234 475 -2233
rect 485 -2234 507 -2233
rect 75 -2236 115 -2235
rect 131 -2236 227 -2235
rect 240 -2236 391 -2235
rect 149 -2238 164 -2237
rect 219 -2238 283 -2237
rect 289 -2238 304 -2237
rect 310 -2238 374 -2237
rect 247 -2240 356 -2239
rect 254 -2242 314 -2241
<< m2contact >>
rect 131 0 132 1
rect 156 0 157 1
rect 163 0 164 1
rect 187 0 188 1
rect 191 0 192 1
rect 233 0 234 1
rect 261 0 262 1
rect 282 0 283 1
rect 177 -2 178 -1
rect 212 -2 213 -1
rect 215 -2 216 -1
rect 247 -2 248 -1
rect 268 -2 269 -1
rect 278 -2 279 -1
rect 226 -4 227 -3
rect 257 -4 258 -3
rect 86 -15 87 -14
rect 163 -15 164 -14
rect 170 -15 171 -14
rect 219 -15 220 -14
rect 240 -15 241 -14
rect 261 -15 262 -14
rect 268 -15 269 -14
rect 345 -15 346 -14
rect 369 -15 370 -14
rect 401 -15 402 -14
rect 93 -17 94 -16
rect 100 -17 101 -16
rect 107 -17 108 -16
rect 110 -17 111 -16
rect 142 -17 143 -16
rect 226 -17 227 -16
rect 247 -17 248 -16
rect 289 -17 290 -16
rect 327 -17 328 -16
rect 331 -17 332 -16
rect 376 -17 377 -16
rect 380 -17 381 -16
rect 110 -19 111 -18
rect 254 -19 255 -18
rect 257 -19 258 -18
rect 387 -19 388 -18
rect 138 -21 139 -20
rect 142 -21 143 -20
rect 149 -21 150 -20
rect 166 -21 167 -20
rect 170 -21 171 -20
rect 177 -21 178 -20
rect 180 -21 181 -20
rect 233 -21 234 -20
rect 243 -21 244 -20
rect 247 -21 248 -20
rect 275 -21 276 -20
rect 418 -21 419 -20
rect 156 -23 157 -22
rect 177 -23 178 -22
rect 184 -23 185 -22
rect 212 -23 213 -22
rect 215 -23 216 -22
rect 296 -23 297 -22
rect 117 -25 118 -24
rect 156 -25 157 -24
rect 191 -25 192 -24
rect 352 -25 353 -24
rect 128 -27 129 -26
rect 191 -27 192 -26
rect 198 -27 199 -26
rect 303 -27 304 -26
rect 198 -29 199 -28
rect 208 -29 209 -28
rect 222 -29 223 -28
rect 261 -29 262 -28
rect 282 -29 283 -28
rect 359 -29 360 -28
rect 205 -31 206 -30
rect 268 -31 269 -30
rect 282 -31 283 -30
rect 317 -31 318 -30
rect 65 -42 66 -41
rect 93 -42 94 -41
rect 100 -42 101 -41
rect 184 -42 185 -41
rect 212 -42 213 -41
rect 359 -42 360 -41
rect 72 -44 73 -43
rect 128 -44 129 -43
rect 149 -44 150 -43
rect 180 -44 181 -43
rect 184 -44 185 -43
rect 198 -44 199 -43
rect 226 -44 227 -43
rect 373 -44 374 -43
rect 75 -46 76 -45
rect 149 -46 150 -45
rect 156 -46 157 -45
rect 198 -46 199 -45
rect 229 -46 230 -45
rect 261 -46 262 -45
rect 275 -46 276 -45
rect 278 -46 279 -45
rect 282 -46 283 -45
rect 408 -46 409 -45
rect 79 -48 80 -47
rect 215 -48 216 -47
rect 233 -48 234 -47
rect 313 -48 314 -47
rect 324 -48 325 -47
rect 387 -48 388 -47
rect 86 -50 87 -49
rect 222 -50 223 -49
rect 233 -50 234 -49
rect 240 -50 241 -49
rect 261 -50 262 -49
rect 268 -50 269 -49
rect 275 -50 276 -49
rect 317 -50 318 -49
rect 44 -52 45 -51
rect 86 -52 87 -51
rect 114 -52 115 -51
rect 156 -52 157 -51
rect 163 -52 164 -51
rect 212 -52 213 -51
rect 240 -52 241 -51
rect 247 -52 248 -51
rect 278 -52 279 -51
rect 317 -52 318 -51
rect 107 -54 108 -53
rect 114 -54 115 -53
rect 117 -54 118 -53
rect 173 -54 174 -53
rect 191 -54 192 -53
rect 247 -54 248 -53
rect 282 -54 283 -53
rect 380 -54 381 -53
rect 121 -56 122 -55
rect 177 -56 178 -55
rect 205 -56 206 -55
rect 380 -56 381 -55
rect 121 -58 122 -57
rect 135 -58 136 -57
rect 170 -58 171 -57
rect 359 -58 360 -57
rect 131 -60 132 -59
rect 387 -60 388 -59
rect 135 -62 136 -61
rect 142 -62 143 -61
rect 170 -62 171 -61
rect 401 -62 402 -61
rect 285 -64 286 -63
rect 345 -64 346 -63
rect 289 -66 290 -65
rect 310 -66 311 -65
rect 331 -66 332 -65
rect 401 -66 402 -65
rect 219 -68 220 -67
rect 289 -68 290 -67
rect 296 -68 297 -67
rect 324 -68 325 -67
rect 338 -68 339 -67
rect 345 -68 346 -67
rect 219 -70 220 -69
rect 366 -70 367 -69
rect 254 -72 255 -71
rect 296 -72 297 -71
rect 338 -72 339 -71
rect 394 -72 395 -71
rect 51 -74 52 -73
rect 254 -74 255 -73
rect 257 -74 258 -73
rect 331 -74 332 -73
rect 352 -74 353 -73
rect 394 -74 395 -73
rect 44 -85 45 -84
rect 100 -85 101 -84
rect 121 -85 122 -84
rect 135 -85 136 -84
rect 159 -85 160 -84
rect 191 -85 192 -84
rect 194 -85 195 -84
rect 226 -85 227 -84
rect 250 -85 251 -84
rect 401 -85 402 -84
rect 51 -87 52 -86
rect 156 -87 157 -86
rect 163 -87 164 -86
rect 170 -87 171 -86
rect 201 -87 202 -86
rect 247 -87 248 -86
rect 254 -87 255 -86
rect 303 -87 304 -86
rect 331 -87 332 -86
rect 383 -87 384 -86
rect 394 -87 395 -86
rect 443 -87 444 -86
rect 58 -89 59 -88
rect 145 -89 146 -88
rect 205 -89 206 -88
rect 240 -89 241 -88
rect 257 -89 258 -88
rect 373 -89 374 -88
rect 401 -89 402 -88
rect 453 -89 454 -88
rect 65 -91 66 -90
rect 114 -91 115 -90
rect 128 -91 129 -90
rect 394 -91 395 -90
rect 65 -93 66 -92
rect 79 -93 80 -92
rect 86 -93 87 -92
rect 107 -93 108 -92
rect 131 -93 132 -92
rect 289 -93 290 -92
rect 317 -93 318 -92
rect 331 -93 332 -92
rect 352 -93 353 -92
rect 408 -93 409 -92
rect 93 -95 94 -94
rect 124 -95 125 -94
rect 142 -95 143 -94
rect 163 -95 164 -94
rect 212 -95 213 -94
rect 261 -95 262 -94
rect 271 -95 272 -94
rect 387 -95 388 -94
rect 408 -95 409 -94
rect 432 -95 433 -94
rect 107 -97 108 -96
rect 247 -97 248 -96
rect 275 -97 276 -96
rect 282 -97 283 -96
rect 289 -97 290 -96
rect 359 -97 360 -96
rect 366 -97 367 -96
rect 415 -97 416 -96
rect 96 -99 97 -98
rect 359 -99 360 -98
rect 149 -101 150 -100
rect 373 -101 374 -100
rect 149 -103 150 -102
rect 184 -103 185 -102
rect 212 -103 213 -102
rect 219 -103 220 -102
rect 222 -103 223 -102
rect 422 -103 423 -102
rect 177 -105 178 -104
rect 261 -105 262 -104
rect 278 -105 279 -104
rect 380 -105 381 -104
rect 184 -107 185 -106
rect 191 -107 192 -106
rect 215 -107 216 -106
rect 324 -107 325 -106
rect 338 -107 339 -106
rect 387 -107 388 -106
rect 79 -109 80 -108
rect 215 -109 216 -108
rect 233 -109 234 -108
rect 254 -109 255 -108
rect 271 -109 272 -108
rect 338 -109 339 -108
rect 345 -109 346 -108
rect 352 -109 353 -108
rect 198 -111 199 -110
rect 345 -111 346 -110
rect 240 -113 241 -112
rect 429 -113 430 -112
rect 278 -115 279 -114
rect 303 -115 304 -114
rect 310 -115 311 -114
rect 324 -115 325 -114
rect 296 -117 297 -116
rect 317 -117 318 -116
rect 296 -119 297 -118
rect 366 -119 367 -118
rect 37 -130 38 -129
rect 149 -130 150 -129
rect 156 -130 157 -129
rect 198 -130 199 -129
rect 215 -130 216 -129
rect 429 -130 430 -129
rect 436 -130 437 -129
rect 481 -130 482 -129
rect 44 -132 45 -131
rect 93 -132 94 -131
rect 110 -132 111 -131
rect 114 -132 115 -131
rect 128 -132 129 -131
rect 205 -132 206 -131
rect 219 -132 220 -131
rect 222 -132 223 -131
rect 226 -132 227 -131
rect 250 -132 251 -131
rect 254 -132 255 -131
rect 268 -132 269 -131
rect 275 -132 276 -131
rect 450 -132 451 -131
rect 51 -134 52 -133
rect 166 -134 167 -133
rect 170 -134 171 -133
rect 429 -134 430 -133
rect 58 -136 59 -135
rect 142 -136 143 -135
rect 145 -136 146 -135
rect 226 -136 227 -135
rect 233 -136 234 -135
rect 236 -136 237 -135
rect 247 -136 248 -135
rect 338 -136 339 -135
rect 359 -136 360 -135
rect 366 -136 367 -135
rect 380 -136 381 -135
rect 471 -136 472 -135
rect 58 -138 59 -137
rect 166 -138 167 -137
rect 170 -138 171 -137
rect 191 -138 192 -137
rect 236 -138 237 -137
rect 415 -138 416 -137
rect 72 -140 73 -139
rect 121 -140 122 -139
rect 131 -140 132 -139
rect 422 -140 423 -139
rect 79 -142 80 -141
rect 93 -142 94 -141
rect 177 -142 178 -141
rect 198 -142 199 -141
rect 254 -142 255 -141
rect 464 -142 465 -141
rect 79 -144 80 -143
rect 121 -144 122 -143
rect 184 -144 185 -143
rect 247 -144 248 -143
rect 261 -144 262 -143
rect 285 -144 286 -143
rect 289 -144 290 -143
rect 380 -144 381 -143
rect 387 -144 388 -143
rect 485 -144 486 -143
rect 89 -146 90 -145
rect 100 -146 101 -145
rect 103 -146 104 -145
rect 177 -146 178 -145
rect 191 -146 192 -145
rect 324 -146 325 -145
rect 352 -146 353 -145
rect 359 -146 360 -145
rect 401 -146 402 -145
rect 457 -146 458 -145
rect 100 -148 101 -147
rect 107 -148 108 -147
rect 117 -148 118 -147
rect 324 -148 325 -147
rect 345 -148 346 -147
rect 352 -148 353 -147
rect 415 -148 416 -147
rect 443 -148 444 -147
rect 138 -150 139 -149
rect 184 -150 185 -149
rect 208 -150 209 -149
rect 401 -150 402 -149
rect 86 -152 87 -151
rect 138 -152 139 -151
rect 282 -152 283 -151
rect 338 -152 339 -151
rect 296 -154 297 -153
rect 313 -154 314 -153
rect 317 -154 318 -153
rect 492 -154 493 -153
rect 296 -156 297 -155
rect 387 -156 388 -155
rect 303 -158 304 -157
rect 345 -158 346 -157
rect 306 -160 307 -159
rect 443 -160 444 -159
rect 310 -162 311 -161
rect 408 -162 409 -161
rect 317 -164 318 -163
rect 408 -164 409 -163
rect 320 -166 321 -165
rect 394 -166 395 -165
rect 373 -168 374 -167
rect 394 -168 395 -167
rect 331 -170 332 -169
rect 373 -170 374 -169
rect 331 -172 332 -171
rect 439 -172 440 -171
rect 16 -183 17 -182
rect 89 -183 90 -182
rect 114 -183 115 -182
rect 152 -183 153 -182
rect 191 -183 192 -182
rect 285 -183 286 -182
rect 292 -183 293 -182
rect 373 -183 374 -182
rect 380 -183 381 -182
rect 555 -183 556 -182
rect 583 -183 584 -182
rect 639 -183 640 -182
rect 30 -185 31 -184
rect 222 -185 223 -184
rect 226 -185 227 -184
rect 478 -185 479 -184
rect 534 -185 535 -184
rect 548 -185 549 -184
rect 37 -187 38 -186
rect 208 -187 209 -186
rect 254 -187 255 -186
rect 334 -187 335 -186
rect 380 -187 381 -186
rect 565 -187 566 -186
rect 37 -189 38 -188
rect 79 -189 80 -188
rect 86 -189 87 -188
rect 107 -189 108 -188
rect 114 -189 115 -188
rect 341 -189 342 -188
rect 387 -189 388 -188
rect 548 -189 549 -188
rect 44 -191 45 -190
rect 145 -191 146 -190
rect 191 -191 192 -190
rect 233 -191 234 -190
rect 257 -191 258 -190
rect 268 -191 269 -190
rect 275 -191 276 -190
rect 338 -191 339 -190
rect 366 -191 367 -190
rect 387 -191 388 -190
rect 464 -191 465 -190
rect 499 -191 500 -190
rect 51 -193 52 -192
rect 289 -193 290 -192
rect 296 -193 297 -192
rect 324 -193 325 -192
rect 450 -193 451 -192
rect 464 -193 465 -192
rect 471 -193 472 -192
rect 506 -193 507 -192
rect 58 -195 59 -194
rect 527 -195 528 -194
rect 58 -197 59 -196
rect 93 -197 94 -196
rect 121 -197 122 -196
rect 247 -197 248 -196
rect 261 -197 262 -196
rect 289 -197 290 -196
rect 306 -197 307 -196
rect 485 -197 486 -196
rect 65 -199 66 -198
rect 68 -199 69 -198
rect 72 -199 73 -198
rect 152 -199 153 -198
rect 156 -199 157 -198
rect 261 -199 262 -198
rect 278 -199 279 -198
rect 429 -199 430 -198
rect 443 -199 444 -198
rect 450 -199 451 -198
rect 457 -199 458 -198
rect 471 -199 472 -198
rect 79 -201 80 -200
rect 422 -201 423 -200
rect 436 -201 437 -200
rect 443 -201 444 -200
rect 89 -203 90 -202
rect 415 -203 416 -202
rect 103 -205 104 -204
rect 429 -205 430 -204
rect 121 -207 122 -206
rect 373 -207 374 -206
rect 408 -207 409 -206
rect 457 -207 458 -206
rect 124 -209 125 -208
rect 240 -209 241 -208
rect 243 -209 244 -208
rect 268 -209 269 -208
rect 282 -209 283 -208
rect 415 -209 416 -208
rect 128 -211 129 -210
rect 184 -211 185 -210
rect 187 -211 188 -210
rect 366 -211 367 -210
rect 408 -211 409 -210
rect 520 -211 521 -210
rect 82 -213 83 -212
rect 128 -213 129 -212
rect 135 -213 136 -212
rect 243 -213 244 -212
rect 317 -213 318 -212
rect 492 -213 493 -212
rect 135 -215 136 -214
rect 163 -215 164 -214
rect 170 -215 171 -214
rect 247 -215 248 -214
rect 324 -215 325 -214
rect 513 -215 514 -214
rect 142 -217 143 -216
rect 226 -217 227 -216
rect 233 -217 234 -216
rect 345 -217 346 -216
rect 401 -217 402 -216
rect 492 -217 493 -216
rect 96 -219 97 -218
rect 401 -219 402 -218
rect 142 -221 143 -220
rect 303 -221 304 -220
rect 331 -221 332 -220
rect 485 -221 486 -220
rect 170 -223 171 -222
rect 177 -223 178 -222
rect 198 -223 199 -222
rect 215 -223 216 -222
rect 310 -223 311 -222
rect 331 -223 332 -222
rect 345 -223 346 -222
rect 394 -223 395 -222
rect 156 -225 157 -224
rect 177 -225 178 -224
rect 198 -225 199 -224
rect 352 -225 353 -224
rect 359 -225 360 -224
rect 394 -225 395 -224
rect 205 -227 206 -226
rect 219 -227 220 -226
rect 359 -227 360 -226
rect 436 -227 437 -226
rect 149 -229 150 -228
rect 219 -229 220 -228
rect 16 -240 17 -239
rect 149 -240 150 -239
rect 180 -240 181 -239
rect 247 -240 248 -239
rect 285 -240 286 -239
rect 492 -240 493 -239
rect 499 -240 500 -239
rect 576 -240 577 -239
rect 586 -240 587 -239
rect 625 -240 626 -239
rect 639 -240 640 -239
rect 660 -240 661 -239
rect 30 -242 31 -241
rect 145 -242 146 -241
rect 205 -242 206 -241
rect 219 -242 220 -241
rect 240 -242 241 -241
rect 604 -242 605 -241
rect 30 -244 31 -243
rect 198 -244 199 -243
rect 205 -244 206 -243
rect 240 -244 241 -243
rect 243 -244 244 -243
rect 275 -244 276 -243
rect 278 -244 279 -243
rect 492 -244 493 -243
rect 506 -244 507 -243
rect 562 -244 563 -243
rect 44 -246 45 -245
rect 79 -246 80 -245
rect 82 -246 83 -245
rect 478 -246 479 -245
rect 481 -246 482 -245
rect 590 -246 591 -245
rect 51 -248 52 -247
rect 527 -248 528 -247
rect 534 -248 535 -247
rect 565 -248 566 -247
rect 58 -250 59 -249
rect 93 -250 94 -249
rect 103 -250 104 -249
rect 345 -250 346 -249
rect 352 -250 353 -249
rect 485 -250 486 -249
rect 513 -250 514 -249
rect 583 -250 584 -249
rect 72 -252 73 -251
rect 135 -252 136 -251
rect 156 -252 157 -251
rect 352 -252 353 -251
rect 362 -252 363 -251
rect 401 -252 402 -251
rect 408 -252 409 -251
rect 506 -252 507 -251
rect 555 -252 556 -251
rect 597 -252 598 -251
rect 86 -254 87 -253
rect 194 -254 195 -253
rect 198 -254 199 -253
rect 359 -254 360 -253
rect 366 -254 367 -253
rect 485 -254 486 -253
rect 558 -254 559 -253
rect 618 -254 619 -253
rect 93 -256 94 -255
rect 100 -256 101 -255
rect 124 -256 125 -255
rect 135 -256 136 -255
rect 156 -256 157 -255
rect 177 -256 178 -255
rect 212 -256 213 -255
rect 226 -256 227 -255
rect 247 -256 248 -255
rect 408 -256 409 -255
rect 422 -256 423 -255
rect 527 -256 528 -255
rect 100 -258 101 -257
rect 166 -258 167 -257
rect 226 -258 227 -257
rect 257 -258 258 -257
rect 268 -258 269 -257
rect 275 -258 276 -257
rect 285 -258 286 -257
rect 632 -258 633 -257
rect 254 -260 255 -259
rect 422 -260 423 -259
rect 429 -260 430 -259
rect 534 -260 535 -259
rect 268 -262 269 -261
rect 324 -262 325 -261
rect 331 -262 332 -261
rect 499 -262 500 -261
rect 233 -264 234 -263
rect 331 -264 332 -263
rect 338 -264 339 -263
rect 513 -264 514 -263
rect 289 -266 290 -265
rect 296 -266 297 -265
rect 303 -266 304 -265
rect 345 -266 346 -265
rect 380 -266 381 -265
rect 439 -266 440 -265
rect 443 -266 444 -265
rect 520 -266 521 -265
rect 114 -268 115 -267
rect 289 -268 290 -267
rect 310 -268 311 -267
rect 401 -268 402 -267
rect 415 -268 416 -267
rect 429 -268 430 -267
rect 457 -268 458 -267
rect 611 -268 612 -267
rect 114 -270 115 -269
rect 261 -270 262 -269
rect 282 -270 283 -269
rect 443 -270 444 -269
rect 457 -270 458 -269
rect 464 -270 465 -269
rect 471 -270 472 -269
rect 569 -270 570 -269
rect 128 -272 129 -271
rect 380 -272 381 -271
rect 387 -272 388 -271
rect 555 -272 556 -271
rect 107 -274 108 -273
rect 128 -274 129 -273
rect 152 -274 153 -273
rect 261 -274 262 -273
rect 299 -274 300 -273
rect 415 -274 416 -273
rect 107 -276 108 -275
rect 191 -276 192 -275
rect 222 -276 223 -275
rect 464 -276 465 -275
rect 152 -278 153 -277
rect 163 -278 164 -277
rect 170 -278 171 -277
rect 303 -278 304 -277
rect 313 -278 314 -277
rect 541 -278 542 -277
rect 40 -280 41 -279
rect 170 -280 171 -279
rect 317 -280 318 -279
rect 324 -280 325 -279
rect 366 -280 367 -279
rect 387 -280 388 -279
rect 394 -280 395 -279
rect 548 -280 549 -279
rect 215 -282 216 -281
rect 394 -282 395 -281
rect 450 -282 451 -281
rect 541 -282 542 -281
rect 215 -284 216 -283
rect 233 -284 234 -283
rect 373 -284 374 -283
rect 471 -284 472 -283
rect 163 -286 164 -285
rect 373 -286 374 -285
rect 436 -286 437 -285
rect 450 -286 451 -285
rect 9 -297 10 -296
rect 317 -297 318 -296
rect 320 -297 321 -296
rect 534 -297 535 -296
rect 653 -297 654 -296
rect 656 -297 657 -296
rect 660 -297 661 -296
rect 674 -297 675 -296
rect 30 -299 31 -298
rect 163 -299 164 -298
rect 191 -299 192 -298
rect 380 -299 381 -298
rect 387 -299 388 -298
rect 569 -299 570 -298
rect 653 -299 654 -298
rect 660 -299 661 -298
rect 30 -301 31 -300
rect 219 -301 220 -300
rect 247 -301 248 -300
rect 352 -301 353 -300
rect 359 -301 360 -300
rect 611 -301 612 -300
rect 44 -303 45 -302
rect 219 -303 220 -302
rect 247 -303 248 -302
rect 296 -303 297 -302
rect 310 -303 311 -302
rect 506 -303 507 -302
rect 534 -303 535 -302
rect 562 -303 563 -302
rect 569 -303 570 -302
rect 604 -303 605 -302
rect 611 -303 612 -302
rect 632 -303 633 -302
rect 51 -305 52 -304
rect 212 -305 213 -304
rect 215 -305 216 -304
rect 485 -305 486 -304
rect 506 -305 507 -304
rect 513 -305 514 -304
rect 562 -305 563 -304
rect 597 -305 598 -304
rect 604 -305 605 -304
rect 618 -305 619 -304
rect 58 -307 59 -306
rect 152 -307 153 -306
rect 156 -307 157 -306
rect 187 -307 188 -306
rect 191 -307 192 -306
rect 226 -307 227 -306
rect 254 -307 255 -306
rect 499 -307 500 -306
rect 597 -307 598 -306
rect 625 -307 626 -306
rect 65 -309 66 -308
rect 268 -309 269 -308
rect 289 -309 290 -308
rect 513 -309 514 -308
rect 79 -311 80 -310
rect 394 -311 395 -310
rect 401 -311 402 -310
rect 404 -311 405 -310
rect 429 -311 430 -310
rect 485 -311 486 -310
rect 79 -313 80 -312
rect 135 -313 136 -312
rect 170 -313 171 -312
rect 268 -313 269 -312
rect 289 -313 290 -312
rect 390 -313 391 -312
rect 401 -313 402 -312
rect 422 -313 423 -312
rect 432 -313 433 -312
rect 576 -313 577 -312
rect 23 -315 24 -314
rect 170 -315 171 -314
rect 205 -315 206 -314
rect 233 -315 234 -314
rect 240 -315 241 -314
rect 254 -315 255 -314
rect 257 -315 258 -314
rect 303 -315 304 -314
rect 310 -315 311 -314
rect 366 -315 367 -314
rect 373 -315 374 -314
rect 383 -315 384 -314
rect 408 -315 409 -314
rect 576 -315 577 -314
rect 86 -317 87 -316
rect 149 -317 150 -316
rect 313 -317 314 -316
rect 527 -317 528 -316
rect 86 -319 87 -318
rect 275 -319 276 -318
rect 317 -319 318 -318
rect 345 -319 346 -318
rect 352 -319 353 -318
rect 555 -319 556 -318
rect 26 -321 27 -320
rect 345 -321 346 -320
rect 373 -321 374 -320
rect 471 -321 472 -320
rect 478 -321 479 -320
rect 492 -321 493 -320
rect 527 -321 528 -320
rect 590 -321 591 -320
rect 93 -323 94 -322
rect 233 -323 234 -322
rect 331 -323 332 -322
rect 555 -323 556 -322
rect 93 -325 94 -324
rect 142 -325 143 -324
rect 261 -325 262 -324
rect 331 -325 332 -324
rect 338 -325 339 -324
rect 548 -325 549 -324
rect 100 -327 101 -326
rect 250 -327 251 -326
rect 324 -327 325 -326
rect 338 -327 339 -326
rect 341 -327 342 -326
rect 394 -327 395 -326
rect 408 -327 409 -326
rect 541 -327 542 -326
rect 548 -327 549 -326
rect 621 -327 622 -326
rect 100 -329 101 -328
rect 226 -329 227 -328
rect 415 -329 416 -328
rect 422 -329 423 -328
rect 436 -329 437 -328
rect 590 -329 591 -328
rect 110 -331 111 -330
rect 177 -331 178 -330
rect 222 -331 223 -330
rect 261 -331 262 -330
rect 404 -331 405 -330
rect 415 -331 416 -330
rect 457 -331 458 -330
rect 471 -331 472 -330
rect 492 -331 493 -330
rect 520 -331 521 -330
rect 541 -331 542 -330
rect 583 -331 584 -330
rect 72 -333 73 -332
rect 177 -333 178 -332
rect 222 -333 223 -332
rect 362 -333 363 -332
rect 450 -333 451 -332
rect 520 -333 521 -332
rect 72 -335 73 -334
rect 198 -335 199 -334
rect 362 -335 363 -334
rect 429 -335 430 -334
rect 457 -335 458 -334
rect 464 -335 465 -334
rect 107 -337 108 -336
rect 198 -337 199 -336
rect 299 -337 300 -336
rect 464 -337 465 -336
rect 107 -339 108 -338
rect 436 -339 437 -338
rect 114 -341 115 -340
rect 282 -341 283 -340
rect 299 -341 300 -340
rect 443 -341 444 -340
rect 114 -343 115 -342
rect 303 -343 304 -342
rect 443 -343 444 -342
rect 453 -343 454 -342
rect 121 -345 122 -344
rect 163 -345 164 -344
rect 166 -345 167 -344
rect 583 -345 584 -344
rect 128 -347 129 -346
rect 240 -347 241 -346
rect 135 -349 136 -348
rect 278 -349 279 -348
rect 58 -351 59 -350
rect 278 -351 279 -350
rect 142 -353 143 -352
rect 184 -353 185 -352
rect 128 -355 129 -354
rect 184 -355 185 -354
rect 9 -366 10 -365
rect 117 -366 118 -365
rect 128 -366 129 -365
rect 285 -366 286 -365
rect 324 -366 325 -365
rect 639 -366 640 -365
rect 653 -366 654 -365
rect 670 -366 671 -365
rect 674 -366 675 -365
rect 681 -366 682 -365
rect 16 -368 17 -367
rect 142 -368 143 -367
rect 170 -368 171 -367
rect 436 -368 437 -367
rect 453 -368 454 -367
rect 569 -368 570 -367
rect 583 -368 584 -367
rect 653 -368 654 -367
rect 660 -368 661 -367
rect 674 -368 675 -367
rect 23 -370 24 -369
rect 121 -370 122 -369
rect 128 -370 129 -369
rect 208 -370 209 -369
rect 219 -370 220 -369
rect 499 -370 500 -369
rect 520 -370 521 -369
rect 667 -370 668 -369
rect 30 -372 31 -371
rect 324 -372 325 -371
rect 341 -372 342 -371
rect 401 -372 402 -371
rect 408 -372 409 -371
rect 569 -372 570 -371
rect 583 -372 584 -371
rect 611 -372 612 -371
rect 44 -374 45 -373
rect 194 -374 195 -373
rect 212 -374 213 -373
rect 408 -374 409 -373
rect 429 -374 430 -373
rect 618 -374 619 -373
rect 51 -376 52 -375
rect 180 -376 181 -375
rect 229 -376 230 -375
rect 632 -376 633 -375
rect 58 -378 59 -377
rect 296 -378 297 -377
rect 359 -378 360 -377
rect 492 -378 493 -377
rect 506 -378 507 -377
rect 520 -378 521 -377
rect 548 -378 549 -377
rect 611 -378 612 -377
rect 33 -380 34 -379
rect 548 -380 549 -379
rect 555 -380 556 -379
rect 646 -380 647 -379
rect 72 -382 73 -381
rect 152 -382 153 -381
rect 177 -382 178 -381
rect 250 -382 251 -381
rect 254 -382 255 -381
rect 296 -382 297 -381
rect 366 -382 367 -381
rect 457 -382 458 -381
rect 464 -382 465 -381
rect 492 -382 493 -381
rect 562 -382 563 -381
rect 625 -382 626 -381
rect 72 -384 73 -383
rect 86 -384 87 -383
rect 100 -384 101 -383
rect 163 -384 164 -383
rect 275 -384 276 -383
rect 373 -384 374 -383
rect 383 -384 384 -383
rect 576 -384 577 -383
rect 604 -384 605 -383
rect 660 -384 661 -383
rect 65 -386 66 -385
rect 163 -386 164 -385
rect 275 -386 276 -385
rect 303 -386 304 -385
rect 345 -386 346 -385
rect 464 -386 465 -385
rect 471 -386 472 -385
rect 576 -386 577 -385
rect 79 -388 80 -387
rect 222 -388 223 -387
rect 240 -388 241 -387
rect 303 -388 304 -387
rect 338 -388 339 -387
rect 345 -388 346 -387
rect 352 -388 353 -387
rect 457 -388 458 -387
rect 478 -388 479 -387
rect 506 -388 507 -387
rect 527 -388 528 -387
rect 604 -388 605 -387
rect 86 -390 87 -389
rect 264 -390 265 -389
rect 282 -390 283 -389
rect 366 -390 367 -389
rect 383 -390 384 -389
rect 527 -390 528 -389
rect 93 -392 94 -391
rect 222 -392 223 -391
rect 261 -392 262 -391
rect 282 -392 283 -391
rect 289 -392 290 -391
rect 373 -392 374 -391
rect 387 -392 388 -391
rect 450 -392 451 -391
rect 481 -392 482 -391
rect 590 -392 591 -391
rect 93 -394 94 -393
rect 159 -394 160 -393
rect 198 -394 199 -393
rect 240 -394 241 -393
rect 331 -394 332 -393
rect 352 -394 353 -393
rect 355 -394 356 -393
rect 590 -394 591 -393
rect 107 -396 108 -395
rect 166 -396 167 -395
rect 233 -396 234 -395
rect 289 -396 290 -395
rect 310 -396 311 -395
rect 331 -396 332 -395
rect 362 -396 363 -395
rect 562 -396 563 -395
rect 107 -398 108 -397
rect 261 -398 262 -397
rect 317 -398 318 -397
rect 362 -398 363 -397
rect 390 -398 391 -397
rect 597 -398 598 -397
rect 114 -400 115 -399
rect 555 -400 556 -399
rect 121 -402 122 -401
rect 327 -402 328 -401
rect 401 -402 402 -401
rect 415 -402 416 -401
rect 422 -402 423 -401
rect 429 -402 430 -401
rect 436 -402 437 -401
rect 443 -402 444 -401
rect 534 -402 535 -401
rect 597 -402 598 -401
rect 135 -404 136 -403
rect 177 -404 178 -403
rect 268 -404 269 -403
rect 422 -404 423 -403
rect 135 -406 136 -405
rect 156 -406 157 -405
rect 170 -406 171 -405
rect 233 -406 234 -405
rect 317 -406 318 -405
rect 513 -406 514 -405
rect 138 -408 139 -407
rect 254 -408 255 -407
rect 387 -408 388 -407
rect 534 -408 535 -407
rect 142 -410 143 -409
rect 215 -410 216 -409
rect 226 -410 227 -409
rect 268 -410 269 -409
rect 394 -410 395 -409
rect 415 -410 416 -409
rect 485 -410 486 -409
rect 513 -410 514 -409
rect 117 -412 118 -411
rect 485 -412 486 -411
rect 149 -414 150 -413
rect 198 -414 199 -413
rect 247 -414 248 -413
rect 394 -414 395 -413
rect 149 -416 150 -415
rect 191 -416 192 -415
rect 247 -416 248 -415
rect 443 -416 444 -415
rect 184 -418 185 -417
rect 226 -418 227 -417
rect 191 -420 192 -419
rect 541 -420 542 -419
rect 474 -422 475 -421
rect 541 -422 542 -421
rect 16 -433 17 -432
rect 243 -433 244 -432
rect 257 -433 258 -432
rect 366 -433 367 -432
rect 380 -433 381 -432
rect 513 -433 514 -432
rect 541 -433 542 -432
rect 544 -433 545 -432
rect 583 -433 584 -432
rect 702 -433 703 -432
rect 33 -435 34 -434
rect 142 -435 143 -434
rect 149 -435 150 -434
rect 166 -435 167 -434
rect 201 -435 202 -434
rect 562 -435 563 -434
rect 646 -435 647 -434
rect 674 -435 675 -434
rect 40 -437 41 -436
rect 212 -437 213 -436
rect 219 -437 220 -436
rect 548 -437 549 -436
rect 653 -437 654 -436
rect 688 -437 689 -436
rect 44 -439 45 -438
rect 513 -439 514 -438
rect 527 -439 528 -438
rect 583 -439 584 -438
rect 639 -439 640 -438
rect 653 -439 654 -438
rect 44 -441 45 -440
rect 156 -441 157 -440
rect 205 -441 206 -440
rect 464 -441 465 -440
rect 471 -441 472 -440
rect 625 -441 626 -440
rect 632 -441 633 -440
rect 639 -441 640 -440
rect 51 -443 52 -442
rect 383 -443 384 -442
rect 390 -443 391 -442
rect 576 -443 577 -442
rect 611 -443 612 -442
rect 625 -443 626 -442
rect 58 -445 59 -444
rect 296 -445 297 -444
rect 320 -445 321 -444
rect 429 -445 430 -444
rect 450 -445 451 -444
rect 611 -445 612 -444
rect 618 -445 619 -444
rect 632 -445 633 -444
rect 65 -447 66 -446
rect 205 -447 206 -446
rect 222 -447 223 -446
rect 562 -447 563 -446
rect 65 -449 66 -448
rect 348 -449 349 -448
rect 352 -449 353 -448
rect 366 -449 367 -448
rect 390 -449 391 -448
rect 667 -449 668 -448
rect 72 -451 73 -450
rect 173 -451 174 -450
rect 177 -451 178 -450
rect 667 -451 668 -450
rect 72 -453 73 -452
rect 198 -453 199 -452
rect 229 -453 230 -452
rect 240 -453 241 -452
rect 257 -453 258 -452
rect 464 -453 465 -452
rect 478 -453 479 -452
rect 646 -453 647 -452
rect 79 -455 80 -454
rect 121 -455 122 -454
rect 128 -455 129 -454
rect 131 -455 132 -454
rect 135 -455 136 -454
rect 254 -455 255 -454
rect 264 -455 265 -454
rect 415 -455 416 -454
rect 425 -455 426 -454
rect 590 -455 591 -454
rect 82 -457 83 -456
rect 149 -457 150 -456
rect 156 -457 157 -456
rect 303 -457 304 -456
rect 331 -457 332 -456
rect 429 -457 430 -456
rect 439 -457 440 -456
rect 478 -457 479 -456
rect 485 -457 486 -456
rect 527 -457 528 -456
rect 534 -457 535 -456
rect 590 -457 591 -456
rect 93 -459 94 -458
rect 163 -459 164 -458
rect 177 -459 178 -458
rect 338 -459 339 -458
rect 345 -459 346 -458
rect 380 -459 381 -458
rect 401 -459 402 -458
rect 471 -459 472 -458
rect 492 -459 493 -458
rect 534 -459 535 -458
rect 541 -459 542 -458
rect 597 -459 598 -458
rect 100 -461 101 -460
rect 331 -461 332 -460
rect 338 -461 339 -460
rect 408 -461 409 -460
rect 443 -461 444 -460
rect 485 -461 486 -460
rect 499 -461 500 -460
rect 618 -461 619 -460
rect 100 -463 101 -462
rect 198 -463 199 -462
rect 215 -463 216 -462
rect 415 -463 416 -462
rect 436 -463 437 -462
rect 499 -463 500 -462
rect 520 -463 521 -462
rect 576 -463 577 -462
rect 107 -465 108 -464
rect 247 -465 248 -464
rect 275 -465 276 -464
rect 520 -465 521 -464
rect 61 -467 62 -466
rect 275 -467 276 -466
rect 310 -467 311 -466
rect 408 -467 409 -466
rect 450 -467 451 -466
rect 709 -467 710 -466
rect 110 -469 111 -468
rect 443 -469 444 -468
rect 457 -469 458 -468
rect 492 -469 493 -468
rect 114 -471 115 -470
rect 569 -471 570 -470
rect 114 -473 115 -472
rect 362 -473 363 -472
rect 117 -475 118 -474
rect 373 -475 374 -474
rect 128 -477 129 -476
rect 289 -477 290 -476
rect 327 -477 328 -476
rect 373 -477 374 -476
rect 184 -479 185 -478
rect 310 -479 311 -478
rect 355 -479 356 -478
rect 569 -479 570 -478
rect 86 -481 87 -480
rect 184 -481 185 -480
rect 191 -481 192 -480
rect 327 -481 328 -480
rect 359 -481 360 -480
rect 506 -481 507 -480
rect 544 -481 545 -480
rect 597 -481 598 -480
rect 86 -483 87 -482
rect 93 -483 94 -482
rect 194 -483 195 -482
rect 506 -483 507 -482
rect 215 -485 216 -484
rect 422 -485 423 -484
rect 226 -487 227 -486
rect 457 -487 458 -486
rect 226 -489 227 -488
rect 268 -489 269 -488
rect 359 -489 360 -488
rect 604 -489 605 -488
rect 229 -491 230 -490
rect 261 -491 262 -490
rect 268 -491 269 -490
rect 303 -491 304 -490
rect 422 -491 423 -490
rect 548 -491 549 -490
rect 555 -491 556 -490
rect 604 -491 605 -490
rect 37 -493 38 -492
rect 555 -493 556 -492
rect 233 -495 234 -494
rect 352 -495 353 -494
rect 233 -497 234 -496
rect 271 -497 272 -496
rect 240 -499 241 -498
rect 394 -499 395 -498
rect 247 -501 248 -500
rect 320 -501 321 -500
rect 387 -501 388 -500
rect 394 -501 395 -500
rect 261 -503 262 -502
rect 317 -503 318 -502
rect 317 -505 318 -504
rect 660 -505 661 -504
rect 282 -507 283 -506
rect 660 -507 661 -506
rect 282 -509 283 -508
rect 695 -509 696 -508
rect 16 -520 17 -519
rect 345 -520 346 -519
rect 348 -520 349 -519
rect 611 -520 612 -519
rect 23 -522 24 -521
rect 499 -522 500 -521
rect 558 -522 559 -521
rect 674 -522 675 -521
rect 26 -524 27 -523
rect 310 -524 311 -523
rect 324 -524 325 -523
rect 471 -524 472 -523
rect 502 -524 503 -523
rect 674 -524 675 -523
rect 30 -526 31 -525
rect 436 -526 437 -525
rect 460 -526 461 -525
rect 618 -526 619 -525
rect 30 -528 31 -527
rect 464 -528 465 -527
rect 611 -528 612 -527
rect 695 -528 696 -527
rect 37 -530 38 -529
rect 299 -530 300 -529
rect 310 -530 311 -529
rect 418 -530 419 -529
rect 464 -530 465 -529
rect 513 -530 514 -529
rect 618 -530 619 -529
rect 639 -530 640 -529
rect 44 -532 45 -531
rect 285 -532 286 -531
rect 296 -532 297 -531
rect 429 -532 430 -531
rect 513 -532 514 -531
rect 667 -532 668 -531
rect 44 -534 45 -533
rect 100 -534 101 -533
rect 107 -534 108 -533
rect 562 -534 563 -533
rect 576 -534 577 -533
rect 667 -534 668 -533
rect 58 -536 59 -535
rect 257 -536 258 -535
rect 282 -536 283 -535
rect 289 -536 290 -535
rect 327 -536 328 -535
rect 485 -536 486 -535
rect 562 -536 563 -535
rect 583 -536 584 -535
rect 639 -536 640 -535
rect 660 -536 661 -535
rect 51 -538 52 -537
rect 660 -538 661 -537
rect 58 -540 59 -539
rect 373 -540 374 -539
rect 387 -540 388 -539
rect 495 -540 496 -539
rect 65 -542 66 -541
rect 324 -542 325 -541
rect 352 -542 353 -541
rect 390 -542 391 -541
rect 401 -542 402 -541
rect 520 -542 521 -541
rect 65 -544 66 -543
rect 296 -544 297 -543
rect 306 -544 307 -543
rect 583 -544 584 -543
rect 68 -546 69 -545
rect 576 -546 577 -545
rect 72 -548 73 -547
rect 124 -548 125 -547
rect 128 -548 129 -547
rect 320 -548 321 -547
rect 355 -548 356 -547
rect 653 -548 654 -547
rect 54 -550 55 -549
rect 72 -550 73 -549
rect 79 -550 80 -549
rect 219 -550 220 -549
rect 240 -550 241 -549
rect 250 -550 251 -549
rect 254 -550 255 -549
rect 415 -550 416 -549
rect 425 -550 426 -549
rect 429 -550 430 -549
rect 520 -550 521 -549
rect 590 -550 591 -549
rect 79 -552 80 -551
rect 117 -552 118 -551
rect 131 -552 132 -551
rect 401 -552 402 -551
rect 404 -552 405 -551
rect 688 -552 689 -551
rect 86 -554 87 -553
rect 184 -554 185 -553
rect 194 -554 195 -553
rect 555 -554 556 -553
rect 114 -556 115 -555
rect 226 -556 227 -555
rect 233 -556 234 -555
rect 254 -556 255 -555
rect 285 -556 286 -555
rect 527 -556 528 -555
rect 541 -556 542 -555
rect 590 -556 591 -555
rect 107 -558 108 -557
rect 527 -558 528 -557
rect 541 -558 542 -557
rect 597 -558 598 -557
rect 114 -560 115 -559
rect 569 -560 570 -559
rect 135 -562 136 -561
rect 359 -562 360 -561
rect 387 -562 388 -561
rect 450 -562 451 -561
rect 478 -562 479 -561
rect 597 -562 598 -561
rect 135 -564 136 -563
rect 492 -564 493 -563
rect 569 -564 570 -563
rect 625 -564 626 -563
rect 145 -566 146 -565
rect 534 -566 535 -565
rect 625 -566 626 -565
rect 646 -566 647 -565
rect 170 -568 171 -567
rect 198 -568 199 -567
rect 201 -568 202 -567
rect 338 -568 339 -567
rect 408 -568 409 -567
rect 439 -568 440 -567
rect 478 -568 479 -567
rect 506 -568 507 -567
rect 534 -568 535 -567
rect 632 -568 633 -567
rect 177 -570 178 -569
rect 201 -570 202 -569
rect 205 -570 206 -569
rect 268 -570 269 -569
rect 289 -570 290 -569
rect 317 -570 318 -569
rect 320 -570 321 -569
rect 450 -570 451 -569
rect 506 -570 507 -569
rect 604 -570 605 -569
rect 163 -572 164 -571
rect 177 -572 178 -571
rect 184 -572 185 -571
rect 362 -572 363 -571
rect 394 -572 395 -571
rect 408 -572 409 -571
rect 411 -572 412 -571
rect 653 -572 654 -571
rect 159 -574 160 -573
rect 163 -574 164 -573
rect 205 -574 206 -573
rect 212 -574 213 -573
rect 215 -574 216 -573
rect 632 -574 633 -573
rect 215 -576 216 -575
rect 457 -576 458 -575
rect 492 -576 493 -575
rect 604 -576 605 -575
rect 219 -578 220 -577
rect 331 -578 332 -577
rect 422 -578 423 -577
rect 439 -578 440 -577
rect 457 -578 458 -577
rect 709 -578 710 -577
rect 233 -580 234 -579
rect 338 -580 339 -579
rect 548 -580 549 -579
rect 646 -580 647 -579
rect 681 -580 682 -579
rect 709 -580 710 -579
rect 121 -582 122 -581
rect 548 -582 549 -581
rect 121 -584 122 -583
rect 142 -584 143 -583
rect 173 -584 174 -583
rect 681 -584 682 -583
rect 142 -586 143 -585
rect 156 -586 157 -585
rect 240 -586 241 -585
rect 261 -586 262 -585
rect 275 -586 276 -585
rect 331 -586 332 -585
rect 243 -588 244 -587
rect 485 -588 486 -587
rect 247 -590 248 -589
rect 394 -590 395 -589
rect 149 -592 150 -591
rect 247 -592 248 -591
rect 250 -592 251 -591
rect 261 -592 262 -591
rect 275 -592 276 -591
rect 443 -592 444 -591
rect 149 -594 150 -593
rect 191 -594 192 -593
rect 317 -594 318 -593
rect 380 -594 381 -593
rect 443 -594 444 -593
rect 702 -594 703 -593
rect 303 -596 304 -595
rect 380 -596 381 -595
rect 23 -607 24 -606
rect 376 -607 377 -606
rect 411 -607 412 -606
rect 583 -607 584 -606
rect 611 -607 612 -606
rect 737 -607 738 -606
rect 30 -609 31 -608
rect 702 -609 703 -608
rect 709 -609 710 -608
rect 765 -609 766 -608
rect 37 -611 38 -610
rect 72 -611 73 -610
rect 93 -611 94 -610
rect 103 -611 104 -610
rect 107 -611 108 -610
rect 562 -611 563 -610
rect 632 -611 633 -610
rect 772 -611 773 -610
rect 37 -613 38 -612
rect 184 -613 185 -612
rect 187 -613 188 -612
rect 201 -613 202 -612
rect 219 -613 220 -612
rect 660 -613 661 -612
rect 674 -613 675 -612
rect 751 -613 752 -612
rect 44 -615 45 -614
rect 65 -615 66 -614
rect 93 -615 94 -614
rect 380 -615 381 -614
rect 415 -615 416 -614
rect 527 -615 528 -614
rect 541 -615 542 -614
rect 688 -615 689 -614
rect 44 -617 45 -616
rect 215 -617 216 -616
rect 222 -617 223 -616
rect 723 -617 724 -616
rect 51 -619 52 -618
rect 352 -619 353 -618
rect 355 -619 356 -618
rect 744 -619 745 -618
rect 58 -621 59 -620
rect 65 -621 66 -620
rect 100 -621 101 -620
rect 198 -621 199 -620
rect 212 -621 213 -620
rect 222 -621 223 -620
rect 233 -621 234 -620
rect 338 -621 339 -620
rect 348 -621 349 -620
rect 562 -621 563 -620
rect 569 -621 570 -620
rect 660 -621 661 -620
rect 681 -621 682 -620
rect 758 -621 759 -620
rect 23 -623 24 -622
rect 58 -623 59 -622
rect 75 -623 76 -622
rect 233 -623 234 -622
rect 275 -623 276 -622
rect 387 -623 388 -622
rect 418 -623 419 -622
rect 506 -623 507 -622
rect 513 -623 514 -622
rect 716 -623 717 -622
rect 79 -625 80 -624
rect 100 -625 101 -624
rect 107 -625 108 -624
rect 142 -625 143 -624
rect 170 -625 171 -624
rect 191 -625 192 -624
rect 282 -625 283 -624
rect 527 -625 528 -624
rect 555 -625 556 -624
rect 695 -625 696 -624
rect 79 -627 80 -626
rect 205 -627 206 -626
rect 303 -627 304 -626
rect 331 -627 332 -626
rect 380 -627 381 -626
rect 401 -627 402 -626
rect 422 -627 423 -626
rect 443 -627 444 -626
rect 450 -627 451 -626
rect 569 -627 570 -626
rect 583 -627 584 -626
rect 632 -627 633 -626
rect 639 -627 640 -626
rect 709 -627 710 -626
rect 114 -629 115 -628
rect 261 -629 262 -628
rect 296 -629 297 -628
rect 331 -629 332 -628
rect 425 -629 426 -628
rect 653 -629 654 -628
rect 117 -631 118 -630
rect 247 -631 248 -630
rect 261 -631 262 -630
rect 408 -631 409 -630
rect 439 -631 440 -630
rect 534 -631 535 -630
rect 590 -631 591 -630
rect 653 -631 654 -630
rect 54 -633 55 -632
rect 439 -633 440 -632
rect 453 -633 454 -632
rect 639 -633 640 -632
rect 121 -635 122 -634
rect 387 -635 388 -634
rect 457 -635 458 -634
rect 611 -635 612 -634
rect 618 -635 619 -634
rect 681 -635 682 -634
rect 124 -637 125 -636
rect 674 -637 675 -636
rect 128 -639 129 -638
rect 359 -639 360 -638
rect 457 -639 458 -638
rect 520 -639 521 -638
rect 135 -641 136 -640
rect 513 -641 514 -640
rect 142 -643 143 -642
rect 401 -643 402 -642
rect 464 -643 465 -642
rect 555 -643 556 -642
rect 163 -645 164 -644
rect 170 -645 171 -644
rect 198 -645 199 -644
rect 590 -645 591 -644
rect 149 -647 150 -646
rect 163 -647 164 -646
rect 247 -647 248 -646
rect 268 -647 269 -646
rect 296 -647 297 -646
rect 422 -647 423 -646
rect 429 -647 430 -646
rect 464 -647 465 -646
rect 471 -647 472 -646
rect 534 -647 535 -646
rect 19 -649 20 -648
rect 149 -649 150 -648
rect 303 -649 304 -648
rect 404 -649 405 -648
rect 478 -649 479 -648
rect 520 -649 521 -648
rect 86 -651 87 -650
rect 268 -651 269 -650
rect 310 -651 311 -650
rect 408 -651 409 -650
rect 478 -651 479 -650
rect 667 -651 668 -650
rect 86 -653 87 -652
rect 285 -653 286 -652
rect 317 -653 318 -652
rect 730 -653 731 -652
rect 177 -655 178 -654
rect 310 -655 311 -654
rect 320 -655 321 -654
rect 576 -655 577 -654
rect 604 -655 605 -654
rect 667 -655 668 -654
rect 177 -657 178 -656
rect 240 -657 241 -656
rect 359 -657 360 -656
rect 446 -657 447 -656
rect 485 -657 486 -656
rect 541 -657 542 -656
rect 548 -657 549 -656
rect 604 -657 605 -656
rect 159 -659 160 -658
rect 240 -659 241 -658
rect 373 -659 374 -658
rect 576 -659 577 -658
rect 194 -661 195 -660
rect 285 -661 286 -660
rect 324 -661 325 -660
rect 373 -661 374 -660
rect 394 -661 395 -660
rect 429 -661 430 -660
rect 467 -661 468 -660
rect 485 -661 486 -660
rect 492 -661 493 -660
rect 646 -661 647 -660
rect 201 -663 202 -662
rect 548 -663 549 -662
rect 205 -665 206 -664
rect 394 -665 395 -664
rect 460 -665 461 -664
rect 646 -665 647 -664
rect 324 -667 325 -666
rect 618 -667 619 -666
rect 499 -669 500 -668
rect 597 -669 598 -668
rect 135 -671 136 -670
rect 597 -671 598 -670
rect 289 -673 290 -672
rect 499 -673 500 -672
rect 289 -675 290 -674
rect 317 -675 318 -674
rect 30 -686 31 -685
rect 457 -686 458 -685
rect 467 -686 468 -685
rect 758 -686 759 -685
rect 765 -686 766 -685
rect 793 -686 794 -685
rect 37 -688 38 -687
rect 324 -688 325 -687
rect 345 -688 346 -687
rect 639 -688 640 -687
rect 730 -688 731 -687
rect 779 -688 780 -687
rect 37 -690 38 -689
rect 107 -690 108 -689
rect 114 -690 115 -689
rect 422 -690 423 -689
rect 443 -690 444 -689
rect 471 -690 472 -689
rect 485 -690 486 -689
rect 492 -690 493 -689
rect 506 -690 507 -689
rect 765 -690 766 -689
rect 772 -690 773 -689
rect 849 -690 850 -689
rect 44 -692 45 -691
rect 355 -692 356 -691
rect 362 -692 363 -691
rect 366 -692 367 -691
rect 380 -692 381 -691
rect 457 -692 458 -691
rect 495 -692 496 -691
rect 772 -692 773 -691
rect 44 -694 45 -693
rect 93 -694 94 -693
rect 107 -694 108 -693
rect 303 -694 304 -693
rect 320 -694 321 -693
rect 555 -694 556 -693
rect 586 -694 587 -693
rect 751 -694 752 -693
rect 51 -696 52 -695
rect 436 -696 437 -695
rect 450 -696 451 -695
rect 590 -696 591 -695
rect 604 -696 605 -695
rect 639 -696 640 -695
rect 744 -696 745 -695
rect 786 -696 787 -695
rect 54 -698 55 -697
rect 352 -698 353 -697
rect 359 -698 360 -697
rect 366 -698 367 -697
rect 383 -698 384 -697
rect 702 -698 703 -697
rect 58 -700 59 -699
rect 61 -700 62 -699
rect 65 -700 66 -699
rect 327 -700 328 -699
rect 345 -700 346 -699
rect 355 -700 356 -699
rect 397 -700 398 -699
rect 681 -700 682 -699
rect 65 -702 66 -701
rect 499 -702 500 -701
rect 506 -702 507 -701
rect 513 -702 514 -701
rect 555 -702 556 -701
rect 562 -702 563 -701
rect 597 -702 598 -701
rect 604 -702 605 -701
rect 632 -702 633 -701
rect 758 -702 759 -701
rect 72 -704 73 -703
rect 744 -704 745 -703
rect 72 -706 73 -705
rect 93 -706 94 -705
rect 124 -706 125 -705
rect 289 -706 290 -705
rect 296 -706 297 -705
rect 464 -706 465 -705
rect 478 -706 479 -705
rect 632 -706 633 -705
rect 646 -706 647 -705
rect 681 -706 682 -705
rect 86 -708 87 -707
rect 187 -708 188 -707
rect 222 -708 223 -707
rect 310 -708 311 -707
rect 320 -708 321 -707
rect 733 -708 734 -707
rect 89 -710 90 -709
rect 404 -710 405 -709
rect 415 -710 416 -709
rect 590 -710 591 -709
rect 625 -710 626 -709
rect 646 -710 647 -709
rect 653 -710 654 -709
rect 702 -710 703 -709
rect 128 -712 129 -711
rect 261 -712 262 -711
rect 268 -712 269 -711
rect 282 -712 283 -711
rect 289 -712 290 -711
rect 509 -712 510 -711
rect 562 -712 563 -711
rect 569 -712 570 -711
rect 611 -712 612 -711
rect 653 -712 654 -711
rect 79 -714 80 -713
rect 268 -714 269 -713
rect 282 -714 283 -713
rect 751 -714 752 -713
rect 79 -716 80 -715
rect 723 -716 724 -715
rect 131 -718 132 -717
rect 387 -718 388 -717
rect 397 -718 398 -717
rect 688 -718 689 -717
rect 695 -718 696 -717
rect 723 -718 724 -717
rect 16 -720 17 -719
rect 688 -720 689 -719
rect 135 -722 136 -721
rect 583 -722 584 -721
rect 618 -722 619 -721
rect 625 -722 626 -721
rect 135 -724 136 -723
rect 205 -724 206 -723
rect 233 -724 234 -723
rect 394 -724 395 -723
rect 401 -724 402 -723
rect 737 -724 738 -723
rect 114 -726 115 -725
rect 401 -726 402 -725
rect 408 -726 409 -725
rect 415 -726 416 -725
rect 429 -726 430 -725
rect 597 -726 598 -725
rect 621 -726 622 -725
rect 695 -726 696 -725
rect 121 -728 122 -727
rect 233 -728 234 -727
rect 247 -728 248 -727
rect 306 -728 307 -727
rect 348 -728 349 -727
rect 481 -728 482 -727
rect 499 -728 500 -727
rect 534 -728 535 -727
rect 142 -730 143 -729
rect 674 -730 675 -729
rect 124 -732 125 -731
rect 142 -732 143 -731
rect 145 -732 146 -731
rect 159 -732 160 -731
rect 163 -732 164 -731
rect 408 -732 409 -731
rect 429 -732 430 -731
rect 660 -732 661 -731
rect 86 -734 87 -733
rect 660 -734 661 -733
rect 156 -736 157 -735
rect 716 -736 717 -735
rect 156 -738 157 -737
rect 222 -738 223 -737
rect 247 -738 248 -737
rect 303 -738 304 -737
rect 348 -738 349 -737
rect 716 -738 717 -737
rect 163 -740 164 -739
rect 278 -740 279 -739
rect 373 -740 374 -739
rect 387 -740 388 -739
rect 394 -740 395 -739
rect 569 -740 570 -739
rect 184 -742 185 -741
rect 737 -742 738 -741
rect 170 -744 171 -743
rect 184 -744 185 -743
rect 191 -744 192 -743
rect 205 -744 206 -743
rect 254 -744 255 -743
rect 275 -744 276 -743
rect 373 -744 374 -743
rect 488 -744 489 -743
rect 149 -746 150 -745
rect 275 -746 276 -745
rect 436 -746 437 -745
rect 674 -746 675 -745
rect 149 -748 150 -747
rect 709 -748 710 -747
rect 170 -750 171 -749
rect 226 -750 227 -749
rect 254 -750 255 -749
rect 313 -750 314 -749
rect 453 -750 454 -749
rect 513 -750 514 -749
rect 576 -750 577 -749
rect 709 -750 710 -749
rect 177 -752 178 -751
rect 191 -752 192 -751
rect 201 -752 202 -751
rect 611 -752 612 -751
rect 96 -754 97 -753
rect 177 -754 178 -753
rect 201 -754 202 -753
rect 296 -754 297 -753
rect 446 -754 447 -753
rect 576 -754 577 -753
rect 226 -756 227 -755
rect 240 -756 241 -755
rect 261 -756 262 -755
rect 331 -756 332 -755
rect 481 -756 482 -755
rect 667 -756 668 -755
rect 100 -758 101 -757
rect 331 -758 332 -757
rect 439 -758 440 -757
rect 667 -758 668 -757
rect 30 -760 31 -759
rect 100 -760 101 -759
rect 240 -760 241 -759
rect 292 -760 293 -759
rect 439 -760 440 -759
rect 534 -760 535 -759
rect 19 -771 20 -770
rect 23 -771 24 -770
rect 30 -771 31 -770
rect 394 -771 395 -770
rect 408 -771 409 -770
rect 485 -771 486 -770
rect 488 -771 489 -770
rect 835 -771 836 -770
rect 849 -771 850 -770
rect 940 -771 941 -770
rect 23 -773 24 -772
rect 149 -773 150 -772
rect 159 -773 160 -772
rect 275 -773 276 -772
rect 289 -773 290 -772
rect 296 -773 297 -772
rect 310 -773 311 -772
rect 513 -773 514 -772
rect 534 -773 535 -772
rect 709 -773 710 -772
rect 751 -773 752 -772
rect 814 -773 815 -772
rect 37 -775 38 -774
rect 152 -775 153 -774
rect 177 -775 178 -774
rect 180 -775 181 -774
rect 201 -775 202 -774
rect 261 -775 262 -774
rect 268 -775 269 -774
rect 282 -775 283 -774
rect 292 -775 293 -774
rect 457 -775 458 -774
rect 460 -775 461 -774
rect 562 -775 563 -774
rect 621 -775 622 -774
rect 772 -775 773 -774
rect 779 -775 780 -774
rect 849 -775 850 -774
rect 37 -777 38 -776
rect 432 -777 433 -776
rect 446 -777 447 -776
rect 702 -777 703 -776
rect 758 -777 759 -776
rect 828 -777 829 -776
rect 40 -779 41 -778
rect 275 -779 276 -778
rect 296 -779 297 -778
rect 618 -779 619 -778
rect 646 -779 647 -778
rect 779 -779 780 -778
rect 793 -779 794 -778
rect 863 -779 864 -778
rect 54 -781 55 -780
rect 65 -781 66 -780
rect 86 -781 87 -780
rect 219 -781 220 -780
rect 222 -781 223 -780
rect 660 -781 661 -780
rect 667 -781 668 -780
rect 709 -781 710 -780
rect 765 -781 766 -780
rect 842 -781 843 -780
rect 44 -783 45 -782
rect 219 -783 220 -782
rect 226 -783 227 -782
rect 282 -783 283 -782
rect 317 -783 318 -782
rect 345 -783 346 -782
rect 352 -783 353 -782
rect 765 -783 766 -782
rect 44 -785 45 -784
rect 156 -785 157 -784
rect 166 -785 167 -784
rect 646 -785 647 -784
rect 674 -785 675 -784
rect 807 -785 808 -784
rect 58 -787 59 -786
rect 96 -787 97 -786
rect 100 -787 101 -786
rect 310 -787 311 -786
rect 320 -787 321 -786
rect 597 -787 598 -786
rect 688 -787 689 -786
rect 856 -787 857 -786
rect 65 -789 66 -788
rect 464 -789 465 -788
rect 467 -789 468 -788
rect 737 -789 738 -788
rect 72 -791 73 -790
rect 667 -791 668 -790
rect 681 -791 682 -790
rect 737 -791 738 -790
rect 79 -793 80 -792
rect 597 -793 598 -792
rect 639 -793 640 -792
rect 681 -793 682 -792
rect 695 -793 696 -792
rect 751 -793 752 -792
rect 79 -795 80 -794
rect 107 -795 108 -794
rect 114 -795 115 -794
rect 135 -795 136 -794
rect 149 -795 150 -794
rect 289 -795 290 -794
rect 327 -795 328 -794
rect 397 -795 398 -794
rect 411 -795 412 -794
rect 716 -795 717 -794
rect 86 -797 87 -796
rect 730 -797 731 -796
rect 93 -799 94 -798
rect 362 -799 363 -798
rect 397 -799 398 -798
rect 786 -799 787 -798
rect 117 -801 118 -800
rect 583 -801 584 -800
rect 604 -801 605 -800
rect 639 -801 640 -800
rect 653 -801 654 -800
rect 688 -801 689 -800
rect 702 -801 703 -800
rect 723 -801 724 -800
rect 121 -803 122 -802
rect 401 -803 402 -802
rect 408 -803 409 -802
rect 604 -803 605 -802
rect 611 -803 612 -802
rect 653 -803 654 -802
rect 723 -803 724 -802
rect 744 -803 745 -802
rect 72 -805 73 -804
rect 121 -805 122 -804
rect 135 -805 136 -804
rect 191 -805 192 -804
rect 198 -805 199 -804
rect 432 -805 433 -804
rect 436 -805 437 -804
rect 786 -805 787 -804
rect 152 -807 153 -806
rect 317 -807 318 -806
rect 338 -807 339 -806
rect 443 -807 444 -806
rect 446 -807 447 -806
rect 772 -807 773 -806
rect 58 -809 59 -808
rect 338 -809 339 -808
rect 352 -809 353 -808
rect 373 -809 374 -808
rect 429 -809 430 -808
rect 660 -809 661 -808
rect 674 -809 675 -808
rect 744 -809 745 -808
rect 156 -811 157 -810
rect 191 -811 192 -810
rect 226 -811 227 -810
rect 380 -811 381 -810
rect 401 -811 402 -810
rect 429 -811 430 -810
rect 464 -811 465 -810
rect 583 -811 584 -810
rect 625 -811 626 -810
rect 695 -811 696 -810
rect 177 -813 178 -812
rect 184 -813 185 -812
rect 233 -813 234 -812
rect 373 -813 374 -812
rect 513 -813 514 -812
rect 870 -813 871 -812
rect 170 -815 171 -814
rect 233 -815 234 -814
rect 240 -815 241 -814
rect 243 -815 244 -814
rect 247 -815 248 -814
rect 250 -815 251 -814
rect 254 -815 255 -814
rect 516 -815 517 -814
rect 520 -815 521 -814
rect 534 -815 535 -814
rect 537 -815 538 -814
rect 716 -815 717 -814
rect 142 -817 143 -816
rect 170 -817 171 -816
rect 184 -817 185 -816
rect 205 -817 206 -816
rect 240 -817 241 -816
rect 387 -817 388 -816
rect 548 -817 549 -816
rect 562 -817 563 -816
rect 569 -817 570 -816
rect 758 -817 759 -816
rect 142 -819 143 -818
rect 590 -819 591 -818
rect 163 -821 164 -820
rect 254 -821 255 -820
rect 268 -821 269 -820
rect 457 -821 458 -820
rect 499 -821 500 -820
rect 548 -821 549 -820
rect 555 -821 556 -820
rect 569 -821 570 -820
rect 576 -821 577 -820
rect 625 -821 626 -820
rect 128 -823 129 -822
rect 576 -823 577 -822
rect 128 -825 129 -824
rect 422 -825 423 -824
rect 471 -825 472 -824
rect 499 -825 500 -824
rect 541 -825 542 -824
rect 555 -825 556 -824
rect 163 -827 164 -826
rect 324 -827 325 -826
rect 331 -827 332 -826
rect 520 -827 521 -826
rect 527 -827 528 -826
rect 541 -827 542 -826
rect 107 -829 108 -828
rect 324 -829 325 -828
rect 331 -829 332 -828
rect 800 -829 801 -828
rect 243 -831 244 -830
rect 387 -831 388 -830
rect 471 -831 472 -830
rect 492 -831 493 -830
rect 506 -831 507 -830
rect 527 -831 528 -830
rect 299 -833 300 -832
rect 422 -833 423 -832
rect 506 -833 507 -832
rect 821 -833 822 -832
rect 306 -835 307 -834
rect 590 -835 591 -834
rect 100 -837 101 -836
rect 306 -837 307 -836
rect 355 -837 356 -836
rect 415 -837 416 -836
rect 359 -839 360 -838
rect 611 -839 612 -838
rect 198 -841 199 -840
rect 359 -841 360 -840
rect 366 -841 367 -840
rect 415 -841 416 -840
rect 366 -843 367 -842
rect 632 -843 633 -842
rect 383 -845 384 -844
rect 492 -845 493 -844
rect 450 -847 451 -846
rect 632 -847 633 -846
rect 450 -849 451 -848
rect 478 -849 479 -848
rect 9 -860 10 -859
rect 593 -860 594 -859
rect 674 -860 675 -859
rect 863 -860 864 -859
rect 16 -862 17 -861
rect 191 -862 192 -861
rect 201 -862 202 -861
rect 278 -862 279 -861
rect 282 -862 283 -861
rect 334 -862 335 -861
rect 338 -862 339 -861
rect 366 -862 367 -861
rect 404 -862 405 -861
rect 562 -862 563 -861
rect 660 -862 661 -861
rect 674 -862 675 -861
rect 831 -862 832 -861
rect 940 -862 941 -861
rect 30 -864 31 -863
rect 222 -864 223 -863
rect 240 -864 241 -863
rect 306 -864 307 -863
rect 317 -864 318 -863
rect 408 -864 409 -863
rect 411 -864 412 -863
rect 786 -864 787 -863
rect 44 -866 45 -865
rect 159 -866 160 -865
rect 163 -866 164 -865
rect 793 -866 794 -865
rect 44 -868 45 -867
rect 352 -868 353 -867
rect 359 -868 360 -867
rect 534 -868 535 -867
rect 562 -868 563 -867
rect 611 -868 612 -867
rect 653 -868 654 -867
rect 660 -868 661 -867
rect 58 -870 59 -869
rect 250 -870 251 -869
rect 261 -870 262 -869
rect 366 -870 367 -869
rect 429 -870 430 -869
rect 814 -870 815 -869
rect 72 -872 73 -871
rect 639 -872 640 -871
rect 653 -872 654 -871
rect 730 -872 731 -871
rect 744 -872 745 -871
rect 814 -872 815 -871
rect 72 -874 73 -873
rect 107 -874 108 -873
rect 121 -874 122 -873
rect 124 -874 125 -873
rect 135 -874 136 -873
rect 264 -874 265 -873
rect 268 -874 269 -873
rect 324 -874 325 -873
rect 327 -874 328 -873
rect 856 -874 857 -873
rect 23 -876 24 -875
rect 135 -876 136 -875
rect 142 -876 143 -875
rect 289 -876 290 -875
rect 317 -876 318 -875
rect 380 -876 381 -875
rect 387 -876 388 -875
rect 429 -876 430 -875
rect 443 -876 444 -875
rect 835 -876 836 -875
rect 23 -878 24 -877
rect 520 -878 521 -877
rect 590 -878 591 -877
rect 786 -878 787 -877
rect 75 -880 76 -879
rect 373 -880 374 -879
rect 387 -880 388 -879
rect 422 -880 423 -879
rect 453 -880 454 -879
rect 527 -880 528 -879
rect 597 -880 598 -879
rect 639 -880 640 -879
rect 730 -880 731 -879
rect 758 -880 759 -879
rect 79 -882 80 -881
rect 296 -882 297 -881
rect 310 -882 311 -881
rect 422 -882 423 -881
rect 457 -882 458 -881
rect 499 -882 500 -881
rect 506 -882 507 -881
rect 709 -882 710 -881
rect 744 -882 745 -881
rect 765 -882 766 -881
rect 79 -884 80 -883
rect 527 -884 528 -883
rect 611 -884 612 -883
rect 625 -884 626 -883
rect 702 -884 703 -883
rect 758 -884 759 -883
rect 765 -884 766 -883
rect 800 -884 801 -883
rect 82 -886 83 -885
rect 485 -886 486 -885
rect 506 -886 507 -885
rect 688 -886 689 -885
rect 709 -886 710 -885
rect 737 -886 738 -885
rect 800 -886 801 -885
rect 828 -886 829 -885
rect 86 -888 87 -887
rect 114 -888 115 -887
rect 142 -888 143 -887
rect 163 -888 164 -887
rect 166 -888 167 -887
rect 177 -888 178 -887
rect 184 -888 185 -887
rect 310 -888 311 -887
rect 345 -888 346 -887
rect 373 -888 374 -887
rect 439 -888 440 -887
rect 499 -888 500 -887
rect 534 -888 535 -887
rect 828 -888 829 -887
rect 30 -890 31 -889
rect 345 -890 346 -889
rect 362 -890 363 -889
rect 436 -890 437 -889
rect 460 -890 461 -889
rect 842 -890 843 -889
rect 51 -892 52 -891
rect 114 -892 115 -891
rect 177 -892 178 -891
rect 226 -892 227 -891
rect 233 -892 234 -891
rect 268 -892 269 -891
rect 464 -892 465 -891
rect 597 -892 598 -891
rect 625 -892 626 -891
rect 695 -892 696 -891
rect 737 -892 738 -891
rect 751 -892 752 -891
rect 842 -892 843 -891
rect 870 -892 871 -891
rect 40 -894 41 -893
rect 233 -894 234 -893
rect 254 -894 255 -893
rect 289 -894 290 -893
rect 467 -894 468 -893
rect 569 -894 570 -893
rect 583 -894 584 -893
rect 702 -894 703 -893
rect 751 -894 752 -893
rect 772 -894 773 -893
rect 51 -896 52 -895
rect 415 -896 416 -895
rect 478 -896 479 -895
rect 516 -896 517 -895
rect 555 -896 556 -895
rect 569 -896 570 -895
rect 681 -896 682 -895
rect 688 -896 689 -895
rect 695 -896 696 -895
rect 779 -896 780 -895
rect 86 -898 87 -897
rect 156 -898 157 -897
rect 170 -898 171 -897
rect 226 -898 227 -897
rect 254 -898 255 -897
rect 299 -898 300 -897
rect 471 -898 472 -897
rect 516 -898 517 -897
rect 541 -898 542 -897
rect 555 -898 556 -897
rect 667 -898 668 -897
rect 681 -898 682 -897
rect 716 -898 717 -897
rect 779 -898 780 -897
rect 93 -900 94 -899
rect 149 -900 150 -899
rect 156 -900 157 -899
rect 282 -900 283 -899
rect 446 -900 447 -899
rect 667 -900 668 -899
rect 716 -900 717 -899
rect 723 -900 724 -899
rect 772 -900 773 -899
rect 821 -900 822 -899
rect 93 -902 94 -901
rect 401 -902 402 -901
rect 471 -902 472 -901
rect 492 -902 493 -901
rect 646 -902 647 -901
rect 723 -902 724 -901
rect 821 -902 822 -901
rect 849 -902 850 -901
rect 54 -904 55 -903
rect 492 -904 493 -903
rect 632 -904 633 -903
rect 646 -904 647 -903
rect 835 -904 836 -903
rect 849 -904 850 -903
rect 100 -906 101 -905
rect 807 -906 808 -905
rect 65 -908 66 -907
rect 100 -908 101 -907
rect 103 -908 104 -907
rect 348 -908 349 -907
rect 401 -908 402 -907
rect 583 -908 584 -907
rect 618 -908 619 -907
rect 632 -908 633 -907
rect 107 -910 108 -909
rect 145 -910 146 -909
rect 191 -910 192 -909
rect 198 -910 199 -909
rect 205 -910 206 -909
rect 359 -910 360 -909
rect 485 -910 486 -909
rect 590 -910 591 -909
rect 604 -910 605 -909
rect 618 -910 619 -909
rect 58 -912 59 -911
rect 198 -912 199 -911
rect 212 -912 213 -911
rect 240 -912 241 -911
rect 261 -912 262 -911
rect 338 -912 339 -911
rect 548 -912 549 -911
rect 604 -912 605 -911
rect 128 -914 129 -913
rect 446 -914 447 -913
rect 128 -916 129 -915
rect 184 -916 185 -915
rect 215 -916 216 -915
rect 520 -916 521 -915
rect 170 -918 171 -917
rect 205 -918 206 -917
rect 219 -918 220 -917
rect 331 -918 332 -917
rect 380 -918 381 -917
rect 548 -918 549 -917
rect 219 -920 220 -919
rect 415 -920 416 -919
rect 275 -922 276 -921
rect 478 -922 479 -921
rect 303 -924 304 -923
rect 807 -924 808 -923
rect 19 -926 20 -925
rect 303 -926 304 -925
rect 331 -926 332 -925
rect 341 -926 342 -925
rect 2 -937 3 -936
rect 233 -937 234 -936
rect 247 -937 248 -936
rect 261 -937 262 -936
rect 275 -937 276 -936
rect 359 -937 360 -936
rect 390 -937 391 -936
rect 723 -937 724 -936
rect 779 -937 780 -936
rect 898 -937 899 -936
rect 9 -939 10 -938
rect 82 -939 83 -938
rect 100 -939 101 -938
rect 338 -939 339 -938
rect 348 -939 349 -938
rect 786 -939 787 -938
rect 814 -939 815 -938
rect 849 -939 850 -938
rect 9 -941 10 -940
rect 128 -941 129 -940
rect 149 -941 150 -940
rect 170 -941 171 -940
rect 173 -941 174 -940
rect 387 -941 388 -940
rect 394 -941 395 -940
rect 436 -941 437 -940
rect 450 -941 451 -940
rect 863 -941 864 -940
rect 16 -943 17 -942
rect 334 -943 335 -942
rect 352 -943 353 -942
rect 499 -943 500 -942
rect 509 -943 510 -942
rect 737 -943 738 -942
rect 786 -943 787 -942
rect 828 -943 829 -942
rect 30 -945 31 -944
rect 296 -945 297 -944
rect 331 -945 332 -944
rect 359 -945 360 -944
rect 397 -945 398 -944
rect 674 -945 675 -944
rect 716 -945 717 -944
rect 779 -945 780 -944
rect 814 -945 815 -944
rect 835 -945 836 -944
rect 37 -947 38 -946
rect 124 -947 125 -946
rect 128 -947 129 -946
rect 222 -947 223 -946
rect 247 -947 248 -946
rect 313 -947 314 -946
rect 331 -947 332 -946
rect 702 -947 703 -946
rect 737 -947 738 -946
rect 744 -947 745 -946
rect 40 -949 41 -948
rect 72 -949 73 -948
rect 79 -949 80 -948
rect 380 -949 381 -948
rect 401 -949 402 -948
rect 667 -949 668 -948
rect 744 -949 745 -948
rect 751 -949 752 -948
rect 44 -951 45 -950
rect 285 -951 286 -950
rect 404 -951 405 -950
rect 408 -951 409 -950
rect 429 -951 430 -950
rect 499 -951 500 -950
rect 513 -951 514 -950
rect 660 -951 661 -950
rect 751 -951 752 -950
rect 807 -951 808 -950
rect 51 -953 52 -952
rect 93 -953 94 -952
rect 117 -953 118 -952
rect 576 -953 577 -952
rect 590 -953 591 -952
rect 821 -953 822 -952
rect 58 -955 59 -954
rect 394 -955 395 -954
rect 408 -955 409 -954
rect 604 -955 605 -954
rect 646 -955 647 -954
rect 667 -955 668 -954
rect 793 -955 794 -954
rect 807 -955 808 -954
rect 58 -957 59 -956
rect 93 -957 94 -956
rect 121 -957 122 -956
rect 194 -957 195 -956
rect 201 -957 202 -956
rect 282 -957 283 -956
rect 303 -957 304 -956
rect 590 -957 591 -956
rect 646 -957 647 -956
rect 688 -957 689 -956
rect 44 -959 45 -958
rect 121 -959 122 -958
rect 152 -959 153 -958
rect 835 -959 836 -958
rect 61 -961 62 -960
rect 411 -961 412 -960
rect 429 -961 430 -960
rect 828 -961 829 -960
rect 65 -963 66 -962
rect 86 -963 87 -962
rect 163 -963 164 -962
rect 485 -963 486 -962
rect 516 -963 517 -962
rect 793 -963 794 -962
rect 65 -965 66 -964
rect 373 -965 374 -964
rect 436 -965 437 -964
rect 632 -965 633 -964
rect 653 -965 654 -964
rect 702 -965 703 -964
rect 72 -967 73 -966
rect 156 -967 157 -966
rect 177 -967 178 -966
rect 303 -967 304 -966
rect 373 -967 374 -966
rect 380 -967 381 -966
rect 443 -967 444 -966
rect 821 -967 822 -966
rect 86 -969 87 -968
rect 317 -969 318 -968
rect 443 -969 444 -968
rect 457 -969 458 -968
rect 464 -969 465 -968
rect 471 -969 472 -968
rect 474 -969 475 -968
rect 723 -969 724 -968
rect 135 -971 136 -970
rect 156 -971 157 -970
rect 177 -971 178 -970
rect 226 -971 227 -970
rect 254 -971 255 -970
rect 296 -971 297 -970
rect 317 -971 318 -970
rect 345 -971 346 -970
rect 446 -971 447 -970
rect 716 -971 717 -970
rect 135 -973 136 -972
rect 201 -973 202 -972
rect 205 -973 206 -972
rect 856 -973 857 -972
rect 170 -975 171 -974
rect 226 -975 227 -974
rect 254 -975 255 -974
rect 453 -975 454 -974
rect 457 -975 458 -974
rect 492 -975 493 -974
rect 541 -975 542 -974
rect 618 -975 619 -974
rect 653 -975 654 -974
rect 681 -975 682 -974
rect 688 -975 689 -974
rect 695 -975 696 -974
rect 191 -977 192 -976
rect 233 -977 234 -976
rect 261 -977 262 -976
rect 268 -977 269 -976
rect 278 -977 279 -976
rect 422 -977 423 -976
rect 450 -977 451 -976
rect 478 -977 479 -976
rect 481 -977 482 -976
rect 541 -977 542 -976
rect 548 -977 549 -976
rect 800 -977 801 -976
rect 208 -979 209 -978
rect 639 -979 640 -978
rect 695 -979 696 -978
rect 730 -979 731 -978
rect 772 -979 773 -978
rect 800 -979 801 -978
rect 212 -981 213 -980
rect 387 -981 388 -980
rect 478 -981 479 -980
rect 660 -981 661 -980
rect 765 -981 766 -980
rect 772 -981 773 -980
rect 215 -983 216 -982
rect 310 -983 311 -982
rect 338 -983 339 -982
rect 548 -983 549 -982
rect 562 -983 563 -982
rect 618 -983 619 -982
rect 639 -983 640 -982
rect 709 -983 710 -982
rect 758 -983 759 -982
rect 765 -983 766 -982
rect 184 -985 185 -984
rect 709 -985 710 -984
rect 758 -985 759 -984
rect 873 -985 874 -984
rect 142 -987 143 -986
rect 184 -987 185 -986
rect 219 -987 220 -986
rect 240 -987 241 -986
rect 268 -987 269 -986
rect 352 -987 353 -986
rect 376 -987 377 -986
rect 730 -987 731 -986
rect 114 -989 115 -988
rect 142 -989 143 -988
rect 240 -989 241 -988
rect 415 -989 416 -988
rect 485 -989 486 -988
rect 569 -989 570 -988
rect 576 -989 577 -988
rect 597 -989 598 -988
rect 114 -991 115 -990
rect 674 -991 675 -990
rect 289 -993 290 -992
rect 632 -993 633 -992
rect 289 -995 290 -994
rect 324 -995 325 -994
rect 345 -995 346 -994
rect 366 -995 367 -994
rect 404 -995 405 -994
rect 415 -995 416 -994
rect 555 -995 556 -994
rect 562 -995 563 -994
rect 583 -995 584 -994
rect 681 -995 682 -994
rect 23 -997 24 -996
rect 366 -997 367 -996
rect 555 -997 556 -996
rect 625 -997 626 -996
rect 23 -999 24 -998
rect 107 -999 108 -998
rect 299 -999 300 -998
rect 492 -999 493 -998
rect 558 -999 559 -998
rect 569 -999 570 -998
rect 597 -999 598 -998
rect 859 -999 860 -998
rect 107 -1001 108 -1000
rect 131 -1001 132 -1000
rect 324 -1001 325 -1000
rect 506 -1001 507 -1000
rect 611 -1001 612 -1000
rect 625 -1001 626 -1000
rect 425 -1003 426 -1002
rect 611 -1003 612 -1002
rect 506 -1005 507 -1004
rect 604 -1005 605 -1004
rect 2 -1016 3 -1015
rect 411 -1016 412 -1015
rect 422 -1016 423 -1015
rect 541 -1016 542 -1015
rect 551 -1016 552 -1015
rect 723 -1016 724 -1015
rect 786 -1016 787 -1015
rect 856 -1016 857 -1015
rect 863 -1016 864 -1015
rect 919 -1016 920 -1015
rect 9 -1018 10 -1017
rect 170 -1018 171 -1017
rect 212 -1018 213 -1017
rect 338 -1018 339 -1017
rect 341 -1018 342 -1017
rect 492 -1018 493 -1017
rect 502 -1018 503 -1017
rect 842 -1018 843 -1017
rect 849 -1018 850 -1017
rect 912 -1018 913 -1017
rect 16 -1020 17 -1019
rect 205 -1020 206 -1019
rect 212 -1020 213 -1019
rect 401 -1020 402 -1019
rect 404 -1020 405 -1019
rect 485 -1020 486 -1019
rect 492 -1020 493 -1019
rect 884 -1020 885 -1019
rect 898 -1020 899 -1019
rect 926 -1020 927 -1019
rect 19 -1022 20 -1021
rect 786 -1022 787 -1021
rect 800 -1022 801 -1021
rect 877 -1022 878 -1021
rect 23 -1024 24 -1023
rect 26 -1024 27 -1023
rect 30 -1024 31 -1023
rect 198 -1024 199 -1023
rect 205 -1024 206 -1023
rect 261 -1024 262 -1023
rect 303 -1024 304 -1023
rect 467 -1024 468 -1023
rect 478 -1024 479 -1023
rect 639 -1024 640 -1023
rect 642 -1024 643 -1023
rect 842 -1024 843 -1023
rect 23 -1026 24 -1025
rect 156 -1026 157 -1025
rect 166 -1026 167 -1025
rect 233 -1026 234 -1025
rect 261 -1026 262 -1025
rect 558 -1026 559 -1025
rect 590 -1026 591 -1025
rect 891 -1026 892 -1025
rect 33 -1028 34 -1027
rect 709 -1028 710 -1027
rect 772 -1028 773 -1027
rect 800 -1028 801 -1027
rect 807 -1028 808 -1027
rect 870 -1028 871 -1027
rect 37 -1030 38 -1029
rect 191 -1030 192 -1029
rect 219 -1030 220 -1029
rect 282 -1030 283 -1029
rect 303 -1030 304 -1029
rect 324 -1030 325 -1029
rect 331 -1030 332 -1029
rect 730 -1030 731 -1029
rect 772 -1030 773 -1029
rect 859 -1030 860 -1029
rect 37 -1032 38 -1031
rect 86 -1032 87 -1031
rect 93 -1032 94 -1031
rect 436 -1032 437 -1031
rect 439 -1032 440 -1031
rect 478 -1032 479 -1031
rect 506 -1032 507 -1031
rect 611 -1032 612 -1031
rect 660 -1032 661 -1031
rect 723 -1032 724 -1031
rect 779 -1032 780 -1031
rect 849 -1032 850 -1031
rect 54 -1034 55 -1033
rect 86 -1034 87 -1033
rect 107 -1034 108 -1033
rect 408 -1034 409 -1033
rect 415 -1034 416 -1033
rect 485 -1034 486 -1033
rect 513 -1034 514 -1033
rect 751 -1034 752 -1033
rect 821 -1034 822 -1033
rect 940 -1034 941 -1033
rect 58 -1036 59 -1035
rect 159 -1036 160 -1035
rect 163 -1036 164 -1035
rect 513 -1036 514 -1035
rect 516 -1036 517 -1035
rect 597 -1036 598 -1035
rect 604 -1036 605 -1035
rect 614 -1036 615 -1035
rect 681 -1036 682 -1035
rect 730 -1036 731 -1035
rect 828 -1036 829 -1035
rect 898 -1036 899 -1035
rect 65 -1038 66 -1037
rect 415 -1038 416 -1037
rect 432 -1038 433 -1037
rect 443 -1038 444 -1037
rect 446 -1038 447 -1037
rect 807 -1038 808 -1037
rect 835 -1038 836 -1037
rect 905 -1038 906 -1037
rect 65 -1040 66 -1039
rect 254 -1040 255 -1039
rect 278 -1040 279 -1039
rect 282 -1040 283 -1039
rect 289 -1040 290 -1039
rect 506 -1040 507 -1039
rect 527 -1040 528 -1039
rect 590 -1040 591 -1039
rect 604 -1040 605 -1039
rect 744 -1040 745 -1039
rect 72 -1042 73 -1041
rect 114 -1042 115 -1041
rect 121 -1042 122 -1041
rect 142 -1042 143 -1041
rect 163 -1042 164 -1041
rect 814 -1042 815 -1041
rect 72 -1044 73 -1043
rect 149 -1044 150 -1043
rect 152 -1044 153 -1043
rect 814 -1044 815 -1043
rect 79 -1046 80 -1045
rect 310 -1046 311 -1045
rect 317 -1046 318 -1045
rect 401 -1046 402 -1045
rect 453 -1046 454 -1045
rect 572 -1046 573 -1045
rect 576 -1046 577 -1045
rect 660 -1046 661 -1045
rect 674 -1046 675 -1045
rect 744 -1046 745 -1045
rect 79 -1048 80 -1047
rect 275 -1048 276 -1047
rect 296 -1048 297 -1047
rect 324 -1048 325 -1047
rect 352 -1048 353 -1047
rect 394 -1048 395 -1047
rect 499 -1048 500 -1047
rect 828 -1048 829 -1047
rect 103 -1050 104 -1049
rect 114 -1050 115 -1049
rect 128 -1050 129 -1049
rect 667 -1050 668 -1049
rect 688 -1050 689 -1049
rect 821 -1050 822 -1049
rect 107 -1052 108 -1051
rect 117 -1052 118 -1051
rect 128 -1052 129 -1051
rect 334 -1052 335 -1051
rect 352 -1052 353 -1051
rect 583 -1052 584 -1051
rect 614 -1052 615 -1051
rect 674 -1052 675 -1051
rect 695 -1052 696 -1051
rect 863 -1052 864 -1051
rect 135 -1054 136 -1053
rect 142 -1054 143 -1053
rect 170 -1054 171 -1053
rect 268 -1054 269 -1053
rect 275 -1054 276 -1053
rect 450 -1054 451 -1053
rect 464 -1054 465 -1053
rect 499 -1054 500 -1053
rect 520 -1054 521 -1053
rect 576 -1054 577 -1053
rect 716 -1054 717 -1053
rect 779 -1054 780 -1053
rect 177 -1056 178 -1055
rect 233 -1056 234 -1055
rect 243 -1056 244 -1055
rect 289 -1056 290 -1055
rect 317 -1056 318 -1055
rect 495 -1056 496 -1055
rect 527 -1056 528 -1055
rect 681 -1056 682 -1055
rect 737 -1056 738 -1055
rect 835 -1056 836 -1055
rect 100 -1058 101 -1057
rect 177 -1058 178 -1057
rect 184 -1058 185 -1057
rect 254 -1058 255 -1057
rect 268 -1058 269 -1057
rect 348 -1058 349 -1057
rect 359 -1058 360 -1057
rect 373 -1058 374 -1057
rect 380 -1058 381 -1057
rect 390 -1058 391 -1057
rect 429 -1058 430 -1057
rect 520 -1058 521 -1057
rect 534 -1058 535 -1057
rect 695 -1058 696 -1057
rect 191 -1060 192 -1059
rect 222 -1060 223 -1059
rect 226 -1060 227 -1059
rect 541 -1060 542 -1059
rect 565 -1060 566 -1059
rect 667 -1060 668 -1059
rect 44 -1062 45 -1061
rect 222 -1062 223 -1061
rect 226 -1062 227 -1061
rect 240 -1062 241 -1061
rect 247 -1062 248 -1061
rect 296 -1062 297 -1061
rect 345 -1062 346 -1061
rect 380 -1062 381 -1061
rect 387 -1062 388 -1061
rect 632 -1062 633 -1061
rect 646 -1062 647 -1061
rect 737 -1062 738 -1061
rect 44 -1064 45 -1063
rect 51 -1064 52 -1063
rect 201 -1064 202 -1063
rect 331 -1064 332 -1063
rect 345 -1064 346 -1063
rect 758 -1064 759 -1063
rect 359 -1066 360 -1065
rect 537 -1066 538 -1065
rect 548 -1066 549 -1065
rect 632 -1066 633 -1065
rect 653 -1066 654 -1065
rect 716 -1066 717 -1065
rect 758 -1066 759 -1065
rect 765 -1066 766 -1065
rect 184 -1068 185 -1067
rect 548 -1068 549 -1067
rect 562 -1068 563 -1067
rect 646 -1068 647 -1067
rect 366 -1070 367 -1069
rect 611 -1070 612 -1069
rect 625 -1070 626 -1069
rect 765 -1070 766 -1069
rect 366 -1072 367 -1071
rect 530 -1072 531 -1071
rect 534 -1072 535 -1071
rect 751 -1072 752 -1071
rect 376 -1074 377 -1073
rect 653 -1074 654 -1073
rect 390 -1076 391 -1075
rect 471 -1076 472 -1075
rect 562 -1076 563 -1075
rect 709 -1076 710 -1075
rect 429 -1078 430 -1077
rect 457 -1078 458 -1077
rect 569 -1078 570 -1077
rect 597 -1078 598 -1077
rect 607 -1078 608 -1077
rect 625 -1078 626 -1077
rect 194 -1080 195 -1079
rect 457 -1080 458 -1079
rect 450 -1082 451 -1081
rect 688 -1082 689 -1081
rect 9 -1093 10 -1092
rect 786 -1093 787 -1092
rect 884 -1093 885 -1092
rect 975 -1093 976 -1092
rect 982 -1093 983 -1092
rect 989 -1093 990 -1092
rect 9 -1095 10 -1094
rect 170 -1095 171 -1094
rect 198 -1095 199 -1094
rect 226 -1095 227 -1094
rect 240 -1095 241 -1094
rect 282 -1095 283 -1094
rect 317 -1095 318 -1094
rect 443 -1095 444 -1094
rect 446 -1095 447 -1094
rect 891 -1095 892 -1094
rect 898 -1095 899 -1094
rect 968 -1095 969 -1094
rect 16 -1097 17 -1096
rect 579 -1097 580 -1096
rect 642 -1097 643 -1096
rect 849 -1097 850 -1096
rect 856 -1097 857 -1096
rect 898 -1097 899 -1096
rect 912 -1097 913 -1096
rect 947 -1097 948 -1096
rect 16 -1099 17 -1098
rect 30 -1099 31 -1098
rect 44 -1099 45 -1098
rect 96 -1099 97 -1098
rect 103 -1099 104 -1098
rect 716 -1099 717 -1098
rect 828 -1099 829 -1098
rect 884 -1099 885 -1098
rect 30 -1101 31 -1100
rect 37 -1101 38 -1100
rect 44 -1101 45 -1100
rect 205 -1101 206 -1100
rect 226 -1101 227 -1100
rect 310 -1101 311 -1100
rect 345 -1101 346 -1100
rect 366 -1101 367 -1100
rect 387 -1101 388 -1100
rect 408 -1101 409 -1100
rect 436 -1101 437 -1100
rect 439 -1101 440 -1100
rect 450 -1101 451 -1100
rect 639 -1101 640 -1100
rect 667 -1101 668 -1100
rect 933 -1101 934 -1100
rect 37 -1103 38 -1102
rect 268 -1103 269 -1102
rect 275 -1103 276 -1102
rect 320 -1103 321 -1102
rect 348 -1103 349 -1102
rect 415 -1103 416 -1102
rect 436 -1103 437 -1102
rect 492 -1103 493 -1102
rect 506 -1103 507 -1102
rect 534 -1103 535 -1102
rect 544 -1103 545 -1102
rect 821 -1103 822 -1102
rect 842 -1103 843 -1102
rect 891 -1103 892 -1102
rect 51 -1105 52 -1104
rect 86 -1105 87 -1104
rect 93 -1105 94 -1104
rect 912 -1105 913 -1104
rect 58 -1107 59 -1106
rect 65 -1107 66 -1106
rect 72 -1107 73 -1106
rect 152 -1107 153 -1106
rect 156 -1107 157 -1106
rect 177 -1107 178 -1106
rect 198 -1107 199 -1106
rect 555 -1107 556 -1106
rect 558 -1107 559 -1106
rect 863 -1107 864 -1106
rect 58 -1109 59 -1108
rect 254 -1109 255 -1108
rect 268 -1109 269 -1108
rect 296 -1109 297 -1108
rect 303 -1109 304 -1108
rect 310 -1109 311 -1108
rect 355 -1109 356 -1108
rect 695 -1109 696 -1108
rect 702 -1109 703 -1108
rect 856 -1109 857 -1108
rect 863 -1109 864 -1108
rect 929 -1109 930 -1108
rect 72 -1111 73 -1110
rect 201 -1111 202 -1110
rect 205 -1111 206 -1110
rect 362 -1111 363 -1110
rect 366 -1111 367 -1110
rect 632 -1111 633 -1110
rect 684 -1111 685 -1110
rect 877 -1111 878 -1110
rect 82 -1113 83 -1112
rect 219 -1113 220 -1112
rect 247 -1113 248 -1112
rect 289 -1113 290 -1112
rect 303 -1113 304 -1112
rect 324 -1113 325 -1112
rect 355 -1113 356 -1112
rect 415 -1113 416 -1112
rect 439 -1113 440 -1112
rect 492 -1113 493 -1112
rect 520 -1113 521 -1112
rect 604 -1113 605 -1112
rect 607 -1113 608 -1112
rect 667 -1113 668 -1112
rect 702 -1113 703 -1112
rect 716 -1113 717 -1112
rect 751 -1113 752 -1112
rect 842 -1113 843 -1112
rect 849 -1113 850 -1112
rect 961 -1113 962 -1112
rect 86 -1115 87 -1114
rect 107 -1115 108 -1114
rect 128 -1115 129 -1114
rect 296 -1115 297 -1114
rect 331 -1115 332 -1114
rect 604 -1115 605 -1114
rect 758 -1115 759 -1114
rect 821 -1115 822 -1114
rect 103 -1117 104 -1116
rect 254 -1117 255 -1116
rect 278 -1117 279 -1116
rect 751 -1117 752 -1116
rect 800 -1117 801 -1116
rect 828 -1117 829 -1116
rect 107 -1119 108 -1118
rect 114 -1119 115 -1118
rect 128 -1119 129 -1118
rect 142 -1119 143 -1118
rect 152 -1119 153 -1118
rect 506 -1119 507 -1118
rect 527 -1119 528 -1118
rect 737 -1119 738 -1118
rect 114 -1121 115 -1120
rect 380 -1121 381 -1120
rect 390 -1121 391 -1120
rect 919 -1121 920 -1120
rect 135 -1123 136 -1122
rect 786 -1123 787 -1122
rect 870 -1123 871 -1122
rect 919 -1123 920 -1122
rect 135 -1125 136 -1124
rect 520 -1125 521 -1124
rect 530 -1125 531 -1124
rect 905 -1125 906 -1124
rect 138 -1127 139 -1126
rect 233 -1127 234 -1126
rect 250 -1127 251 -1126
rect 695 -1127 696 -1126
rect 772 -1127 773 -1126
rect 870 -1127 871 -1126
rect 23 -1129 24 -1128
rect 233 -1129 234 -1128
rect 282 -1129 283 -1128
rect 527 -1129 528 -1128
rect 562 -1129 563 -1128
rect 814 -1129 815 -1128
rect 93 -1131 94 -1130
rect 772 -1131 773 -1130
rect 793 -1131 794 -1130
rect 905 -1131 906 -1130
rect 142 -1133 143 -1132
rect 429 -1133 430 -1132
rect 453 -1133 454 -1132
rect 688 -1133 689 -1132
rect 709 -1133 710 -1132
rect 814 -1133 815 -1132
rect 163 -1135 164 -1134
rect 261 -1135 262 -1134
rect 289 -1135 290 -1134
rect 359 -1135 360 -1134
rect 380 -1135 381 -1134
rect 394 -1135 395 -1134
rect 422 -1135 423 -1134
rect 688 -1135 689 -1134
rect 166 -1137 167 -1136
rect 877 -1137 878 -1136
rect 177 -1139 178 -1138
rect 191 -1139 192 -1138
rect 261 -1139 262 -1138
rect 485 -1139 486 -1138
rect 562 -1139 563 -1138
rect 926 -1139 927 -1138
rect 184 -1141 185 -1140
rect 429 -1141 430 -1140
rect 464 -1141 465 -1140
rect 835 -1141 836 -1140
rect 170 -1143 171 -1142
rect 184 -1143 185 -1142
rect 191 -1143 192 -1142
rect 212 -1143 213 -1142
rect 324 -1143 325 -1142
rect 453 -1143 454 -1142
rect 485 -1143 486 -1142
rect 509 -1143 510 -1142
rect 569 -1143 570 -1142
rect 800 -1143 801 -1142
rect 331 -1145 332 -1144
rect 590 -1145 591 -1144
rect 618 -1145 619 -1144
rect 758 -1145 759 -1144
rect 338 -1147 339 -1146
rect 422 -1147 423 -1146
rect 513 -1147 514 -1146
rect 569 -1147 570 -1146
rect 572 -1147 573 -1146
rect 765 -1147 766 -1146
rect 222 -1149 223 -1148
rect 765 -1149 766 -1148
rect 222 -1151 223 -1150
rect 394 -1151 395 -1150
rect 401 -1151 402 -1150
rect 513 -1151 514 -1150
rect 576 -1151 577 -1150
rect 632 -1151 633 -1150
rect 646 -1151 647 -1150
rect 709 -1151 710 -1150
rect 730 -1151 731 -1150
rect 835 -1151 836 -1150
rect 338 -1153 339 -1152
rect 373 -1153 374 -1152
rect 583 -1153 584 -1152
rect 639 -1153 640 -1152
rect 646 -1153 647 -1152
rect 681 -1153 682 -1152
rect 359 -1155 360 -1154
rect 779 -1155 780 -1154
rect 373 -1157 374 -1156
rect 450 -1157 451 -1156
rect 548 -1157 549 -1156
rect 681 -1157 682 -1156
rect 744 -1157 745 -1156
rect 779 -1157 780 -1156
rect 79 -1159 80 -1158
rect 744 -1159 745 -1158
rect 79 -1161 80 -1160
rect 121 -1161 122 -1160
rect 425 -1161 426 -1160
rect 583 -1161 584 -1160
rect 618 -1161 619 -1160
rect 723 -1161 724 -1160
rect 625 -1163 626 -1162
rect 793 -1163 794 -1162
rect 611 -1165 612 -1164
rect 625 -1165 626 -1164
rect 653 -1165 654 -1164
rect 723 -1165 724 -1164
rect 597 -1167 598 -1166
rect 611 -1167 612 -1166
rect 656 -1167 657 -1166
rect 926 -1167 927 -1166
rect 499 -1169 500 -1168
rect 597 -1169 598 -1168
rect 660 -1169 661 -1168
rect 730 -1169 731 -1168
rect 478 -1171 479 -1170
rect 499 -1171 500 -1170
rect 541 -1171 542 -1170
rect 660 -1171 661 -1170
rect 674 -1171 675 -1170
rect 737 -1171 738 -1170
rect 401 -1173 402 -1172
rect 478 -1173 479 -1172
rect 541 -1173 542 -1172
rect 590 -1173 591 -1172
rect 457 -1175 458 -1174
rect 674 -1175 675 -1174
rect 457 -1177 458 -1176
rect 471 -1177 472 -1176
rect 212 -1179 213 -1178
rect 471 -1179 472 -1178
rect 5 -1190 6 -1189
rect 219 -1190 220 -1189
rect 222 -1190 223 -1189
rect 674 -1190 675 -1189
rect 719 -1190 720 -1189
rect 828 -1190 829 -1189
rect 940 -1190 941 -1189
rect 964 -1190 965 -1189
rect 975 -1190 976 -1189
rect 982 -1190 983 -1189
rect 985 -1190 986 -1189
rect 1010 -1190 1011 -1189
rect 9 -1192 10 -1191
rect 212 -1192 213 -1191
rect 215 -1192 216 -1191
rect 723 -1192 724 -1191
rect 737 -1192 738 -1191
rect 740 -1192 741 -1191
rect 751 -1192 752 -1191
rect 954 -1192 955 -1191
rect 989 -1192 990 -1191
rect 1003 -1192 1004 -1191
rect 16 -1194 17 -1193
rect 215 -1194 216 -1193
rect 254 -1194 255 -1193
rect 306 -1194 307 -1193
rect 341 -1194 342 -1193
rect 618 -1194 619 -1193
rect 625 -1194 626 -1193
rect 716 -1194 717 -1193
rect 723 -1194 724 -1193
rect 744 -1194 745 -1193
rect 800 -1194 801 -1193
rect 828 -1194 829 -1193
rect 968 -1194 969 -1193
rect 989 -1194 990 -1193
rect 16 -1196 17 -1195
rect 177 -1196 178 -1195
rect 201 -1196 202 -1195
rect 765 -1196 766 -1195
rect 800 -1196 801 -1195
rect 884 -1196 885 -1195
rect 912 -1196 913 -1195
rect 968 -1196 969 -1195
rect 44 -1198 45 -1197
rect 313 -1198 314 -1197
rect 352 -1198 353 -1197
rect 485 -1198 486 -1197
rect 506 -1198 507 -1197
rect 898 -1198 899 -1197
rect 58 -1200 59 -1199
rect 173 -1200 174 -1199
rect 254 -1200 255 -1199
rect 362 -1200 363 -1199
rect 373 -1200 374 -1199
rect 422 -1200 423 -1199
rect 429 -1200 430 -1199
rect 765 -1200 766 -1199
rect 814 -1200 815 -1199
rect 996 -1200 997 -1199
rect 58 -1202 59 -1201
rect 460 -1202 461 -1201
rect 464 -1202 465 -1201
rect 793 -1202 794 -1201
rect 814 -1202 815 -1201
rect 926 -1202 927 -1201
rect 72 -1204 73 -1203
rect 198 -1204 199 -1203
rect 268 -1204 269 -1203
rect 317 -1204 318 -1203
rect 355 -1204 356 -1203
rect 366 -1204 367 -1203
rect 411 -1204 412 -1203
rect 688 -1204 689 -1203
rect 737 -1204 738 -1203
rect 856 -1204 857 -1203
rect 65 -1206 66 -1205
rect 366 -1206 367 -1205
rect 411 -1206 412 -1205
rect 681 -1206 682 -1205
rect 842 -1206 843 -1205
rect 856 -1206 857 -1205
rect 65 -1208 66 -1207
rect 499 -1208 500 -1207
rect 534 -1208 535 -1207
rect 688 -1208 689 -1207
rect 786 -1208 787 -1207
rect 842 -1208 843 -1207
rect 849 -1208 850 -1207
rect 912 -1208 913 -1207
rect 86 -1210 87 -1209
rect 121 -1210 122 -1209
rect 135 -1210 136 -1209
rect 226 -1210 227 -1209
rect 268 -1210 269 -1209
rect 303 -1210 304 -1209
rect 310 -1210 311 -1209
rect 373 -1210 374 -1209
rect 429 -1210 430 -1209
rect 562 -1210 563 -1209
rect 579 -1210 580 -1209
rect 975 -1210 976 -1209
rect 79 -1212 80 -1211
rect 135 -1212 136 -1211
rect 142 -1212 143 -1211
rect 320 -1212 321 -1211
rect 359 -1212 360 -1211
rect 807 -1212 808 -1211
rect 30 -1214 31 -1213
rect 142 -1214 143 -1213
rect 149 -1214 150 -1213
rect 331 -1214 332 -1213
rect 446 -1214 447 -1213
rect 709 -1214 710 -1213
rect 772 -1214 773 -1213
rect 786 -1214 787 -1213
rect 30 -1216 31 -1215
rect 408 -1216 409 -1215
rect 450 -1216 451 -1215
rect 597 -1216 598 -1215
rect 604 -1216 605 -1215
rect 674 -1216 675 -1215
rect 740 -1216 741 -1215
rect 772 -1216 773 -1215
rect 779 -1216 780 -1215
rect 849 -1216 850 -1215
rect 12 -1218 13 -1217
rect 408 -1218 409 -1217
rect 436 -1218 437 -1217
rect 450 -1218 451 -1217
rect 453 -1218 454 -1217
rect 758 -1218 759 -1217
rect 79 -1220 80 -1219
rect 324 -1220 325 -1219
rect 464 -1220 465 -1219
rect 933 -1220 934 -1219
rect 86 -1222 87 -1221
rect 152 -1222 153 -1221
rect 163 -1222 164 -1221
rect 198 -1222 199 -1221
rect 226 -1222 227 -1221
rect 495 -1222 496 -1221
rect 520 -1222 521 -1221
rect 562 -1222 563 -1221
rect 583 -1222 584 -1221
rect 926 -1222 927 -1221
rect 93 -1224 94 -1223
rect 205 -1224 206 -1223
rect 233 -1224 234 -1223
rect 324 -1224 325 -1223
rect 467 -1224 468 -1223
rect 653 -1224 654 -1223
rect 656 -1224 657 -1223
rect 905 -1224 906 -1223
rect 37 -1226 38 -1225
rect 205 -1226 206 -1225
rect 233 -1226 234 -1225
rect 401 -1226 402 -1225
rect 474 -1226 475 -1225
rect 520 -1226 521 -1225
rect 527 -1226 528 -1225
rect 534 -1226 535 -1225
rect 541 -1226 542 -1225
rect 957 -1226 958 -1225
rect 93 -1228 94 -1227
rect 632 -1228 633 -1227
rect 635 -1228 636 -1227
rect 807 -1228 808 -1227
rect 877 -1228 878 -1227
rect 933 -1228 934 -1227
rect 96 -1230 97 -1229
rect 163 -1230 164 -1229
rect 170 -1230 171 -1229
rect 177 -1230 178 -1229
rect 275 -1230 276 -1229
rect 744 -1230 745 -1229
rect 758 -1230 759 -1229
rect 870 -1230 871 -1229
rect 877 -1230 878 -1229
rect 947 -1230 948 -1229
rect 96 -1232 97 -1231
rect 331 -1232 332 -1231
rect 401 -1232 402 -1231
rect 467 -1232 468 -1231
rect 471 -1232 472 -1231
rect 541 -1232 542 -1231
rect 544 -1232 545 -1231
rect 898 -1232 899 -1231
rect 100 -1234 101 -1233
rect 156 -1234 157 -1233
rect 285 -1234 286 -1233
rect 492 -1234 493 -1233
rect 555 -1234 556 -1233
rect 625 -1234 626 -1233
rect 639 -1234 640 -1233
rect 709 -1234 710 -1233
rect 863 -1234 864 -1233
rect 870 -1234 871 -1233
rect 103 -1236 104 -1235
rect 695 -1236 696 -1235
rect 107 -1238 108 -1237
rect 121 -1238 122 -1237
rect 128 -1238 129 -1237
rect 156 -1238 157 -1237
rect 296 -1238 297 -1237
rect 436 -1238 437 -1237
rect 457 -1238 458 -1237
rect 527 -1238 528 -1237
rect 583 -1238 584 -1237
rect 590 -1238 591 -1237
rect 597 -1238 598 -1237
rect 695 -1238 696 -1237
rect 44 -1240 45 -1239
rect 128 -1240 129 -1239
rect 149 -1240 150 -1239
rect 184 -1240 185 -1239
rect 296 -1240 297 -1239
rect 345 -1240 346 -1239
rect 394 -1240 395 -1239
rect 639 -1240 640 -1239
rect 646 -1240 647 -1239
rect 793 -1240 794 -1239
rect 110 -1242 111 -1241
rect 191 -1242 192 -1241
rect 303 -1242 304 -1241
rect 425 -1242 426 -1241
rect 457 -1242 458 -1241
rect 730 -1242 731 -1241
rect 114 -1244 115 -1243
rect 576 -1244 577 -1243
rect 604 -1244 605 -1243
rect 751 -1244 752 -1243
rect 51 -1246 52 -1245
rect 114 -1246 115 -1245
rect 184 -1246 185 -1245
rect 275 -1246 276 -1245
rect 338 -1246 339 -1245
rect 394 -1246 395 -1245
rect 471 -1246 472 -1245
rect 961 -1246 962 -1245
rect 51 -1248 52 -1247
rect 261 -1248 262 -1247
rect 345 -1248 346 -1247
rect 380 -1248 381 -1247
rect 478 -1248 479 -1247
rect 905 -1248 906 -1247
rect 191 -1250 192 -1249
rect 222 -1250 223 -1249
rect 261 -1250 262 -1249
rect 289 -1250 290 -1249
rect 380 -1250 381 -1249
rect 590 -1250 591 -1249
rect 607 -1250 608 -1249
rect 821 -1250 822 -1249
rect 891 -1250 892 -1249
rect 961 -1250 962 -1249
rect 212 -1252 213 -1251
rect 730 -1252 731 -1251
rect 835 -1252 836 -1251
rect 891 -1252 892 -1251
rect 289 -1254 290 -1253
rect 387 -1254 388 -1253
rect 443 -1254 444 -1253
rect 478 -1254 479 -1253
rect 492 -1254 493 -1253
rect 779 -1254 780 -1253
rect 310 -1256 311 -1255
rect 835 -1256 836 -1255
rect 387 -1258 388 -1257
rect 415 -1258 416 -1257
rect 443 -1258 444 -1257
rect 485 -1258 486 -1257
rect 513 -1258 514 -1257
rect 555 -1258 556 -1257
rect 600 -1258 601 -1257
rect 821 -1258 822 -1257
rect 282 -1260 283 -1259
rect 415 -1260 416 -1259
rect 513 -1260 514 -1259
rect 548 -1260 549 -1259
rect 646 -1260 647 -1259
rect 943 -1260 944 -1259
rect 240 -1262 241 -1261
rect 282 -1262 283 -1261
rect 548 -1262 549 -1261
rect 569 -1262 570 -1261
rect 656 -1262 657 -1261
rect 919 -1262 920 -1261
rect 40 -1264 41 -1263
rect 240 -1264 241 -1263
rect 569 -1264 570 -1263
rect 919 -1264 920 -1263
rect 660 -1266 661 -1265
rect 863 -1266 864 -1265
rect 660 -1268 661 -1267
rect 702 -1268 703 -1267
rect 124 -1270 125 -1269
rect 702 -1270 703 -1269
rect 667 -1272 668 -1271
rect 884 -1272 885 -1271
rect 670 -1274 671 -1273
rect 947 -1274 948 -1273
rect 9 -1285 10 -1284
rect 30 -1285 31 -1284
rect 37 -1285 38 -1284
rect 149 -1285 150 -1284
rect 170 -1285 171 -1284
rect 219 -1285 220 -1284
rect 222 -1285 223 -1284
rect 289 -1285 290 -1284
rect 310 -1285 311 -1284
rect 576 -1285 577 -1284
rect 579 -1285 580 -1284
rect 926 -1285 927 -1284
rect 943 -1285 944 -1284
rect 1010 -1285 1011 -1284
rect 30 -1287 31 -1286
rect 688 -1287 689 -1286
rect 971 -1287 972 -1286
rect 989 -1287 990 -1286
rect 44 -1289 45 -1288
rect 215 -1289 216 -1288
rect 226 -1289 227 -1288
rect 506 -1289 507 -1288
rect 509 -1289 510 -1288
rect 695 -1289 696 -1288
rect 940 -1289 941 -1288
rect 989 -1289 990 -1288
rect 44 -1291 45 -1290
rect 86 -1291 87 -1290
rect 89 -1291 90 -1290
rect 453 -1291 454 -1290
rect 457 -1291 458 -1290
rect 541 -1291 542 -1290
rect 569 -1291 570 -1290
rect 954 -1291 955 -1290
rect 51 -1293 52 -1292
rect 341 -1293 342 -1292
rect 408 -1293 409 -1292
rect 436 -1293 437 -1292
rect 446 -1293 447 -1292
rect 492 -1293 493 -1292
rect 499 -1293 500 -1292
rect 709 -1293 710 -1292
rect 954 -1293 955 -1292
rect 1003 -1293 1004 -1292
rect 51 -1295 52 -1294
rect 96 -1295 97 -1294
rect 124 -1295 125 -1294
rect 226 -1295 227 -1294
rect 240 -1295 241 -1294
rect 289 -1295 290 -1294
rect 310 -1295 311 -1294
rect 317 -1295 318 -1294
rect 352 -1295 353 -1294
rect 499 -1295 500 -1294
rect 569 -1295 570 -1294
rect 583 -1295 584 -1294
rect 597 -1295 598 -1294
rect 611 -1295 612 -1294
rect 618 -1295 619 -1294
rect 919 -1295 920 -1294
rect 58 -1297 59 -1296
rect 173 -1297 174 -1296
rect 184 -1297 185 -1296
rect 863 -1297 864 -1296
rect 919 -1297 920 -1296
rect 975 -1297 976 -1296
rect 61 -1299 62 -1298
rect 107 -1299 108 -1298
rect 135 -1299 136 -1298
rect 184 -1299 185 -1298
rect 198 -1299 199 -1298
rect 219 -1299 220 -1298
rect 229 -1299 230 -1298
rect 863 -1299 864 -1298
rect 65 -1301 66 -1300
rect 352 -1301 353 -1300
rect 387 -1301 388 -1300
rect 408 -1301 409 -1300
rect 411 -1301 412 -1300
rect 898 -1301 899 -1300
rect 65 -1303 66 -1302
rect 380 -1303 381 -1302
rect 387 -1303 388 -1302
rect 555 -1303 556 -1302
rect 576 -1303 577 -1302
rect 912 -1303 913 -1302
rect 72 -1305 73 -1304
rect 128 -1305 129 -1304
rect 149 -1305 150 -1304
rect 261 -1305 262 -1304
rect 282 -1305 283 -1304
rect 359 -1305 360 -1304
rect 415 -1305 416 -1304
rect 464 -1305 465 -1304
rect 467 -1305 468 -1304
rect 488 -1305 489 -1304
rect 502 -1305 503 -1304
rect 583 -1305 584 -1304
rect 632 -1305 633 -1304
rect 660 -1305 661 -1304
rect 667 -1305 668 -1304
rect 891 -1305 892 -1304
rect 898 -1305 899 -1304
rect 982 -1305 983 -1304
rect 16 -1307 17 -1306
rect 261 -1307 262 -1306
rect 296 -1307 297 -1306
rect 359 -1307 360 -1306
rect 366 -1307 367 -1306
rect 464 -1307 465 -1306
rect 471 -1307 472 -1306
rect 793 -1307 794 -1306
rect 16 -1309 17 -1308
rect 110 -1309 111 -1308
rect 114 -1309 115 -1308
rect 135 -1309 136 -1308
rect 163 -1309 164 -1308
rect 282 -1309 283 -1308
rect 303 -1309 304 -1308
rect 471 -1309 472 -1308
rect 474 -1309 475 -1308
rect 646 -1309 647 -1308
rect 653 -1309 654 -1308
rect 891 -1309 892 -1308
rect 72 -1311 73 -1310
rect 730 -1311 731 -1310
rect 793 -1311 794 -1310
rect 849 -1311 850 -1310
rect 12 -1313 13 -1312
rect 730 -1313 731 -1312
rect 93 -1315 94 -1314
rect 530 -1315 531 -1314
rect 548 -1315 549 -1314
rect 611 -1315 612 -1314
rect 646 -1315 647 -1314
rect 716 -1315 717 -1314
rect 114 -1317 115 -1316
rect 121 -1317 122 -1316
rect 128 -1317 129 -1316
rect 254 -1317 255 -1316
rect 317 -1317 318 -1316
rect 324 -1317 325 -1316
rect 331 -1317 332 -1316
rect 618 -1317 619 -1316
rect 653 -1317 654 -1316
rect 702 -1317 703 -1316
rect 709 -1317 710 -1316
rect 835 -1317 836 -1316
rect 121 -1319 122 -1318
rect 625 -1319 626 -1318
rect 656 -1319 657 -1318
rect 996 -1319 997 -1318
rect 156 -1321 157 -1320
rect 163 -1321 164 -1320
rect 177 -1321 178 -1320
rect 324 -1321 325 -1320
rect 415 -1321 416 -1320
rect 943 -1321 944 -1320
rect 142 -1323 143 -1322
rect 177 -1323 178 -1322
rect 191 -1323 192 -1322
rect 198 -1323 199 -1322
rect 208 -1323 209 -1322
rect 506 -1323 507 -1322
rect 534 -1323 535 -1322
rect 548 -1323 549 -1322
rect 590 -1323 591 -1322
rect 660 -1323 661 -1322
rect 667 -1323 668 -1322
rect 807 -1323 808 -1322
rect 835 -1323 836 -1322
rect 933 -1323 934 -1322
rect 100 -1325 101 -1324
rect 191 -1325 192 -1324
rect 212 -1325 213 -1324
rect 296 -1325 297 -1324
rect 313 -1325 314 -1324
rect 590 -1325 591 -1324
rect 625 -1325 626 -1324
rect 681 -1325 682 -1324
rect 688 -1325 689 -1324
rect 779 -1325 780 -1324
rect 100 -1327 101 -1326
rect 156 -1327 157 -1326
rect 233 -1327 234 -1326
rect 331 -1327 332 -1326
rect 429 -1327 430 -1326
rect 555 -1327 556 -1326
rect 674 -1327 675 -1326
rect 912 -1327 913 -1326
rect 142 -1329 143 -1328
rect 527 -1329 528 -1328
rect 562 -1329 563 -1328
rect 674 -1329 675 -1328
rect 702 -1329 703 -1328
rect 786 -1329 787 -1328
rect 233 -1331 234 -1330
rect 401 -1331 402 -1330
rect 432 -1331 433 -1330
rect 765 -1331 766 -1330
rect 240 -1333 241 -1332
rect 422 -1333 423 -1332
rect 436 -1333 437 -1332
rect 450 -1333 451 -1332
rect 460 -1333 461 -1332
rect 849 -1333 850 -1332
rect 247 -1335 248 -1334
rect 383 -1335 384 -1334
rect 394 -1335 395 -1334
rect 422 -1335 423 -1334
rect 443 -1335 444 -1334
rect 807 -1335 808 -1334
rect 205 -1337 206 -1336
rect 247 -1337 248 -1336
rect 254 -1337 255 -1336
rect 345 -1337 346 -1336
rect 366 -1337 367 -1336
rect 394 -1337 395 -1336
rect 443 -1337 444 -1336
rect 478 -1337 479 -1336
rect 481 -1337 482 -1336
rect 884 -1337 885 -1336
rect 303 -1339 304 -1338
rect 429 -1339 430 -1338
rect 450 -1339 451 -1338
rect 520 -1339 521 -1338
rect 527 -1339 528 -1338
rect 541 -1339 542 -1338
rect 716 -1339 717 -1338
rect 751 -1339 752 -1338
rect 765 -1339 766 -1338
rect 828 -1339 829 -1338
rect 877 -1339 878 -1338
rect 884 -1339 885 -1338
rect 338 -1341 339 -1340
rect 401 -1341 402 -1340
rect 478 -1341 479 -1340
rect 534 -1341 535 -1340
rect 639 -1341 640 -1340
rect 751 -1341 752 -1340
rect 814 -1341 815 -1340
rect 877 -1341 878 -1340
rect 338 -1343 339 -1342
rect 373 -1343 374 -1342
rect 383 -1343 384 -1342
rect 779 -1343 780 -1342
rect 814 -1343 815 -1342
rect 856 -1343 857 -1342
rect 268 -1345 269 -1344
rect 373 -1345 374 -1344
rect 485 -1345 486 -1344
rect 681 -1345 682 -1344
rect 737 -1345 738 -1344
rect 786 -1345 787 -1344
rect 800 -1345 801 -1344
rect 856 -1345 857 -1344
rect 268 -1347 269 -1346
rect 275 -1347 276 -1346
rect 513 -1347 514 -1346
rect 562 -1347 563 -1346
rect 639 -1347 640 -1346
rect 744 -1347 745 -1346
rect 758 -1347 759 -1346
rect 800 -1347 801 -1346
rect 828 -1347 829 -1346
rect 905 -1347 906 -1346
rect 79 -1349 80 -1348
rect 275 -1349 276 -1348
rect 485 -1349 486 -1348
rect 744 -1349 745 -1348
rect 758 -1349 759 -1348
rect 968 -1349 969 -1348
rect 79 -1351 80 -1350
rect 604 -1351 605 -1350
rect 695 -1351 696 -1350
rect 905 -1351 906 -1350
rect 513 -1353 514 -1352
rect 842 -1353 843 -1352
rect 520 -1355 521 -1354
rect 604 -1355 605 -1354
rect 737 -1355 738 -1354
rect 821 -1355 822 -1354
rect 842 -1355 843 -1354
rect 947 -1355 948 -1354
rect 821 -1357 822 -1356
rect 870 -1357 871 -1356
rect 870 -1359 871 -1358
rect 961 -1359 962 -1358
rect 2 -1370 3 -1369
rect 44 -1370 45 -1369
rect 58 -1370 59 -1369
rect 79 -1370 80 -1369
rect 86 -1370 87 -1369
rect 135 -1370 136 -1369
rect 156 -1370 157 -1369
rect 352 -1370 353 -1369
rect 376 -1370 377 -1369
rect 772 -1370 773 -1369
rect 856 -1370 857 -1369
rect 905 -1370 906 -1369
rect 908 -1370 909 -1369
rect 954 -1370 955 -1369
rect 971 -1370 972 -1369
rect 989 -1370 990 -1369
rect 9 -1372 10 -1371
rect 324 -1372 325 -1371
rect 394 -1372 395 -1371
rect 681 -1372 682 -1371
rect 712 -1372 713 -1371
rect 716 -1372 717 -1371
rect 765 -1372 766 -1371
rect 926 -1372 927 -1371
rect 947 -1372 948 -1371
rect 954 -1372 955 -1371
rect 9 -1374 10 -1373
rect 730 -1374 731 -1373
rect 765 -1374 766 -1373
rect 898 -1374 899 -1373
rect 912 -1374 913 -1373
rect 968 -1374 969 -1373
rect 37 -1376 38 -1375
rect 229 -1376 230 -1375
rect 240 -1376 241 -1375
rect 380 -1376 381 -1375
rect 397 -1376 398 -1375
rect 408 -1376 409 -1375
rect 450 -1376 451 -1375
rect 460 -1376 461 -1375
rect 467 -1376 468 -1375
rect 758 -1376 759 -1375
rect 856 -1376 857 -1375
rect 870 -1376 871 -1375
rect 891 -1376 892 -1375
rect 912 -1376 913 -1375
rect 37 -1378 38 -1377
rect 194 -1378 195 -1377
rect 205 -1378 206 -1377
rect 338 -1378 339 -1377
rect 348 -1378 349 -1377
rect 716 -1378 717 -1377
rect 744 -1378 745 -1377
rect 758 -1378 759 -1377
rect 800 -1378 801 -1377
rect 870 -1378 871 -1377
rect 51 -1380 52 -1379
rect 380 -1380 381 -1379
rect 401 -1380 402 -1379
rect 467 -1380 468 -1379
rect 478 -1380 479 -1379
rect 653 -1380 654 -1379
rect 681 -1380 682 -1379
rect 695 -1380 696 -1379
rect 702 -1380 703 -1379
rect 730 -1380 731 -1379
rect 800 -1380 801 -1379
rect 821 -1380 822 -1379
rect 849 -1380 850 -1379
rect 891 -1380 892 -1379
rect 51 -1382 52 -1381
rect 268 -1382 269 -1381
rect 296 -1382 297 -1381
rect 376 -1382 377 -1381
rect 401 -1382 402 -1381
rect 562 -1382 563 -1381
rect 576 -1382 577 -1381
rect 597 -1382 598 -1381
rect 604 -1382 605 -1381
rect 828 -1382 829 -1381
rect 842 -1382 843 -1381
rect 849 -1382 850 -1381
rect 863 -1382 864 -1381
rect 933 -1382 934 -1381
rect 65 -1384 66 -1383
rect 187 -1384 188 -1383
rect 191 -1384 192 -1383
rect 772 -1384 773 -1383
rect 807 -1384 808 -1383
rect 842 -1384 843 -1383
rect 863 -1384 864 -1383
rect 940 -1384 941 -1383
rect 33 -1386 34 -1385
rect 65 -1386 66 -1385
rect 72 -1386 73 -1385
rect 551 -1386 552 -1385
rect 555 -1386 556 -1385
rect 695 -1386 696 -1385
rect 702 -1386 703 -1385
rect 737 -1386 738 -1385
rect 72 -1388 73 -1387
rect 457 -1388 458 -1387
rect 464 -1388 465 -1387
rect 562 -1388 563 -1387
rect 590 -1388 591 -1387
rect 919 -1388 920 -1387
rect 79 -1390 80 -1389
rect 334 -1390 335 -1389
rect 338 -1390 339 -1389
rect 492 -1390 493 -1389
rect 516 -1390 517 -1389
rect 688 -1390 689 -1389
rect 723 -1390 724 -1389
rect 744 -1390 745 -1389
rect 89 -1392 90 -1391
rect 583 -1392 584 -1391
rect 593 -1392 594 -1391
rect 877 -1392 878 -1391
rect 93 -1394 94 -1393
rect 205 -1394 206 -1393
rect 226 -1394 227 -1393
rect 558 -1394 559 -1393
rect 569 -1394 570 -1393
rect 583 -1394 584 -1393
rect 604 -1394 605 -1393
rect 807 -1394 808 -1393
rect 877 -1394 878 -1393
rect 884 -1394 885 -1393
rect 93 -1396 94 -1395
rect 114 -1396 115 -1395
rect 124 -1396 125 -1395
rect 751 -1396 752 -1395
rect 835 -1396 836 -1395
rect 884 -1396 885 -1395
rect 100 -1398 101 -1397
rect 555 -1398 556 -1397
rect 667 -1398 668 -1397
rect 688 -1398 689 -1397
rect 709 -1398 710 -1397
rect 723 -1398 724 -1397
rect 751 -1398 752 -1397
rect 793 -1398 794 -1397
rect 835 -1398 836 -1397
rect 943 -1398 944 -1397
rect 23 -1400 24 -1399
rect 100 -1400 101 -1399
rect 128 -1400 129 -1399
rect 296 -1400 297 -1399
rect 310 -1400 311 -1399
rect 373 -1400 374 -1399
rect 453 -1400 454 -1399
rect 737 -1400 738 -1399
rect 779 -1400 780 -1399
rect 793 -1400 794 -1399
rect 943 -1400 944 -1399
rect 982 -1400 983 -1399
rect 23 -1402 24 -1401
rect 254 -1402 255 -1401
rect 261 -1402 262 -1401
rect 345 -1402 346 -1401
rect 373 -1402 374 -1401
rect 667 -1402 668 -1401
rect 121 -1404 122 -1403
rect 345 -1404 346 -1403
rect 478 -1404 479 -1403
rect 499 -1404 500 -1403
rect 527 -1404 528 -1403
rect 786 -1404 787 -1403
rect 121 -1406 122 -1405
rect 219 -1406 220 -1405
rect 233 -1406 234 -1405
rect 408 -1406 409 -1405
rect 471 -1406 472 -1405
rect 527 -1406 528 -1405
rect 530 -1406 531 -1405
rect 674 -1406 675 -1405
rect 786 -1406 787 -1405
rect 814 -1406 815 -1405
rect 135 -1408 136 -1407
rect 289 -1408 290 -1407
rect 310 -1408 311 -1407
rect 317 -1408 318 -1407
rect 331 -1408 332 -1407
rect 569 -1408 570 -1407
rect 646 -1408 647 -1407
rect 674 -1408 675 -1407
rect 149 -1410 150 -1409
rect 261 -1410 262 -1409
rect 289 -1410 290 -1409
rect 366 -1410 367 -1409
rect 390 -1410 391 -1409
rect 471 -1410 472 -1409
rect 481 -1410 482 -1409
rect 898 -1410 899 -1409
rect 107 -1412 108 -1411
rect 149 -1412 150 -1411
rect 159 -1412 160 -1411
rect 240 -1412 241 -1411
rect 247 -1412 248 -1411
rect 352 -1412 353 -1411
rect 366 -1412 367 -1411
rect 387 -1412 388 -1411
rect 485 -1412 486 -1411
rect 548 -1412 549 -1411
rect 632 -1412 633 -1411
rect 646 -1412 647 -1411
rect 660 -1412 661 -1411
rect 779 -1412 780 -1411
rect 30 -1414 31 -1413
rect 159 -1414 160 -1413
rect 166 -1414 167 -1413
rect 191 -1414 192 -1413
rect 219 -1414 220 -1413
rect 222 -1414 223 -1413
rect 233 -1414 234 -1413
rect 513 -1414 514 -1413
rect 537 -1414 538 -1413
rect 625 -1414 626 -1413
rect 632 -1414 633 -1413
rect 814 -1414 815 -1413
rect 107 -1416 108 -1415
rect 117 -1416 118 -1415
rect 170 -1416 171 -1415
rect 268 -1416 269 -1415
rect 317 -1416 318 -1415
rect 432 -1416 433 -1415
rect 492 -1416 493 -1415
rect 506 -1416 507 -1415
rect 513 -1416 514 -1415
rect 520 -1416 521 -1415
rect 534 -1416 535 -1415
rect 625 -1416 626 -1415
rect 639 -1416 640 -1415
rect 660 -1416 661 -1415
rect 16 -1418 17 -1417
rect 506 -1418 507 -1417
rect 541 -1418 542 -1417
rect 597 -1418 598 -1417
rect 16 -1420 17 -1419
rect 303 -1420 304 -1419
rect 464 -1420 465 -1419
rect 520 -1420 521 -1419
rect 541 -1420 542 -1419
rect 611 -1420 612 -1419
rect 163 -1422 164 -1421
rect 170 -1422 171 -1421
rect 177 -1422 178 -1421
rect 247 -1422 248 -1421
rect 254 -1422 255 -1421
rect 359 -1422 360 -1421
rect 488 -1422 489 -1421
rect 639 -1422 640 -1421
rect 128 -1424 129 -1423
rect 177 -1424 178 -1423
rect 184 -1424 185 -1423
rect 331 -1424 332 -1423
rect 499 -1424 500 -1423
rect 618 -1424 619 -1423
rect 212 -1426 213 -1425
rect 303 -1426 304 -1425
rect 509 -1426 510 -1425
rect 611 -1426 612 -1425
rect 282 -1428 283 -1427
rect 359 -1428 360 -1427
rect 579 -1428 580 -1427
rect 618 -1428 619 -1427
rect 282 -1430 283 -1429
rect 415 -1430 416 -1429
rect 579 -1430 580 -1429
rect 821 -1430 822 -1429
rect 415 -1432 416 -1431
rect 422 -1432 423 -1431
rect 422 -1434 423 -1433
rect 436 -1434 437 -1433
rect 436 -1436 437 -1435
rect 443 -1436 444 -1435
rect 142 -1438 143 -1437
rect 443 -1438 444 -1437
rect 9 -1449 10 -1448
rect 16 -1449 17 -1448
rect 23 -1449 24 -1448
rect 394 -1449 395 -1448
rect 432 -1449 433 -1448
rect 520 -1449 521 -1448
rect 548 -1449 549 -1448
rect 870 -1449 871 -1448
rect 940 -1449 941 -1448
rect 968 -1449 969 -1448
rect 16 -1451 17 -1450
rect 226 -1451 227 -1450
rect 282 -1451 283 -1450
rect 394 -1451 395 -1450
rect 457 -1451 458 -1450
rect 499 -1451 500 -1450
rect 502 -1451 503 -1450
rect 730 -1451 731 -1450
rect 961 -1451 962 -1450
rect 982 -1451 983 -1450
rect 23 -1453 24 -1452
rect 37 -1453 38 -1452
rect 44 -1453 45 -1452
rect 107 -1453 108 -1452
rect 114 -1453 115 -1452
rect 282 -1453 283 -1452
rect 285 -1453 286 -1452
rect 513 -1453 514 -1452
rect 555 -1453 556 -1452
rect 884 -1453 885 -1452
rect 982 -1453 983 -1452
rect 989 -1453 990 -1452
rect 51 -1455 52 -1454
rect 362 -1455 363 -1454
rect 373 -1455 374 -1454
rect 415 -1455 416 -1454
rect 432 -1455 433 -1454
rect 499 -1455 500 -1454
rect 506 -1455 507 -1454
rect 863 -1455 864 -1454
rect 51 -1457 52 -1456
rect 551 -1457 552 -1456
rect 558 -1457 559 -1456
rect 926 -1457 927 -1456
rect 79 -1459 80 -1458
rect 590 -1459 591 -1458
rect 604 -1459 605 -1458
rect 779 -1459 780 -1458
rect 79 -1461 80 -1460
rect 222 -1461 223 -1460
rect 303 -1461 304 -1460
rect 390 -1461 391 -1460
rect 397 -1461 398 -1460
rect 779 -1461 780 -1460
rect 93 -1463 94 -1462
rect 131 -1463 132 -1462
rect 142 -1463 143 -1462
rect 331 -1463 332 -1462
rect 338 -1463 339 -1462
rect 429 -1463 430 -1462
rect 460 -1463 461 -1462
rect 898 -1463 899 -1462
rect 93 -1465 94 -1464
rect 317 -1465 318 -1464
rect 345 -1465 346 -1464
rect 548 -1465 549 -1464
rect 576 -1465 577 -1464
rect 611 -1465 612 -1464
rect 632 -1465 633 -1464
rect 905 -1465 906 -1464
rect 100 -1467 101 -1466
rect 317 -1467 318 -1466
rect 352 -1467 353 -1466
rect 366 -1467 367 -1466
rect 376 -1467 377 -1466
rect 380 -1467 381 -1466
rect 415 -1467 416 -1466
rect 422 -1467 423 -1466
rect 467 -1467 468 -1466
rect 828 -1467 829 -1466
rect 887 -1467 888 -1466
rect 898 -1467 899 -1466
rect 905 -1467 906 -1466
rect 912 -1467 913 -1466
rect 100 -1469 101 -1468
rect 411 -1469 412 -1468
rect 422 -1469 423 -1468
rect 478 -1469 479 -1468
rect 485 -1469 486 -1468
rect 607 -1469 608 -1468
rect 611 -1469 612 -1468
rect 660 -1469 661 -1468
rect 688 -1469 689 -1468
rect 709 -1469 710 -1468
rect 712 -1469 713 -1468
rect 814 -1469 815 -1468
rect 912 -1469 913 -1468
rect 933 -1469 934 -1468
rect 65 -1471 66 -1470
rect 660 -1471 661 -1470
rect 688 -1471 689 -1470
rect 793 -1471 794 -1470
rect 65 -1473 66 -1472
rect 72 -1473 73 -1472
rect 117 -1473 118 -1472
rect 149 -1473 150 -1472
rect 156 -1473 157 -1472
rect 737 -1473 738 -1472
rect 793 -1473 794 -1472
rect 842 -1473 843 -1472
rect 86 -1475 87 -1474
rect 156 -1475 157 -1474
rect 159 -1475 160 -1474
rect 625 -1475 626 -1474
rect 632 -1475 633 -1474
rect 635 -1475 636 -1474
rect 653 -1475 654 -1474
rect 891 -1475 892 -1474
rect 86 -1477 87 -1476
rect 194 -1477 195 -1476
rect 201 -1477 202 -1476
rect 268 -1477 269 -1476
rect 352 -1477 353 -1476
rect 464 -1477 465 -1476
rect 467 -1477 468 -1476
rect 695 -1477 696 -1476
rect 730 -1477 731 -1476
rect 744 -1477 745 -1476
rect 821 -1477 822 -1476
rect 891 -1477 892 -1476
rect 107 -1479 108 -1478
rect 464 -1479 465 -1478
rect 471 -1479 472 -1478
rect 555 -1479 556 -1478
rect 590 -1479 591 -1478
rect 681 -1479 682 -1478
rect 695 -1479 696 -1478
rect 723 -1479 724 -1478
rect 737 -1479 738 -1478
rect 950 -1479 951 -1478
rect 58 -1481 59 -1480
rect 471 -1481 472 -1480
rect 478 -1481 479 -1480
rect 772 -1481 773 -1480
rect 842 -1481 843 -1480
rect 919 -1481 920 -1480
rect 58 -1483 59 -1482
rect 233 -1483 234 -1482
rect 240 -1483 241 -1482
rect 345 -1483 346 -1482
rect 355 -1483 356 -1482
rect 450 -1483 451 -1482
rect 485 -1483 486 -1482
rect 541 -1483 542 -1482
rect 597 -1483 598 -1482
rect 604 -1483 605 -1482
rect 625 -1483 626 -1482
rect 656 -1483 657 -1482
rect 681 -1483 682 -1482
rect 702 -1483 703 -1482
rect 723 -1483 724 -1482
rect 751 -1483 752 -1482
rect 765 -1483 766 -1482
rect 772 -1483 773 -1482
rect 919 -1483 920 -1482
rect 954 -1483 955 -1482
rect 121 -1485 122 -1484
rect 303 -1485 304 -1484
rect 324 -1485 325 -1484
rect 541 -1485 542 -1484
rect 597 -1485 598 -1484
rect 639 -1485 640 -1484
rect 653 -1485 654 -1484
rect 716 -1485 717 -1484
rect 744 -1485 745 -1484
rect 758 -1485 759 -1484
rect 933 -1485 934 -1484
rect 954 -1485 955 -1484
rect 128 -1487 129 -1486
rect 506 -1487 507 -1486
rect 509 -1487 510 -1486
rect 674 -1487 675 -1486
rect 702 -1487 703 -1486
rect 835 -1487 836 -1486
rect 135 -1489 136 -1488
rect 380 -1489 381 -1488
rect 443 -1489 444 -1488
rect 716 -1489 717 -1488
rect 751 -1489 752 -1488
rect 786 -1489 787 -1488
rect 835 -1489 836 -1488
rect 849 -1489 850 -1488
rect 40 -1491 41 -1490
rect 849 -1491 850 -1490
rect 142 -1493 143 -1492
rect 180 -1493 181 -1492
rect 184 -1493 185 -1492
rect 331 -1493 332 -1492
rect 366 -1493 367 -1492
rect 408 -1493 409 -1492
rect 443 -1493 444 -1492
rect 520 -1493 521 -1492
rect 537 -1493 538 -1492
rect 821 -1493 822 -1492
rect 149 -1495 150 -1494
rect 254 -1495 255 -1494
rect 261 -1495 262 -1494
rect 324 -1495 325 -1494
rect 369 -1495 370 -1494
rect 765 -1495 766 -1494
rect 786 -1495 787 -1494
rect 807 -1495 808 -1494
rect 163 -1497 164 -1496
rect 170 -1497 171 -1496
rect 173 -1497 174 -1496
rect 359 -1497 360 -1496
rect 492 -1497 493 -1496
rect 513 -1497 514 -1496
rect 537 -1497 538 -1496
rect 814 -1497 815 -1496
rect 30 -1499 31 -1498
rect 163 -1499 164 -1498
rect 184 -1499 185 -1498
rect 387 -1499 388 -1498
rect 492 -1499 493 -1498
rect 527 -1499 528 -1498
rect 618 -1499 619 -1498
rect 639 -1499 640 -1498
rect 667 -1499 668 -1498
rect 674 -1499 675 -1498
rect 807 -1499 808 -1498
rect 877 -1499 878 -1498
rect 30 -1501 31 -1500
rect 289 -1501 290 -1500
rect 359 -1501 360 -1500
rect 618 -1501 619 -1500
rect 646 -1501 647 -1500
rect 667 -1501 668 -1500
rect 152 -1503 153 -1502
rect 646 -1503 647 -1502
rect 187 -1505 188 -1504
rect 247 -1505 248 -1504
rect 261 -1505 262 -1504
rect 593 -1505 594 -1504
rect 187 -1507 188 -1506
rect 569 -1507 570 -1506
rect 191 -1509 192 -1508
rect 254 -1509 255 -1508
rect 289 -1509 290 -1508
rect 446 -1509 447 -1508
rect 562 -1509 563 -1508
rect 569 -1509 570 -1508
rect 191 -1511 192 -1510
rect 306 -1511 307 -1510
rect 401 -1511 402 -1510
rect 527 -1511 528 -1510
rect 562 -1511 563 -1510
rect 583 -1511 584 -1510
rect 205 -1513 206 -1512
rect 247 -1513 248 -1512
rect 401 -1513 402 -1512
rect 436 -1513 437 -1512
rect 583 -1513 584 -1512
rect 884 -1513 885 -1512
rect 166 -1515 167 -1514
rect 436 -1515 437 -1514
rect 177 -1517 178 -1516
rect 205 -1517 206 -1516
rect 219 -1517 220 -1516
rect 226 -1517 227 -1516
rect 233 -1517 234 -1516
rect 453 -1517 454 -1516
rect 177 -1519 178 -1518
rect 268 -1519 269 -1518
rect 219 -1521 220 -1520
rect 296 -1521 297 -1520
rect 240 -1523 241 -1522
rect 429 -1523 430 -1522
rect 275 -1525 276 -1524
rect 296 -1525 297 -1524
rect 2 -1527 3 -1526
rect 275 -1527 276 -1526
rect 23 -1538 24 -1537
rect 40 -1538 41 -1537
rect 44 -1538 45 -1537
rect 163 -1538 164 -1537
rect 166 -1538 167 -1537
rect 289 -1538 290 -1537
rect 306 -1538 307 -1537
rect 373 -1538 374 -1537
rect 432 -1538 433 -1537
rect 485 -1538 486 -1537
rect 509 -1538 510 -1537
rect 842 -1538 843 -1537
rect 849 -1538 850 -1537
rect 926 -1538 927 -1537
rect 947 -1538 948 -1537
rect 968 -1538 969 -1537
rect 982 -1538 983 -1537
rect 989 -1538 990 -1537
rect 30 -1540 31 -1539
rect 292 -1540 293 -1539
rect 345 -1540 346 -1539
rect 366 -1540 367 -1539
rect 373 -1540 374 -1539
rect 401 -1540 402 -1539
rect 436 -1540 437 -1539
rect 852 -1540 853 -1539
rect 884 -1540 885 -1539
rect 940 -1540 941 -1539
rect 954 -1540 955 -1539
rect 971 -1540 972 -1539
rect 16 -1542 17 -1541
rect 30 -1542 31 -1541
rect 37 -1542 38 -1541
rect 275 -1542 276 -1541
rect 282 -1542 283 -1541
rect 285 -1542 286 -1541
rect 352 -1542 353 -1541
rect 464 -1542 465 -1541
rect 478 -1542 479 -1541
rect 590 -1542 591 -1541
rect 604 -1542 605 -1541
rect 870 -1542 871 -1541
rect 898 -1542 899 -1541
rect 915 -1542 916 -1541
rect 940 -1542 941 -1541
rect 975 -1542 976 -1541
rect 16 -1544 17 -1543
rect 348 -1544 349 -1543
rect 352 -1544 353 -1543
rect 380 -1544 381 -1543
rect 401 -1544 402 -1543
rect 646 -1544 647 -1543
rect 705 -1544 706 -1543
rect 772 -1544 773 -1543
rect 800 -1544 801 -1543
rect 849 -1544 850 -1543
rect 898 -1544 899 -1543
rect 912 -1544 913 -1543
rect 37 -1546 38 -1545
rect 96 -1546 97 -1545
rect 100 -1546 101 -1545
rect 138 -1546 139 -1545
rect 149 -1546 150 -1545
rect 457 -1546 458 -1545
rect 478 -1546 479 -1545
rect 492 -1546 493 -1545
rect 520 -1546 521 -1545
rect 523 -1546 524 -1545
rect 534 -1546 535 -1545
rect 730 -1546 731 -1545
rect 733 -1546 734 -1545
rect 807 -1546 808 -1545
rect 814 -1546 815 -1545
rect 842 -1546 843 -1545
rect 44 -1548 45 -1547
rect 128 -1548 129 -1547
rect 135 -1548 136 -1547
rect 359 -1548 360 -1547
rect 436 -1548 437 -1547
rect 481 -1548 482 -1547
rect 485 -1548 486 -1547
rect 527 -1548 528 -1547
rect 586 -1548 587 -1547
rect 716 -1548 717 -1547
rect 814 -1548 815 -1547
rect 905 -1548 906 -1547
rect 9 -1550 10 -1549
rect 481 -1550 482 -1549
rect 492 -1550 493 -1549
rect 632 -1550 633 -1549
rect 646 -1550 647 -1549
rect 695 -1550 696 -1549
rect 716 -1550 717 -1549
rect 751 -1550 752 -1549
rect 65 -1552 66 -1551
rect 408 -1552 409 -1551
rect 446 -1552 447 -1551
rect 709 -1552 710 -1551
rect 751 -1552 752 -1551
rect 891 -1552 892 -1551
rect 65 -1554 66 -1553
rect 184 -1554 185 -1553
rect 194 -1554 195 -1553
rect 597 -1554 598 -1553
rect 604 -1554 605 -1553
rect 653 -1554 654 -1553
rect 709 -1554 710 -1553
rect 828 -1554 829 -1553
rect 86 -1556 87 -1555
rect 366 -1556 367 -1555
rect 408 -1556 409 -1555
rect 471 -1556 472 -1555
rect 520 -1556 521 -1555
rect 576 -1556 577 -1555
rect 590 -1556 591 -1555
rect 688 -1556 689 -1555
rect 86 -1558 87 -1557
rect 110 -1558 111 -1557
rect 114 -1558 115 -1557
rect 499 -1558 500 -1557
rect 555 -1558 556 -1557
rect 597 -1558 598 -1557
rect 618 -1558 619 -1557
rect 954 -1558 955 -1557
rect 93 -1560 94 -1559
rect 443 -1560 444 -1559
rect 450 -1560 451 -1559
rect 737 -1560 738 -1559
rect 100 -1562 101 -1561
rect 303 -1562 304 -1561
rect 341 -1562 342 -1561
rect 828 -1562 829 -1561
rect 107 -1564 108 -1563
rect 345 -1564 346 -1563
rect 369 -1564 370 -1563
rect 443 -1564 444 -1563
rect 453 -1564 454 -1563
rect 744 -1564 745 -1563
rect 58 -1566 59 -1565
rect 453 -1566 454 -1565
rect 457 -1566 458 -1565
rect 513 -1566 514 -1565
rect 530 -1566 531 -1565
rect 555 -1566 556 -1565
rect 632 -1566 633 -1565
rect 660 -1566 661 -1565
rect 688 -1566 689 -1565
rect 702 -1566 703 -1565
rect 744 -1566 745 -1565
rect 835 -1566 836 -1565
rect 58 -1568 59 -1567
rect 695 -1568 696 -1567
rect 702 -1568 703 -1567
rect 919 -1568 920 -1567
rect 128 -1570 129 -1569
rect 331 -1570 332 -1569
rect 411 -1570 412 -1569
rect 653 -1570 654 -1569
rect 660 -1570 661 -1569
rect 681 -1570 682 -1569
rect 880 -1570 881 -1569
rect 919 -1570 920 -1569
rect 135 -1572 136 -1571
rect 205 -1572 206 -1571
rect 212 -1572 213 -1571
rect 247 -1572 248 -1571
rect 261 -1572 262 -1571
rect 275 -1572 276 -1571
rect 282 -1572 283 -1571
rect 324 -1572 325 -1571
rect 331 -1572 332 -1571
rect 467 -1572 468 -1571
rect 513 -1572 514 -1571
rect 548 -1572 549 -1571
rect 75 -1574 76 -1573
rect 261 -1574 262 -1573
rect 289 -1574 290 -1573
rect 471 -1574 472 -1573
rect 534 -1574 535 -1573
rect 681 -1574 682 -1573
rect 149 -1576 150 -1575
rect 359 -1576 360 -1575
rect 429 -1576 430 -1575
rect 499 -1576 500 -1575
rect 548 -1576 549 -1575
rect 562 -1576 563 -1575
rect 156 -1578 157 -1577
rect 254 -1578 255 -1577
rect 303 -1578 304 -1577
rect 317 -1578 318 -1577
rect 324 -1578 325 -1577
rect 541 -1578 542 -1577
rect 562 -1578 563 -1577
rect 765 -1578 766 -1577
rect 156 -1580 157 -1579
rect 793 -1580 794 -1579
rect 159 -1582 160 -1581
rect 254 -1582 255 -1581
rect 317 -1582 318 -1581
rect 394 -1582 395 -1581
rect 429 -1582 430 -1581
rect 565 -1582 566 -1581
rect 765 -1582 766 -1581
rect 821 -1582 822 -1581
rect 72 -1584 73 -1583
rect 394 -1584 395 -1583
rect 793 -1584 794 -1583
rect 856 -1584 857 -1583
rect 72 -1586 73 -1585
rect 240 -1586 241 -1585
rect 247 -1586 248 -1585
rect 296 -1586 297 -1585
rect 362 -1586 363 -1585
rect 856 -1586 857 -1585
rect 177 -1588 178 -1587
rect 611 -1588 612 -1587
rect 177 -1590 178 -1589
rect 674 -1590 675 -1589
rect 198 -1592 199 -1591
rect 268 -1592 269 -1591
rect 296 -1592 297 -1591
rect 338 -1592 339 -1591
rect 362 -1592 363 -1591
rect 422 -1592 423 -1591
rect 569 -1592 570 -1591
rect 611 -1592 612 -1591
rect 674 -1592 675 -1591
rect 779 -1592 780 -1591
rect 173 -1594 174 -1593
rect 268 -1594 269 -1593
rect 338 -1594 339 -1593
rect 625 -1594 626 -1593
rect 201 -1596 202 -1595
rect 219 -1596 220 -1595
rect 240 -1596 241 -1595
rect 537 -1596 538 -1595
rect 569 -1596 570 -1595
rect 639 -1596 640 -1595
rect 215 -1598 216 -1597
rect 226 -1598 227 -1597
rect 387 -1598 388 -1597
rect 541 -1598 542 -1597
rect 639 -1598 640 -1597
rect 667 -1598 668 -1597
rect 226 -1600 227 -1599
rect 310 -1600 311 -1599
rect 506 -1600 507 -1599
rect 625 -1600 626 -1599
rect 667 -1600 668 -1599
rect 800 -1600 801 -1599
rect 233 -1602 234 -1601
rect 310 -1602 311 -1601
rect 506 -1602 507 -1601
rect 583 -1602 584 -1601
rect 51 -1604 52 -1603
rect 233 -1604 234 -1603
rect 523 -1604 524 -1603
rect 576 -1604 577 -1603
rect 51 -1606 52 -1605
rect 79 -1606 80 -1605
rect 537 -1606 538 -1605
rect 786 -1606 787 -1605
rect 26 -1608 27 -1607
rect 786 -1608 787 -1607
rect 79 -1610 80 -1609
rect 121 -1610 122 -1609
rect 121 -1612 122 -1611
rect 758 -1612 759 -1611
rect 9 -1623 10 -1622
rect 23 -1623 24 -1622
rect 30 -1623 31 -1622
rect 121 -1623 122 -1622
rect 124 -1623 125 -1622
rect 681 -1623 682 -1622
rect 695 -1623 696 -1622
rect 940 -1623 941 -1622
rect 943 -1623 944 -1622
rect 961 -1623 962 -1622
rect 971 -1623 972 -1622
rect 975 -1623 976 -1622
rect 9 -1625 10 -1624
rect 240 -1625 241 -1624
rect 247 -1625 248 -1624
rect 250 -1625 251 -1624
rect 289 -1625 290 -1624
rect 387 -1625 388 -1624
rect 390 -1625 391 -1624
rect 737 -1625 738 -1624
rect 793 -1625 794 -1624
rect 849 -1625 850 -1624
rect 877 -1625 878 -1624
rect 898 -1625 899 -1624
rect 912 -1625 913 -1624
rect 919 -1625 920 -1624
rect 975 -1625 976 -1624
rect 982 -1625 983 -1624
rect 16 -1627 17 -1626
rect 187 -1627 188 -1626
rect 240 -1627 241 -1626
rect 296 -1627 297 -1626
rect 299 -1627 300 -1626
rect 653 -1627 654 -1626
rect 660 -1627 661 -1626
rect 667 -1627 668 -1626
rect 712 -1627 713 -1626
rect 765 -1627 766 -1626
rect 835 -1627 836 -1626
rect 856 -1627 857 -1626
rect 894 -1627 895 -1626
rect 926 -1627 927 -1626
rect 16 -1629 17 -1628
rect 61 -1629 62 -1628
rect 93 -1629 94 -1628
rect 625 -1629 626 -1628
rect 639 -1629 640 -1628
rect 863 -1629 864 -1628
rect 926 -1629 927 -1628
rect 947 -1629 948 -1628
rect 23 -1631 24 -1630
rect 96 -1631 97 -1630
rect 100 -1631 101 -1630
rect 184 -1631 185 -1630
rect 247 -1631 248 -1630
rect 310 -1631 311 -1630
rect 341 -1631 342 -1630
rect 705 -1631 706 -1630
rect 723 -1631 724 -1630
rect 730 -1631 731 -1630
rect 842 -1631 843 -1630
rect 887 -1631 888 -1630
rect 30 -1633 31 -1632
rect 296 -1633 297 -1632
rect 303 -1633 304 -1632
rect 338 -1633 339 -1632
rect 341 -1633 342 -1632
rect 632 -1633 633 -1632
rect 660 -1633 661 -1632
rect 744 -1633 745 -1632
rect 828 -1633 829 -1632
rect 842 -1633 843 -1632
rect 37 -1635 38 -1634
rect 58 -1635 59 -1634
rect 93 -1635 94 -1634
rect 117 -1635 118 -1634
rect 163 -1635 164 -1634
rect 625 -1635 626 -1634
rect 667 -1635 668 -1634
rect 751 -1635 752 -1634
rect 37 -1637 38 -1636
rect 422 -1637 423 -1636
rect 439 -1637 440 -1636
rect 618 -1637 619 -1636
rect 716 -1637 717 -1636
rect 744 -1637 745 -1636
rect 44 -1639 45 -1638
rect 205 -1639 206 -1638
rect 250 -1639 251 -1638
rect 310 -1639 311 -1638
rect 331 -1639 332 -1638
rect 632 -1639 633 -1638
rect 44 -1641 45 -1640
rect 51 -1641 52 -1640
rect 58 -1641 59 -1640
rect 86 -1641 87 -1640
rect 107 -1641 108 -1640
rect 226 -1641 227 -1640
rect 303 -1641 304 -1640
rect 397 -1641 398 -1640
rect 404 -1641 405 -1640
rect 765 -1641 766 -1640
rect 51 -1643 52 -1642
rect 212 -1643 213 -1642
rect 226 -1643 227 -1642
rect 345 -1643 346 -1642
rect 348 -1643 349 -1642
rect 373 -1643 374 -1642
rect 383 -1643 384 -1642
rect 730 -1643 731 -1642
rect 86 -1645 87 -1644
rect 103 -1645 104 -1644
rect 110 -1645 111 -1644
rect 324 -1645 325 -1644
rect 359 -1645 360 -1644
rect 366 -1645 367 -1644
rect 387 -1645 388 -1644
rect 429 -1645 430 -1644
rect 450 -1645 451 -1644
rect 723 -1645 724 -1644
rect 128 -1647 129 -1646
rect 212 -1647 213 -1646
rect 282 -1647 283 -1646
rect 324 -1647 325 -1646
rect 352 -1647 353 -1646
rect 366 -1647 367 -1646
rect 429 -1647 430 -1646
rect 457 -1647 458 -1646
rect 464 -1647 465 -1646
rect 702 -1647 703 -1646
rect 65 -1649 66 -1648
rect 352 -1649 353 -1648
rect 401 -1649 402 -1648
rect 457 -1649 458 -1648
rect 464 -1649 465 -1648
rect 681 -1649 682 -1648
rect 65 -1651 66 -1650
rect 79 -1651 80 -1650
rect 128 -1651 129 -1650
rect 180 -1651 181 -1650
rect 282 -1651 283 -1650
rect 408 -1651 409 -1650
rect 450 -1651 451 -1650
rect 779 -1651 780 -1650
rect 135 -1653 136 -1652
rect 205 -1653 206 -1652
rect 317 -1653 318 -1652
rect 345 -1653 346 -1652
rect 401 -1653 402 -1652
rect 772 -1653 773 -1652
rect 135 -1655 136 -1654
rect 149 -1655 150 -1654
rect 163 -1655 164 -1654
rect 191 -1655 192 -1654
rect 219 -1655 220 -1654
rect 317 -1655 318 -1654
rect 331 -1655 332 -1654
rect 702 -1655 703 -1654
rect 72 -1657 73 -1656
rect 191 -1657 192 -1656
rect 408 -1657 409 -1656
rect 415 -1657 416 -1656
rect 453 -1657 454 -1656
rect 709 -1657 710 -1656
rect 145 -1659 146 -1658
rect 422 -1659 423 -1658
rect 471 -1659 472 -1658
rect 653 -1659 654 -1658
rect 149 -1661 150 -1660
rect 758 -1661 759 -1660
rect 166 -1663 167 -1662
rect 268 -1663 269 -1662
rect 471 -1663 472 -1662
rect 513 -1663 514 -1662
rect 527 -1663 528 -1662
rect 674 -1663 675 -1662
rect 170 -1665 171 -1664
rect 177 -1665 178 -1664
rect 198 -1665 199 -1664
rect 415 -1665 416 -1664
rect 478 -1665 479 -1664
rect 492 -1665 493 -1664
rect 495 -1665 496 -1664
rect 688 -1665 689 -1664
rect 173 -1667 174 -1666
rect 219 -1667 220 -1666
rect 254 -1667 255 -1666
rect 513 -1667 514 -1666
rect 527 -1667 528 -1666
rect 548 -1667 549 -1666
rect 555 -1667 556 -1666
rect 716 -1667 717 -1666
rect 173 -1669 174 -1668
rect 184 -1669 185 -1668
rect 198 -1669 199 -1668
rect 208 -1669 209 -1668
rect 254 -1669 255 -1668
rect 261 -1669 262 -1668
rect 268 -1669 269 -1668
rect 425 -1669 426 -1668
rect 488 -1669 489 -1668
rect 954 -1669 955 -1668
rect 79 -1671 80 -1670
rect 208 -1671 209 -1670
rect 261 -1671 262 -1670
rect 275 -1671 276 -1670
rect 492 -1671 493 -1670
rect 499 -1671 500 -1670
rect 506 -1671 507 -1670
rect 548 -1671 549 -1670
rect 555 -1671 556 -1670
rect 576 -1671 577 -1670
rect 586 -1671 587 -1670
rect 695 -1671 696 -1670
rect 233 -1673 234 -1672
rect 275 -1673 276 -1672
rect 499 -1673 500 -1672
rect 520 -1673 521 -1672
rect 534 -1673 535 -1672
rect 800 -1673 801 -1672
rect 156 -1675 157 -1674
rect 534 -1675 535 -1674
rect 537 -1675 538 -1674
rect 828 -1675 829 -1674
rect 142 -1677 143 -1676
rect 156 -1677 157 -1676
rect 509 -1677 510 -1676
rect 870 -1677 871 -1676
rect 142 -1679 143 -1678
rect 576 -1679 577 -1678
rect 590 -1679 591 -1678
rect 758 -1679 759 -1678
rect 786 -1679 787 -1678
rect 800 -1679 801 -1678
rect 814 -1679 815 -1678
rect 870 -1679 871 -1678
rect 485 -1681 486 -1680
rect 786 -1681 787 -1680
rect 541 -1683 542 -1682
rect 814 -1683 815 -1682
rect 520 -1685 521 -1684
rect 541 -1685 542 -1684
rect 544 -1685 545 -1684
rect 646 -1685 647 -1684
rect 562 -1687 563 -1686
rect 604 -1687 605 -1686
rect 611 -1687 612 -1686
rect 674 -1687 675 -1686
rect 152 -1689 153 -1688
rect 611 -1689 612 -1688
rect 443 -1691 444 -1690
rect 604 -1691 605 -1690
rect 436 -1693 437 -1692
rect 443 -1693 444 -1692
rect 481 -1693 482 -1692
rect 562 -1693 563 -1692
rect 565 -1693 566 -1692
rect 639 -1693 640 -1692
rect 380 -1695 381 -1694
rect 436 -1695 437 -1694
rect 569 -1695 570 -1694
rect 821 -1695 822 -1694
rect 569 -1697 570 -1696
rect 688 -1697 689 -1696
rect 583 -1699 584 -1698
rect 646 -1699 647 -1698
rect 572 -1701 573 -1700
rect 583 -1701 584 -1700
rect 590 -1701 591 -1700
rect 733 -1701 734 -1700
rect 597 -1703 598 -1702
rect 751 -1703 752 -1702
rect 394 -1705 395 -1704
rect 597 -1705 598 -1704
rect 16 -1716 17 -1715
rect 58 -1716 59 -1715
rect 72 -1716 73 -1715
rect 75 -1716 76 -1715
rect 79 -1716 80 -1715
rect 495 -1716 496 -1715
rect 506 -1716 507 -1715
rect 548 -1716 549 -1715
rect 572 -1716 573 -1715
rect 863 -1716 864 -1715
rect 905 -1716 906 -1715
rect 912 -1716 913 -1715
rect 926 -1716 927 -1715
rect 940 -1716 941 -1715
rect 961 -1716 962 -1715
rect 978 -1716 979 -1715
rect 16 -1718 17 -1717
rect 345 -1718 346 -1717
rect 355 -1718 356 -1717
rect 772 -1718 773 -1717
rect 37 -1720 38 -1719
rect 394 -1720 395 -1719
rect 397 -1720 398 -1719
rect 429 -1720 430 -1719
rect 436 -1720 437 -1719
rect 688 -1720 689 -1719
rect 709 -1720 710 -1719
rect 758 -1720 759 -1719
rect 37 -1722 38 -1721
rect 509 -1722 510 -1721
rect 523 -1722 524 -1721
rect 702 -1722 703 -1721
rect 51 -1724 52 -1723
rect 341 -1724 342 -1723
rect 376 -1724 377 -1723
rect 730 -1724 731 -1723
rect 58 -1726 59 -1725
rect 65 -1726 66 -1725
rect 93 -1726 94 -1725
rect 387 -1726 388 -1725
rect 439 -1726 440 -1725
rect 786 -1726 787 -1725
rect 9 -1728 10 -1727
rect 65 -1728 66 -1727
rect 103 -1728 104 -1727
rect 457 -1728 458 -1727
rect 467 -1728 468 -1727
rect 814 -1728 815 -1727
rect 9 -1730 10 -1729
rect 373 -1730 374 -1729
rect 387 -1730 388 -1729
rect 408 -1730 409 -1729
rect 450 -1730 451 -1729
rect 821 -1730 822 -1729
rect 86 -1732 87 -1731
rect 103 -1732 104 -1731
rect 117 -1732 118 -1731
rect 534 -1732 535 -1731
rect 548 -1732 549 -1731
rect 555 -1732 556 -1731
rect 642 -1732 643 -1731
rect 870 -1732 871 -1731
rect 23 -1734 24 -1733
rect 117 -1734 118 -1733
rect 121 -1734 122 -1733
rect 149 -1734 150 -1733
rect 159 -1734 160 -1733
rect 737 -1734 738 -1733
rect 23 -1736 24 -1735
rect 187 -1736 188 -1735
rect 191 -1736 192 -1735
rect 205 -1736 206 -1735
rect 222 -1736 223 -1735
rect 383 -1736 384 -1735
rect 450 -1736 451 -1735
rect 478 -1736 479 -1735
rect 485 -1736 486 -1735
rect 492 -1736 493 -1735
rect 534 -1736 535 -1735
rect 590 -1736 591 -1735
rect 667 -1736 668 -1735
rect 758 -1736 759 -1735
rect 82 -1738 83 -1737
rect 86 -1738 87 -1737
rect 124 -1738 125 -1737
rect 569 -1738 570 -1737
rect 702 -1738 703 -1737
rect 765 -1738 766 -1737
rect 128 -1740 129 -1739
rect 590 -1740 591 -1739
rect 730 -1740 731 -1739
rect 800 -1740 801 -1739
rect 142 -1742 143 -1741
rect 660 -1742 661 -1741
rect 737 -1742 738 -1741
rect 828 -1742 829 -1741
rect 163 -1744 164 -1743
rect 170 -1744 171 -1743
rect 173 -1744 174 -1743
rect 261 -1744 262 -1743
rect 268 -1744 269 -1743
rect 334 -1744 335 -1743
rect 471 -1744 472 -1743
rect 485 -1744 486 -1743
rect 488 -1744 489 -1743
rect 667 -1744 668 -1743
rect 166 -1746 167 -1745
rect 422 -1746 423 -1745
rect 474 -1746 475 -1745
rect 716 -1746 717 -1745
rect 170 -1748 171 -1747
rect 408 -1748 409 -1747
rect 422 -1748 423 -1747
rect 887 -1748 888 -1747
rect 191 -1750 192 -1749
rect 247 -1750 248 -1749
rect 261 -1750 262 -1749
rect 303 -1750 304 -1749
rect 310 -1750 311 -1749
rect 376 -1750 377 -1749
rect 478 -1750 479 -1749
rect 527 -1750 528 -1749
rect 555 -1750 556 -1749
rect 611 -1750 612 -1749
rect 660 -1750 661 -1749
rect 723 -1750 724 -1749
rect 107 -1752 108 -1751
rect 303 -1752 304 -1751
rect 324 -1752 325 -1751
rect 345 -1752 346 -1751
rect 527 -1752 528 -1751
rect 576 -1752 577 -1751
rect 716 -1752 717 -1751
rect 842 -1752 843 -1751
rect 107 -1754 108 -1753
rect 135 -1754 136 -1753
rect 156 -1754 157 -1753
rect 247 -1754 248 -1753
rect 271 -1754 272 -1753
rect 835 -1754 836 -1753
rect 30 -1756 31 -1755
rect 156 -1756 157 -1755
rect 219 -1756 220 -1755
rect 310 -1756 311 -1755
rect 324 -1756 325 -1755
rect 338 -1756 339 -1755
rect 576 -1756 577 -1755
rect 625 -1756 626 -1755
rect 723 -1756 724 -1755
rect 779 -1756 780 -1755
rect 30 -1758 31 -1757
rect 51 -1758 52 -1757
rect 219 -1758 220 -1757
rect 429 -1758 430 -1757
rect 625 -1758 626 -1757
rect 695 -1758 696 -1757
rect 226 -1760 227 -1759
rect 541 -1760 542 -1759
rect 695 -1760 696 -1759
rect 744 -1760 745 -1759
rect 114 -1762 115 -1761
rect 226 -1762 227 -1761
rect 233 -1762 234 -1761
rect 415 -1762 416 -1761
rect 541 -1762 542 -1761
rect 597 -1762 598 -1761
rect 639 -1762 640 -1761
rect 744 -1762 745 -1761
rect 198 -1764 199 -1763
rect 233 -1764 234 -1763
rect 236 -1764 237 -1763
rect 611 -1764 612 -1763
rect 198 -1766 199 -1765
rect 320 -1766 321 -1765
rect 338 -1766 339 -1765
rect 366 -1766 367 -1765
rect 415 -1766 416 -1765
rect 520 -1766 521 -1765
rect 597 -1766 598 -1765
rect 646 -1766 647 -1765
rect 240 -1768 241 -1767
rect 401 -1768 402 -1767
rect 443 -1768 444 -1767
rect 646 -1768 647 -1767
rect 44 -1770 45 -1769
rect 443 -1770 444 -1769
rect 44 -1772 45 -1771
rect 499 -1772 500 -1771
rect 240 -1774 241 -1773
rect 369 -1774 370 -1773
rect 499 -1774 500 -1773
rect 653 -1774 654 -1773
rect 254 -1776 255 -1775
rect 639 -1776 640 -1775
rect 653 -1776 654 -1775
rect 751 -1776 752 -1775
rect 184 -1778 185 -1777
rect 254 -1778 255 -1777
rect 275 -1778 276 -1777
rect 688 -1778 689 -1777
rect 184 -1780 185 -1779
rect 359 -1780 360 -1779
rect 583 -1780 584 -1779
rect 751 -1780 752 -1779
rect 212 -1782 213 -1781
rect 275 -1782 276 -1781
rect 282 -1782 283 -1781
rect 464 -1782 465 -1781
rect 583 -1782 584 -1781
rect 618 -1782 619 -1781
rect 93 -1784 94 -1783
rect 212 -1784 213 -1783
rect 282 -1784 283 -1783
rect 453 -1784 454 -1783
rect 464 -1784 465 -1783
rect 513 -1784 514 -1783
rect 618 -1784 619 -1783
rect 681 -1784 682 -1783
rect 289 -1786 290 -1785
rect 457 -1786 458 -1785
rect 562 -1786 563 -1785
rect 681 -1786 682 -1785
rect 180 -1788 181 -1787
rect 289 -1788 290 -1787
rect 296 -1788 297 -1787
rect 331 -1788 332 -1787
rect 352 -1788 353 -1787
rect 562 -1788 563 -1787
rect 296 -1790 297 -1789
rect 380 -1790 381 -1789
rect 401 -1790 402 -1789
rect 513 -1790 514 -1789
rect 299 -1792 300 -1791
rect 471 -1792 472 -1791
rect 317 -1794 318 -1793
rect 331 -1794 332 -1793
rect 359 -1794 360 -1793
rect 604 -1794 605 -1793
rect 604 -1796 605 -1795
rect 674 -1796 675 -1795
rect 632 -1798 633 -1797
rect 674 -1798 675 -1797
rect 352 -1800 353 -1799
rect 632 -1800 633 -1799
rect 9 -1811 10 -1810
rect 30 -1811 31 -1810
rect 33 -1811 34 -1810
rect 37 -1811 38 -1810
rect 40 -1811 41 -1810
rect 82 -1811 83 -1810
rect 89 -1811 90 -1810
rect 422 -1811 423 -1810
rect 471 -1811 472 -1810
rect 478 -1811 479 -1810
rect 492 -1811 493 -1810
rect 758 -1811 759 -1810
rect 23 -1813 24 -1812
rect 86 -1813 87 -1812
rect 93 -1813 94 -1812
rect 212 -1813 213 -1812
rect 219 -1813 220 -1812
rect 275 -1813 276 -1812
rect 306 -1813 307 -1812
rect 338 -1813 339 -1812
rect 345 -1813 346 -1812
rect 355 -1813 356 -1812
rect 366 -1813 367 -1812
rect 376 -1813 377 -1812
rect 380 -1813 381 -1812
rect 555 -1813 556 -1812
rect 579 -1813 580 -1812
rect 737 -1813 738 -1812
rect 44 -1815 45 -1814
rect 478 -1815 479 -1814
rect 492 -1815 493 -1814
rect 499 -1815 500 -1814
rect 506 -1815 507 -1814
rect 604 -1815 605 -1814
rect 674 -1815 675 -1814
rect 677 -1815 678 -1814
rect 737 -1815 738 -1814
rect 751 -1815 752 -1814
rect 51 -1817 52 -1816
rect 107 -1817 108 -1816
rect 121 -1817 122 -1816
rect 331 -1817 332 -1816
rect 348 -1817 349 -1816
rect 688 -1817 689 -1816
rect 65 -1819 66 -1818
rect 215 -1819 216 -1818
rect 219 -1819 220 -1818
rect 282 -1819 283 -1818
rect 331 -1819 332 -1818
rect 464 -1819 465 -1818
rect 495 -1819 496 -1818
rect 751 -1819 752 -1818
rect 65 -1821 66 -1820
rect 233 -1821 234 -1820
rect 240 -1821 241 -1820
rect 502 -1821 503 -1820
rect 513 -1821 514 -1820
rect 527 -1821 528 -1820
rect 604 -1821 605 -1820
rect 611 -1821 612 -1820
rect 653 -1821 654 -1820
rect 688 -1821 689 -1820
rect 72 -1823 73 -1822
rect 222 -1823 223 -1822
rect 240 -1823 241 -1822
rect 296 -1823 297 -1822
rect 352 -1823 353 -1822
rect 422 -1823 423 -1822
rect 464 -1823 465 -1822
rect 534 -1823 535 -1822
rect 611 -1823 612 -1822
rect 618 -1823 619 -1822
rect 674 -1823 675 -1822
rect 681 -1823 682 -1822
rect 72 -1825 73 -1824
rect 142 -1825 143 -1824
rect 149 -1825 150 -1824
rect 177 -1825 178 -1824
rect 184 -1825 185 -1824
rect 191 -1825 192 -1824
rect 201 -1825 202 -1824
rect 394 -1825 395 -1824
rect 415 -1825 416 -1824
rect 506 -1825 507 -1824
rect 516 -1825 517 -1824
rect 730 -1825 731 -1824
rect 47 -1827 48 -1826
rect 415 -1827 416 -1826
rect 453 -1827 454 -1826
rect 534 -1827 535 -1826
rect 618 -1827 619 -1826
rect 632 -1827 633 -1826
rect 681 -1827 682 -1826
rect 709 -1827 710 -1826
rect 79 -1829 80 -1828
rect 114 -1829 115 -1828
rect 121 -1829 122 -1828
rect 191 -1829 192 -1828
rect 268 -1829 269 -1828
rect 590 -1829 591 -1828
rect 695 -1829 696 -1828
rect 709 -1829 710 -1828
rect 93 -1831 94 -1830
rect 499 -1831 500 -1830
rect 509 -1831 510 -1830
rect 632 -1831 633 -1830
rect 695 -1831 696 -1830
rect 716 -1831 717 -1830
rect 103 -1833 104 -1832
rect 289 -1833 290 -1832
rect 296 -1833 297 -1832
rect 303 -1833 304 -1832
rect 338 -1833 339 -1832
rect 730 -1833 731 -1832
rect 107 -1835 108 -1834
rect 198 -1835 199 -1834
rect 275 -1835 276 -1834
rect 443 -1835 444 -1834
rect 520 -1835 521 -1834
rect 548 -1835 549 -1834
rect 590 -1835 591 -1834
rect 625 -1835 626 -1834
rect 677 -1835 678 -1834
rect 716 -1835 717 -1834
rect 100 -1837 101 -1836
rect 198 -1837 199 -1836
rect 282 -1837 283 -1836
rect 485 -1837 486 -1836
rect 625 -1837 626 -1836
rect 660 -1837 661 -1836
rect 124 -1839 125 -1838
rect 527 -1839 528 -1838
rect 642 -1839 643 -1838
rect 660 -1839 661 -1838
rect 128 -1841 129 -1840
rect 247 -1841 248 -1840
rect 352 -1841 353 -1840
rect 653 -1841 654 -1840
rect 135 -1843 136 -1842
rect 436 -1843 437 -1842
rect 443 -1843 444 -1842
rect 541 -1843 542 -1842
rect 142 -1845 143 -1844
rect 254 -1845 255 -1844
rect 355 -1845 356 -1844
rect 569 -1845 570 -1844
rect 156 -1847 157 -1846
rect 205 -1847 206 -1846
rect 247 -1847 248 -1846
rect 261 -1847 262 -1846
rect 310 -1847 311 -1846
rect 569 -1847 570 -1846
rect 16 -1849 17 -1848
rect 205 -1849 206 -1848
rect 254 -1849 255 -1848
rect 362 -1849 363 -1848
rect 369 -1849 370 -1848
rect 597 -1849 598 -1848
rect 16 -1851 17 -1850
rect 292 -1851 293 -1850
rect 310 -1851 311 -1850
rect 324 -1851 325 -1850
rect 359 -1851 360 -1850
rect 380 -1851 381 -1850
rect 387 -1851 388 -1850
rect 394 -1851 395 -1850
rect 450 -1851 451 -1850
rect 597 -1851 598 -1850
rect 163 -1853 164 -1852
rect 562 -1853 563 -1852
rect 12 -1855 13 -1854
rect 562 -1855 563 -1854
rect 131 -1857 132 -1856
rect 163 -1857 164 -1856
rect 166 -1857 167 -1856
rect 555 -1857 556 -1856
rect 170 -1859 171 -1858
rect 233 -1859 234 -1858
rect 261 -1859 262 -1858
rect 401 -1859 402 -1858
rect 485 -1859 486 -1858
rect 747 -1859 748 -1858
rect 135 -1861 136 -1860
rect 170 -1861 171 -1860
rect 173 -1861 174 -1860
rect 401 -1861 402 -1860
rect 187 -1863 188 -1862
rect 226 -1863 227 -1862
rect 268 -1863 269 -1862
rect 450 -1863 451 -1862
rect 114 -1865 115 -1864
rect 226 -1865 227 -1864
rect 324 -1865 325 -1864
rect 541 -1865 542 -1864
rect 373 -1867 374 -1866
rect 702 -1867 703 -1866
rect 303 -1869 304 -1868
rect 373 -1869 374 -1868
rect 387 -1869 388 -1868
rect 583 -1869 584 -1868
rect 390 -1871 391 -1870
rect 646 -1871 647 -1870
rect 180 -1873 181 -1872
rect 646 -1873 647 -1872
rect 408 -1875 409 -1874
rect 702 -1875 703 -1874
rect 408 -1877 409 -1876
rect 429 -1877 430 -1876
rect 576 -1877 577 -1876
rect 583 -1877 584 -1876
rect 317 -1879 318 -1878
rect 429 -1879 430 -1878
rect 138 -1881 139 -1880
rect 317 -1881 318 -1880
rect 2 -1892 3 -1891
rect 72 -1892 73 -1891
rect 107 -1892 108 -1891
rect 170 -1892 171 -1891
rect 177 -1892 178 -1891
rect 191 -1892 192 -1891
rect 194 -1892 195 -1891
rect 415 -1892 416 -1891
rect 432 -1892 433 -1891
rect 737 -1892 738 -1891
rect 5 -1894 6 -1893
rect 198 -1894 199 -1893
rect 201 -1894 202 -1893
rect 369 -1894 370 -1893
rect 376 -1894 377 -1893
rect 646 -1894 647 -1893
rect 709 -1894 710 -1893
rect 747 -1894 748 -1893
rect 9 -1896 10 -1895
rect 387 -1896 388 -1895
rect 397 -1896 398 -1895
rect 555 -1896 556 -1895
rect 12 -1898 13 -1897
rect 170 -1898 171 -1897
rect 177 -1898 178 -1897
rect 226 -1898 227 -1897
rect 240 -1898 241 -1897
rect 327 -1898 328 -1897
rect 338 -1898 339 -1897
rect 534 -1898 535 -1897
rect 541 -1898 542 -1897
rect 555 -1898 556 -1897
rect 23 -1900 24 -1899
rect 233 -1900 234 -1899
rect 292 -1900 293 -1899
rect 569 -1900 570 -1899
rect 23 -1902 24 -1901
rect 464 -1902 465 -1901
rect 471 -1902 472 -1901
rect 548 -1902 549 -1901
rect 562 -1902 563 -1901
rect 569 -1902 570 -1901
rect 33 -1904 34 -1903
rect 37 -1904 38 -1903
rect 44 -1904 45 -1903
rect 268 -1904 269 -1903
rect 296 -1904 297 -1903
rect 306 -1904 307 -1903
rect 317 -1904 318 -1903
rect 418 -1904 419 -1903
rect 436 -1904 437 -1903
rect 597 -1904 598 -1903
rect 26 -1906 27 -1905
rect 268 -1906 269 -1905
rect 296 -1906 297 -1905
rect 324 -1906 325 -1905
rect 345 -1906 346 -1905
rect 702 -1906 703 -1905
rect 51 -1908 52 -1907
rect 149 -1908 150 -1907
rect 156 -1908 157 -1907
rect 303 -1908 304 -1907
rect 324 -1908 325 -1907
rect 506 -1908 507 -1907
rect 520 -1908 521 -1907
rect 534 -1908 535 -1907
rect 541 -1908 542 -1907
rect 590 -1908 591 -1907
rect 597 -1908 598 -1907
rect 632 -1908 633 -1907
rect 674 -1908 675 -1907
rect 702 -1908 703 -1907
rect 51 -1910 52 -1909
rect 58 -1910 59 -1909
rect 61 -1910 62 -1909
rect 79 -1910 80 -1909
rect 117 -1910 118 -1909
rect 156 -1910 157 -1909
rect 184 -1910 185 -1909
rect 222 -1910 223 -1909
rect 254 -1910 255 -1909
rect 317 -1910 318 -1909
rect 359 -1910 360 -1909
rect 562 -1910 563 -1909
rect 590 -1910 591 -1909
rect 660 -1910 661 -1909
rect 667 -1910 668 -1909
rect 674 -1910 675 -1909
rect 65 -1912 66 -1911
rect 166 -1912 167 -1911
rect 184 -1912 185 -1911
rect 219 -1912 220 -1911
rect 303 -1912 304 -1911
rect 460 -1912 461 -1911
rect 471 -1912 472 -1911
rect 481 -1912 482 -1911
rect 502 -1912 503 -1911
rect 723 -1912 724 -1911
rect 65 -1914 66 -1913
rect 282 -1914 283 -1913
rect 331 -1914 332 -1913
rect 359 -1914 360 -1913
rect 362 -1914 363 -1913
rect 366 -1914 367 -1913
rect 380 -1914 381 -1913
rect 520 -1914 521 -1913
rect 625 -1914 626 -1913
rect 660 -1914 661 -1913
rect 16 -1916 17 -1915
rect 282 -1916 283 -1915
rect 366 -1916 367 -1915
rect 646 -1916 647 -1915
rect 72 -1918 73 -1917
rect 579 -1918 580 -1917
rect 618 -1918 619 -1917
rect 625 -1918 626 -1917
rect 639 -1918 640 -1917
rect 723 -1918 724 -1917
rect 79 -1920 80 -1919
rect 499 -1920 500 -1919
rect 506 -1920 507 -1919
rect 527 -1920 528 -1919
rect 618 -1920 619 -1919
rect 751 -1920 752 -1919
rect 19 -1922 20 -1921
rect 527 -1922 528 -1921
rect 114 -1924 115 -1923
rect 254 -1924 255 -1923
rect 261 -1924 262 -1923
rect 331 -1924 332 -1923
rect 380 -1924 381 -1923
rect 394 -1924 395 -1923
rect 401 -1924 402 -1923
rect 576 -1924 577 -1923
rect 100 -1926 101 -1925
rect 261 -1926 262 -1925
rect 355 -1926 356 -1925
rect 394 -1926 395 -1925
rect 401 -1926 402 -1925
rect 422 -1926 423 -1925
rect 429 -1926 430 -1925
rect 667 -1926 668 -1925
rect 100 -1928 101 -1927
rect 632 -1928 633 -1927
rect 128 -1930 129 -1929
rect 310 -1930 311 -1929
rect 429 -1930 430 -1929
rect 467 -1930 468 -1929
rect 131 -1932 132 -1931
rect 653 -1932 654 -1931
rect 145 -1934 146 -1933
rect 373 -1934 374 -1933
rect 436 -1934 437 -1933
rect 485 -1934 486 -1933
rect 205 -1936 206 -1935
rect 289 -1936 290 -1935
rect 310 -1936 311 -1935
rect 457 -1936 458 -1935
rect 485 -1936 486 -1935
rect 513 -1936 514 -1935
rect 149 -1938 150 -1937
rect 205 -1938 206 -1937
rect 208 -1938 209 -1937
rect 730 -1938 731 -1937
rect 142 -1940 143 -1939
rect 730 -1940 731 -1939
rect 86 -1942 87 -1941
rect 142 -1942 143 -1941
rect 212 -1942 213 -1941
rect 240 -1942 241 -1941
rect 271 -1942 272 -1941
rect 653 -1942 654 -1941
rect 86 -1944 87 -1943
rect 135 -1944 136 -1943
rect 163 -1944 164 -1943
rect 212 -1944 213 -1943
rect 219 -1944 220 -1943
rect 233 -1944 234 -1943
rect 352 -1944 353 -1943
rect 513 -1944 514 -1943
rect 135 -1946 136 -1945
rect 408 -1946 409 -1945
rect 439 -1946 440 -1945
rect 709 -1946 710 -1945
rect 275 -1948 276 -1947
rect 408 -1948 409 -1947
rect 443 -1948 444 -1947
rect 492 -1948 493 -1947
rect 247 -1950 248 -1949
rect 275 -1950 276 -1949
rect 422 -1950 423 -1949
rect 492 -1950 493 -1949
rect 93 -1952 94 -1951
rect 247 -1952 248 -1951
rect 450 -1952 451 -1951
rect 688 -1952 689 -1951
rect 37 -1954 38 -1953
rect 688 -1954 689 -1953
rect 93 -1956 94 -1955
rect 348 -1956 349 -1955
rect 450 -1956 451 -1955
rect 478 -1956 479 -1955
rect 478 -1958 479 -1957
rect 716 -1958 717 -1957
rect 695 -1960 696 -1959
rect 716 -1960 717 -1959
rect 681 -1962 682 -1961
rect 695 -1962 696 -1961
rect 54 -1964 55 -1963
rect 681 -1964 682 -1963
rect 16 -1975 17 -1974
rect 142 -1975 143 -1974
rect 156 -1975 157 -1974
rect 261 -1975 262 -1974
rect 285 -1975 286 -1974
rect 632 -1975 633 -1974
rect 635 -1975 636 -1974
rect 716 -1975 717 -1974
rect 19 -1977 20 -1976
rect 331 -1977 332 -1976
rect 366 -1977 367 -1976
rect 590 -1977 591 -1976
rect 642 -1977 643 -1976
rect 695 -1977 696 -1976
rect 23 -1979 24 -1978
rect 205 -1979 206 -1978
rect 240 -1979 241 -1978
rect 313 -1979 314 -1978
rect 324 -1979 325 -1978
rect 439 -1979 440 -1978
rect 450 -1979 451 -1978
rect 488 -1979 489 -1978
rect 534 -1979 535 -1978
rect 548 -1979 549 -1978
rect 551 -1979 552 -1978
rect 660 -1979 661 -1978
rect 695 -1979 696 -1978
rect 723 -1979 724 -1978
rect 23 -1981 24 -1980
rect 30 -1981 31 -1980
rect 37 -1981 38 -1980
rect 75 -1981 76 -1980
rect 100 -1981 101 -1980
rect 359 -1981 360 -1980
rect 366 -1981 367 -1980
rect 551 -1981 552 -1980
rect 562 -1981 563 -1980
rect 639 -1981 640 -1980
rect 30 -1983 31 -1982
rect 107 -1983 108 -1982
rect 110 -1983 111 -1982
rect 159 -1983 160 -1982
rect 163 -1983 164 -1982
rect 324 -1983 325 -1982
rect 331 -1983 332 -1982
rect 397 -1983 398 -1982
rect 404 -1983 405 -1982
rect 471 -1983 472 -1982
rect 478 -1983 479 -1982
rect 632 -1983 633 -1982
rect 44 -1985 45 -1984
rect 432 -1985 433 -1984
rect 443 -1985 444 -1984
rect 450 -1985 451 -1984
rect 457 -1985 458 -1984
rect 583 -1985 584 -1984
rect 618 -1985 619 -1984
rect 660 -1985 661 -1984
rect 44 -1987 45 -1986
rect 86 -1987 87 -1986
rect 93 -1987 94 -1986
rect 163 -1987 164 -1986
rect 170 -1987 171 -1986
rect 296 -1987 297 -1986
rect 303 -1987 304 -1986
rect 310 -1987 311 -1986
rect 369 -1987 370 -1986
rect 667 -1987 668 -1986
rect 51 -1989 52 -1988
rect 688 -1989 689 -1988
rect 58 -1991 59 -1990
rect 103 -1991 104 -1990
rect 107 -1991 108 -1990
rect 135 -1991 136 -1990
rect 142 -1991 143 -1990
rect 212 -1991 213 -1990
rect 219 -1991 220 -1990
rect 296 -1991 297 -1990
rect 387 -1991 388 -1990
rect 569 -1991 570 -1990
rect 583 -1991 584 -1990
rect 646 -1991 647 -1990
rect 65 -1993 66 -1992
rect 79 -1993 80 -1992
rect 100 -1993 101 -1992
rect 709 -1993 710 -1992
rect 2 -1995 3 -1994
rect 65 -1995 66 -1994
rect 68 -1995 69 -1994
rect 156 -1995 157 -1994
rect 177 -1995 178 -1994
rect 208 -1995 209 -1994
rect 215 -1995 216 -1994
rect 646 -1995 647 -1994
rect 72 -1997 73 -1996
rect 89 -1997 90 -1996
rect 117 -1997 118 -1996
rect 499 -1997 500 -1996
rect 534 -1997 535 -1996
rect 681 -1997 682 -1996
rect 117 -1999 118 -1998
rect 135 -1999 136 -1998
rect 149 -1999 150 -1998
rect 170 -1999 171 -1998
rect 177 -1999 178 -1998
rect 184 -1999 185 -1998
rect 191 -1999 192 -1998
rect 240 -1999 241 -1998
rect 254 -1999 255 -1998
rect 268 -1999 269 -1998
rect 289 -1999 290 -1998
rect 352 -1999 353 -1998
rect 387 -1999 388 -1998
rect 408 -1999 409 -1998
rect 415 -1999 416 -1998
rect 590 -1999 591 -1998
rect 604 -1999 605 -1998
rect 618 -1999 619 -1998
rect 9 -2001 10 -2000
rect 149 -2001 150 -2000
rect 184 -2001 185 -2000
rect 555 -2001 556 -2000
rect 562 -2001 563 -2000
rect 597 -2001 598 -2000
rect 604 -2001 605 -2000
rect 674 -2001 675 -2000
rect 9 -2003 10 -2002
rect 173 -2003 174 -2002
rect 219 -2003 220 -2002
rect 233 -2003 234 -2002
rect 247 -2003 248 -2002
rect 268 -2003 269 -2002
rect 289 -2003 290 -2002
rect 338 -2003 339 -2002
rect 380 -2003 381 -2002
rect 415 -2003 416 -2002
rect 418 -2003 419 -2002
rect 506 -2003 507 -2002
rect 569 -2003 570 -2002
rect 653 -2003 654 -2002
rect 54 -2005 55 -2004
rect 338 -2005 339 -2004
rect 394 -2005 395 -2004
rect 401 -2005 402 -2004
rect 408 -2005 409 -2004
rect 436 -2005 437 -2004
rect 443 -2005 444 -2004
rect 513 -2005 514 -2004
rect 597 -2005 598 -2004
rect 730 -2005 731 -2004
rect 54 -2007 55 -2006
rect 499 -2007 500 -2006
rect 506 -2007 507 -2006
rect 576 -2007 577 -2006
rect 642 -2007 643 -2006
rect 653 -2007 654 -2006
rect 121 -2009 122 -2008
rect 201 -2009 202 -2008
rect 226 -2009 227 -2008
rect 247 -2009 248 -2008
rect 261 -2009 262 -2008
rect 275 -2009 276 -2008
rect 422 -2009 423 -2008
rect 481 -2009 482 -2008
rect 513 -2009 514 -2008
rect 541 -2009 542 -2008
rect 576 -2009 577 -2008
rect 625 -2009 626 -2008
rect 128 -2011 129 -2010
rect 359 -2011 360 -2010
rect 457 -2011 458 -2010
rect 485 -2011 486 -2010
rect 541 -2011 542 -2010
rect 611 -2011 612 -2010
rect 625 -2011 626 -2010
rect 649 -2011 650 -2010
rect 121 -2013 122 -2012
rect 128 -2013 129 -2012
rect 131 -2013 132 -2012
rect 306 -2013 307 -2012
rect 464 -2013 465 -2012
rect 520 -2013 521 -2012
rect 611 -2013 612 -2012
rect 702 -2013 703 -2012
rect 226 -2015 227 -2014
rect 373 -2015 374 -2014
rect 474 -2015 475 -2014
rect 555 -2015 556 -2014
rect 233 -2017 234 -2016
rect 345 -2017 346 -2016
rect 373 -2017 374 -2016
rect 429 -2017 430 -2016
rect 492 -2017 493 -2016
rect 520 -2017 521 -2016
rect 275 -2019 276 -2018
rect 317 -2019 318 -2018
rect 429 -2019 430 -2018
rect 527 -2019 528 -2018
rect 282 -2021 283 -2020
rect 317 -2021 318 -2020
rect 348 -2021 349 -2020
rect 527 -2021 528 -2020
rect 282 -2023 283 -2022
rect 464 -2023 465 -2022
rect 303 -2025 304 -2024
rect 345 -2025 346 -2024
rect 436 -2025 437 -2024
rect 492 -2025 493 -2024
rect 9 -2036 10 -2035
rect 201 -2036 202 -2035
rect 212 -2036 213 -2035
rect 429 -2036 430 -2035
rect 436 -2036 437 -2035
rect 625 -2036 626 -2035
rect 632 -2036 633 -2035
rect 639 -2036 640 -2035
rect 646 -2036 647 -2035
rect 660 -2036 661 -2035
rect 688 -2036 689 -2035
rect 695 -2036 696 -2035
rect 16 -2038 17 -2037
rect 96 -2038 97 -2037
rect 114 -2038 115 -2037
rect 289 -2038 290 -2037
rect 303 -2038 304 -2037
rect 352 -2038 353 -2037
rect 380 -2038 381 -2037
rect 443 -2038 444 -2037
rect 474 -2038 475 -2037
rect 513 -2038 514 -2037
rect 520 -2038 521 -2037
rect 541 -2038 542 -2037
rect 548 -2038 549 -2037
rect 583 -2038 584 -2037
rect 16 -2040 17 -2039
rect 128 -2040 129 -2039
rect 191 -2040 192 -2039
rect 387 -2040 388 -2039
rect 415 -2040 416 -2039
rect 534 -2040 535 -2039
rect 541 -2040 542 -2039
rect 562 -2040 563 -2039
rect 30 -2042 31 -2041
rect 117 -2042 118 -2041
rect 128 -2042 129 -2041
rect 135 -2042 136 -2041
rect 191 -2042 192 -2041
rect 240 -2042 241 -2041
rect 257 -2042 258 -2041
rect 261 -2042 262 -2041
rect 289 -2042 290 -2041
rect 471 -2042 472 -2041
rect 481 -2042 482 -2041
rect 569 -2042 570 -2041
rect 37 -2044 38 -2043
rect 254 -2044 255 -2043
rect 303 -2044 304 -2043
rect 436 -2044 437 -2043
rect 443 -2044 444 -2043
rect 450 -2044 451 -2043
rect 471 -2044 472 -2043
rect 506 -2044 507 -2043
rect 548 -2044 549 -2043
rect 576 -2044 577 -2043
rect 33 -2046 34 -2045
rect 37 -2046 38 -2045
rect 44 -2046 45 -2045
rect 86 -2046 87 -2045
rect 100 -2046 101 -2045
rect 114 -2046 115 -2045
rect 117 -2046 118 -2045
rect 184 -2046 185 -2045
rect 198 -2046 199 -2045
rect 404 -2046 405 -2045
rect 425 -2046 426 -2045
rect 597 -2046 598 -2045
rect 44 -2048 45 -2047
rect 142 -2048 143 -2047
rect 194 -2048 195 -2047
rect 198 -2048 199 -2047
rect 205 -2048 206 -2047
rect 261 -2048 262 -2047
rect 313 -2048 314 -2047
rect 576 -2048 577 -2047
rect 51 -2050 52 -2049
rect 72 -2050 73 -2049
rect 79 -2050 80 -2049
rect 418 -2050 419 -2049
rect 429 -2050 430 -2049
rect 478 -2050 479 -2049
rect 485 -2050 486 -2049
rect 642 -2050 643 -2049
rect 51 -2052 52 -2051
rect 96 -2052 97 -2051
rect 212 -2052 213 -2051
rect 310 -2052 311 -2051
rect 320 -2052 321 -2051
rect 513 -2052 514 -2051
rect 555 -2052 556 -2051
rect 653 -2052 654 -2051
rect 65 -2054 66 -2053
rect 499 -2054 500 -2053
rect 555 -2054 556 -2053
rect 618 -2054 619 -2053
rect 642 -2054 643 -2053
rect 674 -2054 675 -2053
rect 65 -2056 66 -2055
rect 170 -2056 171 -2055
rect 215 -2056 216 -2055
rect 670 -2056 671 -2055
rect 75 -2058 76 -2057
rect 79 -2058 80 -2057
rect 86 -2058 87 -2057
rect 107 -2058 108 -2057
rect 170 -2058 171 -2057
rect 275 -2058 276 -2057
rect 327 -2058 328 -2057
rect 345 -2058 346 -2057
rect 359 -2058 360 -2057
rect 387 -2058 388 -2057
rect 418 -2058 419 -2057
rect 583 -2058 584 -2057
rect 107 -2060 108 -2059
rect 163 -2060 164 -2059
rect 219 -2060 220 -2059
rect 527 -2060 528 -2059
rect 562 -2060 563 -2059
rect 611 -2060 612 -2059
rect 58 -2062 59 -2061
rect 219 -2062 220 -2061
rect 222 -2062 223 -2061
rect 226 -2062 227 -2061
rect 236 -2062 237 -2061
rect 569 -2062 570 -2061
rect 604 -2062 605 -2061
rect 611 -2062 612 -2061
rect 58 -2064 59 -2063
rect 89 -2064 90 -2063
rect 149 -2064 150 -2063
rect 359 -2064 360 -2063
rect 383 -2064 384 -2063
rect 408 -2064 409 -2063
rect 450 -2064 451 -2063
rect 457 -2064 458 -2063
rect 492 -2064 493 -2063
rect 506 -2064 507 -2063
rect 149 -2066 150 -2065
rect 233 -2066 234 -2065
rect 240 -2066 241 -2065
rect 324 -2066 325 -2065
rect 331 -2066 332 -2065
rect 401 -2066 402 -2065
rect 408 -2066 409 -2065
rect 527 -2066 528 -2065
rect 135 -2068 136 -2067
rect 324 -2068 325 -2067
rect 338 -2068 339 -2067
rect 492 -2068 493 -2067
rect 499 -2068 500 -2067
rect 635 -2068 636 -2067
rect 156 -2070 157 -2069
rect 457 -2070 458 -2069
rect 142 -2072 143 -2071
rect 156 -2072 157 -2071
rect 159 -2072 160 -2071
rect 163 -2072 164 -2071
rect 222 -2072 223 -2071
rect 247 -2072 248 -2071
rect 254 -2072 255 -2071
rect 373 -2072 374 -2071
rect 394 -2072 395 -2071
rect 604 -2072 605 -2071
rect 226 -2074 227 -2073
rect 369 -2074 370 -2073
rect 373 -2074 374 -2073
rect 478 -2074 479 -2073
rect 268 -2076 269 -2075
rect 338 -2076 339 -2075
rect 345 -2076 346 -2075
rect 380 -2076 381 -2075
rect 394 -2076 395 -2075
rect 422 -2076 423 -2075
rect 268 -2078 269 -2077
rect 366 -2078 367 -2077
rect 401 -2078 402 -2077
rect 464 -2078 465 -2077
rect 275 -2080 276 -2079
rect 404 -2080 405 -2079
rect 317 -2082 318 -2081
rect 331 -2082 332 -2081
rect 352 -2082 353 -2081
rect 464 -2082 465 -2081
rect 317 -2084 318 -2083
rect 534 -2084 535 -2083
rect 366 -2086 367 -2085
rect 590 -2086 591 -2085
rect 282 -2088 283 -2087
rect 590 -2088 591 -2087
rect 282 -2090 283 -2089
rect 306 -2090 307 -2089
rect 23 -2101 24 -2100
rect 58 -2101 59 -2100
rect 65 -2101 66 -2100
rect 310 -2101 311 -2100
rect 324 -2101 325 -2100
rect 345 -2101 346 -2100
rect 366 -2101 367 -2100
rect 408 -2101 409 -2100
rect 509 -2101 510 -2100
rect 520 -2101 521 -2100
rect 523 -2101 524 -2100
rect 569 -2101 570 -2100
rect 590 -2101 591 -2100
rect 597 -2101 598 -2100
rect 611 -2101 612 -2100
rect 621 -2101 622 -2100
rect 642 -2101 643 -2100
rect 646 -2101 647 -2100
rect 674 -2101 675 -2100
rect 688 -2101 689 -2100
rect 26 -2103 27 -2102
rect 75 -2103 76 -2102
rect 107 -2103 108 -2102
rect 306 -2103 307 -2102
rect 310 -2103 311 -2102
rect 338 -2103 339 -2102
rect 345 -2103 346 -2102
rect 383 -2103 384 -2102
rect 394 -2103 395 -2102
rect 401 -2103 402 -2102
rect 530 -2103 531 -2102
rect 583 -2103 584 -2102
rect 611 -2103 612 -2102
rect 618 -2103 619 -2102
rect 33 -2105 34 -2104
rect 37 -2105 38 -2104
rect 44 -2105 45 -2104
rect 317 -2105 318 -2104
rect 331 -2105 332 -2104
rect 569 -2105 570 -2104
rect 37 -2107 38 -2106
rect 128 -2107 129 -2106
rect 135 -2107 136 -2106
rect 138 -2107 139 -2106
rect 156 -2107 157 -2106
rect 177 -2107 178 -2106
rect 187 -2107 188 -2106
rect 320 -2107 321 -2106
rect 338 -2107 339 -2106
rect 380 -2107 381 -2106
rect 387 -2107 388 -2106
rect 394 -2107 395 -2106
rect 534 -2107 535 -2106
rect 555 -2107 556 -2106
rect 562 -2107 563 -2106
rect 590 -2107 591 -2106
rect 44 -2109 45 -2108
rect 184 -2109 185 -2108
rect 208 -2109 209 -2108
rect 268 -2109 269 -2108
rect 282 -2109 283 -2108
rect 352 -2109 353 -2108
rect 359 -2109 360 -2108
rect 387 -2109 388 -2108
rect 464 -2109 465 -2108
rect 534 -2109 535 -2108
rect 51 -2111 52 -2110
rect 152 -2111 153 -2110
rect 163 -2111 164 -2110
rect 205 -2111 206 -2110
rect 215 -2111 216 -2110
rect 527 -2111 528 -2110
rect 51 -2113 52 -2112
rect 198 -2113 199 -2112
rect 205 -2113 206 -2112
rect 212 -2113 213 -2112
rect 222 -2113 223 -2112
rect 502 -2113 503 -2112
rect 58 -2115 59 -2114
rect 86 -2115 87 -2114
rect 107 -2115 108 -2114
rect 121 -2115 122 -2114
rect 135 -2115 136 -2114
rect 142 -2115 143 -2114
rect 149 -2115 150 -2114
rect 163 -2115 164 -2114
rect 170 -2115 171 -2114
rect 191 -2115 192 -2114
rect 198 -2115 199 -2114
rect 289 -2115 290 -2114
rect 303 -2115 304 -2114
rect 562 -2115 563 -2114
rect 65 -2117 66 -2116
rect 79 -2117 80 -2116
rect 86 -2117 87 -2116
rect 226 -2117 227 -2116
rect 233 -2117 234 -2116
rect 240 -2117 241 -2116
rect 247 -2117 248 -2116
rect 558 -2117 559 -2116
rect 16 -2119 17 -2118
rect 79 -2119 80 -2118
rect 138 -2119 139 -2118
rect 142 -2119 143 -2118
rect 170 -2119 171 -2118
rect 264 -2119 265 -2118
rect 268 -2119 269 -2118
rect 306 -2119 307 -2118
rect 369 -2119 370 -2118
rect 604 -2119 605 -2118
rect 72 -2121 73 -2120
rect 117 -2121 118 -2120
rect 177 -2121 178 -2120
rect 478 -2121 479 -2120
rect 117 -2123 118 -2122
rect 289 -2123 290 -2122
rect 233 -2125 234 -2124
rect 275 -2125 276 -2124
rect 240 -2127 241 -2126
rect 334 -2127 335 -2126
rect 247 -2129 248 -2128
rect 443 -2129 444 -2128
rect 254 -2131 255 -2130
rect 292 -2131 293 -2130
rect 443 -2131 444 -2130
rect 450 -2131 451 -2130
rect 226 -2133 227 -2132
rect 254 -2133 255 -2132
rect 261 -2133 262 -2132
rect 275 -2133 276 -2132
rect 450 -2133 451 -2132
rect 471 -2133 472 -2132
rect 261 -2135 262 -2134
rect 513 -2135 514 -2134
rect 422 -2137 423 -2136
rect 471 -2137 472 -2136
rect 513 -2137 514 -2136
rect 548 -2137 549 -2136
rect 422 -2139 423 -2138
rect 436 -2139 437 -2138
rect 492 -2139 493 -2138
rect 548 -2139 549 -2138
rect 373 -2141 374 -2140
rect 436 -2141 437 -2140
rect 492 -2141 493 -2140
rect 506 -2141 507 -2140
rect 373 -2143 374 -2142
rect 457 -2143 458 -2142
rect 457 -2145 458 -2144
rect 485 -2145 486 -2144
rect 485 -2147 486 -2146
rect 576 -2147 577 -2146
rect 9 -2158 10 -2157
rect 19 -2158 20 -2157
rect 37 -2158 38 -2157
rect 215 -2158 216 -2157
rect 240 -2158 241 -2157
rect 282 -2158 283 -2157
rect 285 -2158 286 -2157
rect 296 -2158 297 -2157
rect 317 -2158 318 -2157
rect 408 -2158 409 -2157
rect 415 -2158 416 -2157
rect 548 -2158 549 -2157
rect 590 -2158 591 -2157
rect 604 -2158 605 -2157
rect 44 -2160 45 -2159
rect 184 -2160 185 -2159
rect 208 -2160 209 -2159
rect 289 -2160 290 -2159
rect 292 -2160 293 -2159
rect 310 -2160 311 -2159
rect 317 -2160 318 -2159
rect 387 -2160 388 -2159
rect 408 -2160 409 -2159
rect 443 -2160 444 -2159
rect 450 -2160 451 -2159
rect 467 -2160 468 -2159
rect 499 -2160 500 -2159
rect 555 -2160 556 -2159
rect 597 -2160 598 -2159
rect 600 -2160 601 -2159
rect 51 -2162 52 -2161
rect 261 -2162 262 -2161
rect 275 -2162 276 -2161
rect 303 -2162 304 -2161
rect 324 -2162 325 -2161
rect 334 -2162 335 -2161
rect 352 -2162 353 -2161
rect 359 -2162 360 -2161
rect 362 -2162 363 -2161
rect 485 -2162 486 -2161
rect 541 -2162 542 -2161
rect 555 -2162 556 -2161
rect 51 -2164 52 -2163
rect 149 -2164 150 -2163
rect 163 -2164 164 -2163
rect 187 -2164 188 -2163
rect 247 -2164 248 -2163
rect 373 -2164 374 -2163
rect 387 -2164 388 -2163
rect 422 -2164 423 -2163
rect 425 -2164 426 -2163
rect 478 -2164 479 -2163
rect 58 -2166 59 -2165
rect 96 -2166 97 -2165
rect 107 -2166 108 -2165
rect 128 -2166 129 -2165
rect 131 -2166 132 -2165
rect 135 -2166 136 -2165
rect 163 -2166 164 -2165
rect 180 -2166 181 -2165
rect 268 -2166 269 -2165
rect 303 -2166 304 -2165
rect 324 -2166 325 -2165
rect 345 -2166 346 -2165
rect 352 -2166 353 -2165
rect 569 -2166 570 -2165
rect 58 -2168 59 -2167
rect 177 -2168 178 -2167
rect 278 -2168 279 -2167
rect 348 -2168 349 -2167
rect 366 -2168 367 -2167
rect 562 -2168 563 -2167
rect 65 -2170 66 -2169
rect 72 -2170 73 -2169
rect 79 -2170 80 -2169
rect 156 -2170 157 -2169
rect 177 -2170 178 -2169
rect 338 -2170 339 -2169
rect 345 -2170 346 -2169
rect 534 -2170 535 -2169
rect 40 -2172 41 -2171
rect 72 -2172 73 -2171
rect 86 -2172 87 -2171
rect 268 -2172 269 -2171
rect 296 -2172 297 -2171
rect 464 -2172 465 -2171
rect 513 -2172 514 -2171
rect 534 -2172 535 -2171
rect 65 -2174 66 -2173
rect 219 -2174 220 -2173
rect 331 -2174 332 -2173
rect 394 -2174 395 -2173
rect 415 -2174 416 -2173
rect 520 -2174 521 -2173
rect 86 -2176 87 -2175
rect 142 -2176 143 -2175
rect 156 -2176 157 -2175
rect 170 -2176 171 -2175
rect 219 -2176 220 -2175
rect 257 -2176 258 -2175
rect 394 -2176 395 -2175
rect 481 -2176 482 -2175
rect 93 -2178 94 -2177
rect 100 -2178 101 -2177
rect 107 -2178 108 -2177
rect 128 -2178 129 -2177
rect 135 -2178 136 -2177
rect 212 -2178 213 -2177
rect 429 -2178 430 -2177
rect 443 -2178 444 -2177
rect 453 -2178 454 -2177
rect 471 -2178 472 -2177
rect 93 -2180 94 -2179
rect 138 -2180 139 -2179
rect 205 -2180 206 -2179
rect 212 -2180 213 -2179
rect 429 -2180 430 -2179
rect 492 -2180 493 -2179
rect 100 -2182 101 -2181
rect 198 -2182 199 -2181
rect 380 -2182 381 -2181
rect 492 -2182 493 -2181
rect 121 -2184 122 -2183
rect 233 -2184 234 -2183
rect 380 -2184 381 -2183
rect 401 -2184 402 -2183
rect 436 -2184 437 -2183
rect 509 -2184 510 -2183
rect 121 -2186 122 -2185
rect 131 -2186 132 -2185
rect 170 -2186 171 -2185
rect 233 -2186 234 -2185
rect 436 -2186 437 -2185
rect 457 -2186 458 -2185
rect 198 -2188 199 -2187
rect 247 -2188 248 -2187
rect 457 -2188 458 -2187
rect 499 -2188 500 -2187
rect 226 -2190 227 -2189
rect 401 -2190 402 -2189
rect 191 -2192 192 -2191
rect 226 -2192 227 -2191
rect 187 -2194 188 -2193
rect 191 -2194 192 -2193
rect 9 -2205 10 -2204
rect 16 -2205 17 -2204
rect 23 -2205 24 -2204
rect 26 -2205 27 -2204
rect 51 -2205 52 -2204
rect 103 -2205 104 -2204
rect 107 -2205 108 -2204
rect 201 -2205 202 -2204
rect 240 -2205 241 -2204
rect 380 -2205 381 -2204
rect 408 -2205 409 -2204
rect 418 -2205 419 -2204
rect 429 -2205 430 -2204
rect 450 -2205 451 -2204
rect 457 -2205 458 -2204
rect 506 -2205 507 -2204
rect 534 -2205 535 -2204
rect 548 -2205 549 -2204
rect 600 -2205 601 -2204
rect 604 -2205 605 -2204
rect 51 -2207 52 -2206
rect 82 -2207 83 -2206
rect 86 -2207 87 -2206
rect 205 -2207 206 -2206
rect 254 -2207 255 -2206
rect 464 -2207 465 -2206
rect 537 -2207 538 -2206
rect 555 -2207 556 -2206
rect 58 -2209 59 -2208
rect 128 -2209 129 -2208
rect 149 -2209 150 -2208
rect 156 -2209 157 -2208
rect 177 -2209 178 -2208
rect 205 -2209 206 -2208
rect 254 -2209 255 -2208
rect 289 -2209 290 -2208
rect 299 -2209 300 -2208
rect 362 -2209 363 -2208
rect 366 -2209 367 -2208
rect 387 -2209 388 -2208
rect 394 -2209 395 -2208
rect 408 -2209 409 -2208
rect 422 -2209 423 -2208
rect 534 -2209 535 -2208
rect 58 -2211 59 -2210
rect 93 -2211 94 -2210
rect 100 -2211 101 -2210
rect 212 -2211 213 -2210
rect 247 -2211 248 -2210
rect 289 -2211 290 -2210
rect 303 -2211 304 -2210
rect 341 -2211 342 -2210
rect 359 -2211 360 -2210
rect 520 -2211 521 -2210
rect 65 -2213 66 -2212
rect 145 -2213 146 -2212
rect 149 -2213 150 -2212
rect 163 -2213 164 -2212
rect 177 -2213 178 -2212
rect 261 -2213 262 -2212
rect 268 -2213 269 -2212
rect 348 -2213 349 -2212
rect 373 -2213 374 -2212
rect 436 -2213 437 -2212
rect 443 -2213 444 -2212
rect 492 -2213 493 -2212
rect 79 -2215 80 -2214
rect 208 -2215 209 -2214
rect 247 -2215 248 -2214
rect 317 -2215 318 -2214
rect 324 -2215 325 -2214
rect 352 -2215 353 -2214
rect 107 -2217 108 -2216
rect 170 -2217 171 -2216
rect 187 -2217 188 -2216
rect 219 -2217 220 -2216
rect 268 -2217 269 -2216
rect 345 -2217 346 -2216
rect 114 -2219 115 -2218
rect 121 -2219 122 -2218
rect 191 -2219 192 -2218
rect 282 -2219 283 -2218
rect 72 -2221 73 -2220
rect 114 -2221 115 -2220
rect 191 -2221 192 -2220
rect 226 -2221 227 -2220
rect 275 -2221 276 -2220
rect 331 -2221 332 -2220
rect 226 -2223 227 -2222
rect 327 -2223 328 -2222
rect 331 -2223 332 -2222
rect 401 -2223 402 -2222
rect 58 -2234 59 -2233
rect 93 -2234 94 -2233
rect 107 -2234 108 -2233
rect 173 -2234 174 -2233
rect 201 -2234 202 -2233
rect 268 -2234 269 -2233
rect 275 -2234 276 -2233
rect 327 -2234 328 -2233
rect 331 -2234 332 -2233
rect 383 -2234 384 -2233
rect 408 -2234 409 -2233
rect 429 -2234 430 -2233
rect 450 -2234 451 -2233
rect 474 -2234 475 -2233
rect 485 -2234 486 -2233
rect 506 -2234 507 -2233
rect 75 -2236 76 -2235
rect 114 -2236 115 -2235
rect 131 -2236 132 -2235
rect 226 -2236 227 -2235
rect 240 -2236 241 -2235
rect 390 -2236 391 -2235
rect 149 -2238 150 -2237
rect 163 -2238 164 -2237
rect 219 -2238 220 -2237
rect 282 -2238 283 -2237
rect 289 -2238 290 -2237
rect 303 -2238 304 -2237
rect 310 -2238 311 -2237
rect 373 -2238 374 -2237
rect 247 -2240 248 -2239
rect 355 -2240 356 -2239
rect 254 -2242 255 -2241
rect 313 -2242 314 -2241
<< metal2 >>
rect 131 -5 132 1
rect 156 -5 157 1
rect 163 -5 164 1
rect 187 -5 188 1
rect 191 -5 192 1
rect 233 -5 234 1
rect 261 -5 262 1
rect 282 -5 283 1
rect 177 -5 178 -1
rect 212 -5 213 -1
rect 215 -5 216 -1
rect 247 -5 248 -1
rect 268 -5 269 -1
rect 278 -5 279 -1
rect 226 -5 227 -3
rect 257 -5 258 -3
rect 26 -15 27 -13
rect 26 -32 27 -14
rect 26 -15 27 -13
rect 26 -32 27 -14
rect 86 -32 87 -14
rect 163 -15 164 -13
rect 170 -15 171 -13
rect 219 -32 220 -14
rect 240 -32 241 -14
rect 261 -15 262 -13
rect 268 -15 269 -13
rect 345 -32 346 -14
rect 369 -32 370 -14
rect 401 -32 402 -14
rect 93 -32 94 -16
rect 100 -32 101 -16
rect 107 -17 108 -13
rect 110 -17 111 -13
rect 142 -17 143 -13
rect 226 -17 227 -13
rect 247 -17 248 -13
rect 289 -32 290 -16
rect 327 -17 328 -13
rect 331 -32 332 -16
rect 376 -32 377 -16
rect 380 -32 381 -16
rect 110 -32 111 -18
rect 254 -32 255 -18
rect 257 -19 258 -13
rect 387 -32 388 -18
rect 138 -21 139 -13
rect 142 -32 143 -20
rect 149 -32 150 -20
rect 166 -32 167 -20
rect 170 -32 171 -20
rect 177 -21 178 -13
rect 180 -32 181 -20
rect 233 -32 234 -20
rect 243 -21 244 -13
rect 247 -32 248 -20
rect 275 -32 276 -20
rect 418 -32 419 -20
rect 156 -23 157 -13
rect 177 -32 178 -22
rect 184 -32 185 -22
rect 212 -32 213 -22
rect 215 -32 216 -22
rect 296 -32 297 -22
rect 117 -25 118 -13
rect 156 -32 157 -24
rect 191 -25 192 -13
rect 352 -32 353 -24
rect 128 -32 129 -26
rect 191 -32 192 -26
rect 198 -27 199 -13
rect 303 -32 304 -26
rect 198 -32 199 -28
rect 208 -32 209 -28
rect 222 -29 223 -13
rect 261 -32 262 -28
rect 282 -29 283 -13
rect 359 -32 360 -28
rect 205 -31 206 -13
rect 268 -32 269 -30
rect 282 -32 283 -30
rect 317 -32 318 -30
rect 65 -75 66 -41
rect 93 -42 94 -40
rect 100 -75 101 -41
rect 184 -42 185 -40
rect 212 -42 213 -40
rect 359 -42 360 -40
rect 72 -44 73 -40
rect 128 -75 129 -43
rect 149 -44 150 -40
rect 180 -44 181 -40
rect 184 -75 185 -43
rect 198 -44 199 -40
rect 226 -75 227 -43
rect 373 -75 374 -43
rect 75 -75 76 -45
rect 149 -75 150 -45
rect 156 -46 157 -40
rect 198 -75 199 -45
rect 229 -46 230 -40
rect 261 -46 262 -40
rect 275 -46 276 -40
rect 278 -52 279 -45
rect 282 -46 283 -40
rect 408 -75 409 -45
rect 79 -75 80 -47
rect 215 -75 216 -47
rect 233 -48 234 -40
rect 313 -48 314 -40
rect 324 -48 325 -40
rect 387 -48 388 -40
rect 86 -50 87 -40
rect 222 -75 223 -49
rect 233 -75 234 -49
rect 240 -50 241 -40
rect 261 -75 262 -49
rect 268 -50 269 -40
rect 275 -75 276 -49
rect 317 -50 318 -40
rect 44 -75 45 -51
rect 86 -75 87 -51
rect 114 -52 115 -40
rect 156 -75 157 -51
rect 163 -75 164 -51
rect 212 -75 213 -51
rect 240 -75 241 -51
rect 247 -52 248 -40
rect 317 -75 318 -51
rect 107 -75 108 -53
rect 114 -75 115 -53
rect 117 -75 118 -53
rect 173 -75 174 -53
rect 191 -54 192 -40
rect 247 -75 248 -53
rect 282 -75 283 -53
rect 380 -54 381 -40
rect 121 -56 122 -40
rect 177 -56 178 -40
rect 205 -75 206 -55
rect 380 -75 381 -55
rect 121 -75 122 -57
rect 135 -58 136 -40
rect 170 -58 171 -40
rect 359 -75 360 -57
rect 131 -75 132 -59
rect 387 -75 388 -59
rect 135 -75 136 -61
rect 142 -62 143 -40
rect 170 -75 171 -61
rect 401 -62 402 -40
rect 285 -64 286 -40
rect 345 -64 346 -40
rect 289 -66 290 -40
rect 310 -75 311 -65
rect 331 -66 332 -40
rect 401 -75 402 -65
rect 219 -68 220 -40
rect 289 -75 290 -67
rect 296 -68 297 -40
rect 324 -75 325 -67
rect 338 -68 339 -40
rect 345 -75 346 -67
rect 219 -75 220 -69
rect 366 -75 367 -69
rect 254 -72 255 -40
rect 296 -75 297 -71
rect 303 -72 304 -40
rect 303 -75 304 -71
rect 303 -72 304 -40
rect 303 -75 304 -71
rect 338 -75 339 -71
rect 394 -72 395 -40
rect 51 -75 52 -73
rect 254 -75 255 -73
rect 257 -75 258 -73
rect 331 -75 332 -73
rect 352 -74 353 -40
rect 394 -75 395 -73
rect 44 -85 45 -83
rect 100 -120 101 -84
rect 121 -120 122 -84
rect 135 -85 136 -83
rect 159 -85 160 -83
rect 191 -85 192 -83
rect 194 -85 195 -83
rect 226 -120 227 -84
rect 250 -120 251 -84
rect 401 -85 402 -83
rect 51 -87 52 -83
rect 156 -120 157 -86
rect 163 -87 164 -83
rect 170 -120 171 -86
rect 201 -120 202 -86
rect 247 -87 248 -83
rect 254 -87 255 -83
rect 303 -87 304 -83
rect 331 -87 332 -83
rect 383 -120 384 -86
rect 394 -87 395 -83
rect 443 -120 444 -86
rect 58 -120 59 -88
rect 145 -89 146 -83
rect 205 -120 206 -88
rect 240 -89 241 -83
rect 257 -89 258 -83
rect 373 -89 374 -83
rect 401 -120 402 -88
rect 453 -120 454 -88
rect 65 -91 66 -83
rect 114 -91 115 -83
rect 128 -120 129 -90
rect 394 -120 395 -90
rect 65 -120 66 -92
rect 79 -93 80 -83
rect 86 -120 87 -92
rect 107 -93 108 -83
rect 131 -120 132 -92
rect 289 -93 290 -83
rect 317 -93 318 -83
rect 331 -120 332 -92
rect 352 -93 353 -83
rect 408 -93 409 -83
rect 93 -120 94 -94
rect 124 -95 125 -83
rect 142 -95 143 -83
rect 163 -120 164 -94
rect 212 -95 213 -83
rect 261 -95 262 -83
rect 271 -95 272 -83
rect 387 -95 388 -83
rect 408 -120 409 -94
rect 432 -95 433 -83
rect 107 -120 108 -96
rect 247 -120 248 -96
rect 275 -120 276 -96
rect 282 -120 283 -96
rect 289 -120 290 -96
rect 359 -97 360 -83
rect 366 -97 367 -83
rect 415 -120 416 -96
rect 96 -99 97 -83
rect 359 -120 360 -98
rect 149 -101 150 -83
rect 373 -120 374 -100
rect 149 -120 150 -102
rect 184 -103 185 -83
rect 212 -120 213 -102
rect 219 -103 220 -83
rect 222 -103 223 -83
rect 422 -120 423 -102
rect 177 -120 178 -104
rect 261 -120 262 -104
rect 278 -105 279 -83
rect 380 -105 381 -83
rect 184 -120 185 -106
rect 191 -120 192 -106
rect 215 -107 216 -83
rect 324 -107 325 -83
rect 338 -107 339 -83
rect 387 -120 388 -106
rect 79 -120 80 -108
rect 215 -120 216 -108
rect 233 -109 234 -83
rect 254 -120 255 -108
rect 271 -120 272 -108
rect 338 -120 339 -108
rect 345 -109 346 -83
rect 352 -120 353 -108
rect 198 -111 199 -83
rect 345 -120 346 -110
rect 240 -120 241 -112
rect 429 -120 430 -112
rect 278 -120 279 -114
rect 303 -120 304 -114
rect 310 -115 311 -83
rect 324 -120 325 -114
rect 296 -117 297 -83
rect 317 -120 318 -116
rect 296 -120 297 -118
rect 366 -120 367 -118
rect 37 -173 38 -129
rect 149 -130 150 -128
rect 156 -173 157 -129
rect 198 -130 199 -128
rect 215 -130 216 -128
rect 429 -130 430 -128
rect 436 -173 437 -129
rect 481 -173 482 -129
rect 44 -173 45 -131
rect 93 -132 94 -128
rect 110 -173 111 -131
rect 114 -173 115 -131
rect 128 -173 129 -131
rect 205 -132 206 -128
rect 219 -173 220 -131
rect 222 -132 223 -128
rect 226 -132 227 -128
rect 250 -132 251 -128
rect 254 -132 255 -128
rect 268 -173 269 -131
rect 275 -173 276 -131
rect 450 -173 451 -131
rect 51 -173 52 -133
rect 166 -134 167 -128
rect 170 -134 171 -128
rect 429 -173 430 -133
rect 58 -136 59 -128
rect 142 -136 143 -128
rect 145 -136 146 -128
rect 226 -173 227 -135
rect 233 -173 234 -135
rect 236 -136 237 -128
rect 247 -136 248 -128
rect 338 -136 339 -128
rect 359 -136 360 -128
rect 366 -173 367 -135
rect 380 -136 381 -128
rect 471 -173 472 -135
rect 58 -173 59 -137
rect 166 -173 167 -137
rect 170 -173 171 -137
rect 191 -138 192 -128
rect 236 -173 237 -137
rect 415 -138 416 -128
rect 72 -173 73 -139
rect 121 -140 122 -128
rect 131 -140 132 -128
rect 422 -140 423 -128
rect 79 -142 80 -128
rect 93 -173 94 -141
rect 177 -142 178 -128
rect 198 -173 199 -141
rect 254 -173 255 -141
rect 464 -173 465 -141
rect 79 -173 80 -143
rect 121 -173 122 -143
rect 184 -144 185 -128
rect 247 -173 248 -143
rect 261 -173 262 -143
rect 285 -173 286 -143
rect 289 -144 290 -128
rect 380 -173 381 -143
rect 387 -144 388 -128
rect 485 -173 486 -143
rect 89 -173 90 -145
rect 100 -146 101 -128
rect 103 -146 104 -128
rect 177 -173 178 -145
rect 191 -173 192 -145
rect 324 -146 325 -128
rect 352 -146 353 -128
rect 359 -173 360 -145
rect 401 -146 402 -128
rect 457 -173 458 -145
rect 100 -173 101 -147
rect 107 -148 108 -128
rect 117 -148 118 -128
rect 324 -173 325 -147
rect 345 -148 346 -128
rect 352 -173 353 -147
rect 415 -173 416 -147
rect 443 -148 444 -128
rect 138 -150 139 -128
rect 184 -173 185 -149
rect 208 -173 209 -149
rect 401 -173 402 -149
rect 86 -152 87 -128
rect 138 -173 139 -151
rect 282 -152 283 -128
rect 338 -173 339 -151
rect 296 -154 297 -128
rect 313 -173 314 -153
rect 317 -154 318 -128
rect 492 -173 493 -153
rect 296 -173 297 -155
rect 387 -173 388 -155
rect 303 -158 304 -128
rect 345 -173 346 -157
rect 306 -173 307 -159
rect 443 -173 444 -159
rect 310 -162 311 -128
rect 408 -162 409 -128
rect 317 -173 318 -163
rect 408 -173 409 -163
rect 320 -173 321 -165
rect 394 -166 395 -128
rect 373 -168 374 -128
rect 394 -173 395 -167
rect 331 -170 332 -128
rect 373 -173 374 -169
rect 331 -173 332 -171
rect 439 -172 440 -128
rect 16 -230 17 -182
rect 89 -183 90 -181
rect 100 -183 101 -181
rect 100 -230 101 -182
rect 100 -183 101 -181
rect 100 -230 101 -182
rect 114 -183 115 -181
rect 152 -183 153 -181
rect 191 -183 192 -181
rect 285 -230 286 -182
rect 292 -183 293 -181
rect 373 -183 374 -181
rect 380 -183 381 -181
rect 555 -230 556 -182
rect 583 -230 584 -182
rect 639 -230 640 -182
rect 30 -230 31 -184
rect 222 -230 223 -184
rect 226 -185 227 -181
rect 478 -230 479 -184
rect 534 -230 535 -184
rect 548 -185 549 -181
rect 37 -187 38 -181
rect 208 -187 209 -181
rect 212 -187 213 -181
rect 212 -230 213 -186
rect 212 -187 213 -181
rect 212 -230 213 -186
rect 254 -230 255 -186
rect 334 -187 335 -181
rect 380 -230 381 -186
rect 565 -230 566 -186
rect 37 -230 38 -188
rect 79 -189 80 -181
rect 86 -230 87 -188
rect 107 -230 108 -188
rect 114 -230 115 -188
rect 341 -230 342 -188
rect 387 -189 388 -181
rect 548 -230 549 -188
rect 44 -191 45 -181
rect 145 -191 146 -181
rect 191 -230 192 -190
rect 233 -191 234 -181
rect 257 -191 258 -181
rect 268 -191 269 -181
rect 275 -230 276 -190
rect 338 -191 339 -181
rect 366 -191 367 -181
rect 387 -230 388 -190
rect 464 -191 465 -181
rect 499 -230 500 -190
rect 51 -193 52 -181
rect 289 -193 290 -181
rect 296 -193 297 -181
rect 324 -193 325 -181
rect 450 -193 451 -181
rect 464 -230 465 -192
rect 471 -193 472 -181
rect 506 -230 507 -192
rect 58 -195 59 -181
rect 527 -230 528 -194
rect 58 -230 59 -196
rect 93 -230 94 -196
rect 121 -197 122 -181
rect 247 -197 248 -181
rect 261 -197 262 -181
rect 289 -230 290 -196
rect 306 -197 307 -181
rect 485 -197 486 -181
rect 65 -230 66 -198
rect 68 -199 69 -181
rect 72 -199 73 -181
rect 152 -230 153 -198
rect 156 -199 157 -181
rect 261 -230 262 -198
rect 278 -199 279 -181
rect 429 -199 430 -181
rect 443 -199 444 -181
rect 450 -230 451 -198
rect 457 -199 458 -181
rect 471 -230 472 -198
rect 79 -230 80 -200
rect 422 -230 423 -200
rect 436 -201 437 -181
rect 443 -230 444 -200
rect 89 -230 90 -202
rect 415 -203 416 -181
rect 103 -230 104 -204
rect 429 -230 430 -204
rect 121 -230 122 -206
rect 373 -230 374 -206
rect 408 -207 409 -181
rect 457 -230 458 -206
rect 124 -230 125 -208
rect 240 -230 241 -208
rect 243 -209 244 -181
rect 268 -230 269 -208
rect 282 -230 283 -208
rect 415 -230 416 -208
rect 128 -211 129 -181
rect 184 -230 185 -210
rect 187 -211 188 -181
rect 366 -230 367 -210
rect 408 -230 409 -210
rect 520 -230 521 -210
rect 82 -230 83 -212
rect 128 -230 129 -212
rect 135 -213 136 -181
rect 243 -230 244 -212
rect 317 -230 318 -212
rect 492 -213 493 -181
rect 135 -230 136 -214
rect 163 -230 164 -214
rect 170 -215 171 -181
rect 247 -230 248 -214
rect 324 -230 325 -214
rect 513 -230 514 -214
rect 142 -217 143 -181
rect 226 -230 227 -216
rect 233 -230 234 -216
rect 345 -217 346 -181
rect 401 -217 402 -181
rect 492 -230 493 -216
rect 96 -219 97 -181
rect 401 -230 402 -218
rect 142 -230 143 -220
rect 303 -230 304 -220
rect 331 -221 332 -181
rect 485 -230 486 -220
rect 170 -230 171 -222
rect 177 -223 178 -181
rect 198 -223 199 -181
rect 215 -223 216 -181
rect 310 -230 311 -222
rect 331 -230 332 -222
rect 345 -230 346 -222
rect 394 -223 395 -181
rect 156 -230 157 -224
rect 177 -230 178 -224
rect 198 -230 199 -224
rect 352 -225 353 -181
rect 359 -225 360 -181
rect 394 -230 395 -224
rect 205 -230 206 -226
rect 219 -227 220 -181
rect 359 -230 360 -226
rect 436 -230 437 -226
rect 149 -229 150 -181
rect 219 -230 220 -228
rect 16 -240 17 -238
rect 149 -240 150 -238
rect 180 -287 181 -239
rect 247 -240 248 -238
rect 285 -240 286 -238
rect 492 -240 493 -238
rect 499 -240 500 -238
rect 576 -287 577 -239
rect 586 -240 587 -238
rect 625 -287 626 -239
rect 639 -240 640 -238
rect 660 -287 661 -239
rect 30 -242 31 -238
rect 145 -287 146 -241
rect 184 -242 185 -238
rect 184 -287 185 -241
rect 184 -242 185 -238
rect 184 -287 185 -241
rect 205 -242 206 -238
rect 219 -287 220 -241
rect 240 -242 241 -238
rect 604 -287 605 -241
rect 653 -242 654 -238
rect 653 -287 654 -241
rect 653 -242 654 -238
rect 653 -287 654 -241
rect 30 -287 31 -243
rect 198 -244 199 -238
rect 205 -287 206 -243
rect 240 -287 241 -243
rect 243 -244 244 -238
rect 275 -244 276 -238
rect 278 -287 279 -243
rect 492 -287 493 -243
rect 506 -244 507 -238
rect 562 -287 563 -243
rect 44 -287 45 -245
rect 79 -287 80 -245
rect 82 -246 83 -238
rect 478 -246 479 -238
rect 481 -287 482 -245
rect 590 -287 591 -245
rect 51 -287 52 -247
rect 527 -248 528 -238
rect 534 -248 535 -238
rect 565 -248 566 -238
rect 58 -287 59 -249
rect 93 -250 94 -238
rect 103 -250 104 -238
rect 345 -250 346 -238
rect 352 -250 353 -238
rect 485 -250 486 -238
rect 513 -250 514 -238
rect 583 -287 584 -249
rect 72 -287 73 -251
rect 135 -252 136 -238
rect 156 -252 157 -238
rect 352 -287 353 -251
rect 362 -252 363 -238
rect 401 -252 402 -238
rect 408 -252 409 -238
rect 506 -287 507 -251
rect 555 -252 556 -238
rect 597 -287 598 -251
rect 86 -287 87 -253
rect 194 -287 195 -253
rect 198 -287 199 -253
rect 359 -287 360 -253
rect 366 -254 367 -238
rect 485 -287 486 -253
rect 558 -254 559 -238
rect 618 -287 619 -253
rect 93 -287 94 -255
rect 100 -256 101 -238
rect 124 -287 125 -255
rect 135 -287 136 -255
rect 156 -287 157 -255
rect 177 -256 178 -238
rect 212 -287 213 -255
rect 226 -256 227 -238
rect 247 -287 248 -255
rect 408 -287 409 -255
rect 422 -256 423 -238
rect 527 -287 528 -255
rect 100 -287 101 -257
rect 166 -258 167 -238
rect 226 -287 227 -257
rect 257 -258 258 -238
rect 268 -258 269 -238
rect 275 -287 276 -257
rect 285 -287 286 -257
rect 632 -287 633 -257
rect 254 -287 255 -259
rect 422 -287 423 -259
rect 429 -260 430 -238
rect 534 -287 535 -259
rect 268 -287 269 -261
rect 324 -262 325 -238
rect 331 -262 332 -238
rect 499 -287 500 -261
rect 233 -264 234 -238
rect 331 -287 332 -263
rect 338 -287 339 -263
rect 513 -287 514 -263
rect 289 -266 290 -238
rect 296 -287 297 -265
rect 303 -266 304 -238
rect 345 -287 346 -265
rect 380 -266 381 -238
rect 439 -287 440 -265
rect 443 -266 444 -238
rect 520 -287 521 -265
rect 114 -268 115 -238
rect 289 -287 290 -267
rect 310 -287 311 -267
rect 401 -287 402 -267
rect 415 -268 416 -238
rect 429 -287 430 -267
rect 457 -268 458 -238
rect 611 -287 612 -267
rect 114 -287 115 -269
rect 261 -270 262 -238
rect 282 -270 283 -238
rect 443 -287 444 -269
rect 457 -287 458 -269
rect 464 -270 465 -238
rect 471 -270 472 -238
rect 569 -287 570 -269
rect 128 -272 129 -238
rect 380 -287 381 -271
rect 387 -272 388 -238
rect 555 -287 556 -271
rect 107 -274 108 -238
rect 128 -287 129 -273
rect 152 -274 153 -238
rect 261 -287 262 -273
rect 299 -287 300 -273
rect 415 -287 416 -273
rect 107 -287 108 -275
rect 191 -276 192 -238
rect 222 -276 223 -238
rect 464 -287 465 -275
rect 152 -287 153 -277
rect 163 -278 164 -238
rect 170 -278 171 -238
rect 303 -287 304 -277
rect 313 -287 314 -277
rect 541 -278 542 -238
rect 40 -287 41 -279
rect 170 -287 171 -279
rect 317 -280 318 -238
rect 324 -287 325 -279
rect 366 -287 367 -279
rect 387 -287 388 -279
rect 394 -280 395 -238
rect 548 -287 549 -279
rect 215 -282 216 -238
rect 394 -287 395 -281
rect 450 -282 451 -238
rect 541 -287 542 -281
rect 215 -287 216 -283
rect 233 -287 234 -283
rect 373 -284 374 -238
rect 471 -287 472 -283
rect 163 -287 164 -285
rect 373 -287 374 -285
rect 436 -286 437 -238
rect 450 -287 451 -285
rect 9 -356 10 -296
rect 317 -297 318 -295
rect 320 -297 321 -295
rect 534 -297 535 -295
rect 653 -297 654 -295
rect 656 -356 657 -296
rect 660 -297 661 -295
rect 674 -356 675 -296
rect 30 -299 31 -295
rect 163 -299 164 -295
rect 191 -299 192 -295
rect 380 -299 381 -295
rect 387 -299 388 -295
rect 569 -299 570 -295
rect 653 -356 654 -298
rect 660 -356 661 -298
rect 30 -356 31 -300
rect 219 -301 220 -295
rect 247 -301 248 -295
rect 352 -301 353 -295
rect 359 -301 360 -295
rect 611 -301 612 -295
rect 44 -303 45 -295
rect 219 -356 220 -302
rect 247 -356 248 -302
rect 296 -356 297 -302
rect 310 -303 311 -295
rect 506 -303 507 -295
rect 534 -356 535 -302
rect 562 -303 563 -295
rect 569 -356 570 -302
rect 604 -303 605 -295
rect 611 -356 612 -302
rect 632 -303 633 -295
rect 51 -305 52 -295
rect 212 -356 213 -304
rect 215 -305 216 -295
rect 485 -305 486 -295
rect 506 -356 507 -304
rect 513 -305 514 -295
rect 562 -356 563 -304
rect 597 -305 598 -295
rect 604 -356 605 -304
rect 618 -305 619 -295
rect 58 -307 59 -295
rect 152 -356 153 -306
rect 156 -307 157 -295
rect 187 -356 188 -306
rect 191 -356 192 -306
rect 226 -307 227 -295
rect 254 -307 255 -295
rect 499 -307 500 -295
rect 597 -356 598 -306
rect 625 -307 626 -295
rect 65 -309 66 -295
rect 268 -309 269 -295
rect 289 -309 290 -295
rect 513 -356 514 -308
rect 79 -311 80 -295
rect 394 -311 395 -295
rect 401 -311 402 -295
rect 404 -331 405 -310
rect 429 -311 430 -295
rect 485 -356 486 -310
rect 79 -356 80 -312
rect 135 -313 136 -295
rect 170 -313 171 -295
rect 268 -356 269 -312
rect 289 -356 290 -312
rect 390 -356 391 -312
rect 401 -356 402 -312
rect 422 -313 423 -295
rect 432 -356 433 -312
rect 576 -313 577 -295
rect 23 -356 24 -314
rect 170 -356 171 -314
rect 205 -315 206 -295
rect 233 -315 234 -295
rect 240 -315 241 -295
rect 254 -356 255 -314
rect 257 -315 258 -295
rect 303 -315 304 -295
rect 310 -356 311 -314
rect 366 -315 367 -295
rect 373 -315 374 -295
rect 383 -356 384 -314
rect 408 -315 409 -295
rect 576 -356 577 -314
rect 86 -317 87 -295
rect 149 -317 150 -295
rect 313 -317 314 -295
rect 527 -317 528 -295
rect 86 -356 87 -318
rect 275 -356 276 -318
rect 317 -356 318 -318
rect 345 -319 346 -295
rect 352 -356 353 -318
rect 555 -319 556 -295
rect 26 -321 27 -295
rect 345 -356 346 -320
rect 373 -356 374 -320
rect 471 -321 472 -295
rect 478 -356 479 -320
rect 492 -321 493 -295
rect 527 -356 528 -320
rect 590 -321 591 -295
rect 93 -323 94 -295
rect 233 -356 234 -322
rect 331 -323 332 -295
rect 555 -356 556 -322
rect 93 -356 94 -324
rect 142 -325 143 -295
rect 261 -325 262 -295
rect 331 -356 332 -324
rect 338 -325 339 -295
rect 548 -325 549 -295
rect 100 -327 101 -295
rect 250 -327 251 -295
rect 324 -327 325 -295
rect 338 -356 339 -326
rect 341 -327 342 -295
rect 394 -356 395 -326
rect 408 -356 409 -326
rect 541 -327 542 -295
rect 548 -356 549 -326
rect 621 -356 622 -326
rect 100 -356 101 -328
rect 226 -356 227 -328
rect 415 -329 416 -295
rect 422 -356 423 -328
rect 436 -329 437 -295
rect 590 -356 591 -328
rect 110 -356 111 -330
rect 177 -331 178 -295
rect 222 -331 223 -295
rect 261 -356 262 -330
rect 415 -356 416 -330
rect 457 -331 458 -295
rect 471 -356 472 -330
rect 492 -356 493 -330
rect 520 -331 521 -295
rect 541 -356 542 -330
rect 583 -331 584 -295
rect 72 -333 73 -295
rect 177 -356 178 -332
rect 222 -356 223 -332
rect 362 -333 363 -295
rect 450 -333 451 -295
rect 520 -356 521 -332
rect 72 -356 73 -334
rect 198 -335 199 -295
rect 362 -356 363 -334
rect 429 -356 430 -334
rect 457 -356 458 -334
rect 464 -335 465 -295
rect 107 -337 108 -295
rect 198 -356 199 -336
rect 299 -337 300 -295
rect 464 -356 465 -336
rect 107 -356 108 -338
rect 436 -356 437 -338
rect 114 -341 115 -295
rect 282 -341 283 -295
rect 299 -356 300 -340
rect 443 -341 444 -295
rect 114 -356 115 -342
rect 303 -356 304 -342
rect 443 -356 444 -342
rect 453 -356 454 -342
rect 121 -356 122 -344
rect 163 -356 164 -344
rect 166 -345 167 -295
rect 583 -356 584 -344
rect 128 -347 129 -295
rect 240 -356 241 -346
rect 135 -356 136 -348
rect 278 -349 279 -295
rect 58 -356 59 -350
rect 278 -356 279 -350
rect 142 -356 143 -352
rect 184 -353 185 -295
rect 128 -356 129 -354
rect 184 -356 185 -354
rect 9 -366 10 -364
rect 117 -366 118 -364
rect 128 -366 129 -364
rect 285 -423 286 -365
rect 324 -366 325 -364
rect 639 -423 640 -365
rect 653 -366 654 -364
rect 670 -366 671 -364
rect 674 -366 675 -364
rect 681 -423 682 -365
rect 16 -423 17 -367
rect 142 -368 143 -364
rect 170 -368 171 -364
rect 436 -368 437 -364
rect 453 -368 454 -364
rect 569 -368 570 -364
rect 583 -368 584 -364
rect 653 -423 654 -367
rect 660 -368 661 -364
rect 674 -423 675 -367
rect 23 -370 24 -364
rect 121 -370 122 -364
rect 128 -423 129 -369
rect 208 -370 209 -364
rect 219 -370 220 -364
rect 499 -423 500 -369
rect 520 -370 521 -364
rect 667 -423 668 -369
rect 30 -372 31 -364
rect 324 -423 325 -371
rect 341 -423 342 -371
rect 401 -372 402 -364
rect 408 -372 409 -364
rect 569 -423 570 -371
rect 583 -423 584 -371
rect 611 -372 612 -364
rect 44 -423 45 -373
rect 194 -374 195 -364
rect 212 -374 213 -364
rect 408 -423 409 -373
rect 429 -374 430 -364
rect 618 -423 619 -373
rect 51 -423 52 -375
rect 180 -376 181 -364
rect 229 -423 230 -375
rect 632 -423 633 -375
rect 58 -378 59 -364
rect 296 -378 297 -364
rect 359 -423 360 -377
rect 492 -378 493 -364
rect 506 -378 507 -364
rect 520 -423 521 -377
rect 548 -378 549 -364
rect 611 -423 612 -377
rect 33 -423 34 -379
rect 548 -423 549 -379
rect 555 -380 556 -364
rect 646 -423 647 -379
rect 72 -382 73 -364
rect 152 -382 153 -364
rect 177 -382 178 -364
rect 250 -423 251 -381
rect 254 -382 255 -364
rect 296 -423 297 -381
rect 366 -382 367 -364
rect 457 -382 458 -364
rect 464 -382 465 -364
rect 492 -423 493 -381
rect 562 -382 563 -364
rect 625 -423 626 -381
rect 72 -423 73 -383
rect 86 -384 87 -364
rect 100 -423 101 -383
rect 163 -384 164 -364
rect 275 -384 276 -364
rect 373 -384 374 -364
rect 383 -384 384 -364
rect 576 -384 577 -364
rect 604 -384 605 -364
rect 660 -423 661 -383
rect 65 -423 66 -385
rect 163 -423 164 -385
rect 275 -423 276 -385
rect 303 -386 304 -364
rect 345 -386 346 -364
rect 464 -423 465 -385
rect 471 -386 472 -364
rect 576 -423 577 -385
rect 79 -388 80 -364
rect 222 -388 223 -364
rect 240 -388 241 -364
rect 303 -423 304 -387
rect 338 -388 339 -364
rect 345 -423 346 -387
rect 352 -388 353 -364
rect 457 -423 458 -387
rect 478 -388 479 -364
rect 506 -423 507 -387
rect 527 -388 528 -364
rect 604 -423 605 -387
rect 86 -423 87 -389
rect 264 -423 265 -389
rect 282 -390 283 -364
rect 366 -423 367 -389
rect 383 -423 384 -389
rect 527 -423 528 -389
rect 93 -392 94 -364
rect 222 -423 223 -391
rect 261 -392 262 -364
rect 282 -423 283 -391
rect 289 -392 290 -364
rect 373 -423 374 -391
rect 387 -392 388 -364
rect 450 -423 451 -391
rect 481 -423 482 -391
rect 590 -392 591 -364
rect 93 -423 94 -393
rect 159 -394 160 -364
rect 198 -394 199 -364
rect 240 -423 241 -393
rect 331 -394 332 -364
rect 352 -423 353 -393
rect 355 -394 356 -364
rect 590 -423 591 -393
rect 107 -396 108 -364
rect 166 -423 167 -395
rect 233 -396 234 -364
rect 289 -423 290 -395
rect 310 -396 311 -364
rect 331 -423 332 -395
rect 362 -396 363 -364
rect 562 -423 563 -395
rect 107 -423 108 -397
rect 261 -423 262 -397
rect 317 -398 318 -364
rect 362 -423 363 -397
rect 390 -398 391 -364
rect 597 -398 598 -364
rect 114 -423 115 -399
rect 555 -423 556 -399
rect 121 -423 122 -401
rect 327 -402 328 -364
rect 401 -423 402 -401
rect 415 -402 416 -364
rect 422 -402 423 -364
rect 429 -423 430 -401
rect 436 -423 437 -401
rect 443 -402 444 -364
rect 534 -402 535 -364
rect 597 -423 598 -401
rect 135 -404 136 -364
rect 177 -423 178 -403
rect 268 -404 269 -364
rect 422 -423 423 -403
rect 135 -423 136 -405
rect 156 -423 157 -405
rect 170 -423 171 -405
rect 233 -423 234 -405
rect 317 -423 318 -405
rect 513 -406 514 -364
rect 138 -423 139 -407
rect 254 -423 255 -407
rect 387 -423 388 -407
rect 534 -423 535 -407
rect 142 -423 143 -409
rect 215 -423 216 -409
rect 226 -410 227 -364
rect 268 -423 269 -409
rect 394 -410 395 -364
rect 415 -423 416 -409
rect 485 -410 486 -364
rect 513 -423 514 -409
rect 117 -423 118 -411
rect 485 -423 486 -411
rect 149 -414 150 -364
rect 198 -423 199 -413
rect 247 -414 248 -364
rect 394 -423 395 -413
rect 149 -423 150 -415
rect 191 -416 192 -364
rect 247 -423 248 -415
rect 443 -423 444 -415
rect 184 -423 185 -417
rect 226 -423 227 -417
rect 191 -423 192 -419
rect 541 -420 542 -364
rect 474 -423 475 -421
rect 541 -423 542 -421
rect 16 -433 17 -431
rect 243 -510 244 -432
rect 257 -433 258 -431
rect 366 -433 367 -431
rect 380 -433 381 -431
rect 513 -433 514 -431
rect 541 -433 542 -431
rect 544 -433 545 -431
rect 583 -433 584 -431
rect 702 -510 703 -432
rect 33 -510 34 -434
rect 142 -435 143 -431
rect 149 -435 150 -431
rect 166 -435 167 -431
rect 201 -435 202 -431
rect 562 -435 563 -431
rect 646 -435 647 -431
rect 674 -510 675 -434
rect 681 -435 682 -431
rect 681 -510 682 -434
rect 681 -435 682 -431
rect 681 -510 682 -434
rect 40 -437 41 -431
rect 212 -510 213 -436
rect 219 -510 220 -436
rect 548 -437 549 -431
rect 653 -437 654 -431
rect 688 -510 689 -436
rect 44 -439 45 -431
rect 513 -510 514 -438
rect 527 -439 528 -431
rect 583 -510 584 -438
rect 639 -439 640 -431
rect 653 -510 654 -438
rect 44 -510 45 -440
rect 156 -441 157 -431
rect 205 -441 206 -431
rect 464 -441 465 -431
rect 471 -441 472 -431
rect 625 -441 626 -431
rect 632 -441 633 -431
rect 639 -510 640 -440
rect 51 -443 52 -431
rect 383 -443 384 -431
rect 390 -443 391 -431
rect 576 -443 577 -431
rect 611 -443 612 -431
rect 625 -510 626 -442
rect 58 -510 59 -444
rect 296 -445 297 -431
rect 320 -445 321 -431
rect 429 -445 430 -431
rect 450 -445 451 -431
rect 611 -510 612 -444
rect 618 -445 619 -431
rect 632 -510 633 -444
rect 65 -447 66 -431
rect 205 -510 206 -446
rect 222 -447 223 -431
rect 562 -510 563 -446
rect 65 -510 66 -448
rect 348 -510 349 -448
rect 352 -449 353 -431
rect 366 -510 367 -448
rect 390 -510 391 -448
rect 667 -449 668 -431
rect 72 -451 73 -431
rect 173 -451 174 -431
rect 177 -451 178 -431
rect 667 -510 668 -450
rect 72 -510 73 -452
rect 198 -453 199 -431
rect 229 -453 230 -431
rect 240 -453 241 -431
rect 257 -510 258 -452
rect 464 -510 465 -452
rect 478 -453 479 -431
rect 646 -510 647 -452
rect 79 -510 80 -454
rect 121 -455 122 -431
rect 128 -455 129 -431
rect 131 -481 132 -454
rect 135 -510 136 -454
rect 254 -510 255 -454
rect 264 -455 265 -431
rect 415 -455 416 -431
rect 425 -510 426 -454
rect 590 -455 591 -431
rect 82 -457 83 -431
rect 149 -510 150 -456
rect 156 -510 157 -456
rect 303 -457 304 -431
rect 331 -457 332 -431
rect 429 -510 430 -456
rect 439 -510 440 -456
rect 478 -510 479 -456
rect 485 -457 486 -431
rect 527 -510 528 -456
rect 534 -457 535 -431
rect 590 -510 591 -456
rect 93 -459 94 -431
rect 163 -510 164 -458
rect 177 -510 178 -458
rect 338 -459 339 -431
rect 345 -459 346 -431
rect 380 -510 381 -458
rect 401 -459 402 -431
rect 471 -510 472 -458
rect 492 -459 493 -431
rect 534 -510 535 -458
rect 541 -510 542 -458
rect 597 -459 598 -431
rect 100 -461 101 -431
rect 331 -510 332 -460
rect 338 -510 339 -460
rect 408 -461 409 -431
rect 443 -461 444 -431
rect 485 -510 486 -460
rect 499 -461 500 -431
rect 618 -510 619 -460
rect 100 -510 101 -462
rect 198 -510 199 -462
rect 215 -463 216 -431
rect 415 -510 416 -462
rect 436 -463 437 -431
rect 499 -510 500 -462
rect 520 -463 521 -431
rect 576 -510 577 -462
rect 107 -465 108 -431
rect 247 -465 248 -431
rect 275 -465 276 -431
rect 520 -510 521 -464
rect 61 -467 62 -431
rect 275 -510 276 -466
rect 310 -467 311 -431
rect 408 -510 409 -466
rect 450 -510 451 -466
rect 709 -510 710 -466
rect 110 -510 111 -468
rect 443 -510 444 -468
rect 457 -469 458 -431
rect 492 -510 493 -468
rect 114 -471 115 -431
rect 569 -471 570 -431
rect 114 -510 115 -472
rect 362 -473 363 -431
rect 117 -475 118 -431
rect 373 -475 374 -431
rect 128 -510 129 -476
rect 327 -477 328 -431
rect 373 -510 374 -476
rect 184 -479 185 -431
rect 310 -510 311 -478
rect 355 -510 356 -478
rect 569 -510 570 -478
rect 86 -481 87 -431
rect 184 -510 185 -480
rect 191 -510 192 -480
rect 327 -510 328 -480
rect 359 -481 360 -431
rect 506 -481 507 -431
rect 544 -510 545 -480
rect 597 -510 598 -480
rect 86 -510 87 -482
rect 93 -510 94 -482
rect 194 -483 195 -431
rect 506 -510 507 -482
rect 215 -510 216 -484
rect 422 -485 423 -431
rect 226 -487 227 -431
rect 457 -510 458 -486
rect 226 -510 227 -488
rect 268 -489 269 -431
rect 359 -510 360 -488
rect 604 -489 605 -431
rect 229 -510 230 -490
rect 261 -491 262 -431
rect 268 -510 269 -490
rect 303 -510 304 -490
rect 422 -510 423 -490
rect 548 -510 549 -490
rect 555 -491 556 -431
rect 604 -510 605 -490
rect 37 -510 38 -492
rect 555 -510 556 -492
rect 233 -495 234 -431
rect 352 -510 353 -494
rect 233 -510 234 -496
rect 271 -510 272 -496
rect 240 -510 241 -498
rect 394 -499 395 -431
rect 247 -510 248 -500
rect 320 -510 321 -500
rect 387 -501 388 -431
rect 394 -510 395 -500
rect 261 -510 262 -502
rect 317 -503 318 -431
rect 317 -510 318 -504
rect 660 -505 661 -431
rect 282 -507 283 -431
rect 660 -510 661 -506
rect 282 -510 283 -508
rect 695 -510 696 -508
rect 16 -597 17 -519
rect 345 -597 346 -519
rect 348 -520 349 -518
rect 611 -520 612 -518
rect 23 -597 24 -521
rect 499 -522 500 -518
rect 558 -597 559 -521
rect 674 -522 675 -518
rect 26 -524 27 -518
rect 310 -524 311 -518
rect 324 -524 325 -518
rect 471 -524 472 -518
rect 502 -597 503 -523
rect 674 -597 675 -523
rect 30 -526 31 -518
rect 436 -597 437 -525
rect 460 -597 461 -525
rect 618 -526 619 -518
rect 30 -597 31 -527
rect 464 -528 465 -518
rect 611 -597 612 -527
rect 695 -528 696 -518
rect 37 -597 38 -529
rect 299 -530 300 -518
rect 310 -597 311 -529
rect 418 -597 419 -529
rect 464 -597 465 -529
rect 513 -530 514 -518
rect 618 -597 619 -529
rect 639 -530 640 -518
rect 44 -532 45 -518
rect 285 -532 286 -518
rect 296 -532 297 -518
rect 429 -532 430 -518
rect 513 -597 514 -531
rect 667 -532 668 -518
rect 44 -597 45 -533
rect 100 -534 101 -518
rect 107 -534 108 -518
rect 562 -534 563 -518
rect 576 -534 577 -518
rect 667 -597 668 -533
rect 58 -536 59 -518
rect 257 -536 258 -518
rect 282 -536 283 -518
rect 289 -536 290 -518
rect 327 -536 328 -518
rect 485 -536 486 -518
rect 562 -597 563 -535
rect 583 -536 584 -518
rect 639 -597 640 -535
rect 660 -536 661 -518
rect 51 -538 52 -518
rect 660 -597 661 -537
rect 58 -597 59 -539
rect 373 -540 374 -518
rect 387 -540 388 -518
rect 495 -597 496 -539
rect 65 -542 66 -518
rect 324 -597 325 -541
rect 352 -597 353 -541
rect 390 -542 391 -518
rect 401 -542 402 -518
rect 520 -542 521 -518
rect 65 -597 66 -543
rect 296 -597 297 -543
rect 306 -597 307 -543
rect 583 -597 584 -543
rect 68 -597 69 -545
rect 576 -597 577 -545
rect 72 -548 73 -518
rect 124 -548 125 -518
rect 128 -548 129 -518
rect 320 -548 321 -518
rect 355 -548 356 -518
rect 653 -548 654 -518
rect 54 -597 55 -549
rect 72 -597 73 -549
rect 79 -550 80 -518
rect 219 -550 220 -518
rect 240 -550 241 -518
rect 250 -592 251 -549
rect 254 -550 255 -518
rect 415 -550 416 -518
rect 425 -550 426 -518
rect 429 -597 430 -549
rect 520 -597 521 -549
rect 590 -550 591 -518
rect 79 -597 80 -551
rect 117 -597 118 -551
rect 131 -597 132 -551
rect 401 -597 402 -551
rect 404 -552 405 -518
rect 688 -552 689 -518
rect 86 -597 87 -553
rect 184 -554 185 -518
rect 194 -597 195 -553
rect 555 -554 556 -518
rect 93 -556 94 -518
rect 93 -597 94 -555
rect 93 -556 94 -518
rect 93 -597 94 -555
rect 114 -556 115 -518
rect 226 -597 227 -555
rect 233 -556 234 -518
rect 254 -597 255 -555
rect 285 -597 286 -555
rect 527 -556 528 -518
rect 541 -556 542 -518
rect 590 -597 591 -555
rect 107 -597 108 -557
rect 527 -597 528 -557
rect 541 -597 542 -557
rect 597 -558 598 -518
rect 114 -597 115 -559
rect 569 -560 570 -518
rect 135 -562 136 -518
rect 359 -597 360 -561
rect 366 -562 367 -518
rect 366 -597 367 -561
rect 366 -562 367 -518
rect 366 -597 367 -561
rect 387 -597 388 -561
rect 450 -562 451 -518
rect 478 -562 479 -518
rect 597 -597 598 -561
rect 135 -597 136 -563
rect 492 -564 493 -518
rect 569 -597 570 -563
rect 625 -564 626 -518
rect 145 -566 146 -518
rect 534 -566 535 -518
rect 625 -597 626 -565
rect 646 -566 647 -518
rect 170 -597 171 -567
rect 198 -597 199 -567
rect 201 -568 202 -518
rect 338 -568 339 -518
rect 408 -568 409 -518
rect 439 -568 440 -518
rect 478 -597 479 -567
rect 506 -568 507 -518
rect 534 -597 535 -567
rect 632 -568 633 -518
rect 177 -570 178 -518
rect 201 -597 202 -569
rect 205 -570 206 -518
rect 268 -597 269 -569
rect 289 -597 290 -569
rect 317 -570 318 -518
rect 320 -597 321 -569
rect 450 -597 451 -569
rect 506 -597 507 -569
rect 604 -570 605 -518
rect 163 -572 164 -518
rect 177 -597 178 -571
rect 184 -597 185 -571
rect 362 -572 363 -518
rect 394 -572 395 -518
rect 408 -597 409 -571
rect 411 -597 412 -571
rect 653 -597 654 -571
rect 159 -597 160 -573
rect 163 -597 164 -573
rect 205 -597 206 -573
rect 212 -597 213 -573
rect 215 -574 216 -518
rect 632 -597 633 -573
rect 215 -597 216 -575
rect 457 -576 458 -518
rect 492 -597 493 -575
rect 604 -597 605 -575
rect 219 -597 220 -577
rect 331 -578 332 -518
rect 422 -597 423 -577
rect 439 -597 440 -577
rect 457 -597 458 -577
rect 709 -578 710 -518
rect 233 -597 234 -579
rect 338 -597 339 -579
rect 548 -580 549 -518
rect 646 -597 647 -579
rect 681 -580 682 -518
rect 709 -597 710 -579
rect 121 -582 122 -518
rect 548 -597 549 -581
rect 121 -597 122 -583
rect 142 -584 143 -518
rect 173 -584 174 -518
rect 681 -597 682 -583
rect 142 -597 143 -585
rect 156 -586 157 -518
rect 240 -597 241 -585
rect 261 -586 262 -518
rect 275 -586 276 -518
rect 331 -597 332 -585
rect 243 -588 244 -518
rect 485 -597 486 -587
rect 247 -590 248 -518
rect 394 -597 395 -589
rect 149 -592 150 -518
rect 247 -597 248 -591
rect 261 -597 262 -591
rect 275 -597 276 -591
rect 443 -592 444 -518
rect 149 -597 150 -593
rect 191 -594 192 -518
rect 317 -597 318 -593
rect 380 -594 381 -518
rect 443 -597 444 -593
rect 702 -594 703 -518
rect 303 -596 304 -518
rect 380 -597 381 -595
rect 23 -607 24 -605
rect 376 -607 377 -605
rect 411 -607 412 -605
rect 583 -607 584 -605
rect 611 -607 612 -605
rect 737 -676 738 -606
rect 30 -609 31 -605
rect 702 -676 703 -608
rect 709 -609 710 -605
rect 765 -676 766 -608
rect 37 -611 38 -605
rect 72 -676 73 -610
rect 93 -611 94 -605
rect 103 -611 104 -605
rect 107 -611 108 -605
rect 562 -611 563 -605
rect 625 -611 626 -605
rect 625 -676 626 -610
rect 625 -611 626 -605
rect 625 -676 626 -610
rect 632 -611 633 -605
rect 772 -676 773 -610
rect 37 -676 38 -612
rect 184 -613 185 -605
rect 187 -676 188 -612
rect 201 -613 202 -605
rect 219 -676 220 -612
rect 660 -613 661 -605
rect 674 -613 675 -605
rect 751 -676 752 -612
rect 44 -615 45 -605
rect 65 -615 66 -605
rect 93 -676 94 -614
rect 380 -615 381 -605
rect 415 -676 416 -614
rect 527 -615 528 -605
rect 541 -615 542 -605
rect 688 -676 689 -614
rect 44 -676 45 -616
rect 215 -617 216 -605
rect 222 -617 223 -605
rect 723 -676 724 -616
rect 51 -676 52 -618
rect 352 -619 353 -605
rect 355 -676 356 -618
rect 744 -676 745 -618
rect 58 -621 59 -605
rect 65 -676 66 -620
rect 100 -621 101 -605
rect 198 -621 199 -605
rect 212 -676 213 -620
rect 222 -676 223 -620
rect 226 -621 227 -605
rect 226 -676 227 -620
rect 226 -621 227 -605
rect 226 -676 227 -620
rect 233 -621 234 -605
rect 338 -676 339 -620
rect 348 -621 349 -605
rect 562 -676 563 -620
rect 569 -621 570 -605
rect 660 -676 661 -620
rect 681 -621 682 -605
rect 758 -676 759 -620
rect 23 -676 24 -622
rect 58 -676 59 -622
rect 75 -676 76 -622
rect 233 -676 234 -622
rect 254 -623 255 -605
rect 254 -676 255 -622
rect 254 -623 255 -605
rect 254 -676 255 -622
rect 275 -676 276 -622
rect 387 -623 388 -605
rect 418 -623 419 -605
rect 506 -623 507 -605
rect 513 -623 514 -605
rect 716 -676 717 -622
rect 79 -625 80 -605
rect 100 -676 101 -624
rect 107 -676 108 -624
rect 142 -625 143 -605
rect 170 -625 171 -605
rect 191 -676 192 -624
rect 282 -676 283 -624
rect 527 -676 528 -624
rect 555 -625 556 -605
rect 695 -676 696 -624
rect 79 -676 80 -626
rect 205 -627 206 -605
rect 303 -627 304 -605
rect 331 -627 332 -605
rect 366 -627 367 -605
rect 366 -676 367 -626
rect 366 -627 367 -605
rect 366 -676 367 -626
rect 380 -676 381 -626
rect 401 -627 402 -605
rect 422 -627 423 -605
rect 443 -676 444 -626
rect 450 -627 451 -605
rect 569 -676 570 -626
rect 583 -676 584 -626
rect 632 -676 633 -626
rect 639 -627 640 -605
rect 709 -676 710 -626
rect 114 -676 115 -628
rect 261 -629 262 -605
rect 296 -629 297 -605
rect 331 -676 332 -628
rect 425 -676 426 -628
rect 653 -629 654 -605
rect 117 -631 118 -605
rect 247 -631 248 -605
rect 261 -676 262 -630
rect 408 -631 409 -605
rect 439 -631 440 -605
rect 534 -631 535 -605
rect 590 -631 591 -605
rect 653 -676 654 -630
rect 54 -633 55 -605
rect 439 -676 440 -632
rect 453 -676 454 -632
rect 639 -676 640 -632
rect 121 -635 122 -605
rect 387 -676 388 -634
rect 457 -635 458 -605
rect 611 -676 612 -634
rect 618 -635 619 -605
rect 681 -676 682 -634
rect 124 -676 125 -636
rect 674 -676 675 -636
rect 128 -639 129 -605
rect 359 -639 360 -605
rect 457 -676 458 -638
rect 520 -639 521 -605
rect 135 -641 136 -605
rect 513 -676 514 -640
rect 142 -676 143 -642
rect 401 -676 402 -642
rect 464 -643 465 -605
rect 555 -676 556 -642
rect 163 -645 164 -605
rect 170 -676 171 -644
rect 198 -676 199 -644
rect 590 -676 591 -644
rect 149 -647 150 -605
rect 163 -676 164 -646
rect 247 -676 248 -646
rect 268 -647 269 -605
rect 296 -676 297 -646
rect 422 -676 423 -646
rect 429 -647 430 -605
rect 464 -676 465 -646
rect 471 -647 472 -605
rect 534 -676 535 -646
rect 19 -676 20 -648
rect 149 -676 150 -648
rect 303 -676 304 -648
rect 404 -676 405 -648
rect 478 -649 479 -605
rect 520 -676 521 -648
rect 86 -651 87 -605
rect 268 -676 269 -650
rect 310 -651 311 -605
rect 408 -676 409 -650
rect 478 -676 479 -650
rect 667 -651 668 -605
rect 86 -676 87 -652
rect 285 -653 286 -605
rect 317 -653 318 -605
rect 730 -676 731 -652
rect 177 -655 178 -605
rect 310 -676 311 -654
rect 320 -655 321 -605
rect 576 -655 577 -605
rect 604 -655 605 -605
rect 667 -676 668 -654
rect 177 -676 178 -656
rect 240 -657 241 -605
rect 359 -676 360 -656
rect 446 -657 447 -605
rect 485 -657 486 -605
rect 541 -676 542 -656
rect 548 -657 549 -605
rect 604 -676 605 -656
rect 159 -676 160 -658
rect 240 -676 241 -658
rect 373 -659 374 -605
rect 576 -676 577 -658
rect 194 -661 195 -605
rect 285 -676 286 -660
rect 324 -661 325 -605
rect 373 -676 374 -660
rect 394 -661 395 -605
rect 429 -676 430 -660
rect 467 -676 468 -660
rect 485 -676 486 -660
rect 492 -661 493 -605
rect 646 -661 647 -605
rect 201 -676 202 -662
rect 548 -676 549 -662
rect 205 -676 206 -664
rect 394 -676 395 -664
rect 460 -676 461 -664
rect 646 -676 647 -664
rect 324 -676 325 -666
rect 618 -676 619 -666
rect 499 -669 500 -605
rect 597 -669 598 -605
rect 135 -676 136 -670
rect 597 -676 598 -670
rect 289 -673 290 -605
rect 499 -676 500 -672
rect 289 -676 290 -674
rect 317 -676 318 -674
rect 30 -686 31 -684
rect 457 -686 458 -684
rect 467 -686 468 -684
rect 758 -686 759 -684
rect 765 -686 766 -684
rect 793 -761 794 -685
rect 37 -688 38 -684
rect 324 -761 325 -687
rect 338 -688 339 -684
rect 338 -761 339 -687
rect 338 -688 339 -684
rect 338 -761 339 -687
rect 345 -688 346 -684
rect 639 -688 640 -684
rect 730 -688 731 -684
rect 779 -761 780 -687
rect 37 -761 38 -689
rect 107 -690 108 -684
rect 114 -690 115 -684
rect 422 -761 423 -689
rect 443 -690 444 -684
rect 471 -761 472 -689
rect 485 -690 486 -684
rect 492 -761 493 -689
rect 506 -690 507 -684
rect 765 -761 766 -689
rect 772 -690 773 -684
rect 849 -761 850 -689
rect 44 -692 45 -684
rect 355 -692 356 -684
rect 362 -761 363 -691
rect 366 -692 367 -684
rect 380 -692 381 -684
rect 457 -761 458 -691
rect 495 -692 496 -684
rect 772 -761 773 -691
rect 44 -761 45 -693
rect 93 -694 94 -684
rect 107 -761 108 -693
rect 303 -694 304 -684
rect 320 -694 321 -684
rect 555 -694 556 -684
rect 586 -694 587 -684
rect 751 -694 752 -684
rect 51 -696 52 -684
rect 436 -696 437 -684
rect 450 -761 451 -695
rect 590 -696 591 -684
rect 604 -696 605 -684
rect 639 -761 640 -695
rect 744 -696 745 -684
rect 786 -761 787 -695
rect 54 -761 55 -697
rect 352 -761 353 -697
rect 359 -698 360 -684
rect 366 -761 367 -697
rect 383 -761 384 -697
rect 702 -698 703 -684
rect 58 -761 59 -699
rect 61 -700 62 -684
rect 65 -700 66 -684
rect 327 -700 328 -684
rect 345 -761 346 -699
rect 355 -761 356 -699
rect 397 -700 398 -684
rect 681 -700 682 -684
rect 65 -761 66 -701
rect 499 -702 500 -684
rect 506 -761 507 -701
rect 513 -702 514 -684
rect 520 -702 521 -684
rect 520 -761 521 -701
rect 520 -702 521 -684
rect 520 -761 521 -701
rect 527 -702 528 -684
rect 527 -761 528 -701
rect 527 -702 528 -684
rect 527 -761 528 -701
rect 541 -702 542 -684
rect 541 -761 542 -701
rect 541 -702 542 -684
rect 541 -761 542 -701
rect 548 -702 549 -684
rect 548 -761 549 -701
rect 548 -702 549 -684
rect 548 -761 549 -701
rect 555 -761 556 -701
rect 562 -702 563 -684
rect 597 -702 598 -684
rect 604 -761 605 -701
rect 632 -702 633 -684
rect 758 -761 759 -701
rect 72 -704 73 -684
rect 744 -761 745 -703
rect 72 -761 73 -705
rect 93 -761 94 -705
rect 124 -706 125 -684
rect 289 -706 290 -684
rect 296 -706 297 -684
rect 464 -761 465 -705
rect 478 -761 479 -705
rect 632 -761 633 -705
rect 646 -706 647 -684
rect 681 -761 682 -705
rect 86 -708 87 -684
rect 187 -708 188 -684
rect 212 -708 213 -684
rect 212 -761 213 -707
rect 212 -708 213 -684
rect 212 -761 213 -707
rect 222 -708 223 -684
rect 310 -708 311 -684
rect 320 -761 321 -707
rect 733 -761 734 -707
rect 89 -761 90 -709
rect 404 -710 405 -684
rect 415 -710 416 -684
rect 590 -761 591 -709
rect 625 -710 626 -684
rect 646 -761 647 -709
rect 653 -710 654 -684
rect 702 -761 703 -709
rect 128 -712 129 -684
rect 261 -712 262 -684
rect 268 -712 269 -684
rect 282 -712 283 -684
rect 289 -761 290 -711
rect 509 -712 510 -684
rect 562 -761 563 -711
rect 569 -712 570 -684
rect 611 -712 612 -684
rect 653 -761 654 -711
rect 79 -714 80 -684
rect 268 -761 269 -713
rect 282 -761 283 -713
rect 751 -761 752 -713
rect 79 -761 80 -715
rect 723 -716 724 -684
rect 131 -761 132 -717
rect 387 -718 388 -684
rect 397 -761 398 -717
rect 688 -718 689 -684
rect 695 -718 696 -684
rect 723 -761 724 -717
rect 16 -761 17 -719
rect 688 -761 689 -719
rect 135 -722 136 -684
rect 583 -761 584 -721
rect 618 -722 619 -684
rect 625 -761 626 -721
rect 135 -761 136 -723
rect 205 -724 206 -684
rect 233 -724 234 -684
rect 394 -724 395 -684
rect 401 -724 402 -684
rect 737 -724 738 -684
rect 114 -761 115 -725
rect 401 -761 402 -725
rect 408 -726 409 -684
rect 415 -761 416 -725
rect 429 -726 430 -684
rect 597 -761 598 -725
rect 621 -761 622 -725
rect 695 -761 696 -725
rect 121 -728 122 -684
rect 233 -761 234 -727
rect 247 -728 248 -684
rect 306 -761 307 -727
rect 348 -728 349 -684
rect 481 -728 482 -684
rect 499 -761 500 -727
rect 534 -728 535 -684
rect 142 -730 143 -684
rect 674 -730 675 -684
rect 124 -761 125 -731
rect 142 -761 143 -731
rect 145 -732 146 -684
rect 159 -732 160 -684
rect 163 -732 164 -684
rect 408 -761 409 -731
rect 429 -761 430 -731
rect 660 -732 661 -684
rect 86 -761 87 -733
rect 660 -761 661 -733
rect 156 -736 157 -684
rect 716 -736 717 -684
rect 156 -761 157 -737
rect 222 -761 223 -737
rect 247 -761 248 -737
rect 303 -761 304 -737
rect 348 -761 349 -737
rect 716 -761 717 -737
rect 163 -761 164 -739
rect 278 -740 279 -684
rect 373 -740 374 -684
rect 387 -761 388 -739
rect 394 -761 395 -739
rect 569 -761 570 -739
rect 184 -742 185 -684
rect 737 -761 738 -741
rect 170 -744 171 -684
rect 184 -761 185 -743
rect 191 -744 192 -684
rect 205 -761 206 -743
rect 254 -744 255 -684
rect 275 -744 276 -684
rect 373 -761 374 -743
rect 488 -761 489 -743
rect 149 -746 150 -684
rect 275 -761 276 -745
rect 436 -761 437 -745
rect 674 -761 675 -745
rect 149 -761 150 -747
rect 709 -748 710 -684
rect 170 -761 171 -749
rect 226 -750 227 -684
rect 254 -761 255 -749
rect 313 -761 314 -749
rect 453 -750 454 -684
rect 513 -761 514 -749
rect 576 -750 577 -684
rect 709 -761 710 -749
rect 177 -752 178 -684
rect 191 -761 192 -751
rect 201 -752 202 -684
rect 611 -761 612 -751
rect 96 -761 97 -753
rect 177 -761 178 -753
rect 201 -761 202 -753
rect 296 -761 297 -753
rect 446 -761 447 -753
rect 576 -761 577 -753
rect 226 -761 227 -755
rect 240 -756 241 -684
rect 261 -761 262 -755
rect 331 -756 332 -684
rect 481 -761 482 -755
rect 667 -756 668 -684
rect 100 -758 101 -684
rect 331 -761 332 -757
rect 439 -758 440 -684
rect 667 -761 668 -757
rect 30 -761 31 -759
rect 100 -761 101 -759
rect 240 -761 241 -759
rect 292 -761 293 -759
rect 439 -761 440 -759
rect 534 -761 535 -759
rect 19 -771 20 -769
rect 23 -771 24 -769
rect 30 -850 31 -770
rect 394 -850 395 -770
rect 408 -771 409 -769
rect 485 -850 486 -770
rect 488 -771 489 -769
rect 835 -850 836 -770
rect 849 -771 850 -769
rect 940 -850 941 -770
rect 23 -850 24 -772
rect 149 -773 150 -769
rect 159 -850 160 -772
rect 275 -773 276 -769
rect 289 -773 290 -769
rect 296 -773 297 -769
rect 310 -773 311 -769
rect 513 -773 514 -769
rect 534 -773 535 -769
rect 709 -773 710 -769
rect 751 -773 752 -769
rect 814 -850 815 -772
rect 37 -775 38 -769
rect 152 -775 153 -769
rect 177 -775 178 -769
rect 180 -831 181 -774
rect 201 -775 202 -769
rect 261 -775 262 -769
rect 268 -775 269 -769
rect 282 -775 283 -769
rect 292 -775 293 -769
rect 457 -775 458 -769
rect 460 -850 461 -774
rect 562 -775 563 -769
rect 621 -775 622 -769
rect 772 -775 773 -769
rect 779 -775 780 -769
rect 849 -850 850 -774
rect 37 -850 38 -776
rect 432 -777 433 -769
rect 446 -777 447 -769
rect 702 -777 703 -769
rect 758 -777 759 -769
rect 828 -850 829 -776
rect 40 -850 41 -778
rect 275 -850 276 -778
rect 296 -850 297 -778
rect 618 -850 619 -778
rect 646 -779 647 -769
rect 779 -850 780 -778
rect 793 -779 794 -769
rect 863 -850 864 -778
rect 54 -850 55 -780
rect 65 -781 66 -769
rect 86 -781 87 -769
rect 219 -781 220 -769
rect 222 -781 223 -769
rect 660 -781 661 -769
rect 667 -781 668 -769
rect 709 -850 710 -780
rect 765 -781 766 -769
rect 842 -850 843 -780
rect 44 -783 45 -769
rect 219 -850 220 -782
rect 226 -783 227 -769
rect 282 -850 283 -782
rect 317 -783 318 -769
rect 345 -850 346 -782
rect 352 -783 353 -769
rect 765 -850 766 -782
rect 44 -850 45 -784
rect 156 -785 157 -769
rect 166 -850 167 -784
rect 646 -850 647 -784
rect 674 -785 675 -769
rect 807 -850 808 -784
rect 58 -787 59 -769
rect 96 -787 97 -769
rect 100 -787 101 -769
rect 310 -850 311 -786
rect 320 -787 321 -769
rect 597 -787 598 -769
rect 688 -787 689 -769
rect 856 -850 857 -786
rect 65 -850 66 -788
rect 464 -789 465 -769
rect 467 -850 468 -788
rect 737 -789 738 -769
rect 72 -791 73 -769
rect 667 -850 668 -790
rect 681 -791 682 -769
rect 737 -850 738 -790
rect 79 -793 80 -769
rect 597 -850 598 -792
rect 639 -793 640 -769
rect 681 -850 682 -792
rect 695 -793 696 -769
rect 751 -850 752 -792
rect 79 -850 80 -794
rect 107 -795 108 -769
rect 114 -850 115 -794
rect 135 -795 136 -769
rect 149 -850 150 -794
rect 289 -850 290 -794
rect 327 -850 328 -794
rect 397 -795 398 -769
rect 411 -850 412 -794
rect 716 -795 717 -769
rect 86 -850 87 -796
rect 730 -850 731 -796
rect 89 -799 90 -769
rect 89 -850 90 -798
rect 89 -799 90 -769
rect 89 -850 90 -798
rect 93 -850 94 -798
rect 362 -850 363 -798
rect 397 -850 398 -798
rect 786 -799 787 -769
rect 117 -801 118 -769
rect 583 -801 584 -769
rect 604 -801 605 -769
rect 639 -850 640 -800
rect 653 -801 654 -769
rect 688 -850 689 -800
rect 702 -850 703 -800
rect 723 -801 724 -769
rect 121 -803 122 -769
rect 401 -803 402 -769
rect 408 -850 409 -802
rect 604 -850 605 -802
rect 611 -803 612 -769
rect 653 -850 654 -802
rect 723 -850 724 -802
rect 744 -803 745 -769
rect 72 -850 73 -804
rect 121 -850 122 -804
rect 135 -850 136 -804
rect 191 -805 192 -769
rect 198 -805 199 -769
rect 432 -850 433 -804
rect 436 -850 437 -804
rect 786 -850 787 -804
rect 152 -850 153 -806
rect 317 -850 318 -806
rect 338 -807 339 -769
rect 443 -807 444 -769
rect 446 -850 447 -806
rect 772 -850 773 -806
rect 58 -850 59 -808
rect 338 -850 339 -808
rect 352 -850 353 -808
rect 373 -809 374 -769
rect 429 -809 430 -769
rect 660 -850 661 -808
rect 674 -850 675 -808
rect 744 -850 745 -808
rect 156 -850 157 -810
rect 191 -850 192 -810
rect 212 -811 213 -769
rect 212 -850 213 -810
rect 212 -811 213 -769
rect 212 -850 213 -810
rect 226 -850 227 -810
rect 380 -811 381 -769
rect 401 -850 402 -810
rect 429 -850 430 -810
rect 464 -850 465 -810
rect 583 -850 584 -810
rect 625 -811 626 -769
rect 695 -850 696 -810
rect 177 -850 178 -812
rect 184 -813 185 -769
rect 233 -813 234 -769
rect 373 -850 374 -812
rect 513 -850 514 -812
rect 870 -850 871 -812
rect 170 -815 171 -769
rect 233 -850 234 -814
rect 240 -815 241 -769
rect 243 -815 244 -769
rect 247 -815 248 -769
rect 250 -850 251 -814
rect 254 -815 255 -769
rect 516 -850 517 -814
rect 520 -815 521 -769
rect 534 -850 535 -814
rect 537 -815 538 -769
rect 716 -850 717 -814
rect 142 -817 143 -769
rect 170 -850 171 -816
rect 184 -850 185 -816
rect 240 -850 241 -816
rect 387 -817 388 -769
rect 548 -817 549 -769
rect 562 -850 563 -816
rect 569 -817 570 -769
rect 758 -850 759 -816
rect 142 -850 143 -818
rect 590 -819 591 -769
rect 163 -821 164 -769
rect 254 -850 255 -820
rect 268 -850 269 -820
rect 457 -850 458 -820
rect 499 -821 500 -769
rect 548 -850 549 -820
rect 555 -821 556 -769
rect 569 -850 570 -820
rect 576 -821 577 -769
rect 625 -850 626 -820
rect 128 -823 129 -769
rect 576 -850 577 -822
rect 128 -850 129 -824
rect 422 -825 423 -769
rect 471 -825 472 -769
rect 499 -850 500 -824
rect 541 -825 542 -769
rect 555 -850 556 -824
rect 163 -850 164 -826
rect 324 -827 325 -769
rect 331 -827 332 -769
rect 520 -850 521 -826
rect 527 -827 528 -769
rect 541 -850 542 -826
rect 107 -850 108 -828
rect 324 -850 325 -828
rect 331 -850 332 -828
rect 800 -850 801 -828
rect 243 -850 244 -830
rect 387 -850 388 -830
rect 471 -850 472 -830
rect 492 -831 493 -769
rect 506 -831 507 -769
rect 527 -850 528 -830
rect 299 -850 300 -832
rect 422 -850 423 -832
rect 506 -850 507 -832
rect 821 -850 822 -832
rect 306 -835 307 -769
rect 590 -850 591 -834
rect 100 -850 101 -836
rect 306 -850 307 -836
rect 355 -837 356 -769
rect 415 -837 416 -769
rect 359 -839 360 -769
rect 611 -850 612 -838
rect 198 -850 199 -840
rect 359 -850 360 -840
rect 366 -841 367 -769
rect 415 -850 416 -840
rect 366 -850 367 -842
rect 632 -843 633 -769
rect 383 -850 384 -844
rect 492 -850 493 -844
rect 450 -847 451 -769
rect 632 -850 633 -846
rect 450 -850 451 -848
rect 478 -850 479 -848
rect 9 -927 10 -859
rect 593 -927 594 -859
rect 674 -860 675 -858
rect 863 -860 864 -858
rect 16 -927 17 -861
rect 191 -862 192 -858
rect 201 -927 202 -861
rect 278 -927 279 -861
rect 282 -862 283 -858
rect 334 -862 335 -858
rect 338 -862 339 -858
rect 366 -862 367 -858
rect 404 -927 405 -861
rect 562 -862 563 -858
rect 576 -862 577 -858
rect 576 -927 577 -861
rect 576 -862 577 -858
rect 576 -927 577 -861
rect 660 -862 661 -858
rect 674 -927 675 -861
rect 831 -927 832 -861
rect 940 -862 941 -858
rect 30 -864 31 -858
rect 222 -927 223 -863
rect 240 -864 241 -858
rect 306 -864 307 -858
rect 317 -864 318 -858
rect 408 -927 409 -863
rect 411 -864 412 -858
rect 786 -864 787 -858
rect 44 -866 45 -858
rect 159 -866 160 -858
rect 163 -866 164 -858
rect 793 -927 794 -865
rect 44 -927 45 -867
rect 352 -868 353 -858
rect 359 -868 360 -858
rect 534 -868 535 -858
rect 562 -927 563 -867
rect 611 -868 612 -858
rect 653 -868 654 -858
rect 660 -927 661 -867
rect 58 -870 59 -858
rect 250 -927 251 -869
rect 261 -870 262 -858
rect 366 -927 367 -869
rect 429 -870 430 -858
rect 814 -870 815 -858
rect 72 -872 73 -858
rect 639 -872 640 -858
rect 653 -927 654 -871
rect 730 -872 731 -858
rect 744 -872 745 -858
rect 814 -927 815 -871
rect 72 -927 73 -873
rect 107 -874 108 -858
rect 121 -874 122 -858
rect 124 -927 125 -873
rect 135 -874 136 -858
rect 264 -874 265 -858
rect 268 -874 269 -858
rect 324 -927 325 -873
rect 327 -874 328 -858
rect 856 -874 857 -858
rect 23 -876 24 -858
rect 135 -927 136 -875
rect 142 -876 143 -858
rect 289 -876 290 -858
rect 317 -927 318 -875
rect 380 -876 381 -858
rect 387 -876 388 -858
rect 429 -927 430 -875
rect 443 -927 444 -875
rect 835 -876 836 -858
rect 23 -927 24 -877
rect 520 -878 521 -858
rect 590 -878 591 -858
rect 786 -927 787 -877
rect 75 -880 76 -858
rect 373 -880 374 -858
rect 387 -927 388 -879
rect 422 -880 423 -858
rect 453 -927 454 -879
rect 527 -880 528 -858
rect 597 -880 598 -858
rect 639 -927 640 -879
rect 730 -927 731 -879
rect 758 -880 759 -858
rect 79 -882 80 -858
rect 296 -882 297 -858
rect 310 -882 311 -858
rect 422 -927 423 -881
rect 457 -927 458 -881
rect 499 -882 500 -858
rect 506 -882 507 -858
rect 709 -882 710 -858
rect 744 -927 745 -881
rect 765 -882 766 -858
rect 79 -927 80 -883
rect 527 -927 528 -883
rect 611 -927 612 -883
rect 625 -884 626 -858
rect 702 -884 703 -858
rect 758 -927 759 -883
rect 765 -927 766 -883
rect 800 -884 801 -858
rect 82 -927 83 -885
rect 485 -886 486 -858
rect 506 -927 507 -885
rect 688 -886 689 -858
rect 709 -927 710 -885
rect 737 -886 738 -858
rect 800 -927 801 -885
rect 828 -886 829 -858
rect 86 -888 87 -858
rect 114 -888 115 -858
rect 142 -927 143 -887
rect 163 -927 164 -887
rect 166 -927 167 -887
rect 177 -888 178 -858
rect 184 -888 185 -858
rect 310 -927 311 -887
rect 345 -888 346 -858
rect 373 -927 374 -887
rect 439 -888 440 -858
rect 499 -927 500 -887
rect 534 -927 535 -887
rect 828 -927 829 -887
rect 30 -927 31 -889
rect 345 -927 346 -889
rect 362 -890 363 -858
rect 436 -927 437 -889
rect 460 -890 461 -858
rect 842 -890 843 -858
rect 51 -892 52 -858
rect 114 -927 115 -891
rect 177 -927 178 -891
rect 226 -892 227 -858
rect 233 -892 234 -858
rect 268 -927 269 -891
rect 464 -927 465 -891
rect 597 -927 598 -891
rect 625 -927 626 -891
rect 695 -892 696 -858
rect 737 -927 738 -891
rect 751 -892 752 -858
rect 842 -927 843 -891
rect 870 -892 871 -858
rect 40 -927 41 -893
rect 233 -927 234 -893
rect 254 -894 255 -858
rect 289 -927 290 -893
rect 467 -927 468 -893
rect 569 -894 570 -858
rect 583 -894 584 -858
rect 702 -927 703 -893
rect 751 -927 752 -893
rect 772 -894 773 -858
rect 51 -927 52 -895
rect 415 -896 416 -858
rect 478 -896 479 -858
rect 516 -896 517 -858
rect 555 -896 556 -858
rect 569 -927 570 -895
rect 681 -896 682 -858
rect 688 -927 689 -895
rect 695 -927 696 -895
rect 779 -896 780 -858
rect 86 -927 87 -897
rect 156 -898 157 -858
rect 170 -898 171 -858
rect 226 -927 227 -897
rect 254 -927 255 -897
rect 299 -927 300 -897
rect 471 -898 472 -858
rect 516 -927 517 -897
rect 541 -898 542 -858
rect 555 -927 556 -897
rect 667 -898 668 -858
rect 681 -927 682 -897
rect 716 -898 717 -858
rect 779 -927 780 -897
rect 93 -900 94 -858
rect 149 -927 150 -899
rect 156 -927 157 -899
rect 282 -927 283 -899
rect 446 -900 447 -858
rect 667 -927 668 -899
rect 716 -927 717 -899
rect 723 -900 724 -858
rect 772 -927 773 -899
rect 821 -900 822 -858
rect 93 -927 94 -901
rect 401 -902 402 -858
rect 471 -927 472 -901
rect 492 -902 493 -858
rect 646 -902 647 -858
rect 723 -927 724 -901
rect 821 -927 822 -901
rect 849 -902 850 -858
rect 54 -927 55 -903
rect 492 -927 493 -903
rect 632 -904 633 -858
rect 646 -927 647 -903
rect 835 -927 836 -903
rect 849 -927 850 -903
rect 100 -906 101 -858
rect 807 -906 808 -858
rect 65 -908 66 -858
rect 100 -927 101 -907
rect 103 -908 104 -858
rect 348 -927 349 -907
rect 401 -927 402 -907
rect 583 -927 584 -907
rect 618 -908 619 -858
rect 632 -927 633 -907
rect 107 -927 108 -909
rect 145 -910 146 -858
rect 191 -927 192 -909
rect 198 -910 199 -858
rect 205 -910 206 -858
rect 359 -927 360 -909
rect 485 -927 486 -909
rect 590 -927 591 -909
rect 604 -910 605 -858
rect 618 -927 619 -909
rect 58 -927 59 -911
rect 198 -927 199 -911
rect 212 -912 213 -858
rect 240 -927 241 -911
rect 261 -927 262 -911
rect 338 -927 339 -911
rect 548 -912 549 -858
rect 604 -927 605 -911
rect 128 -914 129 -858
rect 446 -927 447 -913
rect 128 -927 129 -915
rect 184 -927 185 -915
rect 215 -927 216 -915
rect 520 -927 521 -915
rect 170 -927 171 -917
rect 205 -927 206 -917
rect 219 -918 220 -858
rect 331 -918 332 -858
rect 380 -927 381 -917
rect 548 -927 549 -917
rect 219 -927 220 -919
rect 415 -927 416 -919
rect 275 -922 276 -858
rect 478 -927 479 -921
rect 303 -924 304 -858
rect 807 -927 808 -923
rect 19 -926 20 -858
rect 303 -927 304 -925
rect 331 -927 332 -925
rect 341 -927 342 -925
rect 2 -1006 3 -936
rect 233 -937 234 -935
rect 247 -937 248 -935
rect 261 -937 262 -935
rect 275 -1006 276 -936
rect 359 -937 360 -935
rect 390 -1006 391 -936
rect 723 -937 724 -935
rect 779 -937 780 -935
rect 898 -1006 899 -936
rect 9 -939 10 -935
rect 82 -939 83 -935
rect 100 -939 101 -935
rect 338 -939 339 -935
rect 348 -939 349 -935
rect 786 -939 787 -935
rect 814 -939 815 -935
rect 849 -1006 850 -938
rect 9 -1006 10 -940
rect 128 -941 129 -935
rect 149 -1006 150 -940
rect 170 -941 171 -935
rect 173 -1006 174 -940
rect 387 -941 388 -935
rect 394 -941 395 -935
rect 436 -941 437 -935
rect 450 -941 451 -935
rect 863 -1006 864 -940
rect 16 -943 17 -935
rect 334 -1006 335 -942
rect 352 -943 353 -935
rect 499 -943 500 -935
rect 509 -943 510 -935
rect 737 -943 738 -935
rect 786 -1006 787 -942
rect 828 -943 829 -935
rect 842 -943 843 -935
rect 842 -1006 843 -942
rect 842 -943 843 -935
rect 842 -1006 843 -942
rect 30 -945 31 -935
rect 296 -945 297 -935
rect 331 -945 332 -935
rect 359 -1006 360 -944
rect 397 -1006 398 -944
rect 674 -945 675 -935
rect 716 -945 717 -935
rect 779 -1006 780 -944
rect 814 -1006 815 -944
rect 835 -945 836 -935
rect 37 -1006 38 -946
rect 124 -947 125 -935
rect 128 -1006 129 -946
rect 222 -1006 223 -946
rect 247 -1006 248 -946
rect 313 -1006 314 -946
rect 331 -1006 332 -946
rect 702 -947 703 -935
rect 737 -1006 738 -946
rect 744 -947 745 -935
rect 40 -949 41 -935
rect 72 -949 73 -935
rect 79 -1006 80 -948
rect 380 -949 381 -935
rect 401 -949 402 -935
rect 667 -949 668 -935
rect 744 -1006 745 -948
rect 751 -949 752 -935
rect 44 -951 45 -935
rect 285 -951 286 -935
rect 404 -951 405 -935
rect 408 -951 409 -935
rect 429 -951 430 -935
rect 499 -1006 500 -950
rect 513 -951 514 -935
rect 660 -951 661 -935
rect 751 -1006 752 -950
rect 807 -951 808 -935
rect 51 -1006 52 -952
rect 93 -953 94 -935
rect 117 -1006 118 -952
rect 576 -953 577 -935
rect 590 -953 591 -935
rect 821 -953 822 -935
rect 58 -955 59 -935
rect 394 -1006 395 -954
rect 408 -1006 409 -954
rect 604 -955 605 -935
rect 646 -955 647 -935
rect 667 -1006 668 -954
rect 793 -955 794 -935
rect 807 -1006 808 -954
rect 58 -1006 59 -956
rect 93 -1006 94 -956
rect 121 -957 122 -935
rect 194 -1006 195 -956
rect 201 -957 202 -935
rect 282 -1006 283 -956
rect 303 -957 304 -935
rect 590 -1006 591 -956
rect 646 -1006 647 -956
rect 688 -957 689 -935
rect 44 -1006 45 -958
rect 121 -1006 122 -958
rect 152 -959 153 -935
rect 835 -1006 836 -958
rect 61 -1006 62 -960
rect 411 -1006 412 -960
rect 429 -1006 430 -960
rect 828 -1006 829 -960
rect 65 -963 66 -935
rect 86 -963 87 -935
rect 163 -1006 164 -962
rect 485 -963 486 -935
rect 516 -963 517 -935
rect 793 -1006 794 -962
rect 65 -1006 66 -964
rect 373 -965 374 -935
rect 436 -1006 437 -964
rect 632 -965 633 -935
rect 653 -965 654 -935
rect 702 -1006 703 -964
rect 72 -1006 73 -966
rect 156 -967 157 -935
rect 177 -967 178 -935
rect 303 -1006 304 -966
rect 373 -1006 374 -966
rect 380 -1006 381 -966
rect 443 -967 444 -935
rect 821 -1006 822 -966
rect 86 -1006 87 -968
rect 317 -969 318 -935
rect 443 -1006 444 -968
rect 457 -969 458 -935
rect 464 -1006 465 -968
rect 471 -969 472 -935
rect 474 -1006 475 -968
rect 723 -1006 724 -968
rect 135 -971 136 -935
rect 156 -1006 157 -970
rect 177 -1006 178 -970
rect 226 -971 227 -935
rect 254 -971 255 -935
rect 296 -1006 297 -970
rect 317 -1006 318 -970
rect 345 -971 346 -935
rect 446 -971 447 -935
rect 716 -1006 717 -970
rect 135 -1006 136 -972
rect 201 -1006 202 -972
rect 205 -1006 206 -972
rect 856 -1006 857 -972
rect 170 -1006 171 -974
rect 226 -1006 227 -974
rect 254 -1006 255 -974
rect 453 -975 454 -935
rect 457 -1006 458 -974
rect 492 -975 493 -935
rect 520 -975 521 -935
rect 520 -1006 521 -974
rect 520 -975 521 -935
rect 520 -1006 521 -974
rect 527 -975 528 -935
rect 527 -1006 528 -974
rect 527 -975 528 -935
rect 527 -1006 528 -974
rect 534 -975 535 -935
rect 534 -1006 535 -974
rect 534 -975 535 -935
rect 534 -1006 535 -974
rect 541 -975 542 -935
rect 618 -975 619 -935
rect 653 -1006 654 -974
rect 681 -975 682 -935
rect 688 -1006 689 -974
rect 695 -975 696 -935
rect 191 -977 192 -935
rect 233 -1006 234 -976
rect 261 -1006 262 -976
rect 268 -977 269 -935
rect 278 -977 279 -935
rect 422 -977 423 -935
rect 450 -1006 451 -976
rect 478 -977 479 -935
rect 481 -1006 482 -976
rect 541 -1006 542 -976
rect 548 -977 549 -935
rect 800 -977 801 -935
rect 208 -979 209 -935
rect 639 -979 640 -935
rect 695 -1006 696 -978
rect 730 -979 731 -935
rect 772 -979 773 -935
rect 800 -1006 801 -978
rect 212 -1006 213 -980
rect 387 -1006 388 -980
rect 478 -1006 479 -980
rect 660 -1006 661 -980
rect 765 -981 766 -935
rect 772 -1006 773 -980
rect 215 -983 216 -935
rect 310 -983 311 -935
rect 338 -1006 339 -982
rect 548 -1006 549 -982
rect 562 -983 563 -935
rect 618 -1006 619 -982
rect 639 -1006 640 -982
rect 709 -983 710 -935
rect 758 -983 759 -935
rect 765 -1006 766 -982
rect 184 -985 185 -935
rect 709 -1006 710 -984
rect 758 -1006 759 -984
rect 873 -1006 874 -984
rect 142 -987 143 -935
rect 184 -1006 185 -986
rect 219 -1006 220 -986
rect 240 -987 241 -935
rect 268 -1006 269 -986
rect 352 -1006 353 -986
rect 376 -1006 377 -986
rect 730 -1006 731 -986
rect 114 -989 115 -935
rect 142 -1006 143 -988
rect 240 -1006 241 -988
rect 415 -989 416 -935
rect 485 -1006 486 -988
rect 569 -989 570 -935
rect 576 -1006 577 -988
rect 597 -989 598 -935
rect 114 -1006 115 -990
rect 674 -1006 675 -990
rect 289 -993 290 -935
rect 632 -1006 633 -992
rect 289 -1006 290 -994
rect 324 -995 325 -935
rect 345 -1006 346 -994
rect 366 -995 367 -935
rect 404 -1006 405 -994
rect 415 -1006 416 -994
rect 555 -995 556 -935
rect 562 -1006 563 -994
rect 583 -995 584 -935
rect 681 -1006 682 -994
rect 23 -997 24 -935
rect 366 -1006 367 -996
rect 555 -1006 556 -996
rect 625 -997 626 -935
rect 23 -1006 24 -998
rect 107 -999 108 -935
rect 299 -999 300 -935
rect 492 -1006 493 -998
rect 558 -1006 559 -998
rect 569 -1006 570 -998
rect 597 -1006 598 -998
rect 859 -1006 860 -998
rect 107 -1006 108 -1000
rect 131 -1006 132 -1000
rect 324 -1006 325 -1000
rect 506 -1001 507 -935
rect 611 -1001 612 -935
rect 625 -1006 626 -1000
rect 425 -1006 426 -1002
rect 611 -1006 612 -1002
rect 506 -1006 507 -1004
rect 604 -1006 605 -1004
rect 2 -1016 3 -1014
rect 411 -1016 412 -1014
rect 422 -1083 423 -1015
rect 541 -1016 542 -1014
rect 551 -1083 552 -1015
rect 723 -1016 724 -1014
rect 786 -1016 787 -1014
rect 856 -1083 857 -1015
rect 863 -1016 864 -1014
rect 919 -1083 920 -1015
rect 9 -1018 10 -1014
rect 170 -1018 171 -1014
rect 212 -1018 213 -1014
rect 338 -1083 339 -1017
rect 341 -1018 342 -1014
rect 492 -1018 493 -1014
rect 502 -1018 503 -1014
rect 842 -1018 843 -1014
rect 849 -1018 850 -1014
rect 912 -1083 913 -1017
rect 16 -1083 17 -1019
rect 205 -1020 206 -1014
rect 212 -1083 213 -1019
rect 401 -1020 402 -1014
rect 404 -1020 405 -1014
rect 485 -1020 486 -1014
rect 492 -1083 493 -1019
rect 884 -1083 885 -1019
rect 898 -1020 899 -1014
rect 926 -1083 927 -1019
rect 19 -1022 20 -1014
rect 786 -1083 787 -1021
rect 793 -1022 794 -1014
rect 793 -1083 794 -1021
rect 793 -1022 794 -1014
rect 793 -1083 794 -1021
rect 800 -1022 801 -1014
rect 877 -1083 878 -1021
rect 23 -1024 24 -1014
rect 26 -1052 27 -1023
rect 30 -1083 31 -1023
rect 198 -1083 199 -1023
rect 205 -1083 206 -1023
rect 261 -1024 262 -1014
rect 303 -1024 304 -1014
rect 467 -1083 468 -1023
rect 478 -1024 479 -1014
rect 639 -1024 640 -1014
rect 642 -1083 643 -1023
rect 842 -1083 843 -1023
rect 23 -1083 24 -1025
rect 166 -1083 167 -1025
rect 233 -1026 234 -1014
rect 261 -1083 262 -1025
rect 558 -1083 559 -1025
rect 590 -1026 591 -1014
rect 891 -1083 892 -1025
rect 33 -1028 34 -1014
rect 709 -1028 710 -1014
rect 772 -1028 773 -1014
rect 800 -1083 801 -1027
rect 807 -1028 808 -1014
rect 870 -1083 871 -1027
rect 37 -1030 38 -1014
rect 191 -1030 192 -1014
rect 219 -1030 220 -1014
rect 282 -1030 283 -1014
rect 303 -1083 304 -1029
rect 324 -1030 325 -1014
rect 331 -1030 332 -1014
rect 730 -1030 731 -1014
rect 772 -1083 773 -1029
rect 859 -1030 860 -1014
rect 37 -1083 38 -1031
rect 86 -1032 87 -1014
rect 93 -1032 94 -1014
rect 436 -1083 437 -1031
rect 439 -1032 440 -1014
rect 478 -1083 479 -1031
rect 506 -1032 507 -1014
rect 611 -1032 612 -1014
rect 618 -1032 619 -1014
rect 618 -1083 619 -1031
rect 618 -1032 619 -1014
rect 618 -1083 619 -1031
rect 660 -1032 661 -1014
rect 723 -1083 724 -1031
rect 779 -1032 780 -1014
rect 849 -1083 850 -1031
rect 54 -1083 55 -1033
rect 86 -1083 87 -1033
rect 107 -1034 108 -1014
rect 408 -1083 409 -1033
rect 415 -1034 416 -1014
rect 485 -1083 486 -1033
rect 513 -1034 514 -1014
rect 751 -1034 752 -1014
rect 821 -1034 822 -1014
rect 940 -1083 941 -1033
rect 58 -1083 59 -1035
rect 159 -1083 160 -1035
rect 163 -1036 164 -1014
rect 513 -1083 514 -1035
rect 516 -1036 517 -1014
rect 597 -1036 598 -1014
rect 604 -1036 605 -1014
rect 614 -1036 615 -1014
rect 681 -1036 682 -1014
rect 730 -1083 731 -1035
rect 828 -1036 829 -1014
rect 898 -1083 899 -1035
rect 65 -1038 66 -1014
rect 415 -1083 416 -1037
rect 432 -1038 433 -1014
rect 443 -1038 444 -1014
rect 446 -1083 447 -1037
rect 807 -1083 808 -1037
rect 835 -1038 836 -1014
rect 905 -1083 906 -1037
rect 65 -1083 66 -1039
rect 254 -1040 255 -1014
rect 278 -1083 279 -1039
rect 282 -1083 283 -1039
rect 289 -1040 290 -1014
rect 506 -1083 507 -1039
rect 527 -1040 528 -1014
rect 590 -1083 591 -1039
rect 604 -1083 605 -1039
rect 744 -1040 745 -1014
rect 72 -1042 73 -1014
rect 114 -1042 115 -1014
rect 121 -1083 122 -1041
rect 142 -1042 143 -1014
rect 163 -1083 164 -1041
rect 814 -1042 815 -1014
rect 72 -1083 73 -1043
rect 149 -1044 150 -1014
rect 152 -1083 153 -1043
rect 814 -1083 815 -1043
rect 79 -1046 80 -1014
rect 310 -1083 311 -1045
rect 317 -1046 318 -1014
rect 401 -1083 402 -1045
rect 453 -1083 454 -1045
rect 572 -1083 573 -1045
rect 576 -1046 577 -1014
rect 660 -1083 661 -1045
rect 674 -1046 675 -1014
rect 744 -1083 745 -1045
rect 79 -1083 80 -1047
rect 275 -1048 276 -1014
rect 296 -1048 297 -1014
rect 324 -1083 325 -1047
rect 352 -1048 353 -1014
rect 394 -1083 395 -1047
rect 499 -1048 500 -1014
rect 828 -1083 829 -1047
rect 103 -1083 104 -1049
rect 114 -1083 115 -1049
rect 128 -1050 129 -1014
rect 667 -1050 668 -1014
rect 688 -1050 689 -1014
rect 821 -1083 822 -1049
rect 107 -1083 108 -1051
rect 117 -1052 118 -1014
rect 128 -1083 129 -1051
rect 334 -1052 335 -1014
rect 352 -1083 353 -1051
rect 583 -1083 584 -1051
rect 614 -1083 615 -1051
rect 674 -1083 675 -1051
rect 695 -1052 696 -1014
rect 863 -1083 864 -1051
rect 135 -1054 136 -1014
rect 142 -1083 143 -1053
rect 170 -1083 171 -1053
rect 268 -1054 269 -1014
rect 275 -1083 276 -1053
rect 450 -1054 451 -1014
rect 464 -1054 465 -1014
rect 499 -1083 500 -1053
rect 520 -1054 521 -1014
rect 576 -1083 577 -1053
rect 702 -1054 703 -1014
rect 702 -1083 703 -1053
rect 702 -1054 703 -1014
rect 702 -1083 703 -1053
rect 716 -1054 717 -1014
rect 779 -1083 780 -1053
rect 177 -1056 178 -1014
rect 233 -1083 234 -1055
rect 243 -1083 244 -1055
rect 289 -1083 290 -1055
rect 317 -1083 318 -1055
rect 495 -1083 496 -1055
rect 527 -1083 528 -1055
rect 681 -1083 682 -1055
rect 737 -1056 738 -1014
rect 835 -1083 836 -1055
rect 100 -1058 101 -1014
rect 177 -1083 178 -1057
rect 184 -1058 185 -1014
rect 254 -1083 255 -1057
rect 268 -1083 269 -1057
rect 348 -1083 349 -1057
rect 359 -1058 360 -1014
rect 373 -1083 374 -1057
rect 380 -1058 381 -1014
rect 390 -1058 391 -1014
rect 429 -1058 430 -1014
rect 520 -1083 521 -1057
rect 534 -1058 535 -1014
rect 695 -1083 696 -1057
rect 191 -1083 192 -1059
rect 222 -1060 223 -1014
rect 226 -1060 227 -1014
rect 541 -1083 542 -1059
rect 565 -1083 566 -1059
rect 667 -1083 668 -1059
rect 44 -1062 45 -1014
rect 222 -1083 223 -1061
rect 226 -1083 227 -1061
rect 240 -1062 241 -1014
rect 247 -1062 248 -1014
rect 296 -1083 297 -1061
rect 345 -1062 346 -1014
rect 380 -1083 381 -1061
rect 387 -1083 388 -1061
rect 632 -1062 633 -1014
rect 646 -1062 647 -1014
rect 737 -1083 738 -1061
rect 44 -1083 45 -1063
rect 51 -1064 52 -1014
rect 201 -1064 202 -1014
rect 331 -1083 332 -1063
rect 345 -1083 346 -1063
rect 758 -1064 759 -1014
rect 359 -1083 360 -1065
rect 537 -1083 538 -1065
rect 548 -1066 549 -1014
rect 632 -1083 633 -1065
rect 653 -1066 654 -1014
rect 716 -1083 717 -1065
rect 758 -1083 759 -1065
rect 765 -1066 766 -1014
rect 184 -1083 185 -1067
rect 548 -1083 549 -1067
rect 562 -1068 563 -1014
rect 646 -1083 647 -1067
rect 366 -1070 367 -1014
rect 611 -1083 612 -1069
rect 625 -1070 626 -1014
rect 765 -1083 766 -1069
rect 366 -1083 367 -1071
rect 530 -1083 531 -1071
rect 534 -1083 535 -1071
rect 751 -1083 752 -1071
rect 376 -1074 377 -1014
rect 653 -1083 654 -1073
rect 390 -1083 391 -1075
rect 471 -1083 472 -1075
rect 562 -1083 563 -1075
rect 709 -1083 710 -1075
rect 429 -1083 430 -1077
rect 457 -1078 458 -1014
rect 569 -1078 570 -1014
rect 597 -1083 598 -1077
rect 607 -1083 608 -1077
rect 625 -1083 626 -1077
rect 194 -1080 195 -1014
rect 457 -1083 458 -1079
rect 450 -1083 451 -1081
rect 688 -1083 689 -1081
rect 9 -1093 10 -1091
rect 786 -1093 787 -1091
rect 807 -1093 808 -1091
rect 807 -1180 808 -1092
rect 807 -1093 808 -1091
rect 807 -1180 808 -1092
rect 884 -1093 885 -1091
rect 975 -1180 976 -1092
rect 982 -1180 983 -1092
rect 989 -1180 990 -1092
rect 9 -1180 10 -1094
rect 170 -1095 171 -1091
rect 198 -1095 199 -1091
rect 226 -1095 227 -1091
rect 240 -1180 241 -1094
rect 282 -1095 283 -1091
rect 317 -1095 318 -1091
rect 443 -1180 444 -1094
rect 446 -1095 447 -1091
rect 891 -1095 892 -1091
rect 898 -1095 899 -1091
rect 968 -1180 969 -1094
rect 16 -1097 17 -1091
rect 579 -1180 580 -1096
rect 642 -1097 643 -1091
rect 849 -1097 850 -1091
rect 856 -1097 857 -1091
rect 898 -1180 899 -1096
rect 912 -1097 913 -1091
rect 947 -1180 948 -1096
rect 16 -1180 17 -1098
rect 30 -1099 31 -1091
rect 44 -1099 45 -1091
rect 96 -1099 97 -1091
rect 103 -1099 104 -1091
rect 716 -1099 717 -1091
rect 828 -1099 829 -1091
rect 884 -1180 885 -1098
rect 940 -1099 941 -1091
rect 940 -1180 941 -1098
rect 940 -1099 941 -1091
rect 940 -1180 941 -1098
rect 30 -1180 31 -1100
rect 37 -1101 38 -1091
rect 44 -1180 45 -1100
rect 205 -1101 206 -1091
rect 226 -1180 227 -1100
rect 310 -1101 311 -1091
rect 345 -1180 346 -1100
rect 366 -1101 367 -1091
rect 387 -1180 388 -1100
rect 408 -1101 409 -1091
rect 436 -1101 437 -1091
rect 439 -1113 440 -1100
rect 450 -1101 451 -1091
rect 639 -1101 640 -1091
rect 667 -1101 668 -1091
rect 933 -1180 934 -1100
rect 37 -1180 38 -1102
rect 268 -1103 269 -1091
rect 275 -1180 276 -1102
rect 320 -1180 321 -1102
rect 348 -1103 349 -1091
rect 415 -1103 416 -1091
rect 436 -1180 437 -1102
rect 492 -1103 493 -1091
rect 506 -1103 507 -1091
rect 534 -1180 535 -1102
rect 544 -1180 545 -1102
rect 821 -1103 822 -1091
rect 842 -1103 843 -1091
rect 891 -1180 892 -1102
rect 51 -1180 52 -1104
rect 86 -1105 87 -1091
rect 93 -1105 94 -1091
rect 912 -1180 913 -1104
rect 58 -1107 59 -1091
rect 65 -1180 66 -1106
rect 72 -1107 73 -1091
rect 152 -1107 153 -1091
rect 156 -1180 157 -1106
rect 177 -1107 178 -1091
rect 198 -1180 199 -1106
rect 555 -1180 556 -1106
rect 558 -1107 559 -1091
rect 863 -1107 864 -1091
rect 58 -1180 59 -1108
rect 254 -1109 255 -1091
rect 268 -1180 269 -1108
rect 296 -1109 297 -1091
rect 303 -1109 304 -1091
rect 310 -1180 311 -1108
rect 355 -1109 356 -1091
rect 695 -1109 696 -1091
rect 702 -1109 703 -1091
rect 856 -1180 857 -1108
rect 863 -1180 864 -1108
rect 929 -1109 930 -1091
rect 72 -1180 73 -1110
rect 201 -1180 202 -1110
rect 205 -1180 206 -1110
rect 362 -1180 363 -1110
rect 366 -1180 367 -1110
rect 632 -1111 633 -1091
rect 684 -1180 685 -1110
rect 877 -1111 878 -1091
rect 82 -1113 83 -1091
rect 219 -1113 220 -1091
rect 247 -1180 248 -1112
rect 289 -1113 290 -1091
rect 303 -1180 304 -1112
rect 324 -1113 325 -1091
rect 355 -1180 356 -1112
rect 415 -1180 416 -1112
rect 492 -1180 493 -1112
rect 520 -1113 521 -1091
rect 604 -1113 605 -1091
rect 607 -1113 608 -1091
rect 667 -1180 668 -1112
rect 702 -1180 703 -1112
rect 716 -1180 717 -1112
rect 751 -1113 752 -1091
rect 842 -1180 843 -1112
rect 849 -1180 850 -1112
rect 961 -1180 962 -1112
rect 86 -1180 87 -1114
rect 107 -1115 108 -1091
rect 128 -1115 129 -1091
rect 296 -1180 297 -1114
rect 331 -1115 332 -1091
rect 604 -1180 605 -1114
rect 758 -1115 759 -1091
rect 821 -1180 822 -1114
rect 103 -1180 104 -1116
rect 254 -1180 255 -1116
rect 278 -1117 279 -1091
rect 751 -1180 752 -1116
rect 800 -1117 801 -1091
rect 828 -1180 829 -1116
rect 107 -1180 108 -1118
rect 114 -1119 115 -1091
rect 128 -1180 129 -1118
rect 142 -1119 143 -1091
rect 152 -1180 153 -1118
rect 506 -1180 507 -1118
rect 527 -1119 528 -1091
rect 737 -1119 738 -1091
rect 114 -1180 115 -1120
rect 380 -1121 381 -1091
rect 390 -1121 391 -1091
rect 919 -1121 920 -1091
rect 135 -1123 136 -1091
rect 786 -1180 787 -1122
rect 870 -1123 871 -1091
rect 919 -1180 920 -1122
rect 135 -1180 136 -1124
rect 520 -1180 521 -1124
rect 530 -1125 531 -1091
rect 905 -1125 906 -1091
rect 138 -1127 139 -1091
rect 233 -1127 234 -1091
rect 250 -1127 251 -1091
rect 695 -1180 696 -1126
rect 772 -1127 773 -1091
rect 870 -1180 871 -1126
rect 23 -1129 24 -1091
rect 233 -1180 234 -1128
rect 282 -1180 283 -1128
rect 527 -1180 528 -1128
rect 562 -1129 563 -1091
rect 814 -1129 815 -1091
rect 93 -1180 94 -1130
rect 772 -1180 773 -1130
rect 793 -1131 794 -1091
rect 905 -1180 906 -1130
rect 142 -1180 143 -1132
rect 429 -1133 430 -1091
rect 453 -1133 454 -1091
rect 688 -1133 689 -1091
rect 709 -1133 710 -1091
rect 814 -1180 815 -1132
rect 163 -1180 164 -1134
rect 261 -1135 262 -1091
rect 289 -1180 290 -1134
rect 359 -1135 360 -1091
rect 380 -1180 381 -1134
rect 394 -1135 395 -1091
rect 422 -1135 423 -1091
rect 688 -1180 689 -1134
rect 166 -1137 167 -1091
rect 877 -1180 878 -1136
rect 177 -1180 178 -1138
rect 191 -1139 192 -1091
rect 261 -1180 262 -1138
rect 485 -1139 486 -1091
rect 562 -1180 563 -1138
rect 926 -1139 927 -1091
rect 184 -1141 185 -1091
rect 429 -1180 430 -1140
rect 464 -1141 465 -1091
rect 835 -1141 836 -1091
rect 170 -1180 171 -1142
rect 184 -1180 185 -1142
rect 191 -1180 192 -1142
rect 212 -1143 213 -1091
rect 324 -1180 325 -1142
rect 453 -1180 454 -1142
rect 485 -1180 486 -1142
rect 509 -1180 510 -1142
rect 569 -1143 570 -1091
rect 800 -1180 801 -1142
rect 331 -1180 332 -1144
rect 590 -1145 591 -1091
rect 618 -1145 619 -1091
rect 758 -1180 759 -1144
rect 338 -1147 339 -1091
rect 422 -1180 423 -1146
rect 513 -1147 514 -1091
rect 569 -1180 570 -1146
rect 572 -1147 573 -1091
rect 765 -1147 766 -1091
rect 222 -1149 223 -1091
rect 765 -1180 766 -1148
rect 222 -1180 223 -1150
rect 394 -1180 395 -1150
rect 401 -1151 402 -1091
rect 513 -1180 514 -1150
rect 576 -1151 577 -1091
rect 632 -1180 633 -1150
rect 646 -1151 647 -1091
rect 709 -1180 710 -1150
rect 730 -1151 731 -1091
rect 835 -1180 836 -1150
rect 338 -1180 339 -1152
rect 373 -1153 374 -1091
rect 583 -1153 584 -1091
rect 639 -1180 640 -1152
rect 646 -1180 647 -1152
rect 681 -1153 682 -1091
rect 359 -1180 360 -1154
rect 779 -1155 780 -1091
rect 373 -1180 374 -1156
rect 450 -1180 451 -1156
rect 548 -1180 549 -1156
rect 681 -1180 682 -1156
rect 744 -1157 745 -1091
rect 779 -1180 780 -1156
rect 79 -1159 80 -1091
rect 744 -1180 745 -1158
rect 79 -1180 80 -1160
rect 121 -1161 122 -1091
rect 425 -1180 426 -1160
rect 583 -1180 584 -1160
rect 618 -1180 619 -1160
rect 723 -1161 724 -1091
rect 625 -1163 626 -1091
rect 793 -1180 794 -1162
rect 611 -1165 612 -1091
rect 625 -1180 626 -1164
rect 653 -1165 654 -1091
rect 723 -1180 724 -1164
rect 597 -1167 598 -1091
rect 611 -1180 612 -1166
rect 656 -1180 657 -1166
rect 926 -1180 927 -1166
rect 499 -1169 500 -1091
rect 597 -1180 598 -1168
rect 660 -1169 661 -1091
rect 730 -1180 731 -1168
rect 478 -1171 479 -1091
rect 499 -1180 500 -1170
rect 541 -1171 542 -1091
rect 660 -1180 661 -1170
rect 674 -1171 675 -1091
rect 737 -1180 738 -1170
rect 401 -1180 402 -1172
rect 478 -1180 479 -1172
rect 541 -1180 542 -1172
rect 590 -1180 591 -1172
rect 457 -1175 458 -1091
rect 674 -1180 675 -1174
rect 457 -1180 458 -1176
rect 471 -1177 472 -1091
rect 212 -1180 213 -1178
rect 471 -1180 472 -1178
rect 5 -1190 6 -1188
rect 219 -1190 220 -1188
rect 222 -1190 223 -1188
rect 674 -1190 675 -1188
rect 719 -1190 720 -1188
rect 828 -1190 829 -1188
rect 940 -1190 941 -1188
rect 964 -1190 965 -1188
rect 975 -1190 976 -1188
rect 982 -1275 983 -1189
rect 985 -1190 986 -1188
rect 1010 -1275 1011 -1189
rect 9 -1192 10 -1188
rect 212 -1192 213 -1188
rect 215 -1192 216 -1188
rect 723 -1192 724 -1188
rect 737 -1192 738 -1188
rect 740 -1216 741 -1191
rect 751 -1192 752 -1188
rect 954 -1275 955 -1191
rect 989 -1192 990 -1188
rect 1003 -1275 1004 -1191
rect 16 -1194 17 -1188
rect 215 -1275 216 -1193
rect 247 -1194 248 -1188
rect 247 -1275 248 -1193
rect 247 -1194 248 -1188
rect 247 -1275 248 -1193
rect 254 -1194 255 -1188
rect 306 -1275 307 -1193
rect 341 -1275 342 -1193
rect 618 -1275 619 -1193
rect 625 -1194 626 -1188
rect 716 -1275 717 -1193
rect 723 -1275 724 -1193
rect 744 -1194 745 -1188
rect 800 -1194 801 -1188
rect 828 -1275 829 -1193
rect 968 -1194 969 -1188
rect 989 -1275 990 -1193
rect 16 -1275 17 -1195
rect 177 -1196 178 -1188
rect 201 -1196 202 -1188
rect 765 -1196 766 -1188
rect 800 -1275 801 -1195
rect 884 -1196 885 -1188
rect 912 -1196 913 -1188
rect 968 -1275 969 -1195
rect 26 -1198 27 -1188
rect 26 -1275 27 -1197
rect 26 -1198 27 -1188
rect 26 -1275 27 -1197
rect 44 -1198 45 -1188
rect 313 -1275 314 -1197
rect 352 -1275 353 -1197
rect 485 -1198 486 -1188
rect 506 -1198 507 -1188
rect 898 -1198 899 -1188
rect 58 -1200 59 -1188
rect 173 -1200 174 -1188
rect 254 -1275 255 -1199
rect 362 -1275 363 -1199
rect 373 -1200 374 -1188
rect 422 -1275 423 -1199
rect 429 -1200 430 -1188
rect 765 -1275 766 -1199
rect 814 -1200 815 -1188
rect 996 -1275 997 -1199
rect 58 -1275 59 -1201
rect 460 -1275 461 -1201
rect 464 -1202 465 -1188
rect 793 -1202 794 -1188
rect 814 -1275 815 -1201
rect 926 -1202 927 -1188
rect 72 -1275 73 -1203
rect 198 -1204 199 -1188
rect 268 -1204 269 -1188
rect 317 -1275 318 -1203
rect 355 -1204 356 -1188
rect 366 -1204 367 -1188
rect 411 -1204 412 -1188
rect 688 -1204 689 -1188
rect 737 -1275 738 -1203
rect 856 -1204 857 -1188
rect 65 -1206 66 -1188
rect 366 -1275 367 -1205
rect 411 -1275 412 -1205
rect 681 -1275 682 -1205
rect 842 -1206 843 -1188
rect 856 -1275 857 -1205
rect 65 -1275 66 -1207
rect 499 -1208 500 -1188
rect 534 -1208 535 -1188
rect 688 -1275 689 -1207
rect 786 -1208 787 -1188
rect 842 -1275 843 -1207
rect 849 -1208 850 -1188
rect 912 -1275 913 -1207
rect 86 -1210 87 -1188
rect 121 -1210 122 -1188
rect 135 -1210 136 -1188
rect 226 -1210 227 -1188
rect 268 -1275 269 -1209
rect 303 -1210 304 -1188
rect 310 -1210 311 -1188
rect 373 -1275 374 -1209
rect 429 -1275 430 -1209
rect 562 -1210 563 -1188
rect 579 -1210 580 -1188
rect 975 -1275 976 -1209
rect 79 -1212 80 -1188
rect 135 -1275 136 -1211
rect 142 -1212 143 -1188
rect 320 -1212 321 -1188
rect 359 -1275 360 -1211
rect 807 -1212 808 -1188
rect 30 -1214 31 -1188
rect 142 -1275 143 -1213
rect 149 -1214 150 -1188
rect 331 -1214 332 -1188
rect 446 -1275 447 -1213
rect 709 -1214 710 -1188
rect 772 -1214 773 -1188
rect 786 -1275 787 -1213
rect 30 -1275 31 -1215
rect 408 -1216 409 -1188
rect 450 -1216 451 -1188
rect 597 -1216 598 -1188
rect 604 -1216 605 -1188
rect 674 -1275 675 -1215
rect 772 -1275 773 -1215
rect 779 -1216 780 -1188
rect 849 -1275 850 -1215
rect 12 -1275 13 -1217
rect 408 -1275 409 -1217
rect 436 -1218 437 -1188
rect 450 -1275 451 -1217
rect 453 -1218 454 -1188
rect 758 -1218 759 -1188
rect 79 -1275 80 -1219
rect 324 -1220 325 -1188
rect 464 -1275 465 -1219
rect 933 -1220 934 -1188
rect 86 -1275 87 -1221
rect 152 -1222 153 -1188
rect 163 -1222 164 -1188
rect 198 -1275 199 -1221
rect 226 -1275 227 -1221
rect 495 -1275 496 -1221
rect 520 -1222 521 -1188
rect 562 -1275 563 -1221
rect 583 -1222 584 -1188
rect 926 -1275 927 -1221
rect 93 -1224 94 -1188
rect 205 -1224 206 -1188
rect 233 -1224 234 -1188
rect 324 -1275 325 -1223
rect 467 -1224 468 -1188
rect 653 -1275 654 -1223
rect 656 -1224 657 -1188
rect 905 -1224 906 -1188
rect 37 -1226 38 -1188
rect 205 -1275 206 -1225
rect 233 -1275 234 -1225
rect 401 -1226 402 -1188
rect 474 -1275 475 -1225
rect 520 -1275 521 -1225
rect 527 -1226 528 -1188
rect 534 -1275 535 -1225
rect 541 -1226 542 -1188
rect 957 -1226 958 -1188
rect 93 -1275 94 -1227
rect 632 -1228 633 -1188
rect 635 -1275 636 -1227
rect 807 -1275 808 -1227
rect 877 -1228 878 -1188
rect 933 -1275 934 -1227
rect 96 -1230 97 -1188
rect 163 -1275 164 -1229
rect 170 -1275 171 -1229
rect 177 -1275 178 -1229
rect 275 -1230 276 -1188
rect 744 -1275 745 -1229
rect 758 -1275 759 -1229
rect 870 -1230 871 -1188
rect 877 -1275 878 -1229
rect 947 -1230 948 -1188
rect 96 -1275 97 -1231
rect 331 -1275 332 -1231
rect 401 -1275 402 -1231
rect 467 -1275 468 -1231
rect 471 -1232 472 -1188
rect 541 -1275 542 -1231
rect 544 -1232 545 -1188
rect 898 -1275 899 -1231
rect 100 -1275 101 -1233
rect 156 -1234 157 -1188
rect 285 -1234 286 -1188
rect 492 -1234 493 -1188
rect 555 -1234 556 -1188
rect 625 -1275 626 -1233
rect 639 -1234 640 -1188
rect 709 -1275 710 -1233
rect 863 -1234 864 -1188
rect 870 -1275 871 -1233
rect 103 -1236 104 -1188
rect 695 -1236 696 -1188
rect 107 -1238 108 -1188
rect 121 -1275 122 -1237
rect 128 -1238 129 -1188
rect 156 -1275 157 -1237
rect 296 -1238 297 -1188
rect 436 -1275 437 -1237
rect 457 -1238 458 -1188
rect 527 -1275 528 -1237
rect 583 -1275 584 -1237
rect 590 -1238 591 -1188
rect 597 -1275 598 -1237
rect 695 -1275 696 -1237
rect 44 -1275 45 -1239
rect 128 -1275 129 -1239
rect 149 -1275 150 -1239
rect 184 -1240 185 -1188
rect 296 -1275 297 -1239
rect 345 -1240 346 -1188
rect 394 -1240 395 -1188
rect 639 -1275 640 -1239
rect 646 -1240 647 -1188
rect 793 -1275 794 -1239
rect 110 -1275 111 -1241
rect 191 -1242 192 -1188
rect 303 -1275 304 -1241
rect 425 -1242 426 -1188
rect 457 -1275 458 -1241
rect 730 -1242 731 -1188
rect 114 -1244 115 -1188
rect 576 -1275 577 -1243
rect 604 -1275 605 -1243
rect 751 -1275 752 -1243
rect 51 -1246 52 -1188
rect 114 -1275 115 -1245
rect 184 -1275 185 -1245
rect 275 -1275 276 -1245
rect 338 -1246 339 -1188
rect 394 -1275 395 -1245
rect 471 -1275 472 -1245
rect 961 -1246 962 -1188
rect 51 -1275 52 -1247
rect 261 -1248 262 -1188
rect 345 -1275 346 -1247
rect 380 -1248 381 -1188
rect 478 -1248 479 -1188
rect 905 -1275 906 -1247
rect 191 -1275 192 -1249
rect 222 -1275 223 -1249
rect 261 -1275 262 -1249
rect 289 -1250 290 -1188
rect 380 -1275 381 -1249
rect 590 -1275 591 -1249
rect 607 -1275 608 -1249
rect 821 -1250 822 -1188
rect 891 -1250 892 -1188
rect 961 -1275 962 -1249
rect 212 -1275 213 -1251
rect 730 -1275 731 -1251
rect 835 -1252 836 -1188
rect 891 -1275 892 -1251
rect 289 -1275 290 -1253
rect 387 -1254 388 -1188
rect 443 -1254 444 -1188
rect 478 -1275 479 -1253
rect 492 -1275 493 -1253
rect 779 -1275 780 -1253
rect 310 -1275 311 -1255
rect 835 -1275 836 -1255
rect 387 -1275 388 -1257
rect 415 -1258 416 -1188
rect 443 -1275 444 -1257
rect 485 -1275 486 -1257
rect 513 -1258 514 -1188
rect 555 -1275 556 -1257
rect 600 -1275 601 -1257
rect 821 -1275 822 -1257
rect 282 -1260 283 -1188
rect 415 -1275 416 -1259
rect 513 -1275 514 -1259
rect 548 -1260 549 -1188
rect 611 -1260 612 -1188
rect 611 -1275 612 -1259
rect 611 -1260 612 -1188
rect 611 -1275 612 -1259
rect 646 -1275 647 -1259
rect 943 -1275 944 -1259
rect 240 -1262 241 -1188
rect 282 -1275 283 -1261
rect 548 -1275 549 -1261
rect 569 -1262 570 -1188
rect 656 -1275 657 -1261
rect 919 -1262 920 -1188
rect 40 -1275 41 -1263
rect 240 -1275 241 -1263
rect 569 -1275 570 -1263
rect 919 -1275 920 -1263
rect 660 -1266 661 -1188
rect 863 -1275 864 -1265
rect 660 -1275 661 -1267
rect 702 -1268 703 -1188
rect 124 -1270 125 -1188
rect 702 -1275 703 -1269
rect 667 -1272 668 -1188
rect 884 -1275 885 -1271
rect 670 -1275 671 -1273
rect 947 -1275 948 -1273
rect 9 -1360 10 -1284
rect 30 -1285 31 -1283
rect 37 -1360 38 -1284
rect 149 -1285 150 -1283
rect 170 -1360 171 -1284
rect 219 -1285 220 -1283
rect 222 -1285 223 -1283
rect 289 -1285 290 -1283
rect 310 -1285 311 -1283
rect 576 -1285 577 -1283
rect 579 -1360 580 -1284
rect 926 -1285 927 -1283
rect 943 -1285 944 -1283
rect 1010 -1285 1011 -1283
rect 30 -1360 31 -1286
rect 688 -1287 689 -1283
rect 723 -1287 724 -1283
rect 723 -1360 724 -1286
rect 723 -1287 724 -1283
rect 723 -1360 724 -1286
rect 772 -1287 773 -1283
rect 772 -1360 773 -1286
rect 772 -1287 773 -1283
rect 772 -1360 773 -1286
rect 971 -1360 972 -1286
rect 989 -1287 990 -1283
rect 44 -1289 45 -1283
rect 215 -1360 216 -1288
rect 226 -1289 227 -1283
rect 506 -1289 507 -1283
rect 509 -1289 510 -1283
rect 695 -1289 696 -1283
rect 940 -1360 941 -1288
rect 989 -1360 990 -1288
rect 44 -1360 45 -1290
rect 86 -1291 87 -1283
rect 89 -1360 90 -1290
rect 453 -1360 454 -1290
rect 457 -1360 458 -1290
rect 541 -1291 542 -1283
rect 569 -1291 570 -1283
rect 954 -1291 955 -1283
rect 51 -1293 52 -1283
rect 341 -1293 342 -1283
rect 408 -1293 409 -1283
rect 436 -1293 437 -1283
rect 446 -1293 447 -1283
rect 492 -1360 493 -1292
rect 499 -1293 500 -1283
rect 709 -1293 710 -1283
rect 954 -1360 955 -1292
rect 1003 -1293 1004 -1283
rect 51 -1360 52 -1294
rect 96 -1295 97 -1283
rect 124 -1360 125 -1294
rect 226 -1360 227 -1294
rect 240 -1295 241 -1283
rect 289 -1360 290 -1294
rect 310 -1360 311 -1294
rect 317 -1295 318 -1283
rect 352 -1295 353 -1283
rect 499 -1360 500 -1294
rect 569 -1360 570 -1294
rect 583 -1295 584 -1283
rect 597 -1360 598 -1294
rect 611 -1295 612 -1283
rect 618 -1295 619 -1283
rect 919 -1295 920 -1283
rect 58 -1297 59 -1283
rect 173 -1297 174 -1283
rect 184 -1297 185 -1283
rect 863 -1297 864 -1283
rect 919 -1360 920 -1296
rect 975 -1297 976 -1283
rect 61 -1360 62 -1298
rect 107 -1360 108 -1298
rect 135 -1299 136 -1283
rect 184 -1360 185 -1298
rect 198 -1299 199 -1283
rect 219 -1360 220 -1298
rect 229 -1360 230 -1298
rect 863 -1360 864 -1298
rect 65 -1301 66 -1283
rect 352 -1360 353 -1300
rect 387 -1301 388 -1283
rect 408 -1360 409 -1300
rect 411 -1301 412 -1283
rect 898 -1301 899 -1283
rect 65 -1360 66 -1302
rect 380 -1303 381 -1283
rect 387 -1360 388 -1302
rect 555 -1303 556 -1283
rect 576 -1360 577 -1302
rect 912 -1303 913 -1283
rect 72 -1305 73 -1283
rect 128 -1305 129 -1283
rect 149 -1360 150 -1304
rect 261 -1305 262 -1283
rect 282 -1305 283 -1283
rect 359 -1305 360 -1283
rect 415 -1305 416 -1283
rect 464 -1305 465 -1283
rect 467 -1360 468 -1304
rect 488 -1360 489 -1304
rect 502 -1305 503 -1283
rect 583 -1360 584 -1304
rect 632 -1360 633 -1304
rect 660 -1305 661 -1283
rect 667 -1305 668 -1283
rect 891 -1305 892 -1283
rect 898 -1360 899 -1304
rect 982 -1305 983 -1283
rect 16 -1307 17 -1283
rect 261 -1360 262 -1306
rect 296 -1307 297 -1283
rect 359 -1360 360 -1306
rect 366 -1307 367 -1283
rect 464 -1360 465 -1306
rect 471 -1307 472 -1283
rect 793 -1307 794 -1283
rect 16 -1360 17 -1308
rect 110 -1309 111 -1283
rect 114 -1309 115 -1283
rect 135 -1360 136 -1308
rect 163 -1309 164 -1283
rect 282 -1360 283 -1308
rect 303 -1309 304 -1283
rect 471 -1360 472 -1308
rect 474 -1309 475 -1283
rect 646 -1309 647 -1283
rect 653 -1309 654 -1283
rect 891 -1360 892 -1308
rect 72 -1360 73 -1310
rect 730 -1311 731 -1283
rect 793 -1360 794 -1310
rect 849 -1311 850 -1283
rect 12 -1360 13 -1312
rect 730 -1360 731 -1312
rect 93 -1360 94 -1314
rect 530 -1360 531 -1314
rect 548 -1315 549 -1283
rect 611 -1360 612 -1314
rect 646 -1360 647 -1314
rect 716 -1315 717 -1283
rect 114 -1360 115 -1316
rect 121 -1317 122 -1283
rect 128 -1360 129 -1316
rect 254 -1317 255 -1283
rect 317 -1360 318 -1316
rect 324 -1317 325 -1283
rect 331 -1317 332 -1283
rect 618 -1360 619 -1316
rect 653 -1360 654 -1316
rect 702 -1317 703 -1283
rect 709 -1360 710 -1316
rect 835 -1317 836 -1283
rect 121 -1360 122 -1318
rect 625 -1319 626 -1283
rect 656 -1319 657 -1283
rect 996 -1319 997 -1283
rect 156 -1321 157 -1283
rect 163 -1360 164 -1320
rect 177 -1321 178 -1283
rect 324 -1360 325 -1320
rect 415 -1360 416 -1320
rect 943 -1360 944 -1320
rect 142 -1323 143 -1283
rect 177 -1360 178 -1322
rect 191 -1323 192 -1283
rect 198 -1360 199 -1322
rect 208 -1360 209 -1322
rect 506 -1360 507 -1322
rect 534 -1323 535 -1283
rect 548 -1360 549 -1322
rect 590 -1323 591 -1283
rect 660 -1360 661 -1322
rect 667 -1360 668 -1322
rect 807 -1323 808 -1283
rect 835 -1360 836 -1322
rect 933 -1323 934 -1283
rect 100 -1325 101 -1283
rect 191 -1360 192 -1324
rect 212 -1360 213 -1324
rect 296 -1360 297 -1324
rect 313 -1325 314 -1283
rect 590 -1360 591 -1324
rect 625 -1360 626 -1324
rect 681 -1325 682 -1283
rect 688 -1360 689 -1324
rect 779 -1325 780 -1283
rect 100 -1360 101 -1326
rect 156 -1360 157 -1326
rect 233 -1327 234 -1283
rect 331 -1360 332 -1326
rect 429 -1327 430 -1283
rect 555 -1360 556 -1326
rect 674 -1327 675 -1283
rect 912 -1360 913 -1326
rect 142 -1360 143 -1328
rect 527 -1329 528 -1283
rect 562 -1329 563 -1283
rect 674 -1360 675 -1328
rect 702 -1360 703 -1328
rect 786 -1329 787 -1283
rect 233 -1360 234 -1330
rect 401 -1331 402 -1283
rect 432 -1360 433 -1330
rect 765 -1331 766 -1283
rect 240 -1360 241 -1332
rect 422 -1333 423 -1283
rect 436 -1360 437 -1332
rect 450 -1333 451 -1283
rect 460 -1333 461 -1283
rect 849 -1360 850 -1332
rect 247 -1335 248 -1283
rect 383 -1335 384 -1283
rect 394 -1335 395 -1283
rect 422 -1360 423 -1334
rect 443 -1335 444 -1283
rect 807 -1360 808 -1334
rect 205 -1337 206 -1283
rect 247 -1360 248 -1336
rect 254 -1360 255 -1336
rect 345 -1337 346 -1283
rect 366 -1360 367 -1336
rect 394 -1360 395 -1336
rect 443 -1360 444 -1336
rect 478 -1337 479 -1283
rect 481 -1360 482 -1336
rect 884 -1337 885 -1283
rect 303 -1360 304 -1338
rect 429 -1360 430 -1338
rect 450 -1360 451 -1338
rect 520 -1339 521 -1283
rect 527 -1360 528 -1338
rect 541 -1360 542 -1338
rect 716 -1360 717 -1338
rect 751 -1339 752 -1283
rect 765 -1360 766 -1338
rect 828 -1339 829 -1283
rect 877 -1339 878 -1283
rect 884 -1360 885 -1338
rect 338 -1341 339 -1283
rect 401 -1360 402 -1340
rect 478 -1360 479 -1340
rect 534 -1360 535 -1340
rect 639 -1341 640 -1283
rect 751 -1360 752 -1340
rect 814 -1341 815 -1283
rect 877 -1360 878 -1340
rect 338 -1360 339 -1342
rect 373 -1343 374 -1283
rect 383 -1360 384 -1342
rect 779 -1360 780 -1342
rect 814 -1360 815 -1342
rect 856 -1343 857 -1283
rect 268 -1345 269 -1283
rect 373 -1360 374 -1344
rect 485 -1345 486 -1283
rect 681 -1360 682 -1344
rect 737 -1345 738 -1283
rect 786 -1360 787 -1344
rect 800 -1345 801 -1283
rect 856 -1360 857 -1344
rect 268 -1360 269 -1346
rect 275 -1347 276 -1283
rect 513 -1347 514 -1283
rect 562 -1360 563 -1346
rect 639 -1360 640 -1346
rect 744 -1347 745 -1283
rect 758 -1347 759 -1283
rect 800 -1360 801 -1346
rect 828 -1360 829 -1346
rect 905 -1347 906 -1283
rect 79 -1349 80 -1283
rect 275 -1360 276 -1348
rect 485 -1360 486 -1348
rect 744 -1360 745 -1348
rect 758 -1360 759 -1348
rect 968 -1349 969 -1283
rect 79 -1360 80 -1350
rect 604 -1351 605 -1283
rect 695 -1360 696 -1350
rect 905 -1360 906 -1350
rect 513 -1360 514 -1352
rect 842 -1353 843 -1283
rect 520 -1360 521 -1354
rect 604 -1360 605 -1354
rect 737 -1360 738 -1354
rect 821 -1355 822 -1283
rect 842 -1360 843 -1354
rect 947 -1355 948 -1283
rect 821 -1360 822 -1356
rect 870 -1357 871 -1283
rect 870 -1360 871 -1358
rect 961 -1359 962 -1283
rect 2 -1439 3 -1369
rect 44 -1370 45 -1368
rect 58 -1439 59 -1369
rect 79 -1370 80 -1368
rect 86 -1439 87 -1369
rect 135 -1370 136 -1368
rect 156 -1370 157 -1368
rect 352 -1370 353 -1368
rect 376 -1370 377 -1368
rect 772 -1370 773 -1368
rect 856 -1370 857 -1368
rect 905 -1439 906 -1369
rect 908 -1370 909 -1368
rect 954 -1370 955 -1368
rect 971 -1370 972 -1368
rect 989 -1370 990 -1368
rect 9 -1372 10 -1368
rect 324 -1372 325 -1368
rect 394 -1372 395 -1368
rect 681 -1372 682 -1368
rect 712 -1439 713 -1371
rect 716 -1372 717 -1368
rect 765 -1372 766 -1368
rect 926 -1439 927 -1371
rect 947 -1439 948 -1371
rect 954 -1439 955 -1371
rect 9 -1439 10 -1373
rect 730 -1374 731 -1368
rect 765 -1439 766 -1373
rect 898 -1374 899 -1368
rect 912 -1374 913 -1368
rect 968 -1439 969 -1373
rect 37 -1376 38 -1368
rect 229 -1376 230 -1368
rect 240 -1376 241 -1368
rect 380 -1376 381 -1368
rect 397 -1376 398 -1368
rect 408 -1376 409 -1368
rect 450 -1439 451 -1375
rect 460 -1439 461 -1375
rect 467 -1376 468 -1368
rect 758 -1376 759 -1368
rect 856 -1439 857 -1375
rect 870 -1376 871 -1368
rect 891 -1376 892 -1368
rect 912 -1439 913 -1375
rect 37 -1439 38 -1377
rect 194 -1378 195 -1368
rect 198 -1378 199 -1368
rect 198 -1439 199 -1377
rect 198 -1378 199 -1368
rect 198 -1439 199 -1377
rect 205 -1378 206 -1368
rect 338 -1378 339 -1368
rect 348 -1378 349 -1368
rect 716 -1439 717 -1377
rect 744 -1378 745 -1368
rect 758 -1439 759 -1377
rect 800 -1378 801 -1368
rect 870 -1439 871 -1377
rect 51 -1380 52 -1368
rect 380 -1439 381 -1379
rect 401 -1380 402 -1368
rect 467 -1439 468 -1379
rect 478 -1380 479 -1368
rect 653 -1380 654 -1368
rect 681 -1439 682 -1379
rect 695 -1380 696 -1368
rect 702 -1380 703 -1368
rect 730 -1439 731 -1379
rect 800 -1439 801 -1379
rect 821 -1380 822 -1368
rect 849 -1380 850 -1368
rect 891 -1439 892 -1379
rect 51 -1439 52 -1381
rect 268 -1382 269 -1368
rect 275 -1382 276 -1368
rect 275 -1439 276 -1381
rect 275 -1382 276 -1368
rect 275 -1439 276 -1381
rect 296 -1382 297 -1368
rect 376 -1439 377 -1381
rect 401 -1439 402 -1381
rect 562 -1382 563 -1368
rect 576 -1439 577 -1381
rect 597 -1382 598 -1368
rect 604 -1382 605 -1368
rect 828 -1382 829 -1368
rect 842 -1382 843 -1368
rect 849 -1439 850 -1381
rect 863 -1382 864 -1368
rect 933 -1439 934 -1381
rect 65 -1384 66 -1368
rect 187 -1439 188 -1383
rect 191 -1384 192 -1368
rect 772 -1439 773 -1383
rect 807 -1384 808 -1368
rect 842 -1439 843 -1383
rect 863 -1439 864 -1383
rect 940 -1439 941 -1383
rect 33 -1386 34 -1368
rect 65 -1439 66 -1385
rect 72 -1386 73 -1368
rect 551 -1439 552 -1385
rect 555 -1386 556 -1368
rect 695 -1439 696 -1385
rect 702 -1439 703 -1385
rect 737 -1386 738 -1368
rect 72 -1439 73 -1387
rect 457 -1388 458 -1368
rect 464 -1388 465 -1368
rect 562 -1439 563 -1387
rect 590 -1388 591 -1368
rect 919 -1439 920 -1387
rect 79 -1439 80 -1389
rect 334 -1390 335 -1368
rect 338 -1439 339 -1389
rect 492 -1390 493 -1368
rect 516 -1390 517 -1368
rect 688 -1390 689 -1368
rect 723 -1390 724 -1368
rect 744 -1439 745 -1389
rect 89 -1392 90 -1368
rect 583 -1392 584 -1368
rect 593 -1439 594 -1391
rect 877 -1392 878 -1368
rect 93 -1394 94 -1368
rect 205 -1439 206 -1393
rect 226 -1439 227 -1393
rect 558 -1439 559 -1393
rect 569 -1394 570 -1368
rect 583 -1439 584 -1393
rect 604 -1439 605 -1393
rect 807 -1439 808 -1393
rect 877 -1439 878 -1393
rect 884 -1394 885 -1368
rect 93 -1439 94 -1395
rect 114 -1396 115 -1368
rect 124 -1439 125 -1395
rect 751 -1396 752 -1368
rect 835 -1396 836 -1368
rect 884 -1439 885 -1395
rect 100 -1398 101 -1368
rect 555 -1439 556 -1397
rect 667 -1398 668 -1368
rect 688 -1439 689 -1397
rect 709 -1398 710 -1368
rect 723 -1439 724 -1397
rect 751 -1439 752 -1397
rect 793 -1398 794 -1368
rect 835 -1439 836 -1397
rect 943 -1398 944 -1368
rect 23 -1400 24 -1368
rect 100 -1439 101 -1399
rect 128 -1400 129 -1368
rect 296 -1439 297 -1399
rect 310 -1400 311 -1368
rect 373 -1400 374 -1368
rect 453 -1439 454 -1399
rect 737 -1439 738 -1399
rect 779 -1400 780 -1368
rect 793 -1439 794 -1399
rect 943 -1439 944 -1399
rect 982 -1439 983 -1399
rect 23 -1439 24 -1401
rect 254 -1402 255 -1368
rect 261 -1402 262 -1368
rect 345 -1402 346 -1368
rect 373 -1439 374 -1401
rect 667 -1439 668 -1401
rect 121 -1404 122 -1368
rect 345 -1439 346 -1403
rect 478 -1439 479 -1403
rect 499 -1404 500 -1368
rect 527 -1404 528 -1368
rect 786 -1404 787 -1368
rect 121 -1439 122 -1405
rect 219 -1406 220 -1368
rect 233 -1406 234 -1368
rect 408 -1439 409 -1405
rect 471 -1406 472 -1368
rect 527 -1439 528 -1405
rect 530 -1406 531 -1368
rect 674 -1406 675 -1368
rect 786 -1439 787 -1405
rect 814 -1406 815 -1368
rect 135 -1439 136 -1407
rect 289 -1408 290 -1368
rect 310 -1439 311 -1407
rect 317 -1408 318 -1368
rect 331 -1408 332 -1368
rect 569 -1439 570 -1407
rect 646 -1408 647 -1368
rect 674 -1439 675 -1407
rect 149 -1410 150 -1368
rect 261 -1439 262 -1409
rect 289 -1439 290 -1409
rect 366 -1410 367 -1368
rect 390 -1439 391 -1409
rect 471 -1439 472 -1409
rect 481 -1410 482 -1368
rect 898 -1439 899 -1409
rect 107 -1412 108 -1368
rect 149 -1439 150 -1411
rect 159 -1412 160 -1368
rect 240 -1439 241 -1411
rect 247 -1412 248 -1368
rect 352 -1439 353 -1411
rect 366 -1439 367 -1411
rect 387 -1412 388 -1368
rect 485 -1412 486 -1368
rect 548 -1412 549 -1368
rect 632 -1412 633 -1368
rect 646 -1439 647 -1411
rect 660 -1412 661 -1368
rect 779 -1439 780 -1411
rect 30 -1439 31 -1413
rect 159 -1439 160 -1413
rect 166 -1439 167 -1413
rect 191 -1439 192 -1413
rect 219 -1439 220 -1413
rect 222 -1414 223 -1368
rect 233 -1439 234 -1413
rect 513 -1414 514 -1368
rect 537 -1439 538 -1413
rect 625 -1414 626 -1368
rect 632 -1439 633 -1413
rect 814 -1439 815 -1413
rect 107 -1439 108 -1415
rect 117 -1439 118 -1415
rect 170 -1416 171 -1368
rect 268 -1439 269 -1415
rect 317 -1439 318 -1415
rect 432 -1416 433 -1368
rect 492 -1439 493 -1415
rect 506 -1416 507 -1368
rect 513 -1439 514 -1415
rect 520 -1416 521 -1368
rect 534 -1416 535 -1368
rect 625 -1439 626 -1415
rect 639 -1416 640 -1368
rect 660 -1439 661 -1415
rect 16 -1418 17 -1368
rect 506 -1439 507 -1417
rect 541 -1418 542 -1368
rect 597 -1439 598 -1417
rect 16 -1439 17 -1419
rect 303 -1420 304 -1368
rect 464 -1439 465 -1419
rect 520 -1439 521 -1419
rect 541 -1439 542 -1419
rect 611 -1420 612 -1368
rect 163 -1422 164 -1368
rect 170 -1439 171 -1421
rect 177 -1422 178 -1368
rect 247 -1439 248 -1421
rect 254 -1439 255 -1421
rect 359 -1422 360 -1368
rect 488 -1439 489 -1421
rect 639 -1439 640 -1421
rect 128 -1439 129 -1423
rect 177 -1439 178 -1423
rect 184 -1424 185 -1368
rect 331 -1439 332 -1423
rect 499 -1439 500 -1423
rect 618 -1424 619 -1368
rect 212 -1439 213 -1425
rect 303 -1439 304 -1425
rect 509 -1439 510 -1425
rect 611 -1439 612 -1425
rect 282 -1428 283 -1368
rect 359 -1439 360 -1427
rect 579 -1428 580 -1368
rect 618 -1439 619 -1427
rect 282 -1439 283 -1429
rect 415 -1430 416 -1368
rect 579 -1439 580 -1429
rect 821 -1439 822 -1429
rect 415 -1439 416 -1431
rect 422 -1432 423 -1368
rect 422 -1439 423 -1433
rect 436 -1434 437 -1368
rect 436 -1439 437 -1435
rect 443 -1436 444 -1368
rect 142 -1438 143 -1368
rect 443 -1439 444 -1437
rect 9 -1528 10 -1448
rect 16 -1449 17 -1447
rect 23 -1449 24 -1447
rect 394 -1449 395 -1447
rect 432 -1449 433 -1447
rect 520 -1449 521 -1447
rect 548 -1449 549 -1447
rect 870 -1449 871 -1447
rect 940 -1528 941 -1448
rect 968 -1449 969 -1447
rect 16 -1528 17 -1450
rect 226 -1451 227 -1447
rect 282 -1451 283 -1447
rect 394 -1528 395 -1450
rect 457 -1528 458 -1450
rect 499 -1451 500 -1447
rect 502 -1528 503 -1450
rect 730 -1451 731 -1447
rect 800 -1451 801 -1447
rect 800 -1528 801 -1450
rect 800 -1451 801 -1447
rect 800 -1528 801 -1450
rect 856 -1451 857 -1447
rect 856 -1528 857 -1450
rect 856 -1451 857 -1447
rect 856 -1528 857 -1450
rect 961 -1528 962 -1450
rect 982 -1451 983 -1447
rect 23 -1528 24 -1452
rect 37 -1453 38 -1447
rect 44 -1528 45 -1452
rect 107 -1453 108 -1447
rect 114 -1528 115 -1452
rect 282 -1528 283 -1452
rect 285 -1528 286 -1452
rect 513 -1453 514 -1447
rect 555 -1453 556 -1447
rect 884 -1453 885 -1447
rect 982 -1528 983 -1452
rect 989 -1528 990 -1452
rect 51 -1455 52 -1447
rect 362 -1528 363 -1454
rect 373 -1528 374 -1454
rect 415 -1455 416 -1447
rect 432 -1528 433 -1454
rect 499 -1528 500 -1454
rect 506 -1455 507 -1447
rect 863 -1455 864 -1447
rect 51 -1528 52 -1456
rect 551 -1457 552 -1447
rect 558 -1528 559 -1456
rect 926 -1457 927 -1447
rect 79 -1459 80 -1447
rect 590 -1459 591 -1447
rect 604 -1459 605 -1447
rect 779 -1459 780 -1447
rect 79 -1528 80 -1460
rect 222 -1528 223 -1460
rect 303 -1461 304 -1447
rect 390 -1461 391 -1447
rect 397 -1461 398 -1447
rect 779 -1528 780 -1460
rect 93 -1463 94 -1447
rect 131 -1463 132 -1447
rect 142 -1463 143 -1447
rect 331 -1463 332 -1447
rect 338 -1528 339 -1462
rect 429 -1463 430 -1447
rect 460 -1463 461 -1447
rect 898 -1463 899 -1447
rect 93 -1528 94 -1464
rect 317 -1465 318 -1447
rect 345 -1465 346 -1447
rect 548 -1528 549 -1464
rect 576 -1528 577 -1464
rect 611 -1465 612 -1447
rect 632 -1465 633 -1447
rect 905 -1465 906 -1447
rect 100 -1467 101 -1447
rect 317 -1528 318 -1466
rect 352 -1467 353 -1447
rect 366 -1467 367 -1447
rect 376 -1467 377 -1447
rect 380 -1467 381 -1447
rect 415 -1528 416 -1466
rect 422 -1467 423 -1447
rect 467 -1467 468 -1447
rect 828 -1528 829 -1466
rect 887 -1528 888 -1466
rect 898 -1528 899 -1466
rect 905 -1528 906 -1466
rect 912 -1467 913 -1447
rect 100 -1528 101 -1468
rect 411 -1528 412 -1468
rect 422 -1528 423 -1468
rect 478 -1469 479 -1447
rect 485 -1469 486 -1447
rect 607 -1469 608 -1447
rect 611 -1528 612 -1468
rect 660 -1469 661 -1447
rect 688 -1469 689 -1447
rect 709 -1528 710 -1468
rect 712 -1469 713 -1447
rect 814 -1469 815 -1447
rect 912 -1528 913 -1468
rect 933 -1469 934 -1447
rect 65 -1471 66 -1447
rect 660 -1528 661 -1470
rect 688 -1528 689 -1470
rect 793 -1471 794 -1447
rect 65 -1528 66 -1472
rect 72 -1473 73 -1447
rect 117 -1473 118 -1447
rect 149 -1473 150 -1447
rect 156 -1473 157 -1447
rect 737 -1473 738 -1447
rect 793 -1528 794 -1472
rect 842 -1473 843 -1447
rect 86 -1475 87 -1447
rect 156 -1528 157 -1474
rect 159 -1528 160 -1474
rect 625 -1475 626 -1447
rect 632 -1528 633 -1474
rect 635 -1475 636 -1447
rect 653 -1475 654 -1447
rect 891 -1475 892 -1447
rect 86 -1528 87 -1476
rect 194 -1528 195 -1476
rect 198 -1477 199 -1447
rect 198 -1528 199 -1476
rect 198 -1477 199 -1447
rect 198 -1528 199 -1476
rect 201 -1528 202 -1476
rect 268 -1477 269 -1447
rect 310 -1477 311 -1447
rect 310 -1528 311 -1476
rect 310 -1477 311 -1447
rect 310 -1528 311 -1476
rect 352 -1528 353 -1476
rect 464 -1477 465 -1447
rect 467 -1528 468 -1476
rect 695 -1477 696 -1447
rect 730 -1528 731 -1476
rect 744 -1477 745 -1447
rect 821 -1477 822 -1447
rect 891 -1528 892 -1476
rect 107 -1528 108 -1478
rect 464 -1528 465 -1478
rect 471 -1479 472 -1447
rect 555 -1528 556 -1478
rect 590 -1528 591 -1478
rect 681 -1479 682 -1447
rect 695 -1528 696 -1478
rect 723 -1479 724 -1447
rect 737 -1528 738 -1478
rect 950 -1479 951 -1447
rect 58 -1481 59 -1447
rect 471 -1528 472 -1480
rect 478 -1528 479 -1480
rect 772 -1481 773 -1447
rect 842 -1528 843 -1480
rect 919 -1481 920 -1447
rect 58 -1528 59 -1482
rect 233 -1483 234 -1447
rect 240 -1483 241 -1447
rect 345 -1528 346 -1482
rect 355 -1483 356 -1447
rect 450 -1528 451 -1482
rect 485 -1528 486 -1482
rect 541 -1483 542 -1447
rect 597 -1483 598 -1447
rect 604 -1528 605 -1482
rect 625 -1528 626 -1482
rect 656 -1483 657 -1447
rect 681 -1528 682 -1482
rect 702 -1483 703 -1447
rect 723 -1528 724 -1482
rect 751 -1483 752 -1447
rect 765 -1483 766 -1447
rect 772 -1528 773 -1482
rect 919 -1528 920 -1482
rect 954 -1483 955 -1447
rect 121 -1528 122 -1484
rect 303 -1528 304 -1484
rect 324 -1485 325 -1447
rect 541 -1528 542 -1484
rect 597 -1528 598 -1484
rect 639 -1485 640 -1447
rect 653 -1528 654 -1484
rect 716 -1485 717 -1447
rect 744 -1528 745 -1484
rect 758 -1485 759 -1447
rect 933 -1528 934 -1484
rect 954 -1528 955 -1484
rect 128 -1528 129 -1486
rect 506 -1528 507 -1486
rect 509 -1487 510 -1447
rect 674 -1487 675 -1447
rect 702 -1528 703 -1486
rect 835 -1487 836 -1447
rect 135 -1489 136 -1447
rect 380 -1528 381 -1488
rect 443 -1489 444 -1447
rect 716 -1528 717 -1488
rect 751 -1528 752 -1488
rect 786 -1489 787 -1447
rect 835 -1528 836 -1488
rect 849 -1489 850 -1447
rect 40 -1528 41 -1490
rect 849 -1528 850 -1490
rect 142 -1528 143 -1492
rect 180 -1528 181 -1492
rect 184 -1493 185 -1447
rect 331 -1528 332 -1492
rect 366 -1528 367 -1492
rect 408 -1493 409 -1447
rect 443 -1528 444 -1492
rect 520 -1528 521 -1492
rect 537 -1493 538 -1447
rect 821 -1528 822 -1492
rect 149 -1528 150 -1494
rect 254 -1495 255 -1447
rect 261 -1495 262 -1447
rect 324 -1528 325 -1494
rect 369 -1528 370 -1494
rect 765 -1528 766 -1494
rect 786 -1528 787 -1494
rect 807 -1495 808 -1447
rect 163 -1497 164 -1447
rect 170 -1497 171 -1447
rect 173 -1528 174 -1496
rect 359 -1497 360 -1447
rect 492 -1497 493 -1447
rect 513 -1528 514 -1496
rect 537 -1528 538 -1496
rect 814 -1528 815 -1496
rect 30 -1499 31 -1447
rect 163 -1528 164 -1498
rect 184 -1528 185 -1498
rect 387 -1528 388 -1498
rect 492 -1528 493 -1498
rect 527 -1499 528 -1447
rect 618 -1499 619 -1447
rect 639 -1528 640 -1498
rect 667 -1499 668 -1447
rect 674 -1528 675 -1498
rect 807 -1528 808 -1498
rect 877 -1499 878 -1447
rect 30 -1528 31 -1500
rect 289 -1501 290 -1447
rect 359 -1528 360 -1500
rect 618 -1528 619 -1500
rect 646 -1501 647 -1447
rect 667 -1528 668 -1500
rect 152 -1528 153 -1502
rect 646 -1528 647 -1502
rect 187 -1505 188 -1447
rect 247 -1505 248 -1447
rect 261 -1528 262 -1504
rect 593 -1505 594 -1447
rect 187 -1528 188 -1506
rect 569 -1507 570 -1447
rect 191 -1509 192 -1447
rect 254 -1528 255 -1508
rect 289 -1528 290 -1508
rect 446 -1528 447 -1508
rect 562 -1509 563 -1447
rect 569 -1528 570 -1508
rect 191 -1528 192 -1510
rect 306 -1528 307 -1510
rect 401 -1511 402 -1447
rect 527 -1528 528 -1510
rect 562 -1528 563 -1510
rect 583 -1511 584 -1447
rect 205 -1513 206 -1447
rect 247 -1528 248 -1512
rect 401 -1528 402 -1512
rect 436 -1513 437 -1447
rect 583 -1528 584 -1512
rect 884 -1528 885 -1512
rect 166 -1528 167 -1514
rect 436 -1528 437 -1514
rect 177 -1517 178 -1447
rect 205 -1528 206 -1516
rect 219 -1517 220 -1447
rect 226 -1528 227 -1516
rect 233 -1528 234 -1516
rect 453 -1528 454 -1516
rect 177 -1528 178 -1518
rect 268 -1528 269 -1518
rect 219 -1528 220 -1520
rect 296 -1521 297 -1447
rect 240 -1528 241 -1522
rect 429 -1528 430 -1522
rect 275 -1525 276 -1447
rect 296 -1528 297 -1524
rect 2 -1527 3 -1447
rect 275 -1528 276 -1526
rect 23 -1613 24 -1537
rect 40 -1538 41 -1536
rect 44 -1538 45 -1536
rect 163 -1538 164 -1536
rect 166 -1613 167 -1537
rect 289 -1538 290 -1536
rect 306 -1538 307 -1536
rect 373 -1538 374 -1536
rect 415 -1538 416 -1536
rect 415 -1613 416 -1537
rect 415 -1538 416 -1536
rect 415 -1613 416 -1537
rect 432 -1538 433 -1536
rect 485 -1538 486 -1536
rect 509 -1538 510 -1536
rect 842 -1538 843 -1536
rect 849 -1538 850 -1536
rect 926 -1613 927 -1537
rect 947 -1613 948 -1537
rect 968 -1613 969 -1537
rect 982 -1613 983 -1537
rect 989 -1538 990 -1536
rect 30 -1540 31 -1536
rect 292 -1613 293 -1539
rect 345 -1540 346 -1536
rect 366 -1540 367 -1536
rect 373 -1613 374 -1539
rect 401 -1540 402 -1536
rect 436 -1540 437 -1536
rect 852 -1613 853 -1539
rect 884 -1540 885 -1536
rect 940 -1540 941 -1536
rect 954 -1540 955 -1536
rect 971 -1613 972 -1539
rect 16 -1542 17 -1536
rect 30 -1613 31 -1541
rect 37 -1542 38 -1536
rect 275 -1542 276 -1536
rect 282 -1542 283 -1536
rect 285 -1604 286 -1541
rect 352 -1542 353 -1536
rect 464 -1613 465 -1541
rect 478 -1542 479 -1536
rect 590 -1542 591 -1536
rect 604 -1542 605 -1536
rect 870 -1613 871 -1541
rect 898 -1542 899 -1536
rect 915 -1613 916 -1541
rect 940 -1613 941 -1541
rect 975 -1613 976 -1541
rect 16 -1613 17 -1543
rect 348 -1613 349 -1543
rect 352 -1613 353 -1543
rect 380 -1544 381 -1536
rect 401 -1613 402 -1543
rect 646 -1544 647 -1536
rect 705 -1613 706 -1543
rect 772 -1544 773 -1536
rect 800 -1544 801 -1536
rect 849 -1613 850 -1543
rect 898 -1613 899 -1543
rect 912 -1544 913 -1536
rect 37 -1613 38 -1545
rect 96 -1613 97 -1545
rect 100 -1546 101 -1536
rect 138 -1546 139 -1536
rect 142 -1546 143 -1536
rect 142 -1613 143 -1545
rect 142 -1546 143 -1536
rect 142 -1613 143 -1545
rect 149 -1546 150 -1536
rect 457 -1546 458 -1536
rect 478 -1613 479 -1545
rect 492 -1546 493 -1536
rect 520 -1546 521 -1536
rect 523 -1546 524 -1536
rect 534 -1546 535 -1536
rect 730 -1546 731 -1536
rect 733 -1613 734 -1545
rect 807 -1546 808 -1536
rect 814 -1546 815 -1536
rect 842 -1613 843 -1545
rect 44 -1613 45 -1547
rect 128 -1548 129 -1536
rect 135 -1548 136 -1536
rect 359 -1548 360 -1536
rect 436 -1613 437 -1547
rect 481 -1548 482 -1536
rect 485 -1613 486 -1547
rect 527 -1548 528 -1536
rect 586 -1613 587 -1547
rect 716 -1548 717 -1536
rect 723 -1548 724 -1536
rect 723 -1613 724 -1547
rect 723 -1548 724 -1536
rect 723 -1613 724 -1547
rect 814 -1613 815 -1547
rect 905 -1548 906 -1536
rect 9 -1550 10 -1536
rect 481 -1613 482 -1549
rect 492 -1613 493 -1549
rect 632 -1550 633 -1536
rect 646 -1613 647 -1549
rect 695 -1550 696 -1536
rect 716 -1613 717 -1549
rect 751 -1550 752 -1536
rect 65 -1552 66 -1536
rect 408 -1552 409 -1536
rect 446 -1552 447 -1536
rect 709 -1552 710 -1536
rect 751 -1613 752 -1551
rect 891 -1552 892 -1536
rect 65 -1613 66 -1553
rect 184 -1554 185 -1536
rect 194 -1613 195 -1553
rect 597 -1554 598 -1536
rect 604 -1613 605 -1553
rect 653 -1554 654 -1536
rect 709 -1613 710 -1553
rect 828 -1554 829 -1536
rect 86 -1556 87 -1536
rect 366 -1613 367 -1555
rect 408 -1613 409 -1555
rect 471 -1556 472 -1536
rect 520 -1613 521 -1555
rect 576 -1556 577 -1536
rect 590 -1613 591 -1555
rect 688 -1556 689 -1536
rect 86 -1613 87 -1557
rect 110 -1613 111 -1557
rect 114 -1558 115 -1536
rect 499 -1558 500 -1536
rect 555 -1558 556 -1536
rect 597 -1613 598 -1557
rect 618 -1558 619 -1536
rect 954 -1613 955 -1557
rect 93 -1560 94 -1536
rect 443 -1560 444 -1536
rect 450 -1560 451 -1536
rect 737 -1560 738 -1536
rect 100 -1613 101 -1561
rect 303 -1562 304 -1536
rect 341 -1613 342 -1561
rect 828 -1613 829 -1561
rect 107 -1564 108 -1536
rect 345 -1613 346 -1563
rect 369 -1564 370 -1536
rect 443 -1613 444 -1563
rect 453 -1564 454 -1536
rect 744 -1564 745 -1536
rect 58 -1566 59 -1536
rect 453 -1613 454 -1565
rect 457 -1613 458 -1565
rect 513 -1566 514 -1536
rect 530 -1613 531 -1565
rect 555 -1613 556 -1565
rect 632 -1613 633 -1565
rect 660 -1566 661 -1536
rect 688 -1613 689 -1565
rect 702 -1566 703 -1536
rect 744 -1613 745 -1565
rect 835 -1566 836 -1536
rect 58 -1613 59 -1567
rect 695 -1613 696 -1567
rect 702 -1613 703 -1567
rect 919 -1568 920 -1536
rect 128 -1613 129 -1569
rect 331 -1570 332 -1536
rect 411 -1570 412 -1536
rect 653 -1613 654 -1569
rect 660 -1613 661 -1569
rect 681 -1570 682 -1536
rect 880 -1613 881 -1569
rect 919 -1613 920 -1569
rect 135 -1613 136 -1571
rect 205 -1572 206 -1536
rect 212 -1613 213 -1571
rect 247 -1572 248 -1536
rect 261 -1572 262 -1536
rect 275 -1613 276 -1571
rect 282 -1613 283 -1571
rect 324 -1572 325 -1536
rect 331 -1613 332 -1571
rect 467 -1572 468 -1536
rect 513 -1613 514 -1571
rect 548 -1572 549 -1536
rect 75 -1574 76 -1536
rect 261 -1613 262 -1573
rect 289 -1613 290 -1573
rect 471 -1613 472 -1573
rect 534 -1613 535 -1573
rect 681 -1613 682 -1573
rect 149 -1613 150 -1575
rect 359 -1613 360 -1575
rect 429 -1576 430 -1536
rect 499 -1613 500 -1575
rect 548 -1613 549 -1575
rect 562 -1576 563 -1536
rect 156 -1578 157 -1536
rect 254 -1578 255 -1536
rect 303 -1613 304 -1577
rect 317 -1578 318 -1536
rect 324 -1613 325 -1577
rect 541 -1578 542 -1536
rect 562 -1613 563 -1577
rect 765 -1578 766 -1536
rect 156 -1613 157 -1579
rect 793 -1580 794 -1536
rect 159 -1613 160 -1581
rect 254 -1613 255 -1581
rect 317 -1613 318 -1581
rect 394 -1582 395 -1536
rect 429 -1613 430 -1581
rect 565 -1613 566 -1581
rect 765 -1613 766 -1581
rect 821 -1582 822 -1536
rect 72 -1584 73 -1536
rect 394 -1613 395 -1583
rect 793 -1613 794 -1583
rect 856 -1584 857 -1536
rect 72 -1613 73 -1585
rect 240 -1586 241 -1536
rect 247 -1613 248 -1585
rect 296 -1586 297 -1536
rect 362 -1586 363 -1536
rect 856 -1613 857 -1585
rect 177 -1588 178 -1536
rect 611 -1588 612 -1536
rect 177 -1613 178 -1589
rect 674 -1590 675 -1536
rect 198 -1613 199 -1591
rect 268 -1592 269 -1536
rect 296 -1613 297 -1591
rect 338 -1592 339 -1536
rect 362 -1613 363 -1591
rect 422 -1592 423 -1536
rect 569 -1592 570 -1536
rect 611 -1613 612 -1591
rect 674 -1613 675 -1591
rect 779 -1592 780 -1536
rect 173 -1613 174 -1593
rect 268 -1613 269 -1593
rect 338 -1613 339 -1593
rect 625 -1594 626 -1536
rect 201 -1596 202 -1536
rect 219 -1613 220 -1595
rect 240 -1613 241 -1595
rect 537 -1596 538 -1536
rect 569 -1613 570 -1595
rect 639 -1596 640 -1536
rect 215 -1598 216 -1536
rect 226 -1598 227 -1536
rect 541 -1613 542 -1597
rect 639 -1613 640 -1597
rect 667 -1598 668 -1536
rect 226 -1613 227 -1599
rect 310 -1600 311 -1536
rect 506 -1600 507 -1536
rect 625 -1613 626 -1599
rect 667 -1613 668 -1599
rect 800 -1613 801 -1599
rect 233 -1602 234 -1536
rect 310 -1613 311 -1601
rect 506 -1613 507 -1601
rect 583 -1602 584 -1536
rect 51 -1604 52 -1536
rect 233 -1613 234 -1603
rect 523 -1613 524 -1603
rect 576 -1613 577 -1603
rect 51 -1613 52 -1605
rect 79 -1606 80 -1536
rect 537 -1613 538 -1605
rect 786 -1606 787 -1536
rect 26 -1608 27 -1536
rect 786 -1613 787 -1607
rect 79 -1613 80 -1609
rect 121 -1610 122 -1536
rect 121 -1613 122 -1611
rect 758 -1613 759 -1611
rect 9 -1623 10 -1621
rect 23 -1623 24 -1621
rect 30 -1623 31 -1621
rect 121 -1706 122 -1622
rect 124 -1623 125 -1621
rect 681 -1623 682 -1621
rect 695 -1623 696 -1621
rect 940 -1623 941 -1621
rect 943 -1623 944 -1621
rect 961 -1706 962 -1622
rect 971 -1706 972 -1622
rect 975 -1623 976 -1621
rect 9 -1706 10 -1624
rect 240 -1625 241 -1621
rect 247 -1625 248 -1621
rect 250 -1639 251 -1624
rect 289 -1706 290 -1624
rect 387 -1625 388 -1621
rect 390 -1706 391 -1624
rect 737 -1706 738 -1624
rect 793 -1625 794 -1621
rect 849 -1625 850 -1621
rect 877 -1625 878 -1621
rect 898 -1625 899 -1621
rect 912 -1706 913 -1624
rect 919 -1625 920 -1621
rect 975 -1706 976 -1624
rect 982 -1625 983 -1621
rect 16 -1627 17 -1621
rect 187 -1627 188 -1621
rect 240 -1706 241 -1626
rect 296 -1627 297 -1621
rect 299 -1706 300 -1626
rect 653 -1627 654 -1621
rect 660 -1627 661 -1621
rect 667 -1627 668 -1621
rect 712 -1706 713 -1626
rect 765 -1627 766 -1621
rect 835 -1706 836 -1626
rect 856 -1627 857 -1621
rect 894 -1706 895 -1626
rect 926 -1627 927 -1621
rect 16 -1706 17 -1628
rect 61 -1706 62 -1628
rect 93 -1629 94 -1621
rect 625 -1629 626 -1621
rect 639 -1629 640 -1621
rect 863 -1706 864 -1628
rect 926 -1706 927 -1628
rect 947 -1629 948 -1621
rect 23 -1706 24 -1630
rect 96 -1631 97 -1621
rect 100 -1631 101 -1621
rect 184 -1631 185 -1621
rect 247 -1706 248 -1630
rect 310 -1631 311 -1621
rect 341 -1631 342 -1621
rect 705 -1631 706 -1621
rect 723 -1631 724 -1621
rect 730 -1631 731 -1621
rect 842 -1631 843 -1621
rect 887 -1706 888 -1630
rect 30 -1706 31 -1632
rect 296 -1706 297 -1632
rect 303 -1633 304 -1621
rect 338 -1633 339 -1621
rect 341 -1706 342 -1632
rect 632 -1633 633 -1621
rect 660 -1706 661 -1632
rect 744 -1633 745 -1621
rect 828 -1633 829 -1621
rect 842 -1706 843 -1632
rect 37 -1635 38 -1621
rect 58 -1635 59 -1621
rect 93 -1706 94 -1634
rect 117 -1706 118 -1634
rect 163 -1635 164 -1621
rect 625 -1706 626 -1634
rect 667 -1706 668 -1634
rect 751 -1635 752 -1621
rect 37 -1706 38 -1636
rect 422 -1637 423 -1621
rect 439 -1706 440 -1636
rect 618 -1706 619 -1636
rect 716 -1637 717 -1621
rect 744 -1706 745 -1636
rect 44 -1639 45 -1621
rect 205 -1639 206 -1621
rect 310 -1706 311 -1638
rect 331 -1639 332 -1621
rect 632 -1706 633 -1638
rect 44 -1706 45 -1640
rect 51 -1641 52 -1621
rect 58 -1706 59 -1640
rect 86 -1641 87 -1621
rect 107 -1706 108 -1640
rect 226 -1641 227 -1621
rect 303 -1706 304 -1640
rect 397 -1706 398 -1640
rect 404 -1706 405 -1640
rect 765 -1706 766 -1640
rect 51 -1706 52 -1642
rect 212 -1643 213 -1621
rect 226 -1706 227 -1642
rect 345 -1643 346 -1621
rect 348 -1643 349 -1621
rect 373 -1643 374 -1621
rect 383 -1643 384 -1621
rect 730 -1706 731 -1642
rect 86 -1706 87 -1644
rect 103 -1706 104 -1644
rect 110 -1645 111 -1621
rect 324 -1645 325 -1621
rect 359 -1706 360 -1644
rect 366 -1645 367 -1621
rect 387 -1706 388 -1644
rect 429 -1645 430 -1621
rect 450 -1645 451 -1621
rect 723 -1706 724 -1644
rect 128 -1647 129 -1621
rect 212 -1706 213 -1646
rect 282 -1647 283 -1621
rect 324 -1706 325 -1646
rect 352 -1647 353 -1621
rect 366 -1706 367 -1646
rect 429 -1706 430 -1646
rect 457 -1647 458 -1621
rect 464 -1647 465 -1621
rect 702 -1647 703 -1621
rect 65 -1649 66 -1621
rect 352 -1706 353 -1648
rect 401 -1649 402 -1621
rect 457 -1706 458 -1648
rect 464 -1706 465 -1648
rect 681 -1706 682 -1648
rect 65 -1706 66 -1650
rect 79 -1651 80 -1621
rect 128 -1706 129 -1650
rect 180 -1706 181 -1650
rect 282 -1706 283 -1650
rect 408 -1651 409 -1621
rect 450 -1706 451 -1650
rect 779 -1706 780 -1650
rect 135 -1653 136 -1621
rect 205 -1706 206 -1652
rect 317 -1653 318 -1621
rect 345 -1706 346 -1652
rect 401 -1706 402 -1652
rect 772 -1706 773 -1652
rect 135 -1706 136 -1654
rect 149 -1655 150 -1621
rect 163 -1706 164 -1654
rect 191 -1655 192 -1621
rect 219 -1655 220 -1621
rect 317 -1706 318 -1654
rect 331 -1706 332 -1654
rect 702 -1706 703 -1654
rect 72 -1657 73 -1621
rect 191 -1706 192 -1656
rect 408 -1706 409 -1656
rect 415 -1657 416 -1621
rect 453 -1657 454 -1621
rect 709 -1657 710 -1621
rect 145 -1706 146 -1658
rect 422 -1706 423 -1658
rect 471 -1659 472 -1621
rect 653 -1706 654 -1658
rect 149 -1706 150 -1660
rect 758 -1661 759 -1621
rect 166 -1663 167 -1621
rect 268 -1663 269 -1621
rect 471 -1706 472 -1662
rect 513 -1663 514 -1621
rect 527 -1663 528 -1621
rect 674 -1663 675 -1621
rect 170 -1665 171 -1621
rect 177 -1665 178 -1621
rect 198 -1665 199 -1621
rect 415 -1706 416 -1664
rect 478 -1706 479 -1664
rect 492 -1665 493 -1621
rect 495 -1665 496 -1621
rect 688 -1665 689 -1621
rect 173 -1667 174 -1621
rect 219 -1706 220 -1666
rect 254 -1667 255 -1621
rect 513 -1706 514 -1666
rect 527 -1706 528 -1666
rect 548 -1667 549 -1621
rect 555 -1667 556 -1621
rect 716 -1706 717 -1666
rect 173 -1706 174 -1668
rect 184 -1706 185 -1668
rect 198 -1706 199 -1668
rect 208 -1669 209 -1621
rect 254 -1706 255 -1668
rect 261 -1669 262 -1621
rect 268 -1706 269 -1668
rect 425 -1669 426 -1621
rect 488 -1706 489 -1668
rect 954 -1669 955 -1621
rect 79 -1706 80 -1670
rect 208 -1706 209 -1670
rect 261 -1706 262 -1670
rect 275 -1671 276 -1621
rect 492 -1706 493 -1670
rect 499 -1671 500 -1621
rect 506 -1671 507 -1621
rect 548 -1706 549 -1670
rect 555 -1706 556 -1670
rect 576 -1671 577 -1621
rect 586 -1671 587 -1621
rect 695 -1706 696 -1670
rect 233 -1673 234 -1621
rect 275 -1706 276 -1672
rect 499 -1706 500 -1672
rect 520 -1673 521 -1621
rect 534 -1673 535 -1621
rect 800 -1673 801 -1621
rect 156 -1675 157 -1621
rect 534 -1706 535 -1674
rect 537 -1675 538 -1621
rect 828 -1706 829 -1674
rect 142 -1677 143 -1621
rect 156 -1706 157 -1676
rect 509 -1706 510 -1676
rect 870 -1677 871 -1621
rect 142 -1706 143 -1678
rect 576 -1706 577 -1678
rect 590 -1679 591 -1621
rect 758 -1706 759 -1678
rect 786 -1679 787 -1621
rect 800 -1706 801 -1678
rect 814 -1679 815 -1621
rect 870 -1706 871 -1678
rect 485 -1681 486 -1621
rect 786 -1706 787 -1680
rect 541 -1683 542 -1621
rect 814 -1706 815 -1682
rect 520 -1706 521 -1684
rect 541 -1706 542 -1684
rect 544 -1706 545 -1684
rect 646 -1685 647 -1621
rect 562 -1687 563 -1621
rect 604 -1687 605 -1621
rect 611 -1687 612 -1621
rect 674 -1706 675 -1686
rect 152 -1706 153 -1688
rect 611 -1706 612 -1688
rect 443 -1691 444 -1621
rect 604 -1706 605 -1690
rect 436 -1693 437 -1621
rect 443 -1706 444 -1692
rect 481 -1693 482 -1621
rect 562 -1706 563 -1692
rect 565 -1693 566 -1621
rect 639 -1706 640 -1692
rect 380 -1706 381 -1694
rect 436 -1706 437 -1694
rect 569 -1695 570 -1621
rect 821 -1706 822 -1694
rect 569 -1706 570 -1696
rect 688 -1706 689 -1696
rect 583 -1699 584 -1621
rect 646 -1706 647 -1698
rect 572 -1706 573 -1700
rect 583 -1706 584 -1700
rect 590 -1706 591 -1700
rect 733 -1701 734 -1621
rect 597 -1703 598 -1621
rect 751 -1706 752 -1702
rect 394 -1705 395 -1621
rect 597 -1706 598 -1704
rect 16 -1716 17 -1714
rect 58 -1716 59 -1714
rect 72 -1801 73 -1715
rect 75 -1716 76 -1714
rect 79 -1716 80 -1714
rect 495 -1801 496 -1715
rect 506 -1801 507 -1715
rect 548 -1716 549 -1714
rect 572 -1716 573 -1714
rect 863 -1716 864 -1714
rect 905 -1801 906 -1715
rect 912 -1716 913 -1714
rect 926 -1716 927 -1714
rect 940 -1716 941 -1714
rect 961 -1716 962 -1714
rect 978 -1716 979 -1714
rect 16 -1801 17 -1717
rect 345 -1718 346 -1714
rect 355 -1801 356 -1717
rect 772 -1718 773 -1714
rect 37 -1720 38 -1714
rect 394 -1720 395 -1714
rect 397 -1720 398 -1714
rect 429 -1720 430 -1714
rect 436 -1801 437 -1719
rect 688 -1720 689 -1714
rect 709 -1801 710 -1719
rect 758 -1720 759 -1714
rect 37 -1801 38 -1721
rect 509 -1722 510 -1714
rect 523 -1801 524 -1721
rect 702 -1722 703 -1714
rect 51 -1724 52 -1714
rect 341 -1724 342 -1714
rect 376 -1724 377 -1714
rect 730 -1724 731 -1714
rect 58 -1801 59 -1725
rect 65 -1726 66 -1714
rect 93 -1726 94 -1714
rect 387 -1726 388 -1714
rect 439 -1726 440 -1714
rect 786 -1726 787 -1714
rect 9 -1728 10 -1714
rect 65 -1801 66 -1727
rect 103 -1728 104 -1714
rect 457 -1728 458 -1714
rect 467 -1728 468 -1714
rect 814 -1728 815 -1714
rect 9 -1801 10 -1729
rect 373 -1730 374 -1714
rect 387 -1801 388 -1729
rect 408 -1730 409 -1714
rect 450 -1730 451 -1714
rect 821 -1730 822 -1714
rect 86 -1732 87 -1714
rect 103 -1801 104 -1731
rect 117 -1732 118 -1714
rect 534 -1732 535 -1714
rect 548 -1801 549 -1731
rect 555 -1732 556 -1714
rect 642 -1801 643 -1731
rect 870 -1732 871 -1714
rect 23 -1734 24 -1714
rect 117 -1801 118 -1733
rect 121 -1734 122 -1714
rect 149 -1801 150 -1733
rect 159 -1801 160 -1733
rect 737 -1734 738 -1714
rect 23 -1801 24 -1735
rect 187 -1801 188 -1735
rect 191 -1736 192 -1714
rect 205 -1801 206 -1735
rect 222 -1801 223 -1735
rect 383 -1801 384 -1735
rect 450 -1801 451 -1735
rect 478 -1736 479 -1714
rect 485 -1736 486 -1714
rect 492 -1736 493 -1714
rect 534 -1801 535 -1735
rect 590 -1736 591 -1714
rect 667 -1736 668 -1714
rect 758 -1801 759 -1735
rect 82 -1801 83 -1737
rect 86 -1801 87 -1737
rect 124 -1801 125 -1737
rect 569 -1801 570 -1737
rect 702 -1801 703 -1737
rect 765 -1738 766 -1714
rect 128 -1740 129 -1714
rect 590 -1801 591 -1739
rect 730 -1801 731 -1739
rect 800 -1740 801 -1714
rect 142 -1801 143 -1741
rect 660 -1742 661 -1714
rect 737 -1801 738 -1741
rect 828 -1742 829 -1714
rect 163 -1744 164 -1714
rect 170 -1744 171 -1714
rect 173 -1801 174 -1743
rect 261 -1744 262 -1714
rect 268 -1744 269 -1714
rect 334 -1744 335 -1714
rect 471 -1744 472 -1714
rect 485 -1801 486 -1743
rect 488 -1744 489 -1714
rect 667 -1801 668 -1743
rect 166 -1801 167 -1745
rect 422 -1746 423 -1714
rect 474 -1801 475 -1745
rect 716 -1746 717 -1714
rect 170 -1801 171 -1747
rect 408 -1801 409 -1747
rect 422 -1801 423 -1747
rect 887 -1748 888 -1714
rect 191 -1801 192 -1749
rect 247 -1750 248 -1714
rect 261 -1801 262 -1749
rect 303 -1750 304 -1714
rect 310 -1750 311 -1714
rect 376 -1801 377 -1749
rect 478 -1801 479 -1749
rect 527 -1750 528 -1714
rect 555 -1801 556 -1749
rect 611 -1750 612 -1714
rect 660 -1801 661 -1749
rect 723 -1750 724 -1714
rect 107 -1752 108 -1714
rect 303 -1801 304 -1751
rect 324 -1752 325 -1714
rect 345 -1801 346 -1751
rect 527 -1801 528 -1751
rect 576 -1752 577 -1714
rect 716 -1801 717 -1751
rect 842 -1752 843 -1714
rect 107 -1801 108 -1753
rect 135 -1754 136 -1714
rect 156 -1754 157 -1714
rect 247 -1801 248 -1753
rect 271 -1801 272 -1753
rect 835 -1754 836 -1714
rect 30 -1756 31 -1714
rect 156 -1801 157 -1755
rect 219 -1756 220 -1714
rect 310 -1801 311 -1755
rect 324 -1801 325 -1755
rect 338 -1756 339 -1714
rect 576 -1801 577 -1755
rect 625 -1756 626 -1714
rect 723 -1801 724 -1755
rect 779 -1756 780 -1714
rect 30 -1801 31 -1757
rect 51 -1801 52 -1757
rect 219 -1801 220 -1757
rect 429 -1801 430 -1757
rect 625 -1801 626 -1757
rect 695 -1758 696 -1714
rect 226 -1760 227 -1714
rect 541 -1760 542 -1714
rect 695 -1801 696 -1759
rect 744 -1760 745 -1714
rect 114 -1801 115 -1761
rect 226 -1801 227 -1761
rect 233 -1762 234 -1714
rect 415 -1762 416 -1714
rect 541 -1801 542 -1761
rect 597 -1762 598 -1714
rect 639 -1762 640 -1714
rect 744 -1801 745 -1761
rect 198 -1764 199 -1714
rect 233 -1801 234 -1763
rect 236 -1764 237 -1714
rect 611 -1801 612 -1763
rect 198 -1801 199 -1765
rect 320 -1801 321 -1765
rect 338 -1801 339 -1765
rect 366 -1766 367 -1714
rect 415 -1801 416 -1765
rect 520 -1766 521 -1714
rect 597 -1801 598 -1765
rect 646 -1766 647 -1714
rect 240 -1768 241 -1714
rect 401 -1768 402 -1714
rect 443 -1768 444 -1714
rect 646 -1801 647 -1767
rect 44 -1770 45 -1714
rect 443 -1801 444 -1769
rect 44 -1801 45 -1771
rect 499 -1772 500 -1714
rect 240 -1801 241 -1773
rect 369 -1801 370 -1773
rect 499 -1801 500 -1773
rect 653 -1774 654 -1714
rect 254 -1776 255 -1714
rect 639 -1801 640 -1775
rect 653 -1801 654 -1775
rect 751 -1776 752 -1714
rect 184 -1778 185 -1714
rect 254 -1801 255 -1777
rect 275 -1778 276 -1714
rect 688 -1801 689 -1777
rect 184 -1801 185 -1779
rect 359 -1780 360 -1714
rect 583 -1780 584 -1714
rect 751 -1801 752 -1779
rect 212 -1782 213 -1714
rect 275 -1801 276 -1781
rect 282 -1782 283 -1714
rect 464 -1782 465 -1714
rect 583 -1801 584 -1781
rect 618 -1782 619 -1714
rect 93 -1801 94 -1783
rect 212 -1801 213 -1783
rect 282 -1801 283 -1783
rect 453 -1784 454 -1714
rect 464 -1801 465 -1783
rect 513 -1784 514 -1714
rect 618 -1801 619 -1783
rect 681 -1784 682 -1714
rect 289 -1786 290 -1714
rect 457 -1801 458 -1785
rect 562 -1786 563 -1714
rect 681 -1801 682 -1785
rect 180 -1801 181 -1787
rect 289 -1801 290 -1787
rect 296 -1788 297 -1714
rect 331 -1788 332 -1714
rect 352 -1788 353 -1714
rect 562 -1801 563 -1787
rect 296 -1801 297 -1789
rect 380 -1790 381 -1714
rect 401 -1801 402 -1789
rect 513 -1801 514 -1789
rect 299 -1792 300 -1714
rect 471 -1801 472 -1791
rect 317 -1794 318 -1714
rect 331 -1801 332 -1793
rect 359 -1801 360 -1793
rect 604 -1794 605 -1714
rect 604 -1801 605 -1795
rect 674 -1796 675 -1714
rect 632 -1798 633 -1714
rect 674 -1801 675 -1797
rect 352 -1801 353 -1799
rect 632 -1801 633 -1799
rect 9 -1811 10 -1809
rect 30 -1811 31 -1809
rect 33 -1882 34 -1810
rect 37 -1882 38 -1810
rect 40 -1811 41 -1809
rect 82 -1811 83 -1809
rect 89 -1811 90 -1809
rect 422 -1811 423 -1809
rect 457 -1811 458 -1809
rect 457 -1882 458 -1810
rect 457 -1811 458 -1809
rect 457 -1882 458 -1810
rect 471 -1882 472 -1810
rect 478 -1811 479 -1809
rect 492 -1811 493 -1809
rect 758 -1811 759 -1809
rect 23 -1813 24 -1809
rect 86 -1882 87 -1812
rect 93 -1813 94 -1809
rect 212 -1882 213 -1812
rect 219 -1813 220 -1809
rect 275 -1813 276 -1809
rect 306 -1882 307 -1812
rect 338 -1813 339 -1809
rect 345 -1813 346 -1809
rect 355 -1813 356 -1809
rect 366 -1882 367 -1812
rect 376 -1882 377 -1812
rect 380 -1813 381 -1809
rect 555 -1813 556 -1809
rect 579 -1882 580 -1812
rect 737 -1813 738 -1809
rect 744 -1813 745 -1809
rect 744 -1882 745 -1812
rect 744 -1813 745 -1809
rect 744 -1882 745 -1812
rect 44 -1815 45 -1809
rect 478 -1882 479 -1814
rect 492 -1882 493 -1814
rect 499 -1815 500 -1809
rect 506 -1815 507 -1809
rect 604 -1815 605 -1809
rect 667 -1815 668 -1809
rect 667 -1882 668 -1814
rect 667 -1815 668 -1809
rect 667 -1882 668 -1814
rect 674 -1815 675 -1809
rect 677 -1835 678 -1814
rect 723 -1815 724 -1809
rect 723 -1882 724 -1814
rect 723 -1815 724 -1809
rect 723 -1882 724 -1814
rect 737 -1882 738 -1814
rect 751 -1815 752 -1809
rect 51 -1882 52 -1816
rect 107 -1817 108 -1809
rect 121 -1817 122 -1809
rect 331 -1817 332 -1809
rect 348 -1882 349 -1816
rect 688 -1817 689 -1809
rect 58 -1819 59 -1809
rect 58 -1882 59 -1818
rect 58 -1819 59 -1809
rect 58 -1882 59 -1818
rect 65 -1819 66 -1809
rect 215 -1819 216 -1809
rect 219 -1882 220 -1818
rect 282 -1819 283 -1809
rect 331 -1882 332 -1818
rect 464 -1819 465 -1809
rect 495 -1819 496 -1809
rect 751 -1882 752 -1818
rect 65 -1882 66 -1820
rect 233 -1821 234 -1809
rect 240 -1821 241 -1809
rect 502 -1882 503 -1820
rect 513 -1882 514 -1820
rect 527 -1821 528 -1809
rect 604 -1882 605 -1820
rect 611 -1821 612 -1809
rect 653 -1821 654 -1809
rect 688 -1882 689 -1820
rect 72 -1823 73 -1809
rect 222 -1823 223 -1809
rect 240 -1882 241 -1822
rect 296 -1823 297 -1809
rect 352 -1823 353 -1809
rect 422 -1882 423 -1822
rect 464 -1882 465 -1822
rect 534 -1823 535 -1809
rect 611 -1882 612 -1822
rect 618 -1823 619 -1809
rect 674 -1882 675 -1822
rect 681 -1823 682 -1809
rect 72 -1882 73 -1824
rect 142 -1825 143 -1809
rect 149 -1825 150 -1809
rect 177 -1882 178 -1824
rect 184 -1882 185 -1824
rect 191 -1825 192 -1809
rect 201 -1882 202 -1824
rect 394 -1825 395 -1809
rect 415 -1825 416 -1809
rect 506 -1882 507 -1824
rect 516 -1825 517 -1809
rect 730 -1825 731 -1809
rect 47 -1882 48 -1826
rect 415 -1882 416 -1826
rect 453 -1882 454 -1826
rect 534 -1882 535 -1826
rect 618 -1882 619 -1826
rect 632 -1827 633 -1809
rect 681 -1882 682 -1826
rect 709 -1827 710 -1809
rect 79 -1882 80 -1828
rect 114 -1829 115 -1809
rect 121 -1882 122 -1828
rect 191 -1882 192 -1828
rect 268 -1829 269 -1809
rect 590 -1829 591 -1809
rect 695 -1829 696 -1809
rect 709 -1882 710 -1828
rect 93 -1882 94 -1830
rect 499 -1882 500 -1830
rect 509 -1831 510 -1809
rect 632 -1882 633 -1830
rect 695 -1882 696 -1830
rect 716 -1831 717 -1809
rect 103 -1833 104 -1809
rect 289 -1833 290 -1809
rect 296 -1882 297 -1832
rect 303 -1833 304 -1809
rect 338 -1882 339 -1832
rect 730 -1882 731 -1832
rect 107 -1882 108 -1834
rect 198 -1835 199 -1809
rect 275 -1882 276 -1834
rect 443 -1835 444 -1809
rect 520 -1882 521 -1834
rect 548 -1835 549 -1809
rect 590 -1882 591 -1834
rect 625 -1835 626 -1809
rect 716 -1882 717 -1834
rect 100 -1882 101 -1836
rect 198 -1882 199 -1836
rect 282 -1882 283 -1836
rect 485 -1837 486 -1809
rect 625 -1882 626 -1836
rect 660 -1837 661 -1809
rect 124 -1839 125 -1809
rect 527 -1882 528 -1838
rect 642 -1882 643 -1838
rect 660 -1882 661 -1838
rect 128 -1841 129 -1809
rect 247 -1841 248 -1809
rect 352 -1882 353 -1840
rect 653 -1882 654 -1840
rect 135 -1843 136 -1809
rect 436 -1843 437 -1809
rect 443 -1882 444 -1842
rect 541 -1843 542 -1809
rect 142 -1882 143 -1844
rect 254 -1845 255 -1809
rect 355 -1882 356 -1844
rect 569 -1845 570 -1809
rect 156 -1882 157 -1846
rect 205 -1847 206 -1809
rect 247 -1882 248 -1846
rect 261 -1847 262 -1809
rect 310 -1847 311 -1809
rect 569 -1882 570 -1846
rect 16 -1849 17 -1809
rect 205 -1882 206 -1848
rect 254 -1882 255 -1848
rect 362 -1882 363 -1848
rect 369 -1849 370 -1809
rect 597 -1849 598 -1809
rect 16 -1882 17 -1850
rect 292 -1882 293 -1850
rect 310 -1882 311 -1850
rect 324 -1851 325 -1809
rect 359 -1851 360 -1809
rect 380 -1882 381 -1850
rect 387 -1851 388 -1809
rect 394 -1882 395 -1850
rect 450 -1851 451 -1809
rect 597 -1882 598 -1850
rect 163 -1853 164 -1809
rect 562 -1853 563 -1809
rect 12 -1855 13 -1809
rect 562 -1882 563 -1854
rect 131 -1882 132 -1856
rect 163 -1882 164 -1856
rect 166 -1857 167 -1809
rect 555 -1882 556 -1856
rect 170 -1859 171 -1809
rect 233 -1882 234 -1858
rect 261 -1882 262 -1858
rect 401 -1859 402 -1809
rect 485 -1882 486 -1858
rect 747 -1882 748 -1858
rect 135 -1882 136 -1860
rect 170 -1882 171 -1860
rect 173 -1861 174 -1809
rect 401 -1882 402 -1860
rect 187 -1863 188 -1809
rect 226 -1863 227 -1809
rect 268 -1882 269 -1862
rect 450 -1882 451 -1862
rect 114 -1882 115 -1864
rect 226 -1882 227 -1864
rect 324 -1882 325 -1864
rect 541 -1882 542 -1864
rect 373 -1867 374 -1809
rect 702 -1867 703 -1809
rect 303 -1882 304 -1868
rect 373 -1882 374 -1868
rect 387 -1882 388 -1868
rect 583 -1869 584 -1809
rect 390 -1882 391 -1870
rect 646 -1871 647 -1809
rect 180 -1873 181 -1809
rect 646 -1882 647 -1872
rect 408 -1875 409 -1809
rect 702 -1882 703 -1874
rect 408 -1882 409 -1876
rect 429 -1877 430 -1809
rect 576 -1877 577 -1809
rect 583 -1882 584 -1876
rect 317 -1879 318 -1809
rect 429 -1882 430 -1878
rect 138 -1881 139 -1809
rect 317 -1882 318 -1880
rect 2 -1965 3 -1891
rect 72 -1892 73 -1890
rect 107 -1892 108 -1890
rect 170 -1892 171 -1890
rect 177 -1892 178 -1890
rect 191 -1965 192 -1891
rect 194 -1892 195 -1890
rect 415 -1892 416 -1890
rect 432 -1965 433 -1891
rect 737 -1892 738 -1890
rect 5 -1894 6 -1890
rect 198 -1894 199 -1890
rect 201 -1965 202 -1893
rect 369 -1965 370 -1893
rect 376 -1894 377 -1890
rect 646 -1894 647 -1890
rect 709 -1894 710 -1890
rect 747 -1894 748 -1890
rect 9 -1965 10 -1895
rect 387 -1896 388 -1890
rect 397 -1965 398 -1895
rect 555 -1896 556 -1890
rect 583 -1896 584 -1890
rect 583 -1965 584 -1895
rect 583 -1896 584 -1890
rect 583 -1965 584 -1895
rect 604 -1896 605 -1890
rect 604 -1965 605 -1895
rect 604 -1896 605 -1890
rect 604 -1965 605 -1895
rect 611 -1896 612 -1890
rect 611 -1965 612 -1895
rect 611 -1896 612 -1890
rect 611 -1965 612 -1895
rect 12 -1898 13 -1890
rect 170 -1965 171 -1897
rect 177 -1965 178 -1897
rect 226 -1965 227 -1897
rect 240 -1898 241 -1890
rect 327 -1898 328 -1890
rect 338 -1965 339 -1897
rect 534 -1898 535 -1890
rect 541 -1898 542 -1890
rect 555 -1965 556 -1897
rect 23 -1900 24 -1890
rect 233 -1900 234 -1890
rect 292 -1900 293 -1890
rect 569 -1900 570 -1890
rect 23 -1965 24 -1901
rect 464 -1902 465 -1890
rect 471 -1902 472 -1890
rect 548 -1902 549 -1890
rect 562 -1902 563 -1890
rect 569 -1965 570 -1901
rect 33 -1965 34 -1903
rect 37 -1904 38 -1890
rect 44 -1965 45 -1903
rect 268 -1904 269 -1890
rect 296 -1904 297 -1890
rect 306 -1904 307 -1890
rect 317 -1904 318 -1890
rect 418 -1965 419 -1903
rect 436 -1904 437 -1890
rect 597 -1904 598 -1890
rect 26 -1906 27 -1890
rect 268 -1965 269 -1905
rect 296 -1965 297 -1905
rect 324 -1906 325 -1890
rect 345 -1965 346 -1905
rect 702 -1906 703 -1890
rect 51 -1908 52 -1890
rect 149 -1908 150 -1890
rect 156 -1908 157 -1890
rect 303 -1908 304 -1890
rect 324 -1965 325 -1907
rect 506 -1908 507 -1890
rect 520 -1908 521 -1890
rect 534 -1965 535 -1907
rect 541 -1965 542 -1907
rect 590 -1908 591 -1890
rect 597 -1965 598 -1907
rect 632 -1908 633 -1890
rect 674 -1908 675 -1890
rect 702 -1965 703 -1907
rect 51 -1965 52 -1909
rect 58 -1910 59 -1890
rect 61 -1965 62 -1909
rect 79 -1910 80 -1890
rect 117 -1965 118 -1909
rect 156 -1965 157 -1909
rect 184 -1910 185 -1890
rect 222 -1965 223 -1909
rect 254 -1910 255 -1890
rect 317 -1965 318 -1909
rect 359 -1910 360 -1890
rect 562 -1965 563 -1909
rect 590 -1965 591 -1909
rect 660 -1910 661 -1890
rect 667 -1910 668 -1890
rect 674 -1965 675 -1909
rect 65 -1912 66 -1890
rect 166 -1912 167 -1890
rect 184 -1965 185 -1911
rect 219 -1912 220 -1890
rect 303 -1965 304 -1911
rect 460 -1965 461 -1911
rect 471 -1965 472 -1911
rect 481 -1965 482 -1911
rect 502 -1912 503 -1890
rect 723 -1912 724 -1890
rect 65 -1965 66 -1913
rect 282 -1914 283 -1890
rect 331 -1914 332 -1890
rect 359 -1965 360 -1913
rect 362 -1914 363 -1890
rect 366 -1914 367 -1890
rect 380 -1914 381 -1890
rect 520 -1965 521 -1913
rect 625 -1914 626 -1890
rect 660 -1965 661 -1913
rect 16 -1916 17 -1890
rect 282 -1965 283 -1915
rect 366 -1965 367 -1915
rect 646 -1965 647 -1915
rect 72 -1965 73 -1917
rect 579 -1918 580 -1890
rect 618 -1918 619 -1890
rect 625 -1965 626 -1917
rect 639 -1918 640 -1890
rect 723 -1965 724 -1917
rect 79 -1965 80 -1919
rect 499 -1965 500 -1919
rect 506 -1965 507 -1919
rect 527 -1920 528 -1890
rect 618 -1965 619 -1919
rect 751 -1920 752 -1890
rect 19 -1965 20 -1921
rect 527 -1965 528 -1921
rect 114 -1924 115 -1890
rect 254 -1965 255 -1923
rect 261 -1924 262 -1890
rect 331 -1965 332 -1923
rect 380 -1965 381 -1923
rect 394 -1924 395 -1890
rect 401 -1924 402 -1890
rect 576 -1965 577 -1923
rect 100 -1926 101 -1890
rect 261 -1965 262 -1925
rect 355 -1965 356 -1925
rect 394 -1965 395 -1925
rect 401 -1965 402 -1925
rect 422 -1926 423 -1890
rect 429 -1926 430 -1890
rect 667 -1965 668 -1925
rect 100 -1965 101 -1927
rect 632 -1965 633 -1927
rect 121 -1930 122 -1890
rect 121 -1965 122 -1929
rect 121 -1930 122 -1890
rect 121 -1965 122 -1929
rect 128 -1965 129 -1929
rect 310 -1930 311 -1890
rect 429 -1965 430 -1929
rect 467 -1930 468 -1890
rect 131 -1932 132 -1890
rect 653 -1932 654 -1890
rect 145 -1934 146 -1890
rect 373 -1965 374 -1933
rect 436 -1965 437 -1933
rect 485 -1934 486 -1890
rect 205 -1936 206 -1890
rect 289 -1965 290 -1935
rect 310 -1965 311 -1935
rect 457 -1936 458 -1890
rect 485 -1965 486 -1935
rect 513 -1936 514 -1890
rect 149 -1965 150 -1937
rect 205 -1965 206 -1937
rect 208 -1965 209 -1937
rect 730 -1938 731 -1890
rect 142 -1940 143 -1890
rect 730 -1965 731 -1939
rect 86 -1942 87 -1890
rect 142 -1965 143 -1941
rect 212 -1942 213 -1890
rect 240 -1965 241 -1941
rect 271 -1965 272 -1941
rect 653 -1965 654 -1941
rect 86 -1965 87 -1943
rect 135 -1944 136 -1890
rect 163 -1965 164 -1943
rect 212 -1965 213 -1943
rect 219 -1965 220 -1943
rect 233 -1965 234 -1943
rect 352 -1965 353 -1943
rect 513 -1965 514 -1943
rect 135 -1965 136 -1945
rect 408 -1946 409 -1890
rect 439 -1946 440 -1890
rect 709 -1965 710 -1945
rect 275 -1948 276 -1890
rect 408 -1965 409 -1947
rect 443 -1965 444 -1947
rect 492 -1948 493 -1890
rect 247 -1950 248 -1890
rect 275 -1965 276 -1949
rect 422 -1965 423 -1949
rect 492 -1965 493 -1949
rect 93 -1952 94 -1890
rect 247 -1965 248 -1951
rect 450 -1952 451 -1890
rect 688 -1952 689 -1890
rect 37 -1965 38 -1953
rect 688 -1965 689 -1953
rect 93 -1965 94 -1955
rect 348 -1965 349 -1955
rect 450 -1965 451 -1955
rect 478 -1956 479 -1890
rect 478 -1965 479 -1957
rect 716 -1958 717 -1890
rect 695 -1960 696 -1890
rect 716 -1965 717 -1959
rect 681 -1962 682 -1890
rect 695 -1965 696 -1961
rect 54 -1965 55 -1963
rect 681 -1965 682 -1963
rect 16 -2026 17 -1974
rect 142 -1975 143 -1973
rect 156 -1975 157 -1973
rect 261 -1975 262 -1973
rect 285 -2026 286 -1974
rect 632 -1975 633 -1973
rect 635 -2026 636 -1974
rect 716 -1975 717 -1973
rect 19 -1977 20 -1973
rect 331 -1977 332 -1973
rect 366 -1977 367 -1973
rect 590 -1977 591 -1973
rect 642 -1977 643 -1973
rect 695 -1977 696 -1973
rect 23 -1979 24 -1973
rect 205 -2026 206 -1978
rect 240 -1979 241 -1973
rect 313 -1979 314 -1973
rect 324 -1979 325 -1973
rect 439 -2026 440 -1978
rect 450 -1979 451 -1973
rect 488 -2026 489 -1978
rect 534 -1979 535 -1973
rect 548 -1979 549 -1973
rect 551 -1979 552 -1973
rect 660 -1979 661 -1973
rect 695 -2026 696 -1978
rect 723 -1979 724 -1973
rect 23 -2026 24 -1980
rect 30 -1981 31 -1973
rect 37 -2026 38 -1980
rect 75 -1981 76 -1973
rect 100 -1981 101 -1973
rect 359 -1981 360 -1973
rect 366 -2026 367 -1980
rect 551 -2026 552 -1980
rect 562 -1981 563 -1973
rect 639 -1981 640 -1973
rect 30 -2026 31 -1982
rect 107 -1983 108 -1973
rect 110 -1983 111 -1973
rect 159 -1983 160 -1973
rect 163 -1983 164 -1973
rect 324 -2026 325 -1982
rect 331 -2026 332 -1982
rect 397 -1983 398 -1973
rect 404 -2026 405 -1982
rect 471 -1983 472 -1973
rect 478 -2026 479 -1982
rect 632 -2026 633 -1982
rect 44 -1985 45 -1973
rect 432 -1985 433 -1973
rect 443 -1985 444 -1973
rect 450 -2026 451 -1984
rect 457 -1985 458 -1973
rect 583 -1985 584 -1973
rect 618 -1985 619 -1973
rect 660 -2026 661 -1984
rect 44 -2026 45 -1986
rect 86 -1987 87 -1973
rect 93 -1987 94 -1973
rect 163 -2026 164 -1986
rect 170 -1987 171 -1973
rect 296 -1987 297 -1973
rect 303 -1987 304 -1973
rect 310 -2026 311 -1986
rect 369 -1987 370 -1973
rect 667 -1987 668 -1973
rect 51 -2026 52 -1988
rect 688 -1989 689 -1973
rect 58 -2026 59 -1990
rect 103 -2026 104 -1990
rect 107 -2026 108 -1990
rect 135 -1991 136 -1973
rect 142 -2026 143 -1990
rect 212 -1991 213 -1973
rect 219 -1991 220 -1973
rect 296 -2026 297 -1990
rect 387 -1991 388 -1973
rect 569 -1991 570 -1973
rect 583 -2026 584 -1990
rect 646 -1991 647 -1973
rect 65 -1993 66 -1973
rect 79 -2026 80 -1992
rect 100 -2026 101 -1992
rect 709 -1993 710 -1973
rect 2 -1995 3 -1973
rect 65 -2026 66 -1994
rect 68 -2026 69 -1994
rect 156 -2026 157 -1994
rect 177 -1995 178 -1973
rect 208 -1995 209 -1973
rect 215 -1995 216 -1973
rect 646 -2026 647 -1994
rect 72 -2026 73 -1996
rect 89 -2026 90 -1996
rect 117 -1997 118 -1973
rect 499 -1997 500 -1973
rect 534 -2026 535 -1996
rect 681 -1997 682 -1973
rect 117 -2026 118 -1998
rect 135 -2026 136 -1998
rect 149 -1999 150 -1973
rect 170 -2026 171 -1998
rect 177 -2026 178 -1998
rect 184 -1999 185 -1973
rect 191 -1999 192 -1973
rect 240 -2026 241 -1998
rect 254 -1999 255 -1973
rect 268 -1999 269 -1973
rect 289 -1999 290 -1973
rect 352 -2026 353 -1998
rect 387 -2026 388 -1998
rect 408 -1999 409 -1973
rect 415 -1999 416 -1973
rect 590 -2026 591 -1998
rect 604 -1999 605 -1973
rect 618 -2026 619 -1998
rect 9 -2001 10 -1973
rect 149 -2026 150 -2000
rect 184 -2026 185 -2000
rect 555 -2001 556 -1973
rect 562 -2026 563 -2000
rect 597 -2001 598 -1973
rect 604 -2026 605 -2000
rect 674 -2001 675 -1973
rect 9 -2026 10 -2002
rect 173 -2003 174 -1973
rect 219 -2026 220 -2002
rect 233 -2003 234 -1973
rect 247 -2003 248 -1973
rect 268 -2026 269 -2002
rect 289 -2026 290 -2002
rect 338 -2003 339 -1973
rect 380 -2003 381 -1973
rect 415 -2026 416 -2002
rect 418 -2003 419 -1973
rect 506 -2003 507 -1973
rect 569 -2026 570 -2002
rect 653 -2003 654 -1973
rect 54 -2005 55 -1973
rect 338 -2026 339 -2004
rect 394 -2026 395 -2004
rect 401 -2005 402 -1973
rect 408 -2026 409 -2004
rect 436 -2005 437 -1973
rect 443 -2026 444 -2004
rect 513 -2005 514 -1973
rect 597 -2026 598 -2004
rect 730 -2005 731 -1973
rect 54 -2026 55 -2006
rect 499 -2026 500 -2006
rect 506 -2026 507 -2006
rect 576 -2007 577 -1973
rect 642 -2026 643 -2006
rect 653 -2026 654 -2006
rect 121 -2009 122 -1973
rect 201 -2009 202 -1973
rect 226 -2009 227 -1973
rect 247 -2026 248 -2008
rect 261 -2026 262 -2008
rect 275 -2009 276 -1973
rect 422 -2026 423 -2008
rect 481 -2009 482 -1973
rect 513 -2026 514 -2008
rect 541 -2009 542 -1973
rect 576 -2026 577 -2008
rect 625 -2009 626 -1973
rect 128 -2011 129 -1973
rect 359 -2026 360 -2010
rect 457 -2026 458 -2010
rect 485 -2011 486 -1973
rect 541 -2026 542 -2010
rect 611 -2011 612 -1973
rect 625 -2026 626 -2010
rect 649 -2026 650 -2010
rect 121 -2026 122 -2012
rect 128 -2026 129 -2012
rect 131 -2026 132 -2012
rect 306 -2026 307 -2012
rect 464 -2013 465 -1973
rect 520 -2013 521 -1973
rect 611 -2026 612 -2012
rect 702 -2013 703 -1973
rect 226 -2026 227 -2014
rect 373 -2015 374 -1973
rect 474 -2026 475 -2014
rect 555 -2026 556 -2014
rect 233 -2026 234 -2016
rect 345 -2017 346 -1973
rect 373 -2026 374 -2016
rect 429 -2017 430 -1973
rect 492 -2017 493 -1973
rect 520 -2026 521 -2016
rect 275 -2026 276 -2018
rect 317 -2019 318 -1973
rect 429 -2026 430 -2018
rect 527 -2019 528 -1973
rect 282 -2021 283 -1973
rect 317 -2026 318 -2020
rect 348 -2021 349 -1973
rect 527 -2026 528 -2020
rect 282 -2026 283 -2022
rect 464 -2026 465 -2022
rect 303 -2026 304 -2024
rect 345 -2026 346 -2024
rect 436 -2026 437 -2024
rect 492 -2026 493 -2024
rect 9 -2036 10 -2034
rect 201 -2036 202 -2034
rect 212 -2036 213 -2034
rect 429 -2036 430 -2034
rect 436 -2036 437 -2034
rect 625 -2036 626 -2034
rect 632 -2036 633 -2034
rect 639 -2036 640 -2034
rect 646 -2091 647 -2035
rect 660 -2036 661 -2034
rect 688 -2091 689 -2035
rect 695 -2036 696 -2034
rect 16 -2038 17 -2034
rect 96 -2038 97 -2034
rect 114 -2038 115 -2034
rect 289 -2038 290 -2034
rect 296 -2038 297 -2034
rect 296 -2091 297 -2037
rect 296 -2038 297 -2034
rect 296 -2091 297 -2037
rect 303 -2038 304 -2034
rect 352 -2038 353 -2034
rect 380 -2038 381 -2034
rect 443 -2038 444 -2034
rect 474 -2038 475 -2034
rect 513 -2038 514 -2034
rect 520 -2091 521 -2037
rect 541 -2038 542 -2034
rect 548 -2038 549 -2034
rect 583 -2038 584 -2034
rect 16 -2091 17 -2039
rect 128 -2040 129 -2034
rect 177 -2040 178 -2034
rect 177 -2091 178 -2039
rect 177 -2040 178 -2034
rect 177 -2091 178 -2039
rect 191 -2040 192 -2034
rect 387 -2040 388 -2034
rect 415 -2091 416 -2039
rect 534 -2040 535 -2034
rect 541 -2091 542 -2039
rect 562 -2040 563 -2034
rect 30 -2042 31 -2034
rect 117 -2042 118 -2034
rect 121 -2042 122 -2034
rect 121 -2091 122 -2041
rect 121 -2042 122 -2034
rect 121 -2091 122 -2041
rect 128 -2091 129 -2041
rect 135 -2042 136 -2034
rect 191 -2091 192 -2041
rect 240 -2042 241 -2034
rect 257 -2042 258 -2034
rect 261 -2042 262 -2034
rect 289 -2091 290 -2041
rect 471 -2042 472 -2034
rect 481 -2091 482 -2041
rect 569 -2042 570 -2034
rect 37 -2044 38 -2034
rect 254 -2044 255 -2034
rect 303 -2091 304 -2043
rect 436 -2091 437 -2043
rect 443 -2091 444 -2043
rect 450 -2044 451 -2034
rect 471 -2091 472 -2043
rect 506 -2044 507 -2034
rect 548 -2091 549 -2043
rect 576 -2044 577 -2034
rect 33 -2091 34 -2045
rect 37 -2091 38 -2045
rect 44 -2046 45 -2034
rect 86 -2046 87 -2034
rect 100 -2091 101 -2045
rect 114 -2091 115 -2045
rect 117 -2091 118 -2045
rect 184 -2046 185 -2034
rect 198 -2046 199 -2034
rect 404 -2046 405 -2034
rect 425 -2091 426 -2045
rect 597 -2046 598 -2034
rect 44 -2091 45 -2047
rect 142 -2048 143 -2034
rect 194 -2091 195 -2047
rect 198 -2091 199 -2047
rect 205 -2048 206 -2034
rect 261 -2091 262 -2047
rect 313 -2091 314 -2047
rect 576 -2091 577 -2047
rect 51 -2050 52 -2034
rect 72 -2050 73 -2034
rect 79 -2050 80 -2034
rect 418 -2050 419 -2034
rect 429 -2091 430 -2049
rect 478 -2050 479 -2034
rect 485 -2091 486 -2049
rect 642 -2050 643 -2034
rect 51 -2091 52 -2051
rect 96 -2091 97 -2051
rect 212 -2091 213 -2051
rect 310 -2052 311 -2034
rect 320 -2091 321 -2051
rect 513 -2091 514 -2051
rect 555 -2052 556 -2034
rect 653 -2052 654 -2034
rect 65 -2054 66 -2034
rect 499 -2054 500 -2034
rect 555 -2091 556 -2053
rect 618 -2054 619 -2034
rect 642 -2091 643 -2053
rect 674 -2091 675 -2053
rect 65 -2091 66 -2055
rect 170 -2056 171 -2034
rect 215 -2056 216 -2034
rect 670 -2056 671 -2034
rect 75 -2091 76 -2057
rect 79 -2091 80 -2057
rect 86 -2091 87 -2057
rect 107 -2058 108 -2034
rect 170 -2091 171 -2057
rect 275 -2058 276 -2034
rect 327 -2091 328 -2057
rect 345 -2058 346 -2034
rect 359 -2058 360 -2034
rect 387 -2091 388 -2057
rect 418 -2091 419 -2057
rect 583 -2091 584 -2057
rect 107 -2091 108 -2059
rect 163 -2060 164 -2034
rect 219 -2060 220 -2034
rect 527 -2060 528 -2034
rect 562 -2091 563 -2059
rect 611 -2060 612 -2034
rect 58 -2062 59 -2034
rect 219 -2091 220 -2061
rect 222 -2062 223 -2034
rect 226 -2062 227 -2034
rect 236 -2091 237 -2061
rect 569 -2091 570 -2061
rect 604 -2062 605 -2034
rect 611 -2091 612 -2061
rect 58 -2091 59 -2063
rect 89 -2064 90 -2034
rect 149 -2064 150 -2034
rect 359 -2091 360 -2063
rect 383 -2091 384 -2063
rect 408 -2064 409 -2034
rect 450 -2091 451 -2063
rect 457 -2064 458 -2034
rect 492 -2064 493 -2034
rect 506 -2091 507 -2063
rect 149 -2091 150 -2065
rect 233 -2066 234 -2034
rect 240 -2091 241 -2065
rect 324 -2066 325 -2034
rect 331 -2066 332 -2034
rect 401 -2066 402 -2034
rect 408 -2091 409 -2065
rect 527 -2091 528 -2065
rect 135 -2091 136 -2067
rect 324 -2091 325 -2067
rect 338 -2068 339 -2034
rect 492 -2091 493 -2067
rect 499 -2091 500 -2067
rect 635 -2068 636 -2034
rect 156 -2070 157 -2034
rect 457 -2091 458 -2069
rect 142 -2091 143 -2071
rect 156 -2091 157 -2071
rect 159 -2091 160 -2071
rect 163 -2091 164 -2071
rect 222 -2091 223 -2071
rect 247 -2091 248 -2071
rect 254 -2091 255 -2071
rect 373 -2072 374 -2034
rect 394 -2072 395 -2034
rect 604 -2091 605 -2071
rect 226 -2091 227 -2073
rect 369 -2091 370 -2073
rect 373 -2091 374 -2073
rect 478 -2091 479 -2073
rect 268 -2076 269 -2034
rect 338 -2091 339 -2075
rect 345 -2091 346 -2075
rect 380 -2091 381 -2075
rect 394 -2091 395 -2075
rect 422 -2076 423 -2034
rect 268 -2091 269 -2077
rect 366 -2078 367 -2034
rect 401 -2091 402 -2077
rect 464 -2078 465 -2034
rect 275 -2091 276 -2079
rect 404 -2091 405 -2079
rect 317 -2082 318 -2034
rect 331 -2091 332 -2081
rect 352 -2091 353 -2081
rect 464 -2091 465 -2081
rect 317 -2091 318 -2083
rect 534 -2091 535 -2083
rect 366 -2091 367 -2085
rect 590 -2086 591 -2034
rect 282 -2088 283 -2034
rect 590 -2091 591 -2087
rect 282 -2091 283 -2089
rect 306 -2091 307 -2089
rect 23 -2101 24 -2099
rect 58 -2101 59 -2099
rect 65 -2101 66 -2099
rect 310 -2101 311 -2099
rect 324 -2148 325 -2100
rect 345 -2101 346 -2099
rect 366 -2148 367 -2100
rect 408 -2148 409 -2100
rect 429 -2101 430 -2099
rect 429 -2148 430 -2100
rect 429 -2101 430 -2099
rect 429 -2148 430 -2100
rect 509 -2148 510 -2100
rect 520 -2101 521 -2099
rect 523 -2148 524 -2100
rect 569 -2101 570 -2099
rect 590 -2101 591 -2099
rect 597 -2148 598 -2100
rect 611 -2101 612 -2099
rect 621 -2101 622 -2099
rect 642 -2101 643 -2099
rect 646 -2101 647 -2099
rect 674 -2101 675 -2099
rect 688 -2101 689 -2099
rect 26 -2148 27 -2102
rect 75 -2103 76 -2099
rect 100 -2103 101 -2099
rect 100 -2148 101 -2102
rect 100 -2103 101 -2099
rect 100 -2148 101 -2102
rect 107 -2103 108 -2099
rect 306 -2103 307 -2099
rect 310 -2148 311 -2102
rect 338 -2103 339 -2099
rect 345 -2148 346 -2102
rect 383 -2103 384 -2099
rect 394 -2103 395 -2099
rect 401 -2148 402 -2102
rect 530 -2148 531 -2102
rect 583 -2103 584 -2099
rect 611 -2148 612 -2102
rect 618 -2103 619 -2099
rect 33 -2148 34 -2104
rect 37 -2105 38 -2099
rect 44 -2105 45 -2099
rect 317 -2105 318 -2099
rect 331 -2105 332 -2099
rect 569 -2148 570 -2104
rect 37 -2148 38 -2106
rect 128 -2107 129 -2099
rect 135 -2107 136 -2099
rect 138 -2119 139 -2106
rect 156 -2148 157 -2106
rect 177 -2107 178 -2099
rect 187 -2107 188 -2099
rect 320 -2107 321 -2099
rect 338 -2148 339 -2106
rect 380 -2148 381 -2106
rect 387 -2107 388 -2099
rect 394 -2148 395 -2106
rect 534 -2107 535 -2099
rect 555 -2148 556 -2106
rect 562 -2107 563 -2099
rect 590 -2148 591 -2106
rect 44 -2148 45 -2108
rect 184 -2109 185 -2099
rect 208 -2109 209 -2099
rect 268 -2109 269 -2099
rect 282 -2109 283 -2099
rect 352 -2148 353 -2108
rect 359 -2109 360 -2099
rect 387 -2148 388 -2108
rect 464 -2109 465 -2099
rect 534 -2148 535 -2108
rect 541 -2109 542 -2099
rect 541 -2148 542 -2108
rect 541 -2109 542 -2099
rect 541 -2148 542 -2108
rect 51 -2111 52 -2099
rect 152 -2148 153 -2110
rect 163 -2111 164 -2099
rect 205 -2111 206 -2099
rect 215 -2148 216 -2110
rect 527 -2111 528 -2099
rect 51 -2148 52 -2112
rect 198 -2113 199 -2099
rect 205 -2148 206 -2112
rect 212 -2113 213 -2099
rect 222 -2148 223 -2112
rect 502 -2113 503 -2099
rect 58 -2148 59 -2114
rect 86 -2115 87 -2099
rect 107 -2148 108 -2114
rect 121 -2115 122 -2099
rect 135 -2148 136 -2114
rect 142 -2115 143 -2099
rect 149 -2115 150 -2099
rect 163 -2148 164 -2114
rect 170 -2115 171 -2099
rect 191 -2148 192 -2114
rect 198 -2148 199 -2114
rect 289 -2115 290 -2099
rect 296 -2115 297 -2099
rect 296 -2148 297 -2114
rect 296 -2115 297 -2099
rect 296 -2148 297 -2114
rect 303 -2148 304 -2114
rect 562 -2148 563 -2114
rect 65 -2148 66 -2116
rect 79 -2117 80 -2099
rect 86 -2148 87 -2116
rect 226 -2117 227 -2099
rect 233 -2117 234 -2099
rect 240 -2117 241 -2099
rect 247 -2117 248 -2099
rect 558 -2117 559 -2099
rect 16 -2119 17 -2099
rect 79 -2148 80 -2118
rect 142 -2148 143 -2118
rect 170 -2148 171 -2118
rect 264 -2148 265 -2118
rect 268 -2148 269 -2118
rect 306 -2148 307 -2118
rect 369 -2119 370 -2099
rect 604 -2119 605 -2099
rect 72 -2121 73 -2099
rect 117 -2121 118 -2099
rect 177 -2148 178 -2120
rect 478 -2148 479 -2120
rect 117 -2148 118 -2122
rect 289 -2148 290 -2122
rect 233 -2148 234 -2124
rect 275 -2125 276 -2099
rect 240 -2148 241 -2126
rect 334 -2148 335 -2126
rect 247 -2148 248 -2128
rect 443 -2129 444 -2099
rect 254 -2131 255 -2099
rect 292 -2148 293 -2130
rect 443 -2148 444 -2130
rect 450 -2131 451 -2099
rect 226 -2148 227 -2132
rect 254 -2148 255 -2132
rect 261 -2133 262 -2099
rect 275 -2148 276 -2132
rect 450 -2148 451 -2132
rect 471 -2133 472 -2099
rect 261 -2148 262 -2134
rect 513 -2135 514 -2099
rect 422 -2137 423 -2099
rect 471 -2148 472 -2136
rect 513 -2148 514 -2136
rect 548 -2137 549 -2099
rect 422 -2148 423 -2138
rect 436 -2139 437 -2099
rect 492 -2139 493 -2099
rect 548 -2148 549 -2138
rect 373 -2141 374 -2099
rect 436 -2148 437 -2140
rect 492 -2148 493 -2140
rect 506 -2141 507 -2099
rect 373 -2148 374 -2142
rect 457 -2143 458 -2099
rect 457 -2148 458 -2144
rect 485 -2145 486 -2099
rect 485 -2148 486 -2146
rect 576 -2147 577 -2099
rect 9 -2195 10 -2157
rect 19 -2195 20 -2157
rect 37 -2158 38 -2156
rect 215 -2195 216 -2157
rect 240 -2158 241 -2156
rect 282 -2158 283 -2156
rect 285 -2195 286 -2157
rect 296 -2158 297 -2156
rect 317 -2158 318 -2156
rect 408 -2158 409 -2156
rect 415 -2158 416 -2156
rect 548 -2158 549 -2156
rect 590 -2158 591 -2156
rect 604 -2195 605 -2157
rect 611 -2158 612 -2156
rect 611 -2195 612 -2157
rect 611 -2158 612 -2156
rect 611 -2195 612 -2157
rect 44 -2160 45 -2156
rect 184 -2160 185 -2156
rect 208 -2195 209 -2159
rect 289 -2195 290 -2159
rect 292 -2160 293 -2156
rect 310 -2160 311 -2156
rect 317 -2195 318 -2159
rect 387 -2160 388 -2156
rect 408 -2195 409 -2159
rect 443 -2160 444 -2156
rect 450 -2160 451 -2156
rect 467 -2160 468 -2156
rect 499 -2160 500 -2156
rect 555 -2160 556 -2156
rect 597 -2160 598 -2156
rect 600 -2195 601 -2159
rect 51 -2162 52 -2156
rect 261 -2195 262 -2161
rect 275 -2162 276 -2156
rect 303 -2162 304 -2156
rect 324 -2162 325 -2156
rect 334 -2162 335 -2156
rect 352 -2162 353 -2156
rect 359 -2162 360 -2156
rect 362 -2162 363 -2156
rect 485 -2162 486 -2156
rect 541 -2162 542 -2156
rect 555 -2195 556 -2161
rect 51 -2195 52 -2163
rect 149 -2195 150 -2163
rect 163 -2164 164 -2156
rect 187 -2164 188 -2156
rect 247 -2164 248 -2156
rect 373 -2195 374 -2163
rect 387 -2195 388 -2163
rect 422 -2164 423 -2156
rect 425 -2195 426 -2163
rect 478 -2164 479 -2156
rect 58 -2166 59 -2156
rect 96 -2166 97 -2156
rect 107 -2166 108 -2156
rect 128 -2166 129 -2156
rect 131 -2166 132 -2156
rect 135 -2166 136 -2156
rect 163 -2195 164 -2165
rect 180 -2166 181 -2156
rect 268 -2166 269 -2156
rect 303 -2195 304 -2165
rect 324 -2195 325 -2165
rect 345 -2166 346 -2156
rect 352 -2195 353 -2165
rect 569 -2166 570 -2156
rect 58 -2195 59 -2167
rect 177 -2168 178 -2156
rect 278 -2195 279 -2167
rect 348 -2195 349 -2167
rect 366 -2168 367 -2156
rect 562 -2168 563 -2156
rect 65 -2170 66 -2156
rect 72 -2170 73 -2156
rect 79 -2195 80 -2169
rect 156 -2170 157 -2156
rect 177 -2195 178 -2169
rect 338 -2170 339 -2156
rect 345 -2195 346 -2169
rect 534 -2170 535 -2156
rect 40 -2195 41 -2171
rect 72 -2195 73 -2171
rect 86 -2172 87 -2156
rect 268 -2195 269 -2171
rect 296 -2195 297 -2171
rect 464 -2195 465 -2171
rect 513 -2172 514 -2156
rect 534 -2195 535 -2171
rect 65 -2195 66 -2173
rect 219 -2174 220 -2156
rect 331 -2195 332 -2173
rect 394 -2174 395 -2156
rect 415 -2195 416 -2173
rect 520 -2195 521 -2173
rect 86 -2195 87 -2175
rect 142 -2176 143 -2156
rect 156 -2195 157 -2175
rect 170 -2176 171 -2156
rect 219 -2195 220 -2175
rect 257 -2195 258 -2175
rect 394 -2195 395 -2175
rect 481 -2195 482 -2175
rect 93 -2178 94 -2156
rect 100 -2178 101 -2156
rect 107 -2195 108 -2177
rect 128 -2195 129 -2177
rect 135 -2195 136 -2177
rect 212 -2178 213 -2156
rect 429 -2178 430 -2156
rect 443 -2195 444 -2177
rect 453 -2195 454 -2177
rect 471 -2178 472 -2156
rect 93 -2195 94 -2179
rect 138 -2195 139 -2179
rect 205 -2180 206 -2156
rect 212 -2195 213 -2179
rect 429 -2195 430 -2179
rect 492 -2180 493 -2156
rect 100 -2195 101 -2181
rect 198 -2182 199 -2156
rect 380 -2182 381 -2156
rect 492 -2195 493 -2181
rect 121 -2184 122 -2156
rect 233 -2184 234 -2156
rect 380 -2195 381 -2183
rect 401 -2184 402 -2156
rect 436 -2184 437 -2156
rect 509 -2184 510 -2156
rect 121 -2195 122 -2185
rect 131 -2195 132 -2185
rect 170 -2195 171 -2185
rect 233 -2195 234 -2185
rect 436 -2195 437 -2185
rect 457 -2186 458 -2156
rect 198 -2195 199 -2187
rect 247 -2195 248 -2187
rect 457 -2195 458 -2187
rect 499 -2195 500 -2187
rect 226 -2190 227 -2156
rect 401 -2195 402 -2189
rect 191 -2192 192 -2156
rect 226 -2195 227 -2191
rect 187 -2195 188 -2193
rect 191 -2195 192 -2193
rect 9 -2205 10 -2203
rect 16 -2224 17 -2204
rect 23 -2205 24 -2203
rect 26 -2224 27 -2204
rect 44 -2205 45 -2203
rect 44 -2224 45 -2204
rect 44 -2205 45 -2203
rect 44 -2224 45 -2204
rect 51 -2205 52 -2203
rect 103 -2224 104 -2204
rect 107 -2205 108 -2203
rect 201 -2205 202 -2203
rect 240 -2224 241 -2204
rect 380 -2205 381 -2203
rect 408 -2205 409 -2203
rect 418 -2205 419 -2203
rect 429 -2205 430 -2203
rect 450 -2224 451 -2204
rect 457 -2205 458 -2203
rect 506 -2224 507 -2204
rect 534 -2205 535 -2203
rect 548 -2205 549 -2203
rect 600 -2205 601 -2203
rect 604 -2205 605 -2203
rect 611 -2205 612 -2203
rect 611 -2224 612 -2204
rect 611 -2205 612 -2203
rect 611 -2224 612 -2204
rect 51 -2224 52 -2206
rect 82 -2224 83 -2206
rect 86 -2207 87 -2203
rect 205 -2207 206 -2203
rect 254 -2207 255 -2203
rect 464 -2207 465 -2203
rect 537 -2224 538 -2206
rect 555 -2207 556 -2203
rect 58 -2209 59 -2203
rect 128 -2209 129 -2203
rect 149 -2209 150 -2203
rect 156 -2209 157 -2203
rect 177 -2209 178 -2203
rect 205 -2224 206 -2208
rect 254 -2224 255 -2208
rect 289 -2209 290 -2203
rect 299 -2209 300 -2203
rect 362 -2209 363 -2203
rect 366 -2209 367 -2203
rect 387 -2209 388 -2203
rect 394 -2209 395 -2203
rect 408 -2224 409 -2208
rect 422 -2209 423 -2203
rect 534 -2224 535 -2208
rect 58 -2224 59 -2210
rect 93 -2211 94 -2203
rect 100 -2211 101 -2203
rect 212 -2224 213 -2210
rect 247 -2211 248 -2203
rect 289 -2224 290 -2210
rect 303 -2211 304 -2203
rect 341 -2224 342 -2210
rect 359 -2211 360 -2203
rect 520 -2211 521 -2203
rect 65 -2213 66 -2203
rect 145 -2213 146 -2203
rect 149 -2224 150 -2212
rect 163 -2213 164 -2203
rect 177 -2224 178 -2212
rect 261 -2213 262 -2203
rect 268 -2213 269 -2203
rect 348 -2224 349 -2212
rect 373 -2224 374 -2212
rect 436 -2213 437 -2203
rect 443 -2213 444 -2203
rect 492 -2213 493 -2203
rect 79 -2215 80 -2203
rect 208 -2224 209 -2214
rect 247 -2224 248 -2214
rect 317 -2215 318 -2203
rect 324 -2215 325 -2203
rect 352 -2215 353 -2203
rect 107 -2224 108 -2216
rect 170 -2217 171 -2203
rect 187 -2224 188 -2216
rect 219 -2217 220 -2203
rect 268 -2224 269 -2216
rect 345 -2217 346 -2203
rect 114 -2219 115 -2203
rect 121 -2219 122 -2203
rect 191 -2219 192 -2203
rect 282 -2224 283 -2218
rect 72 -2221 73 -2203
rect 114 -2224 115 -2220
rect 191 -2224 192 -2220
rect 226 -2221 227 -2203
rect 275 -2224 276 -2220
rect 331 -2221 332 -2203
rect 226 -2224 227 -2222
rect 327 -2224 328 -2222
rect 331 -2224 332 -2222
rect 401 -2223 402 -2203
rect 58 -2234 59 -2232
rect 93 -2234 94 -2232
rect 107 -2234 108 -2232
rect 173 -2234 174 -2232
rect 201 -2234 202 -2232
rect 268 -2234 269 -2232
rect 275 -2234 276 -2232
rect 327 -2234 328 -2232
rect 331 -2234 332 -2232
rect 383 -2234 384 -2232
rect 408 -2234 409 -2232
rect 429 -2234 430 -2232
rect 450 -2234 451 -2232
rect 474 -2234 475 -2232
rect 485 -2234 486 -2232
rect 506 -2234 507 -2232
rect 75 -2236 76 -2232
rect 114 -2236 115 -2232
rect 131 -2236 132 -2232
rect 226 -2236 227 -2232
rect 240 -2236 241 -2232
rect 390 -2236 391 -2232
rect 149 -2238 150 -2232
rect 163 -2238 164 -2232
rect 219 -2238 220 -2232
rect 282 -2238 283 -2232
rect 289 -2238 290 -2232
rect 303 -2238 304 -2232
rect 310 -2238 311 -2232
rect 373 -2238 374 -2232
rect 247 -2240 248 -2232
rect 355 -2240 356 -2232
rect 254 -2242 255 -2232
rect 313 -2242 314 -2232
<< labels >>
rlabel pdiffusion 3 -10 3 -10 0 cellNo=55
rlabel pdiffusion 10 -10 10 -10 0 cellNo=456
rlabel pdiffusion 17 -10 17 -10 0 cellNo=496
rlabel pdiffusion 24 -10 24 -10 0 cellNo=330
rlabel pdiffusion 31 -10 31 -10 0 cellNo=470
rlabel pdiffusion 38 -10 38 -10 0 cellNo=100
rlabel pdiffusion 45 -10 45 -10 0 cellNo=292
rlabel pdiffusion 52 -10 52 -10 0 cellNo=357
rlabel pdiffusion 59 -10 59 -10 0 cellNo=377
rlabel pdiffusion 66 -10 66 -10 0 cellNo=418
rlabel pdiffusion 73 -10 73 -10 0 cellNo=934
rlabel pdiffusion 108 -10 108 -10 0 cellNo=16
rlabel pdiffusion 115 -10 115 -10 0 cellNo=870
rlabel pdiffusion 129 -10 129 -10 0 cellNo=229
rlabel pdiffusion 136 -10 136 -10 0 cellNo=621
rlabel pdiffusion 143 -10 143 -10 0 cellNo=466
rlabel pdiffusion 157 -10 157 -10 0 feedthrough
rlabel pdiffusion 164 -10 164 -10 0 feedthrough
rlabel pdiffusion 171 -10 171 -10 0 cellNo=186
rlabel pdiffusion 178 -10 178 -10 0 feedthrough
rlabel pdiffusion 185 -10 185 -10 0 cellNo=93
rlabel pdiffusion 192 -10 192 -10 0 feedthrough
rlabel pdiffusion 199 -10 199 -10 0 cellNo=367
rlabel pdiffusion 206 -10 206 -10 0 cellNo=440
rlabel pdiffusion 213 -10 213 -10 0 cellNo=954
rlabel pdiffusion 220 -10 220 -10 0 cellNo=275
rlabel pdiffusion 227 -10 227 -10 0 feedthrough
rlabel pdiffusion 234 -10 234 -10 0 cellNo=798
rlabel pdiffusion 241 -10 241 -10 0 cellNo=489
rlabel pdiffusion 248 -10 248 -10 0 feedthrough
rlabel pdiffusion 255 -10 255 -10 0 cellNo=343
rlabel pdiffusion 262 -10 262 -10 0 feedthrough
rlabel pdiffusion 269 -10 269 -10 0 feedthrough
rlabel pdiffusion 276 -10 276 -10 0 cellNo=171
rlabel pdiffusion 283 -10 283 -10 0 cellNo=838
rlabel pdiffusion 325 -10 325 -10 0 cellNo=784
rlabel pdiffusion 3 -37 3 -37 0 cellNo=213
rlabel pdiffusion 10 -37 10 -37 0 cellNo=407
rlabel pdiffusion 17 -37 17 -37 0 cellNo=951
rlabel pdiffusion 24 -37 24 -37 0 cellNo=399
rlabel pdiffusion 31 -37 31 -37 0 cellNo=351
rlabel pdiffusion 38 -37 38 -37 0 cellNo=458
rlabel pdiffusion 45 -37 45 -37 0 cellNo=988
rlabel pdiffusion 73 -37 73 -37 0 cellNo=682
rlabel pdiffusion 80 -37 80 -37 0 cellNo=855
rlabel pdiffusion 87 -37 87 -37 0 feedthrough
rlabel pdiffusion 94 -37 94 -37 0 feedthrough
rlabel pdiffusion 101 -37 101 -37 0 cellNo=41
rlabel pdiffusion 108 -37 108 -37 0 cellNo=586
rlabel pdiffusion 115 -37 115 -37 0 cellNo=204
rlabel pdiffusion 122 -37 122 -37 0 cellNo=165
rlabel pdiffusion 129 -37 129 -37 0 cellNo=321
rlabel pdiffusion 136 -37 136 -37 0 cellNo=497
rlabel pdiffusion 143 -37 143 -37 0 feedthrough
rlabel pdiffusion 150 -37 150 -37 0 feedthrough
rlabel pdiffusion 157 -37 157 -37 0 feedthrough
rlabel pdiffusion 164 -37 164 -37 0 cellNo=510
rlabel pdiffusion 171 -37 171 -37 0 feedthrough
rlabel pdiffusion 178 -37 178 -37 0 cellNo=400
rlabel pdiffusion 185 -37 185 -37 0 feedthrough
rlabel pdiffusion 192 -37 192 -37 0 feedthrough
rlabel pdiffusion 199 -37 199 -37 0 feedthrough
rlabel pdiffusion 206 -37 206 -37 0 cellNo=82
rlabel pdiffusion 213 -37 213 -37 0 cellNo=322
rlabel pdiffusion 220 -37 220 -37 0 feedthrough
rlabel pdiffusion 227 -37 227 -37 0 cellNo=243
rlabel pdiffusion 234 -37 234 -37 0 feedthrough
rlabel pdiffusion 241 -37 241 -37 0 feedthrough
rlabel pdiffusion 248 -37 248 -37 0 feedthrough
rlabel pdiffusion 255 -37 255 -37 0 feedthrough
rlabel pdiffusion 262 -37 262 -37 0 feedthrough
rlabel pdiffusion 269 -37 269 -37 0 feedthrough
rlabel pdiffusion 276 -37 276 -37 0 feedthrough
rlabel pdiffusion 283 -37 283 -37 0 cellNo=537
rlabel pdiffusion 290 -37 290 -37 0 feedthrough
rlabel pdiffusion 297 -37 297 -37 0 feedthrough
rlabel pdiffusion 304 -37 304 -37 0 feedthrough
rlabel pdiffusion 311 -37 311 -37 0 cellNo=437
rlabel pdiffusion 318 -37 318 -37 0 feedthrough
rlabel pdiffusion 325 -37 325 -37 0 cellNo=790
rlabel pdiffusion 332 -37 332 -37 0 feedthrough
rlabel pdiffusion 339 -37 339 -37 0 cellNo=221
rlabel pdiffusion 346 -37 346 -37 0 feedthrough
rlabel pdiffusion 353 -37 353 -37 0 feedthrough
rlabel pdiffusion 360 -37 360 -37 0 feedthrough
rlabel pdiffusion 367 -37 367 -37 0 cellNo=2
rlabel pdiffusion 374 -37 374 -37 0 cellNo=26
rlabel pdiffusion 381 -37 381 -37 0 feedthrough
rlabel pdiffusion 388 -37 388 -37 0 feedthrough
rlabel pdiffusion 395 -37 395 -37 0 cellNo=450
rlabel pdiffusion 402 -37 402 -37 0 feedthrough
rlabel pdiffusion 416 -37 416 -37 0 cellNo=785
rlabel pdiffusion 3 -80 3 -80 0 cellNo=95
rlabel pdiffusion 10 -80 10 -80 0 cellNo=301
rlabel pdiffusion 17 -80 17 -80 0 cellNo=539
rlabel pdiffusion 24 -80 24 -80 0 cellNo=394
rlabel pdiffusion 31 -80 31 -80 0 cellNo=531
rlabel pdiffusion 38 -80 38 -80 0 cellNo=339
rlabel pdiffusion 45 -80 45 -80 0 feedthrough
rlabel pdiffusion 52 -80 52 -80 0 feedthrough
rlabel pdiffusion 59 -80 59 -80 0 cellNo=631
rlabel pdiffusion 66 -80 66 -80 0 feedthrough
rlabel pdiffusion 73 -80 73 -80 0 cellNo=43
rlabel pdiffusion 80 -80 80 -80 0 feedthrough
rlabel pdiffusion 87 -80 87 -80 0 cellNo=746
rlabel pdiffusion 94 -80 94 -80 0 cellNo=675
rlabel pdiffusion 101 -80 101 -80 0 cellNo=515
rlabel pdiffusion 108 -80 108 -80 0 feedthrough
rlabel pdiffusion 115 -80 115 -80 0 cellNo=460
rlabel pdiffusion 122 -80 122 -80 0 cellNo=230
rlabel pdiffusion 129 -80 129 -80 0 cellNo=125
rlabel pdiffusion 136 -80 136 -80 0 feedthrough
rlabel pdiffusion 143 -80 143 -80 0 cellNo=410
rlabel pdiffusion 150 -80 150 -80 0 feedthrough
rlabel pdiffusion 157 -80 157 -80 0 cellNo=154
rlabel pdiffusion 164 -80 164 -80 0 feedthrough
rlabel pdiffusion 171 -80 171 -80 0 cellNo=471
rlabel pdiffusion 178 -80 178 -80 0 cellNo=731
rlabel pdiffusion 185 -80 185 -80 0 feedthrough
rlabel pdiffusion 192 -80 192 -80 0 cellNo=188
rlabel pdiffusion 199 -80 199 -80 0 cellNo=472
rlabel pdiffusion 206 -80 206 -80 0 cellNo=416
rlabel pdiffusion 213 -80 213 -80 0 cellNo=465
rlabel pdiffusion 220 -80 220 -80 0 cellNo=955
rlabel pdiffusion 227 -80 227 -80 0 cellNo=14
rlabel pdiffusion 234 -80 234 -80 0 feedthrough
rlabel pdiffusion 241 -80 241 -80 0 feedthrough
rlabel pdiffusion 248 -80 248 -80 0 feedthrough
rlabel pdiffusion 255 -80 255 -80 0 cellNo=27
rlabel pdiffusion 262 -80 262 -80 0 feedthrough
rlabel pdiffusion 269 -80 269 -80 0 cellNo=573
rlabel pdiffusion 276 -80 276 -80 0 cellNo=591
rlabel pdiffusion 283 -80 283 -80 0 cellNo=664
rlabel pdiffusion 290 -80 290 -80 0 feedthrough
rlabel pdiffusion 297 -80 297 -80 0 feedthrough
rlabel pdiffusion 304 -80 304 -80 0 feedthrough
rlabel pdiffusion 311 -80 311 -80 0 feedthrough
rlabel pdiffusion 318 -80 318 -80 0 feedthrough
rlabel pdiffusion 325 -80 325 -80 0 feedthrough
rlabel pdiffusion 332 -80 332 -80 0 feedthrough
rlabel pdiffusion 339 -80 339 -80 0 feedthrough
rlabel pdiffusion 346 -80 346 -80 0 feedthrough
rlabel pdiffusion 353 -80 353 -80 0 cellNo=110
rlabel pdiffusion 360 -80 360 -80 0 feedthrough
rlabel pdiffusion 367 -80 367 -80 0 feedthrough
rlabel pdiffusion 374 -80 374 -80 0 feedthrough
rlabel pdiffusion 381 -80 381 -80 0 feedthrough
rlabel pdiffusion 388 -80 388 -80 0 feedthrough
rlabel pdiffusion 395 -80 395 -80 0 feedthrough
rlabel pdiffusion 402 -80 402 -80 0 feedthrough
rlabel pdiffusion 409 -80 409 -80 0 feedthrough
rlabel pdiffusion 430 -80 430 -80 0 cellNo=316
rlabel pdiffusion 3 -125 3 -125 0 cellNo=8
rlabel pdiffusion 10 -125 10 -125 0 cellNo=725
rlabel pdiffusion 17 -125 17 -125 0 cellNo=151
rlabel pdiffusion 24 -125 24 -125 0 cellNo=245
rlabel pdiffusion 31 -125 31 -125 0 cellNo=315
rlabel pdiffusion 38 -125 38 -125 0 cellNo=761
rlabel pdiffusion 45 -125 45 -125 0 cellNo=464
rlabel pdiffusion 52 -125 52 -125 0 cellNo=180
rlabel pdiffusion 59 -125 59 -125 0 feedthrough
rlabel pdiffusion 66 -125 66 -125 0 cellNo=714
rlabel pdiffusion 80 -125 80 -125 0 feedthrough
rlabel pdiffusion 87 -125 87 -125 0 feedthrough
rlabel pdiffusion 94 -125 94 -125 0 feedthrough
rlabel pdiffusion 101 -125 101 -125 0 cellNo=844
rlabel pdiffusion 108 -125 108 -125 0 feedthrough
rlabel pdiffusion 115 -125 115 -125 0 cellNo=660
rlabel pdiffusion 122 -125 122 -125 0 feedthrough
rlabel pdiffusion 129 -125 129 -125 0 cellNo=548
rlabel pdiffusion 136 -125 136 -125 0 cellNo=195
rlabel pdiffusion 143 -125 143 -125 0 cellNo=409
rlabel pdiffusion 150 -125 150 -125 0 feedthrough
rlabel pdiffusion 157 -125 157 -125 0 cellNo=234
rlabel pdiffusion 164 -125 164 -125 0 cellNo=484
rlabel pdiffusion 171 -125 171 -125 0 feedthrough
rlabel pdiffusion 178 -125 178 -125 0 feedthrough
rlabel pdiffusion 185 -125 185 -125 0 cellNo=854
rlabel pdiffusion 192 -125 192 -125 0 feedthrough
rlabel pdiffusion 199 -125 199 -125 0 cellNo=499
rlabel pdiffusion 206 -125 206 -125 0 feedthrough
rlabel pdiffusion 213 -125 213 -125 0 cellNo=386
rlabel pdiffusion 220 -125 220 -125 0 cellNo=641
rlabel pdiffusion 227 -125 227 -125 0 feedthrough
rlabel pdiffusion 234 -125 234 -125 0 cellNo=888
rlabel pdiffusion 241 -125 241 -125 0 cellNo=425
rlabel pdiffusion 248 -125 248 -125 0 cellNo=517
rlabel pdiffusion 255 -125 255 -125 0 feedthrough
rlabel pdiffusion 262 -125 262 -125 0 cellNo=703
rlabel pdiffusion 269 -125 269 -125 0 cellNo=52
rlabel pdiffusion 276 -125 276 -125 0 cellNo=184
rlabel pdiffusion 283 -125 283 -125 0 feedthrough
rlabel pdiffusion 290 -125 290 -125 0 feedthrough
rlabel pdiffusion 297 -125 297 -125 0 feedthrough
rlabel pdiffusion 304 -125 304 -125 0 feedthrough
rlabel pdiffusion 311 -125 311 -125 0 cellNo=921
rlabel pdiffusion 318 -125 318 -125 0 feedthrough
rlabel pdiffusion 325 -125 325 -125 0 feedthrough
rlabel pdiffusion 332 -125 332 -125 0 feedthrough
rlabel pdiffusion 339 -125 339 -125 0 feedthrough
rlabel pdiffusion 346 -125 346 -125 0 feedthrough
rlabel pdiffusion 353 -125 353 -125 0 feedthrough
rlabel pdiffusion 360 -125 360 -125 0 feedthrough
rlabel pdiffusion 367 -125 367 -125 0 cellNo=112
rlabel pdiffusion 374 -125 374 -125 0 feedthrough
rlabel pdiffusion 381 -125 381 -125 0 cellNo=884
rlabel pdiffusion 388 -125 388 -125 0 feedthrough
rlabel pdiffusion 395 -125 395 -125 0 feedthrough
rlabel pdiffusion 402 -125 402 -125 0 feedthrough
rlabel pdiffusion 409 -125 409 -125 0 feedthrough
rlabel pdiffusion 416 -125 416 -125 0 feedthrough
rlabel pdiffusion 423 -125 423 -125 0 feedthrough
rlabel pdiffusion 430 -125 430 -125 0 feedthrough
rlabel pdiffusion 437 -125 437 -125 0 cellNo=865
rlabel pdiffusion 444 -125 444 -125 0 feedthrough
rlabel pdiffusion 451 -125 451 -125 0 cellNo=300
rlabel pdiffusion 3 -178 3 -178 0 cellNo=68
rlabel pdiffusion 10 -178 10 -178 0 cellNo=473
rlabel pdiffusion 17 -178 17 -178 0 cellNo=109
rlabel pdiffusion 24 -178 24 -178 0 cellNo=294
rlabel pdiffusion 31 -178 31 -178 0 cellNo=947
rlabel pdiffusion 38 -178 38 -178 0 feedthrough
rlabel pdiffusion 45 -178 45 -178 0 feedthrough
rlabel pdiffusion 52 -178 52 -178 0 feedthrough
rlabel pdiffusion 59 -178 59 -178 0 feedthrough
rlabel pdiffusion 66 -178 66 -178 0 cellNo=254
rlabel pdiffusion 73 -178 73 -178 0 feedthrough
rlabel pdiffusion 80 -178 80 -178 0 feedthrough
rlabel pdiffusion 87 -178 87 -178 0 cellNo=426
rlabel pdiffusion 94 -178 94 -178 0 cellNo=429
rlabel pdiffusion 101 -178 101 -178 0 feedthrough
rlabel pdiffusion 108 -178 108 -178 0 cellNo=965
rlabel pdiffusion 115 -178 115 -178 0 feedthrough
rlabel pdiffusion 122 -178 122 -178 0 cellNo=671
rlabel pdiffusion 129 -178 129 -178 0 feedthrough
rlabel pdiffusion 136 -178 136 -178 0 cellNo=4
rlabel pdiffusion 143 -178 143 -178 0 cellNo=144
rlabel pdiffusion 150 -178 150 -178 0 cellNo=393
rlabel pdiffusion 157 -178 157 -178 0 feedthrough
rlabel pdiffusion 164 -178 164 -178 0 cellNo=775
rlabel pdiffusion 171 -178 171 -178 0 feedthrough
rlabel pdiffusion 178 -178 178 -178 0 cellNo=646
rlabel pdiffusion 185 -178 185 -178 0 cellNo=875
rlabel pdiffusion 192 -178 192 -178 0 feedthrough
rlabel pdiffusion 199 -178 199 -178 0 feedthrough
rlabel pdiffusion 206 -178 206 -178 0 cellNo=65
rlabel pdiffusion 213 -178 213 -178 0 cellNo=513
rlabel pdiffusion 220 -178 220 -178 0 feedthrough
rlabel pdiffusion 227 -178 227 -178 0 feedthrough
rlabel pdiffusion 234 -178 234 -178 0 cellNo=24
rlabel pdiffusion 241 -178 241 -178 0 cellNo=659
rlabel pdiffusion 248 -178 248 -178 0 feedthrough
rlabel pdiffusion 255 -178 255 -178 0 cellNo=587
rlabel pdiffusion 262 -178 262 -178 0 feedthrough
rlabel pdiffusion 269 -178 269 -178 0 feedthrough
rlabel pdiffusion 276 -178 276 -178 0 cellNo=406
rlabel pdiffusion 283 -178 283 -178 0 cellNo=268
rlabel pdiffusion 290 -178 290 -178 0 cellNo=384
rlabel pdiffusion 297 -178 297 -178 0 cellNo=799
rlabel pdiffusion 304 -178 304 -178 0 cellNo=770
rlabel pdiffusion 311 -178 311 -178 0 cellNo=687
rlabel pdiffusion 318 -178 318 -178 0 cellNo=845
rlabel pdiffusion 325 -178 325 -178 0 feedthrough
rlabel pdiffusion 332 -178 332 -178 0 cellNo=102
rlabel pdiffusion 339 -178 339 -178 0 feedthrough
rlabel pdiffusion 346 -178 346 -178 0 feedthrough
rlabel pdiffusion 353 -178 353 -178 0 feedthrough
rlabel pdiffusion 360 -178 360 -178 0 feedthrough
rlabel pdiffusion 367 -178 367 -178 0 feedthrough
rlabel pdiffusion 374 -178 374 -178 0 feedthrough
rlabel pdiffusion 381 -178 381 -178 0 feedthrough
rlabel pdiffusion 388 -178 388 -178 0 feedthrough
rlabel pdiffusion 395 -178 395 -178 0 feedthrough
rlabel pdiffusion 402 -178 402 -178 0 feedthrough
rlabel pdiffusion 409 -178 409 -178 0 feedthrough
rlabel pdiffusion 416 -178 416 -178 0 feedthrough
rlabel pdiffusion 430 -178 430 -178 0 feedthrough
rlabel pdiffusion 437 -178 437 -178 0 feedthrough
rlabel pdiffusion 444 -178 444 -178 0 feedthrough
rlabel pdiffusion 451 -178 451 -178 0 feedthrough
rlabel pdiffusion 458 -178 458 -178 0 feedthrough
rlabel pdiffusion 465 -178 465 -178 0 feedthrough
rlabel pdiffusion 472 -178 472 -178 0 feedthrough
rlabel pdiffusion 479 -178 479 -178 0 cellNo=550
rlabel pdiffusion 486 -178 486 -178 0 feedthrough
rlabel pdiffusion 493 -178 493 -178 0 feedthrough
rlabel pdiffusion 549 -178 549 -178 0 cellNo=44
rlabel pdiffusion 3 -235 3 -235 0 cellNo=101
rlabel pdiffusion 17 -235 17 -235 0 feedthrough
rlabel pdiffusion 24 -235 24 -235 0 cellNo=877
rlabel pdiffusion 31 -235 31 -235 0 feedthrough
rlabel pdiffusion 38 -235 38 -235 0 cellNo=575
rlabel pdiffusion 45 -235 45 -235 0 cellNo=161
rlabel pdiffusion 59 -235 59 -235 0 cellNo=200
rlabel pdiffusion 66 -235 66 -235 0 cellNo=117
rlabel pdiffusion 80 -235 80 -235 0 cellNo=707
rlabel pdiffusion 87 -235 87 -235 0 cellNo=787
rlabel pdiffusion 94 -235 94 -235 0 feedthrough
rlabel pdiffusion 101 -235 101 -235 0 cellNo=174
rlabel pdiffusion 108 -235 108 -235 0 feedthrough
rlabel pdiffusion 115 -235 115 -235 0 feedthrough
rlabel pdiffusion 122 -235 122 -235 0 cellNo=627
rlabel pdiffusion 129 -235 129 -235 0 feedthrough
rlabel pdiffusion 136 -235 136 -235 0 feedthrough
rlabel pdiffusion 143 -235 143 -235 0 cellNo=90
rlabel pdiffusion 150 -235 150 -235 0 cellNo=541
rlabel pdiffusion 157 -235 157 -235 0 cellNo=134
rlabel pdiffusion 164 -235 164 -235 0 cellNo=767
rlabel pdiffusion 171 -235 171 -235 0 feedthrough
rlabel pdiffusion 178 -235 178 -235 0 feedthrough
rlabel pdiffusion 185 -235 185 -235 0 feedthrough
rlabel pdiffusion 192 -235 192 -235 0 feedthrough
rlabel pdiffusion 199 -235 199 -235 0 feedthrough
rlabel pdiffusion 206 -235 206 -235 0 feedthrough
rlabel pdiffusion 213 -235 213 -235 0 cellNo=137
rlabel pdiffusion 220 -235 220 -235 0 cellNo=382
rlabel pdiffusion 227 -235 227 -235 0 feedthrough
rlabel pdiffusion 234 -235 234 -235 0 feedthrough
rlabel pdiffusion 241 -235 241 -235 0 cellNo=595
rlabel pdiffusion 248 -235 248 -235 0 feedthrough
rlabel pdiffusion 255 -235 255 -235 0 cellNo=96
rlabel pdiffusion 262 -235 262 -235 0 feedthrough
rlabel pdiffusion 269 -235 269 -235 0 feedthrough
rlabel pdiffusion 276 -235 276 -235 0 feedthrough
rlabel pdiffusion 283 -235 283 -235 0 cellNo=396
rlabel pdiffusion 290 -235 290 -235 0 feedthrough
rlabel pdiffusion 304 -235 304 -235 0 feedthrough
rlabel pdiffusion 311 -235 311 -235 0 cellNo=768
rlabel pdiffusion 318 -235 318 -235 0 feedthrough
rlabel pdiffusion 325 -235 325 -235 0 cellNo=992
rlabel pdiffusion 332 -235 332 -235 0 feedthrough
rlabel pdiffusion 339 -235 339 -235 0 cellNo=891
rlabel pdiffusion 346 -235 346 -235 0 feedthrough
rlabel pdiffusion 353 -235 353 -235 0 cellNo=131
rlabel pdiffusion 360 -235 360 -235 0 cellNo=459
rlabel pdiffusion 367 -235 367 -235 0 feedthrough
rlabel pdiffusion 374 -235 374 -235 0 feedthrough
rlabel pdiffusion 381 -235 381 -235 0 feedthrough
rlabel pdiffusion 388 -235 388 -235 0 feedthrough
rlabel pdiffusion 395 -235 395 -235 0 feedthrough
rlabel pdiffusion 402 -235 402 -235 0 feedthrough
rlabel pdiffusion 409 -235 409 -235 0 feedthrough
rlabel pdiffusion 416 -235 416 -235 0 feedthrough
rlabel pdiffusion 423 -235 423 -235 0 feedthrough
rlabel pdiffusion 430 -235 430 -235 0 feedthrough
rlabel pdiffusion 437 -235 437 -235 0 feedthrough
rlabel pdiffusion 444 -235 444 -235 0 feedthrough
rlabel pdiffusion 451 -235 451 -235 0 feedthrough
rlabel pdiffusion 458 -235 458 -235 0 feedthrough
rlabel pdiffusion 465 -235 465 -235 0 feedthrough
rlabel pdiffusion 472 -235 472 -235 0 feedthrough
rlabel pdiffusion 479 -235 479 -235 0 feedthrough
rlabel pdiffusion 486 -235 486 -235 0 feedthrough
rlabel pdiffusion 493 -235 493 -235 0 feedthrough
rlabel pdiffusion 500 -235 500 -235 0 feedthrough
rlabel pdiffusion 507 -235 507 -235 0 feedthrough
rlabel pdiffusion 514 -235 514 -235 0 feedthrough
rlabel pdiffusion 521 -235 521 -235 0 cellNo=551
rlabel pdiffusion 528 -235 528 -235 0 feedthrough
rlabel pdiffusion 535 -235 535 -235 0 feedthrough
rlabel pdiffusion 542 -235 542 -235 0 cellNo=226
rlabel pdiffusion 549 -235 549 -235 0 cellNo=182
rlabel pdiffusion 556 -235 556 -235 0 cellNo=37
rlabel pdiffusion 563 -235 563 -235 0 cellNo=635
rlabel pdiffusion 584 -235 584 -235 0 cellNo=979
rlabel pdiffusion 640 -235 640 -235 0 feedthrough
rlabel pdiffusion 654 -235 654 -235 0 cellNo=59
rlabel pdiffusion 3 -292 3 -292 0 cellNo=438
rlabel pdiffusion 10 -292 10 -292 0 cellNo=485
rlabel pdiffusion 17 -292 17 -292 0 cellNo=807
rlabel pdiffusion 24 -292 24 -292 0 cellNo=40
rlabel pdiffusion 31 -292 31 -292 0 feedthrough
rlabel pdiffusion 38 -292 38 -292 0 cellNo=237
rlabel pdiffusion 45 -292 45 -292 0 feedthrough
rlabel pdiffusion 52 -292 52 -292 0 cellNo=157
rlabel pdiffusion 59 -292 59 -292 0 feedthrough
rlabel pdiffusion 66 -292 66 -292 0 cellNo=15
rlabel pdiffusion 73 -292 73 -292 0 feedthrough
rlabel pdiffusion 80 -292 80 -292 0 cellNo=160
rlabel pdiffusion 87 -292 87 -292 0 feedthrough
rlabel pdiffusion 94 -292 94 -292 0 feedthrough
rlabel pdiffusion 101 -292 101 -292 0 feedthrough
rlabel pdiffusion 108 -292 108 -292 0 feedthrough
rlabel pdiffusion 115 -292 115 -292 0 feedthrough
rlabel pdiffusion 122 -292 122 -292 0 cellNo=107
rlabel pdiffusion 129 -292 129 -292 0 feedthrough
rlabel pdiffusion 136 -292 136 -292 0 feedthrough
rlabel pdiffusion 143 -292 143 -292 0 cellNo=545
rlabel pdiffusion 150 -292 150 -292 0 cellNo=662
rlabel pdiffusion 157 -292 157 -292 0 feedthrough
rlabel pdiffusion 164 -292 164 -292 0 cellNo=652
rlabel pdiffusion 171 -292 171 -292 0 feedthrough
rlabel pdiffusion 178 -292 178 -292 0 cellNo=383
rlabel pdiffusion 185 -292 185 -292 0 feedthrough
rlabel pdiffusion 192 -292 192 -292 0 cellNo=495
rlabel pdiffusion 199 -292 199 -292 0 feedthrough
rlabel pdiffusion 206 -292 206 -292 0 cellNo=792
rlabel pdiffusion 213 -292 213 -292 0 cellNo=765
rlabel pdiffusion 220 -292 220 -292 0 cellNo=713
rlabel pdiffusion 227 -292 227 -292 0 feedthrough
rlabel pdiffusion 234 -292 234 -292 0 feedthrough
rlabel pdiffusion 241 -292 241 -292 0 feedthrough
rlabel pdiffusion 248 -292 248 -292 0 cellNo=67
rlabel pdiffusion 255 -292 255 -292 0 cellNo=148
rlabel pdiffusion 262 -292 262 -292 0 feedthrough
rlabel pdiffusion 269 -292 269 -292 0 feedthrough
rlabel pdiffusion 276 -292 276 -292 0 cellNo=346
rlabel pdiffusion 283 -292 283 -292 0 cellNo=910
rlabel pdiffusion 290 -292 290 -292 0 feedthrough
rlabel pdiffusion 297 -292 297 -292 0 cellNo=695
rlabel pdiffusion 304 -292 304 -292 0 feedthrough
rlabel pdiffusion 311 -292 311 -292 0 cellNo=566
rlabel pdiffusion 318 -292 318 -292 0 cellNo=443
rlabel pdiffusion 325 -292 325 -292 0 feedthrough
rlabel pdiffusion 332 -292 332 -292 0 cellNo=304
rlabel pdiffusion 339 -292 339 -292 0 cellNo=896
rlabel pdiffusion 346 -292 346 -292 0 feedthrough
rlabel pdiffusion 353 -292 353 -292 0 feedthrough
rlabel pdiffusion 360 -292 360 -292 0 cellNo=325
rlabel pdiffusion 367 -292 367 -292 0 feedthrough
rlabel pdiffusion 374 -292 374 -292 0 feedthrough
rlabel pdiffusion 381 -292 381 -292 0 feedthrough
rlabel pdiffusion 388 -292 388 -292 0 cellNo=433
rlabel pdiffusion 395 -292 395 -292 0 feedthrough
rlabel pdiffusion 402 -292 402 -292 0 feedthrough
rlabel pdiffusion 409 -292 409 -292 0 feedthrough
rlabel pdiffusion 416 -292 416 -292 0 feedthrough
rlabel pdiffusion 423 -292 423 -292 0 feedthrough
rlabel pdiffusion 430 -292 430 -292 0 feedthrough
rlabel pdiffusion 437 -292 437 -292 0 cellNo=201
rlabel pdiffusion 444 -292 444 -292 0 feedthrough
rlabel pdiffusion 451 -292 451 -292 0 feedthrough
rlabel pdiffusion 458 -292 458 -292 0 feedthrough
rlabel pdiffusion 465 -292 465 -292 0 feedthrough
rlabel pdiffusion 472 -292 472 -292 0 feedthrough
rlabel pdiffusion 479 -292 479 -292 0 cellNo=242
rlabel pdiffusion 486 -292 486 -292 0 feedthrough
rlabel pdiffusion 493 -292 493 -292 0 feedthrough
rlabel pdiffusion 500 -292 500 -292 0 feedthrough
rlabel pdiffusion 507 -292 507 -292 0 feedthrough
rlabel pdiffusion 514 -292 514 -292 0 feedthrough
rlabel pdiffusion 521 -292 521 -292 0 feedthrough
rlabel pdiffusion 528 -292 528 -292 0 feedthrough
rlabel pdiffusion 535 -292 535 -292 0 feedthrough
rlabel pdiffusion 542 -292 542 -292 0 feedthrough
rlabel pdiffusion 549 -292 549 -292 0 feedthrough
rlabel pdiffusion 556 -292 556 -292 0 feedthrough
rlabel pdiffusion 563 -292 563 -292 0 feedthrough
rlabel pdiffusion 570 -292 570 -292 0 feedthrough
rlabel pdiffusion 577 -292 577 -292 0 feedthrough
rlabel pdiffusion 584 -292 584 -292 0 feedthrough
rlabel pdiffusion 591 -292 591 -292 0 feedthrough
rlabel pdiffusion 598 -292 598 -292 0 feedthrough
rlabel pdiffusion 605 -292 605 -292 0 feedthrough
rlabel pdiffusion 612 -292 612 -292 0 feedthrough
rlabel pdiffusion 619 -292 619 -292 0 feedthrough
rlabel pdiffusion 626 -292 626 -292 0 feedthrough
rlabel pdiffusion 633 -292 633 -292 0 feedthrough
rlabel pdiffusion 654 -292 654 -292 0 feedthrough
rlabel pdiffusion 661 -292 661 -292 0 feedthrough
rlabel pdiffusion 3 -361 3 -361 0 cellNo=582
rlabel pdiffusion 10 -361 10 -361 0 feedthrough
rlabel pdiffusion 17 -361 17 -361 0 cellNo=643
rlabel pdiffusion 24 -361 24 -361 0 feedthrough
rlabel pdiffusion 31 -361 31 -361 0 feedthrough
rlabel pdiffusion 45 -361 45 -361 0 cellNo=670
rlabel pdiffusion 52 -361 52 -361 0 cellNo=860
rlabel pdiffusion 59 -361 59 -361 0 feedthrough
rlabel pdiffusion 73 -361 73 -361 0 feedthrough
rlabel pdiffusion 80 -361 80 -361 0 feedthrough
rlabel pdiffusion 87 -361 87 -361 0 feedthrough
rlabel pdiffusion 94 -361 94 -361 0 feedthrough
rlabel pdiffusion 101 -361 101 -361 0 cellNo=7
rlabel pdiffusion 108 -361 108 -361 0 cellNo=915
rlabel pdiffusion 115 -361 115 -361 0 cellNo=233
rlabel pdiffusion 122 -361 122 -361 0 cellNo=191
rlabel pdiffusion 129 -361 129 -361 0 feedthrough
rlabel pdiffusion 136 -361 136 -361 0 feedthrough
rlabel pdiffusion 143 -361 143 -361 0 feedthrough
rlabel pdiffusion 150 -361 150 -361 0 cellNo=153
rlabel pdiffusion 157 -361 157 -361 0 cellNo=238
rlabel pdiffusion 164 -361 164 -361 0 cellNo=804
rlabel pdiffusion 171 -361 171 -361 0 cellNo=380
rlabel pdiffusion 178 -361 178 -361 0 cellNo=119
rlabel pdiffusion 185 -361 185 -361 0 cellNo=717
rlabel pdiffusion 192 -361 192 -361 0 cellNo=166
rlabel pdiffusion 199 -361 199 -361 0 feedthrough
rlabel pdiffusion 206 -361 206 -361 0 cellNo=873
rlabel pdiffusion 213 -361 213 -361 0 feedthrough
rlabel pdiffusion 220 -361 220 -361 0 cellNo=239
rlabel pdiffusion 227 -361 227 -361 0 feedthrough
rlabel pdiffusion 234 -361 234 -361 0 feedthrough
rlabel pdiffusion 241 -361 241 -361 0 feedthrough
rlabel pdiffusion 248 -361 248 -361 0 feedthrough
rlabel pdiffusion 255 -361 255 -361 0 feedthrough
rlabel pdiffusion 262 -361 262 -361 0 feedthrough
rlabel pdiffusion 269 -361 269 -361 0 feedthrough
rlabel pdiffusion 276 -361 276 -361 0 cellNo=430
rlabel pdiffusion 283 -361 283 -361 0 cellNo=882
rlabel pdiffusion 290 -361 290 -361 0 feedthrough
rlabel pdiffusion 297 -361 297 -361 0 cellNo=223
rlabel pdiffusion 304 -361 304 -361 0 feedthrough
rlabel pdiffusion 311 -361 311 -361 0 feedthrough
rlabel pdiffusion 318 -361 318 -361 0 feedthrough
rlabel pdiffusion 325 -361 325 -361 0 cellNo=547
rlabel pdiffusion 332 -361 332 -361 0 feedthrough
rlabel pdiffusion 339 -361 339 -361 0 feedthrough
rlabel pdiffusion 346 -361 346 -361 0 feedthrough
rlabel pdiffusion 353 -361 353 -361 0 cellNo=279
rlabel pdiffusion 360 -361 360 -361 0 cellNo=781
rlabel pdiffusion 367 -361 367 -361 0 cellNo=310
rlabel pdiffusion 374 -361 374 -361 0 feedthrough
rlabel pdiffusion 381 -361 381 -361 0 cellNo=176
rlabel pdiffusion 388 -361 388 -361 0 cellNo=319
rlabel pdiffusion 395 -361 395 -361 0 feedthrough
rlabel pdiffusion 402 -361 402 -361 0 feedthrough
rlabel pdiffusion 409 -361 409 -361 0 feedthrough
rlabel pdiffusion 416 -361 416 -361 0 feedthrough
rlabel pdiffusion 423 -361 423 -361 0 feedthrough
rlabel pdiffusion 430 -361 430 -361 0 cellNo=851
rlabel pdiffusion 437 -361 437 -361 0 feedthrough
rlabel pdiffusion 444 -361 444 -361 0 feedthrough
rlabel pdiffusion 451 -361 451 -361 0 cellNo=574
rlabel pdiffusion 458 -361 458 -361 0 feedthrough
rlabel pdiffusion 465 -361 465 -361 0 feedthrough
rlabel pdiffusion 472 -361 472 -361 0 feedthrough
rlabel pdiffusion 479 -361 479 -361 0 feedthrough
rlabel pdiffusion 486 -361 486 -361 0 feedthrough
rlabel pdiffusion 493 -361 493 -361 0 feedthrough
rlabel pdiffusion 507 -361 507 -361 0 feedthrough
rlabel pdiffusion 514 -361 514 -361 0 feedthrough
rlabel pdiffusion 521 -361 521 -361 0 feedthrough
rlabel pdiffusion 528 -361 528 -361 0 feedthrough
rlabel pdiffusion 535 -361 535 -361 0 feedthrough
rlabel pdiffusion 542 -361 542 -361 0 feedthrough
rlabel pdiffusion 549 -361 549 -361 0 feedthrough
rlabel pdiffusion 556 -361 556 -361 0 feedthrough
rlabel pdiffusion 563 -361 563 -361 0 feedthrough
rlabel pdiffusion 570 -361 570 -361 0 feedthrough
rlabel pdiffusion 577 -361 577 -361 0 feedthrough
rlabel pdiffusion 584 -361 584 -361 0 feedthrough
rlabel pdiffusion 591 -361 591 -361 0 feedthrough
rlabel pdiffusion 598 -361 598 -361 0 feedthrough
rlabel pdiffusion 605 -361 605 -361 0 feedthrough
rlabel pdiffusion 612 -361 612 -361 0 feedthrough
rlabel pdiffusion 619 -361 619 -361 0 cellNo=584
rlabel pdiffusion 654 -361 654 -361 0 cellNo=836
rlabel pdiffusion 661 -361 661 -361 0 feedthrough
rlabel pdiffusion 668 -361 668 -361 0 cellNo=177
rlabel pdiffusion 675 -361 675 -361 0 feedthrough
rlabel pdiffusion 3 -428 3 -428 0 cellNo=603
rlabel pdiffusion 10 -428 10 -428 0 cellNo=633
rlabel pdiffusion 17 -428 17 -428 0 feedthrough
rlabel pdiffusion 31 -428 31 -428 0 cellNo=518
rlabel pdiffusion 38 -428 38 -428 0 cellNo=750
rlabel pdiffusion 45 -428 45 -428 0 feedthrough
rlabel pdiffusion 52 -428 52 -428 0 feedthrough
rlabel pdiffusion 59 -428 59 -428 0 cellNo=598
rlabel pdiffusion 66 -428 66 -428 0 feedthrough
rlabel pdiffusion 73 -428 73 -428 0 feedthrough
rlabel pdiffusion 80 -428 80 -428 0 cellNo=210
rlabel pdiffusion 87 -428 87 -428 0 feedthrough
rlabel pdiffusion 94 -428 94 -428 0 feedthrough
rlabel pdiffusion 101 -428 101 -428 0 feedthrough
rlabel pdiffusion 108 -428 108 -428 0 feedthrough
rlabel pdiffusion 115 -428 115 -428 0 cellNo=715
rlabel pdiffusion 122 -428 122 -428 0 feedthrough
rlabel pdiffusion 129 -428 129 -428 0 feedthrough
rlabel pdiffusion 136 -428 136 -428 0 cellNo=690
rlabel pdiffusion 143 -428 143 -428 0 feedthrough
rlabel pdiffusion 150 -428 150 -428 0 feedthrough
rlabel pdiffusion 157 -428 157 -428 0 feedthrough
rlabel pdiffusion 164 -428 164 -428 0 cellNo=813
rlabel pdiffusion 171 -428 171 -428 0 cellNo=348
rlabel pdiffusion 178 -428 178 -428 0 cellNo=442
rlabel pdiffusion 185 -428 185 -428 0 feedthrough
rlabel pdiffusion 192 -428 192 -428 0 cellNo=378
rlabel pdiffusion 199 -428 199 -428 0 cellNo=190
rlabel pdiffusion 206 -428 206 -428 0 cellNo=168
rlabel pdiffusion 213 -428 213 -428 0 cellNo=199
rlabel pdiffusion 220 -428 220 -428 0 cellNo=252
rlabel pdiffusion 227 -428 227 -428 0 cellNo=563
rlabel pdiffusion 234 -428 234 -428 0 cellNo=493
rlabel pdiffusion 241 -428 241 -428 0 feedthrough
rlabel pdiffusion 248 -428 248 -428 0 cellNo=371
rlabel pdiffusion 255 -428 255 -428 0 cellNo=922
rlabel pdiffusion 262 -428 262 -428 0 cellNo=502
rlabel pdiffusion 269 -428 269 -428 0 feedthrough
rlabel pdiffusion 276 -428 276 -428 0 feedthrough
rlabel pdiffusion 283 -428 283 -428 0 cellNo=620
rlabel pdiffusion 290 -428 290 -428 0 feedthrough
rlabel pdiffusion 297 -428 297 -428 0 feedthrough
rlabel pdiffusion 304 -428 304 -428 0 feedthrough
rlabel pdiffusion 311 -428 311 -428 0 cellNo=140
rlabel pdiffusion 318 -428 318 -428 0 cellNo=116
rlabel pdiffusion 325 -428 325 -428 0 cellNo=220
rlabel pdiffusion 332 -428 332 -428 0 feedthrough
rlabel pdiffusion 339 -428 339 -428 0 cellNo=66
rlabel pdiffusion 346 -428 346 -428 0 feedthrough
rlabel pdiffusion 353 -428 353 -428 0 feedthrough
rlabel pdiffusion 360 -428 360 -428 0 cellNo=593
rlabel pdiffusion 367 -428 367 -428 0 feedthrough
rlabel pdiffusion 374 -428 374 -428 0 feedthrough
rlabel pdiffusion 381 -428 381 -428 0 cellNo=542
rlabel pdiffusion 388 -428 388 -428 0 cellNo=262
rlabel pdiffusion 395 -428 395 -428 0 feedthrough
rlabel pdiffusion 402 -428 402 -428 0 feedthrough
rlabel pdiffusion 409 -428 409 -428 0 feedthrough
rlabel pdiffusion 416 -428 416 -428 0 feedthrough
rlabel pdiffusion 423 -428 423 -428 0 feedthrough
rlabel pdiffusion 430 -428 430 -428 0 feedthrough
rlabel pdiffusion 437 -428 437 -428 0 feedthrough
rlabel pdiffusion 444 -428 444 -428 0 feedthrough
rlabel pdiffusion 451 -428 451 -428 0 feedthrough
rlabel pdiffusion 458 -428 458 -428 0 feedthrough
rlabel pdiffusion 465 -428 465 -428 0 feedthrough
rlabel pdiffusion 472 -428 472 -428 0 cellNo=617
rlabel pdiffusion 479 -428 479 -428 0 cellNo=454
rlabel pdiffusion 486 -428 486 -428 0 feedthrough
rlabel pdiffusion 493 -428 493 -428 0 feedthrough
rlabel pdiffusion 500 -428 500 -428 0 feedthrough
rlabel pdiffusion 507 -428 507 -428 0 feedthrough
rlabel pdiffusion 514 -428 514 -428 0 feedthrough
rlabel pdiffusion 521 -428 521 -428 0 feedthrough
rlabel pdiffusion 528 -428 528 -428 0 feedthrough
rlabel pdiffusion 535 -428 535 -428 0 feedthrough
rlabel pdiffusion 542 -428 542 -428 0 feedthrough
rlabel pdiffusion 549 -428 549 -428 0 feedthrough
rlabel pdiffusion 556 -428 556 -428 0 feedthrough
rlabel pdiffusion 563 -428 563 -428 0 feedthrough
rlabel pdiffusion 570 -428 570 -428 0 feedthrough
rlabel pdiffusion 577 -428 577 -428 0 feedthrough
rlabel pdiffusion 584 -428 584 -428 0 feedthrough
rlabel pdiffusion 591 -428 591 -428 0 feedthrough
rlabel pdiffusion 598 -428 598 -428 0 feedthrough
rlabel pdiffusion 605 -428 605 -428 0 feedthrough
rlabel pdiffusion 612 -428 612 -428 0 feedthrough
rlabel pdiffusion 619 -428 619 -428 0 feedthrough
rlabel pdiffusion 626 -428 626 -428 0 feedthrough
rlabel pdiffusion 633 -428 633 -428 0 feedthrough
rlabel pdiffusion 640 -428 640 -428 0 feedthrough
rlabel pdiffusion 647 -428 647 -428 0 feedthrough
rlabel pdiffusion 654 -428 654 -428 0 feedthrough
rlabel pdiffusion 661 -428 661 -428 0 feedthrough
rlabel pdiffusion 668 -428 668 -428 0 feedthrough
rlabel pdiffusion 675 -428 675 -428 0 cellNo=449
rlabel pdiffusion 682 -428 682 -428 0 feedthrough
rlabel pdiffusion 3 -515 3 -515 0 cellNo=388
rlabel pdiffusion 10 -515 10 -515 0 cellNo=650
rlabel pdiffusion 17 -515 17 -515 0 cellNo=498
rlabel pdiffusion 24 -515 24 -515 0 cellNo=264
rlabel pdiffusion 31 -515 31 -515 0 cellNo=533
rlabel pdiffusion 38 -515 38 -515 0 cellNo=415
rlabel pdiffusion 45 -515 45 -515 0 feedthrough
rlabel pdiffusion 52 -515 52 -515 0 cellNo=528
rlabel pdiffusion 59 -515 59 -515 0 feedthrough
rlabel pdiffusion 66 -515 66 -515 0 feedthrough
rlabel pdiffusion 73 -515 73 -515 0 feedthrough
rlabel pdiffusion 80 -515 80 -515 0 feedthrough
rlabel pdiffusion 87 -515 87 -515 0 cellNo=207
rlabel pdiffusion 94 -515 94 -515 0 feedthrough
rlabel pdiffusion 101 -515 101 -515 0 feedthrough
rlabel pdiffusion 108 -515 108 -515 0 cellNo=317
rlabel pdiffusion 115 -515 115 -515 0 feedthrough
rlabel pdiffusion 122 -515 122 -515 0 cellNo=793
rlabel pdiffusion 129 -515 129 -515 0 feedthrough
rlabel pdiffusion 136 -515 136 -515 0 feedthrough
rlabel pdiffusion 143 -515 143 -515 0 cellNo=534
rlabel pdiffusion 150 -515 150 -515 0 feedthrough
rlabel pdiffusion 157 -515 157 -515 0 feedthrough
rlabel pdiffusion 164 -515 164 -515 0 feedthrough
rlabel pdiffusion 171 -515 171 -515 0 cellNo=973
rlabel pdiffusion 178 -515 178 -515 0 feedthrough
rlabel pdiffusion 185 -515 185 -515 0 feedthrough
rlabel pdiffusion 192 -515 192 -515 0 feedthrough
rlabel pdiffusion 199 -515 199 -515 0 cellNo=613
rlabel pdiffusion 206 -515 206 -515 0 feedthrough
rlabel pdiffusion 213 -515 213 -515 0 cellNo=29
rlabel pdiffusion 220 -515 220 -515 0 cellNo=712
rlabel pdiffusion 227 -515 227 -515 0 cellNo=422
rlabel pdiffusion 234 -515 234 -515 0 feedthrough
rlabel pdiffusion 241 -515 241 -515 0 cellNo=258
rlabel pdiffusion 248 -515 248 -515 0 feedthrough
rlabel pdiffusion 255 -515 255 -515 0 cellNo=601
rlabel pdiffusion 262 -515 262 -515 0 feedthrough
rlabel pdiffusion 269 -515 269 -515 0 cellNo=604
rlabel pdiffusion 276 -515 276 -515 0 cellNo=152
rlabel pdiffusion 283 -515 283 -515 0 cellNo=127
rlabel pdiffusion 290 -515 290 -515 0 feedthrough
rlabel pdiffusion 297 -515 297 -515 0 cellNo=211
rlabel pdiffusion 304 -515 304 -515 0 feedthrough
rlabel pdiffusion 311 -515 311 -515 0 feedthrough
rlabel pdiffusion 318 -515 318 -515 0 cellNo=699
rlabel pdiffusion 325 -515 325 -515 0 cellNo=935
rlabel pdiffusion 332 -515 332 -515 0 feedthrough
rlabel pdiffusion 339 -515 339 -515 0 feedthrough
rlabel pdiffusion 346 -515 346 -515 0 cellNo=323
rlabel pdiffusion 353 -515 353 -515 0 cellNo=326
rlabel pdiffusion 360 -515 360 -515 0 cellNo=763
rlabel pdiffusion 367 -515 367 -515 0 feedthrough
rlabel pdiffusion 374 -515 374 -515 0 feedthrough
rlabel pdiffusion 381 -515 381 -515 0 feedthrough
rlabel pdiffusion 388 -515 388 -515 0 cellNo=375
rlabel pdiffusion 395 -515 395 -515 0 feedthrough
rlabel pdiffusion 402 -515 402 -515 0 cellNo=740
rlabel pdiffusion 409 -515 409 -515 0 feedthrough
rlabel pdiffusion 416 -515 416 -515 0 feedthrough
rlabel pdiffusion 423 -515 423 -515 0 cellNo=365
rlabel pdiffusion 430 -515 430 -515 0 feedthrough
rlabel pdiffusion 437 -515 437 -515 0 cellNo=202
rlabel pdiffusion 444 -515 444 -515 0 feedthrough
rlabel pdiffusion 451 -515 451 -515 0 cellNo=260
rlabel pdiffusion 458 -515 458 -515 0 feedthrough
rlabel pdiffusion 465 -515 465 -515 0 feedthrough
rlabel pdiffusion 472 -515 472 -515 0 feedthrough
rlabel pdiffusion 479 -515 479 -515 0 feedthrough
rlabel pdiffusion 486 -515 486 -515 0 feedthrough
rlabel pdiffusion 493 -515 493 -515 0 feedthrough
rlabel pdiffusion 500 -515 500 -515 0 feedthrough
rlabel pdiffusion 507 -515 507 -515 0 feedthrough
rlabel pdiffusion 514 -515 514 -515 0 feedthrough
rlabel pdiffusion 521 -515 521 -515 0 feedthrough
rlabel pdiffusion 528 -515 528 -515 0 feedthrough
rlabel pdiffusion 535 -515 535 -515 0 feedthrough
rlabel pdiffusion 542 -515 542 -515 0 feedthrough
rlabel pdiffusion 549 -515 549 -515 0 feedthrough
rlabel pdiffusion 556 -515 556 -515 0 feedthrough
rlabel pdiffusion 563 -515 563 -515 0 feedthrough
rlabel pdiffusion 570 -515 570 -515 0 feedthrough
rlabel pdiffusion 577 -515 577 -515 0 feedthrough
rlabel pdiffusion 584 -515 584 -515 0 feedthrough
rlabel pdiffusion 591 -515 591 -515 0 feedthrough
rlabel pdiffusion 598 -515 598 -515 0 feedthrough
rlabel pdiffusion 605 -515 605 -515 0 feedthrough
rlabel pdiffusion 612 -515 612 -515 0 feedthrough
rlabel pdiffusion 619 -515 619 -515 0 feedthrough
rlabel pdiffusion 626 -515 626 -515 0 feedthrough
rlabel pdiffusion 633 -515 633 -515 0 feedthrough
rlabel pdiffusion 640 -515 640 -515 0 feedthrough
rlabel pdiffusion 647 -515 647 -515 0 feedthrough
rlabel pdiffusion 654 -515 654 -515 0 feedthrough
rlabel pdiffusion 661 -515 661 -515 0 feedthrough
rlabel pdiffusion 668 -515 668 -515 0 feedthrough
rlabel pdiffusion 675 -515 675 -515 0 feedthrough
rlabel pdiffusion 682 -515 682 -515 0 feedthrough
rlabel pdiffusion 689 -515 689 -515 0 feedthrough
rlabel pdiffusion 696 -515 696 -515 0 feedthrough
rlabel pdiffusion 703 -515 703 -515 0 feedthrough
rlabel pdiffusion 710 -515 710 -515 0 feedthrough
rlabel pdiffusion 3 -602 3 -602 0 cellNo=444
rlabel pdiffusion 10 -602 10 -602 0 cellNo=467
rlabel pdiffusion 17 -602 17 -602 0 cellNo=328
rlabel pdiffusion 24 -602 24 -602 0 feedthrough
rlabel pdiffusion 31 -602 31 -602 0 feedthrough
rlabel pdiffusion 38 -602 38 -602 0 feedthrough
rlabel pdiffusion 45 -602 45 -602 0 feedthrough
rlabel pdiffusion 52 -602 52 -602 0 cellNo=282
rlabel pdiffusion 59 -602 59 -602 0 feedthrough
rlabel pdiffusion 66 -602 66 -602 0 cellNo=138
rlabel pdiffusion 73 -602 73 -602 0 cellNo=724
rlabel pdiffusion 80 -602 80 -602 0 feedthrough
rlabel pdiffusion 87 -602 87 -602 0 feedthrough
rlabel pdiffusion 94 -602 94 -602 0 feedthrough
rlabel pdiffusion 101 -602 101 -602 0 cellNo=331
rlabel pdiffusion 108 -602 108 -602 0 cellNo=208
rlabel pdiffusion 115 -602 115 -602 0 cellNo=789
rlabel pdiffusion 122 -602 122 -602 0 feedthrough
rlabel pdiffusion 129 -602 129 -602 0 cellNo=823
rlabel pdiffusion 136 -602 136 -602 0 cellNo=594
rlabel pdiffusion 143 -602 143 -602 0 feedthrough
rlabel pdiffusion 150 -602 150 -602 0 feedthrough
rlabel pdiffusion 157 -602 157 -602 0 cellNo=261
rlabel pdiffusion 164 -602 164 -602 0 feedthrough
rlabel pdiffusion 171 -602 171 -602 0 feedthrough
rlabel pdiffusion 178 -602 178 -602 0 feedthrough
rlabel pdiffusion 185 -602 185 -602 0 feedthrough
rlabel pdiffusion 192 -602 192 -602 0 cellNo=121
rlabel pdiffusion 199 -602 199 -602 0 cellNo=150
rlabel pdiffusion 206 -602 206 -602 0 feedthrough
rlabel pdiffusion 213 -602 213 -602 0 cellNo=141
rlabel pdiffusion 220 -602 220 -602 0 cellNo=569
rlabel pdiffusion 227 -602 227 -602 0 feedthrough
rlabel pdiffusion 234 -602 234 -602 0 feedthrough
rlabel pdiffusion 241 -602 241 -602 0 feedthrough
rlabel pdiffusion 248 -602 248 -602 0 feedthrough
rlabel pdiffusion 255 -602 255 -602 0 feedthrough
rlabel pdiffusion 262 -602 262 -602 0 feedthrough
rlabel pdiffusion 269 -602 269 -602 0 feedthrough
rlabel pdiffusion 276 -602 276 -602 0 cellNo=379
rlabel pdiffusion 283 -602 283 -602 0 cellNo=431
rlabel pdiffusion 290 -602 290 -602 0 feedthrough
rlabel pdiffusion 297 -602 297 -602 0 feedthrough
rlabel pdiffusion 304 -602 304 -602 0 cellNo=651
rlabel pdiffusion 311 -602 311 -602 0 feedthrough
rlabel pdiffusion 318 -602 318 -602 0 cellNo=745
rlabel pdiffusion 325 -602 325 -602 0 feedthrough
rlabel pdiffusion 332 -602 332 -602 0 feedthrough
rlabel pdiffusion 339 -602 339 -602 0 cellNo=288
rlabel pdiffusion 346 -602 346 -602 0 cellNo=607
rlabel pdiffusion 353 -602 353 -602 0 feedthrough
rlabel pdiffusion 360 -602 360 -602 0 feedthrough
rlabel pdiffusion 367 -602 367 -602 0 feedthrough
rlabel pdiffusion 374 -602 374 -602 0 cellNo=993
rlabel pdiffusion 381 -602 381 -602 0 feedthrough
rlabel pdiffusion 388 -602 388 -602 0 feedthrough
rlabel pdiffusion 395 -602 395 -602 0 feedthrough
rlabel pdiffusion 402 -602 402 -602 0 feedthrough
rlabel pdiffusion 409 -602 409 -602 0 cellNo=861
rlabel pdiffusion 416 -602 416 -602 0 cellNo=329
rlabel pdiffusion 423 -602 423 -602 0 feedthrough
rlabel pdiffusion 430 -602 430 -602 0 feedthrough
rlabel pdiffusion 437 -602 437 -602 0 cellNo=143
rlabel pdiffusion 444 -602 444 -602 0 cellNo=91
rlabel pdiffusion 451 -602 451 -602 0 feedthrough
rlabel pdiffusion 458 -602 458 -602 0 cellNo=514
rlabel pdiffusion 465 -602 465 -602 0 feedthrough
rlabel pdiffusion 472 -602 472 -602 0 cellNo=723
rlabel pdiffusion 479 -602 479 -602 0 feedthrough
rlabel pdiffusion 486 -602 486 -602 0 feedthrough
rlabel pdiffusion 493 -602 493 -602 0 cellNo=126
rlabel pdiffusion 500 -602 500 -602 0 cellNo=147
rlabel pdiffusion 507 -602 507 -602 0 feedthrough
rlabel pdiffusion 514 -602 514 -602 0 feedthrough
rlabel pdiffusion 521 -602 521 -602 0 feedthrough
rlabel pdiffusion 528 -602 528 -602 0 feedthrough
rlabel pdiffusion 535 -602 535 -602 0 feedthrough
rlabel pdiffusion 542 -602 542 -602 0 feedthrough
rlabel pdiffusion 549 -602 549 -602 0 feedthrough
rlabel pdiffusion 556 -602 556 -602 0 cellNo=62
rlabel pdiffusion 563 -602 563 -602 0 feedthrough
rlabel pdiffusion 570 -602 570 -602 0 feedthrough
rlabel pdiffusion 577 -602 577 -602 0 feedthrough
rlabel pdiffusion 584 -602 584 -602 0 feedthrough
rlabel pdiffusion 591 -602 591 -602 0 feedthrough
rlabel pdiffusion 598 -602 598 -602 0 feedthrough
rlabel pdiffusion 605 -602 605 -602 0 feedthrough
rlabel pdiffusion 612 -602 612 -602 0 feedthrough
rlabel pdiffusion 619 -602 619 -602 0 feedthrough
rlabel pdiffusion 626 -602 626 -602 0 feedthrough
rlabel pdiffusion 633 -602 633 -602 0 feedthrough
rlabel pdiffusion 640 -602 640 -602 0 feedthrough
rlabel pdiffusion 647 -602 647 -602 0 feedthrough
rlabel pdiffusion 654 -602 654 -602 0 feedthrough
rlabel pdiffusion 661 -602 661 -602 0 feedthrough
rlabel pdiffusion 668 -602 668 -602 0 feedthrough
rlabel pdiffusion 675 -602 675 -602 0 feedthrough
rlabel pdiffusion 682 -602 682 -602 0 feedthrough
rlabel pdiffusion 710 -602 710 -602 0 feedthrough
rlabel pdiffusion 3 -681 3 -681 0 cellNo=506
rlabel pdiffusion 10 -681 10 -681 0 cellNo=642
rlabel pdiffusion 17 -681 17 -681 0 cellNo=734
rlabel pdiffusion 24 -681 24 -681 0 cellNo=423
rlabel pdiffusion 31 -681 31 -681 0 cellNo=362
rlabel pdiffusion 38 -681 38 -681 0 feedthrough
rlabel pdiffusion 45 -681 45 -681 0 feedthrough
rlabel pdiffusion 52 -681 52 -681 0 feedthrough
rlabel pdiffusion 59 -681 59 -681 0 cellNo=3
rlabel pdiffusion 66 -681 66 -681 0 feedthrough
rlabel pdiffusion 73 -681 73 -681 0 cellNo=53
rlabel pdiffusion 80 -681 80 -681 0 feedthrough
rlabel pdiffusion 87 -681 87 -681 0 feedthrough
rlabel pdiffusion 94 -681 94 -681 0 feedthrough
rlabel pdiffusion 101 -681 101 -681 0 feedthrough
rlabel pdiffusion 108 -681 108 -681 0 feedthrough
rlabel pdiffusion 115 -681 115 -681 0 feedthrough
rlabel pdiffusion 122 -681 122 -681 0 cellNo=421
rlabel pdiffusion 129 -681 129 -681 0 cellNo=306
rlabel pdiffusion 136 -681 136 -681 0 cellNo=10
rlabel pdiffusion 143 -681 143 -681 0 cellNo=108
rlabel pdiffusion 150 -681 150 -681 0 feedthrough
rlabel pdiffusion 157 -681 157 -681 0 cellNo=333
rlabel pdiffusion 164 -681 164 -681 0 feedthrough
rlabel pdiffusion 171 -681 171 -681 0 feedthrough
rlabel pdiffusion 178 -681 178 -681 0 feedthrough
rlabel pdiffusion 185 -681 185 -681 0 cellNo=42
rlabel pdiffusion 192 -681 192 -681 0 feedthrough
rlabel pdiffusion 199 -681 199 -681 0 cellNo=185
rlabel pdiffusion 206 -681 206 -681 0 feedthrough
rlabel pdiffusion 213 -681 213 -681 0 feedthrough
rlabel pdiffusion 220 -681 220 -681 0 cellNo=244
rlabel pdiffusion 227 -681 227 -681 0 feedthrough
rlabel pdiffusion 234 -681 234 -681 0 feedthrough
rlabel pdiffusion 241 -681 241 -681 0 feedthrough
rlabel pdiffusion 248 -681 248 -681 0 feedthrough
rlabel pdiffusion 255 -681 255 -681 0 feedthrough
rlabel pdiffusion 262 -681 262 -681 0 feedthrough
rlabel pdiffusion 269 -681 269 -681 0 feedthrough
rlabel pdiffusion 276 -681 276 -681 0 cellNo=77
rlabel pdiffusion 283 -681 283 -681 0 cellNo=312
rlabel pdiffusion 290 -681 290 -681 0 feedthrough
rlabel pdiffusion 297 -681 297 -681 0 feedthrough
rlabel pdiffusion 304 -681 304 -681 0 feedthrough
rlabel pdiffusion 311 -681 311 -681 0 feedthrough
rlabel pdiffusion 318 -681 318 -681 0 cellNo=754
rlabel pdiffusion 325 -681 325 -681 0 cellNo=413
rlabel pdiffusion 332 -681 332 -681 0 feedthrough
rlabel pdiffusion 339 -681 339 -681 0 feedthrough
rlabel pdiffusion 346 -681 346 -681 0 cellNo=356
rlabel pdiffusion 353 -681 353 -681 0 cellNo=159
rlabel pdiffusion 360 -681 360 -681 0 feedthrough
rlabel pdiffusion 367 -681 367 -681 0 feedthrough
rlabel pdiffusion 374 -681 374 -681 0 feedthrough
rlabel pdiffusion 381 -681 381 -681 0 feedthrough
rlabel pdiffusion 388 -681 388 -681 0 feedthrough
rlabel pdiffusion 395 -681 395 -681 0 cellNo=336
rlabel pdiffusion 402 -681 402 -681 0 cellNo=363
rlabel pdiffusion 409 -681 409 -681 0 feedthrough
rlabel pdiffusion 416 -681 416 -681 0 feedthrough
rlabel pdiffusion 423 -681 423 -681 0 cellNo=30
rlabel pdiffusion 430 -681 430 -681 0 feedthrough
rlabel pdiffusion 437 -681 437 -681 0 cellNo=462
rlabel pdiffusion 444 -681 444 -681 0 feedthrough
rlabel pdiffusion 451 -681 451 -681 0 cellNo=672
rlabel pdiffusion 458 -681 458 -681 0 cellNo=69
rlabel pdiffusion 465 -681 465 -681 0 cellNo=666
rlabel pdiffusion 479 -681 479 -681 0 cellNo=448
rlabel pdiffusion 486 -681 486 -681 0 feedthrough
rlabel pdiffusion 493 -681 493 -681 0 cellNo=352
rlabel pdiffusion 500 -681 500 -681 0 feedthrough
rlabel pdiffusion 507 -681 507 -681 0 cellNo=73
rlabel pdiffusion 514 -681 514 -681 0 feedthrough
rlabel pdiffusion 521 -681 521 -681 0 feedthrough
rlabel pdiffusion 528 -681 528 -681 0 feedthrough
rlabel pdiffusion 535 -681 535 -681 0 feedthrough
rlabel pdiffusion 542 -681 542 -681 0 feedthrough
rlabel pdiffusion 549 -681 549 -681 0 feedthrough
rlabel pdiffusion 556 -681 556 -681 0 feedthrough
rlabel pdiffusion 563 -681 563 -681 0 feedthrough
rlabel pdiffusion 570 -681 570 -681 0 feedthrough
rlabel pdiffusion 577 -681 577 -681 0 feedthrough
rlabel pdiffusion 584 -681 584 -681 0 cellNo=983
rlabel pdiffusion 591 -681 591 -681 0 feedthrough
rlabel pdiffusion 598 -681 598 -681 0 feedthrough
rlabel pdiffusion 605 -681 605 -681 0 feedthrough
rlabel pdiffusion 612 -681 612 -681 0 feedthrough
rlabel pdiffusion 619 -681 619 -681 0 feedthrough
rlabel pdiffusion 626 -681 626 -681 0 feedthrough
rlabel pdiffusion 633 -681 633 -681 0 feedthrough
rlabel pdiffusion 640 -681 640 -681 0 feedthrough
rlabel pdiffusion 647 -681 647 -681 0 feedthrough
rlabel pdiffusion 654 -681 654 -681 0 feedthrough
rlabel pdiffusion 661 -681 661 -681 0 feedthrough
rlabel pdiffusion 668 -681 668 -681 0 feedthrough
rlabel pdiffusion 675 -681 675 -681 0 feedthrough
rlabel pdiffusion 682 -681 682 -681 0 feedthrough
rlabel pdiffusion 689 -681 689 -681 0 feedthrough
rlabel pdiffusion 696 -681 696 -681 0 feedthrough
rlabel pdiffusion 703 -681 703 -681 0 feedthrough
rlabel pdiffusion 710 -681 710 -681 0 feedthrough
rlabel pdiffusion 717 -681 717 -681 0 feedthrough
rlabel pdiffusion 724 -681 724 -681 0 feedthrough
rlabel pdiffusion 731 -681 731 -681 0 feedthrough
rlabel pdiffusion 738 -681 738 -681 0 feedthrough
rlabel pdiffusion 745 -681 745 -681 0 feedthrough
rlabel pdiffusion 752 -681 752 -681 0 feedthrough
rlabel pdiffusion 759 -681 759 -681 0 feedthrough
rlabel pdiffusion 766 -681 766 -681 0 feedthrough
rlabel pdiffusion 773 -681 773 -681 0 feedthrough
rlabel pdiffusion 3 -766 3 -766 0 cellNo=704
rlabel pdiffusion 17 -766 17 -766 0 cellNo=398
rlabel pdiffusion 24 -766 24 -766 0 cellNo=577
rlabel pdiffusion 31 -766 31 -766 0 cellNo=48
rlabel pdiffusion 38 -766 38 -766 0 feedthrough
rlabel pdiffusion 45 -766 45 -766 0 feedthrough
rlabel pdiffusion 52 -766 52 -766 0 cellNo=289
rlabel pdiffusion 59 -766 59 -766 0 feedthrough
rlabel pdiffusion 66 -766 66 -766 0 feedthrough
rlabel pdiffusion 73 -766 73 -766 0 feedthrough
rlabel pdiffusion 80 -766 80 -766 0 cellNo=263
rlabel pdiffusion 87 -766 87 -766 0 cellNo=405
rlabel pdiffusion 94 -766 94 -766 0 cellNo=532
rlabel pdiffusion 101 -766 101 -766 0 feedthrough
rlabel pdiffusion 108 -766 108 -766 0 feedthrough
rlabel pdiffusion 115 -766 115 -766 0 cellNo=224
rlabel pdiffusion 122 -766 122 -766 0 cellNo=673
rlabel pdiffusion 129 -766 129 -766 0 cellNo=271
rlabel pdiffusion 136 -766 136 -766 0 feedthrough
rlabel pdiffusion 143 -766 143 -766 0 feedthrough
rlabel pdiffusion 150 -766 150 -766 0 cellNo=911
rlabel pdiffusion 157 -766 157 -766 0 feedthrough
rlabel pdiffusion 164 -766 164 -766 0 feedthrough
rlabel pdiffusion 171 -766 171 -766 0 feedthrough
rlabel pdiffusion 178 -766 178 -766 0 feedthrough
rlabel pdiffusion 185 -766 185 -766 0 feedthrough
rlabel pdiffusion 192 -766 192 -766 0 feedthrough
rlabel pdiffusion 199 -766 199 -766 0 cellNo=839
rlabel pdiffusion 206 -766 206 -766 0 feedthrough
rlabel pdiffusion 213 -766 213 -766 0 feedthrough
rlabel pdiffusion 220 -766 220 -766 0 cellNo=908
rlabel pdiffusion 227 -766 227 -766 0 feedthrough
rlabel pdiffusion 234 -766 234 -766 0 feedthrough
rlabel pdiffusion 241 -766 241 -766 0 feedthrough
rlabel pdiffusion 248 -766 248 -766 0 feedthrough
rlabel pdiffusion 255 -766 255 -766 0 feedthrough
rlabel pdiffusion 262 -766 262 -766 0 feedthrough
rlabel pdiffusion 269 -766 269 -766 0 feedthrough
rlabel pdiffusion 276 -766 276 -766 0 feedthrough
rlabel pdiffusion 283 -766 283 -766 0 cellNo=277
rlabel pdiffusion 290 -766 290 -766 0 cellNo=205
rlabel pdiffusion 297 -766 297 -766 0 feedthrough
rlabel pdiffusion 304 -766 304 -766 0 cellNo=401
rlabel pdiffusion 311 -766 311 -766 0 cellNo=848
rlabel pdiffusion 318 -766 318 -766 0 cellNo=887
rlabel pdiffusion 325 -766 325 -766 0 feedthrough
rlabel pdiffusion 332 -766 332 -766 0 feedthrough
rlabel pdiffusion 339 -766 339 -766 0 feedthrough
rlabel pdiffusion 346 -766 346 -766 0 cellNo=828
rlabel pdiffusion 353 -766 353 -766 0 cellNo=307
rlabel pdiffusion 360 -766 360 -766 0 cellNo=565
rlabel pdiffusion 367 -766 367 -766 0 feedthrough
rlabel pdiffusion 374 -766 374 -766 0 feedthrough
rlabel pdiffusion 381 -766 381 -766 0 cellNo=249
rlabel pdiffusion 388 -766 388 -766 0 feedthrough
rlabel pdiffusion 395 -766 395 -766 0 cellNo=45
rlabel pdiffusion 402 -766 402 -766 0 feedthrough
rlabel pdiffusion 409 -766 409 -766 0 feedthrough
rlabel pdiffusion 416 -766 416 -766 0 feedthrough
rlabel pdiffusion 423 -766 423 -766 0 feedthrough
rlabel pdiffusion 430 -766 430 -766 0 cellNo=206
rlabel pdiffusion 437 -766 437 -766 0 cellNo=756
rlabel pdiffusion 444 -766 444 -766 0 cellNo=512
rlabel pdiffusion 451 -766 451 -766 0 feedthrough
rlabel pdiffusion 458 -766 458 -766 0 feedthrough
rlabel pdiffusion 465 -766 465 -766 0 feedthrough
rlabel pdiffusion 472 -766 472 -766 0 feedthrough
rlabel pdiffusion 479 -766 479 -766 0 cellNo=397
rlabel pdiffusion 486 -766 486 -766 0 cellNo=81
rlabel pdiffusion 493 -766 493 -766 0 feedthrough
rlabel pdiffusion 500 -766 500 -766 0 feedthrough
rlabel pdiffusion 507 -766 507 -766 0 feedthrough
rlabel pdiffusion 514 -766 514 -766 0 feedthrough
rlabel pdiffusion 521 -766 521 -766 0 feedthrough
rlabel pdiffusion 528 -766 528 -766 0 feedthrough
rlabel pdiffusion 535 -766 535 -766 0 cellNo=553
rlabel pdiffusion 542 -766 542 -766 0 feedthrough
rlabel pdiffusion 549 -766 549 -766 0 feedthrough
rlabel pdiffusion 556 -766 556 -766 0 feedthrough
rlabel pdiffusion 563 -766 563 -766 0 feedthrough
rlabel pdiffusion 570 -766 570 -766 0 feedthrough
rlabel pdiffusion 577 -766 577 -766 0 feedthrough
rlabel pdiffusion 584 -766 584 -766 0 feedthrough
rlabel pdiffusion 591 -766 591 -766 0 feedthrough
rlabel pdiffusion 598 -766 598 -766 0 feedthrough
rlabel pdiffusion 605 -766 605 -766 0 feedthrough
rlabel pdiffusion 612 -766 612 -766 0 feedthrough
rlabel pdiffusion 619 -766 619 -766 0 cellNo=203
rlabel pdiffusion 626 -766 626 -766 0 feedthrough
rlabel pdiffusion 633 -766 633 -766 0 feedthrough
rlabel pdiffusion 640 -766 640 -766 0 feedthrough
rlabel pdiffusion 647 -766 647 -766 0 feedthrough
rlabel pdiffusion 654 -766 654 -766 0 feedthrough
rlabel pdiffusion 661 -766 661 -766 0 feedthrough
rlabel pdiffusion 668 -766 668 -766 0 feedthrough
rlabel pdiffusion 675 -766 675 -766 0 feedthrough
rlabel pdiffusion 682 -766 682 -766 0 feedthrough
rlabel pdiffusion 689 -766 689 -766 0 feedthrough
rlabel pdiffusion 696 -766 696 -766 0 feedthrough
rlabel pdiffusion 703 -766 703 -766 0 feedthrough
rlabel pdiffusion 710 -766 710 -766 0 feedthrough
rlabel pdiffusion 717 -766 717 -766 0 feedthrough
rlabel pdiffusion 724 -766 724 -766 0 feedthrough
rlabel pdiffusion 731 -766 731 -766 0 cellNo=843
rlabel pdiffusion 738 -766 738 -766 0 feedthrough
rlabel pdiffusion 745 -766 745 -766 0 feedthrough
rlabel pdiffusion 752 -766 752 -766 0 feedthrough
rlabel pdiffusion 759 -766 759 -766 0 feedthrough
rlabel pdiffusion 766 -766 766 -766 0 feedthrough
rlabel pdiffusion 773 -766 773 -766 0 feedthrough
rlabel pdiffusion 780 -766 780 -766 0 feedthrough
rlabel pdiffusion 787 -766 787 -766 0 feedthrough
rlabel pdiffusion 794 -766 794 -766 0 feedthrough
rlabel pdiffusion 850 -766 850 -766 0 feedthrough
rlabel pdiffusion 3 -855 3 -855 0 cellNo=697
rlabel pdiffusion 10 -855 10 -855 0 cellNo=758
rlabel pdiffusion 17 -855 17 -855 0 cellNo=287
rlabel pdiffusion 24 -855 24 -855 0 feedthrough
rlabel pdiffusion 31 -855 31 -855 0 feedthrough
rlabel pdiffusion 38 -855 38 -855 0 cellNo=520
rlabel pdiffusion 45 -855 45 -855 0 feedthrough
rlabel pdiffusion 52 -855 52 -855 0 cellNo=649
rlabel pdiffusion 59 -855 59 -855 0 feedthrough
rlabel pdiffusion 66 -855 66 -855 0 feedthrough
rlabel pdiffusion 73 -855 73 -855 0 cellNo=782
rlabel pdiffusion 80 -855 80 -855 0 feedthrough
rlabel pdiffusion 87 -855 87 -855 0 cellNo=914
rlabel pdiffusion 94 -855 94 -855 0 feedthrough
rlabel pdiffusion 101 -855 101 -855 0 cellNo=255
rlabel pdiffusion 108 -855 108 -855 0 feedthrough
rlabel pdiffusion 115 -855 115 -855 0 feedthrough
rlabel pdiffusion 122 -855 122 -855 0 feedthrough
rlabel pdiffusion 129 -855 129 -855 0 feedthrough
rlabel pdiffusion 136 -855 136 -855 0 feedthrough
rlabel pdiffusion 143 -855 143 -855 0 cellNo=863
rlabel pdiffusion 150 -855 150 -855 0 cellNo=503
rlabel pdiffusion 157 -855 157 -855 0 cellNo=801
rlabel pdiffusion 164 -855 164 -855 0 cellNo=501
rlabel pdiffusion 171 -855 171 -855 0 feedthrough
rlabel pdiffusion 178 -855 178 -855 0 feedthrough
rlabel pdiffusion 185 -855 185 -855 0 feedthrough
rlabel pdiffusion 192 -855 192 -855 0 feedthrough
rlabel pdiffusion 199 -855 199 -855 0 feedthrough
rlabel pdiffusion 206 -855 206 -855 0 feedthrough
rlabel pdiffusion 213 -855 213 -855 0 feedthrough
rlabel pdiffusion 220 -855 220 -855 0 feedthrough
rlabel pdiffusion 227 -855 227 -855 0 feedthrough
rlabel pdiffusion 234 -855 234 -855 0 feedthrough
rlabel pdiffusion 241 -855 241 -855 0 feedthrough
rlabel pdiffusion 248 -855 248 -855 0 cellNo=997
rlabel pdiffusion 255 -855 255 -855 0 feedthrough
rlabel pdiffusion 262 -855 262 -855 0 cellNo=816
rlabel pdiffusion 269 -855 269 -855 0 feedthrough
rlabel pdiffusion 276 -855 276 -855 0 feedthrough
rlabel pdiffusion 283 -855 283 -855 0 feedthrough
rlabel pdiffusion 290 -855 290 -855 0 feedthrough
rlabel pdiffusion 297 -855 297 -855 0 cellNo=525
rlabel pdiffusion 304 -855 304 -855 0 cellNo=196
rlabel pdiffusion 311 -855 311 -855 0 feedthrough
rlabel pdiffusion 318 -855 318 -855 0 feedthrough
rlabel pdiffusion 325 -855 325 -855 0 cellNo=474
rlabel pdiffusion 332 -855 332 -855 0 cellNo=588
rlabel pdiffusion 339 -855 339 -855 0 cellNo=241
rlabel pdiffusion 346 -855 346 -855 0 feedthrough
rlabel pdiffusion 353 -855 353 -855 0 feedthrough
rlabel pdiffusion 360 -855 360 -855 0 cellNo=975
rlabel pdiffusion 367 -855 367 -855 0 feedthrough
rlabel pdiffusion 374 -855 374 -855 0 feedthrough
rlabel pdiffusion 381 -855 381 -855 0 cellNo=637
rlabel pdiffusion 388 -855 388 -855 0 feedthrough
rlabel pdiffusion 395 -855 395 -855 0 cellNo=291
rlabel pdiffusion 402 -855 402 -855 0 feedthrough
rlabel pdiffusion 409 -855 409 -855 0 cellNo=28
rlabel pdiffusion 416 -855 416 -855 0 feedthrough
rlabel pdiffusion 423 -855 423 -855 0 feedthrough
rlabel pdiffusion 430 -855 430 -855 0 cellNo=681
rlabel pdiffusion 437 -855 437 -855 0 cellNo=149
rlabel pdiffusion 444 -855 444 -855 0 cellNo=912
rlabel pdiffusion 451 -855 451 -855 0 cellNo=880
rlabel pdiffusion 458 -855 458 -855 0 cellNo=773
rlabel pdiffusion 465 -855 465 -855 0 cellNo=33
rlabel pdiffusion 472 -855 472 -855 0 feedthrough
rlabel pdiffusion 479 -855 479 -855 0 feedthrough
rlabel pdiffusion 486 -855 486 -855 0 feedthrough
rlabel pdiffusion 493 -855 493 -855 0 feedthrough
rlabel pdiffusion 500 -855 500 -855 0 feedthrough
rlabel pdiffusion 507 -855 507 -855 0 cellNo=463
rlabel pdiffusion 514 -855 514 -855 0 cellNo=231
rlabel pdiffusion 521 -855 521 -855 0 feedthrough
rlabel pdiffusion 528 -855 528 -855 0 feedthrough
rlabel pdiffusion 535 -855 535 -855 0 feedthrough
rlabel pdiffusion 542 -855 542 -855 0 feedthrough
rlabel pdiffusion 549 -855 549 -855 0 feedthrough
rlabel pdiffusion 556 -855 556 -855 0 feedthrough
rlabel pdiffusion 563 -855 563 -855 0 feedthrough
rlabel pdiffusion 570 -855 570 -855 0 feedthrough
rlabel pdiffusion 577 -855 577 -855 0 feedthrough
rlabel pdiffusion 584 -855 584 -855 0 feedthrough
rlabel pdiffusion 591 -855 591 -855 0 feedthrough
rlabel pdiffusion 598 -855 598 -855 0 feedthrough
rlabel pdiffusion 605 -855 605 -855 0 feedthrough
rlabel pdiffusion 612 -855 612 -855 0 feedthrough
rlabel pdiffusion 619 -855 619 -855 0 feedthrough
rlabel pdiffusion 626 -855 626 -855 0 feedthrough
rlabel pdiffusion 633 -855 633 -855 0 feedthrough
rlabel pdiffusion 640 -855 640 -855 0 feedthrough
rlabel pdiffusion 647 -855 647 -855 0 feedthrough
rlabel pdiffusion 654 -855 654 -855 0 feedthrough
rlabel pdiffusion 661 -855 661 -855 0 feedthrough
rlabel pdiffusion 668 -855 668 -855 0 feedthrough
rlabel pdiffusion 675 -855 675 -855 0 cellNo=114
rlabel pdiffusion 682 -855 682 -855 0 feedthrough
rlabel pdiffusion 689 -855 689 -855 0 feedthrough
rlabel pdiffusion 696 -855 696 -855 0 feedthrough
rlabel pdiffusion 703 -855 703 -855 0 feedthrough
rlabel pdiffusion 710 -855 710 -855 0 feedthrough
rlabel pdiffusion 717 -855 717 -855 0 feedthrough
rlabel pdiffusion 724 -855 724 -855 0 feedthrough
rlabel pdiffusion 731 -855 731 -855 0 feedthrough
rlabel pdiffusion 738 -855 738 -855 0 feedthrough
rlabel pdiffusion 745 -855 745 -855 0 feedthrough
rlabel pdiffusion 752 -855 752 -855 0 feedthrough
rlabel pdiffusion 759 -855 759 -855 0 feedthrough
rlabel pdiffusion 766 -855 766 -855 0 feedthrough
rlabel pdiffusion 773 -855 773 -855 0 feedthrough
rlabel pdiffusion 780 -855 780 -855 0 feedthrough
rlabel pdiffusion 787 -855 787 -855 0 feedthrough
rlabel pdiffusion 801 -855 801 -855 0 feedthrough
rlabel pdiffusion 808 -855 808 -855 0 feedthrough
rlabel pdiffusion 815 -855 815 -855 0 feedthrough
rlabel pdiffusion 822 -855 822 -855 0 feedthrough
rlabel pdiffusion 829 -855 829 -855 0 feedthrough
rlabel pdiffusion 836 -855 836 -855 0 feedthrough
rlabel pdiffusion 843 -855 843 -855 0 feedthrough
rlabel pdiffusion 850 -855 850 -855 0 feedthrough
rlabel pdiffusion 857 -855 857 -855 0 feedthrough
rlabel pdiffusion 864 -855 864 -855 0 feedthrough
rlabel pdiffusion 871 -855 871 -855 0 feedthrough
rlabel pdiffusion 941 -855 941 -855 0 feedthrough
rlabel pdiffusion 3 -932 3 -932 0 cellNo=741
rlabel pdiffusion 10 -932 10 -932 0 feedthrough
rlabel pdiffusion 17 -932 17 -932 0 feedthrough
rlabel pdiffusion 24 -932 24 -932 0 feedthrough
rlabel pdiffusion 31 -932 31 -932 0 feedthrough
rlabel pdiffusion 38 -932 38 -932 0 cellNo=743
rlabel pdiffusion 45 -932 45 -932 0 feedthrough
rlabel pdiffusion 52 -932 52 -932 0 cellNo=478
rlabel pdiffusion 59 -932 59 -932 0 feedthrough
rlabel pdiffusion 66 -932 66 -932 0 cellNo=387
rlabel pdiffusion 73 -932 73 -932 0 feedthrough
rlabel pdiffusion 80 -932 80 -932 0 cellNo=169
rlabel pdiffusion 87 -932 87 -932 0 feedthrough
rlabel pdiffusion 94 -932 94 -932 0 feedthrough
rlabel pdiffusion 101 -932 101 -932 0 feedthrough
rlabel pdiffusion 108 -932 108 -932 0 feedthrough
rlabel pdiffusion 115 -932 115 -932 0 feedthrough
rlabel pdiffusion 122 -932 122 -932 0 cellNo=324
rlabel pdiffusion 129 -932 129 -932 0 feedthrough
rlabel pdiffusion 136 -932 136 -932 0 feedthrough
rlabel pdiffusion 143 -932 143 -932 0 feedthrough
rlabel pdiffusion 150 -932 150 -932 0 cellNo=729
rlabel pdiffusion 157 -932 157 -932 0 feedthrough
rlabel pdiffusion 164 -932 164 -932 0 cellNo=342
rlabel pdiffusion 171 -932 171 -932 0 feedthrough
rlabel pdiffusion 178 -932 178 -932 0 feedthrough
rlabel pdiffusion 185 -932 185 -932 0 cellNo=360
rlabel pdiffusion 192 -932 192 -932 0 feedthrough
rlabel pdiffusion 199 -932 199 -932 0 cellNo=164
rlabel pdiffusion 206 -932 206 -932 0 cellNo=74
rlabel pdiffusion 213 -932 213 -932 0 cellNo=420
rlabel pdiffusion 220 -932 220 -932 0 cellNo=689
rlabel pdiffusion 227 -932 227 -932 0 feedthrough
rlabel pdiffusion 234 -932 234 -932 0 feedthrough
rlabel pdiffusion 241 -932 241 -932 0 feedthrough
rlabel pdiffusion 248 -932 248 -932 0 cellNo=920
rlabel pdiffusion 255 -932 255 -932 0 feedthrough
rlabel pdiffusion 262 -932 262 -932 0 feedthrough
rlabel pdiffusion 269 -932 269 -932 0 feedthrough
rlabel pdiffusion 276 -932 276 -932 0 cellNo=130
rlabel pdiffusion 283 -932 283 -932 0 cellNo=391
rlabel pdiffusion 290 -932 290 -932 0 feedthrough
rlabel pdiffusion 297 -932 297 -932 0 cellNo=509
rlabel pdiffusion 304 -932 304 -932 0 feedthrough
rlabel pdiffusion 311 -932 311 -932 0 feedthrough
rlabel pdiffusion 318 -932 318 -932 0 feedthrough
rlabel pdiffusion 325 -932 325 -932 0 feedthrough
rlabel pdiffusion 332 -932 332 -932 0 feedthrough
rlabel pdiffusion 339 -932 339 -932 0 cellNo=366
rlabel pdiffusion 346 -932 346 -932 0 cellNo=297
rlabel pdiffusion 353 -932 353 -932 0 cellNo=215
rlabel pdiffusion 360 -932 360 -932 0 feedthrough
rlabel pdiffusion 367 -932 367 -932 0 feedthrough
rlabel pdiffusion 374 -932 374 -932 0 feedthrough
rlabel pdiffusion 381 -932 381 -932 0 feedthrough
rlabel pdiffusion 388 -932 388 -932 0 feedthrough
rlabel pdiffusion 395 -932 395 -932 0 cellNo=759
rlabel pdiffusion 402 -932 402 -932 0 cellNo=51
rlabel pdiffusion 409 -932 409 -932 0 feedthrough
rlabel pdiffusion 416 -932 416 -932 0 feedthrough
rlabel pdiffusion 423 -932 423 -932 0 feedthrough
rlabel pdiffusion 430 -932 430 -932 0 feedthrough
rlabel pdiffusion 437 -932 437 -932 0 feedthrough
rlabel pdiffusion 444 -932 444 -932 0 cellNo=309
rlabel pdiffusion 451 -932 451 -932 0 cellNo=361
rlabel pdiffusion 458 -932 458 -932 0 feedthrough
rlabel pdiffusion 465 -932 465 -932 0 cellNo=97
rlabel pdiffusion 472 -932 472 -932 0 feedthrough
rlabel pdiffusion 479 -932 479 -932 0 feedthrough
rlabel pdiffusion 486 -932 486 -932 0 feedthrough
rlabel pdiffusion 493 -932 493 -932 0 feedthrough
rlabel pdiffusion 500 -932 500 -932 0 feedthrough
rlabel pdiffusion 507 -932 507 -932 0 cellNo=821
rlabel pdiffusion 514 -932 514 -932 0 cellNo=80
rlabel pdiffusion 521 -932 521 -932 0 feedthrough
rlabel pdiffusion 528 -932 528 -932 0 feedthrough
rlabel pdiffusion 535 -932 535 -932 0 feedthrough
rlabel pdiffusion 542 -932 542 -932 0 cellNo=524
rlabel pdiffusion 549 -932 549 -932 0 cellNo=218
rlabel pdiffusion 556 -932 556 -932 0 feedthrough
rlabel pdiffusion 563 -932 563 -932 0 feedthrough
rlabel pdiffusion 570 -932 570 -932 0 feedthrough
rlabel pdiffusion 577 -932 577 -932 0 feedthrough
rlabel pdiffusion 584 -932 584 -932 0 feedthrough
rlabel pdiffusion 591 -932 591 -932 0 cellNo=876
rlabel pdiffusion 598 -932 598 -932 0 feedthrough
rlabel pdiffusion 605 -932 605 -932 0 feedthrough
rlabel pdiffusion 612 -932 612 -932 0 feedthrough
rlabel pdiffusion 619 -932 619 -932 0 feedthrough
rlabel pdiffusion 626 -932 626 -932 0 feedthrough
rlabel pdiffusion 633 -932 633 -932 0 feedthrough
rlabel pdiffusion 640 -932 640 -932 0 feedthrough
rlabel pdiffusion 647 -932 647 -932 0 feedthrough
rlabel pdiffusion 654 -932 654 -932 0 feedthrough
rlabel pdiffusion 661 -932 661 -932 0 feedthrough
rlabel pdiffusion 668 -932 668 -932 0 feedthrough
rlabel pdiffusion 675 -932 675 -932 0 feedthrough
rlabel pdiffusion 682 -932 682 -932 0 feedthrough
rlabel pdiffusion 689 -932 689 -932 0 feedthrough
rlabel pdiffusion 696 -932 696 -932 0 feedthrough
rlabel pdiffusion 703 -932 703 -932 0 feedthrough
rlabel pdiffusion 710 -932 710 -932 0 feedthrough
rlabel pdiffusion 717 -932 717 -932 0 feedthrough
rlabel pdiffusion 724 -932 724 -932 0 feedthrough
rlabel pdiffusion 731 -932 731 -932 0 feedthrough
rlabel pdiffusion 738 -932 738 -932 0 feedthrough
rlabel pdiffusion 745 -932 745 -932 0 feedthrough
rlabel pdiffusion 752 -932 752 -932 0 feedthrough
rlabel pdiffusion 759 -932 759 -932 0 feedthrough
rlabel pdiffusion 766 -932 766 -932 0 feedthrough
rlabel pdiffusion 773 -932 773 -932 0 feedthrough
rlabel pdiffusion 780 -932 780 -932 0 feedthrough
rlabel pdiffusion 787 -932 787 -932 0 feedthrough
rlabel pdiffusion 794 -932 794 -932 0 feedthrough
rlabel pdiffusion 801 -932 801 -932 0 feedthrough
rlabel pdiffusion 808 -932 808 -932 0 feedthrough
rlabel pdiffusion 815 -932 815 -932 0 feedthrough
rlabel pdiffusion 822 -932 822 -932 0 feedthrough
rlabel pdiffusion 829 -932 829 -932 0 cellNo=655
rlabel pdiffusion 836 -932 836 -932 0 feedthrough
rlabel pdiffusion 843 -932 843 -932 0 feedthrough
rlabel pdiffusion 850 -932 850 -932 0 cellNo=303
rlabel pdiffusion 3 -1011 3 -1011 0 feedthrough
rlabel pdiffusion 10 -1011 10 -1011 0 feedthrough
rlabel pdiffusion 17 -1011 17 -1011 0 cellNo=658
rlabel pdiffusion 24 -1011 24 -1011 0 feedthrough
rlabel pdiffusion 31 -1011 31 -1011 0 cellNo=890
rlabel pdiffusion 38 -1011 38 -1011 0 feedthrough
rlabel pdiffusion 45 -1011 45 -1011 0 feedthrough
rlabel pdiffusion 52 -1011 52 -1011 0 feedthrough
rlabel pdiffusion 59 -1011 59 -1011 0 cellNo=217
rlabel pdiffusion 66 -1011 66 -1011 0 feedthrough
rlabel pdiffusion 73 -1011 73 -1011 0 feedthrough
rlabel pdiffusion 80 -1011 80 -1011 0 feedthrough
rlabel pdiffusion 87 -1011 87 -1011 0 feedthrough
rlabel pdiffusion 94 -1011 94 -1011 0 feedthrough
rlabel pdiffusion 101 -1011 101 -1011 0 cellNo=385
rlabel pdiffusion 108 -1011 108 -1011 0 feedthrough
rlabel pdiffusion 115 -1011 115 -1011 0 cellNo=194
rlabel pdiffusion 122 -1011 122 -1011 0 cellNo=557
rlabel pdiffusion 129 -1011 129 -1011 0 cellNo=123
rlabel pdiffusion 136 -1011 136 -1011 0 feedthrough
rlabel pdiffusion 143 -1011 143 -1011 0 feedthrough
rlabel pdiffusion 150 -1011 150 -1011 0 feedthrough
rlabel pdiffusion 157 -1011 157 -1011 0 feedthrough
rlabel pdiffusion 164 -1011 164 -1011 0 feedthrough
rlabel pdiffusion 171 -1011 171 -1011 0 cellNo=209
rlabel pdiffusion 178 -1011 178 -1011 0 feedthrough
rlabel pdiffusion 185 -1011 185 -1011 0 feedthrough
rlabel pdiffusion 192 -1011 192 -1011 0 cellNo=436
rlabel pdiffusion 199 -1011 199 -1011 0 cellNo=881
rlabel pdiffusion 206 -1011 206 -1011 0 feedthrough
rlabel pdiffusion 213 -1011 213 -1011 0 feedthrough
rlabel pdiffusion 220 -1011 220 -1011 0 cellNo=527
rlabel pdiffusion 227 -1011 227 -1011 0 feedthrough
rlabel pdiffusion 234 -1011 234 -1011 0 feedthrough
rlabel pdiffusion 241 -1011 241 -1011 0 feedthrough
rlabel pdiffusion 248 -1011 248 -1011 0 feedthrough
rlabel pdiffusion 255 -1011 255 -1011 0 feedthrough
rlabel pdiffusion 262 -1011 262 -1011 0 feedthrough
rlabel pdiffusion 269 -1011 269 -1011 0 cellNo=476
rlabel pdiffusion 276 -1011 276 -1011 0 feedthrough
rlabel pdiffusion 283 -1011 283 -1011 0 feedthrough
rlabel pdiffusion 290 -1011 290 -1011 0 feedthrough
rlabel pdiffusion 297 -1011 297 -1011 0 feedthrough
rlabel pdiffusion 304 -1011 304 -1011 0 feedthrough
rlabel pdiffusion 311 -1011 311 -1011 0 cellNo=924
rlabel pdiffusion 318 -1011 318 -1011 0 feedthrough
rlabel pdiffusion 325 -1011 325 -1011 0 feedthrough
rlabel pdiffusion 332 -1011 332 -1011 0 cellNo=84
rlabel pdiffusion 339 -1011 339 -1011 0 cellNo=88
rlabel pdiffusion 346 -1011 346 -1011 0 feedthrough
rlabel pdiffusion 353 -1011 353 -1011 0 feedthrough
rlabel pdiffusion 360 -1011 360 -1011 0 feedthrough
rlabel pdiffusion 367 -1011 367 -1011 0 cellNo=49
rlabel pdiffusion 374 -1011 374 -1011 0 cellNo=960
rlabel pdiffusion 381 -1011 381 -1011 0 feedthrough
rlabel pdiffusion 388 -1011 388 -1011 0 cellNo=866
rlabel pdiffusion 395 -1011 395 -1011 0 cellNo=236
rlabel pdiffusion 402 -1011 402 -1011 0 cellNo=158
rlabel pdiffusion 409 -1011 409 -1011 0 cellNo=726
rlabel pdiffusion 416 -1011 416 -1011 0 feedthrough
rlabel pdiffusion 423 -1011 423 -1011 0 cellNo=455
rlabel pdiffusion 430 -1011 430 -1011 0 cellNo=475
rlabel pdiffusion 437 -1011 437 -1011 0 cellNo=85
rlabel pdiffusion 444 -1011 444 -1011 0 feedthrough
rlabel pdiffusion 451 -1011 451 -1011 0 feedthrough
rlabel pdiffusion 458 -1011 458 -1011 0 feedthrough
rlabel pdiffusion 465 -1011 465 -1011 0 feedthrough
rlabel pdiffusion 472 -1011 472 -1011 0 cellNo=991
rlabel pdiffusion 479 -1011 479 -1011 0 cellNo=732
rlabel pdiffusion 486 -1011 486 -1011 0 feedthrough
rlabel pdiffusion 493 -1011 493 -1011 0 feedthrough
rlabel pdiffusion 500 -1011 500 -1011 0 cellNo=253
rlabel pdiffusion 507 -1011 507 -1011 0 cellNo=92
rlabel pdiffusion 514 -1011 514 -1011 0 cellNo=636
rlabel pdiffusion 521 -1011 521 -1011 0 feedthrough
rlabel pdiffusion 528 -1011 528 -1011 0 feedthrough
rlabel pdiffusion 535 -1011 535 -1011 0 feedthrough
rlabel pdiffusion 542 -1011 542 -1011 0 feedthrough
rlabel pdiffusion 549 -1011 549 -1011 0 feedthrough
rlabel pdiffusion 556 -1011 556 -1011 0 cellNo=552
rlabel pdiffusion 563 -1011 563 -1011 0 feedthrough
rlabel pdiffusion 570 -1011 570 -1011 0 feedthrough
rlabel pdiffusion 577 -1011 577 -1011 0 feedthrough
rlabel pdiffusion 591 -1011 591 -1011 0 feedthrough
rlabel pdiffusion 598 -1011 598 -1011 0 feedthrough
rlabel pdiffusion 605 -1011 605 -1011 0 feedthrough
rlabel pdiffusion 612 -1011 612 -1011 0 feedthrough
rlabel pdiffusion 619 -1011 619 -1011 0 feedthrough
rlabel pdiffusion 626 -1011 626 -1011 0 feedthrough
rlabel pdiffusion 633 -1011 633 -1011 0 feedthrough
rlabel pdiffusion 640 -1011 640 -1011 0 feedthrough
rlabel pdiffusion 647 -1011 647 -1011 0 feedthrough
rlabel pdiffusion 654 -1011 654 -1011 0 feedthrough
rlabel pdiffusion 661 -1011 661 -1011 0 feedthrough
rlabel pdiffusion 668 -1011 668 -1011 0 feedthrough
rlabel pdiffusion 675 -1011 675 -1011 0 feedthrough
rlabel pdiffusion 682 -1011 682 -1011 0 feedthrough
rlabel pdiffusion 689 -1011 689 -1011 0 feedthrough
rlabel pdiffusion 696 -1011 696 -1011 0 feedthrough
rlabel pdiffusion 703 -1011 703 -1011 0 feedthrough
rlabel pdiffusion 710 -1011 710 -1011 0 feedthrough
rlabel pdiffusion 717 -1011 717 -1011 0 feedthrough
rlabel pdiffusion 724 -1011 724 -1011 0 feedthrough
rlabel pdiffusion 731 -1011 731 -1011 0 feedthrough
rlabel pdiffusion 738 -1011 738 -1011 0 feedthrough
rlabel pdiffusion 745 -1011 745 -1011 0 feedthrough
rlabel pdiffusion 752 -1011 752 -1011 0 feedthrough
rlabel pdiffusion 759 -1011 759 -1011 0 feedthrough
rlabel pdiffusion 766 -1011 766 -1011 0 feedthrough
rlabel pdiffusion 773 -1011 773 -1011 0 feedthrough
rlabel pdiffusion 780 -1011 780 -1011 0 feedthrough
rlabel pdiffusion 787 -1011 787 -1011 0 feedthrough
rlabel pdiffusion 794 -1011 794 -1011 0 feedthrough
rlabel pdiffusion 801 -1011 801 -1011 0 feedthrough
rlabel pdiffusion 808 -1011 808 -1011 0 feedthrough
rlabel pdiffusion 815 -1011 815 -1011 0 feedthrough
rlabel pdiffusion 822 -1011 822 -1011 0 feedthrough
rlabel pdiffusion 829 -1011 829 -1011 0 feedthrough
rlabel pdiffusion 836 -1011 836 -1011 0 feedthrough
rlabel pdiffusion 843 -1011 843 -1011 0 feedthrough
rlabel pdiffusion 850 -1011 850 -1011 0 feedthrough
rlabel pdiffusion 857 -1011 857 -1011 0 cellNo=833
rlabel pdiffusion 864 -1011 864 -1011 0 feedthrough
rlabel pdiffusion 871 -1011 871 -1011 0 cellNo=492
rlabel pdiffusion 899 -1011 899 -1011 0 feedthrough
rlabel pdiffusion 3 -1088 3 -1088 0 cellNo=897
rlabel pdiffusion 10 -1088 10 -1088 0 cellNo=487
rlabel pdiffusion 17 -1088 17 -1088 0 feedthrough
rlabel pdiffusion 24 -1088 24 -1088 0 feedthrough
rlabel pdiffusion 31 -1088 31 -1088 0 feedthrough
rlabel pdiffusion 38 -1088 38 -1088 0 feedthrough
rlabel pdiffusion 45 -1088 45 -1088 0 feedthrough
rlabel pdiffusion 52 -1088 52 -1088 0 cellNo=189
rlabel pdiffusion 59 -1088 59 -1088 0 feedthrough
rlabel pdiffusion 66 -1088 66 -1088 0 cellNo=918
rlabel pdiffusion 73 -1088 73 -1088 0 feedthrough
rlabel pdiffusion 80 -1088 80 -1088 0 cellNo=867
rlabel pdiffusion 87 -1088 87 -1088 0 feedthrough
rlabel pdiffusion 94 -1088 94 -1088 0 cellNo=461
rlabel pdiffusion 101 -1088 101 -1088 0 cellNo=826
rlabel pdiffusion 108 -1088 108 -1088 0 feedthrough
rlabel pdiffusion 115 -1088 115 -1088 0 feedthrough
rlabel pdiffusion 122 -1088 122 -1088 0 feedthrough
rlabel pdiffusion 129 -1088 129 -1088 0 feedthrough
rlabel pdiffusion 136 -1088 136 -1088 0 cellNo=87
rlabel pdiffusion 143 -1088 143 -1088 0 feedthrough
rlabel pdiffusion 150 -1088 150 -1088 0 cellNo=679
rlabel pdiffusion 157 -1088 157 -1088 0 cellNo=536
rlabel pdiffusion 164 -1088 164 -1088 0 cellNo=780
rlabel pdiffusion 171 -1088 171 -1088 0 feedthrough
rlabel pdiffusion 178 -1088 178 -1088 0 feedthrough
rlabel pdiffusion 185 -1088 185 -1088 0 feedthrough
rlabel pdiffusion 192 -1088 192 -1088 0 feedthrough
rlabel pdiffusion 199 -1088 199 -1088 0 cellNo=940
rlabel pdiffusion 206 -1088 206 -1088 0 feedthrough
rlabel pdiffusion 213 -1088 213 -1088 0 feedthrough
rlabel pdiffusion 220 -1088 220 -1088 0 cellNo=79
rlabel pdiffusion 227 -1088 227 -1088 0 feedthrough
rlabel pdiffusion 234 -1088 234 -1088 0 feedthrough
rlabel pdiffusion 241 -1088 241 -1088 0 cellNo=299
rlabel pdiffusion 248 -1088 248 -1088 0 cellNo=445
rlabel pdiffusion 255 -1088 255 -1088 0 feedthrough
rlabel pdiffusion 262 -1088 262 -1088 0 feedthrough
rlabel pdiffusion 269 -1088 269 -1088 0 feedthrough
rlabel pdiffusion 276 -1088 276 -1088 0 cellNo=558
rlabel pdiffusion 283 -1088 283 -1088 0 feedthrough
rlabel pdiffusion 290 -1088 290 -1088 0 feedthrough
rlabel pdiffusion 297 -1088 297 -1088 0 feedthrough
rlabel pdiffusion 304 -1088 304 -1088 0 feedthrough
rlabel pdiffusion 311 -1088 311 -1088 0 feedthrough
rlabel pdiffusion 318 -1088 318 -1088 0 feedthrough
rlabel pdiffusion 325 -1088 325 -1088 0 feedthrough
rlabel pdiffusion 332 -1088 332 -1088 0 feedthrough
rlabel pdiffusion 339 -1088 339 -1088 0 feedthrough
rlabel pdiffusion 346 -1088 346 -1088 0 cellNo=560
rlabel pdiffusion 353 -1088 353 -1088 0 cellNo=106
rlabel pdiffusion 360 -1088 360 -1088 0 feedthrough
rlabel pdiffusion 367 -1088 367 -1088 0 feedthrough
rlabel pdiffusion 374 -1088 374 -1088 0 feedthrough
rlabel pdiffusion 381 -1088 381 -1088 0 feedthrough
rlabel pdiffusion 388 -1088 388 -1088 0 cellNo=269
rlabel pdiffusion 395 -1088 395 -1088 0 feedthrough
rlabel pdiffusion 402 -1088 402 -1088 0 feedthrough
rlabel pdiffusion 409 -1088 409 -1088 0 feedthrough
rlabel pdiffusion 416 -1088 416 -1088 0 feedthrough
rlabel pdiffusion 423 -1088 423 -1088 0 feedthrough
rlabel pdiffusion 430 -1088 430 -1088 0 feedthrough
rlabel pdiffusion 437 -1088 437 -1088 0 feedthrough
rlabel pdiffusion 444 -1088 444 -1088 0 cellNo=163
rlabel pdiffusion 451 -1088 451 -1088 0 cellNo=21
rlabel pdiffusion 458 -1088 458 -1088 0 feedthrough
rlabel pdiffusion 465 -1088 465 -1088 0 cellNo=504
rlabel pdiffusion 472 -1088 472 -1088 0 feedthrough
rlabel pdiffusion 479 -1088 479 -1088 0 feedthrough
rlabel pdiffusion 486 -1088 486 -1088 0 feedthrough
rlabel pdiffusion 493 -1088 493 -1088 0 cellNo=278
rlabel pdiffusion 500 -1088 500 -1088 0 feedthrough
rlabel pdiffusion 507 -1088 507 -1088 0 feedthrough
rlabel pdiffusion 514 -1088 514 -1088 0 feedthrough
rlabel pdiffusion 521 -1088 521 -1088 0 feedthrough
rlabel pdiffusion 528 -1088 528 -1088 0 cellNo=332
rlabel pdiffusion 535 -1088 535 -1088 0 cellNo=178
rlabel pdiffusion 542 -1088 542 -1088 0 feedthrough
rlabel pdiffusion 549 -1088 549 -1088 0 cellNo=543
rlabel pdiffusion 556 -1088 556 -1088 0 cellNo=111
rlabel pdiffusion 563 -1088 563 -1088 0 cellNo=676
rlabel pdiffusion 570 -1088 570 -1088 0 cellNo=986
rlabel pdiffusion 577 -1088 577 -1088 0 feedthrough
rlabel pdiffusion 584 -1088 584 -1088 0 feedthrough
rlabel pdiffusion 591 -1088 591 -1088 0 feedthrough
rlabel pdiffusion 598 -1088 598 -1088 0 feedthrough
rlabel pdiffusion 605 -1088 605 -1088 0 cellNo=559
rlabel pdiffusion 612 -1088 612 -1088 0 feedthrough
rlabel pdiffusion 619 -1088 619 -1088 0 feedthrough
rlabel pdiffusion 626 -1088 626 -1088 0 feedthrough
rlabel pdiffusion 633 -1088 633 -1088 0 feedthrough
rlabel pdiffusion 640 -1088 640 -1088 0 cellNo=257
rlabel pdiffusion 647 -1088 647 -1088 0 feedthrough
rlabel pdiffusion 654 -1088 654 -1088 0 feedthrough
rlabel pdiffusion 661 -1088 661 -1088 0 feedthrough
rlabel pdiffusion 668 -1088 668 -1088 0 feedthrough
rlabel pdiffusion 675 -1088 675 -1088 0 feedthrough
rlabel pdiffusion 682 -1088 682 -1088 0 feedthrough
rlabel pdiffusion 689 -1088 689 -1088 0 feedthrough
rlabel pdiffusion 696 -1088 696 -1088 0 feedthrough
rlabel pdiffusion 703 -1088 703 -1088 0 feedthrough
rlabel pdiffusion 710 -1088 710 -1088 0 feedthrough
rlabel pdiffusion 717 -1088 717 -1088 0 feedthrough
rlabel pdiffusion 724 -1088 724 -1088 0 feedthrough
rlabel pdiffusion 731 -1088 731 -1088 0 feedthrough
rlabel pdiffusion 738 -1088 738 -1088 0 feedthrough
rlabel pdiffusion 745 -1088 745 -1088 0 feedthrough
rlabel pdiffusion 752 -1088 752 -1088 0 feedthrough
rlabel pdiffusion 759 -1088 759 -1088 0 feedthrough
rlabel pdiffusion 766 -1088 766 -1088 0 feedthrough
rlabel pdiffusion 773 -1088 773 -1088 0 feedthrough
rlabel pdiffusion 780 -1088 780 -1088 0 feedthrough
rlabel pdiffusion 787 -1088 787 -1088 0 feedthrough
rlabel pdiffusion 794 -1088 794 -1088 0 feedthrough
rlabel pdiffusion 801 -1088 801 -1088 0 feedthrough
rlabel pdiffusion 808 -1088 808 -1088 0 feedthrough
rlabel pdiffusion 815 -1088 815 -1088 0 feedthrough
rlabel pdiffusion 822 -1088 822 -1088 0 feedthrough
rlabel pdiffusion 829 -1088 829 -1088 0 feedthrough
rlabel pdiffusion 836 -1088 836 -1088 0 feedthrough
rlabel pdiffusion 843 -1088 843 -1088 0 feedthrough
rlabel pdiffusion 850 -1088 850 -1088 0 feedthrough
rlabel pdiffusion 857 -1088 857 -1088 0 feedthrough
rlabel pdiffusion 864 -1088 864 -1088 0 feedthrough
rlabel pdiffusion 871 -1088 871 -1088 0 feedthrough
rlabel pdiffusion 878 -1088 878 -1088 0 feedthrough
rlabel pdiffusion 885 -1088 885 -1088 0 feedthrough
rlabel pdiffusion 892 -1088 892 -1088 0 feedthrough
rlabel pdiffusion 899 -1088 899 -1088 0 feedthrough
rlabel pdiffusion 906 -1088 906 -1088 0 feedthrough
rlabel pdiffusion 913 -1088 913 -1088 0 feedthrough
rlabel pdiffusion 920 -1088 920 -1088 0 feedthrough
rlabel pdiffusion 927 -1088 927 -1088 0 cellNo=638
rlabel pdiffusion 941 -1088 941 -1088 0 feedthrough
rlabel pdiffusion 3 -1185 3 -1185 0 cellNo=145
rlabel pdiffusion 10 -1185 10 -1185 0 feedthrough
rlabel pdiffusion 17 -1185 17 -1185 0 feedthrough
rlabel pdiffusion 24 -1185 24 -1185 0 cellNo=247
rlabel pdiffusion 31 -1185 31 -1185 0 feedthrough
rlabel pdiffusion 38 -1185 38 -1185 0 feedthrough
rlabel pdiffusion 45 -1185 45 -1185 0 feedthrough
rlabel pdiffusion 52 -1185 52 -1185 0 feedthrough
rlabel pdiffusion 59 -1185 59 -1185 0 feedthrough
rlabel pdiffusion 66 -1185 66 -1185 0 feedthrough
rlabel pdiffusion 73 -1185 73 -1185 0 cellNo=469
rlabel pdiffusion 80 -1185 80 -1185 0 feedthrough
rlabel pdiffusion 87 -1185 87 -1185 0 feedthrough
rlabel pdiffusion 94 -1185 94 -1185 0 cellNo=905
rlabel pdiffusion 101 -1185 101 -1185 0 cellNo=412
rlabel pdiffusion 108 -1185 108 -1185 0 feedthrough
rlabel pdiffusion 115 -1185 115 -1185 0 feedthrough
rlabel pdiffusion 122 -1185 122 -1185 0 cellNo=38
rlabel pdiffusion 129 -1185 129 -1185 0 feedthrough
rlabel pdiffusion 136 -1185 136 -1185 0 cellNo=894
rlabel pdiffusion 143 -1185 143 -1185 0 feedthrough
rlabel pdiffusion 150 -1185 150 -1185 0 cellNo=481
rlabel pdiffusion 157 -1185 157 -1185 0 feedthrough
rlabel pdiffusion 164 -1185 164 -1185 0 feedthrough
rlabel pdiffusion 171 -1185 171 -1185 0 cellNo=54
rlabel pdiffusion 178 -1185 178 -1185 0 feedthrough
rlabel pdiffusion 185 -1185 185 -1185 0 feedthrough
rlabel pdiffusion 192 -1185 192 -1185 0 feedthrough
rlabel pdiffusion 199 -1185 199 -1185 0 cellNo=31
rlabel pdiffusion 206 -1185 206 -1185 0 feedthrough
rlabel pdiffusion 213 -1185 213 -1185 0 cellNo=35
rlabel pdiffusion 220 -1185 220 -1185 0 cellNo=900
rlabel pdiffusion 227 -1185 227 -1185 0 feedthrough
rlabel pdiffusion 234 -1185 234 -1185 0 feedthrough
rlabel pdiffusion 241 -1185 241 -1185 0 feedthrough
rlabel pdiffusion 248 -1185 248 -1185 0 feedthrough
rlabel pdiffusion 255 -1185 255 -1185 0 feedthrough
rlabel pdiffusion 262 -1185 262 -1185 0 feedthrough
rlabel pdiffusion 269 -1185 269 -1185 0 feedthrough
rlabel pdiffusion 276 -1185 276 -1185 0 feedthrough
rlabel pdiffusion 283 -1185 283 -1185 0 cellNo=113
rlabel pdiffusion 290 -1185 290 -1185 0 feedthrough
rlabel pdiffusion 297 -1185 297 -1185 0 feedthrough
rlabel pdiffusion 304 -1185 304 -1185 0 feedthrough
rlabel pdiffusion 311 -1185 311 -1185 0 feedthrough
rlabel pdiffusion 318 -1185 318 -1185 0 cellNo=579
rlabel pdiffusion 325 -1185 325 -1185 0 feedthrough
rlabel pdiffusion 332 -1185 332 -1185 0 feedthrough
rlabel pdiffusion 339 -1185 339 -1185 0 feedthrough
rlabel pdiffusion 346 -1185 346 -1185 0 feedthrough
rlabel pdiffusion 353 -1185 353 -1185 0 cellNo=984
rlabel pdiffusion 360 -1185 360 -1185 0 cellNo=808
rlabel pdiffusion 367 -1185 367 -1185 0 feedthrough
rlabel pdiffusion 374 -1185 374 -1185 0 feedthrough
rlabel pdiffusion 381 -1185 381 -1185 0 feedthrough
rlabel pdiffusion 388 -1185 388 -1185 0 feedthrough
rlabel pdiffusion 395 -1185 395 -1185 0 feedthrough
rlabel pdiffusion 402 -1185 402 -1185 0 feedthrough
rlabel pdiffusion 409 -1185 409 -1185 0 cellNo=483
rlabel pdiffusion 416 -1185 416 -1185 0 feedthrough
rlabel pdiffusion 423 -1185 423 -1185 0 cellNo=103
rlabel pdiffusion 430 -1185 430 -1185 0 feedthrough
rlabel pdiffusion 437 -1185 437 -1185 0 feedthrough
rlabel pdiffusion 444 -1185 444 -1185 0 feedthrough
rlabel pdiffusion 451 -1185 451 -1185 0 cellNo=742
rlabel pdiffusion 458 -1185 458 -1185 0 feedthrough
rlabel pdiffusion 465 -1185 465 -1185 0 cellNo=468
rlabel pdiffusion 472 -1185 472 -1185 0 feedthrough
rlabel pdiffusion 479 -1185 479 -1185 0 cellNo=878
rlabel pdiffusion 486 -1185 486 -1185 0 feedthrough
rlabel pdiffusion 493 -1185 493 -1185 0 feedthrough
rlabel pdiffusion 500 -1185 500 -1185 0 feedthrough
rlabel pdiffusion 507 -1185 507 -1185 0 cellNo=432
rlabel pdiffusion 514 -1185 514 -1185 0 feedthrough
rlabel pdiffusion 521 -1185 521 -1185 0 feedthrough
rlabel pdiffusion 528 -1185 528 -1185 0 feedthrough
rlabel pdiffusion 535 -1185 535 -1185 0 feedthrough
rlabel pdiffusion 542 -1185 542 -1185 0 cellNo=744
rlabel pdiffusion 549 -1185 549 -1185 0 feedthrough
rlabel pdiffusion 556 -1185 556 -1185 0 feedthrough
rlabel pdiffusion 563 -1185 563 -1185 0 feedthrough
rlabel pdiffusion 570 -1185 570 -1185 0 feedthrough
rlabel pdiffusion 577 -1185 577 -1185 0 cellNo=266
rlabel pdiffusion 584 -1185 584 -1185 0 feedthrough
rlabel pdiffusion 591 -1185 591 -1185 0 feedthrough
rlabel pdiffusion 598 -1185 598 -1185 0 feedthrough
rlabel pdiffusion 605 -1185 605 -1185 0 feedthrough
rlabel pdiffusion 612 -1185 612 -1185 0 feedthrough
rlabel pdiffusion 619 -1185 619 -1185 0 cellNo=953
rlabel pdiffusion 626 -1185 626 -1185 0 feedthrough
rlabel pdiffusion 633 -1185 633 -1185 0 feedthrough
rlabel pdiffusion 640 -1185 640 -1185 0 feedthrough
rlabel pdiffusion 647 -1185 647 -1185 0 feedthrough
rlabel pdiffusion 654 -1185 654 -1185 0 cellNo=859
rlabel pdiffusion 661 -1185 661 -1185 0 feedthrough
rlabel pdiffusion 668 -1185 668 -1185 0 feedthrough
rlabel pdiffusion 675 -1185 675 -1185 0 feedthrough
rlabel pdiffusion 682 -1185 682 -1185 0 cellNo=722
rlabel pdiffusion 689 -1185 689 -1185 0 feedthrough
rlabel pdiffusion 696 -1185 696 -1185 0 feedthrough
rlabel pdiffusion 703 -1185 703 -1185 0 feedthrough
rlabel pdiffusion 710 -1185 710 -1185 0 feedthrough
rlabel pdiffusion 717 -1185 717 -1185 0 cellNo=22
rlabel pdiffusion 724 -1185 724 -1185 0 feedthrough
rlabel pdiffusion 731 -1185 731 -1185 0 feedthrough
rlabel pdiffusion 738 -1185 738 -1185 0 feedthrough
rlabel pdiffusion 745 -1185 745 -1185 0 feedthrough
rlabel pdiffusion 752 -1185 752 -1185 0 feedthrough
rlabel pdiffusion 759 -1185 759 -1185 0 feedthrough
rlabel pdiffusion 766 -1185 766 -1185 0 feedthrough
rlabel pdiffusion 773 -1185 773 -1185 0 feedthrough
rlabel pdiffusion 780 -1185 780 -1185 0 feedthrough
rlabel pdiffusion 787 -1185 787 -1185 0 feedthrough
rlabel pdiffusion 794 -1185 794 -1185 0 feedthrough
rlabel pdiffusion 801 -1185 801 -1185 0 feedthrough
rlabel pdiffusion 808 -1185 808 -1185 0 feedthrough
rlabel pdiffusion 815 -1185 815 -1185 0 feedthrough
rlabel pdiffusion 822 -1185 822 -1185 0 feedthrough
rlabel pdiffusion 829 -1185 829 -1185 0 feedthrough
rlabel pdiffusion 836 -1185 836 -1185 0 feedthrough
rlabel pdiffusion 843 -1185 843 -1185 0 feedthrough
rlabel pdiffusion 850 -1185 850 -1185 0 feedthrough
rlabel pdiffusion 857 -1185 857 -1185 0 feedthrough
rlabel pdiffusion 864 -1185 864 -1185 0 feedthrough
rlabel pdiffusion 871 -1185 871 -1185 0 feedthrough
rlabel pdiffusion 878 -1185 878 -1185 0 feedthrough
rlabel pdiffusion 885 -1185 885 -1185 0 feedthrough
rlabel pdiffusion 892 -1185 892 -1185 0 feedthrough
rlabel pdiffusion 899 -1185 899 -1185 0 feedthrough
rlabel pdiffusion 906 -1185 906 -1185 0 feedthrough
rlabel pdiffusion 913 -1185 913 -1185 0 feedthrough
rlabel pdiffusion 920 -1185 920 -1185 0 feedthrough
rlabel pdiffusion 927 -1185 927 -1185 0 feedthrough
rlabel pdiffusion 934 -1185 934 -1185 0 feedthrough
rlabel pdiffusion 941 -1185 941 -1185 0 feedthrough
rlabel pdiffusion 948 -1185 948 -1185 0 feedthrough
rlabel pdiffusion 955 -1185 955 -1185 0 cellNo=451
rlabel pdiffusion 962 -1185 962 -1185 0 cellNo=611
rlabel pdiffusion 969 -1185 969 -1185 0 cellNo=36
rlabel pdiffusion 976 -1185 976 -1185 0 feedthrough
rlabel pdiffusion 983 -1185 983 -1185 0 cellNo=753
rlabel pdiffusion 990 -1185 990 -1185 0 feedthrough
rlabel pdiffusion 3 -1280 3 -1280 0 cellNo=943
rlabel pdiffusion 10 -1280 10 -1280 0 cellNo=737
rlabel pdiffusion 17 -1280 17 -1280 0 feedthrough
rlabel pdiffusion 24 -1280 24 -1280 0 cellNo=694
rlabel pdiffusion 31 -1280 31 -1280 0 feedthrough
rlabel pdiffusion 38 -1280 38 -1280 0 cellNo=869
rlabel pdiffusion 45 -1280 45 -1280 0 feedthrough
rlabel pdiffusion 52 -1280 52 -1280 0 feedthrough
rlabel pdiffusion 59 -1280 59 -1280 0 feedthrough
rlabel pdiffusion 66 -1280 66 -1280 0 feedthrough
rlabel pdiffusion 73 -1280 73 -1280 0 feedthrough
rlabel pdiffusion 80 -1280 80 -1280 0 feedthrough
rlabel pdiffusion 87 -1280 87 -1280 0 feedthrough
rlabel pdiffusion 94 -1280 94 -1280 0 cellNo=519
rlabel pdiffusion 101 -1280 101 -1280 0 feedthrough
rlabel pdiffusion 108 -1280 108 -1280 0 cellNo=286
rlabel pdiffusion 115 -1280 115 -1280 0 feedthrough
rlabel pdiffusion 122 -1280 122 -1280 0 feedthrough
rlabel pdiffusion 129 -1280 129 -1280 0 cellNo=369
rlabel pdiffusion 136 -1280 136 -1280 0 feedthrough
rlabel pdiffusion 143 -1280 143 -1280 0 feedthrough
rlabel pdiffusion 150 -1280 150 -1280 0 feedthrough
rlabel pdiffusion 157 -1280 157 -1280 0 feedthrough
rlabel pdiffusion 164 -1280 164 -1280 0 feedthrough
rlabel pdiffusion 171 -1280 171 -1280 0 cellNo=612
rlabel pdiffusion 178 -1280 178 -1280 0 feedthrough
rlabel pdiffusion 185 -1280 185 -1280 0 cellNo=349
rlabel pdiffusion 192 -1280 192 -1280 0 feedthrough
rlabel pdiffusion 199 -1280 199 -1280 0 feedthrough
rlabel pdiffusion 206 -1280 206 -1280 0 feedthrough
rlabel pdiffusion 213 -1280 213 -1280 0 cellNo=298
rlabel pdiffusion 220 -1280 220 -1280 0 cellNo=795
rlabel pdiffusion 227 -1280 227 -1280 0 feedthrough
rlabel pdiffusion 234 -1280 234 -1280 0 feedthrough
rlabel pdiffusion 241 -1280 241 -1280 0 feedthrough
rlabel pdiffusion 248 -1280 248 -1280 0 feedthrough
rlabel pdiffusion 255 -1280 255 -1280 0 feedthrough
rlabel pdiffusion 262 -1280 262 -1280 0 feedthrough
rlabel pdiffusion 269 -1280 269 -1280 0 feedthrough
rlabel pdiffusion 276 -1280 276 -1280 0 feedthrough
rlabel pdiffusion 283 -1280 283 -1280 0 feedthrough
rlabel pdiffusion 290 -1280 290 -1280 0 feedthrough
rlabel pdiffusion 297 -1280 297 -1280 0 feedthrough
rlabel pdiffusion 304 -1280 304 -1280 0 cellNo=335
rlabel pdiffusion 311 -1280 311 -1280 0 cellNo=246
rlabel pdiffusion 318 -1280 318 -1280 0 feedthrough
rlabel pdiffusion 325 -1280 325 -1280 0 feedthrough
rlabel pdiffusion 332 -1280 332 -1280 0 feedthrough
rlabel pdiffusion 339 -1280 339 -1280 0 cellNo=115
rlabel pdiffusion 346 -1280 346 -1280 0 feedthrough
rlabel pdiffusion 353 -1280 353 -1280 0 feedthrough
rlabel pdiffusion 360 -1280 360 -1280 0 cellNo=755
rlabel pdiffusion 367 -1280 367 -1280 0 feedthrough
rlabel pdiffusion 374 -1280 374 -1280 0 feedthrough
rlabel pdiffusion 381 -1280 381 -1280 0 cellNo=350
rlabel pdiffusion 388 -1280 388 -1280 0 feedthrough
rlabel pdiffusion 395 -1280 395 -1280 0 feedthrough
rlabel pdiffusion 402 -1280 402 -1280 0 feedthrough
rlabel pdiffusion 409 -1280 409 -1280 0 cellNo=822
rlabel pdiffusion 416 -1280 416 -1280 0 feedthrough
rlabel pdiffusion 423 -1280 423 -1280 0 feedthrough
rlabel pdiffusion 430 -1280 430 -1280 0 feedthrough
rlabel pdiffusion 437 -1280 437 -1280 0 feedthrough
rlabel pdiffusion 444 -1280 444 -1280 0 cellNo=494
rlabel pdiffusion 451 -1280 451 -1280 0 feedthrough
rlabel pdiffusion 458 -1280 458 -1280 0 cellNo=771
rlabel pdiffusion 465 -1280 465 -1280 0 cellNo=290
rlabel pdiffusion 472 -1280 472 -1280 0 cellNo=907
rlabel pdiffusion 479 -1280 479 -1280 0 feedthrough
rlabel pdiffusion 486 -1280 486 -1280 0 feedthrough
rlabel pdiffusion 493 -1280 493 -1280 0 cellNo=477
rlabel pdiffusion 500 -1280 500 -1280 0 cellNo=354
rlabel pdiffusion 507 -1280 507 -1280 0 cellNo=318
rlabel pdiffusion 514 -1280 514 -1280 0 feedthrough
rlabel pdiffusion 521 -1280 521 -1280 0 feedthrough
rlabel pdiffusion 528 -1280 528 -1280 0 feedthrough
rlabel pdiffusion 535 -1280 535 -1280 0 feedthrough
rlabel pdiffusion 542 -1280 542 -1280 0 feedthrough
rlabel pdiffusion 549 -1280 549 -1280 0 feedthrough
rlabel pdiffusion 556 -1280 556 -1280 0 feedthrough
rlabel pdiffusion 563 -1280 563 -1280 0 feedthrough
rlabel pdiffusion 570 -1280 570 -1280 0 cellNo=259
rlabel pdiffusion 577 -1280 577 -1280 0 feedthrough
rlabel pdiffusion 584 -1280 584 -1280 0 feedthrough
rlabel pdiffusion 591 -1280 591 -1280 0 feedthrough
rlabel pdiffusion 598 -1280 598 -1280 0 cellNo=776
rlabel pdiffusion 605 -1280 605 -1280 0 cellNo=32
rlabel pdiffusion 612 -1280 612 -1280 0 feedthrough
rlabel pdiffusion 619 -1280 619 -1280 0 cellNo=25
rlabel pdiffusion 626 -1280 626 -1280 0 feedthrough
rlabel pdiffusion 633 -1280 633 -1280 0 cellNo=846
rlabel pdiffusion 640 -1280 640 -1280 0 feedthrough
rlabel pdiffusion 647 -1280 647 -1280 0 feedthrough
rlabel pdiffusion 654 -1280 654 -1280 0 cellNo=989
rlabel pdiffusion 661 -1280 661 -1280 0 feedthrough
rlabel pdiffusion 668 -1280 668 -1280 0 cellNo=227
rlabel pdiffusion 675 -1280 675 -1280 0 feedthrough
rlabel pdiffusion 682 -1280 682 -1280 0 feedthrough
rlabel pdiffusion 689 -1280 689 -1280 0 feedthrough
rlabel pdiffusion 696 -1280 696 -1280 0 feedthrough
rlabel pdiffusion 703 -1280 703 -1280 0 feedthrough
rlabel pdiffusion 710 -1280 710 -1280 0 feedthrough
rlabel pdiffusion 717 -1280 717 -1280 0 feedthrough
rlabel pdiffusion 724 -1280 724 -1280 0 feedthrough
rlabel pdiffusion 731 -1280 731 -1280 0 feedthrough
rlabel pdiffusion 738 -1280 738 -1280 0 feedthrough
rlabel pdiffusion 745 -1280 745 -1280 0 feedthrough
rlabel pdiffusion 752 -1280 752 -1280 0 feedthrough
rlabel pdiffusion 759 -1280 759 -1280 0 feedthrough
rlabel pdiffusion 766 -1280 766 -1280 0 feedthrough
rlabel pdiffusion 773 -1280 773 -1280 0 feedthrough
rlabel pdiffusion 780 -1280 780 -1280 0 feedthrough
rlabel pdiffusion 787 -1280 787 -1280 0 feedthrough
rlabel pdiffusion 794 -1280 794 -1280 0 feedthrough
rlabel pdiffusion 801 -1280 801 -1280 0 feedthrough
rlabel pdiffusion 808 -1280 808 -1280 0 feedthrough
rlabel pdiffusion 815 -1280 815 -1280 0 feedthrough
rlabel pdiffusion 822 -1280 822 -1280 0 feedthrough
rlabel pdiffusion 829 -1280 829 -1280 0 feedthrough
rlabel pdiffusion 836 -1280 836 -1280 0 feedthrough
rlabel pdiffusion 843 -1280 843 -1280 0 feedthrough
rlabel pdiffusion 850 -1280 850 -1280 0 feedthrough
rlabel pdiffusion 857 -1280 857 -1280 0 feedthrough
rlabel pdiffusion 864 -1280 864 -1280 0 feedthrough
rlabel pdiffusion 871 -1280 871 -1280 0 feedthrough
rlabel pdiffusion 878 -1280 878 -1280 0 feedthrough
rlabel pdiffusion 885 -1280 885 -1280 0 feedthrough
rlabel pdiffusion 892 -1280 892 -1280 0 feedthrough
rlabel pdiffusion 899 -1280 899 -1280 0 feedthrough
rlabel pdiffusion 906 -1280 906 -1280 0 feedthrough
rlabel pdiffusion 913 -1280 913 -1280 0 feedthrough
rlabel pdiffusion 920 -1280 920 -1280 0 feedthrough
rlabel pdiffusion 927 -1280 927 -1280 0 feedthrough
rlabel pdiffusion 934 -1280 934 -1280 0 feedthrough
rlabel pdiffusion 941 -1280 941 -1280 0 cellNo=99
rlabel pdiffusion 948 -1280 948 -1280 0 feedthrough
rlabel pdiffusion 955 -1280 955 -1280 0 feedthrough
rlabel pdiffusion 962 -1280 962 -1280 0 feedthrough
rlabel pdiffusion 969 -1280 969 -1280 0 feedthrough
rlabel pdiffusion 976 -1280 976 -1280 0 feedthrough
rlabel pdiffusion 983 -1280 983 -1280 0 feedthrough
rlabel pdiffusion 990 -1280 990 -1280 0 feedthrough
rlabel pdiffusion 997 -1280 997 -1280 0 feedthrough
rlabel pdiffusion 1004 -1280 1004 -1280 0 feedthrough
rlabel pdiffusion 1011 -1280 1011 -1280 0 feedthrough
rlabel pdiffusion 10 -1365 10 -1365 0 cellNo=639
rlabel pdiffusion 17 -1365 17 -1365 0 feedthrough
rlabel pdiffusion 24 -1365 24 -1365 0 cellNo=972
rlabel pdiffusion 31 -1365 31 -1365 0 cellNo=667
rlabel pdiffusion 38 -1365 38 -1365 0 feedthrough
rlabel pdiffusion 45 -1365 45 -1365 0 feedthrough
rlabel pdiffusion 52 -1365 52 -1365 0 feedthrough
rlabel pdiffusion 59 -1365 59 -1365 0 cellNo=830
rlabel pdiffusion 66 -1365 66 -1365 0 cellNo=657
rlabel pdiffusion 73 -1365 73 -1365 0 cellNo=748
rlabel pdiffusion 80 -1365 80 -1365 0 feedthrough
rlabel pdiffusion 87 -1365 87 -1365 0 cellNo=618
rlabel pdiffusion 94 -1365 94 -1365 0 feedthrough
rlabel pdiffusion 101 -1365 101 -1365 0 feedthrough
rlabel pdiffusion 108 -1365 108 -1365 0 feedthrough
rlabel pdiffusion 115 -1365 115 -1365 0 feedthrough
rlabel pdiffusion 122 -1365 122 -1365 0 cellNo=783
rlabel pdiffusion 129 -1365 129 -1365 0 feedthrough
rlabel pdiffusion 136 -1365 136 -1365 0 feedthrough
rlabel pdiffusion 143 -1365 143 -1365 0 feedthrough
rlabel pdiffusion 150 -1365 150 -1365 0 feedthrough
rlabel pdiffusion 157 -1365 157 -1365 0 cellNo=840
rlabel pdiffusion 164 -1365 164 -1365 0 feedthrough
rlabel pdiffusion 171 -1365 171 -1365 0 feedthrough
rlabel pdiffusion 178 -1365 178 -1365 0 feedthrough
rlabel pdiffusion 185 -1365 185 -1365 0 feedthrough
rlabel pdiffusion 192 -1365 192 -1365 0 cellNo=546
rlabel pdiffusion 199 -1365 199 -1365 0 feedthrough
rlabel pdiffusion 206 -1365 206 -1365 0 cellNo=903
rlabel pdiffusion 213 -1365 213 -1365 0 cellNo=736
rlabel pdiffusion 220 -1365 220 -1365 0 cellNo=529
rlabel pdiffusion 227 -1365 227 -1365 0 cellNo=104
rlabel pdiffusion 234 -1365 234 -1365 0 feedthrough
rlabel pdiffusion 241 -1365 241 -1365 0 feedthrough
rlabel pdiffusion 248 -1365 248 -1365 0 feedthrough
rlabel pdiffusion 255 -1365 255 -1365 0 feedthrough
rlabel pdiffusion 262 -1365 262 -1365 0 feedthrough
rlabel pdiffusion 269 -1365 269 -1365 0 feedthrough
rlabel pdiffusion 276 -1365 276 -1365 0 feedthrough
rlabel pdiffusion 283 -1365 283 -1365 0 feedthrough
rlabel pdiffusion 290 -1365 290 -1365 0 feedthrough
rlabel pdiffusion 297 -1365 297 -1365 0 feedthrough
rlabel pdiffusion 304 -1365 304 -1365 0 feedthrough
rlabel pdiffusion 311 -1365 311 -1365 0 feedthrough
rlabel pdiffusion 318 -1365 318 -1365 0 feedthrough
rlabel pdiffusion 325 -1365 325 -1365 0 feedthrough
rlabel pdiffusion 332 -1365 332 -1365 0 cellNo=11
rlabel pdiffusion 339 -1365 339 -1365 0 feedthrough
rlabel pdiffusion 346 -1365 346 -1365 0 cellNo=344
rlabel pdiffusion 353 -1365 353 -1365 0 feedthrough
rlabel pdiffusion 360 -1365 360 -1365 0 feedthrough
rlabel pdiffusion 367 -1365 367 -1365 0 feedthrough
rlabel pdiffusion 374 -1365 374 -1365 0 cellNo=198
rlabel pdiffusion 381 -1365 381 -1365 0 cellNo=686
rlabel pdiffusion 388 -1365 388 -1365 0 feedthrough
rlabel pdiffusion 395 -1365 395 -1365 0 cellNo=98
rlabel pdiffusion 402 -1365 402 -1365 0 feedthrough
rlabel pdiffusion 409 -1365 409 -1365 0 feedthrough
rlabel pdiffusion 416 -1365 416 -1365 0 feedthrough
rlabel pdiffusion 423 -1365 423 -1365 0 feedthrough
rlabel pdiffusion 430 -1365 430 -1365 0 cellNo=327
rlabel pdiffusion 437 -1365 437 -1365 0 feedthrough
rlabel pdiffusion 444 -1365 444 -1365 0 feedthrough
rlabel pdiffusion 451 -1365 451 -1365 0 cellNo=225
rlabel pdiffusion 458 -1365 458 -1365 0 feedthrough
rlabel pdiffusion 465 -1365 465 -1365 0 cellNo=155
rlabel pdiffusion 472 -1365 472 -1365 0 feedthrough
rlabel pdiffusion 479 -1365 479 -1365 0 cellNo=428
rlabel pdiffusion 486 -1365 486 -1365 0 cellNo=606
rlabel pdiffusion 493 -1365 493 -1365 0 feedthrough
rlabel pdiffusion 500 -1365 500 -1365 0 feedthrough
rlabel pdiffusion 507 -1365 507 -1365 0 feedthrough
rlabel pdiffusion 514 -1365 514 -1365 0 cellNo=373
rlabel pdiffusion 521 -1365 521 -1365 0 feedthrough
rlabel pdiffusion 528 -1365 528 -1365 0 cellNo=192
rlabel pdiffusion 535 -1365 535 -1365 0 feedthrough
rlabel pdiffusion 542 -1365 542 -1365 0 feedthrough
rlabel pdiffusion 549 -1365 549 -1365 0 feedthrough
rlabel pdiffusion 556 -1365 556 -1365 0 feedthrough
rlabel pdiffusion 563 -1365 563 -1365 0 feedthrough
rlabel pdiffusion 570 -1365 570 -1365 0 feedthrough
rlabel pdiffusion 577 -1365 577 -1365 0 cellNo=589
rlabel pdiffusion 584 -1365 584 -1365 0 feedthrough
rlabel pdiffusion 591 -1365 591 -1365 0 feedthrough
rlabel pdiffusion 598 -1365 598 -1365 0 feedthrough
rlabel pdiffusion 605 -1365 605 -1365 0 cellNo=18
rlabel pdiffusion 612 -1365 612 -1365 0 feedthrough
rlabel pdiffusion 619 -1365 619 -1365 0 feedthrough
rlabel pdiffusion 626 -1365 626 -1365 0 feedthrough
rlabel pdiffusion 633 -1365 633 -1365 0 feedthrough
rlabel pdiffusion 640 -1365 640 -1365 0 feedthrough
rlabel pdiffusion 647 -1365 647 -1365 0 feedthrough
rlabel pdiffusion 654 -1365 654 -1365 0 feedthrough
rlabel pdiffusion 661 -1365 661 -1365 0 feedthrough
rlabel pdiffusion 668 -1365 668 -1365 0 feedthrough
rlabel pdiffusion 675 -1365 675 -1365 0 feedthrough
rlabel pdiffusion 682 -1365 682 -1365 0 feedthrough
rlabel pdiffusion 689 -1365 689 -1365 0 feedthrough
rlabel pdiffusion 696 -1365 696 -1365 0 feedthrough
rlabel pdiffusion 703 -1365 703 -1365 0 feedthrough
rlabel pdiffusion 710 -1365 710 -1365 0 feedthrough
rlabel pdiffusion 717 -1365 717 -1365 0 feedthrough
rlabel pdiffusion 724 -1365 724 -1365 0 feedthrough
rlabel pdiffusion 731 -1365 731 -1365 0 feedthrough
rlabel pdiffusion 738 -1365 738 -1365 0 feedthrough
rlabel pdiffusion 745 -1365 745 -1365 0 feedthrough
rlabel pdiffusion 752 -1365 752 -1365 0 feedthrough
rlabel pdiffusion 759 -1365 759 -1365 0 feedthrough
rlabel pdiffusion 766 -1365 766 -1365 0 feedthrough
rlabel pdiffusion 773 -1365 773 -1365 0 feedthrough
rlabel pdiffusion 780 -1365 780 -1365 0 feedthrough
rlabel pdiffusion 787 -1365 787 -1365 0 feedthrough
rlabel pdiffusion 794 -1365 794 -1365 0 feedthrough
rlabel pdiffusion 801 -1365 801 -1365 0 feedthrough
rlabel pdiffusion 808 -1365 808 -1365 0 feedthrough
rlabel pdiffusion 815 -1365 815 -1365 0 feedthrough
rlabel pdiffusion 822 -1365 822 -1365 0 feedthrough
rlabel pdiffusion 829 -1365 829 -1365 0 feedthrough
rlabel pdiffusion 836 -1365 836 -1365 0 feedthrough
rlabel pdiffusion 843 -1365 843 -1365 0 feedthrough
rlabel pdiffusion 850 -1365 850 -1365 0 feedthrough
rlabel pdiffusion 857 -1365 857 -1365 0 feedthrough
rlabel pdiffusion 864 -1365 864 -1365 0 feedthrough
rlabel pdiffusion 871 -1365 871 -1365 0 feedthrough
rlabel pdiffusion 878 -1365 878 -1365 0 feedthrough
rlabel pdiffusion 885 -1365 885 -1365 0 feedthrough
rlabel pdiffusion 892 -1365 892 -1365 0 feedthrough
rlabel pdiffusion 899 -1365 899 -1365 0 feedthrough
rlabel pdiffusion 906 -1365 906 -1365 0 cellNo=630
rlabel pdiffusion 913 -1365 913 -1365 0 feedthrough
rlabel pdiffusion 920 -1365 920 -1365 0 cellNo=256
rlabel pdiffusion 941 -1365 941 -1365 0 cellNo=622
rlabel pdiffusion 955 -1365 955 -1365 0 feedthrough
rlabel pdiffusion 969 -1365 969 -1365 0 cellNo=122
rlabel pdiffusion 990 -1365 990 -1365 0 feedthrough
rlabel pdiffusion 3 -1444 3 -1444 0 feedthrough
rlabel pdiffusion 10 -1444 10 -1444 0 cellNo=235
rlabel pdiffusion 17 -1444 17 -1444 0 feedthrough
rlabel pdiffusion 24 -1444 24 -1444 0 feedthrough
rlabel pdiffusion 31 -1444 31 -1444 0 feedthrough
rlabel pdiffusion 38 -1444 38 -1444 0 feedthrough
rlabel pdiffusion 52 -1444 52 -1444 0 feedthrough
rlabel pdiffusion 59 -1444 59 -1444 0 feedthrough
rlabel pdiffusion 66 -1444 66 -1444 0 feedthrough
rlabel pdiffusion 73 -1444 73 -1444 0 feedthrough
rlabel pdiffusion 80 -1444 80 -1444 0 feedthrough
rlabel pdiffusion 87 -1444 87 -1444 0 feedthrough
rlabel pdiffusion 94 -1444 94 -1444 0 feedthrough
rlabel pdiffusion 101 -1444 101 -1444 0 feedthrough
rlabel pdiffusion 108 -1444 108 -1444 0 feedthrough
rlabel pdiffusion 115 -1444 115 -1444 0 cellNo=50
rlabel pdiffusion 122 -1444 122 -1444 0 cellNo=962
rlabel pdiffusion 129 -1444 129 -1444 0 cellNo=567
rlabel pdiffusion 136 -1444 136 -1444 0 feedthrough
rlabel pdiffusion 143 -1444 143 -1444 0 cellNo=899
rlabel pdiffusion 150 -1444 150 -1444 0 feedthrough
rlabel pdiffusion 157 -1444 157 -1444 0 cellNo=674
rlabel pdiffusion 164 -1444 164 -1444 0 cellNo=124
rlabel pdiffusion 171 -1444 171 -1444 0 feedthrough
rlabel pdiffusion 178 -1444 178 -1444 0 feedthrough
rlabel pdiffusion 185 -1444 185 -1444 0 cellNo=829
rlabel pdiffusion 192 -1444 192 -1444 0 feedthrough
rlabel pdiffusion 199 -1444 199 -1444 0 feedthrough
rlabel pdiffusion 206 -1444 206 -1444 0 feedthrough
rlabel pdiffusion 213 -1444 213 -1444 0 cellNo=634
rlabel pdiffusion 220 -1444 220 -1444 0 feedthrough
rlabel pdiffusion 227 -1444 227 -1444 0 feedthrough
rlabel pdiffusion 234 -1444 234 -1444 0 feedthrough
rlabel pdiffusion 241 -1444 241 -1444 0 feedthrough
rlabel pdiffusion 248 -1444 248 -1444 0 feedthrough
rlabel pdiffusion 255 -1444 255 -1444 0 feedthrough
rlabel pdiffusion 262 -1444 262 -1444 0 feedthrough
rlabel pdiffusion 269 -1444 269 -1444 0 feedthrough
rlabel pdiffusion 276 -1444 276 -1444 0 feedthrough
rlabel pdiffusion 283 -1444 283 -1444 0 feedthrough
rlabel pdiffusion 290 -1444 290 -1444 0 feedthrough
rlabel pdiffusion 297 -1444 297 -1444 0 feedthrough
rlabel pdiffusion 304 -1444 304 -1444 0 feedthrough
rlabel pdiffusion 311 -1444 311 -1444 0 feedthrough
rlabel pdiffusion 318 -1444 318 -1444 0 feedthrough
rlabel pdiffusion 325 -1444 325 -1444 0 cellNo=283
rlabel pdiffusion 332 -1444 332 -1444 0 feedthrough
rlabel pdiffusion 339 -1444 339 -1444 0 cellNo=693
rlabel pdiffusion 346 -1444 346 -1444 0 feedthrough
rlabel pdiffusion 353 -1444 353 -1444 0 cellNo=835
rlabel pdiffusion 360 -1444 360 -1444 0 feedthrough
rlabel pdiffusion 367 -1444 367 -1444 0 feedthrough
rlabel pdiffusion 374 -1444 374 -1444 0 cellNo=197
rlabel pdiffusion 381 -1444 381 -1444 0 feedthrough
rlabel pdiffusion 388 -1444 388 -1444 0 cellNo=9
rlabel pdiffusion 395 -1444 395 -1444 0 cellNo=852
rlabel pdiffusion 402 -1444 402 -1444 0 feedthrough
rlabel pdiffusion 409 -1444 409 -1444 0 feedthrough
rlabel pdiffusion 416 -1444 416 -1444 0 feedthrough
rlabel pdiffusion 423 -1444 423 -1444 0 feedthrough
rlabel pdiffusion 430 -1444 430 -1444 0 cellNo=392
rlabel pdiffusion 437 -1444 437 -1444 0 feedthrough
rlabel pdiffusion 444 -1444 444 -1444 0 feedthrough
rlabel pdiffusion 451 -1444 451 -1444 0 cellNo=791
rlabel pdiffusion 458 -1444 458 -1444 0 cellNo=624
rlabel pdiffusion 465 -1444 465 -1444 0 cellNo=146
rlabel pdiffusion 472 -1444 472 -1444 0 feedthrough
rlabel pdiffusion 479 -1444 479 -1444 0 feedthrough
rlabel pdiffusion 486 -1444 486 -1444 0 cellNo=956
rlabel pdiffusion 493 -1444 493 -1444 0 feedthrough
rlabel pdiffusion 500 -1444 500 -1444 0 feedthrough
rlabel pdiffusion 507 -1444 507 -1444 0 cellNo=214
rlabel pdiffusion 514 -1444 514 -1444 0 feedthrough
rlabel pdiffusion 521 -1444 521 -1444 0 feedthrough
rlabel pdiffusion 528 -1444 528 -1444 0 feedthrough
rlabel pdiffusion 535 -1444 535 -1444 0 cellNo=749
rlabel pdiffusion 542 -1444 542 -1444 0 feedthrough
rlabel pdiffusion 549 -1444 549 -1444 0 cellNo=341
rlabel pdiffusion 556 -1444 556 -1444 0 cellNo=83
rlabel pdiffusion 563 -1444 563 -1444 0 feedthrough
rlabel pdiffusion 570 -1444 570 -1444 0 feedthrough
rlabel pdiffusion 577 -1444 577 -1444 0 cellNo=276
rlabel pdiffusion 584 -1444 584 -1444 0 feedthrough
rlabel pdiffusion 591 -1444 591 -1444 0 cellNo=480
rlabel pdiffusion 598 -1444 598 -1444 0 feedthrough
rlabel pdiffusion 605 -1444 605 -1444 0 cellNo=786
rlabel pdiffusion 612 -1444 612 -1444 0 feedthrough
rlabel pdiffusion 619 -1444 619 -1444 0 feedthrough
rlabel pdiffusion 626 -1444 626 -1444 0 feedthrough
rlabel pdiffusion 633 -1444 633 -1444 0 cellNo=945
rlabel pdiffusion 640 -1444 640 -1444 0 feedthrough
rlabel pdiffusion 647 -1444 647 -1444 0 feedthrough
rlabel pdiffusion 654 -1444 654 -1444 0 cellNo=614
rlabel pdiffusion 661 -1444 661 -1444 0 feedthrough
rlabel pdiffusion 668 -1444 668 -1444 0 feedthrough
rlabel pdiffusion 675 -1444 675 -1444 0 feedthrough
rlabel pdiffusion 682 -1444 682 -1444 0 feedthrough
rlabel pdiffusion 689 -1444 689 -1444 0 feedthrough
rlabel pdiffusion 696 -1444 696 -1444 0 feedthrough
rlabel pdiffusion 703 -1444 703 -1444 0 feedthrough
rlabel pdiffusion 710 -1444 710 -1444 0 cellNo=314
rlabel pdiffusion 717 -1444 717 -1444 0 feedthrough
rlabel pdiffusion 724 -1444 724 -1444 0 feedthrough
rlabel pdiffusion 731 -1444 731 -1444 0 feedthrough
rlabel pdiffusion 738 -1444 738 -1444 0 feedthrough
rlabel pdiffusion 745 -1444 745 -1444 0 feedthrough
rlabel pdiffusion 752 -1444 752 -1444 0 feedthrough
rlabel pdiffusion 759 -1444 759 -1444 0 feedthrough
rlabel pdiffusion 766 -1444 766 -1444 0 feedthrough
rlabel pdiffusion 773 -1444 773 -1444 0 feedthrough
rlabel pdiffusion 780 -1444 780 -1444 0 feedthrough
rlabel pdiffusion 787 -1444 787 -1444 0 feedthrough
rlabel pdiffusion 794 -1444 794 -1444 0 feedthrough
rlabel pdiffusion 801 -1444 801 -1444 0 feedthrough
rlabel pdiffusion 808 -1444 808 -1444 0 feedthrough
rlabel pdiffusion 815 -1444 815 -1444 0 feedthrough
rlabel pdiffusion 822 -1444 822 -1444 0 feedthrough
rlabel pdiffusion 836 -1444 836 -1444 0 feedthrough
rlabel pdiffusion 843 -1444 843 -1444 0 feedthrough
rlabel pdiffusion 850 -1444 850 -1444 0 feedthrough
rlabel pdiffusion 857 -1444 857 -1444 0 feedthrough
rlabel pdiffusion 864 -1444 864 -1444 0 feedthrough
rlabel pdiffusion 871 -1444 871 -1444 0 feedthrough
rlabel pdiffusion 878 -1444 878 -1444 0 feedthrough
rlabel pdiffusion 885 -1444 885 -1444 0 feedthrough
rlabel pdiffusion 892 -1444 892 -1444 0 feedthrough
rlabel pdiffusion 899 -1444 899 -1444 0 feedthrough
rlabel pdiffusion 906 -1444 906 -1444 0 feedthrough
rlabel pdiffusion 913 -1444 913 -1444 0 feedthrough
rlabel pdiffusion 920 -1444 920 -1444 0 feedthrough
rlabel pdiffusion 927 -1444 927 -1444 0 feedthrough
rlabel pdiffusion 934 -1444 934 -1444 0 feedthrough
rlabel pdiffusion 941 -1444 941 -1444 0 cellNo=175
rlabel pdiffusion 948 -1444 948 -1444 0 cellNo=885
rlabel pdiffusion 955 -1444 955 -1444 0 feedthrough
rlabel pdiffusion 969 -1444 969 -1444 0 feedthrough
rlabel pdiffusion 983 -1444 983 -1444 0 feedthrough
rlabel pdiffusion 10 -1533 10 -1533 0 feedthrough
rlabel pdiffusion 17 -1533 17 -1533 0 feedthrough
rlabel pdiffusion 24 -1533 24 -1533 0 cellNo=718
rlabel pdiffusion 31 -1533 31 -1533 0 feedthrough
rlabel pdiffusion 38 -1533 38 -1533 0 cellNo=711
rlabel pdiffusion 45 -1533 45 -1533 0 feedthrough
rlabel pdiffusion 52 -1533 52 -1533 0 feedthrough
rlabel pdiffusion 59 -1533 59 -1533 0 feedthrough
rlabel pdiffusion 66 -1533 66 -1533 0 feedthrough
rlabel pdiffusion 73 -1533 73 -1533 0 cellNo=970
rlabel pdiffusion 80 -1533 80 -1533 0 feedthrough
rlabel pdiffusion 87 -1533 87 -1533 0 feedthrough
rlabel pdiffusion 94 -1533 94 -1533 0 feedthrough
rlabel pdiffusion 101 -1533 101 -1533 0 feedthrough
rlabel pdiffusion 108 -1533 108 -1533 0 feedthrough
rlabel pdiffusion 115 -1533 115 -1533 0 feedthrough
rlabel pdiffusion 122 -1533 122 -1533 0 feedthrough
rlabel pdiffusion 129 -1533 129 -1533 0 feedthrough
rlabel pdiffusion 136 -1533 136 -1533 0 cellNo=133
rlabel pdiffusion 143 -1533 143 -1533 0 feedthrough
rlabel pdiffusion 150 -1533 150 -1533 0 cellNo=647
rlabel pdiffusion 157 -1533 157 -1533 0 cellNo=521
rlabel pdiffusion 164 -1533 164 -1533 0 cellNo=849
rlabel pdiffusion 171 -1533 171 -1533 0 cellNo=654
rlabel pdiffusion 178 -1533 178 -1533 0 cellNo=172
rlabel pdiffusion 185 -1533 185 -1533 0 cellNo=17
rlabel pdiffusion 192 -1533 192 -1533 0 cellNo=596
rlabel pdiffusion 199 -1533 199 -1533 0 cellNo=645
rlabel pdiffusion 206 -1533 206 -1533 0 feedthrough
rlabel pdiffusion 213 -1533 213 -1533 0 cellNo=281
rlabel pdiffusion 220 -1533 220 -1533 0 cellNo=187
rlabel pdiffusion 227 -1533 227 -1533 0 feedthrough
rlabel pdiffusion 234 -1533 234 -1533 0 feedthrough
rlabel pdiffusion 241 -1533 241 -1533 0 feedthrough
rlabel pdiffusion 248 -1533 248 -1533 0 feedthrough
rlabel pdiffusion 255 -1533 255 -1533 0 feedthrough
rlabel pdiffusion 262 -1533 262 -1533 0 feedthrough
rlabel pdiffusion 269 -1533 269 -1533 0 feedthrough
rlabel pdiffusion 276 -1533 276 -1533 0 feedthrough
rlabel pdiffusion 283 -1533 283 -1533 0 cellNo=948
rlabel pdiffusion 290 -1533 290 -1533 0 feedthrough
rlabel pdiffusion 297 -1533 297 -1533 0 feedthrough
rlabel pdiffusion 304 -1533 304 -1533 0 cellNo=403
rlabel pdiffusion 311 -1533 311 -1533 0 feedthrough
rlabel pdiffusion 318 -1533 318 -1533 0 feedthrough
rlabel pdiffusion 325 -1533 325 -1533 0 feedthrough
rlabel pdiffusion 332 -1533 332 -1533 0 feedthrough
rlabel pdiffusion 339 -1533 339 -1533 0 feedthrough
rlabel pdiffusion 346 -1533 346 -1533 0 feedthrough
rlabel pdiffusion 353 -1533 353 -1533 0 feedthrough
rlabel pdiffusion 360 -1533 360 -1533 0 cellNo=453
rlabel pdiffusion 367 -1533 367 -1533 0 cellNo=779
rlabel pdiffusion 374 -1533 374 -1533 0 feedthrough
rlabel pdiffusion 381 -1533 381 -1533 0 feedthrough
rlabel pdiffusion 388 -1533 388 -1533 0 feedthrough
rlabel pdiffusion 395 -1533 395 -1533 0 feedthrough
rlabel pdiffusion 402 -1533 402 -1533 0 feedthrough
rlabel pdiffusion 409 -1533 409 -1533 0 cellNo=913
rlabel pdiffusion 416 -1533 416 -1533 0 feedthrough
rlabel pdiffusion 423 -1533 423 -1533 0 feedthrough
rlabel pdiffusion 430 -1533 430 -1533 0 cellNo=680
rlabel pdiffusion 437 -1533 437 -1533 0 feedthrough
rlabel pdiffusion 444 -1533 444 -1533 0 cellNo=692
rlabel pdiffusion 451 -1533 451 -1533 0 cellNo=669
rlabel pdiffusion 458 -1533 458 -1533 0 feedthrough
rlabel pdiffusion 465 -1533 465 -1533 0 cellNo=958
rlabel pdiffusion 472 -1533 472 -1533 0 feedthrough
rlabel pdiffusion 479 -1533 479 -1533 0 cellNo=540
rlabel pdiffusion 486 -1533 486 -1533 0 feedthrough
rlabel pdiffusion 493 -1533 493 -1533 0 feedthrough
rlabel pdiffusion 500 -1533 500 -1533 0 cellNo=752
rlabel pdiffusion 507 -1533 507 -1533 0 cellNo=228
rlabel pdiffusion 514 -1533 514 -1533 0 feedthrough
rlabel pdiffusion 521 -1533 521 -1533 0 feedthrough
rlabel pdiffusion 528 -1533 528 -1533 0 feedthrough
rlabel pdiffusion 535 -1533 535 -1533 0 cellNo=616
rlabel pdiffusion 542 -1533 542 -1533 0 feedthrough
rlabel pdiffusion 549 -1533 549 -1533 0 feedthrough
rlabel pdiffusion 556 -1533 556 -1533 0 cellNo=847
rlabel pdiffusion 563 -1533 563 -1533 0 feedthrough
rlabel pdiffusion 570 -1533 570 -1533 0 feedthrough
rlabel pdiffusion 577 -1533 577 -1533 0 feedthrough
rlabel pdiffusion 584 -1533 584 -1533 0 feedthrough
rlabel pdiffusion 591 -1533 591 -1533 0 feedthrough
rlabel pdiffusion 598 -1533 598 -1533 0 feedthrough
rlabel pdiffusion 605 -1533 605 -1533 0 feedthrough
rlabel pdiffusion 612 -1533 612 -1533 0 feedthrough
rlabel pdiffusion 619 -1533 619 -1533 0 feedthrough
rlabel pdiffusion 626 -1533 626 -1533 0 feedthrough
rlabel pdiffusion 633 -1533 633 -1533 0 feedthrough
rlabel pdiffusion 640 -1533 640 -1533 0 feedthrough
rlabel pdiffusion 647 -1533 647 -1533 0 feedthrough
rlabel pdiffusion 654 -1533 654 -1533 0 feedthrough
rlabel pdiffusion 661 -1533 661 -1533 0 feedthrough
rlabel pdiffusion 668 -1533 668 -1533 0 feedthrough
rlabel pdiffusion 675 -1533 675 -1533 0 feedthrough
rlabel pdiffusion 682 -1533 682 -1533 0 feedthrough
rlabel pdiffusion 689 -1533 689 -1533 0 feedthrough
rlabel pdiffusion 696 -1533 696 -1533 0 feedthrough
rlabel pdiffusion 703 -1533 703 -1533 0 feedthrough
rlabel pdiffusion 710 -1533 710 -1533 0 feedthrough
rlabel pdiffusion 717 -1533 717 -1533 0 feedthrough
rlabel pdiffusion 724 -1533 724 -1533 0 feedthrough
rlabel pdiffusion 731 -1533 731 -1533 0 feedthrough
rlabel pdiffusion 738 -1533 738 -1533 0 feedthrough
rlabel pdiffusion 745 -1533 745 -1533 0 feedthrough
rlabel pdiffusion 752 -1533 752 -1533 0 feedthrough
rlabel pdiffusion 766 -1533 766 -1533 0 feedthrough
rlabel pdiffusion 773 -1533 773 -1533 0 feedthrough
rlabel pdiffusion 780 -1533 780 -1533 0 feedthrough
rlabel pdiffusion 787 -1533 787 -1533 0 feedthrough
rlabel pdiffusion 794 -1533 794 -1533 0 feedthrough
rlabel pdiffusion 801 -1533 801 -1533 0 feedthrough
rlabel pdiffusion 808 -1533 808 -1533 0 feedthrough
rlabel pdiffusion 815 -1533 815 -1533 0 feedthrough
rlabel pdiffusion 822 -1533 822 -1533 0 feedthrough
rlabel pdiffusion 829 -1533 829 -1533 0 feedthrough
rlabel pdiffusion 836 -1533 836 -1533 0 feedthrough
rlabel pdiffusion 843 -1533 843 -1533 0 feedthrough
rlabel pdiffusion 850 -1533 850 -1533 0 feedthrough
rlabel pdiffusion 857 -1533 857 -1533 0 feedthrough
rlabel pdiffusion 885 -1533 885 -1533 0 cellNo=334
rlabel pdiffusion 892 -1533 892 -1533 0 feedthrough
rlabel pdiffusion 899 -1533 899 -1533 0 feedthrough
rlabel pdiffusion 906 -1533 906 -1533 0 feedthrough
rlabel pdiffusion 913 -1533 913 -1533 0 feedthrough
rlabel pdiffusion 920 -1533 920 -1533 0 feedthrough
rlabel pdiffusion 934 -1533 934 -1533 0 cellNo=295
rlabel pdiffusion 941 -1533 941 -1533 0 feedthrough
rlabel pdiffusion 955 -1533 955 -1533 0 feedthrough
rlabel pdiffusion 962 -1533 962 -1533 0 cellNo=957
rlabel pdiffusion 983 -1533 983 -1533 0 cellNo=340
rlabel pdiffusion 990 -1533 990 -1533 0 feedthrough
rlabel pdiffusion 10 -1618 10 -1618 0 cellNo=797
rlabel pdiffusion 17 -1618 17 -1618 0 feedthrough
rlabel pdiffusion 24 -1618 24 -1618 0 feedthrough
rlabel pdiffusion 31 -1618 31 -1618 0 feedthrough
rlabel pdiffusion 38 -1618 38 -1618 0 feedthrough
rlabel pdiffusion 45 -1618 45 -1618 0 feedthrough
rlabel pdiffusion 52 -1618 52 -1618 0 feedthrough
rlabel pdiffusion 59 -1618 59 -1618 0 cellNo=132
rlabel pdiffusion 66 -1618 66 -1618 0 feedthrough
rlabel pdiffusion 73 -1618 73 -1618 0 feedthrough
rlabel pdiffusion 80 -1618 80 -1618 0 feedthrough
rlabel pdiffusion 87 -1618 87 -1618 0 feedthrough
rlabel pdiffusion 94 -1618 94 -1618 0 cellNo=995
rlabel pdiffusion 101 -1618 101 -1618 0 feedthrough
rlabel pdiffusion 108 -1618 108 -1618 0 cellNo=402
rlabel pdiffusion 122 -1618 122 -1618 0 cellNo=128
rlabel pdiffusion 129 -1618 129 -1618 0 feedthrough
rlabel pdiffusion 136 -1618 136 -1618 0 feedthrough
rlabel pdiffusion 143 -1618 143 -1618 0 feedthrough
rlabel pdiffusion 150 -1618 150 -1618 0 feedthrough
rlabel pdiffusion 157 -1618 157 -1618 0 cellNo=987
rlabel pdiffusion 164 -1618 164 -1618 0 cellNo=952
rlabel pdiffusion 171 -1618 171 -1618 0 cellNo=599
rlabel pdiffusion 178 -1618 178 -1618 0 feedthrough
rlabel pdiffusion 185 -1618 185 -1618 0 cellNo=609
rlabel pdiffusion 192 -1618 192 -1618 0 cellNo=1
rlabel pdiffusion 199 -1618 199 -1618 0 feedthrough
rlabel pdiffusion 206 -1618 206 -1618 0 cellNo=698
rlabel pdiffusion 213 -1618 213 -1618 0 feedthrough
rlabel pdiffusion 220 -1618 220 -1618 0 feedthrough
rlabel pdiffusion 227 -1618 227 -1618 0 feedthrough
rlabel pdiffusion 234 -1618 234 -1618 0 feedthrough
rlabel pdiffusion 241 -1618 241 -1618 0 feedthrough
rlabel pdiffusion 248 -1618 248 -1618 0 feedthrough
rlabel pdiffusion 255 -1618 255 -1618 0 feedthrough
rlabel pdiffusion 262 -1618 262 -1618 0 feedthrough
rlabel pdiffusion 269 -1618 269 -1618 0 feedthrough
rlabel pdiffusion 276 -1618 276 -1618 0 feedthrough
rlabel pdiffusion 283 -1618 283 -1618 0 feedthrough
rlabel pdiffusion 290 -1618 290 -1618 0 cellNo=89
rlabel pdiffusion 297 -1618 297 -1618 0 feedthrough
rlabel pdiffusion 304 -1618 304 -1618 0 feedthrough
rlabel pdiffusion 311 -1618 311 -1618 0 feedthrough
rlabel pdiffusion 318 -1618 318 -1618 0 feedthrough
rlabel pdiffusion 325 -1618 325 -1618 0 feedthrough
rlabel pdiffusion 332 -1618 332 -1618 0 feedthrough
rlabel pdiffusion 339 -1618 339 -1618 0 cellNo=447
rlabel pdiffusion 346 -1618 346 -1618 0 cellNo=46
rlabel pdiffusion 353 -1618 353 -1618 0 feedthrough
rlabel pdiffusion 360 -1618 360 -1618 0 cellNo=488
rlabel pdiffusion 367 -1618 367 -1618 0 feedthrough
rlabel pdiffusion 374 -1618 374 -1618 0 feedthrough
rlabel pdiffusion 381 -1618 381 -1618 0 cellNo=688
rlabel pdiffusion 388 -1618 388 -1618 0 feedthrough
rlabel pdiffusion 395 -1618 395 -1618 0 feedthrough
rlabel pdiffusion 402 -1618 402 -1618 0 feedthrough
rlabel pdiffusion 409 -1618 409 -1618 0 feedthrough
rlabel pdiffusion 416 -1618 416 -1618 0 feedthrough
rlabel pdiffusion 423 -1618 423 -1618 0 cellNo=61
rlabel pdiffusion 430 -1618 430 -1618 0 feedthrough
rlabel pdiffusion 437 -1618 437 -1618 0 feedthrough
rlabel pdiffusion 444 -1618 444 -1618 0 feedthrough
rlabel pdiffusion 451 -1618 451 -1618 0 cellNo=76
rlabel pdiffusion 458 -1618 458 -1618 0 feedthrough
rlabel pdiffusion 465 -1618 465 -1618 0 feedthrough
rlabel pdiffusion 472 -1618 472 -1618 0 feedthrough
rlabel pdiffusion 479 -1618 479 -1618 0 cellNo=414
rlabel pdiffusion 486 -1618 486 -1618 0 feedthrough
rlabel pdiffusion 493 -1618 493 -1618 0 cellNo=71
rlabel pdiffusion 500 -1618 500 -1618 0 feedthrough
rlabel pdiffusion 507 -1618 507 -1618 0 feedthrough
rlabel pdiffusion 514 -1618 514 -1618 0 feedthrough
rlabel pdiffusion 521 -1618 521 -1618 0 feedthrough
rlabel pdiffusion 528 -1618 528 -1618 0 cellNo=820
rlabel pdiffusion 535 -1618 535 -1618 0 cellNo=824
rlabel pdiffusion 542 -1618 542 -1618 0 feedthrough
rlabel pdiffusion 549 -1618 549 -1618 0 feedthrough
rlabel pdiffusion 556 -1618 556 -1618 0 feedthrough
rlabel pdiffusion 563 -1618 563 -1618 0 cellNo=170
rlabel pdiffusion 570 -1618 570 -1618 0 feedthrough
rlabel pdiffusion 577 -1618 577 -1618 0 feedthrough
rlabel pdiffusion 584 -1618 584 -1618 0 cellNo=815
rlabel pdiffusion 591 -1618 591 -1618 0 feedthrough
rlabel pdiffusion 598 -1618 598 -1618 0 feedthrough
rlabel pdiffusion 605 -1618 605 -1618 0 feedthrough
rlabel pdiffusion 612 -1618 612 -1618 0 feedthrough
rlabel pdiffusion 626 -1618 626 -1618 0 feedthrough
rlabel pdiffusion 633 -1618 633 -1618 0 feedthrough
rlabel pdiffusion 640 -1618 640 -1618 0 feedthrough
rlabel pdiffusion 647 -1618 647 -1618 0 feedthrough
rlabel pdiffusion 654 -1618 654 -1618 0 feedthrough
rlabel pdiffusion 661 -1618 661 -1618 0 feedthrough
rlabel pdiffusion 668 -1618 668 -1618 0 cellNo=395
rlabel pdiffusion 675 -1618 675 -1618 0 feedthrough
rlabel pdiffusion 682 -1618 682 -1618 0 feedthrough
rlabel pdiffusion 689 -1618 689 -1618 0 feedthrough
rlabel pdiffusion 696 -1618 696 -1618 0 feedthrough
rlabel pdiffusion 703 -1618 703 -1618 0 cellNo=337
rlabel pdiffusion 710 -1618 710 -1618 0 feedthrough
rlabel pdiffusion 717 -1618 717 -1618 0 feedthrough
rlabel pdiffusion 724 -1618 724 -1618 0 feedthrough
rlabel pdiffusion 731 -1618 731 -1618 0 cellNo=135
rlabel pdiffusion 745 -1618 745 -1618 0 feedthrough
rlabel pdiffusion 752 -1618 752 -1618 0 feedthrough
rlabel pdiffusion 759 -1618 759 -1618 0 feedthrough
rlabel pdiffusion 766 -1618 766 -1618 0 feedthrough
rlabel pdiffusion 787 -1618 787 -1618 0 feedthrough
rlabel pdiffusion 794 -1618 794 -1618 0 feedthrough
rlabel pdiffusion 801 -1618 801 -1618 0 feedthrough
rlabel pdiffusion 815 -1618 815 -1618 0 feedthrough
rlabel pdiffusion 829 -1618 829 -1618 0 feedthrough
rlabel pdiffusion 843 -1618 843 -1618 0 feedthrough
rlabel pdiffusion 850 -1618 850 -1618 0 cellNo=446
rlabel pdiffusion 857 -1618 857 -1618 0 feedthrough
rlabel pdiffusion 871 -1618 871 -1618 0 feedthrough
rlabel pdiffusion 878 -1618 878 -1618 0 cellNo=964
rlabel pdiffusion 899 -1618 899 -1618 0 feedthrough
rlabel pdiffusion 913 -1618 913 -1618 0 cellNo=75
rlabel pdiffusion 920 -1618 920 -1618 0 feedthrough
rlabel pdiffusion 927 -1618 927 -1618 0 feedthrough
rlabel pdiffusion 941 -1618 941 -1618 0 cellNo=212
rlabel pdiffusion 948 -1618 948 -1618 0 feedthrough
rlabel pdiffusion 955 -1618 955 -1618 0 feedthrough
rlabel pdiffusion 969 -1618 969 -1618 0 cellNo=810
rlabel pdiffusion 976 -1618 976 -1618 0 feedthrough
rlabel pdiffusion 983 -1618 983 -1618 0 feedthrough
rlabel pdiffusion 10 -1711 10 -1711 0 feedthrough
rlabel pdiffusion 17 -1711 17 -1711 0 cellNo=720
rlabel pdiffusion 24 -1711 24 -1711 0 feedthrough
rlabel pdiffusion 31 -1711 31 -1711 0 feedthrough
rlabel pdiffusion 38 -1711 38 -1711 0 feedthrough
rlabel pdiffusion 45 -1711 45 -1711 0 feedthrough
rlabel pdiffusion 52 -1711 52 -1711 0 feedthrough
rlabel pdiffusion 59 -1711 59 -1711 0 cellNo=904
rlabel pdiffusion 66 -1711 66 -1711 0 feedthrough
rlabel pdiffusion 73 -1711 73 -1711 0 cellNo=156
rlabel pdiffusion 80 -1711 80 -1711 0 feedthrough
rlabel pdiffusion 87 -1711 87 -1711 0 feedthrough
rlabel pdiffusion 94 -1711 94 -1711 0 feedthrough
rlabel pdiffusion 101 -1711 101 -1711 0 cellNo=837
rlabel pdiffusion 108 -1711 108 -1711 0 feedthrough
rlabel pdiffusion 115 -1711 115 -1711 0 cellNo=592
rlabel pdiffusion 122 -1711 122 -1711 0 feedthrough
rlabel pdiffusion 129 -1711 129 -1711 0 feedthrough
rlabel pdiffusion 136 -1711 136 -1711 0 feedthrough
rlabel pdiffusion 143 -1711 143 -1711 0 cellNo=571
rlabel pdiffusion 150 -1711 150 -1711 0 cellNo=142
rlabel pdiffusion 157 -1711 157 -1711 0 feedthrough
rlabel pdiffusion 164 -1711 164 -1711 0 feedthrough
rlabel pdiffusion 171 -1711 171 -1711 0 cellNo=895
rlabel pdiffusion 178 -1711 178 -1711 0 cellNo=976
rlabel pdiffusion 185 -1711 185 -1711 0 feedthrough
rlabel pdiffusion 192 -1711 192 -1711 0 feedthrough
rlabel pdiffusion 199 -1711 199 -1711 0 feedthrough
rlabel pdiffusion 206 -1711 206 -1711 0 cellNo=530
rlabel pdiffusion 213 -1711 213 -1711 0 feedthrough
rlabel pdiffusion 220 -1711 220 -1711 0 feedthrough
rlabel pdiffusion 227 -1711 227 -1711 0 feedthrough
rlabel pdiffusion 234 -1711 234 -1711 0 cellNo=981
rlabel pdiffusion 241 -1711 241 -1711 0 feedthrough
rlabel pdiffusion 248 -1711 248 -1711 0 feedthrough
rlabel pdiffusion 255 -1711 255 -1711 0 feedthrough
rlabel pdiffusion 262 -1711 262 -1711 0 feedthrough
rlabel pdiffusion 269 -1711 269 -1711 0 feedthrough
rlabel pdiffusion 276 -1711 276 -1711 0 feedthrough
rlabel pdiffusion 283 -1711 283 -1711 0 feedthrough
rlabel pdiffusion 290 -1711 290 -1711 0 feedthrough
rlabel pdiffusion 297 -1711 297 -1711 0 cellNo=544
rlabel pdiffusion 304 -1711 304 -1711 0 feedthrough
rlabel pdiffusion 311 -1711 311 -1711 0 feedthrough
rlabel pdiffusion 318 -1711 318 -1711 0 feedthrough
rlabel pdiffusion 325 -1711 325 -1711 0 feedthrough
rlabel pdiffusion 332 -1711 332 -1711 0 cellNo=663
rlabel pdiffusion 339 -1711 339 -1711 0 cellNo=872
rlabel pdiffusion 346 -1711 346 -1711 0 feedthrough
rlabel pdiffusion 353 -1711 353 -1711 0 feedthrough
rlabel pdiffusion 360 -1711 360 -1711 0 feedthrough
rlabel pdiffusion 367 -1711 367 -1711 0 feedthrough
rlabel pdiffusion 374 -1711 374 -1711 0 cellNo=929
rlabel pdiffusion 381 -1711 381 -1711 0 feedthrough
rlabel pdiffusion 388 -1711 388 -1711 0 cellNo=868
rlabel pdiffusion 395 -1711 395 -1711 0 cellNo=58
rlabel pdiffusion 402 -1711 402 -1711 0 cellNo=561
rlabel pdiffusion 409 -1711 409 -1711 0 feedthrough
rlabel pdiffusion 416 -1711 416 -1711 0 feedthrough
rlabel pdiffusion 423 -1711 423 -1711 0 feedthrough
rlabel pdiffusion 430 -1711 430 -1711 0 feedthrough
rlabel pdiffusion 437 -1711 437 -1711 0 cellNo=57
rlabel pdiffusion 444 -1711 444 -1711 0 feedthrough
rlabel pdiffusion 451 -1711 451 -1711 0 cellNo=590
rlabel pdiffusion 458 -1711 458 -1711 0 feedthrough
rlabel pdiffusion 465 -1711 465 -1711 0 cellNo=64
rlabel pdiffusion 472 -1711 472 -1711 0 feedthrough
rlabel pdiffusion 479 -1711 479 -1711 0 feedthrough
rlabel pdiffusion 486 -1711 486 -1711 0 cellNo=628
rlabel pdiffusion 493 -1711 493 -1711 0 feedthrough
rlabel pdiffusion 500 -1711 500 -1711 0 feedthrough
rlabel pdiffusion 507 -1711 507 -1711 0 cellNo=961
rlabel pdiffusion 514 -1711 514 -1711 0 feedthrough
rlabel pdiffusion 521 -1711 521 -1711 0 feedthrough
rlabel pdiffusion 528 -1711 528 -1711 0 feedthrough
rlabel pdiffusion 535 -1711 535 -1711 0 feedthrough
rlabel pdiffusion 542 -1711 542 -1711 0 cellNo=251
rlabel pdiffusion 549 -1711 549 -1711 0 feedthrough
rlabel pdiffusion 556 -1711 556 -1711 0 feedthrough
rlabel pdiffusion 563 -1711 563 -1711 0 feedthrough
rlabel pdiffusion 570 -1711 570 -1711 0 cellNo=766
rlabel pdiffusion 577 -1711 577 -1711 0 feedthrough
rlabel pdiffusion 584 -1711 584 -1711 0 feedthrough
rlabel pdiffusion 591 -1711 591 -1711 0 feedthrough
rlabel pdiffusion 598 -1711 598 -1711 0 feedthrough
rlabel pdiffusion 605 -1711 605 -1711 0 feedthrough
rlabel pdiffusion 612 -1711 612 -1711 0 feedthrough
rlabel pdiffusion 619 -1711 619 -1711 0 feedthrough
rlabel pdiffusion 626 -1711 626 -1711 0 feedthrough
rlabel pdiffusion 633 -1711 633 -1711 0 feedthrough
rlabel pdiffusion 640 -1711 640 -1711 0 feedthrough
rlabel pdiffusion 647 -1711 647 -1711 0 feedthrough
rlabel pdiffusion 654 -1711 654 -1711 0 feedthrough
rlabel pdiffusion 661 -1711 661 -1711 0 cellNo=938
rlabel pdiffusion 668 -1711 668 -1711 0 feedthrough
rlabel pdiffusion 675 -1711 675 -1711 0 feedthrough
rlabel pdiffusion 682 -1711 682 -1711 0 feedthrough
rlabel pdiffusion 689 -1711 689 -1711 0 feedthrough
rlabel pdiffusion 696 -1711 696 -1711 0 feedthrough
rlabel pdiffusion 703 -1711 703 -1711 0 feedthrough
rlabel pdiffusion 710 -1711 710 -1711 0 cellNo=293
rlabel pdiffusion 717 -1711 717 -1711 0 feedthrough
rlabel pdiffusion 724 -1711 724 -1711 0 feedthrough
rlabel pdiffusion 731 -1711 731 -1711 0 feedthrough
rlabel pdiffusion 738 -1711 738 -1711 0 feedthrough
rlabel pdiffusion 745 -1711 745 -1711 0 feedthrough
rlabel pdiffusion 752 -1711 752 -1711 0 feedthrough
rlabel pdiffusion 759 -1711 759 -1711 0 feedthrough
rlabel pdiffusion 766 -1711 766 -1711 0 feedthrough
rlabel pdiffusion 773 -1711 773 -1711 0 feedthrough
rlabel pdiffusion 780 -1711 780 -1711 0 feedthrough
rlabel pdiffusion 787 -1711 787 -1711 0 feedthrough
rlabel pdiffusion 801 -1711 801 -1711 0 feedthrough
rlabel pdiffusion 815 -1711 815 -1711 0 feedthrough
rlabel pdiffusion 822 -1711 822 -1711 0 feedthrough
rlabel pdiffusion 829 -1711 829 -1711 0 feedthrough
rlabel pdiffusion 836 -1711 836 -1711 0 feedthrough
rlabel pdiffusion 843 -1711 843 -1711 0 feedthrough
rlabel pdiffusion 864 -1711 864 -1711 0 feedthrough
rlabel pdiffusion 871 -1711 871 -1711 0 feedthrough
rlabel pdiffusion 885 -1711 885 -1711 0 cellNo=136
rlabel pdiffusion 892 -1711 892 -1711 0 cellNo=535
rlabel pdiffusion 913 -1711 913 -1711 0 feedthrough
rlabel pdiffusion 927 -1711 927 -1711 0 feedthrough
rlabel pdiffusion 941 -1711 941 -1711 0 cellNo=930
rlabel pdiffusion 962 -1711 962 -1711 0 feedthrough
rlabel pdiffusion 969 -1711 969 -1711 0 cellNo=937
rlabel pdiffusion 976 -1711 976 -1711 0 cellNo=376
rlabel pdiffusion 10 -1806 10 -1806 0 cellNo=404
rlabel pdiffusion 17 -1806 17 -1806 0 feedthrough
rlabel pdiffusion 24 -1806 24 -1806 0 feedthrough
rlabel pdiffusion 31 -1806 31 -1806 0 feedthrough
rlabel pdiffusion 38 -1806 38 -1806 0 cellNo=971
rlabel pdiffusion 45 -1806 45 -1806 0 feedthrough
rlabel pdiffusion 52 -1806 52 -1806 0 cellNo=364
rlabel pdiffusion 59 -1806 59 -1806 0 feedthrough
rlabel pdiffusion 66 -1806 66 -1806 0 feedthrough
rlabel pdiffusion 73 -1806 73 -1806 0 feedthrough
rlabel pdiffusion 80 -1806 80 -1806 0 cellNo=181
rlabel pdiffusion 87 -1806 87 -1806 0 cellNo=6
rlabel pdiffusion 94 -1806 94 -1806 0 feedthrough
rlabel pdiffusion 101 -1806 101 -1806 0 cellNo=811
rlabel pdiffusion 108 -1806 108 -1806 0 feedthrough
rlabel pdiffusion 115 -1806 115 -1806 0 cellNo=419
rlabel pdiffusion 122 -1806 122 -1806 0 cellNo=549
rlabel pdiffusion 129 -1806 129 -1806 0 cellNo=20
rlabel pdiffusion 136 -1806 136 -1806 0 cellNo=640
rlabel pdiffusion 143 -1806 143 -1806 0 feedthrough
rlabel pdiffusion 150 -1806 150 -1806 0 feedthrough
rlabel pdiffusion 157 -1806 157 -1806 0 cellNo=389
rlabel pdiffusion 164 -1806 164 -1806 0 cellNo=764
rlabel pdiffusion 171 -1806 171 -1806 0 cellNo=556
rlabel pdiffusion 178 -1806 178 -1806 0 cellNo=338
rlabel pdiffusion 185 -1806 185 -1806 0 cellNo=656
rlabel pdiffusion 192 -1806 192 -1806 0 feedthrough
rlabel pdiffusion 199 -1806 199 -1806 0 feedthrough
rlabel pdiffusion 206 -1806 206 -1806 0 feedthrough
rlabel pdiffusion 213 -1806 213 -1806 0 cellNo=248
rlabel pdiffusion 220 -1806 220 -1806 0 cellNo=167
rlabel pdiffusion 227 -1806 227 -1806 0 feedthrough
rlabel pdiffusion 234 -1806 234 -1806 0 feedthrough
rlabel pdiffusion 241 -1806 241 -1806 0 feedthrough
rlabel pdiffusion 248 -1806 248 -1806 0 feedthrough
rlabel pdiffusion 255 -1806 255 -1806 0 feedthrough
rlabel pdiffusion 262 -1806 262 -1806 0 feedthrough
rlabel pdiffusion 269 -1806 269 -1806 0 cellNo=916
rlabel pdiffusion 276 -1806 276 -1806 0 feedthrough
rlabel pdiffusion 283 -1806 283 -1806 0 feedthrough
rlabel pdiffusion 290 -1806 290 -1806 0 feedthrough
rlabel pdiffusion 297 -1806 297 -1806 0 feedthrough
rlabel pdiffusion 304 -1806 304 -1806 0 feedthrough
rlabel pdiffusion 311 -1806 311 -1806 0 feedthrough
rlabel pdiffusion 318 -1806 318 -1806 0 cellNo=996
rlabel pdiffusion 325 -1806 325 -1806 0 feedthrough
rlabel pdiffusion 332 -1806 332 -1806 0 feedthrough
rlabel pdiffusion 339 -1806 339 -1806 0 feedthrough
rlabel pdiffusion 346 -1806 346 -1806 0 feedthrough
rlabel pdiffusion 353 -1806 353 -1806 0 cellNo=939
rlabel pdiffusion 360 -1806 360 -1806 0 feedthrough
rlabel pdiffusion 367 -1806 367 -1806 0 cellNo=516
rlabel pdiffusion 374 -1806 374 -1806 0 cellNo=267
rlabel pdiffusion 381 -1806 381 -1806 0 cellNo=570
rlabel pdiffusion 388 -1806 388 -1806 0 feedthrough
rlabel pdiffusion 395 -1806 395 -1806 0 cellNo=491
rlabel pdiffusion 402 -1806 402 -1806 0 feedthrough
rlabel pdiffusion 409 -1806 409 -1806 0 feedthrough
rlabel pdiffusion 416 -1806 416 -1806 0 feedthrough
rlabel pdiffusion 423 -1806 423 -1806 0 feedthrough
rlabel pdiffusion 430 -1806 430 -1806 0 feedthrough
rlabel pdiffusion 437 -1806 437 -1806 0 feedthrough
rlabel pdiffusion 444 -1806 444 -1806 0 feedthrough
rlabel pdiffusion 451 -1806 451 -1806 0 feedthrough
rlabel pdiffusion 458 -1806 458 -1806 0 feedthrough
rlabel pdiffusion 465 -1806 465 -1806 0 feedthrough
rlabel pdiffusion 472 -1806 472 -1806 0 cellNo=265
rlabel pdiffusion 479 -1806 479 -1806 0 feedthrough
rlabel pdiffusion 486 -1806 486 -1806 0 feedthrough
rlabel pdiffusion 493 -1806 493 -1806 0 cellNo=183
rlabel pdiffusion 500 -1806 500 -1806 0 cellNo=805
rlabel pdiffusion 507 -1806 507 -1806 0 cellNo=368
rlabel pdiffusion 514 -1806 514 -1806 0 cellNo=769
rlabel pdiffusion 521 -1806 521 -1806 0 cellNo=817
rlabel pdiffusion 528 -1806 528 -1806 0 feedthrough
rlabel pdiffusion 535 -1806 535 -1806 0 feedthrough
rlabel pdiffusion 542 -1806 542 -1806 0 feedthrough
rlabel pdiffusion 549 -1806 549 -1806 0 feedthrough
rlabel pdiffusion 556 -1806 556 -1806 0 feedthrough
rlabel pdiffusion 563 -1806 563 -1806 0 feedthrough
rlabel pdiffusion 570 -1806 570 -1806 0 feedthrough
rlabel pdiffusion 577 -1806 577 -1806 0 feedthrough
rlabel pdiffusion 584 -1806 584 -1806 0 feedthrough
rlabel pdiffusion 591 -1806 591 -1806 0 feedthrough
rlabel pdiffusion 598 -1806 598 -1806 0 feedthrough
rlabel pdiffusion 605 -1806 605 -1806 0 feedthrough
rlabel pdiffusion 612 -1806 612 -1806 0 feedthrough
rlabel pdiffusion 619 -1806 619 -1806 0 feedthrough
rlabel pdiffusion 626 -1806 626 -1806 0 feedthrough
rlabel pdiffusion 633 -1806 633 -1806 0 feedthrough
rlabel pdiffusion 640 -1806 640 -1806 0 cellNo=353
rlabel pdiffusion 647 -1806 647 -1806 0 feedthrough
rlabel pdiffusion 654 -1806 654 -1806 0 feedthrough
rlabel pdiffusion 661 -1806 661 -1806 0 feedthrough
rlabel pdiffusion 668 -1806 668 -1806 0 feedthrough
rlabel pdiffusion 675 -1806 675 -1806 0 feedthrough
rlabel pdiffusion 682 -1806 682 -1806 0 feedthrough
rlabel pdiffusion 689 -1806 689 -1806 0 feedthrough
rlabel pdiffusion 696 -1806 696 -1806 0 feedthrough
rlabel pdiffusion 703 -1806 703 -1806 0 feedthrough
rlabel pdiffusion 710 -1806 710 -1806 0 feedthrough
rlabel pdiffusion 717 -1806 717 -1806 0 feedthrough
rlabel pdiffusion 724 -1806 724 -1806 0 feedthrough
rlabel pdiffusion 731 -1806 731 -1806 0 feedthrough
rlabel pdiffusion 738 -1806 738 -1806 0 feedthrough
rlabel pdiffusion 745 -1806 745 -1806 0 feedthrough
rlabel pdiffusion 752 -1806 752 -1806 0 feedthrough
rlabel pdiffusion 759 -1806 759 -1806 0 feedthrough
rlabel pdiffusion 906 -1806 906 -1806 0 cellNo=653
rlabel pdiffusion 3 -1887 3 -1887 0 cellNo=486
rlabel pdiffusion 10 -1887 10 -1887 0 cellNo=677
rlabel pdiffusion 17 -1887 17 -1887 0 feedthrough
rlabel pdiffusion 24 -1887 24 -1887 0 cellNo=284
rlabel pdiffusion 31 -1887 31 -1887 0 cellNo=629
rlabel pdiffusion 38 -1887 38 -1887 0 feedthrough
rlabel pdiffusion 45 -1887 45 -1887 0 cellNo=280
rlabel pdiffusion 52 -1887 52 -1887 0 feedthrough
rlabel pdiffusion 59 -1887 59 -1887 0 feedthrough
rlabel pdiffusion 66 -1887 66 -1887 0 feedthrough
rlabel pdiffusion 73 -1887 73 -1887 0 feedthrough
rlabel pdiffusion 80 -1887 80 -1887 0 feedthrough
rlabel pdiffusion 87 -1887 87 -1887 0 feedthrough
rlabel pdiffusion 94 -1887 94 -1887 0 feedthrough
rlabel pdiffusion 101 -1887 101 -1887 0 feedthrough
rlabel pdiffusion 108 -1887 108 -1887 0 feedthrough
rlabel pdiffusion 115 -1887 115 -1887 0 feedthrough
rlabel pdiffusion 122 -1887 122 -1887 0 feedthrough
rlabel pdiffusion 129 -1887 129 -1887 0 cellNo=358
rlabel pdiffusion 136 -1887 136 -1887 0 feedthrough
rlabel pdiffusion 143 -1887 143 -1887 0 cellNo=706
rlabel pdiffusion 150 -1887 150 -1887 0 cellNo=932
rlabel pdiffusion 157 -1887 157 -1887 0 feedthrough
rlabel pdiffusion 164 -1887 164 -1887 0 cellNo=526
rlabel pdiffusion 171 -1887 171 -1887 0 cellNo=974
rlabel pdiffusion 178 -1887 178 -1887 0 feedthrough
rlabel pdiffusion 185 -1887 185 -1887 0 feedthrough
rlabel pdiffusion 192 -1887 192 -1887 0 cellNo=179
rlabel pdiffusion 199 -1887 199 -1887 0 cellNo=78
rlabel pdiffusion 206 -1887 206 -1887 0 feedthrough
rlabel pdiffusion 213 -1887 213 -1887 0 feedthrough
rlabel pdiffusion 220 -1887 220 -1887 0 feedthrough
rlabel pdiffusion 227 -1887 227 -1887 0 cellNo=834
rlabel pdiffusion 234 -1887 234 -1887 0 feedthrough
rlabel pdiffusion 241 -1887 241 -1887 0 feedthrough
rlabel pdiffusion 248 -1887 248 -1887 0 feedthrough
rlabel pdiffusion 255 -1887 255 -1887 0 feedthrough
rlabel pdiffusion 262 -1887 262 -1887 0 feedthrough
rlabel pdiffusion 269 -1887 269 -1887 0 feedthrough
rlabel pdiffusion 276 -1887 276 -1887 0 feedthrough
rlabel pdiffusion 283 -1887 283 -1887 0 feedthrough
rlabel pdiffusion 290 -1887 290 -1887 0 cellNo=296
rlabel pdiffusion 297 -1887 297 -1887 0 feedthrough
rlabel pdiffusion 304 -1887 304 -1887 0 cellNo=578
rlabel pdiffusion 311 -1887 311 -1887 0 feedthrough
rlabel pdiffusion 318 -1887 318 -1887 0 feedthrough
rlabel pdiffusion 325 -1887 325 -1887 0 cellNo=222
rlabel pdiffusion 332 -1887 332 -1887 0 feedthrough
rlabel pdiffusion 339 -1887 339 -1887 0 cellNo=320
rlabel pdiffusion 346 -1887 346 -1887 0 cellNo=709
rlabel pdiffusion 353 -1887 353 -1887 0 cellNo=802
rlabel pdiffusion 360 -1887 360 -1887 0 cellNo=417
rlabel pdiffusion 367 -1887 367 -1887 0 feedthrough
rlabel pdiffusion 374 -1887 374 -1887 0 cellNo=47
rlabel pdiffusion 381 -1887 381 -1887 0 feedthrough
rlabel pdiffusion 388 -1887 388 -1887 0 cellNo=747
rlabel pdiffusion 395 -1887 395 -1887 0 feedthrough
rlabel pdiffusion 402 -1887 402 -1887 0 feedthrough
rlabel pdiffusion 409 -1887 409 -1887 0 feedthrough
rlabel pdiffusion 416 -1887 416 -1887 0 feedthrough
rlabel pdiffusion 423 -1887 423 -1887 0 feedthrough
rlabel pdiffusion 430 -1887 430 -1887 0 feedthrough
rlabel pdiffusion 437 -1887 437 -1887 0 cellNo=19
rlabel pdiffusion 444 -1887 444 -1887 0 cellNo=684
rlabel pdiffusion 451 -1887 451 -1887 0 cellNo=632
rlabel pdiffusion 458 -1887 458 -1887 0 feedthrough
rlabel pdiffusion 465 -1887 465 -1887 0 cellNo=978
rlabel pdiffusion 472 -1887 472 -1887 0 feedthrough
rlabel pdiffusion 479 -1887 479 -1887 0 feedthrough
rlabel pdiffusion 486 -1887 486 -1887 0 feedthrough
rlabel pdiffusion 493 -1887 493 -1887 0 feedthrough
rlabel pdiffusion 500 -1887 500 -1887 0 cellNo=408
rlabel pdiffusion 507 -1887 507 -1887 0 feedthrough
rlabel pdiffusion 514 -1887 514 -1887 0 feedthrough
rlabel pdiffusion 521 -1887 521 -1887 0 feedthrough
rlabel pdiffusion 528 -1887 528 -1887 0 feedthrough
rlabel pdiffusion 535 -1887 535 -1887 0 feedthrough
rlabel pdiffusion 542 -1887 542 -1887 0 feedthrough
rlabel pdiffusion 549 -1887 549 -1887 0 cellNo=708
rlabel pdiffusion 556 -1887 556 -1887 0 feedthrough
rlabel pdiffusion 563 -1887 563 -1887 0 feedthrough
rlabel pdiffusion 570 -1887 570 -1887 0 feedthrough
rlabel pdiffusion 577 -1887 577 -1887 0 cellNo=778
rlabel pdiffusion 584 -1887 584 -1887 0 feedthrough
rlabel pdiffusion 591 -1887 591 -1887 0 feedthrough
rlabel pdiffusion 598 -1887 598 -1887 0 feedthrough
rlabel pdiffusion 605 -1887 605 -1887 0 feedthrough
rlabel pdiffusion 612 -1887 612 -1887 0 feedthrough
rlabel pdiffusion 619 -1887 619 -1887 0 feedthrough
rlabel pdiffusion 626 -1887 626 -1887 0 feedthrough
rlabel pdiffusion 633 -1887 633 -1887 0 feedthrough
rlabel pdiffusion 640 -1887 640 -1887 0 cellNo=270
rlabel pdiffusion 647 -1887 647 -1887 0 feedthrough
rlabel pdiffusion 654 -1887 654 -1887 0 feedthrough
rlabel pdiffusion 661 -1887 661 -1887 0 feedthrough
rlabel pdiffusion 668 -1887 668 -1887 0 feedthrough
rlabel pdiffusion 675 -1887 675 -1887 0 feedthrough
rlabel pdiffusion 682 -1887 682 -1887 0 feedthrough
rlabel pdiffusion 689 -1887 689 -1887 0 feedthrough
rlabel pdiffusion 696 -1887 696 -1887 0 feedthrough
rlabel pdiffusion 703 -1887 703 -1887 0 feedthrough
rlabel pdiffusion 710 -1887 710 -1887 0 feedthrough
rlabel pdiffusion 717 -1887 717 -1887 0 feedthrough
rlabel pdiffusion 724 -1887 724 -1887 0 feedthrough
rlabel pdiffusion 731 -1887 731 -1887 0 feedthrough
rlabel pdiffusion 738 -1887 738 -1887 0 feedthrough
rlabel pdiffusion 745 -1887 745 -1887 0 cellNo=583
rlabel pdiffusion 752 -1887 752 -1887 0 feedthrough
rlabel pdiffusion 3 -1970 3 -1970 0 feedthrough
rlabel pdiffusion 10 -1970 10 -1970 0 feedthrough
rlabel pdiffusion 17 -1970 17 -1970 0 cellNo=434
rlabel pdiffusion 24 -1970 24 -1970 0 feedthrough
rlabel pdiffusion 31 -1970 31 -1970 0 cellNo=871
rlabel pdiffusion 38 -1970 38 -1970 0 cellNo=902
rlabel pdiffusion 45 -1970 45 -1970 0 feedthrough
rlabel pdiffusion 52 -1970 52 -1970 0 cellNo=842
rlabel pdiffusion 59 -1970 59 -1970 0 cellNo=60
rlabel pdiffusion 66 -1970 66 -1970 0 feedthrough
rlabel pdiffusion 73 -1970 73 -1970 0 cellNo=678
rlabel pdiffusion 80 -1970 80 -1970 0 cellNo=345
rlabel pdiffusion 87 -1970 87 -1970 0 feedthrough
rlabel pdiffusion 94 -1970 94 -1970 0 feedthrough
rlabel pdiffusion 101 -1970 101 -1970 0 cellNo=883
rlabel pdiffusion 108 -1970 108 -1970 0 cellNo=705
rlabel pdiffusion 115 -1970 115 -1970 0 cellNo=777
rlabel pdiffusion 122 -1970 122 -1970 0 feedthrough
rlabel pdiffusion 129 -1970 129 -1970 0 feedthrough
rlabel pdiffusion 136 -1970 136 -1970 0 feedthrough
rlabel pdiffusion 143 -1970 143 -1970 0 feedthrough
rlabel pdiffusion 150 -1970 150 -1970 0 feedthrough
rlabel pdiffusion 157 -1970 157 -1970 0 cellNo=34
rlabel pdiffusion 164 -1970 164 -1970 0 feedthrough
rlabel pdiffusion 171 -1970 171 -1970 0 cellNo=864
rlabel pdiffusion 178 -1970 178 -1970 0 cellNo=505
rlabel pdiffusion 185 -1970 185 -1970 0 feedthrough
rlabel pdiffusion 192 -1970 192 -1970 0 feedthrough
rlabel pdiffusion 199 -1970 199 -1970 0 cellNo=685
rlabel pdiffusion 206 -1970 206 -1970 0 cellNo=850
rlabel pdiffusion 213 -1970 213 -1970 0 cellNo=825
rlabel pdiffusion 220 -1970 220 -1970 0 cellNo=105
rlabel pdiffusion 227 -1970 227 -1970 0 feedthrough
rlabel pdiffusion 234 -1970 234 -1970 0 feedthrough
rlabel pdiffusion 241 -1970 241 -1970 0 feedthrough
rlabel pdiffusion 248 -1970 248 -1970 0 feedthrough
rlabel pdiffusion 255 -1970 255 -1970 0 feedthrough
rlabel pdiffusion 262 -1970 262 -1970 0 feedthrough
rlabel pdiffusion 269 -1970 269 -1970 0 cellNo=5
rlabel pdiffusion 276 -1970 276 -1970 0 feedthrough
rlabel pdiffusion 283 -1970 283 -1970 0 feedthrough
rlabel pdiffusion 290 -1970 290 -1970 0 feedthrough
rlabel pdiffusion 297 -1970 297 -1970 0 feedthrough
rlabel pdiffusion 304 -1970 304 -1970 0 feedthrough
rlabel pdiffusion 311 -1970 311 -1970 0 cellNo=608
rlabel pdiffusion 318 -1970 318 -1970 0 feedthrough
rlabel pdiffusion 325 -1970 325 -1970 0 feedthrough
rlabel pdiffusion 332 -1970 332 -1970 0 feedthrough
rlabel pdiffusion 339 -1970 339 -1970 0 feedthrough
rlabel pdiffusion 346 -1970 346 -1970 0 cellNo=162
rlabel pdiffusion 353 -1970 353 -1970 0 cellNo=219
rlabel pdiffusion 360 -1970 360 -1970 0 feedthrough
rlabel pdiffusion 367 -1970 367 -1970 0 cellNo=967
rlabel pdiffusion 374 -1970 374 -1970 0 feedthrough
rlabel pdiffusion 381 -1970 381 -1970 0 feedthrough
rlabel pdiffusion 388 -1970 388 -1970 0 cellNo=457
rlabel pdiffusion 395 -1970 395 -1970 0 cellNo=841
rlabel pdiffusion 402 -1970 402 -1970 0 feedthrough
rlabel pdiffusion 409 -1970 409 -1970 0 feedthrough
rlabel pdiffusion 416 -1970 416 -1970 0 cellNo=240
rlabel pdiffusion 423 -1970 423 -1970 0 cellNo=926
rlabel pdiffusion 430 -1970 430 -1970 0 cellNo=977
rlabel pdiffusion 437 -1970 437 -1970 0 feedthrough
rlabel pdiffusion 444 -1970 444 -1970 0 feedthrough
rlabel pdiffusion 451 -1970 451 -1970 0 feedthrough
rlabel pdiffusion 458 -1970 458 -1970 0 cellNo=928
rlabel pdiffusion 465 -1970 465 -1970 0 cellNo=806
rlabel pdiffusion 472 -1970 472 -1970 0 feedthrough
rlabel pdiffusion 479 -1970 479 -1970 0 cellNo=968
rlabel pdiffusion 486 -1970 486 -1970 0 feedthrough
rlabel pdiffusion 493 -1970 493 -1970 0 feedthrough
rlabel pdiffusion 500 -1970 500 -1970 0 feedthrough
rlabel pdiffusion 507 -1970 507 -1970 0 feedthrough
rlabel pdiffusion 514 -1970 514 -1970 0 feedthrough
rlabel pdiffusion 521 -1970 521 -1970 0 feedthrough
rlabel pdiffusion 528 -1970 528 -1970 0 feedthrough
rlabel pdiffusion 535 -1970 535 -1970 0 feedthrough
rlabel pdiffusion 542 -1970 542 -1970 0 feedthrough
rlabel pdiffusion 549 -1970 549 -1970 0 cellNo=832
rlabel pdiffusion 556 -1970 556 -1970 0 feedthrough
rlabel pdiffusion 563 -1970 563 -1970 0 feedthrough
rlabel pdiffusion 570 -1970 570 -1970 0 feedthrough
rlabel pdiffusion 577 -1970 577 -1970 0 feedthrough
rlabel pdiffusion 584 -1970 584 -1970 0 feedthrough
rlabel pdiffusion 591 -1970 591 -1970 0 feedthrough
rlabel pdiffusion 598 -1970 598 -1970 0 feedthrough
rlabel pdiffusion 605 -1970 605 -1970 0 feedthrough
rlabel pdiffusion 612 -1970 612 -1970 0 feedthrough
rlabel pdiffusion 619 -1970 619 -1970 0 feedthrough
rlabel pdiffusion 626 -1970 626 -1970 0 feedthrough
rlabel pdiffusion 633 -1970 633 -1970 0 feedthrough
rlabel pdiffusion 640 -1970 640 -1970 0 cellNo=576
rlabel pdiffusion 647 -1970 647 -1970 0 feedthrough
rlabel pdiffusion 654 -1970 654 -1970 0 feedthrough
rlabel pdiffusion 661 -1970 661 -1970 0 feedthrough
rlabel pdiffusion 668 -1970 668 -1970 0 feedthrough
rlabel pdiffusion 675 -1970 675 -1970 0 feedthrough
rlabel pdiffusion 682 -1970 682 -1970 0 feedthrough
rlabel pdiffusion 689 -1970 689 -1970 0 feedthrough
rlabel pdiffusion 696 -1970 696 -1970 0 feedthrough
rlabel pdiffusion 703 -1970 703 -1970 0 feedthrough
rlabel pdiffusion 710 -1970 710 -1970 0 feedthrough
rlabel pdiffusion 717 -1970 717 -1970 0 feedthrough
rlabel pdiffusion 724 -1970 724 -1970 0 feedthrough
rlabel pdiffusion 731 -1970 731 -1970 0 feedthrough
rlabel pdiffusion 10 -2031 10 -2031 0 feedthrough
rlabel pdiffusion 17 -2031 17 -2031 0 feedthrough
rlabel pdiffusion 24 -2031 24 -2031 0 cellNo=118
rlabel pdiffusion 31 -2031 31 -2031 0 feedthrough
rlabel pdiffusion 38 -2031 38 -2031 0 feedthrough
rlabel pdiffusion 45 -2031 45 -2031 0 feedthrough
rlabel pdiffusion 52 -2031 52 -2031 0 cellNo=120
rlabel pdiffusion 59 -2031 59 -2031 0 feedthrough
rlabel pdiffusion 66 -2031 66 -2031 0 cellNo=72
rlabel pdiffusion 73 -2031 73 -2031 0 feedthrough
rlabel pdiffusion 80 -2031 80 -2031 0 feedthrough
rlabel pdiffusion 87 -2031 87 -2031 0 cellNo=696
rlabel pdiffusion 94 -2031 94 -2031 0 cellNo=12
rlabel pdiffusion 101 -2031 101 -2031 0 cellNo=889
rlabel pdiffusion 108 -2031 108 -2031 0 cellNo=831
rlabel pdiffusion 115 -2031 115 -2031 0 cellNo=710
rlabel pdiffusion 122 -2031 122 -2031 0 feedthrough
rlabel pdiffusion 129 -2031 129 -2031 0 cellNo=555
rlabel pdiffusion 136 -2031 136 -2031 0 feedthrough
rlabel pdiffusion 143 -2031 143 -2031 0 feedthrough
rlabel pdiffusion 150 -2031 150 -2031 0 feedthrough
rlabel pdiffusion 157 -2031 157 -2031 0 feedthrough
rlabel pdiffusion 164 -2031 164 -2031 0 feedthrough
rlabel pdiffusion 171 -2031 171 -2031 0 feedthrough
rlabel pdiffusion 178 -2031 178 -2031 0 feedthrough
rlabel pdiffusion 185 -2031 185 -2031 0 cellNo=716
rlabel pdiffusion 192 -2031 192 -2031 0 cellNo=969
rlabel pdiffusion 199 -2031 199 -2031 0 cellNo=800
rlabel pdiffusion 206 -2031 206 -2031 0 feedthrough
rlabel pdiffusion 213 -2031 213 -2031 0 cellNo=936
rlabel pdiffusion 220 -2031 220 -2031 0 cellNo=272
rlabel pdiffusion 227 -2031 227 -2031 0 feedthrough
rlabel pdiffusion 234 -2031 234 -2031 0 feedthrough
rlabel pdiffusion 241 -2031 241 -2031 0 feedthrough
rlabel pdiffusion 248 -2031 248 -2031 0 cellNo=730
rlabel pdiffusion 255 -2031 255 -2031 0 cellNo=944
rlabel pdiffusion 262 -2031 262 -2031 0 feedthrough
rlabel pdiffusion 269 -2031 269 -2031 0 feedthrough
rlabel pdiffusion 276 -2031 276 -2031 0 feedthrough
rlabel pdiffusion 283 -2031 283 -2031 0 cellNo=39
rlabel pdiffusion 290 -2031 290 -2031 0 feedthrough
rlabel pdiffusion 297 -2031 297 -2031 0 feedthrough
rlabel pdiffusion 304 -2031 304 -2031 0 cellNo=700
rlabel pdiffusion 311 -2031 311 -2031 0 feedthrough
rlabel pdiffusion 318 -2031 318 -2031 0 feedthrough
rlabel pdiffusion 325 -2031 325 -2031 0 feedthrough
rlabel pdiffusion 332 -2031 332 -2031 0 feedthrough
rlabel pdiffusion 339 -2031 339 -2031 0 feedthrough
rlabel pdiffusion 346 -2031 346 -2031 0 feedthrough
rlabel pdiffusion 353 -2031 353 -2031 0 feedthrough
rlabel pdiffusion 360 -2031 360 -2031 0 feedthrough
rlabel pdiffusion 367 -2031 367 -2031 0 feedthrough
rlabel pdiffusion 374 -2031 374 -2031 0 feedthrough
rlabel pdiffusion 381 -2031 381 -2031 0 cellNo=794
rlabel pdiffusion 388 -2031 388 -2031 0 feedthrough
rlabel pdiffusion 395 -2031 395 -2031 0 feedthrough
rlabel pdiffusion 402 -2031 402 -2031 0 cellNo=374
rlabel pdiffusion 409 -2031 409 -2031 0 feedthrough
rlabel pdiffusion 416 -2031 416 -2031 0 cellNo=564
rlabel pdiffusion 423 -2031 423 -2031 0 feedthrough
rlabel pdiffusion 430 -2031 430 -2031 0 feedthrough
rlabel pdiffusion 437 -2031 437 -2031 0 cellNo=949
rlabel pdiffusion 444 -2031 444 -2031 0 feedthrough
rlabel pdiffusion 451 -2031 451 -2031 0 feedthrough
rlabel pdiffusion 458 -2031 458 -2031 0 feedthrough
rlabel pdiffusion 465 -2031 465 -2031 0 feedthrough
rlabel pdiffusion 472 -2031 472 -2031 0 cellNo=411
rlabel pdiffusion 479 -2031 479 -2031 0 feedthrough
rlabel pdiffusion 486 -2031 486 -2031 0 cellNo=302
rlabel pdiffusion 493 -2031 493 -2031 0 feedthrough
rlabel pdiffusion 500 -2031 500 -2031 0 feedthrough
rlabel pdiffusion 507 -2031 507 -2031 0 feedthrough
rlabel pdiffusion 514 -2031 514 -2031 0 feedthrough
rlabel pdiffusion 521 -2031 521 -2031 0 cellNo=728
rlabel pdiffusion 528 -2031 528 -2031 0 feedthrough
rlabel pdiffusion 535 -2031 535 -2031 0 feedthrough
rlabel pdiffusion 542 -2031 542 -2031 0 feedthrough
rlabel pdiffusion 549 -2031 549 -2031 0 cellNo=507
rlabel pdiffusion 556 -2031 556 -2031 0 feedthrough
rlabel pdiffusion 563 -2031 563 -2031 0 feedthrough
rlabel pdiffusion 570 -2031 570 -2031 0 feedthrough
rlabel pdiffusion 577 -2031 577 -2031 0 feedthrough
rlabel pdiffusion 584 -2031 584 -2031 0 feedthrough
rlabel pdiffusion 591 -2031 591 -2031 0 feedthrough
rlabel pdiffusion 598 -2031 598 -2031 0 feedthrough
rlabel pdiffusion 605 -2031 605 -2031 0 feedthrough
rlabel pdiffusion 612 -2031 612 -2031 0 feedthrough
rlabel pdiffusion 619 -2031 619 -2031 0 feedthrough
rlabel pdiffusion 626 -2031 626 -2031 0 feedthrough
rlabel pdiffusion 633 -2031 633 -2031 0 cellNo=819
rlabel pdiffusion 640 -2031 640 -2031 0 cellNo=568
rlabel pdiffusion 647 -2031 647 -2031 0 cellNo=762
rlabel pdiffusion 654 -2031 654 -2031 0 cellNo=853
rlabel pdiffusion 661 -2031 661 -2031 0 feedthrough
rlabel pdiffusion 668 -2031 668 -2031 0 cellNo=129
rlabel pdiffusion 696 -2031 696 -2031 0 feedthrough
rlabel pdiffusion 17 -2096 17 -2096 0 feedthrough
rlabel pdiffusion 24 -2096 24 -2096 0 cellNo=874
rlabel pdiffusion 31 -2096 31 -2096 0 cellNo=886
rlabel pdiffusion 38 -2096 38 -2096 0 feedthrough
rlabel pdiffusion 45 -2096 45 -2096 0 feedthrough
rlabel pdiffusion 52 -2096 52 -2096 0 feedthrough
rlabel pdiffusion 59 -2096 59 -2096 0 cellNo=623
rlabel pdiffusion 66 -2096 66 -2096 0 feedthrough
rlabel pdiffusion 73 -2096 73 -2096 0 cellNo=572
rlabel pdiffusion 80 -2096 80 -2096 0 feedthrough
rlabel pdiffusion 87 -2096 87 -2096 0 feedthrough
rlabel pdiffusion 94 -2096 94 -2096 0 cellNo=511
rlabel pdiffusion 101 -2096 101 -2096 0 feedthrough
rlabel pdiffusion 108 -2096 108 -2096 0 feedthrough
rlabel pdiffusion 115 -2096 115 -2096 0 cellNo=959
rlabel pdiffusion 122 -2096 122 -2096 0 feedthrough
rlabel pdiffusion 129 -2096 129 -2096 0 feedthrough
rlabel pdiffusion 136 -2096 136 -2096 0 feedthrough
rlabel pdiffusion 143 -2096 143 -2096 0 feedthrough
rlabel pdiffusion 150 -2096 150 -2096 0 feedthrough
rlabel pdiffusion 157 -2096 157 -2096 0 cellNo=906
rlabel pdiffusion 164 -2096 164 -2096 0 feedthrough
rlabel pdiffusion 171 -2096 171 -2096 0 feedthrough
rlabel pdiffusion 178 -2096 178 -2096 0 feedthrough
rlabel pdiffusion 185 -2096 185 -2096 0 cellNo=923
rlabel pdiffusion 192 -2096 192 -2096 0 cellNo=796
rlabel pdiffusion 199 -2096 199 -2096 0 feedthrough
rlabel pdiffusion 206 -2096 206 -2096 0 cellNo=562
rlabel pdiffusion 213 -2096 213 -2096 0 feedthrough
rlabel pdiffusion 220 -2096 220 -2096 0 cellNo=626
rlabel pdiffusion 227 -2096 227 -2096 0 feedthrough
rlabel pdiffusion 234 -2096 234 -2096 0 cellNo=648
rlabel pdiffusion 241 -2096 241 -2096 0 feedthrough
rlabel pdiffusion 248 -2096 248 -2096 0 feedthrough
rlabel pdiffusion 255 -2096 255 -2096 0 feedthrough
rlabel pdiffusion 262 -2096 262 -2096 0 feedthrough
rlabel pdiffusion 269 -2096 269 -2096 0 feedthrough
rlabel pdiffusion 276 -2096 276 -2096 0 feedthrough
rlabel pdiffusion 283 -2096 283 -2096 0 feedthrough
rlabel pdiffusion 290 -2096 290 -2096 0 feedthrough
rlabel pdiffusion 297 -2096 297 -2096 0 feedthrough
rlabel pdiffusion 304 -2096 304 -2096 0 cellNo=814
rlabel pdiffusion 311 -2096 311 -2096 0 cellNo=311
rlabel pdiffusion 318 -2096 318 -2096 0 cellNo=602
rlabel pdiffusion 325 -2096 325 -2096 0 cellNo=774
rlabel pdiffusion 332 -2096 332 -2096 0 feedthrough
rlabel pdiffusion 339 -2096 339 -2096 0 feedthrough
rlabel pdiffusion 346 -2096 346 -2096 0 feedthrough
rlabel pdiffusion 353 -2096 353 -2096 0 cellNo=619
rlabel pdiffusion 360 -2096 360 -2096 0 feedthrough
rlabel pdiffusion 367 -2096 367 -2096 0 cellNo=173
rlabel pdiffusion 374 -2096 374 -2096 0 feedthrough
rlabel pdiffusion 381 -2096 381 -2096 0 cellNo=751
rlabel pdiffusion 388 -2096 388 -2096 0 feedthrough
rlabel pdiffusion 395 -2096 395 -2096 0 feedthrough
rlabel pdiffusion 402 -2096 402 -2096 0 cellNo=523
rlabel pdiffusion 409 -2096 409 -2096 0 cellNo=273
rlabel pdiffusion 416 -2096 416 -2096 0 cellNo=691
rlabel pdiffusion 423 -2096 423 -2096 0 cellNo=862
rlabel pdiffusion 430 -2096 430 -2096 0 feedthrough
rlabel pdiffusion 437 -2096 437 -2096 0 feedthrough
rlabel pdiffusion 444 -2096 444 -2096 0 feedthrough
rlabel pdiffusion 451 -2096 451 -2096 0 feedthrough
rlabel pdiffusion 458 -2096 458 -2096 0 feedthrough
rlabel pdiffusion 465 -2096 465 -2096 0 feedthrough
rlabel pdiffusion 472 -2096 472 -2096 0 feedthrough
rlabel pdiffusion 479 -2096 479 -2096 0 cellNo=479
rlabel pdiffusion 486 -2096 486 -2096 0 feedthrough
rlabel pdiffusion 493 -2096 493 -2096 0 feedthrough
rlabel pdiffusion 500 -2096 500 -2096 0 cellNo=63
rlabel pdiffusion 507 -2096 507 -2096 0 feedthrough
rlabel pdiffusion 514 -2096 514 -2096 0 feedthrough
rlabel pdiffusion 521 -2096 521 -2096 0 feedthrough
rlabel pdiffusion 528 -2096 528 -2096 0 feedthrough
rlabel pdiffusion 535 -2096 535 -2096 0 feedthrough
rlabel pdiffusion 542 -2096 542 -2096 0 feedthrough
rlabel pdiffusion 549 -2096 549 -2096 0 feedthrough
rlabel pdiffusion 556 -2096 556 -2096 0 cellNo=193
rlabel pdiffusion 563 -2096 563 -2096 0 feedthrough
rlabel pdiffusion 570 -2096 570 -2096 0 feedthrough
rlabel pdiffusion 577 -2096 577 -2096 0 feedthrough
rlabel pdiffusion 584 -2096 584 -2096 0 feedthrough
rlabel pdiffusion 591 -2096 591 -2096 0 cellNo=452
rlabel pdiffusion 605 -2096 605 -2096 0 feedthrough
rlabel pdiffusion 612 -2096 612 -2096 0 feedthrough
rlabel pdiffusion 619 -2096 619 -2096 0 cellNo=757
rlabel pdiffusion 640 -2096 640 -2096 0 cellNo=857
rlabel pdiffusion 647 -2096 647 -2096 0 feedthrough
rlabel pdiffusion 675 -2096 675 -2096 0 cellNo=893
rlabel pdiffusion 689 -2096 689 -2096 0 feedthrough
rlabel pdiffusion 24 -2153 24 -2153 0 cellNo=600
rlabel pdiffusion 31 -2153 31 -2153 0 cellNo=359
rlabel pdiffusion 38 -2153 38 -2153 0 feedthrough
rlabel pdiffusion 45 -2153 45 -2153 0 feedthrough
rlabel pdiffusion 52 -2153 52 -2153 0 feedthrough
rlabel pdiffusion 59 -2153 59 -2153 0 feedthrough
rlabel pdiffusion 66 -2153 66 -2153 0 feedthrough
rlabel pdiffusion 73 -2153 73 -2153 0 cellNo=585
rlabel pdiffusion 80 -2153 80 -2153 0 cellNo=701
rlabel pdiffusion 87 -2153 87 -2153 0 feedthrough
rlabel pdiffusion 94 -2153 94 -2153 0 cellNo=917
rlabel pdiffusion 101 -2153 101 -2153 0 feedthrough
rlabel pdiffusion 108 -2153 108 -2153 0 feedthrough
rlabel pdiffusion 115 -2153 115 -2153 0 cellNo=70
rlabel pdiffusion 122 -2153 122 -2153 0 cellNo=661
rlabel pdiffusion 129 -2153 129 -2153 0 cellNo=739
rlabel pdiffusion 136 -2153 136 -2153 0 feedthrough
rlabel pdiffusion 143 -2153 143 -2153 0 feedthrough
rlabel pdiffusion 150 -2153 150 -2153 0 cellNo=250
rlabel pdiffusion 157 -2153 157 -2153 0 feedthrough
rlabel pdiffusion 164 -2153 164 -2153 0 feedthrough
rlabel pdiffusion 171 -2153 171 -2153 0 feedthrough
rlabel pdiffusion 178 -2153 178 -2153 0 cellNo=879
rlabel pdiffusion 185 -2153 185 -2153 0 cellNo=644
rlabel pdiffusion 192 -2153 192 -2153 0 feedthrough
rlabel pdiffusion 199 -2153 199 -2153 0 feedthrough
rlabel pdiffusion 206 -2153 206 -2153 0 feedthrough
rlabel pdiffusion 213 -2153 213 -2153 0 cellNo=554
rlabel pdiffusion 220 -2153 220 -2153 0 cellNo=856
rlabel pdiffusion 227 -2153 227 -2153 0 feedthrough
rlabel pdiffusion 234 -2153 234 -2153 0 feedthrough
rlabel pdiffusion 241 -2153 241 -2153 0 feedthrough
rlabel pdiffusion 248 -2153 248 -2153 0 feedthrough
rlabel pdiffusion 255 -2153 255 -2153 0 cellNo=721
rlabel pdiffusion 262 -2153 262 -2153 0 cellNo=963
rlabel pdiffusion 269 -2153 269 -2153 0 feedthrough
rlabel pdiffusion 276 -2153 276 -2153 0 feedthrough
rlabel pdiffusion 283 -2153 283 -2153 0 cellNo=818
rlabel pdiffusion 290 -2153 290 -2153 0 cellNo=994
rlabel pdiffusion 297 -2153 297 -2153 0 feedthrough
rlabel pdiffusion 304 -2153 304 -2153 0 cellNo=858
rlabel pdiffusion 311 -2153 311 -2153 0 feedthrough
rlabel pdiffusion 318 -2153 318 -2153 0 cellNo=605
rlabel pdiffusion 325 -2153 325 -2153 0 feedthrough
rlabel pdiffusion 332 -2153 332 -2153 0 cellNo=827
rlabel pdiffusion 339 -2153 339 -2153 0 cellNo=441
rlabel pdiffusion 346 -2153 346 -2153 0 feedthrough
rlabel pdiffusion 353 -2153 353 -2153 0 feedthrough
rlabel pdiffusion 360 -2153 360 -2153 0 cellNo=683
rlabel pdiffusion 367 -2153 367 -2153 0 cellNo=427
rlabel pdiffusion 374 -2153 374 -2153 0 cellNo=370
rlabel pdiffusion 381 -2153 381 -2153 0 feedthrough
rlabel pdiffusion 388 -2153 388 -2153 0 feedthrough
rlabel pdiffusion 395 -2153 395 -2153 0 feedthrough
rlabel pdiffusion 402 -2153 402 -2153 0 feedthrough
rlabel pdiffusion 409 -2153 409 -2153 0 feedthrough
rlabel pdiffusion 416 -2153 416 -2153 0 cellNo=372
rlabel pdiffusion 423 -2153 423 -2153 0 feedthrough
rlabel pdiffusion 430 -2153 430 -2153 0 feedthrough
rlabel pdiffusion 437 -2153 437 -2153 0 feedthrough
rlabel pdiffusion 444 -2153 444 -2153 0 feedthrough
rlabel pdiffusion 451 -2153 451 -2153 0 feedthrough
rlabel pdiffusion 458 -2153 458 -2153 0 feedthrough
rlabel pdiffusion 465 -2153 465 -2153 0 cellNo=381
rlabel pdiffusion 472 -2153 472 -2153 0 feedthrough
rlabel pdiffusion 479 -2153 479 -2153 0 feedthrough
rlabel pdiffusion 486 -2153 486 -2153 0 feedthrough
rlabel pdiffusion 493 -2153 493 -2153 0 feedthrough
rlabel pdiffusion 500 -2153 500 -2153 0 cellNo=610
rlabel pdiffusion 507 -2153 507 -2153 0 cellNo=933
rlabel pdiffusion 514 -2153 514 -2153 0 feedthrough
rlabel pdiffusion 521 -2153 521 -2153 0 cellNo=313
rlabel pdiffusion 528 -2153 528 -2153 0 cellNo=500
rlabel pdiffusion 535 -2153 535 -2153 0 feedthrough
rlabel pdiffusion 542 -2153 542 -2153 0 feedthrough
rlabel pdiffusion 549 -2153 549 -2153 0 feedthrough
rlabel pdiffusion 556 -2153 556 -2153 0 feedthrough
rlabel pdiffusion 563 -2153 563 -2153 0 feedthrough
rlabel pdiffusion 570 -2153 570 -2153 0 feedthrough
rlabel pdiffusion 591 -2153 591 -2153 0 feedthrough
rlabel pdiffusion 598 -2153 598 -2153 0 feedthrough
rlabel pdiffusion 612 -2153 612 -2153 0 feedthrough
rlabel pdiffusion 10 -2200 10 -2200 0 feedthrough
rlabel pdiffusion 17 -2200 17 -2200 0 cellNo=274
rlabel pdiffusion 24 -2200 24 -2200 0 cellNo=931
rlabel pdiffusion 38 -2200 38 -2200 0 cellNo=522
rlabel pdiffusion 45 -2200 45 -2200 0 cellNo=625
rlabel pdiffusion 52 -2200 52 -2200 0 feedthrough
rlabel pdiffusion 59 -2200 59 -2200 0 feedthrough
rlabel pdiffusion 66 -2200 66 -2200 0 feedthrough
rlabel pdiffusion 73 -2200 73 -2200 0 feedthrough
rlabel pdiffusion 80 -2200 80 -2200 0 feedthrough
rlabel pdiffusion 87 -2200 87 -2200 0 feedthrough
rlabel pdiffusion 94 -2200 94 -2200 0 feedthrough
rlabel pdiffusion 101 -2200 101 -2200 0 feedthrough
rlabel pdiffusion 108 -2200 108 -2200 0 feedthrough
rlabel pdiffusion 115 -2200 115 -2200 0 cellNo=946
rlabel pdiffusion 122 -2200 122 -2200 0 feedthrough
rlabel pdiffusion 129 -2200 129 -2200 0 cellNo=719
rlabel pdiffusion 136 -2200 136 -2200 0 cellNo=597
rlabel pdiffusion 143 -2200 143 -2200 0 cellNo=13
rlabel pdiffusion 150 -2200 150 -2200 0 cellNo=390
rlabel pdiffusion 157 -2200 157 -2200 0 feedthrough
rlabel pdiffusion 164 -2200 164 -2200 0 feedthrough
rlabel pdiffusion 171 -2200 171 -2200 0 feedthrough
rlabel pdiffusion 178 -2200 178 -2200 0 feedthrough
rlabel pdiffusion 185 -2200 185 -2200 0 cellNo=665
rlabel pdiffusion 192 -2200 192 -2200 0 feedthrough
rlabel pdiffusion 199 -2200 199 -2200 0 cellNo=490
rlabel pdiffusion 206 -2200 206 -2200 0 cellNo=901
rlabel pdiffusion 213 -2200 213 -2200 0 cellNo=942
rlabel pdiffusion 220 -2200 220 -2200 0 feedthrough
rlabel pdiffusion 227 -2200 227 -2200 0 feedthrough
rlabel pdiffusion 234 -2200 234 -2200 0 cellNo=985
rlabel pdiffusion 248 -2200 248 -2200 0 feedthrough
rlabel pdiffusion 255 -2200 255 -2200 0 cellNo=435
rlabel pdiffusion 262 -2200 262 -2200 0 feedthrough
rlabel pdiffusion 269 -2200 269 -2200 0 feedthrough
rlabel pdiffusion 276 -2200 276 -2200 0 cellNo=966
rlabel pdiffusion 283 -2200 283 -2200 0 cellNo=305
rlabel pdiffusion 290 -2200 290 -2200 0 feedthrough
rlabel pdiffusion 297 -2200 297 -2200 0 cellNo=615
rlabel pdiffusion 304 -2200 304 -2200 0 feedthrough
rlabel pdiffusion 318 -2200 318 -2200 0 feedthrough
rlabel pdiffusion 325 -2200 325 -2200 0 cellNo=982
rlabel pdiffusion 332 -2200 332 -2200 0 feedthrough
rlabel pdiffusion 346 -2200 346 -2200 0 cellNo=508
rlabel pdiffusion 353 -2200 353 -2200 0 feedthrough
rlabel pdiffusion 360 -2200 360 -2200 0 cellNo=308
rlabel pdiffusion 367 -2200 367 -2200 0 cellNo=733
rlabel pdiffusion 374 -2200 374 -2200 0 cellNo=580
rlabel pdiffusion 381 -2200 381 -2200 0 feedthrough
rlabel pdiffusion 388 -2200 388 -2200 0 feedthrough
rlabel pdiffusion 395 -2200 395 -2200 0 feedthrough
rlabel pdiffusion 402 -2200 402 -2200 0 feedthrough
rlabel pdiffusion 409 -2200 409 -2200 0 feedthrough
rlabel pdiffusion 416 -2200 416 -2200 0 cellNo=812
rlabel pdiffusion 423 -2200 423 -2200 0 cellNo=482
rlabel pdiffusion 430 -2200 430 -2200 0 feedthrough
rlabel pdiffusion 437 -2200 437 -2200 0 feedthrough
rlabel pdiffusion 444 -2200 444 -2200 0 feedthrough
rlabel pdiffusion 451 -2200 451 -2200 0 cellNo=998
rlabel pdiffusion 458 -2200 458 -2200 0 feedthrough
rlabel pdiffusion 465 -2200 465 -2200 0 feedthrough
rlabel pdiffusion 479 -2200 479 -2200 0 cellNo=285
rlabel pdiffusion 493 -2200 493 -2200 0 cellNo=925
rlabel pdiffusion 500 -2200 500 -2200 0 cellNo=892
rlabel pdiffusion 521 -2200 521 -2200 0 feedthrough
rlabel pdiffusion 535 -2200 535 -2200 0 feedthrough
rlabel pdiffusion 549 -2200 549 -2200 0 cellNo=735
rlabel pdiffusion 556 -2200 556 -2200 0 feedthrough
rlabel pdiffusion 598 -2200 598 -2200 0 cellNo=86
rlabel pdiffusion 605 -2200 605 -2200 0 feedthrough
rlabel pdiffusion 612 -2200 612 -2200 0 feedthrough
rlabel pdiffusion 17 -2229 17 -2229 0 cellNo=581
rlabel pdiffusion 24 -2229 24 -2229 0 cellNo=23
rlabel pdiffusion 45 -2229 45 -2229 0 cellNo=439
rlabel pdiffusion 52 -2229 52 -2229 0 cellNo=1000
rlabel pdiffusion 59 -2229 59 -2229 0 feedthrough
rlabel pdiffusion 73 -2229 73 -2229 0 cellNo=999
rlabel pdiffusion 80 -2229 80 -2229 0 cellNo=809
rlabel pdiffusion 94 -2229 94 -2229 0 cellNo=980
rlabel pdiffusion 101 -2229 101 -2229 0 cellNo=772
rlabel pdiffusion 108 -2229 108 -2229 0 feedthrough
rlabel pdiffusion 115 -2229 115 -2229 0 feedthrough
rlabel pdiffusion 129 -2229 129 -2229 0 cellNo=347
rlabel pdiffusion 150 -2229 150 -2229 0 feedthrough
rlabel pdiffusion 164 -2229 164 -2229 0 cellNo=941
rlabel pdiffusion 171 -2229 171 -2229 0 cellNo=538
rlabel pdiffusion 178 -2229 178 -2229 0 cellNo=94
rlabel pdiffusion 185 -2229 185 -2229 0 cellNo=803
rlabel pdiffusion 192 -2229 192 -2229 0 cellNo=56
rlabel pdiffusion 199 -2229 199 -2229 0 cellNo=668
rlabel pdiffusion 206 -2229 206 -2229 0 cellNo=760
rlabel pdiffusion 213 -2229 213 -2229 0 cellNo=788
rlabel pdiffusion 220 -2229 220 -2229 0 cellNo=990
rlabel pdiffusion 227 -2229 227 -2229 0 feedthrough
rlabel pdiffusion 241 -2229 241 -2229 0 feedthrough
rlabel pdiffusion 248 -2229 248 -2229 0 feedthrough
rlabel pdiffusion 255 -2229 255 -2229 0 feedthrough
rlabel pdiffusion 269 -2229 269 -2229 0 feedthrough
rlabel pdiffusion 276 -2229 276 -2229 0 feedthrough
rlabel pdiffusion 283 -2229 283 -2229 0 feedthrough
rlabel pdiffusion 290 -2229 290 -2229 0 feedthrough
rlabel pdiffusion 304 -2229 304 -2229 0 cellNo=727
rlabel pdiffusion 311 -2229 311 -2229 0 cellNo=927
rlabel pdiffusion 325 -2229 325 -2229 0 cellNo=919
rlabel pdiffusion 332 -2229 332 -2229 0 feedthrough
rlabel pdiffusion 339 -2229 339 -2229 0 cellNo=702
rlabel pdiffusion 346 -2229 346 -2229 0 cellNo=139
rlabel pdiffusion 353 -2229 353 -2229 0 cellNo=232
rlabel pdiffusion 374 -2229 374 -2229 0 feedthrough
rlabel pdiffusion 381 -2229 381 -2229 0 cellNo=950
rlabel pdiffusion 388 -2229 388 -2229 0 cellNo=738
rlabel pdiffusion 409 -2229 409 -2229 0 feedthrough
rlabel pdiffusion 430 -2229 430 -2229 0 cellNo=909
rlabel pdiffusion 451 -2229 451 -2229 0 feedthrough
rlabel pdiffusion 472 -2229 472 -2229 0 cellNo=355
rlabel pdiffusion 486 -2229 486 -2229 0 cellNo=424
rlabel pdiffusion 507 -2229 507 -2229 0 feedthrough
rlabel pdiffusion 535 -2229 535 -2229 0 cellNo=898
rlabel pdiffusion 612 -2229 612 -2229 0 cellNo=216
rlabel polysilicon 26 -12 26 -12 0 4
rlabel polysilicon 107 -12 107 -12 0 3
rlabel polysilicon 110 -12 110 -12 0 4
rlabel polysilicon 117 -12 117 -12 0 4
rlabel polysilicon 131 -6 131 -6 0 2
rlabel polysilicon 138 -12 138 -12 0 4
rlabel polysilicon 142 -12 142 -12 0 3
rlabel polysilicon 156 -6 156 -6 0 1
rlabel polysilicon 156 -12 156 -12 0 3
rlabel polysilicon 163 -6 163 -6 0 1
rlabel polysilicon 163 -12 163 -12 0 3
rlabel polysilicon 170 -12 170 -12 0 3
rlabel polysilicon 177 -6 177 -6 0 1
rlabel polysilicon 177 -12 177 -12 0 3
rlabel polysilicon 187 -6 187 -6 0 2
rlabel polysilicon 191 -6 191 -6 0 1
rlabel polysilicon 191 -12 191 -12 0 3
rlabel polysilicon 198 -12 198 -12 0 3
rlabel polysilicon 205 -12 205 -12 0 3
rlabel polysilicon 212 -6 212 -6 0 1
rlabel polysilicon 215 -6 215 -6 0 2
rlabel polysilicon 222 -12 222 -12 0 4
rlabel polysilicon 226 -6 226 -6 0 1
rlabel polysilicon 226 -12 226 -12 0 3
rlabel polysilicon 233 -6 233 -6 0 1
rlabel polysilicon 243 -12 243 -12 0 4
rlabel polysilicon 247 -6 247 -6 0 1
rlabel polysilicon 247 -12 247 -12 0 3
rlabel polysilicon 257 -6 257 -6 0 2
rlabel polysilicon 257 -12 257 -12 0 4
rlabel polysilicon 261 -6 261 -6 0 1
rlabel polysilicon 261 -12 261 -12 0 3
rlabel polysilicon 268 -6 268 -6 0 1
rlabel polysilicon 268 -12 268 -12 0 3
rlabel polysilicon 278 -6 278 -6 0 2
rlabel polysilicon 282 -6 282 -6 0 1
rlabel polysilicon 282 -12 282 -12 0 3
rlabel polysilicon 327 -12 327 -12 0 4
rlabel polysilicon 26 -33 26 -33 0 2
rlabel polysilicon 72 -39 72 -39 0 3
rlabel polysilicon 86 -33 86 -33 0 1
rlabel polysilicon 86 -39 86 -39 0 3
rlabel polysilicon 93 -33 93 -33 0 1
rlabel polysilicon 93 -39 93 -39 0 3
rlabel polysilicon 100 -33 100 -33 0 1
rlabel polysilicon 110 -33 110 -33 0 2
rlabel polysilicon 114 -39 114 -39 0 3
rlabel polysilicon 121 -39 121 -39 0 3
rlabel polysilicon 128 -33 128 -33 0 1
rlabel polysilicon 135 -39 135 -39 0 3
rlabel polysilicon 142 -33 142 -33 0 1
rlabel polysilicon 142 -39 142 -39 0 3
rlabel polysilicon 149 -33 149 -33 0 1
rlabel polysilicon 149 -39 149 -39 0 3
rlabel polysilicon 156 -33 156 -33 0 1
rlabel polysilicon 156 -39 156 -39 0 3
rlabel polysilicon 166 -33 166 -33 0 2
rlabel polysilicon 170 -33 170 -33 0 1
rlabel polysilicon 170 -39 170 -39 0 3
rlabel polysilicon 177 -33 177 -33 0 1
rlabel polysilicon 180 -33 180 -33 0 2
rlabel polysilicon 177 -39 177 -39 0 3
rlabel polysilicon 180 -39 180 -39 0 4
rlabel polysilicon 184 -33 184 -33 0 1
rlabel polysilicon 184 -39 184 -39 0 3
rlabel polysilicon 191 -33 191 -33 0 1
rlabel polysilicon 191 -39 191 -39 0 3
rlabel polysilicon 198 -33 198 -33 0 1
rlabel polysilicon 198 -39 198 -39 0 3
rlabel polysilicon 208 -33 208 -33 0 2
rlabel polysilicon 212 -33 212 -33 0 1
rlabel polysilicon 215 -33 215 -33 0 2
rlabel polysilicon 212 -39 212 -39 0 3
rlabel polysilicon 219 -33 219 -33 0 1
rlabel polysilicon 219 -39 219 -39 0 3
rlabel polysilicon 229 -39 229 -39 0 4
rlabel polysilicon 233 -33 233 -33 0 1
rlabel polysilicon 233 -39 233 -39 0 3
rlabel polysilicon 240 -33 240 -33 0 1
rlabel polysilicon 240 -39 240 -39 0 3
rlabel polysilicon 247 -33 247 -33 0 1
rlabel polysilicon 247 -39 247 -39 0 3
rlabel polysilicon 254 -33 254 -33 0 1
rlabel polysilicon 254 -39 254 -39 0 3
rlabel polysilicon 261 -33 261 -33 0 1
rlabel polysilicon 261 -39 261 -39 0 3
rlabel polysilicon 268 -33 268 -33 0 1
rlabel polysilicon 268 -39 268 -39 0 3
rlabel polysilicon 275 -33 275 -33 0 1
rlabel polysilicon 275 -39 275 -39 0 3
rlabel polysilicon 282 -33 282 -33 0 1
rlabel polysilicon 282 -39 282 -39 0 3
rlabel polysilicon 285 -39 285 -39 0 4
rlabel polysilicon 289 -33 289 -33 0 1
rlabel polysilicon 289 -39 289 -39 0 3
rlabel polysilicon 296 -33 296 -33 0 1
rlabel polysilicon 296 -39 296 -39 0 3
rlabel polysilicon 303 -33 303 -33 0 1
rlabel polysilicon 303 -39 303 -39 0 3
rlabel polysilicon 313 -39 313 -39 0 4
rlabel polysilicon 317 -33 317 -33 0 1
rlabel polysilicon 317 -39 317 -39 0 3
rlabel polysilicon 324 -39 324 -39 0 3
rlabel polysilicon 331 -33 331 -33 0 1
rlabel polysilicon 331 -39 331 -39 0 3
rlabel polysilicon 338 -39 338 -39 0 3
rlabel polysilicon 345 -33 345 -33 0 1
rlabel polysilicon 345 -39 345 -39 0 3
rlabel polysilicon 352 -33 352 -33 0 1
rlabel polysilicon 352 -39 352 -39 0 3
rlabel polysilicon 359 -33 359 -33 0 1
rlabel polysilicon 359 -39 359 -39 0 3
rlabel polysilicon 369 -33 369 -33 0 2
rlabel polysilicon 376 -33 376 -33 0 2
rlabel polysilicon 380 -33 380 -33 0 1
rlabel polysilicon 380 -39 380 -39 0 3
rlabel polysilicon 387 -33 387 -33 0 1
rlabel polysilicon 387 -39 387 -39 0 3
rlabel polysilicon 394 -39 394 -39 0 3
rlabel polysilicon 401 -33 401 -33 0 1
rlabel polysilicon 401 -39 401 -39 0 3
rlabel polysilicon 418 -33 418 -33 0 2
rlabel polysilicon 44 -76 44 -76 0 1
rlabel polysilicon 44 -82 44 -82 0 3
rlabel polysilicon 51 -76 51 -76 0 1
rlabel polysilicon 51 -82 51 -82 0 3
rlabel polysilicon 65 -76 65 -76 0 1
rlabel polysilicon 65 -82 65 -82 0 3
rlabel polysilicon 75 -76 75 -76 0 2
rlabel polysilicon 79 -76 79 -76 0 1
rlabel polysilicon 79 -82 79 -82 0 3
rlabel polysilicon 86 -76 86 -76 0 1
rlabel polysilicon 96 -82 96 -82 0 4
rlabel polysilicon 100 -76 100 -76 0 1
rlabel polysilicon 107 -76 107 -76 0 1
rlabel polysilicon 107 -82 107 -82 0 3
rlabel polysilicon 114 -76 114 -76 0 1
rlabel polysilicon 117 -76 117 -76 0 2
rlabel polysilicon 114 -82 114 -82 0 3
rlabel polysilicon 121 -76 121 -76 0 1
rlabel polysilicon 124 -82 124 -82 0 4
rlabel polysilicon 128 -76 128 -76 0 1
rlabel polysilicon 131 -76 131 -76 0 2
rlabel polysilicon 135 -76 135 -76 0 1
rlabel polysilicon 135 -82 135 -82 0 3
rlabel polysilicon 142 -82 142 -82 0 3
rlabel polysilicon 145 -82 145 -82 0 4
rlabel polysilicon 149 -76 149 -76 0 1
rlabel polysilicon 149 -82 149 -82 0 3
rlabel polysilicon 156 -76 156 -76 0 1
rlabel polysilicon 159 -82 159 -82 0 4
rlabel polysilicon 163 -76 163 -76 0 1
rlabel polysilicon 163 -82 163 -82 0 3
rlabel polysilicon 170 -76 170 -76 0 1
rlabel polysilicon 173 -76 173 -76 0 2
rlabel polysilicon 184 -76 184 -76 0 1
rlabel polysilicon 184 -82 184 -82 0 3
rlabel polysilicon 191 -82 191 -82 0 3
rlabel polysilicon 194 -82 194 -82 0 4
rlabel polysilicon 198 -76 198 -76 0 1
rlabel polysilicon 198 -82 198 -82 0 3
rlabel polysilicon 205 -76 205 -76 0 1
rlabel polysilicon 212 -76 212 -76 0 1
rlabel polysilicon 215 -76 215 -76 0 2
rlabel polysilicon 212 -82 212 -82 0 3
rlabel polysilicon 215 -82 215 -82 0 4
rlabel polysilicon 219 -76 219 -76 0 1
rlabel polysilicon 222 -76 222 -76 0 2
rlabel polysilicon 219 -82 219 -82 0 3
rlabel polysilicon 222 -82 222 -82 0 4
rlabel polysilicon 226 -76 226 -76 0 1
rlabel polysilicon 233 -76 233 -76 0 1
rlabel polysilicon 233 -82 233 -82 0 3
rlabel polysilicon 240 -76 240 -76 0 1
rlabel polysilicon 240 -82 240 -82 0 3
rlabel polysilicon 247 -76 247 -76 0 1
rlabel polysilicon 247 -82 247 -82 0 3
rlabel polysilicon 254 -76 254 -76 0 1
rlabel polysilicon 257 -76 257 -76 0 2
rlabel polysilicon 254 -82 254 -82 0 3
rlabel polysilicon 257 -82 257 -82 0 4
rlabel polysilicon 261 -76 261 -76 0 1
rlabel polysilicon 261 -82 261 -82 0 3
rlabel polysilicon 271 -82 271 -82 0 4
rlabel polysilicon 275 -76 275 -76 0 1
rlabel polysilicon 278 -82 278 -82 0 4
rlabel polysilicon 282 -76 282 -76 0 1
rlabel polysilicon 289 -76 289 -76 0 1
rlabel polysilicon 289 -82 289 -82 0 3
rlabel polysilicon 296 -76 296 -76 0 1
rlabel polysilicon 296 -82 296 -82 0 3
rlabel polysilicon 303 -76 303 -76 0 1
rlabel polysilicon 303 -82 303 -82 0 3
rlabel polysilicon 310 -76 310 -76 0 1
rlabel polysilicon 310 -82 310 -82 0 3
rlabel polysilicon 317 -76 317 -76 0 1
rlabel polysilicon 317 -82 317 -82 0 3
rlabel polysilicon 324 -76 324 -76 0 1
rlabel polysilicon 324 -82 324 -82 0 3
rlabel polysilicon 331 -76 331 -76 0 1
rlabel polysilicon 331 -82 331 -82 0 3
rlabel polysilicon 338 -76 338 -76 0 1
rlabel polysilicon 338 -82 338 -82 0 3
rlabel polysilicon 345 -76 345 -76 0 1
rlabel polysilicon 345 -82 345 -82 0 3
rlabel polysilicon 352 -82 352 -82 0 3
rlabel polysilicon 359 -76 359 -76 0 1
rlabel polysilicon 359 -82 359 -82 0 3
rlabel polysilicon 366 -76 366 -76 0 1
rlabel polysilicon 366 -82 366 -82 0 3
rlabel polysilicon 373 -76 373 -76 0 1
rlabel polysilicon 373 -82 373 -82 0 3
rlabel polysilicon 380 -76 380 -76 0 1
rlabel polysilicon 380 -82 380 -82 0 3
rlabel polysilicon 387 -76 387 -76 0 1
rlabel polysilicon 387 -82 387 -82 0 3
rlabel polysilicon 394 -76 394 -76 0 1
rlabel polysilicon 394 -82 394 -82 0 3
rlabel polysilicon 401 -76 401 -76 0 1
rlabel polysilicon 401 -82 401 -82 0 3
rlabel polysilicon 408 -76 408 -76 0 1
rlabel polysilicon 408 -82 408 -82 0 3
rlabel polysilicon 432 -82 432 -82 0 4
rlabel polysilicon 58 -121 58 -121 0 1
rlabel polysilicon 58 -127 58 -127 0 3
rlabel polysilicon 65 -121 65 -121 0 1
rlabel polysilicon 79 -121 79 -121 0 1
rlabel polysilicon 79 -127 79 -127 0 3
rlabel polysilicon 86 -121 86 -121 0 1
rlabel polysilicon 86 -127 86 -127 0 3
rlabel polysilicon 93 -121 93 -121 0 1
rlabel polysilicon 93 -127 93 -127 0 3
rlabel polysilicon 100 -121 100 -121 0 1
rlabel polysilicon 100 -127 100 -127 0 3
rlabel polysilicon 103 -127 103 -127 0 4
rlabel polysilicon 107 -121 107 -121 0 1
rlabel polysilicon 107 -127 107 -127 0 3
rlabel polysilicon 117 -127 117 -127 0 4
rlabel polysilicon 121 -121 121 -121 0 1
rlabel polysilicon 121 -127 121 -127 0 3
rlabel polysilicon 128 -121 128 -121 0 1
rlabel polysilicon 131 -121 131 -121 0 2
rlabel polysilicon 131 -127 131 -127 0 4
rlabel polysilicon 138 -127 138 -127 0 4
rlabel polysilicon 142 -127 142 -127 0 3
rlabel polysilicon 145 -127 145 -127 0 4
rlabel polysilicon 149 -121 149 -121 0 1
rlabel polysilicon 149 -127 149 -127 0 3
rlabel polysilicon 156 -121 156 -121 0 1
rlabel polysilicon 163 -121 163 -121 0 1
rlabel polysilicon 166 -127 166 -127 0 4
rlabel polysilicon 170 -121 170 -121 0 1
rlabel polysilicon 170 -127 170 -127 0 3
rlabel polysilicon 177 -121 177 -121 0 1
rlabel polysilicon 177 -127 177 -127 0 3
rlabel polysilicon 184 -121 184 -121 0 1
rlabel polysilicon 184 -127 184 -127 0 3
rlabel polysilicon 191 -121 191 -121 0 1
rlabel polysilicon 191 -127 191 -127 0 3
rlabel polysilicon 201 -121 201 -121 0 2
rlabel polysilicon 198 -127 198 -127 0 3
rlabel polysilicon 205 -121 205 -121 0 1
rlabel polysilicon 205 -127 205 -127 0 3
rlabel polysilicon 212 -121 212 -121 0 1
rlabel polysilicon 215 -121 215 -121 0 2
rlabel polysilicon 215 -127 215 -127 0 4
rlabel polysilicon 222 -127 222 -127 0 4
rlabel polysilicon 226 -121 226 -121 0 1
rlabel polysilicon 226 -127 226 -127 0 3
rlabel polysilicon 236 -127 236 -127 0 4
rlabel polysilicon 240 -121 240 -121 0 1
rlabel polysilicon 247 -121 247 -121 0 1
rlabel polysilicon 250 -121 250 -121 0 2
rlabel polysilicon 247 -127 247 -127 0 3
rlabel polysilicon 250 -127 250 -127 0 4
rlabel polysilicon 254 -121 254 -121 0 1
rlabel polysilicon 254 -127 254 -127 0 3
rlabel polysilicon 261 -121 261 -121 0 1
rlabel polysilicon 271 -121 271 -121 0 2
rlabel polysilicon 275 -121 275 -121 0 1
rlabel polysilicon 278 -121 278 -121 0 2
rlabel polysilicon 282 -121 282 -121 0 1
rlabel polysilicon 282 -127 282 -127 0 3
rlabel polysilicon 289 -121 289 -121 0 1
rlabel polysilicon 289 -127 289 -127 0 3
rlabel polysilicon 296 -121 296 -121 0 1
rlabel polysilicon 296 -127 296 -127 0 3
rlabel polysilicon 303 -121 303 -121 0 1
rlabel polysilicon 303 -127 303 -127 0 3
rlabel polysilicon 310 -127 310 -127 0 3
rlabel polysilicon 317 -121 317 -121 0 1
rlabel polysilicon 317 -127 317 -127 0 3
rlabel polysilicon 324 -121 324 -121 0 1
rlabel polysilicon 324 -127 324 -127 0 3
rlabel polysilicon 331 -121 331 -121 0 1
rlabel polysilicon 331 -127 331 -127 0 3
rlabel polysilicon 338 -121 338 -121 0 1
rlabel polysilicon 338 -127 338 -127 0 3
rlabel polysilicon 345 -121 345 -121 0 1
rlabel polysilicon 345 -127 345 -127 0 3
rlabel polysilicon 352 -121 352 -121 0 1
rlabel polysilicon 352 -127 352 -127 0 3
rlabel polysilicon 359 -121 359 -121 0 1
rlabel polysilicon 359 -127 359 -127 0 3
rlabel polysilicon 366 -121 366 -121 0 1
rlabel polysilicon 373 -121 373 -121 0 1
rlabel polysilicon 373 -127 373 -127 0 3
rlabel polysilicon 383 -121 383 -121 0 2
rlabel polysilicon 380 -127 380 -127 0 3
rlabel polysilicon 387 -121 387 -121 0 1
rlabel polysilicon 387 -127 387 -127 0 3
rlabel polysilicon 394 -121 394 -121 0 1
rlabel polysilicon 394 -127 394 -127 0 3
rlabel polysilicon 401 -121 401 -121 0 1
rlabel polysilicon 401 -127 401 -127 0 3
rlabel polysilicon 408 -121 408 -121 0 1
rlabel polysilicon 408 -127 408 -127 0 3
rlabel polysilicon 415 -121 415 -121 0 1
rlabel polysilicon 415 -127 415 -127 0 3
rlabel polysilicon 422 -121 422 -121 0 1
rlabel polysilicon 422 -127 422 -127 0 3
rlabel polysilicon 429 -121 429 -121 0 1
rlabel polysilicon 429 -127 429 -127 0 3
rlabel polysilicon 439 -127 439 -127 0 4
rlabel polysilicon 443 -121 443 -121 0 1
rlabel polysilicon 443 -127 443 -127 0 3
rlabel polysilicon 453 -121 453 -121 0 2
rlabel polysilicon 37 -174 37 -174 0 1
rlabel polysilicon 37 -180 37 -180 0 3
rlabel polysilicon 44 -174 44 -174 0 1
rlabel polysilicon 44 -180 44 -180 0 3
rlabel polysilicon 51 -174 51 -174 0 1
rlabel polysilicon 51 -180 51 -180 0 3
rlabel polysilicon 58 -174 58 -174 0 1
rlabel polysilicon 58 -180 58 -180 0 3
rlabel polysilicon 68 -180 68 -180 0 4
rlabel polysilicon 72 -174 72 -174 0 1
rlabel polysilicon 72 -180 72 -180 0 3
rlabel polysilicon 79 -174 79 -174 0 1
rlabel polysilicon 79 -180 79 -180 0 3
rlabel polysilicon 89 -174 89 -174 0 2
rlabel polysilicon 89 -180 89 -180 0 4
rlabel polysilicon 93 -174 93 -174 0 1
rlabel polysilicon 96 -180 96 -180 0 4
rlabel polysilicon 100 -174 100 -174 0 1
rlabel polysilicon 100 -180 100 -180 0 3
rlabel polysilicon 110 -174 110 -174 0 2
rlabel polysilicon 114 -174 114 -174 0 1
rlabel polysilicon 114 -180 114 -180 0 3
rlabel polysilicon 121 -174 121 -174 0 1
rlabel polysilicon 121 -180 121 -180 0 3
rlabel polysilicon 128 -174 128 -174 0 1
rlabel polysilicon 128 -180 128 -180 0 3
rlabel polysilicon 138 -174 138 -174 0 2
rlabel polysilicon 135 -180 135 -180 0 3
rlabel polysilicon 142 -180 142 -180 0 3
rlabel polysilicon 145 -180 145 -180 0 4
rlabel polysilicon 149 -180 149 -180 0 3
rlabel polysilicon 152 -180 152 -180 0 4
rlabel polysilicon 156 -174 156 -174 0 1
rlabel polysilicon 156 -180 156 -180 0 3
rlabel polysilicon 166 -174 166 -174 0 2
rlabel polysilicon 170 -174 170 -174 0 1
rlabel polysilicon 170 -180 170 -180 0 3
rlabel polysilicon 177 -174 177 -174 0 1
rlabel polysilicon 177 -180 177 -180 0 3
rlabel polysilicon 184 -174 184 -174 0 1
rlabel polysilicon 187 -180 187 -180 0 4
rlabel polysilicon 191 -174 191 -174 0 1
rlabel polysilicon 191 -180 191 -180 0 3
rlabel polysilicon 198 -174 198 -174 0 1
rlabel polysilicon 198 -180 198 -180 0 3
rlabel polysilicon 208 -174 208 -174 0 2
rlabel polysilicon 208 -180 208 -180 0 4
rlabel polysilicon 212 -180 212 -180 0 3
rlabel polysilicon 215 -180 215 -180 0 4
rlabel polysilicon 219 -174 219 -174 0 1
rlabel polysilicon 219 -180 219 -180 0 3
rlabel polysilicon 226 -174 226 -174 0 1
rlabel polysilicon 226 -180 226 -180 0 3
rlabel polysilicon 233 -174 233 -174 0 1
rlabel polysilicon 236 -174 236 -174 0 2
rlabel polysilicon 233 -180 233 -180 0 3
rlabel polysilicon 243 -180 243 -180 0 4
rlabel polysilicon 247 -174 247 -174 0 1
rlabel polysilicon 247 -180 247 -180 0 3
rlabel polysilicon 254 -174 254 -174 0 1
rlabel polysilicon 257 -180 257 -180 0 4
rlabel polysilicon 261 -174 261 -174 0 1
rlabel polysilicon 261 -180 261 -180 0 3
rlabel polysilicon 268 -174 268 -174 0 1
rlabel polysilicon 268 -180 268 -180 0 3
rlabel polysilicon 275 -174 275 -174 0 1
rlabel polysilicon 278 -180 278 -180 0 4
rlabel polysilicon 285 -174 285 -174 0 2
rlabel polysilicon 289 -180 289 -180 0 3
rlabel polysilicon 292 -180 292 -180 0 4
rlabel polysilicon 296 -174 296 -174 0 1
rlabel polysilicon 296 -180 296 -180 0 3
rlabel polysilicon 306 -174 306 -174 0 2
rlabel polysilicon 306 -180 306 -180 0 4
rlabel polysilicon 313 -174 313 -174 0 2
rlabel polysilicon 317 -174 317 -174 0 1
rlabel polysilicon 320 -174 320 -174 0 2
rlabel polysilicon 324 -174 324 -174 0 1
rlabel polysilicon 324 -180 324 -180 0 3
rlabel polysilicon 331 -174 331 -174 0 1
rlabel polysilicon 331 -180 331 -180 0 3
rlabel polysilicon 334 -180 334 -180 0 4
rlabel polysilicon 338 -174 338 -174 0 1
rlabel polysilicon 338 -180 338 -180 0 3
rlabel polysilicon 345 -174 345 -174 0 1
rlabel polysilicon 345 -180 345 -180 0 3
rlabel polysilicon 352 -174 352 -174 0 1
rlabel polysilicon 352 -180 352 -180 0 3
rlabel polysilicon 359 -174 359 -174 0 1
rlabel polysilicon 359 -180 359 -180 0 3
rlabel polysilicon 366 -174 366 -174 0 1
rlabel polysilicon 366 -180 366 -180 0 3
rlabel polysilicon 373 -174 373 -174 0 1
rlabel polysilicon 373 -180 373 -180 0 3
rlabel polysilicon 380 -174 380 -174 0 1
rlabel polysilicon 380 -180 380 -180 0 3
rlabel polysilicon 387 -174 387 -174 0 1
rlabel polysilicon 387 -180 387 -180 0 3
rlabel polysilicon 394 -174 394 -174 0 1
rlabel polysilicon 394 -180 394 -180 0 3
rlabel polysilicon 401 -174 401 -174 0 1
rlabel polysilicon 401 -180 401 -180 0 3
rlabel polysilicon 408 -174 408 -174 0 1
rlabel polysilicon 408 -180 408 -180 0 3
rlabel polysilicon 415 -174 415 -174 0 1
rlabel polysilicon 415 -180 415 -180 0 3
rlabel polysilicon 429 -174 429 -174 0 1
rlabel polysilicon 429 -180 429 -180 0 3
rlabel polysilicon 436 -174 436 -174 0 1
rlabel polysilicon 436 -180 436 -180 0 3
rlabel polysilicon 443 -174 443 -174 0 1
rlabel polysilicon 443 -180 443 -180 0 3
rlabel polysilicon 450 -174 450 -174 0 1
rlabel polysilicon 450 -180 450 -180 0 3
rlabel polysilicon 457 -174 457 -174 0 1
rlabel polysilicon 457 -180 457 -180 0 3
rlabel polysilicon 464 -174 464 -174 0 1
rlabel polysilicon 464 -180 464 -180 0 3
rlabel polysilicon 471 -174 471 -174 0 1
rlabel polysilicon 471 -180 471 -180 0 3
rlabel polysilicon 481 -174 481 -174 0 2
rlabel polysilicon 485 -174 485 -174 0 1
rlabel polysilicon 485 -180 485 -180 0 3
rlabel polysilicon 492 -174 492 -174 0 1
rlabel polysilicon 492 -180 492 -180 0 3
rlabel polysilicon 548 -180 548 -180 0 3
rlabel polysilicon 16 -231 16 -231 0 1
rlabel polysilicon 16 -237 16 -237 0 3
rlabel polysilicon 30 -231 30 -231 0 1
rlabel polysilicon 30 -237 30 -237 0 3
rlabel polysilicon 37 -231 37 -231 0 1
rlabel polysilicon 58 -231 58 -231 0 1
rlabel polysilicon 65 -231 65 -231 0 1
rlabel polysilicon 79 -231 79 -231 0 1
rlabel polysilicon 82 -231 82 -231 0 2
rlabel polysilicon 82 -237 82 -237 0 4
rlabel polysilicon 86 -231 86 -231 0 1
rlabel polysilicon 89 -231 89 -231 0 2
rlabel polysilicon 93 -231 93 -231 0 1
rlabel polysilicon 93 -237 93 -237 0 3
rlabel polysilicon 100 -231 100 -231 0 1
rlabel polysilicon 103 -231 103 -231 0 2
rlabel polysilicon 100 -237 100 -237 0 3
rlabel polysilicon 103 -237 103 -237 0 4
rlabel polysilicon 107 -231 107 -231 0 1
rlabel polysilicon 107 -237 107 -237 0 3
rlabel polysilicon 114 -231 114 -231 0 1
rlabel polysilicon 114 -237 114 -237 0 3
rlabel polysilicon 121 -231 121 -231 0 1
rlabel polysilicon 124 -231 124 -231 0 2
rlabel polysilicon 128 -231 128 -231 0 1
rlabel polysilicon 128 -237 128 -237 0 3
rlabel polysilicon 135 -231 135 -231 0 1
rlabel polysilicon 135 -237 135 -237 0 3
rlabel polysilicon 142 -231 142 -231 0 1
rlabel polysilicon 152 -231 152 -231 0 2
rlabel polysilicon 149 -237 149 -237 0 3
rlabel polysilicon 152 -237 152 -237 0 4
rlabel polysilicon 156 -231 156 -231 0 1
rlabel polysilicon 156 -237 156 -237 0 3
rlabel polysilicon 163 -231 163 -231 0 1
rlabel polysilicon 163 -237 163 -237 0 3
rlabel polysilicon 166 -237 166 -237 0 4
rlabel polysilicon 170 -231 170 -231 0 1
rlabel polysilicon 170 -237 170 -237 0 3
rlabel polysilicon 177 -231 177 -231 0 1
rlabel polysilicon 177 -237 177 -237 0 3
rlabel polysilicon 184 -231 184 -231 0 1
rlabel polysilicon 184 -237 184 -237 0 3
rlabel polysilicon 191 -231 191 -231 0 1
rlabel polysilicon 191 -237 191 -237 0 3
rlabel polysilicon 198 -231 198 -231 0 1
rlabel polysilicon 198 -237 198 -237 0 3
rlabel polysilicon 205 -231 205 -231 0 1
rlabel polysilicon 205 -237 205 -237 0 3
rlabel polysilicon 212 -231 212 -231 0 1
rlabel polysilicon 215 -237 215 -237 0 4
rlabel polysilicon 219 -231 219 -231 0 1
rlabel polysilicon 222 -231 222 -231 0 2
rlabel polysilicon 222 -237 222 -237 0 4
rlabel polysilicon 226 -231 226 -231 0 1
rlabel polysilicon 226 -237 226 -237 0 3
rlabel polysilicon 233 -231 233 -231 0 1
rlabel polysilicon 233 -237 233 -237 0 3
rlabel polysilicon 240 -231 240 -231 0 1
rlabel polysilicon 243 -231 243 -231 0 2
rlabel polysilicon 240 -237 240 -237 0 3
rlabel polysilicon 243 -237 243 -237 0 4
rlabel polysilicon 247 -231 247 -231 0 1
rlabel polysilicon 247 -237 247 -237 0 3
rlabel polysilicon 254 -231 254 -231 0 1
rlabel polysilicon 257 -237 257 -237 0 4
rlabel polysilicon 261 -231 261 -231 0 1
rlabel polysilicon 261 -237 261 -237 0 3
rlabel polysilicon 268 -231 268 -231 0 1
rlabel polysilicon 268 -237 268 -237 0 3
rlabel polysilicon 275 -231 275 -231 0 1
rlabel polysilicon 275 -237 275 -237 0 3
rlabel polysilicon 282 -231 282 -231 0 1
rlabel polysilicon 285 -231 285 -231 0 2
rlabel polysilicon 282 -237 282 -237 0 3
rlabel polysilicon 285 -237 285 -237 0 4
rlabel polysilicon 289 -231 289 -231 0 1
rlabel polysilicon 289 -237 289 -237 0 3
rlabel polysilicon 303 -231 303 -231 0 1
rlabel polysilicon 303 -237 303 -237 0 3
rlabel polysilicon 310 -231 310 -231 0 1
rlabel polysilicon 317 -231 317 -231 0 1
rlabel polysilicon 317 -237 317 -237 0 3
rlabel polysilicon 324 -231 324 -231 0 1
rlabel polysilicon 324 -237 324 -237 0 3
rlabel polysilicon 331 -231 331 -231 0 1
rlabel polysilicon 331 -237 331 -237 0 3
rlabel polysilicon 341 -231 341 -231 0 2
rlabel polysilicon 345 -231 345 -231 0 1
rlabel polysilicon 345 -237 345 -237 0 3
rlabel polysilicon 352 -237 352 -237 0 3
rlabel polysilicon 359 -231 359 -231 0 1
rlabel polysilicon 362 -237 362 -237 0 4
rlabel polysilicon 366 -231 366 -231 0 1
rlabel polysilicon 366 -237 366 -237 0 3
rlabel polysilicon 373 -231 373 -231 0 1
rlabel polysilicon 373 -237 373 -237 0 3
rlabel polysilicon 380 -231 380 -231 0 1
rlabel polysilicon 380 -237 380 -237 0 3
rlabel polysilicon 387 -231 387 -231 0 1
rlabel polysilicon 387 -237 387 -237 0 3
rlabel polysilicon 394 -231 394 -231 0 1
rlabel polysilicon 394 -237 394 -237 0 3
rlabel polysilicon 401 -231 401 -231 0 1
rlabel polysilicon 401 -237 401 -237 0 3
rlabel polysilicon 408 -231 408 -231 0 1
rlabel polysilicon 408 -237 408 -237 0 3
rlabel polysilicon 415 -231 415 -231 0 1
rlabel polysilicon 415 -237 415 -237 0 3
rlabel polysilicon 422 -231 422 -231 0 1
rlabel polysilicon 422 -237 422 -237 0 3
rlabel polysilicon 429 -231 429 -231 0 1
rlabel polysilicon 429 -237 429 -237 0 3
rlabel polysilicon 436 -231 436 -231 0 1
rlabel polysilicon 436 -237 436 -237 0 3
rlabel polysilicon 443 -231 443 -231 0 1
rlabel polysilicon 443 -237 443 -237 0 3
rlabel polysilicon 450 -231 450 -231 0 1
rlabel polysilicon 450 -237 450 -237 0 3
rlabel polysilicon 457 -231 457 -231 0 1
rlabel polysilicon 457 -237 457 -237 0 3
rlabel polysilicon 464 -231 464 -231 0 1
rlabel polysilicon 464 -237 464 -237 0 3
rlabel polysilicon 471 -231 471 -231 0 1
rlabel polysilicon 471 -237 471 -237 0 3
rlabel polysilicon 478 -231 478 -231 0 1
rlabel polysilicon 478 -237 478 -237 0 3
rlabel polysilicon 485 -231 485 -231 0 1
rlabel polysilicon 485 -237 485 -237 0 3
rlabel polysilicon 492 -231 492 -231 0 1
rlabel polysilicon 492 -237 492 -237 0 3
rlabel polysilicon 499 -231 499 -231 0 1
rlabel polysilicon 499 -237 499 -237 0 3
rlabel polysilicon 506 -231 506 -231 0 1
rlabel polysilicon 506 -237 506 -237 0 3
rlabel polysilicon 513 -231 513 -231 0 1
rlabel polysilicon 513 -237 513 -237 0 3
rlabel polysilicon 520 -231 520 -231 0 1
rlabel polysilicon 527 -231 527 -231 0 1
rlabel polysilicon 527 -237 527 -237 0 3
rlabel polysilicon 534 -231 534 -231 0 1
rlabel polysilicon 534 -237 534 -237 0 3
rlabel polysilicon 541 -237 541 -237 0 3
rlabel polysilicon 548 -231 548 -231 0 1
rlabel polysilicon 555 -231 555 -231 0 1
rlabel polysilicon 555 -237 555 -237 0 3
rlabel polysilicon 558 -237 558 -237 0 4
rlabel polysilicon 565 -231 565 -231 0 2
rlabel polysilicon 565 -237 565 -237 0 4
rlabel polysilicon 583 -231 583 -231 0 1
rlabel polysilicon 586 -237 586 -237 0 4
rlabel polysilicon 639 -231 639 -231 0 1
rlabel polysilicon 639 -237 639 -237 0 3
rlabel polysilicon 653 -237 653 -237 0 3
rlabel polysilicon 26 -294 26 -294 0 4
rlabel polysilicon 30 -288 30 -288 0 1
rlabel polysilicon 30 -294 30 -294 0 3
rlabel polysilicon 40 -288 40 -288 0 2
rlabel polysilicon 44 -288 44 -288 0 1
rlabel polysilicon 44 -294 44 -294 0 3
rlabel polysilicon 51 -288 51 -288 0 1
rlabel polysilicon 51 -294 51 -294 0 3
rlabel polysilicon 58 -288 58 -288 0 1
rlabel polysilicon 58 -294 58 -294 0 3
rlabel polysilicon 65 -294 65 -294 0 3
rlabel polysilicon 72 -288 72 -288 0 1
rlabel polysilicon 72 -294 72 -294 0 3
rlabel polysilicon 79 -288 79 -288 0 1
rlabel polysilicon 79 -294 79 -294 0 3
rlabel polysilicon 86 -288 86 -288 0 1
rlabel polysilicon 86 -294 86 -294 0 3
rlabel polysilicon 93 -288 93 -288 0 1
rlabel polysilicon 93 -294 93 -294 0 3
rlabel polysilicon 100 -288 100 -288 0 1
rlabel polysilicon 100 -294 100 -294 0 3
rlabel polysilicon 107 -288 107 -288 0 1
rlabel polysilicon 107 -294 107 -294 0 3
rlabel polysilicon 114 -288 114 -288 0 1
rlabel polysilicon 114 -294 114 -294 0 3
rlabel polysilicon 124 -288 124 -288 0 2
rlabel polysilicon 128 -288 128 -288 0 1
rlabel polysilicon 128 -294 128 -294 0 3
rlabel polysilicon 135 -288 135 -288 0 1
rlabel polysilicon 135 -294 135 -294 0 3
rlabel polysilicon 145 -288 145 -288 0 2
rlabel polysilicon 142 -294 142 -294 0 3
rlabel polysilicon 152 -288 152 -288 0 2
rlabel polysilicon 149 -294 149 -294 0 3
rlabel polysilicon 156 -288 156 -288 0 1
rlabel polysilicon 156 -294 156 -294 0 3
rlabel polysilicon 163 -288 163 -288 0 1
rlabel polysilicon 163 -294 163 -294 0 3
rlabel polysilicon 166 -294 166 -294 0 4
rlabel polysilicon 170 -288 170 -288 0 1
rlabel polysilicon 170 -294 170 -294 0 3
rlabel polysilicon 180 -288 180 -288 0 2
rlabel polysilicon 177 -294 177 -294 0 3
rlabel polysilicon 184 -288 184 -288 0 1
rlabel polysilicon 184 -294 184 -294 0 3
rlabel polysilicon 194 -288 194 -288 0 2
rlabel polysilicon 191 -294 191 -294 0 3
rlabel polysilicon 198 -288 198 -288 0 1
rlabel polysilicon 198 -294 198 -294 0 3
rlabel polysilicon 205 -288 205 -288 0 1
rlabel polysilicon 205 -294 205 -294 0 3
rlabel polysilicon 212 -288 212 -288 0 1
rlabel polysilicon 215 -288 215 -288 0 2
rlabel polysilicon 215 -294 215 -294 0 4
rlabel polysilicon 219 -288 219 -288 0 1
rlabel polysilicon 219 -294 219 -294 0 3
rlabel polysilicon 222 -294 222 -294 0 4
rlabel polysilicon 226 -288 226 -288 0 1
rlabel polysilicon 226 -294 226 -294 0 3
rlabel polysilicon 233 -288 233 -288 0 1
rlabel polysilicon 233 -294 233 -294 0 3
rlabel polysilicon 240 -288 240 -288 0 1
rlabel polysilicon 240 -294 240 -294 0 3
rlabel polysilicon 247 -288 247 -288 0 1
rlabel polysilicon 247 -294 247 -294 0 3
rlabel polysilicon 250 -294 250 -294 0 4
rlabel polysilicon 254 -288 254 -288 0 1
rlabel polysilicon 254 -294 254 -294 0 3
rlabel polysilicon 257 -294 257 -294 0 4
rlabel polysilicon 261 -288 261 -288 0 1
rlabel polysilicon 261 -294 261 -294 0 3
rlabel polysilicon 268 -288 268 -288 0 1
rlabel polysilicon 268 -294 268 -294 0 3
rlabel polysilicon 275 -288 275 -288 0 1
rlabel polysilicon 278 -288 278 -288 0 2
rlabel polysilicon 278 -294 278 -294 0 4
rlabel polysilicon 285 -288 285 -288 0 2
rlabel polysilicon 282 -294 282 -294 0 3
rlabel polysilicon 289 -288 289 -288 0 1
rlabel polysilicon 289 -294 289 -294 0 3
rlabel polysilicon 296 -288 296 -288 0 1
rlabel polysilicon 299 -288 299 -288 0 2
rlabel polysilicon 299 -294 299 -294 0 4
rlabel polysilicon 303 -288 303 -288 0 1
rlabel polysilicon 303 -294 303 -294 0 3
rlabel polysilicon 310 -288 310 -288 0 1
rlabel polysilicon 313 -288 313 -288 0 2
rlabel polysilicon 310 -294 310 -294 0 3
rlabel polysilicon 313 -294 313 -294 0 4
rlabel polysilicon 317 -294 317 -294 0 3
rlabel polysilicon 320 -294 320 -294 0 4
rlabel polysilicon 324 -288 324 -288 0 1
rlabel polysilicon 324 -294 324 -294 0 3
rlabel polysilicon 331 -288 331 -288 0 1
rlabel polysilicon 331 -294 331 -294 0 3
rlabel polysilicon 338 -288 338 -288 0 1
rlabel polysilicon 338 -294 338 -294 0 3
rlabel polysilicon 341 -294 341 -294 0 4
rlabel polysilicon 345 -288 345 -288 0 1
rlabel polysilicon 345 -294 345 -294 0 3
rlabel polysilicon 352 -288 352 -288 0 1
rlabel polysilicon 352 -294 352 -294 0 3
rlabel polysilicon 359 -288 359 -288 0 1
rlabel polysilicon 359 -294 359 -294 0 3
rlabel polysilicon 362 -294 362 -294 0 4
rlabel polysilicon 366 -288 366 -288 0 1
rlabel polysilicon 366 -294 366 -294 0 3
rlabel polysilicon 373 -288 373 -288 0 1
rlabel polysilicon 373 -294 373 -294 0 3
rlabel polysilicon 380 -288 380 -288 0 1
rlabel polysilicon 380 -294 380 -294 0 3
rlabel polysilicon 387 -288 387 -288 0 1
rlabel polysilicon 387 -294 387 -294 0 3
rlabel polysilicon 394 -288 394 -288 0 1
rlabel polysilicon 394 -294 394 -294 0 3
rlabel polysilicon 401 -288 401 -288 0 1
rlabel polysilicon 401 -294 401 -294 0 3
rlabel polysilicon 408 -288 408 -288 0 1
rlabel polysilicon 408 -294 408 -294 0 3
rlabel polysilicon 415 -288 415 -288 0 1
rlabel polysilicon 415 -294 415 -294 0 3
rlabel polysilicon 422 -288 422 -288 0 1
rlabel polysilicon 422 -294 422 -294 0 3
rlabel polysilicon 429 -288 429 -288 0 1
rlabel polysilicon 429 -294 429 -294 0 3
rlabel polysilicon 439 -288 439 -288 0 2
rlabel polysilicon 436 -294 436 -294 0 3
rlabel polysilicon 443 -288 443 -288 0 1
rlabel polysilicon 443 -294 443 -294 0 3
rlabel polysilicon 450 -288 450 -288 0 1
rlabel polysilicon 450 -294 450 -294 0 3
rlabel polysilicon 457 -288 457 -288 0 1
rlabel polysilicon 457 -294 457 -294 0 3
rlabel polysilicon 464 -288 464 -288 0 1
rlabel polysilicon 464 -294 464 -294 0 3
rlabel polysilicon 471 -288 471 -288 0 1
rlabel polysilicon 471 -294 471 -294 0 3
rlabel polysilicon 481 -288 481 -288 0 2
rlabel polysilicon 485 -288 485 -288 0 1
rlabel polysilicon 485 -294 485 -294 0 3
rlabel polysilicon 492 -288 492 -288 0 1
rlabel polysilicon 492 -294 492 -294 0 3
rlabel polysilicon 499 -288 499 -288 0 1
rlabel polysilicon 499 -294 499 -294 0 3
rlabel polysilicon 506 -288 506 -288 0 1
rlabel polysilicon 506 -294 506 -294 0 3
rlabel polysilicon 513 -288 513 -288 0 1
rlabel polysilicon 513 -294 513 -294 0 3
rlabel polysilicon 520 -288 520 -288 0 1
rlabel polysilicon 520 -294 520 -294 0 3
rlabel polysilicon 527 -288 527 -288 0 1
rlabel polysilicon 527 -294 527 -294 0 3
rlabel polysilicon 534 -288 534 -288 0 1
rlabel polysilicon 534 -294 534 -294 0 3
rlabel polysilicon 541 -288 541 -288 0 1
rlabel polysilicon 541 -294 541 -294 0 3
rlabel polysilicon 548 -288 548 -288 0 1
rlabel polysilicon 548 -294 548 -294 0 3
rlabel polysilicon 555 -288 555 -288 0 1
rlabel polysilicon 555 -294 555 -294 0 3
rlabel polysilicon 562 -288 562 -288 0 1
rlabel polysilicon 562 -294 562 -294 0 3
rlabel polysilicon 569 -288 569 -288 0 1
rlabel polysilicon 569 -294 569 -294 0 3
rlabel polysilicon 576 -288 576 -288 0 1
rlabel polysilicon 576 -294 576 -294 0 3
rlabel polysilicon 583 -288 583 -288 0 1
rlabel polysilicon 583 -294 583 -294 0 3
rlabel polysilicon 590 -288 590 -288 0 1
rlabel polysilicon 590 -294 590 -294 0 3
rlabel polysilicon 597 -288 597 -288 0 1
rlabel polysilicon 597 -294 597 -294 0 3
rlabel polysilicon 604 -288 604 -288 0 1
rlabel polysilicon 604 -294 604 -294 0 3
rlabel polysilicon 611 -288 611 -288 0 1
rlabel polysilicon 611 -294 611 -294 0 3
rlabel polysilicon 618 -288 618 -288 0 1
rlabel polysilicon 618 -294 618 -294 0 3
rlabel polysilicon 625 -288 625 -288 0 1
rlabel polysilicon 625 -294 625 -294 0 3
rlabel polysilicon 632 -288 632 -288 0 1
rlabel polysilicon 632 -294 632 -294 0 3
rlabel polysilicon 653 -288 653 -288 0 1
rlabel polysilicon 653 -294 653 -294 0 3
rlabel polysilicon 660 -288 660 -288 0 1
rlabel polysilicon 660 -294 660 -294 0 3
rlabel polysilicon 9 -357 9 -357 0 1
rlabel polysilicon 9 -363 9 -363 0 3
rlabel polysilicon 23 -357 23 -357 0 1
rlabel polysilicon 23 -363 23 -363 0 3
rlabel polysilicon 30 -357 30 -357 0 1
rlabel polysilicon 30 -363 30 -363 0 3
rlabel polysilicon 58 -357 58 -357 0 1
rlabel polysilicon 58 -363 58 -363 0 3
rlabel polysilicon 72 -357 72 -357 0 1
rlabel polysilicon 72 -363 72 -363 0 3
rlabel polysilicon 79 -357 79 -357 0 1
rlabel polysilicon 79 -363 79 -363 0 3
rlabel polysilicon 86 -357 86 -357 0 1
rlabel polysilicon 86 -363 86 -363 0 3
rlabel polysilicon 93 -357 93 -357 0 1
rlabel polysilicon 93 -363 93 -363 0 3
rlabel polysilicon 100 -357 100 -357 0 1
rlabel polysilicon 107 -357 107 -357 0 1
rlabel polysilicon 110 -357 110 -357 0 2
rlabel polysilicon 107 -363 107 -363 0 3
rlabel polysilicon 114 -357 114 -357 0 1
rlabel polysilicon 117 -363 117 -363 0 4
rlabel polysilicon 121 -357 121 -357 0 1
rlabel polysilicon 121 -363 121 -363 0 3
rlabel polysilicon 128 -357 128 -357 0 1
rlabel polysilicon 128 -363 128 -363 0 3
rlabel polysilicon 135 -357 135 -357 0 1
rlabel polysilicon 135 -363 135 -363 0 3
rlabel polysilicon 142 -357 142 -357 0 1
rlabel polysilicon 142 -363 142 -363 0 3
rlabel polysilicon 152 -357 152 -357 0 2
rlabel polysilicon 149 -363 149 -363 0 3
rlabel polysilicon 152 -363 152 -363 0 4
rlabel polysilicon 159 -363 159 -363 0 4
rlabel polysilicon 163 -357 163 -357 0 1
rlabel polysilicon 163 -363 163 -363 0 3
rlabel polysilicon 170 -357 170 -357 0 1
rlabel polysilicon 170 -363 170 -363 0 3
rlabel polysilicon 177 -357 177 -357 0 1
rlabel polysilicon 177 -363 177 -363 0 3
rlabel polysilicon 180 -363 180 -363 0 4
rlabel polysilicon 184 -357 184 -357 0 1
rlabel polysilicon 187 -357 187 -357 0 2
rlabel polysilicon 191 -357 191 -357 0 1
rlabel polysilicon 191 -363 191 -363 0 3
rlabel polysilicon 194 -363 194 -363 0 4
rlabel polysilicon 198 -357 198 -357 0 1
rlabel polysilicon 198 -363 198 -363 0 3
rlabel polysilicon 208 -363 208 -363 0 4
rlabel polysilicon 212 -357 212 -357 0 1
rlabel polysilicon 212 -363 212 -363 0 3
rlabel polysilicon 219 -357 219 -357 0 1
rlabel polysilicon 222 -357 222 -357 0 2
rlabel polysilicon 219 -363 219 -363 0 3
rlabel polysilicon 222 -363 222 -363 0 4
rlabel polysilicon 226 -357 226 -357 0 1
rlabel polysilicon 226 -363 226 -363 0 3
rlabel polysilicon 233 -357 233 -357 0 1
rlabel polysilicon 233 -363 233 -363 0 3
rlabel polysilicon 240 -357 240 -357 0 1
rlabel polysilicon 240 -363 240 -363 0 3
rlabel polysilicon 247 -357 247 -357 0 1
rlabel polysilicon 247 -363 247 -363 0 3
rlabel polysilicon 254 -357 254 -357 0 1
rlabel polysilicon 254 -363 254 -363 0 3
rlabel polysilicon 261 -357 261 -357 0 1
rlabel polysilicon 261 -363 261 -363 0 3
rlabel polysilicon 268 -357 268 -357 0 1
rlabel polysilicon 268 -363 268 -363 0 3
rlabel polysilicon 275 -357 275 -357 0 1
rlabel polysilicon 278 -357 278 -357 0 2
rlabel polysilicon 275 -363 275 -363 0 3
rlabel polysilicon 282 -363 282 -363 0 3
rlabel polysilicon 289 -357 289 -357 0 1
rlabel polysilicon 289 -363 289 -363 0 3
rlabel polysilicon 296 -357 296 -357 0 1
rlabel polysilicon 299 -357 299 -357 0 2
rlabel polysilicon 296 -363 296 -363 0 3
rlabel polysilicon 303 -357 303 -357 0 1
rlabel polysilicon 303 -363 303 -363 0 3
rlabel polysilicon 310 -357 310 -357 0 1
rlabel polysilicon 310 -363 310 -363 0 3
rlabel polysilicon 317 -357 317 -357 0 1
rlabel polysilicon 317 -363 317 -363 0 3
rlabel polysilicon 324 -363 324 -363 0 3
rlabel polysilicon 327 -363 327 -363 0 4
rlabel polysilicon 331 -357 331 -357 0 1
rlabel polysilicon 331 -363 331 -363 0 3
rlabel polysilicon 338 -357 338 -357 0 1
rlabel polysilicon 338 -363 338 -363 0 3
rlabel polysilicon 345 -357 345 -357 0 1
rlabel polysilicon 345 -363 345 -363 0 3
rlabel polysilicon 352 -357 352 -357 0 1
rlabel polysilicon 352 -363 352 -363 0 3
rlabel polysilicon 355 -363 355 -363 0 4
rlabel polysilicon 362 -357 362 -357 0 2
rlabel polysilicon 362 -363 362 -363 0 4
rlabel polysilicon 366 -363 366 -363 0 3
rlabel polysilicon 373 -357 373 -357 0 1
rlabel polysilicon 373 -363 373 -363 0 3
rlabel polysilicon 383 -357 383 -357 0 2
rlabel polysilicon 383 -363 383 -363 0 4
rlabel polysilicon 390 -357 390 -357 0 2
rlabel polysilicon 387 -363 387 -363 0 3
rlabel polysilicon 390 -363 390 -363 0 4
rlabel polysilicon 394 -357 394 -357 0 1
rlabel polysilicon 394 -363 394 -363 0 3
rlabel polysilicon 401 -357 401 -357 0 1
rlabel polysilicon 401 -363 401 -363 0 3
rlabel polysilicon 408 -357 408 -357 0 1
rlabel polysilicon 408 -363 408 -363 0 3
rlabel polysilicon 415 -357 415 -357 0 1
rlabel polysilicon 415 -363 415 -363 0 3
rlabel polysilicon 422 -357 422 -357 0 1
rlabel polysilicon 422 -363 422 -363 0 3
rlabel polysilicon 429 -357 429 -357 0 1
rlabel polysilicon 432 -357 432 -357 0 2
rlabel polysilicon 429 -363 429 -363 0 3
rlabel polysilicon 436 -357 436 -357 0 1
rlabel polysilicon 436 -363 436 -363 0 3
rlabel polysilicon 443 -357 443 -357 0 1
rlabel polysilicon 443 -363 443 -363 0 3
rlabel polysilicon 453 -357 453 -357 0 2
rlabel polysilicon 453 -363 453 -363 0 4
rlabel polysilicon 457 -357 457 -357 0 1
rlabel polysilicon 457 -363 457 -363 0 3
rlabel polysilicon 464 -357 464 -357 0 1
rlabel polysilicon 464 -363 464 -363 0 3
rlabel polysilicon 471 -357 471 -357 0 1
rlabel polysilicon 471 -363 471 -363 0 3
rlabel polysilicon 478 -357 478 -357 0 1
rlabel polysilicon 478 -363 478 -363 0 3
rlabel polysilicon 485 -357 485 -357 0 1
rlabel polysilicon 485 -363 485 -363 0 3
rlabel polysilicon 492 -357 492 -357 0 1
rlabel polysilicon 492 -363 492 -363 0 3
rlabel polysilicon 506 -357 506 -357 0 1
rlabel polysilicon 506 -363 506 -363 0 3
rlabel polysilicon 513 -357 513 -357 0 1
rlabel polysilicon 513 -363 513 -363 0 3
rlabel polysilicon 520 -357 520 -357 0 1
rlabel polysilicon 520 -363 520 -363 0 3
rlabel polysilicon 527 -357 527 -357 0 1
rlabel polysilicon 527 -363 527 -363 0 3
rlabel polysilicon 534 -357 534 -357 0 1
rlabel polysilicon 534 -363 534 -363 0 3
rlabel polysilicon 541 -357 541 -357 0 1
rlabel polysilicon 541 -363 541 -363 0 3
rlabel polysilicon 548 -357 548 -357 0 1
rlabel polysilicon 548 -363 548 -363 0 3
rlabel polysilicon 555 -357 555 -357 0 1
rlabel polysilicon 555 -363 555 -363 0 3
rlabel polysilicon 562 -357 562 -357 0 1
rlabel polysilicon 562 -363 562 -363 0 3
rlabel polysilicon 569 -357 569 -357 0 1
rlabel polysilicon 569 -363 569 -363 0 3
rlabel polysilicon 576 -357 576 -357 0 1
rlabel polysilicon 576 -363 576 -363 0 3
rlabel polysilicon 583 -357 583 -357 0 1
rlabel polysilicon 583 -363 583 -363 0 3
rlabel polysilicon 590 -357 590 -357 0 1
rlabel polysilicon 590 -363 590 -363 0 3
rlabel polysilicon 597 -357 597 -357 0 1
rlabel polysilicon 597 -363 597 -363 0 3
rlabel polysilicon 604 -357 604 -357 0 1
rlabel polysilicon 604 -363 604 -363 0 3
rlabel polysilicon 611 -357 611 -357 0 1
rlabel polysilicon 611 -363 611 -363 0 3
rlabel polysilicon 621 -357 621 -357 0 2
rlabel polysilicon 653 -357 653 -357 0 1
rlabel polysilicon 656 -357 656 -357 0 2
rlabel polysilicon 653 -363 653 -363 0 3
rlabel polysilicon 660 -357 660 -357 0 1
rlabel polysilicon 660 -363 660 -363 0 3
rlabel polysilicon 670 -363 670 -363 0 4
rlabel polysilicon 674 -357 674 -357 0 1
rlabel polysilicon 674 -363 674 -363 0 3
rlabel polysilicon 16 -424 16 -424 0 1
rlabel polysilicon 16 -430 16 -430 0 3
rlabel polysilicon 33 -424 33 -424 0 2
rlabel polysilicon 40 -430 40 -430 0 4
rlabel polysilicon 44 -424 44 -424 0 1
rlabel polysilicon 44 -430 44 -430 0 3
rlabel polysilicon 51 -424 51 -424 0 1
rlabel polysilicon 51 -430 51 -430 0 3
rlabel polysilicon 61 -430 61 -430 0 4
rlabel polysilicon 65 -424 65 -424 0 1
rlabel polysilicon 65 -430 65 -430 0 3
rlabel polysilicon 72 -424 72 -424 0 1
rlabel polysilicon 72 -430 72 -430 0 3
rlabel polysilicon 82 -430 82 -430 0 4
rlabel polysilicon 86 -424 86 -424 0 1
rlabel polysilicon 86 -430 86 -430 0 3
rlabel polysilicon 93 -424 93 -424 0 1
rlabel polysilicon 93 -430 93 -430 0 3
rlabel polysilicon 100 -424 100 -424 0 1
rlabel polysilicon 100 -430 100 -430 0 3
rlabel polysilicon 107 -424 107 -424 0 1
rlabel polysilicon 107 -430 107 -430 0 3
rlabel polysilicon 114 -424 114 -424 0 1
rlabel polysilicon 117 -424 117 -424 0 2
rlabel polysilicon 114 -430 114 -430 0 3
rlabel polysilicon 117 -430 117 -430 0 4
rlabel polysilicon 121 -424 121 -424 0 1
rlabel polysilicon 121 -430 121 -430 0 3
rlabel polysilicon 128 -424 128 -424 0 1
rlabel polysilicon 128 -430 128 -430 0 3
rlabel polysilicon 135 -424 135 -424 0 1
rlabel polysilicon 138 -424 138 -424 0 2
rlabel polysilicon 142 -424 142 -424 0 1
rlabel polysilicon 142 -430 142 -430 0 3
rlabel polysilicon 149 -424 149 -424 0 1
rlabel polysilicon 149 -430 149 -430 0 3
rlabel polysilicon 156 -424 156 -424 0 1
rlabel polysilicon 156 -430 156 -430 0 3
rlabel polysilicon 163 -424 163 -424 0 1
rlabel polysilicon 166 -424 166 -424 0 2
rlabel polysilicon 166 -430 166 -430 0 4
rlabel polysilicon 170 -424 170 -424 0 1
rlabel polysilicon 173 -430 173 -430 0 4
rlabel polysilicon 177 -424 177 -424 0 1
rlabel polysilicon 177 -430 177 -430 0 3
rlabel polysilicon 184 -424 184 -424 0 1
rlabel polysilicon 184 -430 184 -430 0 3
rlabel polysilicon 191 -424 191 -424 0 1
rlabel polysilicon 194 -430 194 -430 0 4
rlabel polysilicon 198 -424 198 -424 0 1
rlabel polysilicon 198 -430 198 -430 0 3
rlabel polysilicon 201 -430 201 -430 0 4
rlabel polysilicon 205 -430 205 -430 0 3
rlabel polysilicon 215 -424 215 -424 0 2
rlabel polysilicon 215 -430 215 -430 0 4
rlabel polysilicon 222 -424 222 -424 0 2
rlabel polysilicon 222 -430 222 -430 0 4
rlabel polysilicon 226 -424 226 -424 0 1
rlabel polysilicon 229 -424 229 -424 0 2
rlabel polysilicon 226 -430 226 -430 0 3
rlabel polysilicon 229 -430 229 -430 0 4
rlabel polysilicon 233 -424 233 -424 0 1
rlabel polysilicon 233 -430 233 -430 0 3
rlabel polysilicon 240 -424 240 -424 0 1
rlabel polysilicon 240 -430 240 -430 0 3
rlabel polysilicon 247 -424 247 -424 0 1
rlabel polysilicon 250 -424 250 -424 0 2
rlabel polysilicon 247 -430 247 -430 0 3
rlabel polysilicon 254 -424 254 -424 0 1
rlabel polysilicon 257 -430 257 -430 0 4
rlabel polysilicon 261 -424 261 -424 0 1
rlabel polysilicon 264 -424 264 -424 0 2
rlabel polysilicon 261 -430 261 -430 0 3
rlabel polysilicon 264 -430 264 -430 0 4
rlabel polysilicon 268 -424 268 -424 0 1
rlabel polysilicon 268 -430 268 -430 0 3
rlabel polysilicon 275 -424 275 -424 0 1
rlabel polysilicon 275 -430 275 -430 0 3
rlabel polysilicon 282 -424 282 -424 0 1
rlabel polysilicon 285 -424 285 -424 0 2
rlabel polysilicon 282 -430 282 -430 0 3
rlabel polysilicon 289 -424 289 -424 0 1
rlabel polysilicon 296 -424 296 -424 0 1
rlabel polysilicon 296 -430 296 -430 0 3
rlabel polysilicon 303 -424 303 -424 0 1
rlabel polysilicon 303 -430 303 -430 0 3
rlabel polysilicon 310 -430 310 -430 0 3
rlabel polysilicon 317 -424 317 -424 0 1
rlabel polysilicon 317 -430 317 -430 0 3
rlabel polysilicon 320 -430 320 -430 0 4
rlabel polysilicon 324 -424 324 -424 0 1
rlabel polysilicon 327 -430 327 -430 0 4
rlabel polysilicon 331 -424 331 -424 0 1
rlabel polysilicon 331 -430 331 -430 0 3
rlabel polysilicon 341 -424 341 -424 0 2
rlabel polysilicon 338 -430 338 -430 0 3
rlabel polysilicon 345 -424 345 -424 0 1
rlabel polysilicon 345 -430 345 -430 0 3
rlabel polysilicon 352 -424 352 -424 0 1
rlabel polysilicon 352 -430 352 -430 0 3
rlabel polysilicon 359 -424 359 -424 0 1
rlabel polysilicon 362 -424 362 -424 0 2
rlabel polysilicon 359 -430 359 -430 0 3
rlabel polysilicon 362 -430 362 -430 0 4
rlabel polysilicon 366 -424 366 -424 0 1
rlabel polysilicon 366 -430 366 -430 0 3
rlabel polysilicon 373 -424 373 -424 0 1
rlabel polysilicon 373 -430 373 -430 0 3
rlabel polysilicon 383 -424 383 -424 0 2
rlabel polysilicon 380 -430 380 -430 0 3
rlabel polysilicon 383 -430 383 -430 0 4
rlabel polysilicon 387 -424 387 -424 0 1
rlabel polysilicon 387 -430 387 -430 0 3
rlabel polysilicon 390 -430 390 -430 0 4
rlabel polysilicon 394 -424 394 -424 0 1
rlabel polysilicon 394 -430 394 -430 0 3
rlabel polysilicon 401 -424 401 -424 0 1
rlabel polysilicon 401 -430 401 -430 0 3
rlabel polysilicon 408 -424 408 -424 0 1
rlabel polysilicon 408 -430 408 -430 0 3
rlabel polysilicon 415 -424 415 -424 0 1
rlabel polysilicon 415 -430 415 -430 0 3
rlabel polysilicon 422 -424 422 -424 0 1
rlabel polysilicon 422 -430 422 -430 0 3
rlabel polysilicon 429 -424 429 -424 0 1
rlabel polysilicon 429 -430 429 -430 0 3
rlabel polysilicon 436 -424 436 -424 0 1
rlabel polysilicon 436 -430 436 -430 0 3
rlabel polysilicon 443 -424 443 -424 0 1
rlabel polysilicon 443 -430 443 -430 0 3
rlabel polysilicon 450 -424 450 -424 0 1
rlabel polysilicon 450 -430 450 -430 0 3
rlabel polysilicon 457 -424 457 -424 0 1
rlabel polysilicon 457 -430 457 -430 0 3
rlabel polysilicon 464 -424 464 -424 0 1
rlabel polysilicon 464 -430 464 -430 0 3
rlabel polysilicon 474 -424 474 -424 0 2
rlabel polysilicon 471 -430 471 -430 0 3
rlabel polysilicon 481 -424 481 -424 0 2
rlabel polysilicon 478 -430 478 -430 0 3
rlabel polysilicon 485 -424 485 -424 0 1
rlabel polysilicon 485 -430 485 -430 0 3
rlabel polysilicon 492 -424 492 -424 0 1
rlabel polysilicon 492 -430 492 -430 0 3
rlabel polysilicon 499 -424 499 -424 0 1
rlabel polysilicon 499 -430 499 -430 0 3
rlabel polysilicon 506 -424 506 -424 0 1
rlabel polysilicon 506 -430 506 -430 0 3
rlabel polysilicon 513 -424 513 -424 0 1
rlabel polysilicon 513 -430 513 -430 0 3
rlabel polysilicon 520 -424 520 -424 0 1
rlabel polysilicon 520 -430 520 -430 0 3
rlabel polysilicon 527 -424 527 -424 0 1
rlabel polysilicon 527 -430 527 -430 0 3
rlabel polysilicon 534 -424 534 -424 0 1
rlabel polysilicon 534 -430 534 -430 0 3
rlabel polysilicon 541 -424 541 -424 0 1
rlabel polysilicon 541 -430 541 -430 0 3
rlabel polysilicon 544 -430 544 -430 0 4
rlabel polysilicon 548 -424 548 -424 0 1
rlabel polysilicon 548 -430 548 -430 0 3
rlabel polysilicon 555 -424 555 -424 0 1
rlabel polysilicon 555 -430 555 -430 0 3
rlabel polysilicon 562 -424 562 -424 0 1
rlabel polysilicon 562 -430 562 -430 0 3
rlabel polysilicon 569 -424 569 -424 0 1
rlabel polysilicon 569 -430 569 -430 0 3
rlabel polysilicon 576 -424 576 -424 0 1
rlabel polysilicon 576 -430 576 -430 0 3
rlabel polysilicon 583 -424 583 -424 0 1
rlabel polysilicon 583 -430 583 -430 0 3
rlabel polysilicon 590 -424 590 -424 0 1
rlabel polysilicon 590 -430 590 -430 0 3
rlabel polysilicon 597 -424 597 -424 0 1
rlabel polysilicon 597 -430 597 -430 0 3
rlabel polysilicon 604 -424 604 -424 0 1
rlabel polysilicon 604 -430 604 -430 0 3
rlabel polysilicon 611 -424 611 -424 0 1
rlabel polysilicon 611 -430 611 -430 0 3
rlabel polysilicon 618 -424 618 -424 0 1
rlabel polysilicon 618 -430 618 -430 0 3
rlabel polysilicon 625 -424 625 -424 0 1
rlabel polysilicon 625 -430 625 -430 0 3
rlabel polysilicon 632 -424 632 -424 0 1
rlabel polysilicon 632 -430 632 -430 0 3
rlabel polysilicon 639 -424 639 -424 0 1
rlabel polysilicon 639 -430 639 -430 0 3
rlabel polysilicon 646 -424 646 -424 0 1
rlabel polysilicon 646 -430 646 -430 0 3
rlabel polysilicon 653 -424 653 -424 0 1
rlabel polysilicon 653 -430 653 -430 0 3
rlabel polysilicon 660 -424 660 -424 0 1
rlabel polysilicon 660 -430 660 -430 0 3
rlabel polysilicon 667 -424 667 -424 0 1
rlabel polysilicon 667 -430 667 -430 0 3
rlabel polysilicon 674 -424 674 -424 0 1
rlabel polysilicon 681 -424 681 -424 0 1
rlabel polysilicon 681 -430 681 -430 0 3
rlabel polysilicon 26 -517 26 -517 0 4
rlabel polysilicon 33 -511 33 -511 0 2
rlabel polysilicon 30 -517 30 -517 0 3
rlabel polysilicon 37 -511 37 -511 0 1
rlabel polysilicon 44 -511 44 -511 0 1
rlabel polysilicon 44 -517 44 -517 0 3
rlabel polysilicon 51 -517 51 -517 0 3
rlabel polysilicon 58 -511 58 -511 0 1
rlabel polysilicon 58 -517 58 -517 0 3
rlabel polysilicon 65 -511 65 -511 0 1
rlabel polysilicon 65 -517 65 -517 0 3
rlabel polysilicon 72 -511 72 -511 0 1
rlabel polysilicon 72 -517 72 -517 0 3
rlabel polysilicon 79 -511 79 -511 0 1
rlabel polysilicon 79 -517 79 -517 0 3
rlabel polysilicon 86 -511 86 -511 0 1
rlabel polysilicon 93 -511 93 -511 0 1
rlabel polysilicon 93 -517 93 -517 0 3
rlabel polysilicon 100 -511 100 -511 0 1
rlabel polysilicon 100 -517 100 -517 0 3
rlabel polysilicon 110 -511 110 -511 0 2
rlabel polysilicon 107 -517 107 -517 0 3
rlabel polysilicon 114 -511 114 -511 0 1
rlabel polysilicon 114 -517 114 -517 0 3
rlabel polysilicon 121 -517 121 -517 0 3
rlabel polysilicon 124 -517 124 -517 0 4
rlabel polysilicon 128 -511 128 -511 0 1
rlabel polysilicon 128 -517 128 -517 0 3
rlabel polysilicon 135 -511 135 -511 0 1
rlabel polysilicon 135 -517 135 -517 0 3
rlabel polysilicon 142 -517 142 -517 0 3
rlabel polysilicon 145 -517 145 -517 0 4
rlabel polysilicon 149 -511 149 -511 0 1
rlabel polysilicon 149 -517 149 -517 0 3
rlabel polysilicon 156 -511 156 -511 0 1
rlabel polysilicon 156 -517 156 -517 0 3
rlabel polysilicon 163 -511 163 -511 0 1
rlabel polysilicon 163 -517 163 -517 0 3
rlabel polysilicon 173 -517 173 -517 0 4
rlabel polysilicon 177 -511 177 -511 0 1
rlabel polysilicon 177 -517 177 -517 0 3
rlabel polysilicon 184 -511 184 -511 0 1
rlabel polysilicon 184 -517 184 -517 0 3
rlabel polysilicon 191 -511 191 -511 0 1
rlabel polysilicon 191 -517 191 -517 0 3
rlabel polysilicon 198 -511 198 -511 0 1
rlabel polysilicon 201 -517 201 -517 0 4
rlabel polysilicon 205 -511 205 -511 0 1
rlabel polysilicon 205 -517 205 -517 0 3
rlabel polysilicon 212 -511 212 -511 0 1
rlabel polysilicon 215 -511 215 -511 0 2
rlabel polysilicon 215 -517 215 -517 0 4
rlabel polysilicon 219 -511 219 -511 0 1
rlabel polysilicon 219 -517 219 -517 0 3
rlabel polysilicon 226 -511 226 -511 0 1
rlabel polysilicon 229 -511 229 -511 0 2
rlabel polysilicon 233 -511 233 -511 0 1
rlabel polysilicon 233 -517 233 -517 0 3
rlabel polysilicon 240 -511 240 -511 0 1
rlabel polysilicon 243 -511 243 -511 0 2
rlabel polysilicon 240 -517 240 -517 0 3
rlabel polysilicon 243 -517 243 -517 0 4
rlabel polysilicon 247 -511 247 -511 0 1
rlabel polysilicon 247 -517 247 -517 0 3
rlabel polysilicon 254 -511 254 -511 0 1
rlabel polysilicon 257 -511 257 -511 0 2
rlabel polysilicon 254 -517 254 -517 0 3
rlabel polysilicon 257 -517 257 -517 0 4
rlabel polysilicon 261 -511 261 -511 0 1
rlabel polysilicon 261 -517 261 -517 0 3
rlabel polysilicon 268 -511 268 -511 0 1
rlabel polysilicon 271 -511 271 -511 0 2
rlabel polysilicon 275 -511 275 -511 0 1
rlabel polysilicon 275 -517 275 -517 0 3
rlabel polysilicon 282 -511 282 -511 0 1
rlabel polysilicon 282 -517 282 -517 0 3
rlabel polysilicon 285 -517 285 -517 0 4
rlabel polysilicon 289 -517 289 -517 0 3
rlabel polysilicon 296 -517 296 -517 0 3
rlabel polysilicon 299 -517 299 -517 0 4
rlabel polysilicon 303 -511 303 -511 0 1
rlabel polysilicon 303 -517 303 -517 0 3
rlabel polysilicon 310 -511 310 -511 0 1
rlabel polysilicon 310 -517 310 -517 0 3
rlabel polysilicon 317 -511 317 -511 0 1
rlabel polysilicon 320 -511 320 -511 0 2
rlabel polysilicon 317 -517 317 -517 0 3
rlabel polysilicon 320 -517 320 -517 0 4
rlabel polysilicon 327 -511 327 -511 0 2
rlabel polysilicon 324 -517 324 -517 0 3
rlabel polysilicon 327 -517 327 -517 0 4
rlabel polysilicon 331 -511 331 -511 0 1
rlabel polysilicon 331 -517 331 -517 0 3
rlabel polysilicon 338 -511 338 -511 0 1
rlabel polysilicon 338 -517 338 -517 0 3
rlabel polysilicon 348 -511 348 -511 0 2
rlabel polysilicon 348 -517 348 -517 0 4
rlabel polysilicon 352 -511 352 -511 0 1
rlabel polysilicon 355 -511 355 -511 0 2
rlabel polysilicon 355 -517 355 -517 0 4
rlabel polysilicon 359 -511 359 -511 0 1
rlabel polysilicon 362 -517 362 -517 0 4
rlabel polysilicon 366 -511 366 -511 0 1
rlabel polysilicon 366 -517 366 -517 0 3
rlabel polysilicon 373 -511 373 -511 0 1
rlabel polysilicon 373 -517 373 -517 0 3
rlabel polysilicon 380 -511 380 -511 0 1
rlabel polysilicon 380 -517 380 -517 0 3
rlabel polysilicon 390 -511 390 -511 0 2
rlabel polysilicon 387 -517 387 -517 0 3
rlabel polysilicon 390 -517 390 -517 0 4
rlabel polysilicon 394 -511 394 -511 0 1
rlabel polysilicon 394 -517 394 -517 0 3
rlabel polysilicon 401 -517 401 -517 0 3
rlabel polysilicon 404 -517 404 -517 0 4
rlabel polysilicon 408 -511 408 -511 0 1
rlabel polysilicon 408 -517 408 -517 0 3
rlabel polysilicon 415 -511 415 -511 0 1
rlabel polysilicon 415 -517 415 -517 0 3
rlabel polysilicon 422 -511 422 -511 0 1
rlabel polysilicon 425 -511 425 -511 0 2
rlabel polysilicon 425 -517 425 -517 0 4
rlabel polysilicon 429 -511 429 -511 0 1
rlabel polysilicon 429 -517 429 -517 0 3
rlabel polysilicon 439 -511 439 -511 0 2
rlabel polysilicon 439 -517 439 -517 0 4
rlabel polysilicon 443 -511 443 -511 0 1
rlabel polysilicon 443 -517 443 -517 0 3
rlabel polysilicon 450 -511 450 -511 0 1
rlabel polysilicon 450 -517 450 -517 0 3
rlabel polysilicon 457 -511 457 -511 0 1
rlabel polysilicon 457 -517 457 -517 0 3
rlabel polysilicon 464 -511 464 -511 0 1
rlabel polysilicon 464 -517 464 -517 0 3
rlabel polysilicon 471 -511 471 -511 0 1
rlabel polysilicon 471 -517 471 -517 0 3
rlabel polysilicon 478 -511 478 -511 0 1
rlabel polysilicon 478 -517 478 -517 0 3
rlabel polysilicon 485 -511 485 -511 0 1
rlabel polysilicon 485 -517 485 -517 0 3
rlabel polysilicon 492 -511 492 -511 0 1
rlabel polysilicon 492 -517 492 -517 0 3
rlabel polysilicon 499 -511 499 -511 0 1
rlabel polysilicon 499 -517 499 -517 0 3
rlabel polysilicon 506 -511 506 -511 0 1
rlabel polysilicon 506 -517 506 -517 0 3
rlabel polysilicon 513 -511 513 -511 0 1
rlabel polysilicon 513 -517 513 -517 0 3
rlabel polysilicon 520 -511 520 -511 0 1
rlabel polysilicon 520 -517 520 -517 0 3
rlabel polysilicon 527 -511 527 -511 0 1
rlabel polysilicon 527 -517 527 -517 0 3
rlabel polysilicon 534 -511 534 -511 0 1
rlabel polysilicon 534 -517 534 -517 0 3
rlabel polysilicon 541 -511 541 -511 0 1
rlabel polysilicon 544 -511 544 -511 0 2
rlabel polysilicon 541 -517 541 -517 0 3
rlabel polysilicon 548 -511 548 -511 0 1
rlabel polysilicon 548 -517 548 -517 0 3
rlabel polysilicon 555 -511 555 -511 0 1
rlabel polysilicon 555 -517 555 -517 0 3
rlabel polysilicon 562 -511 562 -511 0 1
rlabel polysilicon 562 -517 562 -517 0 3
rlabel polysilicon 569 -511 569 -511 0 1
rlabel polysilicon 569 -517 569 -517 0 3
rlabel polysilicon 576 -511 576 -511 0 1
rlabel polysilicon 576 -517 576 -517 0 3
rlabel polysilicon 583 -511 583 -511 0 1
rlabel polysilicon 583 -517 583 -517 0 3
rlabel polysilicon 590 -511 590 -511 0 1
rlabel polysilicon 590 -517 590 -517 0 3
rlabel polysilicon 597 -511 597 -511 0 1
rlabel polysilicon 597 -517 597 -517 0 3
rlabel polysilicon 604 -511 604 -511 0 1
rlabel polysilicon 604 -517 604 -517 0 3
rlabel polysilicon 611 -511 611 -511 0 1
rlabel polysilicon 611 -517 611 -517 0 3
rlabel polysilicon 618 -511 618 -511 0 1
rlabel polysilicon 618 -517 618 -517 0 3
rlabel polysilicon 625 -511 625 -511 0 1
rlabel polysilicon 625 -517 625 -517 0 3
rlabel polysilicon 632 -511 632 -511 0 1
rlabel polysilicon 632 -517 632 -517 0 3
rlabel polysilicon 639 -511 639 -511 0 1
rlabel polysilicon 639 -517 639 -517 0 3
rlabel polysilicon 646 -511 646 -511 0 1
rlabel polysilicon 646 -517 646 -517 0 3
rlabel polysilicon 653 -511 653 -511 0 1
rlabel polysilicon 653 -517 653 -517 0 3
rlabel polysilicon 660 -511 660 -511 0 1
rlabel polysilicon 660 -517 660 -517 0 3
rlabel polysilicon 667 -511 667 -511 0 1
rlabel polysilicon 667 -517 667 -517 0 3
rlabel polysilicon 674 -511 674 -511 0 1
rlabel polysilicon 674 -517 674 -517 0 3
rlabel polysilicon 681 -511 681 -511 0 1
rlabel polysilicon 681 -517 681 -517 0 3
rlabel polysilicon 688 -511 688 -511 0 1
rlabel polysilicon 688 -517 688 -517 0 3
rlabel polysilicon 695 -511 695 -511 0 1
rlabel polysilicon 695 -517 695 -517 0 3
rlabel polysilicon 702 -511 702 -511 0 1
rlabel polysilicon 702 -517 702 -517 0 3
rlabel polysilicon 709 -511 709 -511 0 1
rlabel polysilicon 709 -517 709 -517 0 3
rlabel polysilicon 16 -598 16 -598 0 1
rlabel polysilicon 23 -598 23 -598 0 1
rlabel polysilicon 23 -604 23 -604 0 3
rlabel polysilicon 30 -598 30 -598 0 1
rlabel polysilicon 30 -604 30 -604 0 3
rlabel polysilicon 37 -598 37 -598 0 1
rlabel polysilicon 37 -604 37 -604 0 3
rlabel polysilicon 44 -598 44 -598 0 1
rlabel polysilicon 44 -604 44 -604 0 3
rlabel polysilicon 54 -598 54 -598 0 2
rlabel polysilicon 54 -604 54 -604 0 4
rlabel polysilicon 58 -598 58 -598 0 1
rlabel polysilicon 58 -604 58 -604 0 3
rlabel polysilicon 65 -598 65 -598 0 1
rlabel polysilicon 68 -598 68 -598 0 2
rlabel polysilicon 65 -604 65 -604 0 3
rlabel polysilicon 72 -598 72 -598 0 1
rlabel polysilicon 79 -598 79 -598 0 1
rlabel polysilicon 79 -604 79 -604 0 3
rlabel polysilicon 86 -598 86 -598 0 1
rlabel polysilicon 86 -604 86 -604 0 3
rlabel polysilicon 93 -598 93 -598 0 1
rlabel polysilicon 93 -604 93 -604 0 3
rlabel polysilicon 100 -604 100 -604 0 3
rlabel polysilicon 103 -604 103 -604 0 4
rlabel polysilicon 107 -598 107 -598 0 1
rlabel polysilicon 107 -604 107 -604 0 3
rlabel polysilicon 114 -598 114 -598 0 1
rlabel polysilicon 117 -598 117 -598 0 2
rlabel polysilicon 117 -604 117 -604 0 4
rlabel polysilicon 121 -598 121 -598 0 1
rlabel polysilicon 121 -604 121 -604 0 3
rlabel polysilicon 131 -598 131 -598 0 2
rlabel polysilicon 128 -604 128 -604 0 3
rlabel polysilicon 135 -598 135 -598 0 1
rlabel polysilicon 135 -604 135 -604 0 3
rlabel polysilicon 142 -598 142 -598 0 1
rlabel polysilicon 142 -604 142 -604 0 3
rlabel polysilicon 149 -598 149 -598 0 1
rlabel polysilicon 149 -604 149 -604 0 3
rlabel polysilicon 159 -598 159 -598 0 2
rlabel polysilicon 163 -598 163 -598 0 1
rlabel polysilicon 163 -604 163 -604 0 3
rlabel polysilicon 170 -598 170 -598 0 1
rlabel polysilicon 170 -604 170 -604 0 3
rlabel polysilicon 177 -598 177 -598 0 1
rlabel polysilicon 177 -604 177 -604 0 3
rlabel polysilicon 184 -598 184 -598 0 1
rlabel polysilicon 184 -604 184 -604 0 3
rlabel polysilicon 194 -598 194 -598 0 2
rlabel polysilicon 194 -604 194 -604 0 4
rlabel polysilicon 198 -598 198 -598 0 1
rlabel polysilicon 201 -598 201 -598 0 2
rlabel polysilicon 198 -604 198 -604 0 3
rlabel polysilicon 201 -604 201 -604 0 4
rlabel polysilicon 205 -598 205 -598 0 1
rlabel polysilicon 205 -604 205 -604 0 3
rlabel polysilicon 212 -598 212 -598 0 1
rlabel polysilicon 215 -598 215 -598 0 2
rlabel polysilicon 215 -604 215 -604 0 4
rlabel polysilicon 219 -598 219 -598 0 1
rlabel polysilicon 222 -604 222 -604 0 4
rlabel polysilicon 226 -598 226 -598 0 1
rlabel polysilicon 226 -604 226 -604 0 3
rlabel polysilicon 233 -598 233 -598 0 1
rlabel polysilicon 233 -604 233 -604 0 3
rlabel polysilicon 240 -598 240 -598 0 1
rlabel polysilicon 240 -604 240 -604 0 3
rlabel polysilicon 247 -598 247 -598 0 1
rlabel polysilicon 247 -604 247 -604 0 3
rlabel polysilicon 254 -598 254 -598 0 1
rlabel polysilicon 254 -604 254 -604 0 3
rlabel polysilicon 261 -598 261 -598 0 1
rlabel polysilicon 261 -604 261 -604 0 3
rlabel polysilicon 268 -598 268 -598 0 1
rlabel polysilicon 268 -604 268 -604 0 3
rlabel polysilicon 275 -598 275 -598 0 1
rlabel polysilicon 285 -598 285 -598 0 2
rlabel polysilicon 285 -604 285 -604 0 4
rlabel polysilicon 289 -598 289 -598 0 1
rlabel polysilicon 289 -604 289 -604 0 3
rlabel polysilicon 296 -598 296 -598 0 1
rlabel polysilicon 296 -604 296 -604 0 3
rlabel polysilicon 306 -598 306 -598 0 2
rlabel polysilicon 303 -604 303 -604 0 3
rlabel polysilicon 310 -598 310 -598 0 1
rlabel polysilicon 310 -604 310 -604 0 3
rlabel polysilicon 317 -598 317 -598 0 1
rlabel polysilicon 320 -598 320 -598 0 2
rlabel polysilicon 317 -604 317 -604 0 3
rlabel polysilicon 320 -604 320 -604 0 4
rlabel polysilicon 324 -598 324 -598 0 1
rlabel polysilicon 324 -604 324 -604 0 3
rlabel polysilicon 331 -598 331 -598 0 1
rlabel polysilicon 331 -604 331 -604 0 3
rlabel polysilicon 338 -598 338 -598 0 1
rlabel polysilicon 345 -598 345 -598 0 1
rlabel polysilicon 348 -604 348 -604 0 4
rlabel polysilicon 352 -598 352 -598 0 1
rlabel polysilicon 352 -604 352 -604 0 3
rlabel polysilicon 359 -598 359 -598 0 1
rlabel polysilicon 359 -604 359 -604 0 3
rlabel polysilicon 366 -598 366 -598 0 1
rlabel polysilicon 366 -604 366 -604 0 3
rlabel polysilicon 373 -604 373 -604 0 3
rlabel polysilicon 376 -604 376 -604 0 4
rlabel polysilicon 380 -598 380 -598 0 1
rlabel polysilicon 380 -604 380 -604 0 3
rlabel polysilicon 387 -598 387 -598 0 1
rlabel polysilicon 387 -604 387 -604 0 3
rlabel polysilicon 394 -598 394 -598 0 1
rlabel polysilicon 394 -604 394 -604 0 3
rlabel polysilicon 401 -598 401 -598 0 1
rlabel polysilicon 401 -604 401 -604 0 3
rlabel polysilicon 408 -598 408 -598 0 1
rlabel polysilicon 411 -598 411 -598 0 2
rlabel polysilicon 408 -604 408 -604 0 3
rlabel polysilicon 411 -604 411 -604 0 4
rlabel polysilicon 418 -598 418 -598 0 2
rlabel polysilicon 418 -604 418 -604 0 4
rlabel polysilicon 422 -598 422 -598 0 1
rlabel polysilicon 422 -604 422 -604 0 3
rlabel polysilicon 429 -598 429 -598 0 1
rlabel polysilicon 429 -604 429 -604 0 3
rlabel polysilicon 436 -598 436 -598 0 1
rlabel polysilicon 439 -598 439 -598 0 2
rlabel polysilicon 439 -604 439 -604 0 4
rlabel polysilicon 443 -598 443 -598 0 1
rlabel polysilicon 446 -604 446 -604 0 4
rlabel polysilicon 450 -598 450 -598 0 1
rlabel polysilicon 450 -604 450 -604 0 3
rlabel polysilicon 457 -598 457 -598 0 1
rlabel polysilicon 460 -598 460 -598 0 2
rlabel polysilicon 457 -604 457 -604 0 3
rlabel polysilicon 464 -598 464 -598 0 1
rlabel polysilicon 464 -604 464 -604 0 3
rlabel polysilicon 471 -604 471 -604 0 3
rlabel polysilicon 478 -598 478 -598 0 1
rlabel polysilicon 478 -604 478 -604 0 3
rlabel polysilicon 485 -598 485 -598 0 1
rlabel polysilicon 485 -604 485 -604 0 3
rlabel polysilicon 492 -598 492 -598 0 1
rlabel polysilicon 495 -598 495 -598 0 2
rlabel polysilicon 492 -604 492 -604 0 3
rlabel polysilicon 502 -598 502 -598 0 2
rlabel polysilicon 499 -604 499 -604 0 3
rlabel polysilicon 506 -598 506 -598 0 1
rlabel polysilicon 506 -604 506 -604 0 3
rlabel polysilicon 513 -598 513 -598 0 1
rlabel polysilicon 513 -604 513 -604 0 3
rlabel polysilicon 520 -598 520 -598 0 1
rlabel polysilicon 520 -604 520 -604 0 3
rlabel polysilicon 527 -598 527 -598 0 1
rlabel polysilicon 527 -604 527 -604 0 3
rlabel polysilicon 534 -598 534 -598 0 1
rlabel polysilicon 534 -604 534 -604 0 3
rlabel polysilicon 541 -598 541 -598 0 1
rlabel polysilicon 541 -604 541 -604 0 3
rlabel polysilicon 548 -598 548 -598 0 1
rlabel polysilicon 548 -604 548 -604 0 3
rlabel polysilicon 558 -598 558 -598 0 2
rlabel polysilicon 555 -604 555 -604 0 3
rlabel polysilicon 562 -598 562 -598 0 1
rlabel polysilicon 562 -604 562 -604 0 3
rlabel polysilicon 569 -598 569 -598 0 1
rlabel polysilicon 569 -604 569 -604 0 3
rlabel polysilicon 576 -598 576 -598 0 1
rlabel polysilicon 576 -604 576 -604 0 3
rlabel polysilicon 583 -598 583 -598 0 1
rlabel polysilicon 583 -604 583 -604 0 3
rlabel polysilicon 590 -598 590 -598 0 1
rlabel polysilicon 590 -604 590 -604 0 3
rlabel polysilicon 597 -598 597 -598 0 1
rlabel polysilicon 597 -604 597 -604 0 3
rlabel polysilicon 604 -598 604 -598 0 1
rlabel polysilicon 604 -604 604 -604 0 3
rlabel polysilicon 611 -598 611 -598 0 1
rlabel polysilicon 611 -604 611 -604 0 3
rlabel polysilicon 618 -598 618 -598 0 1
rlabel polysilicon 618 -604 618 -604 0 3
rlabel polysilicon 625 -598 625 -598 0 1
rlabel polysilicon 625 -604 625 -604 0 3
rlabel polysilicon 632 -598 632 -598 0 1
rlabel polysilicon 632 -604 632 -604 0 3
rlabel polysilicon 639 -598 639 -598 0 1
rlabel polysilicon 639 -604 639 -604 0 3
rlabel polysilicon 646 -598 646 -598 0 1
rlabel polysilicon 646 -604 646 -604 0 3
rlabel polysilicon 653 -598 653 -598 0 1
rlabel polysilicon 653 -604 653 -604 0 3
rlabel polysilicon 660 -598 660 -598 0 1
rlabel polysilicon 660 -604 660 -604 0 3
rlabel polysilicon 667 -598 667 -598 0 1
rlabel polysilicon 667 -604 667 -604 0 3
rlabel polysilicon 674 -598 674 -598 0 1
rlabel polysilicon 674 -604 674 -604 0 3
rlabel polysilicon 681 -598 681 -598 0 1
rlabel polysilicon 681 -604 681 -604 0 3
rlabel polysilicon 709 -598 709 -598 0 1
rlabel polysilicon 709 -604 709 -604 0 3
rlabel polysilicon 19 -677 19 -677 0 2
rlabel polysilicon 23 -677 23 -677 0 1
rlabel polysilicon 30 -683 30 -683 0 3
rlabel polysilicon 37 -677 37 -677 0 1
rlabel polysilicon 37 -683 37 -683 0 3
rlabel polysilicon 44 -677 44 -677 0 1
rlabel polysilicon 44 -683 44 -683 0 3
rlabel polysilicon 51 -677 51 -677 0 1
rlabel polysilicon 51 -683 51 -683 0 3
rlabel polysilicon 58 -677 58 -677 0 1
rlabel polysilicon 61 -683 61 -683 0 4
rlabel polysilicon 65 -677 65 -677 0 1
rlabel polysilicon 65 -683 65 -683 0 3
rlabel polysilicon 72 -677 72 -677 0 1
rlabel polysilicon 75 -677 75 -677 0 2
rlabel polysilicon 72 -683 72 -683 0 3
rlabel polysilicon 79 -677 79 -677 0 1
rlabel polysilicon 79 -683 79 -683 0 3
rlabel polysilicon 86 -677 86 -677 0 1
rlabel polysilicon 86 -683 86 -683 0 3
rlabel polysilicon 93 -677 93 -677 0 1
rlabel polysilicon 93 -683 93 -683 0 3
rlabel polysilicon 100 -677 100 -677 0 1
rlabel polysilicon 100 -683 100 -683 0 3
rlabel polysilicon 107 -677 107 -677 0 1
rlabel polysilicon 107 -683 107 -683 0 3
rlabel polysilicon 114 -677 114 -677 0 1
rlabel polysilicon 114 -683 114 -683 0 3
rlabel polysilicon 124 -677 124 -677 0 2
rlabel polysilicon 121 -683 121 -683 0 3
rlabel polysilicon 124 -683 124 -683 0 4
rlabel polysilicon 128 -683 128 -683 0 3
rlabel polysilicon 135 -677 135 -677 0 1
rlabel polysilicon 135 -683 135 -683 0 3
rlabel polysilicon 142 -677 142 -677 0 1
rlabel polysilicon 142 -683 142 -683 0 3
rlabel polysilicon 145 -683 145 -683 0 4
rlabel polysilicon 149 -677 149 -677 0 1
rlabel polysilicon 149 -683 149 -683 0 3
rlabel polysilicon 159 -677 159 -677 0 2
rlabel polysilicon 156 -683 156 -683 0 3
rlabel polysilicon 159 -683 159 -683 0 4
rlabel polysilicon 163 -677 163 -677 0 1
rlabel polysilicon 163 -683 163 -683 0 3
rlabel polysilicon 170 -677 170 -677 0 1
rlabel polysilicon 170 -683 170 -683 0 3
rlabel polysilicon 177 -677 177 -677 0 1
rlabel polysilicon 177 -683 177 -683 0 3
rlabel polysilicon 187 -677 187 -677 0 2
rlabel polysilicon 184 -683 184 -683 0 3
rlabel polysilicon 187 -683 187 -683 0 4
rlabel polysilicon 191 -677 191 -677 0 1
rlabel polysilicon 191 -683 191 -683 0 3
rlabel polysilicon 198 -677 198 -677 0 1
rlabel polysilicon 201 -677 201 -677 0 2
rlabel polysilicon 201 -683 201 -683 0 4
rlabel polysilicon 205 -677 205 -677 0 1
rlabel polysilicon 205 -683 205 -683 0 3
rlabel polysilicon 212 -677 212 -677 0 1
rlabel polysilicon 212 -683 212 -683 0 3
rlabel polysilicon 219 -677 219 -677 0 1
rlabel polysilicon 222 -677 222 -677 0 2
rlabel polysilicon 222 -683 222 -683 0 4
rlabel polysilicon 226 -677 226 -677 0 1
rlabel polysilicon 226 -683 226 -683 0 3
rlabel polysilicon 233 -677 233 -677 0 1
rlabel polysilicon 233 -683 233 -683 0 3
rlabel polysilicon 240 -677 240 -677 0 1
rlabel polysilicon 240 -683 240 -683 0 3
rlabel polysilicon 247 -677 247 -677 0 1
rlabel polysilicon 247 -683 247 -683 0 3
rlabel polysilicon 254 -677 254 -677 0 1
rlabel polysilicon 254 -683 254 -683 0 3
rlabel polysilicon 261 -677 261 -677 0 1
rlabel polysilicon 261 -683 261 -683 0 3
rlabel polysilicon 268 -677 268 -677 0 1
rlabel polysilicon 268 -683 268 -683 0 3
rlabel polysilicon 275 -677 275 -677 0 1
rlabel polysilicon 275 -683 275 -683 0 3
rlabel polysilicon 278 -683 278 -683 0 4
rlabel polysilicon 282 -677 282 -677 0 1
rlabel polysilicon 285 -677 285 -677 0 2
rlabel polysilicon 282 -683 282 -683 0 3
rlabel polysilicon 289 -677 289 -677 0 1
rlabel polysilicon 289 -683 289 -683 0 3
rlabel polysilicon 296 -677 296 -677 0 1
rlabel polysilicon 296 -683 296 -683 0 3
rlabel polysilicon 303 -677 303 -677 0 1
rlabel polysilicon 303 -683 303 -683 0 3
rlabel polysilicon 310 -677 310 -677 0 1
rlabel polysilicon 310 -683 310 -683 0 3
rlabel polysilicon 317 -677 317 -677 0 1
rlabel polysilicon 320 -683 320 -683 0 4
rlabel polysilicon 324 -677 324 -677 0 1
rlabel polysilicon 327 -683 327 -683 0 4
rlabel polysilicon 331 -677 331 -677 0 1
rlabel polysilicon 331 -683 331 -683 0 3
rlabel polysilicon 338 -677 338 -677 0 1
rlabel polysilicon 338 -683 338 -683 0 3
rlabel polysilicon 345 -683 345 -683 0 3
rlabel polysilicon 348 -683 348 -683 0 4
rlabel polysilicon 355 -677 355 -677 0 2
rlabel polysilicon 355 -683 355 -683 0 4
rlabel polysilicon 359 -677 359 -677 0 1
rlabel polysilicon 359 -683 359 -683 0 3
rlabel polysilicon 366 -677 366 -677 0 1
rlabel polysilicon 366 -683 366 -683 0 3
rlabel polysilicon 373 -677 373 -677 0 1
rlabel polysilicon 373 -683 373 -683 0 3
rlabel polysilicon 380 -677 380 -677 0 1
rlabel polysilicon 380 -683 380 -683 0 3
rlabel polysilicon 387 -677 387 -677 0 1
rlabel polysilicon 387 -683 387 -683 0 3
rlabel polysilicon 394 -677 394 -677 0 1
rlabel polysilicon 394 -683 394 -683 0 3
rlabel polysilicon 397 -683 397 -683 0 4
rlabel polysilicon 401 -677 401 -677 0 1
rlabel polysilicon 404 -677 404 -677 0 2
rlabel polysilicon 401 -683 401 -683 0 3
rlabel polysilicon 404 -683 404 -683 0 4
rlabel polysilicon 408 -677 408 -677 0 1
rlabel polysilicon 408 -683 408 -683 0 3
rlabel polysilicon 415 -677 415 -677 0 1
rlabel polysilicon 415 -683 415 -683 0 3
rlabel polysilicon 422 -677 422 -677 0 1
rlabel polysilicon 425 -677 425 -677 0 2
rlabel polysilicon 429 -677 429 -677 0 1
rlabel polysilicon 429 -683 429 -683 0 3
rlabel polysilicon 439 -677 439 -677 0 2
rlabel polysilicon 436 -683 436 -683 0 3
rlabel polysilicon 439 -683 439 -683 0 4
rlabel polysilicon 443 -677 443 -677 0 1
rlabel polysilicon 443 -683 443 -683 0 3
rlabel polysilicon 453 -677 453 -677 0 2
rlabel polysilicon 453 -683 453 -683 0 4
rlabel polysilicon 457 -677 457 -677 0 1
rlabel polysilicon 460 -677 460 -677 0 2
rlabel polysilicon 457 -683 457 -683 0 3
rlabel polysilicon 464 -677 464 -677 0 1
rlabel polysilicon 467 -677 467 -677 0 2
rlabel polysilicon 467 -683 467 -683 0 4
rlabel polysilicon 478 -677 478 -677 0 1
rlabel polysilicon 481 -683 481 -683 0 4
rlabel polysilicon 485 -677 485 -677 0 1
rlabel polysilicon 485 -683 485 -683 0 3
rlabel polysilicon 495 -683 495 -683 0 4
rlabel polysilicon 499 -677 499 -677 0 1
rlabel polysilicon 499 -683 499 -683 0 3
rlabel polysilicon 506 -683 506 -683 0 3
rlabel polysilicon 509 -683 509 -683 0 4
rlabel polysilicon 513 -677 513 -677 0 1
rlabel polysilicon 513 -683 513 -683 0 3
rlabel polysilicon 520 -677 520 -677 0 1
rlabel polysilicon 520 -683 520 -683 0 3
rlabel polysilicon 527 -677 527 -677 0 1
rlabel polysilicon 527 -683 527 -683 0 3
rlabel polysilicon 534 -677 534 -677 0 1
rlabel polysilicon 534 -683 534 -683 0 3
rlabel polysilicon 541 -677 541 -677 0 1
rlabel polysilicon 541 -683 541 -683 0 3
rlabel polysilicon 548 -677 548 -677 0 1
rlabel polysilicon 548 -683 548 -683 0 3
rlabel polysilicon 555 -677 555 -677 0 1
rlabel polysilicon 555 -683 555 -683 0 3
rlabel polysilicon 562 -677 562 -677 0 1
rlabel polysilicon 562 -683 562 -683 0 3
rlabel polysilicon 569 -677 569 -677 0 1
rlabel polysilicon 569 -683 569 -683 0 3
rlabel polysilicon 576 -677 576 -677 0 1
rlabel polysilicon 576 -683 576 -683 0 3
rlabel polysilicon 583 -677 583 -677 0 1
rlabel polysilicon 586 -683 586 -683 0 4
rlabel polysilicon 590 -677 590 -677 0 1
rlabel polysilicon 590 -683 590 -683 0 3
rlabel polysilicon 597 -677 597 -677 0 1
rlabel polysilicon 597 -683 597 -683 0 3
rlabel polysilicon 604 -677 604 -677 0 1
rlabel polysilicon 604 -683 604 -683 0 3
rlabel polysilicon 611 -677 611 -677 0 1
rlabel polysilicon 611 -683 611 -683 0 3
rlabel polysilicon 618 -677 618 -677 0 1
rlabel polysilicon 618 -683 618 -683 0 3
rlabel polysilicon 625 -677 625 -677 0 1
rlabel polysilicon 625 -683 625 -683 0 3
rlabel polysilicon 632 -677 632 -677 0 1
rlabel polysilicon 632 -683 632 -683 0 3
rlabel polysilicon 639 -677 639 -677 0 1
rlabel polysilicon 639 -683 639 -683 0 3
rlabel polysilicon 646 -677 646 -677 0 1
rlabel polysilicon 646 -683 646 -683 0 3
rlabel polysilicon 653 -677 653 -677 0 1
rlabel polysilicon 653 -683 653 -683 0 3
rlabel polysilicon 660 -677 660 -677 0 1
rlabel polysilicon 660 -683 660 -683 0 3
rlabel polysilicon 667 -677 667 -677 0 1
rlabel polysilicon 667 -683 667 -683 0 3
rlabel polysilicon 674 -677 674 -677 0 1
rlabel polysilicon 674 -683 674 -683 0 3
rlabel polysilicon 681 -677 681 -677 0 1
rlabel polysilicon 681 -683 681 -683 0 3
rlabel polysilicon 688 -677 688 -677 0 1
rlabel polysilicon 688 -683 688 -683 0 3
rlabel polysilicon 695 -677 695 -677 0 1
rlabel polysilicon 695 -683 695 -683 0 3
rlabel polysilicon 702 -677 702 -677 0 1
rlabel polysilicon 702 -683 702 -683 0 3
rlabel polysilicon 709 -677 709 -677 0 1
rlabel polysilicon 709 -683 709 -683 0 3
rlabel polysilicon 716 -677 716 -677 0 1
rlabel polysilicon 716 -683 716 -683 0 3
rlabel polysilicon 723 -677 723 -677 0 1
rlabel polysilicon 723 -683 723 -683 0 3
rlabel polysilicon 730 -677 730 -677 0 1
rlabel polysilicon 730 -683 730 -683 0 3
rlabel polysilicon 737 -677 737 -677 0 1
rlabel polysilicon 737 -683 737 -683 0 3
rlabel polysilicon 744 -677 744 -677 0 1
rlabel polysilicon 744 -683 744 -683 0 3
rlabel polysilicon 751 -677 751 -677 0 1
rlabel polysilicon 751 -683 751 -683 0 3
rlabel polysilicon 758 -677 758 -677 0 1
rlabel polysilicon 758 -683 758 -683 0 3
rlabel polysilicon 765 -677 765 -677 0 1
rlabel polysilicon 765 -683 765 -683 0 3
rlabel polysilicon 772 -677 772 -677 0 1
rlabel polysilicon 772 -683 772 -683 0 3
rlabel polysilicon 16 -762 16 -762 0 1
rlabel polysilicon 19 -768 19 -768 0 4
rlabel polysilicon 23 -768 23 -768 0 3
rlabel polysilicon 30 -762 30 -762 0 1
rlabel polysilicon 37 -762 37 -762 0 1
rlabel polysilicon 37 -768 37 -768 0 3
rlabel polysilicon 44 -762 44 -762 0 1
rlabel polysilicon 44 -768 44 -768 0 3
rlabel polysilicon 54 -762 54 -762 0 2
rlabel polysilicon 58 -762 58 -762 0 1
rlabel polysilicon 58 -768 58 -768 0 3
rlabel polysilicon 65 -762 65 -762 0 1
rlabel polysilicon 65 -768 65 -768 0 3
rlabel polysilicon 72 -762 72 -762 0 1
rlabel polysilicon 72 -768 72 -768 0 3
rlabel polysilicon 79 -762 79 -762 0 1
rlabel polysilicon 79 -768 79 -768 0 3
rlabel polysilicon 86 -762 86 -762 0 1
rlabel polysilicon 89 -762 89 -762 0 2
rlabel polysilicon 86 -768 86 -768 0 3
rlabel polysilicon 89 -768 89 -768 0 4
rlabel polysilicon 93 -762 93 -762 0 1
rlabel polysilicon 96 -762 96 -762 0 2
rlabel polysilicon 96 -768 96 -768 0 4
rlabel polysilicon 100 -762 100 -762 0 1
rlabel polysilicon 100 -768 100 -768 0 3
rlabel polysilicon 107 -762 107 -762 0 1
rlabel polysilicon 107 -768 107 -768 0 3
rlabel polysilicon 114 -762 114 -762 0 1
rlabel polysilicon 117 -768 117 -768 0 4
rlabel polysilicon 124 -762 124 -762 0 2
rlabel polysilicon 121 -768 121 -768 0 3
rlabel polysilicon 131 -762 131 -762 0 2
rlabel polysilicon 128 -768 128 -768 0 3
rlabel polysilicon 135 -762 135 -762 0 1
rlabel polysilicon 135 -768 135 -768 0 3
rlabel polysilicon 142 -762 142 -762 0 1
rlabel polysilicon 142 -768 142 -768 0 3
rlabel polysilicon 149 -762 149 -762 0 1
rlabel polysilicon 149 -768 149 -768 0 3
rlabel polysilicon 152 -768 152 -768 0 4
rlabel polysilicon 156 -762 156 -762 0 1
rlabel polysilicon 156 -768 156 -768 0 3
rlabel polysilicon 163 -762 163 -762 0 1
rlabel polysilicon 163 -768 163 -768 0 3
rlabel polysilicon 170 -762 170 -762 0 1
rlabel polysilicon 170 -768 170 -768 0 3
rlabel polysilicon 177 -762 177 -762 0 1
rlabel polysilicon 177 -768 177 -768 0 3
rlabel polysilicon 184 -762 184 -762 0 1
rlabel polysilicon 184 -768 184 -768 0 3
rlabel polysilicon 191 -762 191 -762 0 1
rlabel polysilicon 191 -768 191 -768 0 3
rlabel polysilicon 201 -762 201 -762 0 2
rlabel polysilicon 198 -768 198 -768 0 3
rlabel polysilicon 201 -768 201 -768 0 4
rlabel polysilicon 205 -762 205 -762 0 1
rlabel polysilicon 212 -762 212 -762 0 1
rlabel polysilicon 212 -768 212 -768 0 3
rlabel polysilicon 222 -762 222 -762 0 2
rlabel polysilicon 219 -768 219 -768 0 3
rlabel polysilicon 222 -768 222 -768 0 4
rlabel polysilicon 226 -762 226 -762 0 1
rlabel polysilicon 226 -768 226 -768 0 3
rlabel polysilicon 233 -762 233 -762 0 1
rlabel polysilicon 233 -768 233 -768 0 3
rlabel polysilicon 240 -762 240 -762 0 1
rlabel polysilicon 240 -768 240 -768 0 3
rlabel polysilicon 243 -768 243 -768 0 4
rlabel polysilicon 247 -762 247 -762 0 1
rlabel polysilicon 247 -768 247 -768 0 3
rlabel polysilicon 254 -762 254 -762 0 1
rlabel polysilicon 254 -768 254 -768 0 3
rlabel polysilicon 261 -762 261 -762 0 1
rlabel polysilicon 261 -768 261 -768 0 3
rlabel polysilicon 268 -762 268 -762 0 1
rlabel polysilicon 268 -768 268 -768 0 3
rlabel polysilicon 275 -762 275 -762 0 1
rlabel polysilicon 275 -768 275 -768 0 3
rlabel polysilicon 282 -762 282 -762 0 1
rlabel polysilicon 282 -768 282 -768 0 3
rlabel polysilicon 289 -762 289 -762 0 1
rlabel polysilicon 292 -762 292 -762 0 2
rlabel polysilicon 289 -768 289 -768 0 3
rlabel polysilicon 292 -768 292 -768 0 4
rlabel polysilicon 296 -762 296 -762 0 1
rlabel polysilicon 296 -768 296 -768 0 3
rlabel polysilicon 303 -762 303 -762 0 1
rlabel polysilicon 306 -762 306 -762 0 2
rlabel polysilicon 306 -768 306 -768 0 4
rlabel polysilicon 313 -762 313 -762 0 2
rlabel polysilicon 310 -768 310 -768 0 3
rlabel polysilicon 320 -762 320 -762 0 2
rlabel polysilicon 317 -768 317 -768 0 3
rlabel polysilicon 320 -768 320 -768 0 4
rlabel polysilicon 324 -762 324 -762 0 1
rlabel polysilicon 324 -768 324 -768 0 3
rlabel polysilicon 331 -762 331 -762 0 1
rlabel polysilicon 331 -768 331 -768 0 3
rlabel polysilicon 338 -762 338 -762 0 1
rlabel polysilicon 338 -768 338 -768 0 3
rlabel polysilicon 345 -762 345 -762 0 1
rlabel polysilicon 348 -762 348 -762 0 2
rlabel polysilicon 352 -762 352 -762 0 1
rlabel polysilicon 355 -762 355 -762 0 2
rlabel polysilicon 352 -768 352 -768 0 3
rlabel polysilicon 355 -768 355 -768 0 4
rlabel polysilicon 362 -762 362 -762 0 2
rlabel polysilicon 359 -768 359 -768 0 3
rlabel polysilicon 366 -762 366 -762 0 1
rlabel polysilicon 366 -768 366 -768 0 3
rlabel polysilicon 373 -762 373 -762 0 1
rlabel polysilicon 373 -768 373 -768 0 3
rlabel polysilicon 383 -762 383 -762 0 2
rlabel polysilicon 380 -768 380 -768 0 3
rlabel polysilicon 387 -762 387 -762 0 1
rlabel polysilicon 387 -768 387 -768 0 3
rlabel polysilicon 394 -762 394 -762 0 1
rlabel polysilicon 397 -762 397 -762 0 2
rlabel polysilicon 397 -768 397 -768 0 4
rlabel polysilicon 401 -762 401 -762 0 1
rlabel polysilicon 401 -768 401 -768 0 3
rlabel polysilicon 408 -762 408 -762 0 1
rlabel polysilicon 408 -768 408 -768 0 3
rlabel polysilicon 415 -762 415 -762 0 1
rlabel polysilicon 415 -768 415 -768 0 3
rlabel polysilicon 422 -762 422 -762 0 1
rlabel polysilicon 422 -768 422 -768 0 3
rlabel polysilicon 429 -762 429 -762 0 1
rlabel polysilicon 429 -768 429 -768 0 3
rlabel polysilicon 432 -768 432 -768 0 4
rlabel polysilicon 436 -762 436 -762 0 1
rlabel polysilicon 439 -762 439 -762 0 2
rlabel polysilicon 446 -762 446 -762 0 2
rlabel polysilicon 443 -768 443 -768 0 3
rlabel polysilicon 446 -768 446 -768 0 4
rlabel polysilicon 450 -762 450 -762 0 1
rlabel polysilicon 450 -768 450 -768 0 3
rlabel polysilicon 457 -762 457 -762 0 1
rlabel polysilicon 457 -768 457 -768 0 3
rlabel polysilicon 464 -762 464 -762 0 1
rlabel polysilicon 464 -768 464 -768 0 3
rlabel polysilicon 471 -762 471 -762 0 1
rlabel polysilicon 471 -768 471 -768 0 3
rlabel polysilicon 478 -762 478 -762 0 1
rlabel polysilicon 481 -762 481 -762 0 2
rlabel polysilicon 488 -762 488 -762 0 2
rlabel polysilicon 488 -768 488 -768 0 4
rlabel polysilicon 492 -762 492 -762 0 1
rlabel polysilicon 492 -768 492 -768 0 3
rlabel polysilicon 499 -762 499 -762 0 1
rlabel polysilicon 499 -768 499 -768 0 3
rlabel polysilicon 506 -762 506 -762 0 1
rlabel polysilicon 506 -768 506 -768 0 3
rlabel polysilicon 513 -762 513 -762 0 1
rlabel polysilicon 513 -768 513 -768 0 3
rlabel polysilicon 520 -762 520 -762 0 1
rlabel polysilicon 520 -768 520 -768 0 3
rlabel polysilicon 527 -762 527 -762 0 1
rlabel polysilicon 527 -768 527 -768 0 3
rlabel polysilicon 534 -762 534 -762 0 1
rlabel polysilicon 534 -768 534 -768 0 3
rlabel polysilicon 537 -768 537 -768 0 4
rlabel polysilicon 541 -762 541 -762 0 1
rlabel polysilicon 541 -768 541 -768 0 3
rlabel polysilicon 548 -762 548 -762 0 1
rlabel polysilicon 548 -768 548 -768 0 3
rlabel polysilicon 555 -762 555 -762 0 1
rlabel polysilicon 555 -768 555 -768 0 3
rlabel polysilicon 562 -762 562 -762 0 1
rlabel polysilicon 562 -768 562 -768 0 3
rlabel polysilicon 569 -762 569 -762 0 1
rlabel polysilicon 569 -768 569 -768 0 3
rlabel polysilicon 576 -762 576 -762 0 1
rlabel polysilicon 576 -768 576 -768 0 3
rlabel polysilicon 583 -762 583 -762 0 1
rlabel polysilicon 583 -768 583 -768 0 3
rlabel polysilicon 590 -762 590 -762 0 1
rlabel polysilicon 590 -768 590 -768 0 3
rlabel polysilicon 597 -762 597 -762 0 1
rlabel polysilicon 597 -768 597 -768 0 3
rlabel polysilicon 604 -762 604 -762 0 1
rlabel polysilicon 604 -768 604 -768 0 3
rlabel polysilicon 611 -762 611 -762 0 1
rlabel polysilicon 611 -768 611 -768 0 3
rlabel polysilicon 621 -762 621 -762 0 2
rlabel polysilicon 621 -768 621 -768 0 4
rlabel polysilicon 625 -762 625 -762 0 1
rlabel polysilicon 625 -768 625 -768 0 3
rlabel polysilicon 632 -762 632 -762 0 1
rlabel polysilicon 632 -768 632 -768 0 3
rlabel polysilicon 639 -762 639 -762 0 1
rlabel polysilicon 639 -768 639 -768 0 3
rlabel polysilicon 646 -762 646 -762 0 1
rlabel polysilicon 646 -768 646 -768 0 3
rlabel polysilicon 653 -762 653 -762 0 1
rlabel polysilicon 653 -768 653 -768 0 3
rlabel polysilicon 660 -762 660 -762 0 1
rlabel polysilicon 660 -768 660 -768 0 3
rlabel polysilicon 667 -762 667 -762 0 1
rlabel polysilicon 667 -768 667 -768 0 3
rlabel polysilicon 674 -762 674 -762 0 1
rlabel polysilicon 674 -768 674 -768 0 3
rlabel polysilicon 681 -762 681 -762 0 1
rlabel polysilicon 681 -768 681 -768 0 3
rlabel polysilicon 688 -762 688 -762 0 1
rlabel polysilicon 688 -768 688 -768 0 3
rlabel polysilicon 695 -762 695 -762 0 1
rlabel polysilicon 695 -768 695 -768 0 3
rlabel polysilicon 702 -762 702 -762 0 1
rlabel polysilicon 702 -768 702 -768 0 3
rlabel polysilicon 709 -762 709 -762 0 1
rlabel polysilicon 709 -768 709 -768 0 3
rlabel polysilicon 716 -762 716 -762 0 1
rlabel polysilicon 716 -768 716 -768 0 3
rlabel polysilicon 723 -762 723 -762 0 1
rlabel polysilicon 723 -768 723 -768 0 3
rlabel polysilicon 733 -762 733 -762 0 2
rlabel polysilicon 737 -762 737 -762 0 1
rlabel polysilicon 737 -768 737 -768 0 3
rlabel polysilicon 744 -762 744 -762 0 1
rlabel polysilicon 744 -768 744 -768 0 3
rlabel polysilicon 751 -762 751 -762 0 1
rlabel polysilicon 751 -768 751 -768 0 3
rlabel polysilicon 758 -762 758 -762 0 1
rlabel polysilicon 758 -768 758 -768 0 3
rlabel polysilicon 765 -762 765 -762 0 1
rlabel polysilicon 765 -768 765 -768 0 3
rlabel polysilicon 772 -762 772 -762 0 1
rlabel polysilicon 772 -768 772 -768 0 3
rlabel polysilicon 779 -762 779 -762 0 1
rlabel polysilicon 779 -768 779 -768 0 3
rlabel polysilicon 786 -762 786 -762 0 1
rlabel polysilicon 786 -768 786 -768 0 3
rlabel polysilicon 793 -762 793 -762 0 1
rlabel polysilicon 793 -768 793 -768 0 3
rlabel polysilicon 849 -762 849 -762 0 1
rlabel polysilicon 849 -768 849 -768 0 3
rlabel polysilicon 19 -857 19 -857 0 4
rlabel polysilicon 23 -851 23 -851 0 1
rlabel polysilicon 23 -857 23 -857 0 3
rlabel polysilicon 30 -851 30 -851 0 1
rlabel polysilicon 30 -857 30 -857 0 3
rlabel polysilicon 37 -851 37 -851 0 1
rlabel polysilicon 40 -851 40 -851 0 2
rlabel polysilicon 44 -851 44 -851 0 1
rlabel polysilicon 44 -857 44 -857 0 3
rlabel polysilicon 54 -851 54 -851 0 2
rlabel polysilicon 51 -857 51 -857 0 3
rlabel polysilicon 58 -851 58 -851 0 1
rlabel polysilicon 58 -857 58 -857 0 3
rlabel polysilicon 65 -851 65 -851 0 1
rlabel polysilicon 65 -857 65 -857 0 3
rlabel polysilicon 72 -851 72 -851 0 1
rlabel polysilicon 72 -857 72 -857 0 3
rlabel polysilicon 75 -857 75 -857 0 4
rlabel polysilicon 79 -851 79 -851 0 1
rlabel polysilicon 79 -857 79 -857 0 3
rlabel polysilicon 86 -851 86 -851 0 1
rlabel polysilicon 89 -851 89 -851 0 2
rlabel polysilicon 86 -857 86 -857 0 3
rlabel polysilicon 93 -851 93 -851 0 1
rlabel polysilicon 93 -857 93 -857 0 3
rlabel polysilicon 100 -851 100 -851 0 1
rlabel polysilicon 100 -857 100 -857 0 3
rlabel polysilicon 103 -857 103 -857 0 4
rlabel polysilicon 107 -851 107 -851 0 1
rlabel polysilicon 107 -857 107 -857 0 3
rlabel polysilicon 114 -851 114 -851 0 1
rlabel polysilicon 114 -857 114 -857 0 3
rlabel polysilicon 121 -851 121 -851 0 1
rlabel polysilicon 121 -857 121 -857 0 3
rlabel polysilicon 128 -851 128 -851 0 1
rlabel polysilicon 128 -857 128 -857 0 3
rlabel polysilicon 135 -851 135 -851 0 1
rlabel polysilicon 135 -857 135 -857 0 3
rlabel polysilicon 142 -851 142 -851 0 1
rlabel polysilicon 142 -857 142 -857 0 3
rlabel polysilicon 145 -857 145 -857 0 4
rlabel polysilicon 149 -851 149 -851 0 1
rlabel polysilicon 152 -851 152 -851 0 2
rlabel polysilicon 156 -851 156 -851 0 1
rlabel polysilicon 159 -851 159 -851 0 2
rlabel polysilicon 156 -857 156 -857 0 3
rlabel polysilicon 159 -857 159 -857 0 4
rlabel polysilicon 163 -851 163 -851 0 1
rlabel polysilicon 166 -851 166 -851 0 2
rlabel polysilicon 163 -857 163 -857 0 3
rlabel polysilicon 170 -851 170 -851 0 1
rlabel polysilicon 170 -857 170 -857 0 3
rlabel polysilicon 177 -851 177 -851 0 1
rlabel polysilicon 177 -857 177 -857 0 3
rlabel polysilicon 184 -851 184 -851 0 1
rlabel polysilicon 184 -857 184 -857 0 3
rlabel polysilicon 191 -851 191 -851 0 1
rlabel polysilicon 191 -857 191 -857 0 3
rlabel polysilicon 198 -851 198 -851 0 1
rlabel polysilicon 198 -857 198 -857 0 3
rlabel polysilicon 205 -857 205 -857 0 3
rlabel polysilicon 212 -851 212 -851 0 1
rlabel polysilicon 212 -857 212 -857 0 3
rlabel polysilicon 219 -851 219 -851 0 1
rlabel polysilicon 219 -857 219 -857 0 3
rlabel polysilicon 226 -851 226 -851 0 1
rlabel polysilicon 226 -857 226 -857 0 3
rlabel polysilicon 233 -851 233 -851 0 1
rlabel polysilicon 233 -857 233 -857 0 3
rlabel polysilicon 240 -851 240 -851 0 1
rlabel polysilicon 243 -851 243 -851 0 2
rlabel polysilicon 240 -857 240 -857 0 3
rlabel polysilicon 250 -851 250 -851 0 2
rlabel polysilicon 254 -851 254 -851 0 1
rlabel polysilicon 254 -857 254 -857 0 3
rlabel polysilicon 261 -857 261 -857 0 3
rlabel polysilicon 264 -857 264 -857 0 4
rlabel polysilicon 268 -851 268 -851 0 1
rlabel polysilicon 268 -857 268 -857 0 3
rlabel polysilicon 275 -851 275 -851 0 1
rlabel polysilicon 275 -857 275 -857 0 3
rlabel polysilicon 282 -851 282 -851 0 1
rlabel polysilicon 282 -857 282 -857 0 3
rlabel polysilicon 289 -851 289 -851 0 1
rlabel polysilicon 289 -857 289 -857 0 3
rlabel polysilicon 296 -851 296 -851 0 1
rlabel polysilicon 299 -851 299 -851 0 2
rlabel polysilicon 296 -857 296 -857 0 3
rlabel polysilicon 306 -851 306 -851 0 2
rlabel polysilicon 303 -857 303 -857 0 3
rlabel polysilicon 306 -857 306 -857 0 4
rlabel polysilicon 310 -851 310 -851 0 1
rlabel polysilicon 310 -857 310 -857 0 3
rlabel polysilicon 317 -851 317 -851 0 1
rlabel polysilicon 317 -857 317 -857 0 3
rlabel polysilicon 324 -851 324 -851 0 1
rlabel polysilicon 327 -851 327 -851 0 2
rlabel polysilicon 327 -857 327 -857 0 4
rlabel polysilicon 331 -851 331 -851 0 1
rlabel polysilicon 331 -857 331 -857 0 3
rlabel polysilicon 334 -857 334 -857 0 4
rlabel polysilicon 338 -851 338 -851 0 1
rlabel polysilicon 338 -857 338 -857 0 3
rlabel polysilicon 345 -851 345 -851 0 1
rlabel polysilicon 345 -857 345 -857 0 3
rlabel polysilicon 352 -851 352 -851 0 1
rlabel polysilicon 352 -857 352 -857 0 3
rlabel polysilicon 359 -851 359 -851 0 1
rlabel polysilicon 362 -851 362 -851 0 2
rlabel polysilicon 359 -857 359 -857 0 3
rlabel polysilicon 362 -857 362 -857 0 4
rlabel polysilicon 366 -851 366 -851 0 1
rlabel polysilicon 366 -857 366 -857 0 3
rlabel polysilicon 373 -851 373 -851 0 1
rlabel polysilicon 373 -857 373 -857 0 3
rlabel polysilicon 383 -851 383 -851 0 2
rlabel polysilicon 380 -857 380 -857 0 3
rlabel polysilicon 387 -851 387 -851 0 1
rlabel polysilicon 387 -857 387 -857 0 3
rlabel polysilicon 394 -851 394 -851 0 1
rlabel polysilicon 397 -851 397 -851 0 2
rlabel polysilicon 401 -851 401 -851 0 1
rlabel polysilicon 401 -857 401 -857 0 3
rlabel polysilicon 408 -851 408 -851 0 1
rlabel polysilicon 411 -851 411 -851 0 2
rlabel polysilicon 411 -857 411 -857 0 4
rlabel polysilicon 415 -851 415 -851 0 1
rlabel polysilicon 415 -857 415 -857 0 3
rlabel polysilicon 422 -851 422 -851 0 1
rlabel polysilicon 422 -857 422 -857 0 3
rlabel polysilicon 429 -851 429 -851 0 1
rlabel polysilicon 432 -851 432 -851 0 2
rlabel polysilicon 429 -857 429 -857 0 3
rlabel polysilicon 436 -851 436 -851 0 1
rlabel polysilicon 439 -857 439 -857 0 4
rlabel polysilicon 446 -851 446 -851 0 2
rlabel polysilicon 446 -857 446 -857 0 4
rlabel polysilicon 450 -851 450 -851 0 1
rlabel polysilicon 457 -851 457 -851 0 1
rlabel polysilicon 460 -851 460 -851 0 2
rlabel polysilicon 460 -857 460 -857 0 4
rlabel polysilicon 464 -851 464 -851 0 1
rlabel polysilicon 467 -851 467 -851 0 2
rlabel polysilicon 471 -851 471 -851 0 1
rlabel polysilicon 471 -857 471 -857 0 3
rlabel polysilicon 478 -851 478 -851 0 1
rlabel polysilicon 478 -857 478 -857 0 3
rlabel polysilicon 485 -851 485 -851 0 1
rlabel polysilicon 485 -857 485 -857 0 3
rlabel polysilicon 492 -851 492 -851 0 1
rlabel polysilicon 492 -857 492 -857 0 3
rlabel polysilicon 499 -851 499 -851 0 1
rlabel polysilicon 499 -857 499 -857 0 3
rlabel polysilicon 506 -851 506 -851 0 1
rlabel polysilicon 506 -857 506 -857 0 3
rlabel polysilicon 513 -851 513 -851 0 1
rlabel polysilicon 516 -851 516 -851 0 2
rlabel polysilicon 516 -857 516 -857 0 4
rlabel polysilicon 520 -851 520 -851 0 1
rlabel polysilicon 520 -857 520 -857 0 3
rlabel polysilicon 527 -851 527 -851 0 1
rlabel polysilicon 527 -857 527 -857 0 3
rlabel polysilicon 534 -851 534 -851 0 1
rlabel polysilicon 534 -857 534 -857 0 3
rlabel polysilicon 541 -851 541 -851 0 1
rlabel polysilicon 541 -857 541 -857 0 3
rlabel polysilicon 548 -851 548 -851 0 1
rlabel polysilicon 548 -857 548 -857 0 3
rlabel polysilicon 555 -851 555 -851 0 1
rlabel polysilicon 555 -857 555 -857 0 3
rlabel polysilicon 562 -851 562 -851 0 1
rlabel polysilicon 562 -857 562 -857 0 3
rlabel polysilicon 569 -851 569 -851 0 1
rlabel polysilicon 569 -857 569 -857 0 3
rlabel polysilicon 576 -851 576 -851 0 1
rlabel polysilicon 576 -857 576 -857 0 3
rlabel polysilicon 583 -851 583 -851 0 1
rlabel polysilicon 583 -857 583 -857 0 3
rlabel polysilicon 590 -851 590 -851 0 1
rlabel polysilicon 590 -857 590 -857 0 3
rlabel polysilicon 597 -851 597 -851 0 1
rlabel polysilicon 597 -857 597 -857 0 3
rlabel polysilicon 604 -851 604 -851 0 1
rlabel polysilicon 604 -857 604 -857 0 3
rlabel polysilicon 611 -851 611 -851 0 1
rlabel polysilicon 611 -857 611 -857 0 3
rlabel polysilicon 618 -851 618 -851 0 1
rlabel polysilicon 618 -857 618 -857 0 3
rlabel polysilicon 625 -851 625 -851 0 1
rlabel polysilicon 625 -857 625 -857 0 3
rlabel polysilicon 632 -851 632 -851 0 1
rlabel polysilicon 632 -857 632 -857 0 3
rlabel polysilicon 639 -851 639 -851 0 1
rlabel polysilicon 639 -857 639 -857 0 3
rlabel polysilicon 646 -851 646 -851 0 1
rlabel polysilicon 646 -857 646 -857 0 3
rlabel polysilicon 653 -851 653 -851 0 1
rlabel polysilicon 653 -857 653 -857 0 3
rlabel polysilicon 660 -851 660 -851 0 1
rlabel polysilicon 660 -857 660 -857 0 3
rlabel polysilicon 667 -851 667 -851 0 1
rlabel polysilicon 667 -857 667 -857 0 3
rlabel polysilicon 674 -851 674 -851 0 1
rlabel polysilicon 674 -857 674 -857 0 3
rlabel polysilicon 681 -851 681 -851 0 1
rlabel polysilicon 681 -857 681 -857 0 3
rlabel polysilicon 688 -851 688 -851 0 1
rlabel polysilicon 688 -857 688 -857 0 3
rlabel polysilicon 695 -851 695 -851 0 1
rlabel polysilicon 695 -857 695 -857 0 3
rlabel polysilicon 702 -851 702 -851 0 1
rlabel polysilicon 702 -857 702 -857 0 3
rlabel polysilicon 709 -851 709 -851 0 1
rlabel polysilicon 709 -857 709 -857 0 3
rlabel polysilicon 716 -851 716 -851 0 1
rlabel polysilicon 716 -857 716 -857 0 3
rlabel polysilicon 723 -851 723 -851 0 1
rlabel polysilicon 723 -857 723 -857 0 3
rlabel polysilicon 730 -851 730 -851 0 1
rlabel polysilicon 730 -857 730 -857 0 3
rlabel polysilicon 737 -851 737 -851 0 1
rlabel polysilicon 737 -857 737 -857 0 3
rlabel polysilicon 744 -851 744 -851 0 1
rlabel polysilicon 744 -857 744 -857 0 3
rlabel polysilicon 751 -851 751 -851 0 1
rlabel polysilicon 751 -857 751 -857 0 3
rlabel polysilicon 758 -851 758 -851 0 1
rlabel polysilicon 758 -857 758 -857 0 3
rlabel polysilicon 765 -851 765 -851 0 1
rlabel polysilicon 765 -857 765 -857 0 3
rlabel polysilicon 772 -851 772 -851 0 1
rlabel polysilicon 772 -857 772 -857 0 3
rlabel polysilicon 779 -851 779 -851 0 1
rlabel polysilicon 779 -857 779 -857 0 3
rlabel polysilicon 786 -851 786 -851 0 1
rlabel polysilicon 786 -857 786 -857 0 3
rlabel polysilicon 800 -851 800 -851 0 1
rlabel polysilicon 800 -857 800 -857 0 3
rlabel polysilicon 807 -851 807 -851 0 1
rlabel polysilicon 807 -857 807 -857 0 3
rlabel polysilicon 814 -851 814 -851 0 1
rlabel polysilicon 814 -857 814 -857 0 3
rlabel polysilicon 821 -851 821 -851 0 1
rlabel polysilicon 821 -857 821 -857 0 3
rlabel polysilicon 828 -851 828 -851 0 1
rlabel polysilicon 828 -857 828 -857 0 3
rlabel polysilicon 835 -851 835 -851 0 1
rlabel polysilicon 835 -857 835 -857 0 3
rlabel polysilicon 842 -851 842 -851 0 1
rlabel polysilicon 842 -857 842 -857 0 3
rlabel polysilicon 849 -851 849 -851 0 1
rlabel polysilicon 849 -857 849 -857 0 3
rlabel polysilicon 856 -851 856 -851 0 1
rlabel polysilicon 856 -857 856 -857 0 3
rlabel polysilicon 863 -851 863 -851 0 1
rlabel polysilicon 863 -857 863 -857 0 3
rlabel polysilicon 870 -851 870 -851 0 1
rlabel polysilicon 870 -857 870 -857 0 3
rlabel polysilicon 940 -851 940 -851 0 1
rlabel polysilicon 940 -857 940 -857 0 3
rlabel polysilicon 9 -928 9 -928 0 1
rlabel polysilicon 9 -934 9 -934 0 3
rlabel polysilicon 16 -928 16 -928 0 1
rlabel polysilicon 16 -934 16 -934 0 3
rlabel polysilicon 23 -928 23 -928 0 1
rlabel polysilicon 23 -934 23 -934 0 3
rlabel polysilicon 30 -928 30 -928 0 1
rlabel polysilicon 30 -934 30 -934 0 3
rlabel polysilicon 40 -928 40 -928 0 2
rlabel polysilicon 40 -934 40 -934 0 4
rlabel polysilicon 44 -928 44 -928 0 1
rlabel polysilicon 44 -934 44 -934 0 3
rlabel polysilicon 51 -928 51 -928 0 1
rlabel polysilicon 54 -928 54 -928 0 2
rlabel polysilicon 58 -928 58 -928 0 1
rlabel polysilicon 58 -934 58 -934 0 3
rlabel polysilicon 65 -934 65 -934 0 3
rlabel polysilicon 72 -928 72 -928 0 1
rlabel polysilicon 72 -934 72 -934 0 3
rlabel polysilicon 79 -928 79 -928 0 1
rlabel polysilicon 82 -928 82 -928 0 2
rlabel polysilicon 82 -934 82 -934 0 4
rlabel polysilicon 86 -928 86 -928 0 1
rlabel polysilicon 86 -934 86 -934 0 3
rlabel polysilicon 93 -928 93 -928 0 1
rlabel polysilicon 93 -934 93 -934 0 3
rlabel polysilicon 100 -928 100 -928 0 1
rlabel polysilicon 100 -934 100 -934 0 3
rlabel polysilicon 107 -928 107 -928 0 1
rlabel polysilicon 107 -934 107 -934 0 3
rlabel polysilicon 114 -928 114 -928 0 1
rlabel polysilicon 114 -934 114 -934 0 3
rlabel polysilicon 124 -928 124 -928 0 2
rlabel polysilicon 121 -934 121 -934 0 3
rlabel polysilicon 124 -934 124 -934 0 4
rlabel polysilicon 128 -928 128 -928 0 1
rlabel polysilicon 128 -934 128 -934 0 3
rlabel polysilicon 135 -928 135 -928 0 1
rlabel polysilicon 135 -934 135 -934 0 3
rlabel polysilicon 142 -928 142 -928 0 1
rlabel polysilicon 142 -934 142 -934 0 3
rlabel polysilicon 149 -928 149 -928 0 1
rlabel polysilicon 152 -934 152 -934 0 4
rlabel polysilicon 156 -928 156 -928 0 1
rlabel polysilicon 156 -934 156 -934 0 3
rlabel polysilicon 163 -928 163 -928 0 1
rlabel polysilicon 166 -928 166 -928 0 2
rlabel polysilicon 170 -928 170 -928 0 1
rlabel polysilicon 170 -934 170 -934 0 3
rlabel polysilicon 177 -928 177 -928 0 1
rlabel polysilicon 177 -934 177 -934 0 3
rlabel polysilicon 184 -928 184 -928 0 1
rlabel polysilicon 184 -934 184 -934 0 3
rlabel polysilicon 191 -928 191 -928 0 1
rlabel polysilicon 191 -934 191 -934 0 3
rlabel polysilicon 198 -928 198 -928 0 1
rlabel polysilicon 201 -928 201 -928 0 2
rlabel polysilicon 201 -934 201 -934 0 4
rlabel polysilicon 205 -928 205 -928 0 1
rlabel polysilicon 208 -934 208 -934 0 4
rlabel polysilicon 215 -928 215 -928 0 2
rlabel polysilicon 215 -934 215 -934 0 4
rlabel polysilicon 219 -928 219 -928 0 1
rlabel polysilicon 222 -928 222 -928 0 2
rlabel polysilicon 226 -928 226 -928 0 1
rlabel polysilicon 226 -934 226 -934 0 3
rlabel polysilicon 233 -928 233 -928 0 1
rlabel polysilicon 233 -934 233 -934 0 3
rlabel polysilicon 240 -928 240 -928 0 1
rlabel polysilicon 240 -934 240 -934 0 3
rlabel polysilicon 250 -928 250 -928 0 2
rlabel polysilicon 247 -934 247 -934 0 3
rlabel polysilicon 254 -928 254 -928 0 1
rlabel polysilicon 254 -934 254 -934 0 3
rlabel polysilicon 261 -928 261 -928 0 1
rlabel polysilicon 261 -934 261 -934 0 3
rlabel polysilicon 268 -928 268 -928 0 1
rlabel polysilicon 268 -934 268 -934 0 3
rlabel polysilicon 278 -928 278 -928 0 2
rlabel polysilicon 278 -934 278 -934 0 4
rlabel polysilicon 282 -928 282 -928 0 1
rlabel polysilicon 285 -934 285 -934 0 4
rlabel polysilicon 289 -928 289 -928 0 1
rlabel polysilicon 289 -934 289 -934 0 3
rlabel polysilicon 299 -928 299 -928 0 2
rlabel polysilicon 296 -934 296 -934 0 3
rlabel polysilicon 299 -934 299 -934 0 4
rlabel polysilicon 303 -928 303 -928 0 1
rlabel polysilicon 303 -934 303 -934 0 3
rlabel polysilicon 310 -928 310 -928 0 1
rlabel polysilicon 310 -934 310 -934 0 3
rlabel polysilicon 317 -928 317 -928 0 1
rlabel polysilicon 317 -934 317 -934 0 3
rlabel polysilicon 324 -928 324 -928 0 1
rlabel polysilicon 324 -934 324 -934 0 3
rlabel polysilicon 331 -928 331 -928 0 1
rlabel polysilicon 331 -934 331 -934 0 3
rlabel polysilicon 338 -928 338 -928 0 1
rlabel polysilicon 341 -928 341 -928 0 2
rlabel polysilicon 338 -934 338 -934 0 3
rlabel polysilicon 345 -928 345 -928 0 1
rlabel polysilicon 348 -928 348 -928 0 2
rlabel polysilicon 345 -934 345 -934 0 3
rlabel polysilicon 348 -934 348 -934 0 4
rlabel polysilicon 352 -934 352 -934 0 3
rlabel polysilicon 359 -928 359 -928 0 1
rlabel polysilicon 359 -934 359 -934 0 3
rlabel polysilicon 366 -928 366 -928 0 1
rlabel polysilicon 366 -934 366 -934 0 3
rlabel polysilicon 373 -928 373 -928 0 1
rlabel polysilicon 373 -934 373 -934 0 3
rlabel polysilicon 380 -928 380 -928 0 1
rlabel polysilicon 380 -934 380 -934 0 3
rlabel polysilicon 387 -928 387 -928 0 1
rlabel polysilicon 387 -934 387 -934 0 3
rlabel polysilicon 394 -934 394 -934 0 3
rlabel polysilicon 401 -928 401 -928 0 1
rlabel polysilicon 404 -928 404 -928 0 2
rlabel polysilicon 401 -934 401 -934 0 3
rlabel polysilicon 404 -934 404 -934 0 4
rlabel polysilicon 408 -928 408 -928 0 1
rlabel polysilicon 408 -934 408 -934 0 3
rlabel polysilicon 415 -928 415 -928 0 1
rlabel polysilicon 415 -934 415 -934 0 3
rlabel polysilicon 422 -928 422 -928 0 1
rlabel polysilicon 422 -934 422 -934 0 3
rlabel polysilicon 429 -928 429 -928 0 1
rlabel polysilicon 429 -934 429 -934 0 3
rlabel polysilicon 436 -928 436 -928 0 1
rlabel polysilicon 436 -934 436 -934 0 3
rlabel polysilicon 443 -928 443 -928 0 1
rlabel polysilicon 446 -928 446 -928 0 2
rlabel polysilicon 443 -934 443 -934 0 3
rlabel polysilicon 446 -934 446 -934 0 4
rlabel polysilicon 453 -928 453 -928 0 2
rlabel polysilicon 450 -934 450 -934 0 3
rlabel polysilicon 453 -934 453 -934 0 4
rlabel polysilicon 457 -928 457 -928 0 1
rlabel polysilicon 457 -934 457 -934 0 3
rlabel polysilicon 464 -928 464 -928 0 1
rlabel polysilicon 467 -928 467 -928 0 2
rlabel polysilicon 471 -928 471 -928 0 1
rlabel polysilicon 471 -934 471 -934 0 3
rlabel polysilicon 478 -928 478 -928 0 1
rlabel polysilicon 478 -934 478 -934 0 3
rlabel polysilicon 485 -928 485 -928 0 1
rlabel polysilicon 485 -934 485 -934 0 3
rlabel polysilicon 492 -928 492 -928 0 1
rlabel polysilicon 492 -934 492 -934 0 3
rlabel polysilicon 499 -928 499 -928 0 1
rlabel polysilicon 499 -934 499 -934 0 3
rlabel polysilicon 506 -928 506 -928 0 1
rlabel polysilicon 506 -934 506 -934 0 3
rlabel polysilicon 509 -934 509 -934 0 4
rlabel polysilicon 516 -928 516 -928 0 2
rlabel polysilicon 513 -934 513 -934 0 3
rlabel polysilicon 516 -934 516 -934 0 4
rlabel polysilicon 520 -928 520 -928 0 1
rlabel polysilicon 520 -934 520 -934 0 3
rlabel polysilicon 527 -928 527 -928 0 1
rlabel polysilicon 527 -934 527 -934 0 3
rlabel polysilicon 534 -928 534 -928 0 1
rlabel polysilicon 534 -934 534 -934 0 3
rlabel polysilicon 541 -934 541 -934 0 3
rlabel polysilicon 548 -928 548 -928 0 1
rlabel polysilicon 548 -934 548 -934 0 3
rlabel polysilicon 555 -928 555 -928 0 1
rlabel polysilicon 555 -934 555 -934 0 3
rlabel polysilicon 562 -928 562 -928 0 1
rlabel polysilicon 562 -934 562 -934 0 3
rlabel polysilicon 569 -928 569 -928 0 1
rlabel polysilicon 569 -934 569 -934 0 3
rlabel polysilicon 576 -928 576 -928 0 1
rlabel polysilicon 576 -934 576 -934 0 3
rlabel polysilicon 583 -928 583 -928 0 1
rlabel polysilicon 583 -934 583 -934 0 3
rlabel polysilicon 590 -928 590 -928 0 1
rlabel polysilicon 593 -928 593 -928 0 2
rlabel polysilicon 590 -934 590 -934 0 3
rlabel polysilicon 597 -928 597 -928 0 1
rlabel polysilicon 597 -934 597 -934 0 3
rlabel polysilicon 604 -928 604 -928 0 1
rlabel polysilicon 604 -934 604 -934 0 3
rlabel polysilicon 611 -928 611 -928 0 1
rlabel polysilicon 611 -934 611 -934 0 3
rlabel polysilicon 618 -928 618 -928 0 1
rlabel polysilicon 618 -934 618 -934 0 3
rlabel polysilicon 625 -928 625 -928 0 1
rlabel polysilicon 625 -934 625 -934 0 3
rlabel polysilicon 632 -928 632 -928 0 1
rlabel polysilicon 632 -934 632 -934 0 3
rlabel polysilicon 639 -928 639 -928 0 1
rlabel polysilicon 639 -934 639 -934 0 3
rlabel polysilicon 646 -928 646 -928 0 1
rlabel polysilicon 646 -934 646 -934 0 3
rlabel polysilicon 653 -928 653 -928 0 1
rlabel polysilicon 653 -934 653 -934 0 3
rlabel polysilicon 660 -928 660 -928 0 1
rlabel polysilicon 660 -934 660 -934 0 3
rlabel polysilicon 667 -928 667 -928 0 1
rlabel polysilicon 667 -934 667 -934 0 3
rlabel polysilicon 674 -928 674 -928 0 1
rlabel polysilicon 674 -934 674 -934 0 3
rlabel polysilicon 681 -928 681 -928 0 1
rlabel polysilicon 681 -934 681 -934 0 3
rlabel polysilicon 688 -928 688 -928 0 1
rlabel polysilicon 688 -934 688 -934 0 3
rlabel polysilicon 695 -928 695 -928 0 1
rlabel polysilicon 695 -934 695 -934 0 3
rlabel polysilicon 702 -928 702 -928 0 1
rlabel polysilicon 702 -934 702 -934 0 3
rlabel polysilicon 709 -928 709 -928 0 1
rlabel polysilicon 709 -934 709 -934 0 3
rlabel polysilicon 716 -928 716 -928 0 1
rlabel polysilicon 716 -934 716 -934 0 3
rlabel polysilicon 723 -928 723 -928 0 1
rlabel polysilicon 723 -934 723 -934 0 3
rlabel polysilicon 730 -928 730 -928 0 1
rlabel polysilicon 730 -934 730 -934 0 3
rlabel polysilicon 737 -928 737 -928 0 1
rlabel polysilicon 737 -934 737 -934 0 3
rlabel polysilicon 744 -928 744 -928 0 1
rlabel polysilicon 744 -934 744 -934 0 3
rlabel polysilicon 751 -928 751 -928 0 1
rlabel polysilicon 751 -934 751 -934 0 3
rlabel polysilicon 758 -928 758 -928 0 1
rlabel polysilicon 758 -934 758 -934 0 3
rlabel polysilicon 765 -928 765 -928 0 1
rlabel polysilicon 765 -934 765 -934 0 3
rlabel polysilicon 772 -928 772 -928 0 1
rlabel polysilicon 772 -934 772 -934 0 3
rlabel polysilicon 779 -928 779 -928 0 1
rlabel polysilicon 779 -934 779 -934 0 3
rlabel polysilicon 786 -928 786 -928 0 1
rlabel polysilicon 786 -934 786 -934 0 3
rlabel polysilicon 793 -928 793 -928 0 1
rlabel polysilicon 793 -934 793 -934 0 3
rlabel polysilicon 800 -928 800 -928 0 1
rlabel polysilicon 800 -934 800 -934 0 3
rlabel polysilicon 807 -928 807 -928 0 1
rlabel polysilicon 807 -934 807 -934 0 3
rlabel polysilicon 814 -928 814 -928 0 1
rlabel polysilicon 814 -934 814 -934 0 3
rlabel polysilicon 821 -928 821 -928 0 1
rlabel polysilicon 821 -934 821 -934 0 3
rlabel polysilicon 828 -928 828 -928 0 1
rlabel polysilicon 831 -928 831 -928 0 2
rlabel polysilicon 828 -934 828 -934 0 3
rlabel polysilicon 835 -928 835 -928 0 1
rlabel polysilicon 835 -934 835 -934 0 3
rlabel polysilicon 842 -928 842 -928 0 1
rlabel polysilicon 842 -934 842 -934 0 3
rlabel polysilicon 849 -928 849 -928 0 1
rlabel polysilicon 2 -1007 2 -1007 0 1
rlabel polysilicon 2 -1013 2 -1013 0 3
rlabel polysilicon 9 -1007 9 -1007 0 1
rlabel polysilicon 9 -1013 9 -1013 0 3
rlabel polysilicon 19 -1013 19 -1013 0 4
rlabel polysilicon 23 -1007 23 -1007 0 1
rlabel polysilicon 23 -1013 23 -1013 0 3
rlabel polysilicon 33 -1013 33 -1013 0 4
rlabel polysilicon 37 -1007 37 -1007 0 1
rlabel polysilicon 37 -1013 37 -1013 0 3
rlabel polysilicon 44 -1007 44 -1007 0 1
rlabel polysilicon 44 -1013 44 -1013 0 3
rlabel polysilicon 51 -1007 51 -1007 0 1
rlabel polysilicon 51 -1013 51 -1013 0 3
rlabel polysilicon 58 -1007 58 -1007 0 1
rlabel polysilicon 61 -1007 61 -1007 0 2
rlabel polysilicon 65 -1007 65 -1007 0 1
rlabel polysilicon 65 -1013 65 -1013 0 3
rlabel polysilicon 72 -1007 72 -1007 0 1
rlabel polysilicon 72 -1013 72 -1013 0 3
rlabel polysilicon 79 -1007 79 -1007 0 1
rlabel polysilicon 79 -1013 79 -1013 0 3
rlabel polysilicon 86 -1007 86 -1007 0 1
rlabel polysilicon 86 -1013 86 -1013 0 3
rlabel polysilicon 93 -1007 93 -1007 0 1
rlabel polysilicon 93 -1013 93 -1013 0 3
rlabel polysilicon 100 -1013 100 -1013 0 3
rlabel polysilicon 107 -1007 107 -1007 0 1
rlabel polysilicon 107 -1013 107 -1013 0 3
rlabel polysilicon 114 -1007 114 -1007 0 1
rlabel polysilicon 117 -1007 117 -1007 0 2
rlabel polysilicon 114 -1013 114 -1013 0 3
rlabel polysilicon 117 -1013 117 -1013 0 4
rlabel polysilicon 121 -1007 121 -1007 0 1
rlabel polysilicon 128 -1007 128 -1007 0 1
rlabel polysilicon 131 -1007 131 -1007 0 2
rlabel polysilicon 128 -1013 128 -1013 0 3
rlabel polysilicon 135 -1007 135 -1007 0 1
rlabel polysilicon 135 -1013 135 -1013 0 3
rlabel polysilicon 142 -1007 142 -1007 0 1
rlabel polysilicon 142 -1013 142 -1013 0 3
rlabel polysilicon 149 -1007 149 -1007 0 1
rlabel polysilicon 149 -1013 149 -1013 0 3
rlabel polysilicon 156 -1007 156 -1007 0 1
rlabel polysilicon 163 -1007 163 -1007 0 1
rlabel polysilicon 163 -1013 163 -1013 0 3
rlabel polysilicon 170 -1007 170 -1007 0 1
rlabel polysilicon 173 -1007 173 -1007 0 2
rlabel polysilicon 170 -1013 170 -1013 0 3
rlabel polysilicon 177 -1007 177 -1007 0 1
rlabel polysilicon 177 -1013 177 -1013 0 3
rlabel polysilicon 184 -1007 184 -1007 0 1
rlabel polysilicon 184 -1013 184 -1013 0 3
rlabel polysilicon 194 -1007 194 -1007 0 2
rlabel polysilicon 191 -1013 191 -1013 0 3
rlabel polysilicon 194 -1013 194 -1013 0 4
rlabel polysilicon 201 -1007 201 -1007 0 2
rlabel polysilicon 201 -1013 201 -1013 0 4
rlabel polysilicon 205 -1007 205 -1007 0 1
rlabel polysilicon 205 -1013 205 -1013 0 3
rlabel polysilicon 212 -1007 212 -1007 0 1
rlabel polysilicon 212 -1013 212 -1013 0 3
rlabel polysilicon 219 -1007 219 -1007 0 1
rlabel polysilicon 222 -1007 222 -1007 0 2
rlabel polysilicon 219 -1013 219 -1013 0 3
rlabel polysilicon 222 -1013 222 -1013 0 4
rlabel polysilicon 226 -1007 226 -1007 0 1
rlabel polysilicon 226 -1013 226 -1013 0 3
rlabel polysilicon 233 -1007 233 -1007 0 1
rlabel polysilicon 233 -1013 233 -1013 0 3
rlabel polysilicon 240 -1007 240 -1007 0 1
rlabel polysilicon 240 -1013 240 -1013 0 3
rlabel polysilicon 247 -1007 247 -1007 0 1
rlabel polysilicon 247 -1013 247 -1013 0 3
rlabel polysilicon 254 -1007 254 -1007 0 1
rlabel polysilicon 254 -1013 254 -1013 0 3
rlabel polysilicon 261 -1007 261 -1007 0 1
rlabel polysilicon 261 -1013 261 -1013 0 3
rlabel polysilicon 268 -1007 268 -1007 0 1
rlabel polysilicon 268 -1013 268 -1013 0 3
rlabel polysilicon 275 -1007 275 -1007 0 1
rlabel polysilicon 275 -1013 275 -1013 0 3
rlabel polysilicon 282 -1007 282 -1007 0 1
rlabel polysilicon 282 -1013 282 -1013 0 3
rlabel polysilicon 289 -1007 289 -1007 0 1
rlabel polysilicon 289 -1013 289 -1013 0 3
rlabel polysilicon 296 -1007 296 -1007 0 1
rlabel polysilicon 296 -1013 296 -1013 0 3
rlabel polysilicon 303 -1007 303 -1007 0 1
rlabel polysilicon 303 -1013 303 -1013 0 3
rlabel polysilicon 313 -1007 313 -1007 0 2
rlabel polysilicon 317 -1007 317 -1007 0 1
rlabel polysilicon 317 -1013 317 -1013 0 3
rlabel polysilicon 324 -1007 324 -1007 0 1
rlabel polysilicon 324 -1013 324 -1013 0 3
rlabel polysilicon 331 -1007 331 -1007 0 1
rlabel polysilicon 334 -1007 334 -1007 0 2
rlabel polysilicon 331 -1013 331 -1013 0 3
rlabel polysilicon 334 -1013 334 -1013 0 4
rlabel polysilicon 338 -1007 338 -1007 0 1
rlabel polysilicon 341 -1013 341 -1013 0 4
rlabel polysilicon 345 -1007 345 -1007 0 1
rlabel polysilicon 345 -1013 345 -1013 0 3
rlabel polysilicon 352 -1007 352 -1007 0 1
rlabel polysilicon 352 -1013 352 -1013 0 3
rlabel polysilicon 359 -1007 359 -1007 0 1
rlabel polysilicon 359 -1013 359 -1013 0 3
rlabel polysilicon 366 -1007 366 -1007 0 1
rlabel polysilicon 366 -1013 366 -1013 0 3
rlabel polysilicon 373 -1007 373 -1007 0 1
rlabel polysilicon 376 -1007 376 -1007 0 2
rlabel polysilicon 376 -1013 376 -1013 0 4
rlabel polysilicon 380 -1007 380 -1007 0 1
rlabel polysilicon 380 -1013 380 -1013 0 3
rlabel polysilicon 387 -1007 387 -1007 0 1
rlabel polysilicon 390 -1007 390 -1007 0 2
rlabel polysilicon 390 -1013 390 -1013 0 4
rlabel polysilicon 394 -1007 394 -1007 0 1
rlabel polysilicon 397 -1007 397 -1007 0 2
rlabel polysilicon 404 -1007 404 -1007 0 2
rlabel polysilicon 401 -1013 401 -1013 0 3
rlabel polysilicon 404 -1013 404 -1013 0 4
rlabel polysilicon 408 -1007 408 -1007 0 1
rlabel polysilicon 411 -1007 411 -1007 0 2
rlabel polysilicon 411 -1013 411 -1013 0 4
rlabel polysilicon 415 -1007 415 -1007 0 1
rlabel polysilicon 415 -1013 415 -1013 0 3
rlabel polysilicon 425 -1007 425 -1007 0 2
rlabel polysilicon 429 -1007 429 -1007 0 1
rlabel polysilicon 429 -1013 429 -1013 0 3
rlabel polysilicon 432 -1013 432 -1013 0 4
rlabel polysilicon 436 -1007 436 -1007 0 1
rlabel polysilicon 439 -1013 439 -1013 0 4
rlabel polysilicon 443 -1007 443 -1007 0 1
rlabel polysilicon 443 -1013 443 -1013 0 3
rlabel polysilicon 450 -1007 450 -1007 0 1
rlabel polysilicon 450 -1013 450 -1013 0 3
rlabel polysilicon 457 -1007 457 -1007 0 1
rlabel polysilicon 457 -1013 457 -1013 0 3
rlabel polysilicon 464 -1007 464 -1007 0 1
rlabel polysilicon 464 -1013 464 -1013 0 3
rlabel polysilicon 474 -1007 474 -1007 0 2
rlabel polysilicon 478 -1007 478 -1007 0 1
rlabel polysilicon 481 -1007 481 -1007 0 2
rlabel polysilicon 478 -1013 478 -1013 0 3
rlabel polysilicon 485 -1007 485 -1007 0 1
rlabel polysilicon 485 -1013 485 -1013 0 3
rlabel polysilicon 492 -1007 492 -1007 0 1
rlabel polysilicon 492 -1013 492 -1013 0 3
rlabel polysilicon 499 -1007 499 -1007 0 1
rlabel polysilicon 499 -1013 499 -1013 0 3
rlabel polysilicon 502 -1013 502 -1013 0 4
rlabel polysilicon 506 -1007 506 -1007 0 1
rlabel polysilicon 506 -1013 506 -1013 0 3
rlabel polysilicon 513 -1013 513 -1013 0 3
rlabel polysilicon 516 -1013 516 -1013 0 4
rlabel polysilicon 520 -1007 520 -1007 0 1
rlabel polysilicon 520 -1013 520 -1013 0 3
rlabel polysilicon 527 -1007 527 -1007 0 1
rlabel polysilicon 527 -1013 527 -1013 0 3
rlabel polysilicon 534 -1007 534 -1007 0 1
rlabel polysilicon 534 -1013 534 -1013 0 3
rlabel polysilicon 541 -1007 541 -1007 0 1
rlabel polysilicon 541 -1013 541 -1013 0 3
rlabel polysilicon 548 -1007 548 -1007 0 1
rlabel polysilicon 548 -1013 548 -1013 0 3
rlabel polysilicon 555 -1007 555 -1007 0 1
rlabel polysilicon 558 -1007 558 -1007 0 2
rlabel polysilicon 562 -1007 562 -1007 0 1
rlabel polysilicon 562 -1013 562 -1013 0 3
rlabel polysilicon 569 -1007 569 -1007 0 1
rlabel polysilicon 569 -1013 569 -1013 0 3
rlabel polysilicon 576 -1007 576 -1007 0 1
rlabel polysilicon 576 -1013 576 -1013 0 3
rlabel polysilicon 590 -1007 590 -1007 0 1
rlabel polysilicon 590 -1013 590 -1013 0 3
rlabel polysilicon 597 -1007 597 -1007 0 1
rlabel polysilicon 597 -1013 597 -1013 0 3
rlabel polysilicon 604 -1007 604 -1007 0 1
rlabel polysilicon 604 -1013 604 -1013 0 3
rlabel polysilicon 611 -1007 611 -1007 0 1
rlabel polysilicon 611 -1013 611 -1013 0 3
rlabel polysilicon 614 -1013 614 -1013 0 4
rlabel polysilicon 618 -1007 618 -1007 0 1
rlabel polysilicon 618 -1013 618 -1013 0 3
rlabel polysilicon 625 -1007 625 -1007 0 1
rlabel polysilicon 625 -1013 625 -1013 0 3
rlabel polysilicon 632 -1007 632 -1007 0 1
rlabel polysilicon 632 -1013 632 -1013 0 3
rlabel polysilicon 639 -1007 639 -1007 0 1
rlabel polysilicon 639 -1013 639 -1013 0 3
rlabel polysilicon 646 -1007 646 -1007 0 1
rlabel polysilicon 646 -1013 646 -1013 0 3
rlabel polysilicon 653 -1007 653 -1007 0 1
rlabel polysilicon 653 -1013 653 -1013 0 3
rlabel polysilicon 660 -1007 660 -1007 0 1
rlabel polysilicon 660 -1013 660 -1013 0 3
rlabel polysilicon 667 -1007 667 -1007 0 1
rlabel polysilicon 667 -1013 667 -1013 0 3
rlabel polysilicon 674 -1007 674 -1007 0 1
rlabel polysilicon 674 -1013 674 -1013 0 3
rlabel polysilicon 681 -1007 681 -1007 0 1
rlabel polysilicon 681 -1013 681 -1013 0 3
rlabel polysilicon 688 -1007 688 -1007 0 1
rlabel polysilicon 688 -1013 688 -1013 0 3
rlabel polysilicon 695 -1007 695 -1007 0 1
rlabel polysilicon 695 -1013 695 -1013 0 3
rlabel polysilicon 702 -1007 702 -1007 0 1
rlabel polysilicon 702 -1013 702 -1013 0 3
rlabel polysilicon 709 -1007 709 -1007 0 1
rlabel polysilicon 709 -1013 709 -1013 0 3
rlabel polysilicon 716 -1007 716 -1007 0 1
rlabel polysilicon 716 -1013 716 -1013 0 3
rlabel polysilicon 723 -1007 723 -1007 0 1
rlabel polysilicon 723 -1013 723 -1013 0 3
rlabel polysilicon 730 -1007 730 -1007 0 1
rlabel polysilicon 730 -1013 730 -1013 0 3
rlabel polysilicon 737 -1007 737 -1007 0 1
rlabel polysilicon 737 -1013 737 -1013 0 3
rlabel polysilicon 744 -1007 744 -1007 0 1
rlabel polysilicon 744 -1013 744 -1013 0 3
rlabel polysilicon 751 -1007 751 -1007 0 1
rlabel polysilicon 751 -1013 751 -1013 0 3
rlabel polysilicon 758 -1007 758 -1007 0 1
rlabel polysilicon 758 -1013 758 -1013 0 3
rlabel polysilicon 765 -1007 765 -1007 0 1
rlabel polysilicon 765 -1013 765 -1013 0 3
rlabel polysilicon 772 -1007 772 -1007 0 1
rlabel polysilicon 772 -1013 772 -1013 0 3
rlabel polysilicon 779 -1007 779 -1007 0 1
rlabel polysilicon 779 -1013 779 -1013 0 3
rlabel polysilicon 786 -1007 786 -1007 0 1
rlabel polysilicon 786 -1013 786 -1013 0 3
rlabel polysilicon 793 -1007 793 -1007 0 1
rlabel polysilicon 793 -1013 793 -1013 0 3
rlabel polysilicon 800 -1007 800 -1007 0 1
rlabel polysilicon 800 -1013 800 -1013 0 3
rlabel polysilicon 807 -1007 807 -1007 0 1
rlabel polysilicon 807 -1013 807 -1013 0 3
rlabel polysilicon 814 -1007 814 -1007 0 1
rlabel polysilicon 814 -1013 814 -1013 0 3
rlabel polysilicon 821 -1007 821 -1007 0 1
rlabel polysilicon 821 -1013 821 -1013 0 3
rlabel polysilicon 828 -1007 828 -1007 0 1
rlabel polysilicon 828 -1013 828 -1013 0 3
rlabel polysilicon 835 -1007 835 -1007 0 1
rlabel polysilicon 835 -1013 835 -1013 0 3
rlabel polysilicon 842 -1007 842 -1007 0 1
rlabel polysilicon 842 -1013 842 -1013 0 3
rlabel polysilicon 849 -1007 849 -1007 0 1
rlabel polysilicon 849 -1013 849 -1013 0 3
rlabel polysilicon 856 -1007 856 -1007 0 1
rlabel polysilicon 859 -1007 859 -1007 0 2
rlabel polysilicon 859 -1013 859 -1013 0 4
rlabel polysilicon 863 -1007 863 -1007 0 1
rlabel polysilicon 863 -1013 863 -1013 0 3
rlabel polysilicon 873 -1007 873 -1007 0 2
rlabel polysilicon 898 -1007 898 -1007 0 1
rlabel polysilicon 898 -1013 898 -1013 0 3
rlabel polysilicon 9 -1090 9 -1090 0 3
rlabel polysilicon 16 -1084 16 -1084 0 1
rlabel polysilicon 16 -1090 16 -1090 0 3
rlabel polysilicon 23 -1084 23 -1084 0 1
rlabel polysilicon 23 -1090 23 -1090 0 3
rlabel polysilicon 30 -1084 30 -1084 0 1
rlabel polysilicon 30 -1090 30 -1090 0 3
rlabel polysilicon 37 -1084 37 -1084 0 1
rlabel polysilicon 37 -1090 37 -1090 0 3
rlabel polysilicon 44 -1084 44 -1084 0 1
rlabel polysilicon 44 -1090 44 -1090 0 3
rlabel polysilicon 54 -1084 54 -1084 0 2
rlabel polysilicon 58 -1084 58 -1084 0 1
rlabel polysilicon 58 -1090 58 -1090 0 3
rlabel polysilicon 65 -1084 65 -1084 0 1
rlabel polysilicon 72 -1084 72 -1084 0 1
rlabel polysilicon 72 -1090 72 -1090 0 3
rlabel polysilicon 79 -1084 79 -1084 0 1
rlabel polysilicon 79 -1090 79 -1090 0 3
rlabel polysilicon 82 -1090 82 -1090 0 4
rlabel polysilicon 86 -1084 86 -1084 0 1
rlabel polysilicon 86 -1090 86 -1090 0 3
rlabel polysilicon 93 -1090 93 -1090 0 3
rlabel polysilicon 96 -1090 96 -1090 0 4
rlabel polysilicon 103 -1084 103 -1084 0 2
rlabel polysilicon 103 -1090 103 -1090 0 4
rlabel polysilicon 107 -1084 107 -1084 0 1
rlabel polysilicon 107 -1090 107 -1090 0 3
rlabel polysilicon 114 -1084 114 -1084 0 1
rlabel polysilicon 114 -1090 114 -1090 0 3
rlabel polysilicon 121 -1084 121 -1084 0 1
rlabel polysilicon 121 -1090 121 -1090 0 3
rlabel polysilicon 128 -1084 128 -1084 0 1
rlabel polysilicon 128 -1090 128 -1090 0 3
rlabel polysilicon 135 -1090 135 -1090 0 3
rlabel polysilicon 138 -1090 138 -1090 0 4
rlabel polysilicon 142 -1084 142 -1084 0 1
rlabel polysilicon 142 -1090 142 -1090 0 3
rlabel polysilicon 152 -1084 152 -1084 0 2
rlabel polysilicon 152 -1090 152 -1090 0 4
rlabel polysilicon 159 -1084 159 -1084 0 2
rlabel polysilicon 163 -1084 163 -1084 0 1
rlabel polysilicon 166 -1084 166 -1084 0 2
rlabel polysilicon 166 -1090 166 -1090 0 4
rlabel polysilicon 170 -1084 170 -1084 0 1
rlabel polysilicon 170 -1090 170 -1090 0 3
rlabel polysilicon 177 -1084 177 -1084 0 1
rlabel polysilicon 177 -1090 177 -1090 0 3
rlabel polysilicon 184 -1084 184 -1084 0 1
rlabel polysilicon 184 -1090 184 -1090 0 3
rlabel polysilicon 191 -1084 191 -1084 0 1
rlabel polysilicon 191 -1090 191 -1090 0 3
rlabel polysilicon 198 -1084 198 -1084 0 1
rlabel polysilicon 198 -1090 198 -1090 0 3
rlabel polysilicon 205 -1084 205 -1084 0 1
rlabel polysilicon 205 -1090 205 -1090 0 3
rlabel polysilicon 212 -1084 212 -1084 0 1
rlabel polysilicon 212 -1090 212 -1090 0 3
rlabel polysilicon 222 -1084 222 -1084 0 2
rlabel polysilicon 219 -1090 219 -1090 0 3
rlabel polysilicon 222 -1090 222 -1090 0 4
rlabel polysilicon 226 -1084 226 -1084 0 1
rlabel polysilicon 226 -1090 226 -1090 0 3
rlabel polysilicon 233 -1084 233 -1084 0 1
rlabel polysilicon 233 -1090 233 -1090 0 3
rlabel polysilicon 243 -1084 243 -1084 0 2
rlabel polysilicon 250 -1090 250 -1090 0 4
rlabel polysilicon 254 -1084 254 -1084 0 1
rlabel polysilicon 254 -1090 254 -1090 0 3
rlabel polysilicon 261 -1084 261 -1084 0 1
rlabel polysilicon 261 -1090 261 -1090 0 3
rlabel polysilicon 268 -1084 268 -1084 0 1
rlabel polysilicon 268 -1090 268 -1090 0 3
rlabel polysilicon 275 -1084 275 -1084 0 1
rlabel polysilicon 278 -1084 278 -1084 0 2
rlabel polysilicon 278 -1090 278 -1090 0 4
rlabel polysilicon 282 -1084 282 -1084 0 1
rlabel polysilicon 282 -1090 282 -1090 0 3
rlabel polysilicon 289 -1084 289 -1084 0 1
rlabel polysilicon 289 -1090 289 -1090 0 3
rlabel polysilicon 296 -1084 296 -1084 0 1
rlabel polysilicon 296 -1090 296 -1090 0 3
rlabel polysilicon 303 -1084 303 -1084 0 1
rlabel polysilicon 303 -1090 303 -1090 0 3
rlabel polysilicon 310 -1084 310 -1084 0 1
rlabel polysilicon 310 -1090 310 -1090 0 3
rlabel polysilicon 317 -1084 317 -1084 0 1
rlabel polysilicon 317 -1090 317 -1090 0 3
rlabel polysilicon 324 -1084 324 -1084 0 1
rlabel polysilicon 324 -1090 324 -1090 0 3
rlabel polysilicon 331 -1084 331 -1084 0 1
rlabel polysilicon 331 -1090 331 -1090 0 3
rlabel polysilicon 338 -1084 338 -1084 0 1
rlabel polysilicon 338 -1090 338 -1090 0 3
rlabel polysilicon 345 -1084 345 -1084 0 1
rlabel polysilicon 348 -1084 348 -1084 0 2
rlabel polysilicon 348 -1090 348 -1090 0 4
rlabel polysilicon 352 -1084 352 -1084 0 1
rlabel polysilicon 355 -1090 355 -1090 0 4
rlabel polysilicon 359 -1084 359 -1084 0 1
rlabel polysilicon 359 -1090 359 -1090 0 3
rlabel polysilicon 366 -1084 366 -1084 0 1
rlabel polysilicon 366 -1090 366 -1090 0 3
rlabel polysilicon 373 -1084 373 -1084 0 1
rlabel polysilicon 373 -1090 373 -1090 0 3
rlabel polysilicon 380 -1084 380 -1084 0 1
rlabel polysilicon 380 -1090 380 -1090 0 3
rlabel polysilicon 387 -1084 387 -1084 0 1
rlabel polysilicon 390 -1084 390 -1084 0 2
rlabel polysilicon 390 -1090 390 -1090 0 4
rlabel polysilicon 394 -1084 394 -1084 0 1
rlabel polysilicon 394 -1090 394 -1090 0 3
rlabel polysilicon 401 -1084 401 -1084 0 1
rlabel polysilicon 401 -1090 401 -1090 0 3
rlabel polysilicon 408 -1084 408 -1084 0 1
rlabel polysilicon 408 -1090 408 -1090 0 3
rlabel polysilicon 415 -1084 415 -1084 0 1
rlabel polysilicon 415 -1090 415 -1090 0 3
rlabel polysilicon 422 -1084 422 -1084 0 1
rlabel polysilicon 422 -1090 422 -1090 0 3
rlabel polysilicon 429 -1084 429 -1084 0 1
rlabel polysilicon 429 -1090 429 -1090 0 3
rlabel polysilicon 436 -1084 436 -1084 0 1
rlabel polysilicon 436 -1090 436 -1090 0 3
rlabel polysilicon 446 -1084 446 -1084 0 2
rlabel polysilicon 446 -1090 446 -1090 0 4
rlabel polysilicon 450 -1084 450 -1084 0 1
rlabel polysilicon 453 -1084 453 -1084 0 2
rlabel polysilicon 450 -1090 450 -1090 0 3
rlabel polysilicon 453 -1090 453 -1090 0 4
rlabel polysilicon 457 -1084 457 -1084 0 1
rlabel polysilicon 457 -1090 457 -1090 0 3
rlabel polysilicon 467 -1084 467 -1084 0 2
rlabel polysilicon 464 -1090 464 -1090 0 3
rlabel polysilicon 471 -1084 471 -1084 0 1
rlabel polysilicon 471 -1090 471 -1090 0 3
rlabel polysilicon 478 -1084 478 -1084 0 1
rlabel polysilicon 478 -1090 478 -1090 0 3
rlabel polysilicon 485 -1084 485 -1084 0 1
rlabel polysilicon 485 -1090 485 -1090 0 3
rlabel polysilicon 492 -1084 492 -1084 0 1
rlabel polysilicon 495 -1084 495 -1084 0 2
rlabel polysilicon 492 -1090 492 -1090 0 3
rlabel polysilicon 499 -1084 499 -1084 0 1
rlabel polysilicon 499 -1090 499 -1090 0 3
rlabel polysilicon 506 -1084 506 -1084 0 1
rlabel polysilicon 506 -1090 506 -1090 0 3
rlabel polysilicon 513 -1084 513 -1084 0 1
rlabel polysilicon 513 -1090 513 -1090 0 3
rlabel polysilicon 520 -1084 520 -1084 0 1
rlabel polysilicon 520 -1090 520 -1090 0 3
rlabel polysilicon 527 -1084 527 -1084 0 1
rlabel polysilicon 530 -1084 530 -1084 0 2
rlabel polysilicon 527 -1090 527 -1090 0 3
rlabel polysilicon 530 -1090 530 -1090 0 4
rlabel polysilicon 534 -1084 534 -1084 0 1
rlabel polysilicon 537 -1084 537 -1084 0 2
rlabel polysilicon 541 -1084 541 -1084 0 1
rlabel polysilicon 541 -1090 541 -1090 0 3
rlabel polysilicon 548 -1084 548 -1084 0 1
rlabel polysilicon 551 -1084 551 -1084 0 2
rlabel polysilicon 558 -1084 558 -1084 0 2
rlabel polysilicon 558 -1090 558 -1090 0 4
rlabel polysilicon 562 -1084 562 -1084 0 1
rlabel polysilicon 565 -1084 565 -1084 0 2
rlabel polysilicon 562 -1090 562 -1090 0 3
rlabel polysilicon 572 -1084 572 -1084 0 2
rlabel polysilicon 569 -1090 569 -1090 0 3
rlabel polysilicon 572 -1090 572 -1090 0 4
rlabel polysilicon 576 -1084 576 -1084 0 1
rlabel polysilicon 576 -1090 576 -1090 0 3
rlabel polysilicon 583 -1084 583 -1084 0 1
rlabel polysilicon 583 -1090 583 -1090 0 3
rlabel polysilicon 590 -1084 590 -1084 0 1
rlabel polysilicon 590 -1090 590 -1090 0 3
rlabel polysilicon 597 -1084 597 -1084 0 1
rlabel polysilicon 597 -1090 597 -1090 0 3
rlabel polysilicon 604 -1084 604 -1084 0 1
rlabel polysilicon 607 -1084 607 -1084 0 2
rlabel polysilicon 604 -1090 604 -1090 0 3
rlabel polysilicon 607 -1090 607 -1090 0 4
rlabel polysilicon 611 -1084 611 -1084 0 1
rlabel polysilicon 614 -1084 614 -1084 0 2
rlabel polysilicon 611 -1090 611 -1090 0 3
rlabel polysilicon 618 -1084 618 -1084 0 1
rlabel polysilicon 618 -1090 618 -1090 0 3
rlabel polysilicon 625 -1084 625 -1084 0 1
rlabel polysilicon 625 -1090 625 -1090 0 3
rlabel polysilicon 632 -1084 632 -1084 0 1
rlabel polysilicon 632 -1090 632 -1090 0 3
rlabel polysilicon 642 -1084 642 -1084 0 2
rlabel polysilicon 639 -1090 639 -1090 0 3
rlabel polysilicon 642 -1090 642 -1090 0 4
rlabel polysilicon 646 -1084 646 -1084 0 1
rlabel polysilicon 646 -1090 646 -1090 0 3
rlabel polysilicon 653 -1084 653 -1084 0 1
rlabel polysilicon 653 -1090 653 -1090 0 3
rlabel polysilicon 660 -1084 660 -1084 0 1
rlabel polysilicon 660 -1090 660 -1090 0 3
rlabel polysilicon 667 -1084 667 -1084 0 1
rlabel polysilicon 667 -1090 667 -1090 0 3
rlabel polysilicon 674 -1084 674 -1084 0 1
rlabel polysilicon 674 -1090 674 -1090 0 3
rlabel polysilicon 681 -1084 681 -1084 0 1
rlabel polysilicon 681 -1090 681 -1090 0 3
rlabel polysilicon 688 -1084 688 -1084 0 1
rlabel polysilicon 688 -1090 688 -1090 0 3
rlabel polysilicon 695 -1084 695 -1084 0 1
rlabel polysilicon 695 -1090 695 -1090 0 3
rlabel polysilicon 702 -1084 702 -1084 0 1
rlabel polysilicon 702 -1090 702 -1090 0 3
rlabel polysilicon 709 -1084 709 -1084 0 1
rlabel polysilicon 709 -1090 709 -1090 0 3
rlabel polysilicon 716 -1084 716 -1084 0 1
rlabel polysilicon 716 -1090 716 -1090 0 3
rlabel polysilicon 723 -1084 723 -1084 0 1
rlabel polysilicon 723 -1090 723 -1090 0 3
rlabel polysilicon 730 -1084 730 -1084 0 1
rlabel polysilicon 730 -1090 730 -1090 0 3
rlabel polysilicon 737 -1084 737 -1084 0 1
rlabel polysilicon 737 -1090 737 -1090 0 3
rlabel polysilicon 744 -1084 744 -1084 0 1
rlabel polysilicon 744 -1090 744 -1090 0 3
rlabel polysilicon 751 -1084 751 -1084 0 1
rlabel polysilicon 751 -1090 751 -1090 0 3
rlabel polysilicon 758 -1084 758 -1084 0 1
rlabel polysilicon 758 -1090 758 -1090 0 3
rlabel polysilicon 765 -1084 765 -1084 0 1
rlabel polysilicon 765 -1090 765 -1090 0 3
rlabel polysilicon 772 -1084 772 -1084 0 1
rlabel polysilicon 772 -1090 772 -1090 0 3
rlabel polysilicon 779 -1084 779 -1084 0 1
rlabel polysilicon 779 -1090 779 -1090 0 3
rlabel polysilicon 786 -1084 786 -1084 0 1
rlabel polysilicon 786 -1090 786 -1090 0 3
rlabel polysilicon 793 -1084 793 -1084 0 1
rlabel polysilicon 793 -1090 793 -1090 0 3
rlabel polysilicon 800 -1084 800 -1084 0 1
rlabel polysilicon 800 -1090 800 -1090 0 3
rlabel polysilicon 807 -1084 807 -1084 0 1
rlabel polysilicon 807 -1090 807 -1090 0 3
rlabel polysilicon 814 -1084 814 -1084 0 1
rlabel polysilicon 814 -1090 814 -1090 0 3
rlabel polysilicon 821 -1084 821 -1084 0 1
rlabel polysilicon 821 -1090 821 -1090 0 3
rlabel polysilicon 828 -1084 828 -1084 0 1
rlabel polysilicon 828 -1090 828 -1090 0 3
rlabel polysilicon 835 -1084 835 -1084 0 1
rlabel polysilicon 835 -1090 835 -1090 0 3
rlabel polysilicon 842 -1084 842 -1084 0 1
rlabel polysilicon 842 -1090 842 -1090 0 3
rlabel polysilicon 849 -1084 849 -1084 0 1
rlabel polysilicon 849 -1090 849 -1090 0 3
rlabel polysilicon 856 -1084 856 -1084 0 1
rlabel polysilicon 856 -1090 856 -1090 0 3
rlabel polysilicon 863 -1084 863 -1084 0 1
rlabel polysilicon 863 -1090 863 -1090 0 3
rlabel polysilicon 870 -1084 870 -1084 0 1
rlabel polysilicon 870 -1090 870 -1090 0 3
rlabel polysilicon 877 -1084 877 -1084 0 1
rlabel polysilicon 877 -1090 877 -1090 0 3
rlabel polysilicon 884 -1084 884 -1084 0 1
rlabel polysilicon 884 -1090 884 -1090 0 3
rlabel polysilicon 891 -1084 891 -1084 0 1
rlabel polysilicon 891 -1090 891 -1090 0 3
rlabel polysilicon 898 -1084 898 -1084 0 1
rlabel polysilicon 898 -1090 898 -1090 0 3
rlabel polysilicon 905 -1084 905 -1084 0 1
rlabel polysilicon 905 -1090 905 -1090 0 3
rlabel polysilicon 912 -1084 912 -1084 0 1
rlabel polysilicon 912 -1090 912 -1090 0 3
rlabel polysilicon 919 -1084 919 -1084 0 1
rlabel polysilicon 919 -1090 919 -1090 0 3
rlabel polysilicon 926 -1084 926 -1084 0 1
rlabel polysilicon 926 -1090 926 -1090 0 3
rlabel polysilicon 929 -1090 929 -1090 0 4
rlabel polysilicon 940 -1084 940 -1084 0 1
rlabel polysilicon 940 -1090 940 -1090 0 3
rlabel polysilicon 5 -1187 5 -1187 0 4
rlabel polysilicon 9 -1181 9 -1181 0 1
rlabel polysilicon 9 -1187 9 -1187 0 3
rlabel polysilicon 16 -1181 16 -1181 0 1
rlabel polysilicon 16 -1187 16 -1187 0 3
rlabel polysilicon 26 -1187 26 -1187 0 4
rlabel polysilicon 30 -1181 30 -1181 0 1
rlabel polysilicon 30 -1187 30 -1187 0 3
rlabel polysilicon 37 -1181 37 -1181 0 1
rlabel polysilicon 37 -1187 37 -1187 0 3
rlabel polysilicon 44 -1181 44 -1181 0 1
rlabel polysilicon 44 -1187 44 -1187 0 3
rlabel polysilicon 51 -1181 51 -1181 0 1
rlabel polysilicon 51 -1187 51 -1187 0 3
rlabel polysilicon 58 -1181 58 -1181 0 1
rlabel polysilicon 58 -1187 58 -1187 0 3
rlabel polysilicon 65 -1181 65 -1181 0 1
rlabel polysilicon 65 -1187 65 -1187 0 3
rlabel polysilicon 72 -1181 72 -1181 0 1
rlabel polysilicon 79 -1181 79 -1181 0 1
rlabel polysilicon 79 -1187 79 -1187 0 3
rlabel polysilicon 86 -1181 86 -1181 0 1
rlabel polysilicon 86 -1187 86 -1187 0 3
rlabel polysilicon 93 -1181 93 -1181 0 1
rlabel polysilicon 93 -1187 93 -1187 0 3
rlabel polysilicon 96 -1187 96 -1187 0 4
rlabel polysilicon 103 -1181 103 -1181 0 2
rlabel polysilicon 103 -1187 103 -1187 0 4
rlabel polysilicon 107 -1181 107 -1181 0 1
rlabel polysilicon 107 -1187 107 -1187 0 3
rlabel polysilicon 114 -1181 114 -1181 0 1
rlabel polysilicon 114 -1187 114 -1187 0 3
rlabel polysilicon 121 -1187 121 -1187 0 3
rlabel polysilicon 124 -1187 124 -1187 0 4
rlabel polysilicon 128 -1181 128 -1181 0 1
rlabel polysilicon 128 -1187 128 -1187 0 3
rlabel polysilicon 135 -1181 135 -1181 0 1
rlabel polysilicon 135 -1187 135 -1187 0 3
rlabel polysilicon 142 -1181 142 -1181 0 1
rlabel polysilicon 142 -1187 142 -1187 0 3
rlabel polysilicon 152 -1181 152 -1181 0 2
rlabel polysilicon 149 -1187 149 -1187 0 3
rlabel polysilicon 152 -1187 152 -1187 0 4
rlabel polysilicon 156 -1181 156 -1181 0 1
rlabel polysilicon 156 -1187 156 -1187 0 3
rlabel polysilicon 163 -1181 163 -1181 0 1
rlabel polysilicon 163 -1187 163 -1187 0 3
rlabel polysilicon 170 -1181 170 -1181 0 1
rlabel polysilicon 173 -1187 173 -1187 0 4
rlabel polysilicon 177 -1181 177 -1181 0 1
rlabel polysilicon 177 -1187 177 -1187 0 3
rlabel polysilicon 184 -1181 184 -1181 0 1
rlabel polysilicon 184 -1187 184 -1187 0 3
rlabel polysilicon 191 -1181 191 -1181 0 1
rlabel polysilicon 191 -1187 191 -1187 0 3
rlabel polysilicon 198 -1181 198 -1181 0 1
rlabel polysilicon 201 -1181 201 -1181 0 2
rlabel polysilicon 198 -1187 198 -1187 0 3
rlabel polysilicon 201 -1187 201 -1187 0 4
rlabel polysilicon 205 -1181 205 -1181 0 1
rlabel polysilicon 205 -1187 205 -1187 0 3
rlabel polysilicon 212 -1181 212 -1181 0 1
rlabel polysilicon 212 -1187 212 -1187 0 3
rlabel polysilicon 215 -1187 215 -1187 0 4
rlabel polysilicon 222 -1181 222 -1181 0 2
rlabel polysilicon 219 -1187 219 -1187 0 3
rlabel polysilicon 222 -1187 222 -1187 0 4
rlabel polysilicon 226 -1181 226 -1181 0 1
rlabel polysilicon 226 -1187 226 -1187 0 3
rlabel polysilicon 233 -1181 233 -1181 0 1
rlabel polysilicon 233 -1187 233 -1187 0 3
rlabel polysilicon 240 -1181 240 -1181 0 1
rlabel polysilicon 240 -1187 240 -1187 0 3
rlabel polysilicon 247 -1181 247 -1181 0 1
rlabel polysilicon 247 -1187 247 -1187 0 3
rlabel polysilicon 254 -1181 254 -1181 0 1
rlabel polysilicon 254 -1187 254 -1187 0 3
rlabel polysilicon 261 -1181 261 -1181 0 1
rlabel polysilicon 261 -1187 261 -1187 0 3
rlabel polysilicon 268 -1181 268 -1181 0 1
rlabel polysilicon 268 -1187 268 -1187 0 3
rlabel polysilicon 275 -1181 275 -1181 0 1
rlabel polysilicon 275 -1187 275 -1187 0 3
rlabel polysilicon 282 -1181 282 -1181 0 1
rlabel polysilicon 282 -1187 282 -1187 0 3
rlabel polysilicon 285 -1187 285 -1187 0 4
rlabel polysilicon 289 -1181 289 -1181 0 1
rlabel polysilicon 289 -1187 289 -1187 0 3
rlabel polysilicon 296 -1181 296 -1181 0 1
rlabel polysilicon 296 -1187 296 -1187 0 3
rlabel polysilicon 303 -1181 303 -1181 0 1
rlabel polysilicon 303 -1187 303 -1187 0 3
rlabel polysilicon 310 -1181 310 -1181 0 1
rlabel polysilicon 310 -1187 310 -1187 0 3
rlabel polysilicon 320 -1181 320 -1181 0 2
rlabel polysilicon 320 -1187 320 -1187 0 4
rlabel polysilicon 324 -1181 324 -1181 0 1
rlabel polysilicon 324 -1187 324 -1187 0 3
rlabel polysilicon 331 -1181 331 -1181 0 1
rlabel polysilicon 331 -1187 331 -1187 0 3
rlabel polysilicon 338 -1181 338 -1181 0 1
rlabel polysilicon 338 -1187 338 -1187 0 3
rlabel polysilicon 345 -1181 345 -1181 0 1
rlabel polysilicon 345 -1187 345 -1187 0 3
rlabel polysilicon 355 -1181 355 -1181 0 2
rlabel polysilicon 355 -1187 355 -1187 0 4
rlabel polysilicon 359 -1181 359 -1181 0 1
rlabel polysilicon 362 -1181 362 -1181 0 2
rlabel polysilicon 366 -1181 366 -1181 0 1
rlabel polysilicon 366 -1187 366 -1187 0 3
rlabel polysilicon 373 -1181 373 -1181 0 1
rlabel polysilicon 373 -1187 373 -1187 0 3
rlabel polysilicon 380 -1181 380 -1181 0 1
rlabel polysilicon 380 -1187 380 -1187 0 3
rlabel polysilicon 387 -1181 387 -1181 0 1
rlabel polysilicon 387 -1187 387 -1187 0 3
rlabel polysilicon 394 -1181 394 -1181 0 1
rlabel polysilicon 394 -1187 394 -1187 0 3
rlabel polysilicon 401 -1181 401 -1181 0 1
rlabel polysilicon 401 -1187 401 -1187 0 3
rlabel polysilicon 408 -1187 408 -1187 0 3
rlabel polysilicon 411 -1187 411 -1187 0 4
rlabel polysilicon 415 -1181 415 -1181 0 1
rlabel polysilicon 415 -1187 415 -1187 0 3
rlabel polysilicon 422 -1181 422 -1181 0 1
rlabel polysilicon 425 -1181 425 -1181 0 2
rlabel polysilicon 425 -1187 425 -1187 0 4
rlabel polysilicon 429 -1181 429 -1181 0 1
rlabel polysilicon 429 -1187 429 -1187 0 3
rlabel polysilicon 436 -1181 436 -1181 0 1
rlabel polysilicon 436 -1187 436 -1187 0 3
rlabel polysilicon 443 -1181 443 -1181 0 1
rlabel polysilicon 443 -1187 443 -1187 0 3
rlabel polysilicon 450 -1181 450 -1181 0 1
rlabel polysilicon 453 -1181 453 -1181 0 2
rlabel polysilicon 450 -1187 450 -1187 0 3
rlabel polysilicon 453 -1187 453 -1187 0 4
rlabel polysilicon 457 -1181 457 -1181 0 1
rlabel polysilicon 457 -1187 457 -1187 0 3
rlabel polysilicon 464 -1187 464 -1187 0 3
rlabel polysilicon 467 -1187 467 -1187 0 4
rlabel polysilicon 471 -1181 471 -1181 0 1
rlabel polysilicon 471 -1187 471 -1187 0 3
rlabel polysilicon 478 -1181 478 -1181 0 1
rlabel polysilicon 478 -1187 478 -1187 0 3
rlabel polysilicon 485 -1181 485 -1181 0 1
rlabel polysilicon 485 -1187 485 -1187 0 3
rlabel polysilicon 492 -1181 492 -1181 0 1
rlabel polysilicon 492 -1187 492 -1187 0 3
rlabel polysilicon 499 -1181 499 -1181 0 1
rlabel polysilicon 499 -1187 499 -1187 0 3
rlabel polysilicon 506 -1181 506 -1181 0 1
rlabel polysilicon 509 -1181 509 -1181 0 2
rlabel polysilicon 506 -1187 506 -1187 0 3
rlabel polysilicon 513 -1181 513 -1181 0 1
rlabel polysilicon 513 -1187 513 -1187 0 3
rlabel polysilicon 520 -1181 520 -1181 0 1
rlabel polysilicon 520 -1187 520 -1187 0 3
rlabel polysilicon 527 -1181 527 -1181 0 1
rlabel polysilicon 527 -1187 527 -1187 0 3
rlabel polysilicon 534 -1181 534 -1181 0 1
rlabel polysilicon 534 -1187 534 -1187 0 3
rlabel polysilicon 541 -1181 541 -1181 0 1
rlabel polysilicon 544 -1181 544 -1181 0 2
rlabel polysilicon 541 -1187 541 -1187 0 3
rlabel polysilicon 544 -1187 544 -1187 0 4
rlabel polysilicon 548 -1181 548 -1181 0 1
rlabel polysilicon 548 -1187 548 -1187 0 3
rlabel polysilicon 555 -1181 555 -1181 0 1
rlabel polysilicon 555 -1187 555 -1187 0 3
rlabel polysilicon 562 -1181 562 -1181 0 1
rlabel polysilicon 562 -1187 562 -1187 0 3
rlabel polysilicon 569 -1181 569 -1181 0 1
rlabel polysilicon 569 -1187 569 -1187 0 3
rlabel polysilicon 579 -1181 579 -1181 0 2
rlabel polysilicon 579 -1187 579 -1187 0 4
rlabel polysilicon 583 -1181 583 -1181 0 1
rlabel polysilicon 583 -1187 583 -1187 0 3
rlabel polysilicon 590 -1181 590 -1181 0 1
rlabel polysilicon 590 -1187 590 -1187 0 3
rlabel polysilicon 597 -1181 597 -1181 0 1
rlabel polysilicon 597 -1187 597 -1187 0 3
rlabel polysilicon 604 -1181 604 -1181 0 1
rlabel polysilicon 604 -1187 604 -1187 0 3
rlabel polysilicon 611 -1181 611 -1181 0 1
rlabel polysilicon 611 -1187 611 -1187 0 3
rlabel polysilicon 618 -1181 618 -1181 0 1
rlabel polysilicon 625 -1181 625 -1181 0 1
rlabel polysilicon 625 -1187 625 -1187 0 3
rlabel polysilicon 632 -1181 632 -1181 0 1
rlabel polysilicon 632 -1187 632 -1187 0 3
rlabel polysilicon 639 -1181 639 -1181 0 1
rlabel polysilicon 639 -1187 639 -1187 0 3
rlabel polysilicon 646 -1181 646 -1181 0 1
rlabel polysilicon 646 -1187 646 -1187 0 3
rlabel polysilicon 656 -1181 656 -1181 0 2
rlabel polysilicon 656 -1187 656 -1187 0 4
rlabel polysilicon 660 -1181 660 -1181 0 1
rlabel polysilicon 660 -1187 660 -1187 0 3
rlabel polysilicon 667 -1181 667 -1181 0 1
rlabel polysilicon 667 -1187 667 -1187 0 3
rlabel polysilicon 674 -1181 674 -1181 0 1
rlabel polysilicon 674 -1187 674 -1187 0 3
rlabel polysilicon 681 -1181 681 -1181 0 1
rlabel polysilicon 684 -1181 684 -1181 0 2
rlabel polysilicon 688 -1181 688 -1181 0 1
rlabel polysilicon 688 -1187 688 -1187 0 3
rlabel polysilicon 695 -1181 695 -1181 0 1
rlabel polysilicon 695 -1187 695 -1187 0 3
rlabel polysilicon 702 -1181 702 -1181 0 1
rlabel polysilicon 702 -1187 702 -1187 0 3
rlabel polysilicon 709 -1181 709 -1181 0 1
rlabel polysilicon 709 -1187 709 -1187 0 3
rlabel polysilicon 716 -1181 716 -1181 0 1
rlabel polysilicon 719 -1187 719 -1187 0 4
rlabel polysilicon 723 -1181 723 -1181 0 1
rlabel polysilicon 723 -1187 723 -1187 0 3
rlabel polysilicon 730 -1181 730 -1181 0 1
rlabel polysilicon 730 -1187 730 -1187 0 3
rlabel polysilicon 737 -1181 737 -1181 0 1
rlabel polysilicon 737 -1187 737 -1187 0 3
rlabel polysilicon 744 -1181 744 -1181 0 1
rlabel polysilicon 744 -1187 744 -1187 0 3
rlabel polysilicon 751 -1181 751 -1181 0 1
rlabel polysilicon 751 -1187 751 -1187 0 3
rlabel polysilicon 758 -1181 758 -1181 0 1
rlabel polysilicon 758 -1187 758 -1187 0 3
rlabel polysilicon 765 -1181 765 -1181 0 1
rlabel polysilicon 765 -1187 765 -1187 0 3
rlabel polysilicon 772 -1181 772 -1181 0 1
rlabel polysilicon 772 -1187 772 -1187 0 3
rlabel polysilicon 779 -1181 779 -1181 0 1
rlabel polysilicon 779 -1187 779 -1187 0 3
rlabel polysilicon 786 -1181 786 -1181 0 1
rlabel polysilicon 786 -1187 786 -1187 0 3
rlabel polysilicon 793 -1181 793 -1181 0 1
rlabel polysilicon 793 -1187 793 -1187 0 3
rlabel polysilicon 800 -1181 800 -1181 0 1
rlabel polysilicon 800 -1187 800 -1187 0 3
rlabel polysilicon 807 -1181 807 -1181 0 1
rlabel polysilicon 807 -1187 807 -1187 0 3
rlabel polysilicon 814 -1181 814 -1181 0 1
rlabel polysilicon 814 -1187 814 -1187 0 3
rlabel polysilicon 821 -1181 821 -1181 0 1
rlabel polysilicon 821 -1187 821 -1187 0 3
rlabel polysilicon 828 -1181 828 -1181 0 1
rlabel polysilicon 828 -1187 828 -1187 0 3
rlabel polysilicon 835 -1181 835 -1181 0 1
rlabel polysilicon 835 -1187 835 -1187 0 3
rlabel polysilicon 842 -1181 842 -1181 0 1
rlabel polysilicon 842 -1187 842 -1187 0 3
rlabel polysilicon 849 -1181 849 -1181 0 1
rlabel polysilicon 849 -1187 849 -1187 0 3
rlabel polysilicon 856 -1181 856 -1181 0 1
rlabel polysilicon 856 -1187 856 -1187 0 3
rlabel polysilicon 863 -1181 863 -1181 0 1
rlabel polysilicon 863 -1187 863 -1187 0 3
rlabel polysilicon 870 -1181 870 -1181 0 1
rlabel polysilicon 870 -1187 870 -1187 0 3
rlabel polysilicon 877 -1181 877 -1181 0 1
rlabel polysilicon 877 -1187 877 -1187 0 3
rlabel polysilicon 884 -1181 884 -1181 0 1
rlabel polysilicon 884 -1187 884 -1187 0 3
rlabel polysilicon 891 -1181 891 -1181 0 1
rlabel polysilicon 891 -1187 891 -1187 0 3
rlabel polysilicon 898 -1181 898 -1181 0 1
rlabel polysilicon 898 -1187 898 -1187 0 3
rlabel polysilicon 905 -1181 905 -1181 0 1
rlabel polysilicon 905 -1187 905 -1187 0 3
rlabel polysilicon 912 -1181 912 -1181 0 1
rlabel polysilicon 912 -1187 912 -1187 0 3
rlabel polysilicon 919 -1181 919 -1181 0 1
rlabel polysilicon 919 -1187 919 -1187 0 3
rlabel polysilicon 926 -1181 926 -1181 0 1
rlabel polysilicon 926 -1187 926 -1187 0 3
rlabel polysilicon 933 -1181 933 -1181 0 1
rlabel polysilicon 933 -1187 933 -1187 0 3
rlabel polysilicon 940 -1181 940 -1181 0 1
rlabel polysilicon 940 -1187 940 -1187 0 3
rlabel polysilicon 947 -1181 947 -1181 0 1
rlabel polysilicon 947 -1187 947 -1187 0 3
rlabel polysilicon 957 -1187 957 -1187 0 4
rlabel polysilicon 961 -1181 961 -1181 0 1
rlabel polysilicon 961 -1187 961 -1187 0 3
rlabel polysilicon 964 -1187 964 -1187 0 4
rlabel polysilicon 968 -1181 968 -1181 0 1
rlabel polysilicon 968 -1187 968 -1187 0 3
rlabel polysilicon 975 -1181 975 -1181 0 1
rlabel polysilicon 975 -1187 975 -1187 0 3
rlabel polysilicon 982 -1181 982 -1181 0 1
rlabel polysilicon 985 -1187 985 -1187 0 4
rlabel polysilicon 989 -1181 989 -1181 0 1
rlabel polysilicon 989 -1187 989 -1187 0 3
rlabel polysilicon 12 -1276 12 -1276 0 2
rlabel polysilicon 16 -1276 16 -1276 0 1
rlabel polysilicon 16 -1282 16 -1282 0 3
rlabel polysilicon 26 -1276 26 -1276 0 2
rlabel polysilicon 30 -1276 30 -1276 0 1
rlabel polysilicon 30 -1282 30 -1282 0 3
rlabel polysilicon 40 -1276 40 -1276 0 2
rlabel polysilicon 44 -1276 44 -1276 0 1
rlabel polysilicon 44 -1282 44 -1282 0 3
rlabel polysilicon 51 -1276 51 -1276 0 1
rlabel polysilicon 51 -1282 51 -1282 0 3
rlabel polysilicon 58 -1276 58 -1276 0 1
rlabel polysilicon 58 -1282 58 -1282 0 3
rlabel polysilicon 65 -1276 65 -1276 0 1
rlabel polysilicon 65 -1282 65 -1282 0 3
rlabel polysilicon 72 -1276 72 -1276 0 1
rlabel polysilicon 72 -1282 72 -1282 0 3
rlabel polysilicon 79 -1276 79 -1276 0 1
rlabel polysilicon 79 -1282 79 -1282 0 3
rlabel polysilicon 86 -1276 86 -1276 0 1
rlabel polysilicon 86 -1282 86 -1282 0 3
rlabel polysilicon 93 -1276 93 -1276 0 1
rlabel polysilicon 96 -1276 96 -1276 0 2
rlabel polysilicon 96 -1282 96 -1282 0 4
rlabel polysilicon 100 -1276 100 -1276 0 1
rlabel polysilicon 100 -1282 100 -1282 0 3
rlabel polysilicon 110 -1276 110 -1276 0 2
rlabel polysilicon 110 -1282 110 -1282 0 4
rlabel polysilicon 114 -1276 114 -1276 0 1
rlabel polysilicon 114 -1282 114 -1282 0 3
rlabel polysilicon 121 -1276 121 -1276 0 1
rlabel polysilicon 121 -1282 121 -1282 0 3
rlabel polysilicon 128 -1276 128 -1276 0 1
rlabel polysilicon 128 -1282 128 -1282 0 3
rlabel polysilicon 135 -1276 135 -1276 0 1
rlabel polysilicon 135 -1282 135 -1282 0 3
rlabel polysilicon 142 -1276 142 -1276 0 1
rlabel polysilicon 142 -1282 142 -1282 0 3
rlabel polysilicon 149 -1276 149 -1276 0 1
rlabel polysilicon 149 -1282 149 -1282 0 3
rlabel polysilicon 156 -1276 156 -1276 0 1
rlabel polysilicon 156 -1282 156 -1282 0 3
rlabel polysilicon 163 -1276 163 -1276 0 1
rlabel polysilicon 163 -1282 163 -1282 0 3
rlabel polysilicon 170 -1276 170 -1276 0 1
rlabel polysilicon 173 -1282 173 -1282 0 4
rlabel polysilicon 177 -1276 177 -1276 0 1
rlabel polysilicon 177 -1282 177 -1282 0 3
rlabel polysilicon 184 -1276 184 -1276 0 1
rlabel polysilicon 184 -1282 184 -1282 0 3
rlabel polysilicon 191 -1276 191 -1276 0 1
rlabel polysilicon 191 -1282 191 -1282 0 3
rlabel polysilicon 198 -1276 198 -1276 0 1
rlabel polysilicon 198 -1282 198 -1282 0 3
rlabel polysilicon 205 -1276 205 -1276 0 1
rlabel polysilicon 205 -1282 205 -1282 0 3
rlabel polysilicon 212 -1276 212 -1276 0 1
rlabel polysilicon 215 -1276 215 -1276 0 2
rlabel polysilicon 222 -1276 222 -1276 0 2
rlabel polysilicon 219 -1282 219 -1282 0 3
rlabel polysilicon 222 -1282 222 -1282 0 4
rlabel polysilicon 226 -1276 226 -1276 0 1
rlabel polysilicon 226 -1282 226 -1282 0 3
rlabel polysilicon 233 -1276 233 -1276 0 1
rlabel polysilicon 233 -1282 233 -1282 0 3
rlabel polysilicon 240 -1276 240 -1276 0 1
rlabel polysilicon 240 -1282 240 -1282 0 3
rlabel polysilicon 247 -1276 247 -1276 0 1
rlabel polysilicon 247 -1282 247 -1282 0 3
rlabel polysilicon 254 -1276 254 -1276 0 1
rlabel polysilicon 254 -1282 254 -1282 0 3
rlabel polysilicon 261 -1276 261 -1276 0 1
rlabel polysilicon 261 -1282 261 -1282 0 3
rlabel polysilicon 268 -1276 268 -1276 0 1
rlabel polysilicon 268 -1282 268 -1282 0 3
rlabel polysilicon 275 -1276 275 -1276 0 1
rlabel polysilicon 275 -1282 275 -1282 0 3
rlabel polysilicon 282 -1276 282 -1276 0 1
rlabel polysilicon 282 -1282 282 -1282 0 3
rlabel polysilicon 289 -1276 289 -1276 0 1
rlabel polysilicon 289 -1282 289 -1282 0 3
rlabel polysilicon 296 -1276 296 -1276 0 1
rlabel polysilicon 296 -1282 296 -1282 0 3
rlabel polysilicon 303 -1276 303 -1276 0 1
rlabel polysilicon 306 -1276 306 -1276 0 2
rlabel polysilicon 303 -1282 303 -1282 0 3
rlabel polysilicon 310 -1276 310 -1276 0 1
rlabel polysilicon 313 -1276 313 -1276 0 2
rlabel polysilicon 310 -1282 310 -1282 0 3
rlabel polysilicon 313 -1282 313 -1282 0 4
rlabel polysilicon 317 -1276 317 -1276 0 1
rlabel polysilicon 317 -1282 317 -1282 0 3
rlabel polysilicon 324 -1276 324 -1276 0 1
rlabel polysilicon 324 -1282 324 -1282 0 3
rlabel polysilicon 331 -1276 331 -1276 0 1
rlabel polysilicon 331 -1282 331 -1282 0 3
rlabel polysilicon 341 -1276 341 -1276 0 2
rlabel polysilicon 338 -1282 338 -1282 0 3
rlabel polysilicon 341 -1282 341 -1282 0 4
rlabel polysilicon 345 -1276 345 -1276 0 1
rlabel polysilicon 345 -1282 345 -1282 0 3
rlabel polysilicon 352 -1276 352 -1276 0 1
rlabel polysilicon 352 -1282 352 -1282 0 3
rlabel polysilicon 359 -1276 359 -1276 0 1
rlabel polysilicon 362 -1276 362 -1276 0 2
rlabel polysilicon 359 -1282 359 -1282 0 3
rlabel polysilicon 366 -1276 366 -1276 0 1
rlabel polysilicon 366 -1282 366 -1282 0 3
rlabel polysilicon 373 -1276 373 -1276 0 1
rlabel polysilicon 373 -1282 373 -1282 0 3
rlabel polysilicon 380 -1276 380 -1276 0 1
rlabel polysilicon 380 -1282 380 -1282 0 3
rlabel polysilicon 383 -1282 383 -1282 0 4
rlabel polysilicon 387 -1276 387 -1276 0 1
rlabel polysilicon 387 -1282 387 -1282 0 3
rlabel polysilicon 394 -1276 394 -1276 0 1
rlabel polysilicon 394 -1282 394 -1282 0 3
rlabel polysilicon 401 -1276 401 -1276 0 1
rlabel polysilicon 401 -1282 401 -1282 0 3
rlabel polysilicon 408 -1276 408 -1276 0 1
rlabel polysilicon 411 -1276 411 -1276 0 2
rlabel polysilicon 408 -1282 408 -1282 0 3
rlabel polysilicon 411 -1282 411 -1282 0 4
rlabel polysilicon 415 -1276 415 -1276 0 1
rlabel polysilicon 415 -1282 415 -1282 0 3
rlabel polysilicon 422 -1276 422 -1276 0 1
rlabel polysilicon 422 -1282 422 -1282 0 3
rlabel polysilicon 429 -1276 429 -1276 0 1
rlabel polysilicon 429 -1282 429 -1282 0 3
rlabel polysilicon 436 -1276 436 -1276 0 1
rlabel polysilicon 436 -1282 436 -1282 0 3
rlabel polysilicon 443 -1276 443 -1276 0 1
rlabel polysilicon 446 -1276 446 -1276 0 2
rlabel polysilicon 443 -1282 443 -1282 0 3
rlabel polysilicon 446 -1282 446 -1282 0 4
rlabel polysilicon 450 -1276 450 -1276 0 1
rlabel polysilicon 450 -1282 450 -1282 0 3
rlabel polysilicon 457 -1276 457 -1276 0 1
rlabel polysilicon 460 -1276 460 -1276 0 2
rlabel polysilicon 460 -1282 460 -1282 0 4
rlabel polysilicon 464 -1276 464 -1276 0 1
rlabel polysilicon 467 -1276 467 -1276 0 2
rlabel polysilicon 464 -1282 464 -1282 0 3
rlabel polysilicon 471 -1276 471 -1276 0 1
rlabel polysilicon 474 -1276 474 -1276 0 2
rlabel polysilicon 471 -1282 471 -1282 0 3
rlabel polysilicon 474 -1282 474 -1282 0 4
rlabel polysilicon 478 -1276 478 -1276 0 1
rlabel polysilicon 478 -1282 478 -1282 0 3
rlabel polysilicon 485 -1276 485 -1276 0 1
rlabel polysilicon 485 -1282 485 -1282 0 3
rlabel polysilicon 492 -1276 492 -1276 0 1
rlabel polysilicon 495 -1276 495 -1276 0 2
rlabel polysilicon 499 -1282 499 -1282 0 3
rlabel polysilicon 502 -1282 502 -1282 0 4
rlabel polysilicon 506 -1282 506 -1282 0 3
rlabel polysilicon 509 -1282 509 -1282 0 4
rlabel polysilicon 513 -1276 513 -1276 0 1
rlabel polysilicon 513 -1282 513 -1282 0 3
rlabel polysilicon 520 -1276 520 -1276 0 1
rlabel polysilicon 520 -1282 520 -1282 0 3
rlabel polysilicon 527 -1276 527 -1276 0 1
rlabel polysilicon 527 -1282 527 -1282 0 3
rlabel polysilicon 534 -1276 534 -1276 0 1
rlabel polysilicon 534 -1282 534 -1282 0 3
rlabel polysilicon 541 -1276 541 -1276 0 1
rlabel polysilicon 541 -1282 541 -1282 0 3
rlabel polysilicon 548 -1276 548 -1276 0 1
rlabel polysilicon 548 -1282 548 -1282 0 3
rlabel polysilicon 555 -1276 555 -1276 0 1
rlabel polysilicon 555 -1282 555 -1282 0 3
rlabel polysilicon 562 -1276 562 -1276 0 1
rlabel polysilicon 562 -1282 562 -1282 0 3
rlabel polysilicon 569 -1276 569 -1276 0 1
rlabel polysilicon 569 -1282 569 -1282 0 3
rlabel polysilicon 576 -1276 576 -1276 0 1
rlabel polysilicon 576 -1282 576 -1282 0 3
rlabel polysilicon 583 -1276 583 -1276 0 1
rlabel polysilicon 583 -1282 583 -1282 0 3
rlabel polysilicon 590 -1276 590 -1276 0 1
rlabel polysilicon 590 -1282 590 -1282 0 3
rlabel polysilicon 597 -1276 597 -1276 0 1
rlabel polysilicon 600 -1276 600 -1276 0 2
rlabel polysilicon 604 -1276 604 -1276 0 1
rlabel polysilicon 607 -1276 607 -1276 0 2
rlabel polysilicon 604 -1282 604 -1282 0 3
rlabel polysilicon 611 -1276 611 -1276 0 1
rlabel polysilicon 611 -1282 611 -1282 0 3
rlabel polysilicon 618 -1276 618 -1276 0 1
rlabel polysilicon 618 -1282 618 -1282 0 3
rlabel polysilicon 625 -1276 625 -1276 0 1
rlabel polysilicon 625 -1282 625 -1282 0 3
rlabel polysilicon 635 -1276 635 -1276 0 2
rlabel polysilicon 639 -1276 639 -1276 0 1
rlabel polysilicon 639 -1282 639 -1282 0 3
rlabel polysilicon 646 -1276 646 -1276 0 1
rlabel polysilicon 646 -1282 646 -1282 0 3
rlabel polysilicon 653 -1276 653 -1276 0 1
rlabel polysilicon 656 -1276 656 -1276 0 2
rlabel polysilicon 653 -1282 653 -1282 0 3
rlabel polysilicon 656 -1282 656 -1282 0 4
rlabel polysilicon 660 -1276 660 -1276 0 1
rlabel polysilicon 660 -1282 660 -1282 0 3
rlabel polysilicon 670 -1276 670 -1276 0 2
rlabel polysilicon 667 -1282 667 -1282 0 3
rlabel polysilicon 674 -1276 674 -1276 0 1
rlabel polysilicon 674 -1282 674 -1282 0 3
rlabel polysilicon 681 -1276 681 -1276 0 1
rlabel polysilicon 681 -1282 681 -1282 0 3
rlabel polysilicon 688 -1276 688 -1276 0 1
rlabel polysilicon 688 -1282 688 -1282 0 3
rlabel polysilicon 695 -1276 695 -1276 0 1
rlabel polysilicon 695 -1282 695 -1282 0 3
rlabel polysilicon 702 -1276 702 -1276 0 1
rlabel polysilicon 702 -1282 702 -1282 0 3
rlabel polysilicon 709 -1276 709 -1276 0 1
rlabel polysilicon 709 -1282 709 -1282 0 3
rlabel polysilicon 716 -1276 716 -1276 0 1
rlabel polysilicon 716 -1282 716 -1282 0 3
rlabel polysilicon 723 -1276 723 -1276 0 1
rlabel polysilicon 723 -1282 723 -1282 0 3
rlabel polysilicon 730 -1276 730 -1276 0 1
rlabel polysilicon 730 -1282 730 -1282 0 3
rlabel polysilicon 737 -1276 737 -1276 0 1
rlabel polysilicon 737 -1282 737 -1282 0 3
rlabel polysilicon 744 -1276 744 -1276 0 1
rlabel polysilicon 744 -1282 744 -1282 0 3
rlabel polysilicon 751 -1276 751 -1276 0 1
rlabel polysilicon 751 -1282 751 -1282 0 3
rlabel polysilicon 758 -1276 758 -1276 0 1
rlabel polysilicon 758 -1282 758 -1282 0 3
rlabel polysilicon 765 -1276 765 -1276 0 1
rlabel polysilicon 765 -1282 765 -1282 0 3
rlabel polysilicon 772 -1276 772 -1276 0 1
rlabel polysilicon 772 -1282 772 -1282 0 3
rlabel polysilicon 779 -1276 779 -1276 0 1
rlabel polysilicon 779 -1282 779 -1282 0 3
rlabel polysilicon 786 -1276 786 -1276 0 1
rlabel polysilicon 786 -1282 786 -1282 0 3
rlabel polysilicon 793 -1276 793 -1276 0 1
rlabel polysilicon 793 -1282 793 -1282 0 3
rlabel polysilicon 800 -1276 800 -1276 0 1
rlabel polysilicon 800 -1282 800 -1282 0 3
rlabel polysilicon 807 -1276 807 -1276 0 1
rlabel polysilicon 807 -1282 807 -1282 0 3
rlabel polysilicon 814 -1276 814 -1276 0 1
rlabel polysilicon 814 -1282 814 -1282 0 3
rlabel polysilicon 821 -1276 821 -1276 0 1
rlabel polysilicon 821 -1282 821 -1282 0 3
rlabel polysilicon 828 -1276 828 -1276 0 1
rlabel polysilicon 828 -1282 828 -1282 0 3
rlabel polysilicon 835 -1276 835 -1276 0 1
rlabel polysilicon 835 -1282 835 -1282 0 3
rlabel polysilicon 842 -1276 842 -1276 0 1
rlabel polysilicon 842 -1282 842 -1282 0 3
rlabel polysilicon 849 -1276 849 -1276 0 1
rlabel polysilicon 849 -1282 849 -1282 0 3
rlabel polysilicon 856 -1276 856 -1276 0 1
rlabel polysilicon 856 -1282 856 -1282 0 3
rlabel polysilicon 863 -1276 863 -1276 0 1
rlabel polysilicon 863 -1282 863 -1282 0 3
rlabel polysilicon 870 -1276 870 -1276 0 1
rlabel polysilicon 870 -1282 870 -1282 0 3
rlabel polysilicon 877 -1276 877 -1276 0 1
rlabel polysilicon 877 -1282 877 -1282 0 3
rlabel polysilicon 884 -1276 884 -1276 0 1
rlabel polysilicon 884 -1282 884 -1282 0 3
rlabel polysilicon 891 -1276 891 -1276 0 1
rlabel polysilicon 891 -1282 891 -1282 0 3
rlabel polysilicon 898 -1276 898 -1276 0 1
rlabel polysilicon 898 -1282 898 -1282 0 3
rlabel polysilicon 905 -1276 905 -1276 0 1
rlabel polysilicon 905 -1282 905 -1282 0 3
rlabel polysilicon 912 -1276 912 -1276 0 1
rlabel polysilicon 912 -1282 912 -1282 0 3
rlabel polysilicon 919 -1276 919 -1276 0 1
rlabel polysilicon 919 -1282 919 -1282 0 3
rlabel polysilicon 926 -1276 926 -1276 0 1
rlabel polysilicon 926 -1282 926 -1282 0 3
rlabel polysilicon 933 -1276 933 -1276 0 1
rlabel polysilicon 933 -1282 933 -1282 0 3
rlabel polysilicon 943 -1276 943 -1276 0 2
rlabel polysilicon 943 -1282 943 -1282 0 4
rlabel polysilicon 947 -1276 947 -1276 0 1
rlabel polysilicon 947 -1282 947 -1282 0 3
rlabel polysilicon 954 -1276 954 -1276 0 1
rlabel polysilicon 954 -1282 954 -1282 0 3
rlabel polysilicon 961 -1276 961 -1276 0 1
rlabel polysilicon 961 -1282 961 -1282 0 3
rlabel polysilicon 968 -1276 968 -1276 0 1
rlabel polysilicon 968 -1282 968 -1282 0 3
rlabel polysilicon 975 -1276 975 -1276 0 1
rlabel polysilicon 975 -1282 975 -1282 0 3
rlabel polysilicon 982 -1276 982 -1276 0 1
rlabel polysilicon 982 -1282 982 -1282 0 3
rlabel polysilicon 989 -1276 989 -1276 0 1
rlabel polysilicon 989 -1282 989 -1282 0 3
rlabel polysilicon 996 -1276 996 -1276 0 1
rlabel polysilicon 996 -1282 996 -1282 0 3
rlabel polysilicon 1003 -1276 1003 -1276 0 1
rlabel polysilicon 1003 -1282 1003 -1282 0 3
rlabel polysilicon 1010 -1276 1010 -1276 0 1
rlabel polysilicon 1010 -1282 1010 -1282 0 3
rlabel polysilicon 9 -1361 9 -1361 0 1
rlabel polysilicon 12 -1361 12 -1361 0 2
rlabel polysilicon 9 -1367 9 -1367 0 3
rlabel polysilicon 16 -1361 16 -1361 0 1
rlabel polysilicon 16 -1367 16 -1367 0 3
rlabel polysilicon 23 -1367 23 -1367 0 3
rlabel polysilicon 30 -1361 30 -1361 0 1
rlabel polysilicon 33 -1367 33 -1367 0 4
rlabel polysilicon 37 -1361 37 -1361 0 1
rlabel polysilicon 37 -1367 37 -1367 0 3
rlabel polysilicon 44 -1361 44 -1361 0 1
rlabel polysilicon 44 -1367 44 -1367 0 3
rlabel polysilicon 51 -1361 51 -1361 0 1
rlabel polysilicon 51 -1367 51 -1367 0 3
rlabel polysilicon 61 -1361 61 -1361 0 2
rlabel polysilicon 65 -1361 65 -1361 0 1
rlabel polysilicon 65 -1367 65 -1367 0 3
rlabel polysilicon 72 -1361 72 -1361 0 1
rlabel polysilicon 72 -1367 72 -1367 0 3
rlabel polysilicon 79 -1361 79 -1361 0 1
rlabel polysilicon 79 -1367 79 -1367 0 3
rlabel polysilicon 89 -1361 89 -1361 0 2
rlabel polysilicon 89 -1367 89 -1367 0 4
rlabel polysilicon 93 -1361 93 -1361 0 1
rlabel polysilicon 93 -1367 93 -1367 0 3
rlabel polysilicon 100 -1361 100 -1361 0 1
rlabel polysilicon 100 -1367 100 -1367 0 3
rlabel polysilicon 107 -1361 107 -1361 0 1
rlabel polysilicon 107 -1367 107 -1367 0 3
rlabel polysilicon 114 -1361 114 -1361 0 1
rlabel polysilicon 114 -1367 114 -1367 0 3
rlabel polysilicon 121 -1361 121 -1361 0 1
rlabel polysilicon 124 -1361 124 -1361 0 2
rlabel polysilicon 121 -1367 121 -1367 0 3
rlabel polysilicon 128 -1361 128 -1361 0 1
rlabel polysilicon 128 -1367 128 -1367 0 3
rlabel polysilicon 135 -1361 135 -1361 0 1
rlabel polysilicon 135 -1367 135 -1367 0 3
rlabel polysilicon 142 -1361 142 -1361 0 1
rlabel polysilicon 142 -1367 142 -1367 0 3
rlabel polysilicon 149 -1361 149 -1361 0 1
rlabel polysilicon 149 -1367 149 -1367 0 3
rlabel polysilicon 156 -1361 156 -1361 0 1
rlabel polysilicon 156 -1367 156 -1367 0 3
rlabel polysilicon 159 -1367 159 -1367 0 4
rlabel polysilicon 163 -1361 163 -1361 0 1
rlabel polysilicon 163 -1367 163 -1367 0 3
rlabel polysilicon 170 -1361 170 -1361 0 1
rlabel polysilicon 170 -1367 170 -1367 0 3
rlabel polysilicon 177 -1361 177 -1361 0 1
rlabel polysilicon 177 -1367 177 -1367 0 3
rlabel polysilicon 184 -1361 184 -1361 0 1
rlabel polysilicon 184 -1367 184 -1367 0 3
rlabel polysilicon 191 -1361 191 -1361 0 1
rlabel polysilicon 191 -1367 191 -1367 0 3
rlabel polysilicon 194 -1367 194 -1367 0 4
rlabel polysilicon 198 -1361 198 -1361 0 1
rlabel polysilicon 198 -1367 198 -1367 0 3
rlabel polysilicon 208 -1361 208 -1361 0 2
rlabel polysilicon 205 -1367 205 -1367 0 3
rlabel polysilicon 212 -1361 212 -1361 0 1
rlabel polysilicon 215 -1361 215 -1361 0 2
rlabel polysilicon 219 -1361 219 -1361 0 1
rlabel polysilicon 219 -1367 219 -1367 0 3
rlabel polysilicon 222 -1367 222 -1367 0 4
rlabel polysilicon 226 -1361 226 -1361 0 1
rlabel polysilicon 229 -1361 229 -1361 0 2
rlabel polysilicon 229 -1367 229 -1367 0 4
rlabel polysilicon 233 -1361 233 -1361 0 1
rlabel polysilicon 233 -1367 233 -1367 0 3
rlabel polysilicon 240 -1361 240 -1361 0 1
rlabel polysilicon 240 -1367 240 -1367 0 3
rlabel polysilicon 247 -1361 247 -1361 0 1
rlabel polysilicon 247 -1367 247 -1367 0 3
rlabel polysilicon 254 -1361 254 -1361 0 1
rlabel polysilicon 254 -1367 254 -1367 0 3
rlabel polysilicon 261 -1361 261 -1361 0 1
rlabel polysilicon 261 -1367 261 -1367 0 3
rlabel polysilicon 268 -1361 268 -1361 0 1
rlabel polysilicon 268 -1367 268 -1367 0 3
rlabel polysilicon 275 -1361 275 -1361 0 1
rlabel polysilicon 275 -1367 275 -1367 0 3
rlabel polysilicon 282 -1361 282 -1361 0 1
rlabel polysilicon 282 -1367 282 -1367 0 3
rlabel polysilicon 289 -1361 289 -1361 0 1
rlabel polysilicon 289 -1367 289 -1367 0 3
rlabel polysilicon 296 -1361 296 -1361 0 1
rlabel polysilicon 296 -1367 296 -1367 0 3
rlabel polysilicon 303 -1361 303 -1361 0 1
rlabel polysilicon 303 -1367 303 -1367 0 3
rlabel polysilicon 310 -1361 310 -1361 0 1
rlabel polysilicon 310 -1367 310 -1367 0 3
rlabel polysilicon 317 -1361 317 -1361 0 1
rlabel polysilicon 317 -1367 317 -1367 0 3
rlabel polysilicon 324 -1361 324 -1361 0 1
rlabel polysilicon 324 -1367 324 -1367 0 3
rlabel polysilicon 331 -1361 331 -1361 0 1
rlabel polysilicon 331 -1367 331 -1367 0 3
rlabel polysilicon 334 -1367 334 -1367 0 4
rlabel polysilicon 338 -1361 338 -1361 0 1
rlabel polysilicon 338 -1367 338 -1367 0 3
rlabel polysilicon 345 -1367 345 -1367 0 3
rlabel polysilicon 348 -1367 348 -1367 0 4
rlabel polysilicon 352 -1361 352 -1361 0 1
rlabel polysilicon 352 -1367 352 -1367 0 3
rlabel polysilicon 359 -1361 359 -1361 0 1
rlabel polysilicon 359 -1367 359 -1367 0 3
rlabel polysilicon 366 -1361 366 -1361 0 1
rlabel polysilicon 366 -1367 366 -1367 0 3
rlabel polysilicon 373 -1361 373 -1361 0 1
rlabel polysilicon 373 -1367 373 -1367 0 3
rlabel polysilicon 376 -1367 376 -1367 0 4
rlabel polysilicon 383 -1361 383 -1361 0 2
rlabel polysilicon 380 -1367 380 -1367 0 3
rlabel polysilicon 387 -1361 387 -1361 0 1
rlabel polysilicon 387 -1367 387 -1367 0 3
rlabel polysilicon 394 -1361 394 -1361 0 1
rlabel polysilicon 394 -1367 394 -1367 0 3
rlabel polysilicon 397 -1367 397 -1367 0 4
rlabel polysilicon 401 -1361 401 -1361 0 1
rlabel polysilicon 401 -1367 401 -1367 0 3
rlabel polysilicon 408 -1361 408 -1361 0 1
rlabel polysilicon 408 -1367 408 -1367 0 3
rlabel polysilicon 415 -1361 415 -1361 0 1
rlabel polysilicon 415 -1367 415 -1367 0 3
rlabel polysilicon 422 -1361 422 -1361 0 1
rlabel polysilicon 422 -1367 422 -1367 0 3
rlabel polysilicon 429 -1361 429 -1361 0 1
rlabel polysilicon 432 -1361 432 -1361 0 2
rlabel polysilicon 432 -1367 432 -1367 0 4
rlabel polysilicon 436 -1361 436 -1361 0 1
rlabel polysilicon 436 -1367 436 -1367 0 3
rlabel polysilicon 443 -1361 443 -1361 0 1
rlabel polysilicon 443 -1367 443 -1367 0 3
rlabel polysilicon 450 -1361 450 -1361 0 1
rlabel polysilicon 453 -1361 453 -1361 0 2
rlabel polysilicon 457 -1361 457 -1361 0 1
rlabel polysilicon 457 -1367 457 -1367 0 3
rlabel polysilicon 464 -1361 464 -1361 0 1
rlabel polysilicon 467 -1361 467 -1361 0 2
rlabel polysilicon 464 -1367 464 -1367 0 3
rlabel polysilicon 467 -1367 467 -1367 0 4
rlabel polysilicon 471 -1361 471 -1361 0 1
rlabel polysilicon 471 -1367 471 -1367 0 3
rlabel polysilicon 478 -1361 478 -1361 0 1
rlabel polysilicon 481 -1361 481 -1361 0 2
rlabel polysilicon 478 -1367 478 -1367 0 3
rlabel polysilicon 481 -1367 481 -1367 0 4
rlabel polysilicon 485 -1361 485 -1361 0 1
rlabel polysilicon 488 -1361 488 -1361 0 2
rlabel polysilicon 485 -1367 485 -1367 0 3
rlabel polysilicon 492 -1361 492 -1361 0 1
rlabel polysilicon 492 -1367 492 -1367 0 3
rlabel polysilicon 499 -1361 499 -1361 0 1
rlabel polysilicon 499 -1367 499 -1367 0 3
rlabel polysilicon 506 -1361 506 -1361 0 1
rlabel polysilicon 506 -1367 506 -1367 0 3
rlabel polysilicon 513 -1361 513 -1361 0 1
rlabel polysilicon 513 -1367 513 -1367 0 3
rlabel polysilicon 516 -1367 516 -1367 0 4
rlabel polysilicon 520 -1361 520 -1361 0 1
rlabel polysilicon 520 -1367 520 -1367 0 3
rlabel polysilicon 527 -1361 527 -1361 0 1
rlabel polysilicon 530 -1361 530 -1361 0 2
rlabel polysilicon 527 -1367 527 -1367 0 3
rlabel polysilicon 530 -1367 530 -1367 0 4
rlabel polysilicon 534 -1361 534 -1361 0 1
rlabel polysilicon 534 -1367 534 -1367 0 3
rlabel polysilicon 541 -1361 541 -1361 0 1
rlabel polysilicon 541 -1367 541 -1367 0 3
rlabel polysilicon 548 -1361 548 -1361 0 1
rlabel polysilicon 548 -1367 548 -1367 0 3
rlabel polysilicon 555 -1361 555 -1361 0 1
rlabel polysilicon 555 -1367 555 -1367 0 3
rlabel polysilicon 562 -1361 562 -1361 0 1
rlabel polysilicon 562 -1367 562 -1367 0 3
rlabel polysilicon 569 -1361 569 -1361 0 1
rlabel polysilicon 569 -1367 569 -1367 0 3
rlabel polysilicon 576 -1361 576 -1361 0 1
rlabel polysilicon 579 -1361 579 -1361 0 2
rlabel polysilicon 579 -1367 579 -1367 0 4
rlabel polysilicon 583 -1361 583 -1361 0 1
rlabel polysilicon 583 -1367 583 -1367 0 3
rlabel polysilicon 590 -1361 590 -1361 0 1
rlabel polysilicon 590 -1367 590 -1367 0 3
rlabel polysilicon 597 -1361 597 -1361 0 1
rlabel polysilicon 597 -1367 597 -1367 0 3
rlabel polysilicon 604 -1361 604 -1361 0 1
rlabel polysilicon 604 -1367 604 -1367 0 3
rlabel polysilicon 611 -1361 611 -1361 0 1
rlabel polysilicon 611 -1367 611 -1367 0 3
rlabel polysilicon 618 -1361 618 -1361 0 1
rlabel polysilicon 618 -1367 618 -1367 0 3
rlabel polysilicon 625 -1361 625 -1361 0 1
rlabel polysilicon 625 -1367 625 -1367 0 3
rlabel polysilicon 632 -1361 632 -1361 0 1
rlabel polysilicon 632 -1367 632 -1367 0 3
rlabel polysilicon 639 -1361 639 -1361 0 1
rlabel polysilicon 639 -1367 639 -1367 0 3
rlabel polysilicon 646 -1361 646 -1361 0 1
rlabel polysilicon 646 -1367 646 -1367 0 3
rlabel polysilicon 653 -1361 653 -1361 0 1
rlabel polysilicon 653 -1367 653 -1367 0 3
rlabel polysilicon 660 -1361 660 -1361 0 1
rlabel polysilicon 660 -1367 660 -1367 0 3
rlabel polysilicon 667 -1361 667 -1361 0 1
rlabel polysilicon 667 -1367 667 -1367 0 3
rlabel polysilicon 674 -1361 674 -1361 0 1
rlabel polysilicon 674 -1367 674 -1367 0 3
rlabel polysilicon 681 -1361 681 -1361 0 1
rlabel polysilicon 681 -1367 681 -1367 0 3
rlabel polysilicon 688 -1361 688 -1361 0 1
rlabel polysilicon 688 -1367 688 -1367 0 3
rlabel polysilicon 695 -1361 695 -1361 0 1
rlabel polysilicon 695 -1367 695 -1367 0 3
rlabel polysilicon 702 -1361 702 -1361 0 1
rlabel polysilicon 702 -1367 702 -1367 0 3
rlabel polysilicon 709 -1361 709 -1361 0 1
rlabel polysilicon 709 -1367 709 -1367 0 3
rlabel polysilicon 716 -1361 716 -1361 0 1
rlabel polysilicon 716 -1367 716 -1367 0 3
rlabel polysilicon 723 -1361 723 -1361 0 1
rlabel polysilicon 723 -1367 723 -1367 0 3
rlabel polysilicon 730 -1361 730 -1361 0 1
rlabel polysilicon 730 -1367 730 -1367 0 3
rlabel polysilicon 737 -1361 737 -1361 0 1
rlabel polysilicon 737 -1367 737 -1367 0 3
rlabel polysilicon 744 -1361 744 -1361 0 1
rlabel polysilicon 744 -1367 744 -1367 0 3
rlabel polysilicon 751 -1361 751 -1361 0 1
rlabel polysilicon 751 -1367 751 -1367 0 3
rlabel polysilicon 758 -1361 758 -1361 0 1
rlabel polysilicon 758 -1367 758 -1367 0 3
rlabel polysilicon 765 -1361 765 -1361 0 1
rlabel polysilicon 765 -1367 765 -1367 0 3
rlabel polysilicon 772 -1361 772 -1361 0 1
rlabel polysilicon 772 -1367 772 -1367 0 3
rlabel polysilicon 779 -1361 779 -1361 0 1
rlabel polysilicon 779 -1367 779 -1367 0 3
rlabel polysilicon 786 -1361 786 -1361 0 1
rlabel polysilicon 786 -1367 786 -1367 0 3
rlabel polysilicon 793 -1361 793 -1361 0 1
rlabel polysilicon 793 -1367 793 -1367 0 3
rlabel polysilicon 800 -1361 800 -1361 0 1
rlabel polysilicon 800 -1367 800 -1367 0 3
rlabel polysilicon 807 -1361 807 -1361 0 1
rlabel polysilicon 807 -1367 807 -1367 0 3
rlabel polysilicon 814 -1361 814 -1361 0 1
rlabel polysilicon 814 -1367 814 -1367 0 3
rlabel polysilicon 821 -1361 821 -1361 0 1
rlabel polysilicon 821 -1367 821 -1367 0 3
rlabel polysilicon 828 -1361 828 -1361 0 1
rlabel polysilicon 828 -1367 828 -1367 0 3
rlabel polysilicon 835 -1361 835 -1361 0 1
rlabel polysilicon 835 -1367 835 -1367 0 3
rlabel polysilicon 842 -1361 842 -1361 0 1
rlabel polysilicon 842 -1367 842 -1367 0 3
rlabel polysilicon 849 -1361 849 -1361 0 1
rlabel polysilicon 849 -1367 849 -1367 0 3
rlabel polysilicon 856 -1361 856 -1361 0 1
rlabel polysilicon 856 -1367 856 -1367 0 3
rlabel polysilicon 863 -1361 863 -1361 0 1
rlabel polysilicon 863 -1367 863 -1367 0 3
rlabel polysilicon 870 -1361 870 -1361 0 1
rlabel polysilicon 870 -1367 870 -1367 0 3
rlabel polysilicon 877 -1361 877 -1361 0 1
rlabel polysilicon 877 -1367 877 -1367 0 3
rlabel polysilicon 884 -1361 884 -1361 0 1
rlabel polysilicon 884 -1367 884 -1367 0 3
rlabel polysilicon 891 -1361 891 -1361 0 1
rlabel polysilicon 891 -1367 891 -1367 0 3
rlabel polysilicon 898 -1361 898 -1361 0 1
rlabel polysilicon 898 -1367 898 -1367 0 3
rlabel polysilicon 905 -1361 905 -1361 0 1
rlabel polysilicon 908 -1367 908 -1367 0 4
rlabel polysilicon 912 -1361 912 -1361 0 1
rlabel polysilicon 912 -1367 912 -1367 0 3
rlabel polysilicon 919 -1361 919 -1361 0 1
rlabel polysilicon 940 -1361 940 -1361 0 1
rlabel polysilicon 943 -1361 943 -1361 0 2
rlabel polysilicon 943 -1367 943 -1367 0 4
rlabel polysilicon 954 -1361 954 -1361 0 1
rlabel polysilicon 954 -1367 954 -1367 0 3
rlabel polysilicon 971 -1361 971 -1361 0 2
rlabel polysilicon 971 -1367 971 -1367 0 4
rlabel polysilicon 989 -1361 989 -1361 0 1
rlabel polysilicon 989 -1367 989 -1367 0 3
rlabel polysilicon 2 -1440 2 -1440 0 1
rlabel polysilicon 2 -1446 2 -1446 0 3
rlabel polysilicon 9 -1440 9 -1440 0 1
rlabel polysilicon 16 -1440 16 -1440 0 1
rlabel polysilicon 16 -1446 16 -1446 0 3
rlabel polysilicon 23 -1440 23 -1440 0 1
rlabel polysilicon 23 -1446 23 -1446 0 3
rlabel polysilicon 30 -1440 30 -1440 0 1
rlabel polysilicon 30 -1446 30 -1446 0 3
rlabel polysilicon 37 -1440 37 -1440 0 1
rlabel polysilicon 37 -1446 37 -1446 0 3
rlabel polysilicon 51 -1440 51 -1440 0 1
rlabel polysilicon 51 -1446 51 -1446 0 3
rlabel polysilicon 58 -1440 58 -1440 0 1
rlabel polysilicon 58 -1446 58 -1446 0 3
rlabel polysilicon 65 -1440 65 -1440 0 1
rlabel polysilicon 65 -1446 65 -1446 0 3
rlabel polysilicon 72 -1440 72 -1440 0 1
rlabel polysilicon 72 -1446 72 -1446 0 3
rlabel polysilicon 79 -1440 79 -1440 0 1
rlabel polysilicon 79 -1446 79 -1446 0 3
rlabel polysilicon 86 -1440 86 -1440 0 1
rlabel polysilicon 86 -1446 86 -1446 0 3
rlabel polysilicon 93 -1440 93 -1440 0 1
rlabel polysilicon 93 -1446 93 -1446 0 3
rlabel polysilicon 100 -1440 100 -1440 0 1
rlabel polysilicon 100 -1446 100 -1446 0 3
rlabel polysilicon 107 -1440 107 -1440 0 1
rlabel polysilicon 107 -1446 107 -1446 0 3
rlabel polysilicon 117 -1440 117 -1440 0 2
rlabel polysilicon 117 -1446 117 -1446 0 4
rlabel polysilicon 121 -1440 121 -1440 0 1
rlabel polysilicon 124 -1440 124 -1440 0 2
rlabel polysilicon 128 -1440 128 -1440 0 1
rlabel polysilicon 131 -1446 131 -1446 0 4
rlabel polysilicon 135 -1440 135 -1440 0 1
rlabel polysilicon 135 -1446 135 -1446 0 3
rlabel polysilicon 142 -1446 142 -1446 0 3
rlabel polysilicon 149 -1440 149 -1440 0 1
rlabel polysilicon 149 -1446 149 -1446 0 3
rlabel polysilicon 159 -1440 159 -1440 0 2
rlabel polysilicon 156 -1446 156 -1446 0 3
rlabel polysilicon 166 -1440 166 -1440 0 2
rlabel polysilicon 163 -1446 163 -1446 0 3
rlabel polysilicon 170 -1440 170 -1440 0 1
rlabel polysilicon 170 -1446 170 -1446 0 3
rlabel polysilicon 177 -1440 177 -1440 0 1
rlabel polysilicon 177 -1446 177 -1446 0 3
rlabel polysilicon 187 -1440 187 -1440 0 2
rlabel polysilicon 184 -1446 184 -1446 0 3
rlabel polysilicon 187 -1446 187 -1446 0 4
rlabel polysilicon 191 -1440 191 -1440 0 1
rlabel polysilicon 191 -1446 191 -1446 0 3
rlabel polysilicon 198 -1440 198 -1440 0 1
rlabel polysilicon 198 -1446 198 -1446 0 3
rlabel polysilicon 205 -1440 205 -1440 0 1
rlabel polysilicon 205 -1446 205 -1446 0 3
rlabel polysilicon 212 -1440 212 -1440 0 1
rlabel polysilicon 219 -1440 219 -1440 0 1
rlabel polysilicon 219 -1446 219 -1446 0 3
rlabel polysilicon 226 -1440 226 -1440 0 1
rlabel polysilicon 226 -1446 226 -1446 0 3
rlabel polysilicon 233 -1440 233 -1440 0 1
rlabel polysilicon 233 -1446 233 -1446 0 3
rlabel polysilicon 240 -1440 240 -1440 0 1
rlabel polysilicon 240 -1446 240 -1446 0 3
rlabel polysilicon 247 -1440 247 -1440 0 1
rlabel polysilicon 247 -1446 247 -1446 0 3
rlabel polysilicon 254 -1440 254 -1440 0 1
rlabel polysilicon 254 -1446 254 -1446 0 3
rlabel polysilicon 261 -1440 261 -1440 0 1
rlabel polysilicon 261 -1446 261 -1446 0 3
rlabel polysilicon 268 -1440 268 -1440 0 1
rlabel polysilicon 268 -1446 268 -1446 0 3
rlabel polysilicon 275 -1440 275 -1440 0 1
rlabel polysilicon 275 -1446 275 -1446 0 3
rlabel polysilicon 282 -1440 282 -1440 0 1
rlabel polysilicon 282 -1446 282 -1446 0 3
rlabel polysilicon 289 -1440 289 -1440 0 1
rlabel polysilicon 289 -1446 289 -1446 0 3
rlabel polysilicon 296 -1440 296 -1440 0 1
rlabel polysilicon 296 -1446 296 -1446 0 3
rlabel polysilicon 303 -1440 303 -1440 0 1
rlabel polysilicon 303 -1446 303 -1446 0 3
rlabel polysilicon 310 -1440 310 -1440 0 1
rlabel polysilicon 310 -1446 310 -1446 0 3
rlabel polysilicon 317 -1440 317 -1440 0 1
rlabel polysilicon 317 -1446 317 -1446 0 3
rlabel polysilicon 324 -1446 324 -1446 0 3
rlabel polysilicon 331 -1440 331 -1440 0 1
rlabel polysilicon 331 -1446 331 -1446 0 3
rlabel polysilicon 338 -1440 338 -1440 0 1
rlabel polysilicon 345 -1440 345 -1440 0 1
rlabel polysilicon 345 -1446 345 -1446 0 3
rlabel polysilicon 352 -1440 352 -1440 0 1
rlabel polysilicon 352 -1446 352 -1446 0 3
rlabel polysilicon 355 -1446 355 -1446 0 4
rlabel polysilicon 359 -1440 359 -1440 0 1
rlabel polysilicon 359 -1446 359 -1446 0 3
rlabel polysilicon 366 -1440 366 -1440 0 1
rlabel polysilicon 366 -1446 366 -1446 0 3
rlabel polysilicon 373 -1440 373 -1440 0 1
rlabel polysilicon 376 -1440 376 -1440 0 2
rlabel polysilicon 376 -1446 376 -1446 0 4
rlabel polysilicon 380 -1440 380 -1440 0 1
rlabel polysilicon 380 -1446 380 -1446 0 3
rlabel polysilicon 390 -1440 390 -1440 0 2
rlabel polysilicon 390 -1446 390 -1446 0 4
rlabel polysilicon 394 -1446 394 -1446 0 3
rlabel polysilicon 397 -1446 397 -1446 0 4
rlabel polysilicon 401 -1440 401 -1440 0 1
rlabel polysilicon 401 -1446 401 -1446 0 3
rlabel polysilicon 408 -1440 408 -1440 0 1
rlabel polysilicon 408 -1446 408 -1446 0 3
rlabel polysilicon 415 -1440 415 -1440 0 1
rlabel polysilicon 415 -1446 415 -1446 0 3
rlabel polysilicon 422 -1440 422 -1440 0 1
rlabel polysilicon 422 -1446 422 -1446 0 3
rlabel polysilicon 429 -1446 429 -1446 0 3
rlabel polysilicon 432 -1446 432 -1446 0 4
rlabel polysilicon 436 -1440 436 -1440 0 1
rlabel polysilicon 436 -1446 436 -1446 0 3
rlabel polysilicon 443 -1440 443 -1440 0 1
rlabel polysilicon 443 -1446 443 -1446 0 3
rlabel polysilicon 450 -1440 450 -1440 0 1
rlabel polysilicon 453 -1440 453 -1440 0 2
rlabel polysilicon 460 -1440 460 -1440 0 2
rlabel polysilicon 460 -1446 460 -1446 0 4
rlabel polysilicon 464 -1440 464 -1440 0 1
rlabel polysilicon 467 -1440 467 -1440 0 2
rlabel polysilicon 464 -1446 464 -1446 0 3
rlabel polysilicon 467 -1446 467 -1446 0 4
rlabel polysilicon 471 -1440 471 -1440 0 1
rlabel polysilicon 471 -1446 471 -1446 0 3
rlabel polysilicon 478 -1440 478 -1440 0 1
rlabel polysilicon 478 -1446 478 -1446 0 3
rlabel polysilicon 488 -1440 488 -1440 0 2
rlabel polysilicon 485 -1446 485 -1446 0 3
rlabel polysilicon 492 -1440 492 -1440 0 1
rlabel polysilicon 492 -1446 492 -1446 0 3
rlabel polysilicon 499 -1440 499 -1440 0 1
rlabel polysilicon 499 -1446 499 -1446 0 3
rlabel polysilicon 506 -1440 506 -1440 0 1
rlabel polysilicon 509 -1440 509 -1440 0 2
rlabel polysilicon 506 -1446 506 -1446 0 3
rlabel polysilicon 509 -1446 509 -1446 0 4
rlabel polysilicon 513 -1440 513 -1440 0 1
rlabel polysilicon 513 -1446 513 -1446 0 3
rlabel polysilicon 520 -1440 520 -1440 0 1
rlabel polysilicon 520 -1446 520 -1446 0 3
rlabel polysilicon 527 -1440 527 -1440 0 1
rlabel polysilicon 527 -1446 527 -1446 0 3
rlabel polysilicon 537 -1440 537 -1440 0 2
rlabel polysilicon 537 -1446 537 -1446 0 4
rlabel polysilicon 541 -1440 541 -1440 0 1
rlabel polysilicon 541 -1446 541 -1446 0 3
rlabel polysilicon 551 -1440 551 -1440 0 2
rlabel polysilicon 548 -1446 548 -1446 0 3
rlabel polysilicon 551 -1446 551 -1446 0 4
rlabel polysilicon 555 -1440 555 -1440 0 1
rlabel polysilicon 558 -1440 558 -1440 0 2
rlabel polysilicon 555 -1446 555 -1446 0 3
rlabel polysilicon 562 -1440 562 -1440 0 1
rlabel polysilicon 562 -1446 562 -1446 0 3
rlabel polysilicon 569 -1440 569 -1440 0 1
rlabel polysilicon 569 -1446 569 -1446 0 3
rlabel polysilicon 576 -1440 576 -1440 0 1
rlabel polysilicon 579 -1440 579 -1440 0 2
rlabel polysilicon 583 -1440 583 -1440 0 1
rlabel polysilicon 583 -1446 583 -1446 0 3
rlabel polysilicon 593 -1440 593 -1440 0 2
rlabel polysilicon 590 -1446 590 -1446 0 3
rlabel polysilicon 593 -1446 593 -1446 0 4
rlabel polysilicon 597 -1440 597 -1440 0 1
rlabel polysilicon 597 -1446 597 -1446 0 3
rlabel polysilicon 604 -1440 604 -1440 0 1
rlabel polysilicon 604 -1446 604 -1446 0 3
rlabel polysilicon 607 -1446 607 -1446 0 4
rlabel polysilicon 611 -1440 611 -1440 0 1
rlabel polysilicon 611 -1446 611 -1446 0 3
rlabel polysilicon 618 -1440 618 -1440 0 1
rlabel polysilicon 618 -1446 618 -1446 0 3
rlabel polysilicon 625 -1440 625 -1440 0 1
rlabel polysilicon 625 -1446 625 -1446 0 3
rlabel polysilicon 632 -1440 632 -1440 0 1
rlabel polysilicon 632 -1446 632 -1446 0 3
rlabel polysilicon 635 -1446 635 -1446 0 4
rlabel polysilicon 639 -1440 639 -1440 0 1
rlabel polysilicon 639 -1446 639 -1446 0 3
rlabel polysilicon 646 -1440 646 -1440 0 1
rlabel polysilicon 646 -1446 646 -1446 0 3
rlabel polysilicon 653 -1446 653 -1446 0 3
rlabel polysilicon 656 -1446 656 -1446 0 4
rlabel polysilicon 660 -1440 660 -1440 0 1
rlabel polysilicon 660 -1446 660 -1446 0 3
rlabel polysilicon 667 -1440 667 -1440 0 1
rlabel polysilicon 667 -1446 667 -1446 0 3
rlabel polysilicon 674 -1440 674 -1440 0 1
rlabel polysilicon 674 -1446 674 -1446 0 3
rlabel polysilicon 681 -1440 681 -1440 0 1
rlabel polysilicon 681 -1446 681 -1446 0 3
rlabel polysilicon 688 -1440 688 -1440 0 1
rlabel polysilicon 688 -1446 688 -1446 0 3
rlabel polysilicon 695 -1440 695 -1440 0 1
rlabel polysilicon 695 -1446 695 -1446 0 3
rlabel polysilicon 702 -1440 702 -1440 0 1
rlabel polysilicon 702 -1446 702 -1446 0 3
rlabel polysilicon 712 -1440 712 -1440 0 2
rlabel polysilicon 712 -1446 712 -1446 0 4
rlabel polysilicon 716 -1440 716 -1440 0 1
rlabel polysilicon 716 -1446 716 -1446 0 3
rlabel polysilicon 723 -1440 723 -1440 0 1
rlabel polysilicon 723 -1446 723 -1446 0 3
rlabel polysilicon 730 -1440 730 -1440 0 1
rlabel polysilicon 730 -1446 730 -1446 0 3
rlabel polysilicon 737 -1440 737 -1440 0 1
rlabel polysilicon 737 -1446 737 -1446 0 3
rlabel polysilicon 744 -1440 744 -1440 0 1
rlabel polysilicon 744 -1446 744 -1446 0 3
rlabel polysilicon 751 -1440 751 -1440 0 1
rlabel polysilicon 751 -1446 751 -1446 0 3
rlabel polysilicon 758 -1440 758 -1440 0 1
rlabel polysilicon 758 -1446 758 -1446 0 3
rlabel polysilicon 765 -1440 765 -1440 0 1
rlabel polysilicon 765 -1446 765 -1446 0 3
rlabel polysilicon 772 -1440 772 -1440 0 1
rlabel polysilicon 772 -1446 772 -1446 0 3
rlabel polysilicon 779 -1440 779 -1440 0 1
rlabel polysilicon 779 -1446 779 -1446 0 3
rlabel polysilicon 786 -1440 786 -1440 0 1
rlabel polysilicon 786 -1446 786 -1446 0 3
rlabel polysilicon 793 -1440 793 -1440 0 1
rlabel polysilicon 793 -1446 793 -1446 0 3
rlabel polysilicon 800 -1440 800 -1440 0 1
rlabel polysilicon 800 -1446 800 -1446 0 3
rlabel polysilicon 807 -1440 807 -1440 0 1
rlabel polysilicon 807 -1446 807 -1446 0 3
rlabel polysilicon 814 -1440 814 -1440 0 1
rlabel polysilicon 814 -1446 814 -1446 0 3
rlabel polysilicon 821 -1440 821 -1440 0 1
rlabel polysilicon 821 -1446 821 -1446 0 3
rlabel polysilicon 835 -1440 835 -1440 0 1
rlabel polysilicon 835 -1446 835 -1446 0 3
rlabel polysilicon 842 -1440 842 -1440 0 1
rlabel polysilicon 842 -1446 842 -1446 0 3
rlabel polysilicon 849 -1440 849 -1440 0 1
rlabel polysilicon 849 -1446 849 -1446 0 3
rlabel polysilicon 856 -1440 856 -1440 0 1
rlabel polysilicon 856 -1446 856 -1446 0 3
rlabel polysilicon 863 -1440 863 -1440 0 1
rlabel polysilicon 863 -1446 863 -1446 0 3
rlabel polysilicon 870 -1440 870 -1440 0 1
rlabel polysilicon 870 -1446 870 -1446 0 3
rlabel polysilicon 877 -1440 877 -1440 0 1
rlabel polysilicon 877 -1446 877 -1446 0 3
rlabel polysilicon 884 -1440 884 -1440 0 1
rlabel polysilicon 884 -1446 884 -1446 0 3
rlabel polysilicon 891 -1440 891 -1440 0 1
rlabel polysilicon 891 -1446 891 -1446 0 3
rlabel polysilicon 898 -1440 898 -1440 0 1
rlabel polysilicon 898 -1446 898 -1446 0 3
rlabel polysilicon 905 -1440 905 -1440 0 1
rlabel polysilicon 905 -1446 905 -1446 0 3
rlabel polysilicon 912 -1440 912 -1440 0 1
rlabel polysilicon 912 -1446 912 -1446 0 3
rlabel polysilicon 919 -1440 919 -1440 0 1
rlabel polysilicon 919 -1446 919 -1446 0 3
rlabel polysilicon 926 -1440 926 -1440 0 1
rlabel polysilicon 926 -1446 926 -1446 0 3
rlabel polysilicon 933 -1440 933 -1440 0 1
rlabel polysilicon 933 -1446 933 -1446 0 3
rlabel polysilicon 940 -1440 940 -1440 0 1
rlabel polysilicon 943 -1440 943 -1440 0 2
rlabel polysilicon 947 -1440 947 -1440 0 1
rlabel polysilicon 950 -1446 950 -1446 0 4
rlabel polysilicon 954 -1440 954 -1440 0 1
rlabel polysilicon 954 -1446 954 -1446 0 3
rlabel polysilicon 968 -1440 968 -1440 0 1
rlabel polysilicon 968 -1446 968 -1446 0 3
rlabel polysilicon 982 -1440 982 -1440 0 1
rlabel polysilicon 982 -1446 982 -1446 0 3
rlabel polysilicon 9 -1529 9 -1529 0 1
rlabel polysilicon 9 -1535 9 -1535 0 3
rlabel polysilicon 16 -1529 16 -1529 0 1
rlabel polysilicon 16 -1535 16 -1535 0 3
rlabel polysilicon 23 -1529 23 -1529 0 1
rlabel polysilicon 26 -1535 26 -1535 0 4
rlabel polysilicon 30 -1529 30 -1529 0 1
rlabel polysilicon 30 -1535 30 -1535 0 3
rlabel polysilicon 40 -1529 40 -1529 0 2
rlabel polysilicon 37 -1535 37 -1535 0 3
rlabel polysilicon 40 -1535 40 -1535 0 4
rlabel polysilicon 44 -1529 44 -1529 0 1
rlabel polysilicon 44 -1535 44 -1535 0 3
rlabel polysilicon 51 -1529 51 -1529 0 1
rlabel polysilicon 51 -1535 51 -1535 0 3
rlabel polysilicon 58 -1529 58 -1529 0 1
rlabel polysilicon 58 -1535 58 -1535 0 3
rlabel polysilicon 65 -1529 65 -1529 0 1
rlabel polysilicon 65 -1535 65 -1535 0 3
rlabel polysilicon 72 -1535 72 -1535 0 3
rlabel polysilicon 75 -1535 75 -1535 0 4
rlabel polysilicon 79 -1529 79 -1529 0 1
rlabel polysilicon 79 -1535 79 -1535 0 3
rlabel polysilicon 86 -1529 86 -1529 0 1
rlabel polysilicon 86 -1535 86 -1535 0 3
rlabel polysilicon 93 -1529 93 -1529 0 1
rlabel polysilicon 93 -1535 93 -1535 0 3
rlabel polysilicon 100 -1529 100 -1529 0 1
rlabel polysilicon 100 -1535 100 -1535 0 3
rlabel polysilicon 107 -1529 107 -1529 0 1
rlabel polysilicon 107 -1535 107 -1535 0 3
rlabel polysilicon 114 -1529 114 -1529 0 1
rlabel polysilicon 114 -1535 114 -1535 0 3
rlabel polysilicon 121 -1529 121 -1529 0 1
rlabel polysilicon 121 -1535 121 -1535 0 3
rlabel polysilicon 128 -1529 128 -1529 0 1
rlabel polysilicon 128 -1535 128 -1535 0 3
rlabel polysilicon 135 -1535 135 -1535 0 3
rlabel polysilicon 138 -1535 138 -1535 0 4
rlabel polysilicon 142 -1529 142 -1529 0 1
rlabel polysilicon 142 -1535 142 -1535 0 3
rlabel polysilicon 149 -1529 149 -1529 0 1
rlabel polysilicon 152 -1529 152 -1529 0 2
rlabel polysilicon 149 -1535 149 -1535 0 3
rlabel polysilicon 156 -1529 156 -1529 0 1
rlabel polysilicon 159 -1529 159 -1529 0 2
rlabel polysilicon 156 -1535 156 -1535 0 3
rlabel polysilicon 163 -1529 163 -1529 0 1
rlabel polysilicon 166 -1529 166 -1529 0 2
rlabel polysilicon 163 -1535 163 -1535 0 3
rlabel polysilicon 173 -1529 173 -1529 0 2
rlabel polysilicon 177 -1529 177 -1529 0 1
rlabel polysilicon 180 -1529 180 -1529 0 2
rlabel polysilicon 177 -1535 177 -1535 0 3
rlabel polysilicon 184 -1529 184 -1529 0 1
rlabel polysilicon 187 -1529 187 -1529 0 2
rlabel polysilicon 184 -1535 184 -1535 0 3
rlabel polysilicon 191 -1529 191 -1529 0 1
rlabel polysilicon 194 -1529 194 -1529 0 2
rlabel polysilicon 198 -1529 198 -1529 0 1
rlabel polysilicon 201 -1529 201 -1529 0 2
rlabel polysilicon 201 -1535 201 -1535 0 4
rlabel polysilicon 205 -1529 205 -1529 0 1
rlabel polysilicon 205 -1535 205 -1535 0 3
rlabel polysilicon 215 -1535 215 -1535 0 4
rlabel polysilicon 219 -1529 219 -1529 0 1
rlabel polysilicon 222 -1529 222 -1529 0 2
rlabel polysilicon 226 -1529 226 -1529 0 1
rlabel polysilicon 226 -1535 226 -1535 0 3
rlabel polysilicon 233 -1529 233 -1529 0 1
rlabel polysilicon 233 -1535 233 -1535 0 3
rlabel polysilicon 240 -1529 240 -1529 0 1
rlabel polysilicon 240 -1535 240 -1535 0 3
rlabel polysilicon 247 -1529 247 -1529 0 1
rlabel polysilicon 247 -1535 247 -1535 0 3
rlabel polysilicon 254 -1529 254 -1529 0 1
rlabel polysilicon 254 -1535 254 -1535 0 3
rlabel polysilicon 261 -1529 261 -1529 0 1
rlabel polysilicon 261 -1535 261 -1535 0 3
rlabel polysilicon 268 -1529 268 -1529 0 1
rlabel polysilicon 268 -1535 268 -1535 0 3
rlabel polysilicon 275 -1529 275 -1529 0 1
rlabel polysilicon 275 -1535 275 -1535 0 3
rlabel polysilicon 282 -1529 282 -1529 0 1
rlabel polysilicon 285 -1529 285 -1529 0 2
rlabel polysilicon 282 -1535 282 -1535 0 3
rlabel polysilicon 289 -1529 289 -1529 0 1
rlabel polysilicon 289 -1535 289 -1535 0 3
rlabel polysilicon 296 -1529 296 -1529 0 1
rlabel polysilicon 296 -1535 296 -1535 0 3
rlabel polysilicon 303 -1529 303 -1529 0 1
rlabel polysilicon 306 -1529 306 -1529 0 2
rlabel polysilicon 303 -1535 303 -1535 0 3
rlabel polysilicon 306 -1535 306 -1535 0 4
rlabel polysilicon 310 -1529 310 -1529 0 1
rlabel polysilicon 310 -1535 310 -1535 0 3
rlabel polysilicon 317 -1529 317 -1529 0 1
rlabel polysilicon 317 -1535 317 -1535 0 3
rlabel polysilicon 324 -1529 324 -1529 0 1
rlabel polysilicon 324 -1535 324 -1535 0 3
rlabel polysilicon 331 -1529 331 -1529 0 1
rlabel polysilicon 331 -1535 331 -1535 0 3
rlabel polysilicon 338 -1529 338 -1529 0 1
rlabel polysilicon 338 -1535 338 -1535 0 3
rlabel polysilicon 345 -1529 345 -1529 0 1
rlabel polysilicon 345 -1535 345 -1535 0 3
rlabel polysilicon 352 -1529 352 -1529 0 1
rlabel polysilicon 352 -1535 352 -1535 0 3
rlabel polysilicon 359 -1529 359 -1529 0 1
rlabel polysilicon 362 -1529 362 -1529 0 2
rlabel polysilicon 359 -1535 359 -1535 0 3
rlabel polysilicon 362 -1535 362 -1535 0 4
rlabel polysilicon 366 -1529 366 -1529 0 1
rlabel polysilicon 369 -1529 369 -1529 0 2
rlabel polysilicon 366 -1535 366 -1535 0 3
rlabel polysilicon 369 -1535 369 -1535 0 4
rlabel polysilicon 373 -1529 373 -1529 0 1
rlabel polysilicon 373 -1535 373 -1535 0 3
rlabel polysilicon 380 -1529 380 -1529 0 1
rlabel polysilicon 380 -1535 380 -1535 0 3
rlabel polysilicon 387 -1529 387 -1529 0 1
rlabel polysilicon 394 -1529 394 -1529 0 1
rlabel polysilicon 394 -1535 394 -1535 0 3
rlabel polysilicon 401 -1529 401 -1529 0 1
rlabel polysilicon 401 -1535 401 -1535 0 3
rlabel polysilicon 411 -1529 411 -1529 0 2
rlabel polysilicon 408 -1535 408 -1535 0 3
rlabel polysilicon 411 -1535 411 -1535 0 4
rlabel polysilicon 415 -1529 415 -1529 0 1
rlabel polysilicon 415 -1535 415 -1535 0 3
rlabel polysilicon 422 -1529 422 -1529 0 1
rlabel polysilicon 422 -1535 422 -1535 0 3
rlabel polysilicon 429 -1529 429 -1529 0 1
rlabel polysilicon 432 -1529 432 -1529 0 2
rlabel polysilicon 429 -1535 429 -1535 0 3
rlabel polysilicon 432 -1535 432 -1535 0 4
rlabel polysilicon 436 -1529 436 -1529 0 1
rlabel polysilicon 436 -1535 436 -1535 0 3
rlabel polysilicon 443 -1529 443 -1529 0 1
rlabel polysilicon 446 -1529 446 -1529 0 2
rlabel polysilicon 443 -1535 443 -1535 0 3
rlabel polysilicon 446 -1535 446 -1535 0 4
rlabel polysilicon 450 -1529 450 -1529 0 1
rlabel polysilicon 453 -1529 453 -1529 0 2
rlabel polysilicon 450 -1535 450 -1535 0 3
rlabel polysilicon 453 -1535 453 -1535 0 4
rlabel polysilicon 457 -1529 457 -1529 0 1
rlabel polysilicon 457 -1535 457 -1535 0 3
rlabel polysilicon 464 -1529 464 -1529 0 1
rlabel polysilicon 467 -1529 467 -1529 0 2
rlabel polysilicon 467 -1535 467 -1535 0 4
rlabel polysilicon 471 -1529 471 -1529 0 1
rlabel polysilicon 471 -1535 471 -1535 0 3
rlabel polysilicon 478 -1529 478 -1529 0 1
rlabel polysilicon 478 -1535 478 -1535 0 3
rlabel polysilicon 481 -1535 481 -1535 0 4
rlabel polysilicon 485 -1529 485 -1529 0 1
rlabel polysilicon 485 -1535 485 -1535 0 3
rlabel polysilicon 492 -1529 492 -1529 0 1
rlabel polysilicon 492 -1535 492 -1535 0 3
rlabel polysilicon 499 -1529 499 -1529 0 1
rlabel polysilicon 502 -1529 502 -1529 0 2
rlabel polysilicon 499 -1535 499 -1535 0 3
rlabel polysilicon 506 -1529 506 -1529 0 1
rlabel polysilicon 506 -1535 506 -1535 0 3
rlabel polysilicon 509 -1535 509 -1535 0 4
rlabel polysilicon 513 -1529 513 -1529 0 1
rlabel polysilicon 513 -1535 513 -1535 0 3
rlabel polysilicon 520 -1529 520 -1529 0 1
rlabel polysilicon 520 -1535 520 -1535 0 3
rlabel polysilicon 523 -1535 523 -1535 0 4
rlabel polysilicon 527 -1529 527 -1529 0 1
rlabel polysilicon 527 -1535 527 -1535 0 3
rlabel polysilicon 537 -1529 537 -1529 0 2
rlabel polysilicon 534 -1535 534 -1535 0 3
rlabel polysilicon 537 -1535 537 -1535 0 4
rlabel polysilicon 541 -1529 541 -1529 0 1
rlabel polysilicon 541 -1535 541 -1535 0 3
rlabel polysilicon 548 -1529 548 -1529 0 1
rlabel polysilicon 548 -1535 548 -1535 0 3
rlabel polysilicon 555 -1529 555 -1529 0 1
rlabel polysilicon 558 -1529 558 -1529 0 2
rlabel polysilicon 555 -1535 555 -1535 0 3
rlabel polysilicon 562 -1529 562 -1529 0 1
rlabel polysilicon 562 -1535 562 -1535 0 3
rlabel polysilicon 569 -1529 569 -1529 0 1
rlabel polysilicon 569 -1535 569 -1535 0 3
rlabel polysilicon 576 -1529 576 -1529 0 1
rlabel polysilicon 576 -1535 576 -1535 0 3
rlabel polysilicon 583 -1529 583 -1529 0 1
rlabel polysilicon 583 -1535 583 -1535 0 3
rlabel polysilicon 590 -1529 590 -1529 0 1
rlabel polysilicon 590 -1535 590 -1535 0 3
rlabel polysilicon 597 -1529 597 -1529 0 1
rlabel polysilicon 597 -1535 597 -1535 0 3
rlabel polysilicon 604 -1529 604 -1529 0 1
rlabel polysilicon 604 -1535 604 -1535 0 3
rlabel polysilicon 611 -1529 611 -1529 0 1
rlabel polysilicon 611 -1535 611 -1535 0 3
rlabel polysilicon 618 -1529 618 -1529 0 1
rlabel polysilicon 618 -1535 618 -1535 0 3
rlabel polysilicon 625 -1529 625 -1529 0 1
rlabel polysilicon 625 -1535 625 -1535 0 3
rlabel polysilicon 632 -1529 632 -1529 0 1
rlabel polysilicon 632 -1535 632 -1535 0 3
rlabel polysilicon 639 -1529 639 -1529 0 1
rlabel polysilicon 639 -1535 639 -1535 0 3
rlabel polysilicon 646 -1529 646 -1529 0 1
rlabel polysilicon 646 -1535 646 -1535 0 3
rlabel polysilicon 653 -1529 653 -1529 0 1
rlabel polysilicon 653 -1535 653 -1535 0 3
rlabel polysilicon 660 -1529 660 -1529 0 1
rlabel polysilicon 660 -1535 660 -1535 0 3
rlabel polysilicon 667 -1529 667 -1529 0 1
rlabel polysilicon 667 -1535 667 -1535 0 3
rlabel polysilicon 674 -1529 674 -1529 0 1
rlabel polysilicon 674 -1535 674 -1535 0 3
rlabel polysilicon 681 -1529 681 -1529 0 1
rlabel polysilicon 681 -1535 681 -1535 0 3
rlabel polysilicon 688 -1529 688 -1529 0 1
rlabel polysilicon 688 -1535 688 -1535 0 3
rlabel polysilicon 695 -1529 695 -1529 0 1
rlabel polysilicon 695 -1535 695 -1535 0 3
rlabel polysilicon 702 -1529 702 -1529 0 1
rlabel polysilicon 702 -1535 702 -1535 0 3
rlabel polysilicon 709 -1529 709 -1529 0 1
rlabel polysilicon 709 -1535 709 -1535 0 3
rlabel polysilicon 716 -1529 716 -1529 0 1
rlabel polysilicon 716 -1535 716 -1535 0 3
rlabel polysilicon 723 -1529 723 -1529 0 1
rlabel polysilicon 723 -1535 723 -1535 0 3
rlabel polysilicon 730 -1529 730 -1529 0 1
rlabel polysilicon 730 -1535 730 -1535 0 3
rlabel polysilicon 737 -1529 737 -1529 0 1
rlabel polysilicon 737 -1535 737 -1535 0 3
rlabel polysilicon 744 -1529 744 -1529 0 1
rlabel polysilicon 744 -1535 744 -1535 0 3
rlabel polysilicon 751 -1529 751 -1529 0 1
rlabel polysilicon 751 -1535 751 -1535 0 3
rlabel polysilicon 765 -1529 765 -1529 0 1
rlabel polysilicon 765 -1535 765 -1535 0 3
rlabel polysilicon 772 -1529 772 -1529 0 1
rlabel polysilicon 772 -1535 772 -1535 0 3
rlabel polysilicon 779 -1529 779 -1529 0 1
rlabel polysilicon 779 -1535 779 -1535 0 3
rlabel polysilicon 786 -1529 786 -1529 0 1
rlabel polysilicon 786 -1535 786 -1535 0 3
rlabel polysilicon 793 -1529 793 -1529 0 1
rlabel polysilicon 793 -1535 793 -1535 0 3
rlabel polysilicon 800 -1529 800 -1529 0 1
rlabel polysilicon 800 -1535 800 -1535 0 3
rlabel polysilicon 807 -1529 807 -1529 0 1
rlabel polysilicon 807 -1535 807 -1535 0 3
rlabel polysilicon 814 -1529 814 -1529 0 1
rlabel polysilicon 814 -1535 814 -1535 0 3
rlabel polysilicon 821 -1529 821 -1529 0 1
rlabel polysilicon 821 -1535 821 -1535 0 3
rlabel polysilicon 828 -1529 828 -1529 0 1
rlabel polysilicon 828 -1535 828 -1535 0 3
rlabel polysilicon 835 -1529 835 -1529 0 1
rlabel polysilicon 835 -1535 835 -1535 0 3
rlabel polysilicon 842 -1529 842 -1529 0 1
rlabel polysilicon 842 -1535 842 -1535 0 3
rlabel polysilicon 849 -1529 849 -1529 0 1
rlabel polysilicon 849 -1535 849 -1535 0 3
rlabel polysilicon 856 -1529 856 -1529 0 1
rlabel polysilicon 856 -1535 856 -1535 0 3
rlabel polysilicon 884 -1529 884 -1529 0 1
rlabel polysilicon 887 -1529 887 -1529 0 2
rlabel polysilicon 884 -1535 884 -1535 0 3
rlabel polysilicon 891 -1529 891 -1529 0 1
rlabel polysilicon 891 -1535 891 -1535 0 3
rlabel polysilicon 898 -1529 898 -1529 0 1
rlabel polysilicon 898 -1535 898 -1535 0 3
rlabel polysilicon 905 -1529 905 -1529 0 1
rlabel polysilicon 905 -1535 905 -1535 0 3
rlabel polysilicon 912 -1529 912 -1529 0 1
rlabel polysilicon 912 -1535 912 -1535 0 3
rlabel polysilicon 919 -1529 919 -1529 0 1
rlabel polysilicon 919 -1535 919 -1535 0 3
rlabel polysilicon 933 -1529 933 -1529 0 1
rlabel polysilicon 940 -1529 940 -1529 0 1
rlabel polysilicon 940 -1535 940 -1535 0 3
rlabel polysilicon 954 -1529 954 -1529 0 1
rlabel polysilicon 954 -1535 954 -1535 0 3
rlabel polysilicon 961 -1529 961 -1529 0 1
rlabel polysilicon 982 -1529 982 -1529 0 1
rlabel polysilicon 989 -1529 989 -1529 0 1
rlabel polysilicon 989 -1535 989 -1535 0 3
rlabel polysilicon 9 -1620 9 -1620 0 3
rlabel polysilicon 16 -1614 16 -1614 0 1
rlabel polysilicon 16 -1620 16 -1620 0 3
rlabel polysilicon 23 -1614 23 -1614 0 1
rlabel polysilicon 23 -1620 23 -1620 0 3
rlabel polysilicon 30 -1614 30 -1614 0 1
rlabel polysilicon 30 -1620 30 -1620 0 3
rlabel polysilicon 37 -1614 37 -1614 0 1
rlabel polysilicon 37 -1620 37 -1620 0 3
rlabel polysilicon 44 -1614 44 -1614 0 1
rlabel polysilicon 44 -1620 44 -1620 0 3
rlabel polysilicon 51 -1614 51 -1614 0 1
rlabel polysilicon 51 -1620 51 -1620 0 3
rlabel polysilicon 58 -1614 58 -1614 0 1
rlabel polysilicon 58 -1620 58 -1620 0 3
rlabel polysilicon 65 -1614 65 -1614 0 1
rlabel polysilicon 65 -1620 65 -1620 0 3
rlabel polysilicon 72 -1614 72 -1614 0 1
rlabel polysilicon 72 -1620 72 -1620 0 3
rlabel polysilicon 79 -1614 79 -1614 0 1
rlabel polysilicon 79 -1620 79 -1620 0 3
rlabel polysilicon 86 -1614 86 -1614 0 1
rlabel polysilicon 86 -1620 86 -1620 0 3
rlabel polysilicon 96 -1614 96 -1614 0 2
rlabel polysilicon 93 -1620 93 -1620 0 3
rlabel polysilicon 96 -1620 96 -1620 0 4
rlabel polysilicon 100 -1614 100 -1614 0 1
rlabel polysilicon 100 -1620 100 -1620 0 3
rlabel polysilicon 110 -1614 110 -1614 0 2
rlabel polysilicon 110 -1620 110 -1620 0 4
rlabel polysilicon 121 -1614 121 -1614 0 1
rlabel polysilicon 124 -1620 124 -1620 0 4
rlabel polysilicon 128 -1614 128 -1614 0 1
rlabel polysilicon 128 -1620 128 -1620 0 3
rlabel polysilicon 135 -1614 135 -1614 0 1
rlabel polysilicon 135 -1620 135 -1620 0 3
rlabel polysilicon 142 -1614 142 -1614 0 1
rlabel polysilicon 142 -1620 142 -1620 0 3
rlabel polysilicon 149 -1614 149 -1614 0 1
rlabel polysilicon 149 -1620 149 -1620 0 3
rlabel polysilicon 156 -1614 156 -1614 0 1
rlabel polysilicon 159 -1614 159 -1614 0 2
rlabel polysilicon 156 -1620 156 -1620 0 3
rlabel polysilicon 166 -1614 166 -1614 0 2
rlabel polysilicon 163 -1620 163 -1620 0 3
rlabel polysilicon 166 -1620 166 -1620 0 4
rlabel polysilicon 173 -1614 173 -1614 0 2
rlabel polysilicon 170 -1620 170 -1620 0 3
rlabel polysilicon 173 -1620 173 -1620 0 4
rlabel polysilicon 177 -1614 177 -1614 0 1
rlabel polysilicon 177 -1620 177 -1620 0 3
rlabel polysilicon 184 -1620 184 -1620 0 3
rlabel polysilicon 187 -1620 187 -1620 0 4
rlabel polysilicon 194 -1614 194 -1614 0 2
rlabel polysilicon 191 -1620 191 -1620 0 3
rlabel polysilicon 198 -1614 198 -1614 0 1
rlabel polysilicon 198 -1620 198 -1620 0 3
rlabel polysilicon 205 -1620 205 -1620 0 3
rlabel polysilicon 208 -1620 208 -1620 0 4
rlabel polysilicon 212 -1614 212 -1614 0 1
rlabel polysilicon 212 -1620 212 -1620 0 3
rlabel polysilicon 219 -1614 219 -1614 0 1
rlabel polysilicon 219 -1620 219 -1620 0 3
rlabel polysilicon 226 -1614 226 -1614 0 1
rlabel polysilicon 226 -1620 226 -1620 0 3
rlabel polysilicon 233 -1614 233 -1614 0 1
rlabel polysilicon 233 -1620 233 -1620 0 3
rlabel polysilicon 240 -1614 240 -1614 0 1
rlabel polysilicon 240 -1620 240 -1620 0 3
rlabel polysilicon 247 -1614 247 -1614 0 1
rlabel polysilicon 247 -1620 247 -1620 0 3
rlabel polysilicon 254 -1614 254 -1614 0 1
rlabel polysilicon 254 -1620 254 -1620 0 3
rlabel polysilicon 261 -1614 261 -1614 0 1
rlabel polysilicon 261 -1620 261 -1620 0 3
rlabel polysilicon 268 -1614 268 -1614 0 1
rlabel polysilicon 268 -1620 268 -1620 0 3
rlabel polysilicon 275 -1614 275 -1614 0 1
rlabel polysilicon 275 -1620 275 -1620 0 3
rlabel polysilicon 282 -1614 282 -1614 0 1
rlabel polysilicon 282 -1620 282 -1620 0 3
rlabel polysilicon 289 -1614 289 -1614 0 1
rlabel polysilicon 292 -1614 292 -1614 0 2
rlabel polysilicon 296 -1614 296 -1614 0 1
rlabel polysilicon 296 -1620 296 -1620 0 3
rlabel polysilicon 303 -1614 303 -1614 0 1
rlabel polysilicon 303 -1620 303 -1620 0 3
rlabel polysilicon 310 -1614 310 -1614 0 1
rlabel polysilicon 310 -1620 310 -1620 0 3
rlabel polysilicon 317 -1614 317 -1614 0 1
rlabel polysilicon 317 -1620 317 -1620 0 3
rlabel polysilicon 324 -1614 324 -1614 0 1
rlabel polysilicon 324 -1620 324 -1620 0 3
rlabel polysilicon 331 -1614 331 -1614 0 1
rlabel polysilicon 331 -1620 331 -1620 0 3
rlabel polysilicon 338 -1614 338 -1614 0 1
rlabel polysilicon 341 -1614 341 -1614 0 2
rlabel polysilicon 338 -1620 338 -1620 0 3
rlabel polysilicon 341 -1620 341 -1620 0 4
rlabel polysilicon 345 -1614 345 -1614 0 1
rlabel polysilicon 348 -1614 348 -1614 0 2
rlabel polysilicon 345 -1620 345 -1620 0 3
rlabel polysilicon 348 -1620 348 -1620 0 4
rlabel polysilicon 352 -1614 352 -1614 0 1
rlabel polysilicon 352 -1620 352 -1620 0 3
rlabel polysilicon 359 -1614 359 -1614 0 1
rlabel polysilicon 362 -1614 362 -1614 0 2
rlabel polysilicon 366 -1614 366 -1614 0 1
rlabel polysilicon 366 -1620 366 -1620 0 3
rlabel polysilicon 373 -1614 373 -1614 0 1
rlabel polysilicon 373 -1620 373 -1620 0 3
rlabel polysilicon 383 -1620 383 -1620 0 4
rlabel polysilicon 387 -1620 387 -1620 0 3
rlabel polysilicon 394 -1614 394 -1614 0 1
rlabel polysilicon 394 -1620 394 -1620 0 3
rlabel polysilicon 401 -1614 401 -1614 0 1
rlabel polysilicon 401 -1620 401 -1620 0 3
rlabel polysilicon 408 -1614 408 -1614 0 1
rlabel polysilicon 408 -1620 408 -1620 0 3
rlabel polysilicon 415 -1614 415 -1614 0 1
rlabel polysilicon 415 -1620 415 -1620 0 3
rlabel polysilicon 422 -1620 422 -1620 0 3
rlabel polysilicon 425 -1620 425 -1620 0 4
rlabel polysilicon 429 -1614 429 -1614 0 1
rlabel polysilicon 429 -1620 429 -1620 0 3
rlabel polysilicon 436 -1614 436 -1614 0 1
rlabel polysilicon 436 -1620 436 -1620 0 3
rlabel polysilicon 443 -1614 443 -1614 0 1
rlabel polysilicon 443 -1620 443 -1620 0 3
rlabel polysilicon 453 -1614 453 -1614 0 2
rlabel polysilicon 450 -1620 450 -1620 0 3
rlabel polysilicon 453 -1620 453 -1620 0 4
rlabel polysilicon 457 -1614 457 -1614 0 1
rlabel polysilicon 457 -1620 457 -1620 0 3
rlabel polysilicon 464 -1614 464 -1614 0 1
rlabel polysilicon 464 -1620 464 -1620 0 3
rlabel polysilicon 471 -1614 471 -1614 0 1
rlabel polysilicon 471 -1620 471 -1620 0 3
rlabel polysilicon 478 -1614 478 -1614 0 1
rlabel polysilicon 481 -1614 481 -1614 0 2
rlabel polysilicon 481 -1620 481 -1620 0 4
rlabel polysilicon 485 -1614 485 -1614 0 1
rlabel polysilicon 485 -1620 485 -1620 0 3
rlabel polysilicon 492 -1614 492 -1614 0 1
rlabel polysilicon 492 -1620 492 -1620 0 3
rlabel polysilicon 495 -1620 495 -1620 0 4
rlabel polysilicon 499 -1614 499 -1614 0 1
rlabel polysilicon 499 -1620 499 -1620 0 3
rlabel polysilicon 506 -1614 506 -1614 0 1
rlabel polysilicon 506 -1620 506 -1620 0 3
rlabel polysilicon 513 -1614 513 -1614 0 1
rlabel polysilicon 513 -1620 513 -1620 0 3
rlabel polysilicon 520 -1614 520 -1614 0 1
rlabel polysilicon 523 -1614 523 -1614 0 2
rlabel polysilicon 520 -1620 520 -1620 0 3
rlabel polysilicon 530 -1614 530 -1614 0 2
rlabel polysilicon 527 -1620 527 -1620 0 3
rlabel polysilicon 534 -1614 534 -1614 0 1
rlabel polysilicon 537 -1614 537 -1614 0 2
rlabel polysilicon 534 -1620 534 -1620 0 3
rlabel polysilicon 537 -1620 537 -1620 0 4
rlabel polysilicon 541 -1614 541 -1614 0 1
rlabel polysilicon 541 -1620 541 -1620 0 3
rlabel polysilicon 548 -1614 548 -1614 0 1
rlabel polysilicon 548 -1620 548 -1620 0 3
rlabel polysilicon 555 -1614 555 -1614 0 1
rlabel polysilicon 555 -1620 555 -1620 0 3
rlabel polysilicon 562 -1614 562 -1614 0 1
rlabel polysilicon 565 -1614 565 -1614 0 2
rlabel polysilicon 562 -1620 562 -1620 0 3
rlabel polysilicon 565 -1620 565 -1620 0 4
rlabel polysilicon 569 -1614 569 -1614 0 1
rlabel polysilicon 569 -1620 569 -1620 0 3
rlabel polysilicon 576 -1614 576 -1614 0 1
rlabel polysilicon 576 -1620 576 -1620 0 3
rlabel polysilicon 586 -1614 586 -1614 0 2
rlabel polysilicon 583 -1620 583 -1620 0 3
rlabel polysilicon 586 -1620 586 -1620 0 4
rlabel polysilicon 590 -1614 590 -1614 0 1
rlabel polysilicon 590 -1620 590 -1620 0 3
rlabel polysilicon 597 -1614 597 -1614 0 1
rlabel polysilicon 597 -1620 597 -1620 0 3
rlabel polysilicon 604 -1614 604 -1614 0 1
rlabel polysilicon 604 -1620 604 -1620 0 3
rlabel polysilicon 611 -1614 611 -1614 0 1
rlabel polysilicon 611 -1620 611 -1620 0 3
rlabel polysilicon 625 -1614 625 -1614 0 1
rlabel polysilicon 625 -1620 625 -1620 0 3
rlabel polysilicon 632 -1614 632 -1614 0 1
rlabel polysilicon 632 -1620 632 -1620 0 3
rlabel polysilicon 639 -1614 639 -1614 0 1
rlabel polysilicon 639 -1620 639 -1620 0 3
rlabel polysilicon 646 -1614 646 -1614 0 1
rlabel polysilicon 646 -1620 646 -1620 0 3
rlabel polysilicon 653 -1614 653 -1614 0 1
rlabel polysilicon 653 -1620 653 -1620 0 3
rlabel polysilicon 660 -1614 660 -1614 0 1
rlabel polysilicon 660 -1620 660 -1620 0 3
rlabel polysilicon 667 -1614 667 -1614 0 1
rlabel polysilicon 667 -1620 667 -1620 0 3
rlabel polysilicon 674 -1614 674 -1614 0 1
rlabel polysilicon 674 -1620 674 -1620 0 3
rlabel polysilicon 681 -1614 681 -1614 0 1
rlabel polysilicon 681 -1620 681 -1620 0 3
rlabel polysilicon 688 -1614 688 -1614 0 1
rlabel polysilicon 688 -1620 688 -1620 0 3
rlabel polysilicon 695 -1614 695 -1614 0 1
rlabel polysilicon 695 -1620 695 -1620 0 3
rlabel polysilicon 702 -1614 702 -1614 0 1
rlabel polysilicon 705 -1614 705 -1614 0 2
rlabel polysilicon 702 -1620 702 -1620 0 3
rlabel polysilicon 705 -1620 705 -1620 0 4
rlabel polysilicon 709 -1614 709 -1614 0 1
rlabel polysilicon 709 -1620 709 -1620 0 3
rlabel polysilicon 716 -1614 716 -1614 0 1
rlabel polysilicon 716 -1620 716 -1620 0 3
rlabel polysilicon 723 -1614 723 -1614 0 1
rlabel polysilicon 723 -1620 723 -1620 0 3
rlabel polysilicon 733 -1614 733 -1614 0 2
rlabel polysilicon 730 -1620 730 -1620 0 3
rlabel polysilicon 733 -1620 733 -1620 0 4
rlabel polysilicon 744 -1614 744 -1614 0 1
rlabel polysilicon 744 -1620 744 -1620 0 3
rlabel polysilicon 751 -1614 751 -1614 0 1
rlabel polysilicon 751 -1620 751 -1620 0 3
rlabel polysilicon 758 -1614 758 -1614 0 1
rlabel polysilicon 758 -1620 758 -1620 0 3
rlabel polysilicon 765 -1614 765 -1614 0 1
rlabel polysilicon 765 -1620 765 -1620 0 3
rlabel polysilicon 786 -1614 786 -1614 0 1
rlabel polysilicon 786 -1620 786 -1620 0 3
rlabel polysilicon 793 -1614 793 -1614 0 1
rlabel polysilicon 793 -1620 793 -1620 0 3
rlabel polysilicon 800 -1614 800 -1614 0 1
rlabel polysilicon 800 -1620 800 -1620 0 3
rlabel polysilicon 814 -1614 814 -1614 0 1
rlabel polysilicon 814 -1620 814 -1620 0 3
rlabel polysilicon 828 -1614 828 -1614 0 1
rlabel polysilicon 828 -1620 828 -1620 0 3
rlabel polysilicon 842 -1614 842 -1614 0 1
rlabel polysilicon 842 -1620 842 -1620 0 3
rlabel polysilicon 849 -1614 849 -1614 0 1
rlabel polysilicon 852 -1614 852 -1614 0 2
rlabel polysilicon 849 -1620 849 -1620 0 3
rlabel polysilicon 856 -1614 856 -1614 0 1
rlabel polysilicon 856 -1620 856 -1620 0 3
rlabel polysilicon 870 -1614 870 -1614 0 1
rlabel polysilicon 870 -1620 870 -1620 0 3
rlabel polysilicon 880 -1614 880 -1614 0 2
rlabel polysilicon 877 -1620 877 -1620 0 3
rlabel polysilicon 898 -1614 898 -1614 0 1
rlabel polysilicon 898 -1620 898 -1620 0 3
rlabel polysilicon 915 -1614 915 -1614 0 2
rlabel polysilicon 919 -1614 919 -1614 0 1
rlabel polysilicon 919 -1620 919 -1620 0 3
rlabel polysilicon 926 -1614 926 -1614 0 1
rlabel polysilicon 926 -1620 926 -1620 0 3
rlabel polysilicon 940 -1614 940 -1614 0 1
rlabel polysilicon 940 -1620 940 -1620 0 3
rlabel polysilicon 943 -1620 943 -1620 0 4
rlabel polysilicon 947 -1614 947 -1614 0 1
rlabel polysilicon 947 -1620 947 -1620 0 3
rlabel polysilicon 954 -1614 954 -1614 0 1
rlabel polysilicon 954 -1620 954 -1620 0 3
rlabel polysilicon 968 -1614 968 -1614 0 1
rlabel polysilicon 971 -1614 971 -1614 0 2
rlabel polysilicon 975 -1614 975 -1614 0 1
rlabel polysilicon 975 -1620 975 -1620 0 3
rlabel polysilicon 982 -1614 982 -1614 0 1
rlabel polysilicon 982 -1620 982 -1620 0 3
rlabel polysilicon 9 -1707 9 -1707 0 1
rlabel polysilicon 9 -1713 9 -1713 0 3
rlabel polysilicon 16 -1707 16 -1707 0 1
rlabel polysilicon 16 -1713 16 -1713 0 3
rlabel polysilicon 23 -1707 23 -1707 0 1
rlabel polysilicon 23 -1713 23 -1713 0 3
rlabel polysilicon 30 -1707 30 -1707 0 1
rlabel polysilicon 30 -1713 30 -1713 0 3
rlabel polysilicon 37 -1707 37 -1707 0 1
rlabel polysilicon 37 -1713 37 -1713 0 3
rlabel polysilicon 44 -1707 44 -1707 0 1
rlabel polysilicon 44 -1713 44 -1713 0 3
rlabel polysilicon 51 -1707 51 -1707 0 1
rlabel polysilicon 51 -1713 51 -1713 0 3
rlabel polysilicon 58 -1707 58 -1707 0 1
rlabel polysilicon 61 -1707 61 -1707 0 2
rlabel polysilicon 58 -1713 58 -1713 0 3
rlabel polysilicon 65 -1707 65 -1707 0 1
rlabel polysilicon 65 -1713 65 -1713 0 3
rlabel polysilicon 75 -1713 75 -1713 0 4
rlabel polysilicon 79 -1707 79 -1707 0 1
rlabel polysilicon 79 -1713 79 -1713 0 3
rlabel polysilicon 86 -1707 86 -1707 0 1
rlabel polysilicon 86 -1713 86 -1713 0 3
rlabel polysilicon 93 -1707 93 -1707 0 1
rlabel polysilicon 93 -1713 93 -1713 0 3
rlabel polysilicon 103 -1707 103 -1707 0 2
rlabel polysilicon 103 -1713 103 -1713 0 4
rlabel polysilicon 107 -1707 107 -1707 0 1
rlabel polysilicon 107 -1713 107 -1713 0 3
rlabel polysilicon 117 -1707 117 -1707 0 2
rlabel polysilicon 117 -1713 117 -1713 0 4
rlabel polysilicon 121 -1707 121 -1707 0 1
rlabel polysilicon 121 -1713 121 -1713 0 3
rlabel polysilicon 128 -1707 128 -1707 0 1
rlabel polysilicon 128 -1713 128 -1713 0 3
rlabel polysilicon 135 -1707 135 -1707 0 1
rlabel polysilicon 135 -1713 135 -1713 0 3
rlabel polysilicon 142 -1707 142 -1707 0 1
rlabel polysilicon 145 -1707 145 -1707 0 2
rlabel polysilicon 149 -1707 149 -1707 0 1
rlabel polysilicon 152 -1707 152 -1707 0 2
rlabel polysilicon 156 -1707 156 -1707 0 1
rlabel polysilicon 156 -1713 156 -1713 0 3
rlabel polysilicon 163 -1707 163 -1707 0 1
rlabel polysilicon 163 -1713 163 -1713 0 3
rlabel polysilicon 173 -1707 173 -1707 0 2
rlabel polysilicon 170 -1713 170 -1713 0 3
rlabel polysilicon 180 -1707 180 -1707 0 2
rlabel polysilicon 184 -1707 184 -1707 0 1
rlabel polysilicon 184 -1713 184 -1713 0 3
rlabel polysilicon 191 -1707 191 -1707 0 1
rlabel polysilicon 191 -1713 191 -1713 0 3
rlabel polysilicon 198 -1707 198 -1707 0 1
rlabel polysilicon 198 -1713 198 -1713 0 3
rlabel polysilicon 205 -1707 205 -1707 0 1
rlabel polysilicon 208 -1707 208 -1707 0 2
rlabel polysilicon 212 -1707 212 -1707 0 1
rlabel polysilicon 212 -1713 212 -1713 0 3
rlabel polysilicon 219 -1707 219 -1707 0 1
rlabel polysilicon 219 -1713 219 -1713 0 3
rlabel polysilicon 226 -1707 226 -1707 0 1
rlabel polysilicon 226 -1713 226 -1713 0 3
rlabel polysilicon 233 -1713 233 -1713 0 3
rlabel polysilicon 236 -1713 236 -1713 0 4
rlabel polysilicon 240 -1707 240 -1707 0 1
rlabel polysilicon 240 -1713 240 -1713 0 3
rlabel polysilicon 247 -1707 247 -1707 0 1
rlabel polysilicon 247 -1713 247 -1713 0 3
rlabel polysilicon 254 -1707 254 -1707 0 1
rlabel polysilicon 254 -1713 254 -1713 0 3
rlabel polysilicon 261 -1707 261 -1707 0 1
rlabel polysilicon 261 -1713 261 -1713 0 3
rlabel polysilicon 268 -1707 268 -1707 0 1
rlabel polysilicon 268 -1713 268 -1713 0 3
rlabel polysilicon 275 -1707 275 -1707 0 1
rlabel polysilicon 275 -1713 275 -1713 0 3
rlabel polysilicon 282 -1707 282 -1707 0 1
rlabel polysilicon 282 -1713 282 -1713 0 3
rlabel polysilicon 289 -1707 289 -1707 0 1
rlabel polysilicon 289 -1713 289 -1713 0 3
rlabel polysilicon 296 -1707 296 -1707 0 1
rlabel polysilicon 299 -1707 299 -1707 0 2
rlabel polysilicon 296 -1713 296 -1713 0 3
rlabel polysilicon 299 -1713 299 -1713 0 4
rlabel polysilicon 303 -1707 303 -1707 0 1
rlabel polysilicon 303 -1713 303 -1713 0 3
rlabel polysilicon 310 -1707 310 -1707 0 1
rlabel polysilicon 310 -1713 310 -1713 0 3
rlabel polysilicon 317 -1707 317 -1707 0 1
rlabel polysilicon 317 -1713 317 -1713 0 3
rlabel polysilicon 324 -1707 324 -1707 0 1
rlabel polysilicon 324 -1713 324 -1713 0 3
rlabel polysilicon 331 -1707 331 -1707 0 1
rlabel polysilicon 331 -1713 331 -1713 0 3
rlabel polysilicon 334 -1713 334 -1713 0 4
rlabel polysilicon 341 -1707 341 -1707 0 2
rlabel polysilicon 338 -1713 338 -1713 0 3
rlabel polysilicon 341 -1713 341 -1713 0 4
rlabel polysilicon 345 -1707 345 -1707 0 1
rlabel polysilicon 345 -1713 345 -1713 0 3
rlabel polysilicon 352 -1707 352 -1707 0 1
rlabel polysilicon 352 -1713 352 -1713 0 3
rlabel polysilicon 359 -1707 359 -1707 0 1
rlabel polysilicon 359 -1713 359 -1713 0 3
rlabel polysilicon 366 -1707 366 -1707 0 1
rlabel polysilicon 366 -1713 366 -1713 0 3
rlabel polysilicon 373 -1713 373 -1713 0 3
rlabel polysilicon 376 -1713 376 -1713 0 4
rlabel polysilicon 380 -1707 380 -1707 0 1
rlabel polysilicon 380 -1713 380 -1713 0 3
rlabel polysilicon 387 -1707 387 -1707 0 1
rlabel polysilicon 390 -1707 390 -1707 0 2
rlabel polysilicon 387 -1713 387 -1713 0 3
rlabel polysilicon 397 -1707 397 -1707 0 2
rlabel polysilicon 394 -1713 394 -1713 0 3
rlabel polysilicon 397 -1713 397 -1713 0 4
rlabel polysilicon 401 -1707 401 -1707 0 1
rlabel polysilicon 404 -1707 404 -1707 0 2
rlabel polysilicon 401 -1713 401 -1713 0 3
rlabel polysilicon 408 -1707 408 -1707 0 1
rlabel polysilicon 408 -1713 408 -1713 0 3
rlabel polysilicon 415 -1707 415 -1707 0 1
rlabel polysilicon 415 -1713 415 -1713 0 3
rlabel polysilicon 422 -1707 422 -1707 0 1
rlabel polysilicon 422 -1713 422 -1713 0 3
rlabel polysilicon 429 -1707 429 -1707 0 1
rlabel polysilicon 429 -1713 429 -1713 0 3
rlabel polysilicon 436 -1707 436 -1707 0 1
rlabel polysilicon 439 -1707 439 -1707 0 2
rlabel polysilicon 439 -1713 439 -1713 0 4
rlabel polysilicon 443 -1707 443 -1707 0 1
rlabel polysilicon 443 -1713 443 -1713 0 3
rlabel polysilicon 450 -1707 450 -1707 0 1
rlabel polysilicon 450 -1713 450 -1713 0 3
rlabel polysilicon 453 -1713 453 -1713 0 4
rlabel polysilicon 457 -1707 457 -1707 0 1
rlabel polysilicon 457 -1713 457 -1713 0 3
rlabel polysilicon 464 -1707 464 -1707 0 1
rlabel polysilicon 464 -1713 464 -1713 0 3
rlabel polysilicon 467 -1713 467 -1713 0 4
rlabel polysilicon 471 -1707 471 -1707 0 1
rlabel polysilicon 471 -1713 471 -1713 0 3
rlabel polysilicon 478 -1707 478 -1707 0 1
rlabel polysilicon 478 -1713 478 -1713 0 3
rlabel polysilicon 488 -1707 488 -1707 0 2
rlabel polysilicon 485 -1713 485 -1713 0 3
rlabel polysilicon 488 -1713 488 -1713 0 4
rlabel polysilicon 492 -1707 492 -1707 0 1
rlabel polysilicon 492 -1713 492 -1713 0 3
rlabel polysilicon 499 -1707 499 -1707 0 1
rlabel polysilicon 499 -1713 499 -1713 0 3
rlabel polysilicon 509 -1707 509 -1707 0 2
rlabel polysilicon 509 -1713 509 -1713 0 4
rlabel polysilicon 513 -1707 513 -1707 0 1
rlabel polysilicon 513 -1713 513 -1713 0 3
rlabel polysilicon 520 -1707 520 -1707 0 1
rlabel polysilicon 520 -1713 520 -1713 0 3
rlabel polysilicon 527 -1707 527 -1707 0 1
rlabel polysilicon 527 -1713 527 -1713 0 3
rlabel polysilicon 534 -1707 534 -1707 0 1
rlabel polysilicon 534 -1713 534 -1713 0 3
rlabel polysilicon 541 -1707 541 -1707 0 1
rlabel polysilicon 544 -1707 544 -1707 0 2
rlabel polysilicon 541 -1713 541 -1713 0 3
rlabel polysilicon 548 -1707 548 -1707 0 1
rlabel polysilicon 548 -1713 548 -1713 0 3
rlabel polysilicon 555 -1707 555 -1707 0 1
rlabel polysilicon 555 -1713 555 -1713 0 3
rlabel polysilicon 562 -1707 562 -1707 0 1
rlabel polysilicon 562 -1713 562 -1713 0 3
rlabel polysilicon 569 -1707 569 -1707 0 1
rlabel polysilicon 572 -1707 572 -1707 0 2
rlabel polysilicon 572 -1713 572 -1713 0 4
rlabel polysilicon 576 -1707 576 -1707 0 1
rlabel polysilicon 576 -1713 576 -1713 0 3
rlabel polysilicon 583 -1707 583 -1707 0 1
rlabel polysilicon 583 -1713 583 -1713 0 3
rlabel polysilicon 590 -1707 590 -1707 0 1
rlabel polysilicon 590 -1713 590 -1713 0 3
rlabel polysilicon 597 -1707 597 -1707 0 1
rlabel polysilicon 597 -1713 597 -1713 0 3
rlabel polysilicon 604 -1707 604 -1707 0 1
rlabel polysilicon 604 -1713 604 -1713 0 3
rlabel polysilicon 611 -1707 611 -1707 0 1
rlabel polysilicon 611 -1713 611 -1713 0 3
rlabel polysilicon 618 -1707 618 -1707 0 1
rlabel polysilicon 618 -1713 618 -1713 0 3
rlabel polysilicon 625 -1707 625 -1707 0 1
rlabel polysilicon 625 -1713 625 -1713 0 3
rlabel polysilicon 632 -1707 632 -1707 0 1
rlabel polysilicon 632 -1713 632 -1713 0 3
rlabel polysilicon 639 -1707 639 -1707 0 1
rlabel polysilicon 639 -1713 639 -1713 0 3
rlabel polysilicon 646 -1707 646 -1707 0 1
rlabel polysilicon 646 -1713 646 -1713 0 3
rlabel polysilicon 653 -1707 653 -1707 0 1
rlabel polysilicon 653 -1713 653 -1713 0 3
rlabel polysilicon 660 -1707 660 -1707 0 1
rlabel polysilicon 660 -1713 660 -1713 0 3
rlabel polysilicon 667 -1707 667 -1707 0 1
rlabel polysilicon 667 -1713 667 -1713 0 3
rlabel polysilicon 674 -1707 674 -1707 0 1
rlabel polysilicon 674 -1713 674 -1713 0 3
rlabel polysilicon 681 -1707 681 -1707 0 1
rlabel polysilicon 681 -1713 681 -1713 0 3
rlabel polysilicon 688 -1707 688 -1707 0 1
rlabel polysilicon 688 -1713 688 -1713 0 3
rlabel polysilicon 695 -1707 695 -1707 0 1
rlabel polysilicon 695 -1713 695 -1713 0 3
rlabel polysilicon 702 -1707 702 -1707 0 1
rlabel polysilicon 702 -1713 702 -1713 0 3
rlabel polysilicon 712 -1707 712 -1707 0 2
rlabel polysilicon 716 -1707 716 -1707 0 1
rlabel polysilicon 716 -1713 716 -1713 0 3
rlabel polysilicon 723 -1707 723 -1707 0 1
rlabel polysilicon 723 -1713 723 -1713 0 3
rlabel polysilicon 730 -1707 730 -1707 0 1
rlabel polysilicon 730 -1713 730 -1713 0 3
rlabel polysilicon 737 -1707 737 -1707 0 1
rlabel polysilicon 737 -1713 737 -1713 0 3
rlabel polysilicon 744 -1707 744 -1707 0 1
rlabel polysilicon 744 -1713 744 -1713 0 3
rlabel polysilicon 751 -1707 751 -1707 0 1
rlabel polysilicon 751 -1713 751 -1713 0 3
rlabel polysilicon 758 -1707 758 -1707 0 1
rlabel polysilicon 758 -1713 758 -1713 0 3
rlabel polysilicon 765 -1707 765 -1707 0 1
rlabel polysilicon 765 -1713 765 -1713 0 3
rlabel polysilicon 772 -1707 772 -1707 0 1
rlabel polysilicon 772 -1713 772 -1713 0 3
rlabel polysilicon 779 -1707 779 -1707 0 1
rlabel polysilicon 779 -1713 779 -1713 0 3
rlabel polysilicon 786 -1707 786 -1707 0 1
rlabel polysilicon 786 -1713 786 -1713 0 3
rlabel polysilicon 800 -1707 800 -1707 0 1
rlabel polysilicon 800 -1713 800 -1713 0 3
rlabel polysilicon 814 -1707 814 -1707 0 1
rlabel polysilicon 814 -1713 814 -1713 0 3
rlabel polysilicon 821 -1707 821 -1707 0 1
rlabel polysilicon 821 -1713 821 -1713 0 3
rlabel polysilicon 828 -1707 828 -1707 0 1
rlabel polysilicon 828 -1713 828 -1713 0 3
rlabel polysilicon 835 -1707 835 -1707 0 1
rlabel polysilicon 835 -1713 835 -1713 0 3
rlabel polysilicon 842 -1707 842 -1707 0 1
rlabel polysilicon 842 -1713 842 -1713 0 3
rlabel polysilicon 863 -1707 863 -1707 0 1
rlabel polysilicon 863 -1713 863 -1713 0 3
rlabel polysilicon 870 -1707 870 -1707 0 1
rlabel polysilicon 870 -1713 870 -1713 0 3
rlabel polysilicon 887 -1707 887 -1707 0 2
rlabel polysilicon 887 -1713 887 -1713 0 4
rlabel polysilicon 894 -1707 894 -1707 0 2
rlabel polysilicon 912 -1707 912 -1707 0 1
rlabel polysilicon 912 -1713 912 -1713 0 3
rlabel polysilicon 926 -1707 926 -1707 0 1
rlabel polysilicon 926 -1713 926 -1713 0 3
rlabel polysilicon 940 -1713 940 -1713 0 3
rlabel polysilicon 961 -1707 961 -1707 0 1
rlabel polysilicon 961 -1713 961 -1713 0 3
rlabel polysilicon 971 -1707 971 -1707 0 2
rlabel polysilicon 975 -1707 975 -1707 0 1
rlabel polysilicon 978 -1713 978 -1713 0 4
rlabel polysilicon 9 -1802 9 -1802 0 1
rlabel polysilicon 9 -1808 9 -1808 0 3
rlabel polysilicon 12 -1808 12 -1808 0 4
rlabel polysilicon 16 -1802 16 -1802 0 1
rlabel polysilicon 16 -1808 16 -1808 0 3
rlabel polysilicon 23 -1802 23 -1802 0 1
rlabel polysilicon 23 -1808 23 -1808 0 3
rlabel polysilicon 30 -1802 30 -1802 0 1
rlabel polysilicon 30 -1808 30 -1808 0 3
rlabel polysilicon 37 -1802 37 -1802 0 1
rlabel polysilicon 40 -1808 40 -1808 0 4
rlabel polysilicon 44 -1802 44 -1802 0 1
rlabel polysilicon 44 -1808 44 -1808 0 3
rlabel polysilicon 51 -1802 51 -1802 0 1
rlabel polysilicon 58 -1802 58 -1802 0 1
rlabel polysilicon 58 -1808 58 -1808 0 3
rlabel polysilicon 65 -1802 65 -1802 0 1
rlabel polysilicon 65 -1808 65 -1808 0 3
rlabel polysilicon 72 -1802 72 -1802 0 1
rlabel polysilicon 72 -1808 72 -1808 0 3
rlabel polysilicon 82 -1802 82 -1802 0 2
rlabel polysilicon 82 -1808 82 -1808 0 4
rlabel polysilicon 86 -1802 86 -1802 0 1
rlabel polysilicon 89 -1808 89 -1808 0 4
rlabel polysilicon 93 -1802 93 -1802 0 1
rlabel polysilicon 93 -1808 93 -1808 0 3
rlabel polysilicon 103 -1802 103 -1802 0 2
rlabel polysilicon 103 -1808 103 -1808 0 4
rlabel polysilicon 107 -1802 107 -1802 0 1
rlabel polysilicon 107 -1808 107 -1808 0 3
rlabel polysilicon 114 -1802 114 -1802 0 1
rlabel polysilicon 117 -1802 117 -1802 0 2
rlabel polysilicon 114 -1808 114 -1808 0 3
rlabel polysilicon 124 -1802 124 -1802 0 2
rlabel polysilicon 121 -1808 121 -1808 0 3
rlabel polysilicon 124 -1808 124 -1808 0 4
rlabel polysilicon 128 -1808 128 -1808 0 3
rlabel polysilicon 135 -1808 135 -1808 0 3
rlabel polysilicon 138 -1808 138 -1808 0 4
rlabel polysilicon 142 -1802 142 -1802 0 1
rlabel polysilicon 142 -1808 142 -1808 0 3
rlabel polysilicon 149 -1802 149 -1802 0 1
rlabel polysilicon 149 -1808 149 -1808 0 3
rlabel polysilicon 156 -1802 156 -1802 0 1
rlabel polysilicon 159 -1802 159 -1802 0 2
rlabel polysilicon 166 -1802 166 -1802 0 2
rlabel polysilicon 163 -1808 163 -1808 0 3
rlabel polysilicon 166 -1808 166 -1808 0 4
rlabel polysilicon 170 -1802 170 -1802 0 1
rlabel polysilicon 173 -1802 173 -1802 0 2
rlabel polysilicon 170 -1808 170 -1808 0 3
rlabel polysilicon 173 -1808 173 -1808 0 4
rlabel polysilicon 180 -1802 180 -1802 0 2
rlabel polysilicon 180 -1808 180 -1808 0 4
rlabel polysilicon 184 -1802 184 -1802 0 1
rlabel polysilicon 187 -1802 187 -1802 0 2
rlabel polysilicon 187 -1808 187 -1808 0 4
rlabel polysilicon 191 -1802 191 -1802 0 1
rlabel polysilicon 191 -1808 191 -1808 0 3
rlabel polysilicon 198 -1802 198 -1802 0 1
rlabel polysilicon 198 -1808 198 -1808 0 3
rlabel polysilicon 205 -1802 205 -1802 0 1
rlabel polysilicon 205 -1808 205 -1808 0 3
rlabel polysilicon 212 -1802 212 -1802 0 1
rlabel polysilicon 215 -1808 215 -1808 0 4
rlabel polysilicon 219 -1802 219 -1802 0 1
rlabel polysilicon 222 -1802 222 -1802 0 2
rlabel polysilicon 219 -1808 219 -1808 0 3
rlabel polysilicon 222 -1808 222 -1808 0 4
rlabel polysilicon 226 -1802 226 -1802 0 1
rlabel polysilicon 226 -1808 226 -1808 0 3
rlabel polysilicon 233 -1802 233 -1802 0 1
rlabel polysilicon 233 -1808 233 -1808 0 3
rlabel polysilicon 240 -1802 240 -1802 0 1
rlabel polysilicon 240 -1808 240 -1808 0 3
rlabel polysilicon 247 -1802 247 -1802 0 1
rlabel polysilicon 247 -1808 247 -1808 0 3
rlabel polysilicon 254 -1802 254 -1802 0 1
rlabel polysilicon 254 -1808 254 -1808 0 3
rlabel polysilicon 261 -1802 261 -1802 0 1
rlabel polysilicon 261 -1808 261 -1808 0 3
rlabel polysilicon 271 -1802 271 -1802 0 2
rlabel polysilicon 268 -1808 268 -1808 0 3
rlabel polysilicon 275 -1802 275 -1802 0 1
rlabel polysilicon 275 -1808 275 -1808 0 3
rlabel polysilicon 282 -1802 282 -1802 0 1
rlabel polysilicon 282 -1808 282 -1808 0 3
rlabel polysilicon 289 -1802 289 -1802 0 1
rlabel polysilicon 289 -1808 289 -1808 0 3
rlabel polysilicon 296 -1802 296 -1802 0 1
rlabel polysilicon 296 -1808 296 -1808 0 3
rlabel polysilicon 303 -1802 303 -1802 0 1
rlabel polysilicon 303 -1808 303 -1808 0 3
rlabel polysilicon 310 -1802 310 -1802 0 1
rlabel polysilicon 310 -1808 310 -1808 0 3
rlabel polysilicon 320 -1802 320 -1802 0 2
rlabel polysilicon 317 -1808 317 -1808 0 3
rlabel polysilicon 324 -1802 324 -1802 0 1
rlabel polysilicon 324 -1808 324 -1808 0 3
rlabel polysilicon 331 -1802 331 -1802 0 1
rlabel polysilicon 331 -1808 331 -1808 0 3
rlabel polysilicon 338 -1802 338 -1802 0 1
rlabel polysilicon 338 -1808 338 -1808 0 3
rlabel polysilicon 345 -1802 345 -1802 0 1
rlabel polysilicon 345 -1808 345 -1808 0 3
rlabel polysilicon 352 -1802 352 -1802 0 1
rlabel polysilicon 355 -1802 355 -1802 0 2
rlabel polysilicon 352 -1808 352 -1808 0 3
rlabel polysilicon 355 -1808 355 -1808 0 4
rlabel polysilicon 359 -1802 359 -1802 0 1
rlabel polysilicon 359 -1808 359 -1808 0 3
rlabel polysilicon 369 -1802 369 -1802 0 2
rlabel polysilicon 369 -1808 369 -1808 0 4
rlabel polysilicon 376 -1802 376 -1802 0 2
rlabel polysilicon 373 -1808 373 -1808 0 3
rlabel polysilicon 383 -1802 383 -1802 0 2
rlabel polysilicon 380 -1808 380 -1808 0 3
rlabel polysilicon 387 -1802 387 -1802 0 1
rlabel polysilicon 387 -1808 387 -1808 0 3
rlabel polysilicon 394 -1808 394 -1808 0 3
rlabel polysilicon 401 -1802 401 -1802 0 1
rlabel polysilicon 401 -1808 401 -1808 0 3
rlabel polysilicon 408 -1802 408 -1802 0 1
rlabel polysilicon 408 -1808 408 -1808 0 3
rlabel polysilicon 415 -1802 415 -1802 0 1
rlabel polysilicon 415 -1808 415 -1808 0 3
rlabel polysilicon 422 -1802 422 -1802 0 1
rlabel polysilicon 422 -1808 422 -1808 0 3
rlabel polysilicon 429 -1802 429 -1802 0 1
rlabel polysilicon 429 -1808 429 -1808 0 3
rlabel polysilicon 436 -1802 436 -1802 0 1
rlabel polysilicon 436 -1808 436 -1808 0 3
rlabel polysilicon 443 -1802 443 -1802 0 1
rlabel polysilicon 443 -1808 443 -1808 0 3
rlabel polysilicon 450 -1802 450 -1802 0 1
rlabel polysilicon 450 -1808 450 -1808 0 3
rlabel polysilicon 457 -1802 457 -1802 0 1
rlabel polysilicon 457 -1808 457 -1808 0 3
rlabel polysilicon 464 -1802 464 -1802 0 1
rlabel polysilicon 464 -1808 464 -1808 0 3
rlabel polysilicon 471 -1802 471 -1802 0 1
rlabel polysilicon 474 -1802 474 -1802 0 2
rlabel polysilicon 478 -1802 478 -1802 0 1
rlabel polysilicon 478 -1808 478 -1808 0 3
rlabel polysilicon 485 -1802 485 -1802 0 1
rlabel polysilicon 485 -1808 485 -1808 0 3
rlabel polysilicon 495 -1802 495 -1802 0 2
rlabel polysilicon 492 -1808 492 -1808 0 3
rlabel polysilicon 495 -1808 495 -1808 0 4
rlabel polysilicon 499 -1802 499 -1802 0 1
rlabel polysilicon 499 -1808 499 -1808 0 3
rlabel polysilicon 506 -1802 506 -1802 0 1
rlabel polysilicon 506 -1808 506 -1808 0 3
rlabel polysilicon 509 -1808 509 -1808 0 4
rlabel polysilicon 513 -1802 513 -1802 0 1
rlabel polysilicon 516 -1808 516 -1808 0 4
rlabel polysilicon 523 -1802 523 -1802 0 2
rlabel polysilicon 527 -1802 527 -1802 0 1
rlabel polysilicon 527 -1808 527 -1808 0 3
rlabel polysilicon 534 -1802 534 -1802 0 1
rlabel polysilicon 534 -1808 534 -1808 0 3
rlabel polysilicon 541 -1802 541 -1802 0 1
rlabel polysilicon 541 -1808 541 -1808 0 3
rlabel polysilicon 548 -1802 548 -1802 0 1
rlabel polysilicon 548 -1808 548 -1808 0 3
rlabel polysilicon 555 -1802 555 -1802 0 1
rlabel polysilicon 555 -1808 555 -1808 0 3
rlabel polysilicon 562 -1802 562 -1802 0 1
rlabel polysilicon 562 -1808 562 -1808 0 3
rlabel polysilicon 569 -1802 569 -1802 0 1
rlabel polysilicon 569 -1808 569 -1808 0 3
rlabel polysilicon 576 -1802 576 -1802 0 1
rlabel polysilicon 576 -1808 576 -1808 0 3
rlabel polysilicon 583 -1802 583 -1802 0 1
rlabel polysilicon 583 -1808 583 -1808 0 3
rlabel polysilicon 590 -1802 590 -1802 0 1
rlabel polysilicon 590 -1808 590 -1808 0 3
rlabel polysilicon 597 -1802 597 -1802 0 1
rlabel polysilicon 597 -1808 597 -1808 0 3
rlabel polysilicon 604 -1802 604 -1802 0 1
rlabel polysilicon 604 -1808 604 -1808 0 3
rlabel polysilicon 611 -1802 611 -1802 0 1
rlabel polysilicon 611 -1808 611 -1808 0 3
rlabel polysilicon 618 -1802 618 -1802 0 1
rlabel polysilicon 618 -1808 618 -1808 0 3
rlabel polysilicon 625 -1802 625 -1802 0 1
rlabel polysilicon 625 -1808 625 -1808 0 3
rlabel polysilicon 632 -1802 632 -1802 0 1
rlabel polysilicon 632 -1808 632 -1808 0 3
rlabel polysilicon 639 -1802 639 -1802 0 1
rlabel polysilicon 642 -1802 642 -1802 0 2
rlabel polysilicon 646 -1802 646 -1802 0 1
rlabel polysilicon 646 -1808 646 -1808 0 3
rlabel polysilicon 653 -1802 653 -1802 0 1
rlabel polysilicon 653 -1808 653 -1808 0 3
rlabel polysilicon 660 -1802 660 -1802 0 1
rlabel polysilicon 660 -1808 660 -1808 0 3
rlabel polysilicon 667 -1802 667 -1802 0 1
rlabel polysilicon 667 -1808 667 -1808 0 3
rlabel polysilicon 674 -1802 674 -1802 0 1
rlabel polysilicon 674 -1808 674 -1808 0 3
rlabel polysilicon 681 -1802 681 -1802 0 1
rlabel polysilicon 681 -1808 681 -1808 0 3
rlabel polysilicon 688 -1802 688 -1802 0 1
rlabel polysilicon 688 -1808 688 -1808 0 3
rlabel polysilicon 695 -1802 695 -1802 0 1
rlabel polysilicon 695 -1808 695 -1808 0 3
rlabel polysilicon 702 -1802 702 -1802 0 1
rlabel polysilicon 702 -1808 702 -1808 0 3
rlabel polysilicon 709 -1802 709 -1802 0 1
rlabel polysilicon 709 -1808 709 -1808 0 3
rlabel polysilicon 716 -1802 716 -1802 0 1
rlabel polysilicon 716 -1808 716 -1808 0 3
rlabel polysilicon 723 -1802 723 -1802 0 1
rlabel polysilicon 723 -1808 723 -1808 0 3
rlabel polysilicon 730 -1802 730 -1802 0 1
rlabel polysilicon 730 -1808 730 -1808 0 3
rlabel polysilicon 737 -1802 737 -1802 0 1
rlabel polysilicon 737 -1808 737 -1808 0 3
rlabel polysilicon 744 -1802 744 -1802 0 1
rlabel polysilicon 744 -1808 744 -1808 0 3
rlabel polysilicon 751 -1802 751 -1802 0 1
rlabel polysilicon 751 -1808 751 -1808 0 3
rlabel polysilicon 758 -1802 758 -1802 0 1
rlabel polysilicon 758 -1808 758 -1808 0 3
rlabel polysilicon 905 -1802 905 -1802 0 1
rlabel polysilicon 5 -1889 5 -1889 0 4
rlabel polysilicon 12 -1889 12 -1889 0 4
rlabel polysilicon 16 -1883 16 -1883 0 1
rlabel polysilicon 16 -1889 16 -1889 0 3
rlabel polysilicon 23 -1889 23 -1889 0 3
rlabel polysilicon 26 -1889 26 -1889 0 4
rlabel polysilicon 33 -1883 33 -1883 0 2
rlabel polysilicon 37 -1883 37 -1883 0 1
rlabel polysilicon 37 -1889 37 -1889 0 3
rlabel polysilicon 47 -1883 47 -1883 0 2
rlabel polysilicon 51 -1883 51 -1883 0 1
rlabel polysilicon 51 -1889 51 -1889 0 3
rlabel polysilicon 58 -1883 58 -1883 0 1
rlabel polysilicon 58 -1889 58 -1889 0 3
rlabel polysilicon 65 -1883 65 -1883 0 1
rlabel polysilicon 65 -1889 65 -1889 0 3
rlabel polysilicon 72 -1883 72 -1883 0 1
rlabel polysilicon 72 -1889 72 -1889 0 3
rlabel polysilicon 79 -1883 79 -1883 0 1
rlabel polysilicon 79 -1889 79 -1889 0 3
rlabel polysilicon 86 -1883 86 -1883 0 1
rlabel polysilicon 86 -1889 86 -1889 0 3
rlabel polysilicon 93 -1883 93 -1883 0 1
rlabel polysilicon 93 -1889 93 -1889 0 3
rlabel polysilicon 100 -1883 100 -1883 0 1
rlabel polysilicon 100 -1889 100 -1889 0 3
rlabel polysilicon 107 -1883 107 -1883 0 1
rlabel polysilicon 107 -1889 107 -1889 0 3
rlabel polysilicon 114 -1883 114 -1883 0 1
rlabel polysilicon 114 -1889 114 -1889 0 3
rlabel polysilicon 121 -1883 121 -1883 0 1
rlabel polysilicon 121 -1889 121 -1889 0 3
rlabel polysilicon 131 -1883 131 -1883 0 2
rlabel polysilicon 131 -1889 131 -1889 0 4
rlabel polysilicon 135 -1883 135 -1883 0 1
rlabel polysilicon 135 -1889 135 -1889 0 3
rlabel polysilicon 142 -1883 142 -1883 0 1
rlabel polysilicon 142 -1889 142 -1889 0 3
rlabel polysilicon 145 -1889 145 -1889 0 4
rlabel polysilicon 149 -1889 149 -1889 0 3
rlabel polysilicon 156 -1883 156 -1883 0 1
rlabel polysilicon 156 -1889 156 -1889 0 3
rlabel polysilicon 163 -1883 163 -1883 0 1
rlabel polysilicon 166 -1889 166 -1889 0 4
rlabel polysilicon 170 -1883 170 -1883 0 1
rlabel polysilicon 170 -1889 170 -1889 0 3
rlabel polysilicon 177 -1883 177 -1883 0 1
rlabel polysilicon 177 -1889 177 -1889 0 3
rlabel polysilicon 184 -1883 184 -1883 0 1
rlabel polysilicon 184 -1889 184 -1889 0 3
rlabel polysilicon 191 -1883 191 -1883 0 1
rlabel polysilicon 194 -1889 194 -1889 0 4
rlabel polysilicon 198 -1883 198 -1883 0 1
rlabel polysilicon 201 -1883 201 -1883 0 2
rlabel polysilicon 198 -1889 198 -1889 0 3
rlabel polysilicon 205 -1883 205 -1883 0 1
rlabel polysilicon 205 -1889 205 -1889 0 3
rlabel polysilicon 212 -1883 212 -1883 0 1
rlabel polysilicon 212 -1889 212 -1889 0 3
rlabel polysilicon 219 -1883 219 -1883 0 1
rlabel polysilicon 219 -1889 219 -1889 0 3
rlabel polysilicon 226 -1883 226 -1883 0 1
rlabel polysilicon 233 -1883 233 -1883 0 1
rlabel polysilicon 233 -1889 233 -1889 0 3
rlabel polysilicon 240 -1883 240 -1883 0 1
rlabel polysilicon 240 -1889 240 -1889 0 3
rlabel polysilicon 247 -1883 247 -1883 0 1
rlabel polysilicon 247 -1889 247 -1889 0 3
rlabel polysilicon 254 -1883 254 -1883 0 1
rlabel polysilicon 254 -1889 254 -1889 0 3
rlabel polysilicon 261 -1883 261 -1883 0 1
rlabel polysilicon 261 -1889 261 -1889 0 3
rlabel polysilicon 268 -1883 268 -1883 0 1
rlabel polysilicon 268 -1889 268 -1889 0 3
rlabel polysilicon 275 -1883 275 -1883 0 1
rlabel polysilicon 275 -1889 275 -1889 0 3
rlabel polysilicon 282 -1883 282 -1883 0 1
rlabel polysilicon 282 -1889 282 -1889 0 3
rlabel polysilicon 292 -1883 292 -1883 0 2
rlabel polysilicon 292 -1889 292 -1889 0 4
rlabel polysilicon 296 -1883 296 -1883 0 1
rlabel polysilicon 296 -1889 296 -1889 0 3
rlabel polysilicon 303 -1883 303 -1883 0 1
rlabel polysilicon 306 -1883 306 -1883 0 2
rlabel polysilicon 303 -1889 303 -1889 0 3
rlabel polysilicon 306 -1889 306 -1889 0 4
rlabel polysilicon 310 -1883 310 -1883 0 1
rlabel polysilicon 310 -1889 310 -1889 0 3
rlabel polysilicon 317 -1883 317 -1883 0 1
rlabel polysilicon 317 -1889 317 -1889 0 3
rlabel polysilicon 324 -1883 324 -1883 0 1
rlabel polysilicon 324 -1889 324 -1889 0 3
rlabel polysilicon 327 -1889 327 -1889 0 4
rlabel polysilicon 331 -1883 331 -1883 0 1
rlabel polysilicon 331 -1889 331 -1889 0 3
rlabel polysilicon 338 -1883 338 -1883 0 1
rlabel polysilicon 348 -1883 348 -1883 0 2
rlabel polysilicon 352 -1883 352 -1883 0 1
rlabel polysilicon 355 -1883 355 -1883 0 2
rlabel polysilicon 362 -1883 362 -1883 0 2
rlabel polysilicon 359 -1889 359 -1889 0 3
rlabel polysilicon 362 -1889 362 -1889 0 4
rlabel polysilicon 366 -1883 366 -1883 0 1
rlabel polysilicon 366 -1889 366 -1889 0 3
rlabel polysilicon 373 -1883 373 -1883 0 1
rlabel polysilicon 376 -1883 376 -1883 0 2
rlabel polysilicon 376 -1889 376 -1889 0 4
rlabel polysilicon 380 -1883 380 -1883 0 1
rlabel polysilicon 380 -1889 380 -1889 0 3
rlabel polysilicon 387 -1883 387 -1883 0 1
rlabel polysilicon 390 -1883 390 -1883 0 2
rlabel polysilicon 387 -1889 387 -1889 0 3
rlabel polysilicon 394 -1883 394 -1883 0 1
rlabel polysilicon 394 -1889 394 -1889 0 3
rlabel polysilicon 401 -1883 401 -1883 0 1
rlabel polysilicon 401 -1889 401 -1889 0 3
rlabel polysilicon 408 -1883 408 -1883 0 1
rlabel polysilicon 408 -1889 408 -1889 0 3
rlabel polysilicon 415 -1883 415 -1883 0 1
rlabel polysilicon 415 -1889 415 -1889 0 3
rlabel polysilicon 422 -1883 422 -1883 0 1
rlabel polysilicon 422 -1889 422 -1889 0 3
rlabel polysilicon 429 -1883 429 -1883 0 1
rlabel polysilicon 429 -1889 429 -1889 0 3
rlabel polysilicon 436 -1889 436 -1889 0 3
rlabel polysilicon 439 -1889 439 -1889 0 4
rlabel polysilicon 443 -1883 443 -1883 0 1
rlabel polysilicon 450 -1883 450 -1883 0 1
rlabel polysilicon 453 -1883 453 -1883 0 2
rlabel polysilicon 450 -1889 450 -1889 0 3
rlabel polysilicon 457 -1883 457 -1883 0 1
rlabel polysilicon 457 -1889 457 -1889 0 3
rlabel polysilicon 464 -1883 464 -1883 0 1
rlabel polysilicon 464 -1889 464 -1889 0 3
rlabel polysilicon 467 -1889 467 -1889 0 4
rlabel polysilicon 471 -1883 471 -1883 0 1
rlabel polysilicon 471 -1889 471 -1889 0 3
rlabel polysilicon 478 -1883 478 -1883 0 1
rlabel polysilicon 478 -1889 478 -1889 0 3
rlabel polysilicon 485 -1883 485 -1883 0 1
rlabel polysilicon 485 -1889 485 -1889 0 3
rlabel polysilicon 492 -1883 492 -1883 0 1
rlabel polysilicon 492 -1889 492 -1889 0 3
rlabel polysilicon 499 -1883 499 -1883 0 1
rlabel polysilicon 502 -1883 502 -1883 0 2
rlabel polysilicon 502 -1889 502 -1889 0 4
rlabel polysilicon 506 -1883 506 -1883 0 1
rlabel polysilicon 506 -1889 506 -1889 0 3
rlabel polysilicon 513 -1883 513 -1883 0 1
rlabel polysilicon 513 -1889 513 -1889 0 3
rlabel polysilicon 520 -1883 520 -1883 0 1
rlabel polysilicon 520 -1889 520 -1889 0 3
rlabel polysilicon 527 -1883 527 -1883 0 1
rlabel polysilicon 527 -1889 527 -1889 0 3
rlabel polysilicon 534 -1883 534 -1883 0 1
rlabel polysilicon 534 -1889 534 -1889 0 3
rlabel polysilicon 541 -1883 541 -1883 0 1
rlabel polysilicon 541 -1889 541 -1889 0 3
rlabel polysilicon 548 -1889 548 -1889 0 3
rlabel polysilicon 555 -1883 555 -1883 0 1
rlabel polysilicon 555 -1889 555 -1889 0 3
rlabel polysilicon 562 -1883 562 -1883 0 1
rlabel polysilicon 562 -1889 562 -1889 0 3
rlabel polysilicon 569 -1883 569 -1883 0 1
rlabel polysilicon 569 -1889 569 -1889 0 3
rlabel polysilicon 579 -1883 579 -1883 0 2
rlabel polysilicon 579 -1889 579 -1889 0 4
rlabel polysilicon 583 -1883 583 -1883 0 1
rlabel polysilicon 583 -1889 583 -1889 0 3
rlabel polysilicon 590 -1883 590 -1883 0 1
rlabel polysilicon 590 -1889 590 -1889 0 3
rlabel polysilicon 597 -1883 597 -1883 0 1
rlabel polysilicon 597 -1889 597 -1889 0 3
rlabel polysilicon 604 -1883 604 -1883 0 1
rlabel polysilicon 604 -1889 604 -1889 0 3
rlabel polysilicon 611 -1883 611 -1883 0 1
rlabel polysilicon 611 -1889 611 -1889 0 3
rlabel polysilicon 618 -1883 618 -1883 0 1
rlabel polysilicon 618 -1889 618 -1889 0 3
rlabel polysilicon 625 -1883 625 -1883 0 1
rlabel polysilicon 625 -1889 625 -1889 0 3
rlabel polysilicon 632 -1883 632 -1883 0 1
rlabel polysilicon 632 -1889 632 -1889 0 3
rlabel polysilicon 642 -1883 642 -1883 0 2
rlabel polysilicon 639 -1889 639 -1889 0 3
rlabel polysilicon 646 -1883 646 -1883 0 1
rlabel polysilicon 646 -1889 646 -1889 0 3
rlabel polysilicon 653 -1883 653 -1883 0 1
rlabel polysilicon 653 -1889 653 -1889 0 3
rlabel polysilicon 660 -1883 660 -1883 0 1
rlabel polysilicon 660 -1889 660 -1889 0 3
rlabel polysilicon 667 -1883 667 -1883 0 1
rlabel polysilicon 667 -1889 667 -1889 0 3
rlabel polysilicon 674 -1883 674 -1883 0 1
rlabel polysilicon 674 -1889 674 -1889 0 3
rlabel polysilicon 681 -1883 681 -1883 0 1
rlabel polysilicon 681 -1889 681 -1889 0 3
rlabel polysilicon 688 -1883 688 -1883 0 1
rlabel polysilicon 688 -1889 688 -1889 0 3
rlabel polysilicon 695 -1883 695 -1883 0 1
rlabel polysilicon 695 -1889 695 -1889 0 3
rlabel polysilicon 702 -1883 702 -1883 0 1
rlabel polysilicon 702 -1889 702 -1889 0 3
rlabel polysilicon 709 -1883 709 -1883 0 1
rlabel polysilicon 709 -1889 709 -1889 0 3
rlabel polysilicon 716 -1883 716 -1883 0 1
rlabel polysilicon 716 -1889 716 -1889 0 3
rlabel polysilicon 723 -1883 723 -1883 0 1
rlabel polysilicon 723 -1889 723 -1889 0 3
rlabel polysilicon 730 -1883 730 -1883 0 1
rlabel polysilicon 730 -1889 730 -1889 0 3
rlabel polysilicon 737 -1883 737 -1883 0 1
rlabel polysilicon 737 -1889 737 -1889 0 3
rlabel polysilicon 744 -1883 744 -1883 0 1
rlabel polysilicon 747 -1883 747 -1883 0 2
rlabel polysilicon 747 -1889 747 -1889 0 4
rlabel polysilicon 751 -1883 751 -1883 0 1
rlabel polysilicon 751 -1889 751 -1889 0 3
rlabel polysilicon 2 -1966 2 -1966 0 1
rlabel polysilicon 2 -1972 2 -1972 0 3
rlabel polysilicon 9 -1966 9 -1966 0 1
rlabel polysilicon 9 -1972 9 -1972 0 3
rlabel polysilicon 19 -1966 19 -1966 0 2
rlabel polysilicon 19 -1972 19 -1972 0 4
rlabel polysilicon 23 -1966 23 -1966 0 1
rlabel polysilicon 23 -1972 23 -1972 0 3
rlabel polysilicon 33 -1966 33 -1966 0 2
rlabel polysilicon 30 -1972 30 -1972 0 3
rlabel polysilicon 37 -1966 37 -1966 0 1
rlabel polysilicon 44 -1966 44 -1966 0 1
rlabel polysilicon 44 -1972 44 -1972 0 3
rlabel polysilicon 51 -1966 51 -1966 0 1
rlabel polysilicon 54 -1966 54 -1966 0 2
rlabel polysilicon 54 -1972 54 -1972 0 4
rlabel polysilicon 61 -1966 61 -1966 0 2
rlabel polysilicon 65 -1966 65 -1966 0 1
rlabel polysilicon 65 -1972 65 -1972 0 3
rlabel polysilicon 72 -1966 72 -1966 0 1
rlabel polysilicon 75 -1972 75 -1972 0 4
rlabel polysilicon 79 -1966 79 -1966 0 1
rlabel polysilicon 86 -1966 86 -1966 0 1
rlabel polysilicon 86 -1972 86 -1972 0 3
rlabel polysilicon 93 -1966 93 -1966 0 1
rlabel polysilicon 93 -1972 93 -1972 0 3
rlabel polysilicon 100 -1966 100 -1966 0 1
rlabel polysilicon 100 -1972 100 -1972 0 3
rlabel polysilicon 107 -1972 107 -1972 0 3
rlabel polysilicon 110 -1972 110 -1972 0 4
rlabel polysilicon 117 -1966 117 -1966 0 2
rlabel polysilicon 117 -1972 117 -1972 0 4
rlabel polysilicon 121 -1966 121 -1966 0 1
rlabel polysilicon 121 -1972 121 -1972 0 3
rlabel polysilicon 128 -1966 128 -1966 0 1
rlabel polysilicon 128 -1972 128 -1972 0 3
rlabel polysilicon 135 -1966 135 -1966 0 1
rlabel polysilicon 135 -1972 135 -1972 0 3
rlabel polysilicon 142 -1966 142 -1966 0 1
rlabel polysilicon 142 -1972 142 -1972 0 3
rlabel polysilicon 149 -1966 149 -1966 0 1
rlabel polysilicon 149 -1972 149 -1972 0 3
rlabel polysilicon 156 -1966 156 -1966 0 1
rlabel polysilicon 156 -1972 156 -1972 0 3
rlabel polysilicon 159 -1972 159 -1972 0 4
rlabel polysilicon 163 -1966 163 -1966 0 1
rlabel polysilicon 163 -1972 163 -1972 0 3
rlabel polysilicon 170 -1966 170 -1966 0 1
rlabel polysilicon 170 -1972 170 -1972 0 3
rlabel polysilicon 173 -1972 173 -1972 0 4
rlabel polysilicon 177 -1966 177 -1966 0 1
rlabel polysilicon 177 -1972 177 -1972 0 3
rlabel polysilicon 184 -1966 184 -1966 0 1
rlabel polysilicon 184 -1972 184 -1972 0 3
rlabel polysilicon 191 -1966 191 -1966 0 1
rlabel polysilicon 191 -1972 191 -1972 0 3
rlabel polysilicon 201 -1966 201 -1966 0 2
rlabel polysilicon 201 -1972 201 -1972 0 4
rlabel polysilicon 205 -1966 205 -1966 0 1
rlabel polysilicon 208 -1966 208 -1966 0 2
rlabel polysilicon 208 -1972 208 -1972 0 4
rlabel polysilicon 212 -1966 212 -1966 0 1
rlabel polysilicon 212 -1972 212 -1972 0 3
rlabel polysilicon 215 -1972 215 -1972 0 4
rlabel polysilicon 219 -1966 219 -1966 0 1
rlabel polysilicon 222 -1966 222 -1966 0 2
rlabel polysilicon 219 -1972 219 -1972 0 3
rlabel polysilicon 226 -1966 226 -1966 0 1
rlabel polysilicon 226 -1972 226 -1972 0 3
rlabel polysilicon 233 -1966 233 -1966 0 1
rlabel polysilicon 233 -1972 233 -1972 0 3
rlabel polysilicon 240 -1966 240 -1966 0 1
rlabel polysilicon 240 -1972 240 -1972 0 3
rlabel polysilicon 247 -1966 247 -1966 0 1
rlabel polysilicon 247 -1972 247 -1972 0 3
rlabel polysilicon 254 -1966 254 -1966 0 1
rlabel polysilicon 254 -1972 254 -1972 0 3
rlabel polysilicon 261 -1966 261 -1966 0 1
rlabel polysilicon 261 -1972 261 -1972 0 3
rlabel polysilicon 268 -1966 268 -1966 0 1
rlabel polysilicon 271 -1966 271 -1966 0 2
rlabel polysilicon 268 -1972 268 -1972 0 3
rlabel polysilicon 275 -1966 275 -1966 0 1
rlabel polysilicon 275 -1972 275 -1972 0 3
rlabel polysilicon 282 -1966 282 -1966 0 1
rlabel polysilicon 282 -1972 282 -1972 0 3
rlabel polysilicon 289 -1966 289 -1966 0 1
rlabel polysilicon 289 -1972 289 -1972 0 3
rlabel polysilicon 296 -1966 296 -1966 0 1
rlabel polysilicon 296 -1972 296 -1972 0 3
rlabel polysilicon 303 -1966 303 -1966 0 1
rlabel polysilicon 303 -1972 303 -1972 0 3
rlabel polysilicon 310 -1966 310 -1966 0 1
rlabel polysilicon 313 -1972 313 -1972 0 4
rlabel polysilicon 317 -1966 317 -1966 0 1
rlabel polysilicon 317 -1972 317 -1972 0 3
rlabel polysilicon 324 -1966 324 -1966 0 1
rlabel polysilicon 324 -1972 324 -1972 0 3
rlabel polysilicon 331 -1966 331 -1966 0 1
rlabel polysilicon 331 -1972 331 -1972 0 3
rlabel polysilicon 338 -1966 338 -1966 0 1
rlabel polysilicon 338 -1972 338 -1972 0 3
rlabel polysilicon 345 -1966 345 -1966 0 1
rlabel polysilicon 348 -1966 348 -1966 0 2
rlabel polysilicon 345 -1972 345 -1972 0 3
rlabel polysilicon 348 -1972 348 -1972 0 4
rlabel polysilicon 352 -1966 352 -1966 0 1
rlabel polysilicon 355 -1966 355 -1966 0 2
rlabel polysilicon 359 -1966 359 -1966 0 1
rlabel polysilicon 359 -1972 359 -1972 0 3
rlabel polysilicon 366 -1966 366 -1966 0 1
rlabel polysilicon 369 -1966 369 -1966 0 2
rlabel polysilicon 366 -1972 366 -1972 0 3
rlabel polysilicon 369 -1972 369 -1972 0 4
rlabel polysilicon 373 -1966 373 -1966 0 1
rlabel polysilicon 373 -1972 373 -1972 0 3
rlabel polysilicon 380 -1966 380 -1966 0 1
rlabel polysilicon 380 -1972 380 -1972 0 3
rlabel polysilicon 387 -1972 387 -1972 0 3
rlabel polysilicon 394 -1966 394 -1966 0 1
rlabel polysilicon 397 -1966 397 -1966 0 2
rlabel polysilicon 397 -1972 397 -1972 0 4
rlabel polysilicon 401 -1966 401 -1966 0 1
rlabel polysilicon 401 -1972 401 -1972 0 3
rlabel polysilicon 408 -1966 408 -1966 0 1
rlabel polysilicon 408 -1972 408 -1972 0 3
rlabel polysilicon 418 -1966 418 -1966 0 2
rlabel polysilicon 415 -1972 415 -1972 0 3
rlabel polysilicon 418 -1972 418 -1972 0 4
rlabel polysilicon 422 -1966 422 -1966 0 1
rlabel polysilicon 429 -1966 429 -1966 0 1
rlabel polysilicon 432 -1966 432 -1966 0 2
rlabel polysilicon 429 -1972 429 -1972 0 3
rlabel polysilicon 432 -1972 432 -1972 0 4
rlabel polysilicon 436 -1966 436 -1966 0 1
rlabel polysilicon 436 -1972 436 -1972 0 3
rlabel polysilicon 443 -1966 443 -1966 0 1
rlabel polysilicon 443 -1972 443 -1972 0 3
rlabel polysilicon 450 -1966 450 -1966 0 1
rlabel polysilicon 450 -1972 450 -1972 0 3
rlabel polysilicon 460 -1966 460 -1966 0 2
rlabel polysilicon 457 -1972 457 -1972 0 3
rlabel polysilicon 464 -1972 464 -1972 0 3
rlabel polysilicon 471 -1966 471 -1966 0 1
rlabel polysilicon 471 -1972 471 -1972 0 3
rlabel polysilicon 478 -1966 478 -1966 0 1
rlabel polysilicon 481 -1966 481 -1966 0 2
rlabel polysilicon 481 -1972 481 -1972 0 4
rlabel polysilicon 485 -1966 485 -1966 0 1
rlabel polysilicon 485 -1972 485 -1972 0 3
rlabel polysilicon 492 -1966 492 -1966 0 1
rlabel polysilicon 492 -1972 492 -1972 0 3
rlabel polysilicon 499 -1966 499 -1966 0 1
rlabel polysilicon 499 -1972 499 -1972 0 3
rlabel polysilicon 506 -1966 506 -1966 0 1
rlabel polysilicon 506 -1972 506 -1972 0 3
rlabel polysilicon 513 -1966 513 -1966 0 1
rlabel polysilicon 513 -1972 513 -1972 0 3
rlabel polysilicon 520 -1966 520 -1966 0 1
rlabel polysilicon 520 -1972 520 -1972 0 3
rlabel polysilicon 527 -1966 527 -1966 0 1
rlabel polysilicon 527 -1972 527 -1972 0 3
rlabel polysilicon 534 -1966 534 -1966 0 1
rlabel polysilicon 534 -1972 534 -1972 0 3
rlabel polysilicon 541 -1966 541 -1966 0 1
rlabel polysilicon 541 -1972 541 -1972 0 3
rlabel polysilicon 548 -1972 548 -1972 0 3
rlabel polysilicon 551 -1972 551 -1972 0 4
rlabel polysilicon 555 -1966 555 -1966 0 1
rlabel polysilicon 555 -1972 555 -1972 0 3
rlabel polysilicon 562 -1966 562 -1966 0 1
rlabel polysilicon 562 -1972 562 -1972 0 3
rlabel polysilicon 569 -1966 569 -1966 0 1
rlabel polysilicon 569 -1972 569 -1972 0 3
rlabel polysilicon 576 -1966 576 -1966 0 1
rlabel polysilicon 576 -1972 576 -1972 0 3
rlabel polysilicon 583 -1966 583 -1966 0 1
rlabel polysilicon 583 -1972 583 -1972 0 3
rlabel polysilicon 590 -1966 590 -1966 0 1
rlabel polysilicon 590 -1972 590 -1972 0 3
rlabel polysilicon 597 -1966 597 -1966 0 1
rlabel polysilicon 597 -1972 597 -1972 0 3
rlabel polysilicon 604 -1966 604 -1966 0 1
rlabel polysilicon 604 -1972 604 -1972 0 3
rlabel polysilicon 611 -1966 611 -1966 0 1
rlabel polysilicon 611 -1972 611 -1972 0 3
rlabel polysilicon 618 -1966 618 -1966 0 1
rlabel polysilicon 618 -1972 618 -1972 0 3
rlabel polysilicon 625 -1966 625 -1966 0 1
rlabel polysilicon 625 -1972 625 -1972 0 3
rlabel polysilicon 632 -1966 632 -1966 0 1
rlabel polysilicon 632 -1972 632 -1972 0 3
rlabel polysilicon 639 -1972 639 -1972 0 3
rlabel polysilicon 642 -1972 642 -1972 0 4
rlabel polysilicon 646 -1966 646 -1966 0 1
rlabel polysilicon 646 -1972 646 -1972 0 3
rlabel polysilicon 653 -1966 653 -1966 0 1
rlabel polysilicon 653 -1972 653 -1972 0 3
rlabel polysilicon 660 -1966 660 -1966 0 1
rlabel polysilicon 660 -1972 660 -1972 0 3
rlabel polysilicon 667 -1966 667 -1966 0 1
rlabel polysilicon 667 -1972 667 -1972 0 3
rlabel polysilicon 674 -1966 674 -1966 0 1
rlabel polysilicon 674 -1972 674 -1972 0 3
rlabel polysilicon 681 -1966 681 -1966 0 1
rlabel polysilicon 681 -1972 681 -1972 0 3
rlabel polysilicon 688 -1966 688 -1966 0 1
rlabel polysilicon 688 -1972 688 -1972 0 3
rlabel polysilicon 695 -1966 695 -1966 0 1
rlabel polysilicon 695 -1972 695 -1972 0 3
rlabel polysilicon 702 -1966 702 -1966 0 1
rlabel polysilicon 702 -1972 702 -1972 0 3
rlabel polysilicon 709 -1966 709 -1966 0 1
rlabel polysilicon 709 -1972 709 -1972 0 3
rlabel polysilicon 716 -1966 716 -1966 0 1
rlabel polysilicon 716 -1972 716 -1972 0 3
rlabel polysilicon 723 -1966 723 -1966 0 1
rlabel polysilicon 723 -1972 723 -1972 0 3
rlabel polysilicon 730 -1966 730 -1966 0 1
rlabel polysilicon 730 -1972 730 -1972 0 3
rlabel polysilicon 9 -2027 9 -2027 0 1
rlabel polysilicon 9 -2033 9 -2033 0 3
rlabel polysilicon 16 -2027 16 -2027 0 1
rlabel polysilicon 16 -2033 16 -2033 0 3
rlabel polysilicon 23 -2027 23 -2027 0 1
rlabel polysilicon 30 -2027 30 -2027 0 1
rlabel polysilicon 30 -2033 30 -2033 0 3
rlabel polysilicon 37 -2027 37 -2027 0 1
rlabel polysilicon 37 -2033 37 -2033 0 3
rlabel polysilicon 44 -2027 44 -2027 0 1
rlabel polysilicon 44 -2033 44 -2033 0 3
rlabel polysilicon 51 -2027 51 -2027 0 1
rlabel polysilicon 54 -2027 54 -2027 0 2
rlabel polysilicon 51 -2033 51 -2033 0 3
rlabel polysilicon 58 -2027 58 -2027 0 1
rlabel polysilicon 58 -2033 58 -2033 0 3
rlabel polysilicon 65 -2027 65 -2027 0 1
rlabel polysilicon 68 -2027 68 -2027 0 2
rlabel polysilicon 65 -2033 65 -2033 0 3
rlabel polysilicon 72 -2027 72 -2027 0 1
rlabel polysilicon 72 -2033 72 -2033 0 3
rlabel polysilicon 79 -2027 79 -2027 0 1
rlabel polysilicon 79 -2033 79 -2033 0 3
rlabel polysilicon 89 -2027 89 -2027 0 2
rlabel polysilicon 86 -2033 86 -2033 0 3
rlabel polysilicon 89 -2033 89 -2033 0 4
rlabel polysilicon 96 -2033 96 -2033 0 4
rlabel polysilicon 100 -2027 100 -2027 0 1
rlabel polysilicon 103 -2027 103 -2027 0 2
rlabel polysilicon 107 -2027 107 -2027 0 1
rlabel polysilicon 107 -2033 107 -2033 0 3
rlabel polysilicon 117 -2027 117 -2027 0 2
rlabel polysilicon 114 -2033 114 -2033 0 3
rlabel polysilicon 117 -2033 117 -2033 0 4
rlabel polysilicon 121 -2027 121 -2027 0 1
rlabel polysilicon 121 -2033 121 -2033 0 3
rlabel polysilicon 128 -2027 128 -2027 0 1
rlabel polysilicon 131 -2027 131 -2027 0 2
rlabel polysilicon 128 -2033 128 -2033 0 3
rlabel polysilicon 135 -2027 135 -2027 0 1
rlabel polysilicon 135 -2033 135 -2033 0 3
rlabel polysilicon 142 -2027 142 -2027 0 1
rlabel polysilicon 142 -2033 142 -2033 0 3
rlabel polysilicon 149 -2027 149 -2027 0 1
rlabel polysilicon 149 -2033 149 -2033 0 3
rlabel polysilicon 156 -2027 156 -2027 0 1
rlabel polysilicon 156 -2033 156 -2033 0 3
rlabel polysilicon 163 -2027 163 -2027 0 1
rlabel polysilicon 163 -2033 163 -2033 0 3
rlabel polysilicon 170 -2027 170 -2027 0 1
rlabel polysilicon 170 -2033 170 -2033 0 3
rlabel polysilicon 177 -2027 177 -2027 0 1
rlabel polysilicon 177 -2033 177 -2033 0 3
rlabel polysilicon 184 -2027 184 -2027 0 1
rlabel polysilicon 184 -2033 184 -2033 0 3
rlabel polysilicon 191 -2033 191 -2033 0 3
rlabel polysilicon 198 -2033 198 -2033 0 3
rlabel polysilicon 201 -2033 201 -2033 0 4
rlabel polysilicon 205 -2027 205 -2027 0 1
rlabel polysilicon 205 -2033 205 -2033 0 3
rlabel polysilicon 212 -2033 212 -2033 0 3
rlabel polysilicon 215 -2033 215 -2033 0 4
rlabel polysilicon 219 -2027 219 -2027 0 1
rlabel polysilicon 219 -2033 219 -2033 0 3
rlabel polysilicon 222 -2033 222 -2033 0 4
rlabel polysilicon 226 -2027 226 -2027 0 1
rlabel polysilicon 226 -2033 226 -2033 0 3
rlabel polysilicon 233 -2027 233 -2027 0 1
rlabel polysilicon 233 -2033 233 -2033 0 3
rlabel polysilicon 240 -2027 240 -2027 0 1
rlabel polysilicon 240 -2033 240 -2033 0 3
rlabel polysilicon 247 -2027 247 -2027 0 1
rlabel polysilicon 254 -2033 254 -2033 0 3
rlabel polysilicon 257 -2033 257 -2033 0 4
rlabel polysilicon 261 -2027 261 -2027 0 1
rlabel polysilicon 261 -2033 261 -2033 0 3
rlabel polysilicon 268 -2027 268 -2027 0 1
rlabel polysilicon 268 -2033 268 -2033 0 3
rlabel polysilicon 275 -2027 275 -2027 0 1
rlabel polysilicon 275 -2033 275 -2033 0 3
rlabel polysilicon 282 -2027 282 -2027 0 1
rlabel polysilicon 285 -2027 285 -2027 0 2
rlabel polysilicon 282 -2033 282 -2033 0 3
rlabel polysilicon 289 -2027 289 -2027 0 1
rlabel polysilicon 289 -2033 289 -2033 0 3
rlabel polysilicon 296 -2027 296 -2027 0 1
rlabel polysilicon 296 -2033 296 -2033 0 3
rlabel polysilicon 303 -2027 303 -2027 0 1
rlabel polysilicon 306 -2027 306 -2027 0 2
rlabel polysilicon 303 -2033 303 -2033 0 3
rlabel polysilicon 310 -2027 310 -2027 0 1
rlabel polysilicon 310 -2033 310 -2033 0 3
rlabel polysilicon 317 -2027 317 -2027 0 1
rlabel polysilicon 317 -2033 317 -2033 0 3
rlabel polysilicon 324 -2027 324 -2027 0 1
rlabel polysilicon 324 -2033 324 -2033 0 3
rlabel polysilicon 331 -2027 331 -2027 0 1
rlabel polysilicon 331 -2033 331 -2033 0 3
rlabel polysilicon 338 -2027 338 -2027 0 1
rlabel polysilicon 338 -2033 338 -2033 0 3
rlabel polysilicon 345 -2027 345 -2027 0 1
rlabel polysilicon 345 -2033 345 -2033 0 3
rlabel polysilicon 352 -2027 352 -2027 0 1
rlabel polysilicon 352 -2033 352 -2033 0 3
rlabel polysilicon 359 -2027 359 -2027 0 1
rlabel polysilicon 359 -2033 359 -2033 0 3
rlabel polysilicon 366 -2027 366 -2027 0 1
rlabel polysilicon 366 -2033 366 -2033 0 3
rlabel polysilicon 373 -2027 373 -2027 0 1
rlabel polysilicon 373 -2033 373 -2033 0 3
rlabel polysilicon 380 -2033 380 -2033 0 3
rlabel polysilicon 387 -2027 387 -2027 0 1
rlabel polysilicon 387 -2033 387 -2033 0 3
rlabel polysilicon 394 -2027 394 -2027 0 1
rlabel polysilicon 394 -2033 394 -2033 0 3
rlabel polysilicon 404 -2027 404 -2027 0 2
rlabel polysilicon 401 -2033 401 -2033 0 3
rlabel polysilicon 404 -2033 404 -2033 0 4
rlabel polysilicon 408 -2027 408 -2027 0 1
rlabel polysilicon 408 -2033 408 -2033 0 3
rlabel polysilicon 415 -2027 415 -2027 0 1
rlabel polysilicon 418 -2033 418 -2033 0 4
rlabel polysilicon 422 -2027 422 -2027 0 1
rlabel polysilicon 422 -2033 422 -2033 0 3
rlabel polysilicon 429 -2027 429 -2027 0 1
rlabel polysilicon 429 -2033 429 -2033 0 3
rlabel polysilicon 436 -2027 436 -2027 0 1
rlabel polysilicon 439 -2027 439 -2027 0 2
rlabel polysilicon 436 -2033 436 -2033 0 3
rlabel polysilicon 443 -2027 443 -2027 0 1
rlabel polysilicon 443 -2033 443 -2033 0 3
rlabel polysilicon 450 -2027 450 -2027 0 1
rlabel polysilicon 450 -2033 450 -2033 0 3
rlabel polysilicon 457 -2027 457 -2027 0 1
rlabel polysilicon 457 -2033 457 -2033 0 3
rlabel polysilicon 464 -2027 464 -2027 0 1
rlabel polysilicon 464 -2033 464 -2033 0 3
rlabel polysilicon 474 -2027 474 -2027 0 2
rlabel polysilicon 471 -2033 471 -2033 0 3
rlabel polysilicon 474 -2033 474 -2033 0 4
rlabel polysilicon 478 -2027 478 -2027 0 1
rlabel polysilicon 478 -2033 478 -2033 0 3
rlabel polysilicon 488 -2027 488 -2027 0 2
rlabel polysilicon 492 -2027 492 -2027 0 1
rlabel polysilicon 492 -2033 492 -2033 0 3
rlabel polysilicon 499 -2027 499 -2027 0 1
rlabel polysilicon 499 -2033 499 -2033 0 3
rlabel polysilicon 506 -2027 506 -2027 0 1
rlabel polysilicon 506 -2033 506 -2033 0 3
rlabel polysilicon 513 -2027 513 -2027 0 1
rlabel polysilicon 513 -2033 513 -2033 0 3
rlabel polysilicon 520 -2027 520 -2027 0 1
rlabel polysilicon 527 -2027 527 -2027 0 1
rlabel polysilicon 527 -2033 527 -2033 0 3
rlabel polysilicon 534 -2027 534 -2027 0 1
rlabel polysilicon 534 -2033 534 -2033 0 3
rlabel polysilicon 541 -2027 541 -2027 0 1
rlabel polysilicon 541 -2033 541 -2033 0 3
rlabel polysilicon 551 -2027 551 -2027 0 2
rlabel polysilicon 548 -2033 548 -2033 0 3
rlabel polysilicon 555 -2027 555 -2027 0 1
rlabel polysilicon 555 -2033 555 -2033 0 3
rlabel polysilicon 562 -2027 562 -2027 0 1
rlabel polysilicon 562 -2033 562 -2033 0 3
rlabel polysilicon 569 -2027 569 -2027 0 1
rlabel polysilicon 569 -2033 569 -2033 0 3
rlabel polysilicon 576 -2027 576 -2027 0 1
rlabel polysilicon 576 -2033 576 -2033 0 3
rlabel polysilicon 583 -2027 583 -2027 0 1
rlabel polysilicon 583 -2033 583 -2033 0 3
rlabel polysilicon 590 -2027 590 -2027 0 1
rlabel polysilicon 590 -2033 590 -2033 0 3
rlabel polysilicon 597 -2027 597 -2027 0 1
rlabel polysilicon 597 -2033 597 -2033 0 3
rlabel polysilicon 604 -2027 604 -2027 0 1
rlabel polysilicon 604 -2033 604 -2033 0 3
rlabel polysilicon 611 -2027 611 -2027 0 1
rlabel polysilicon 611 -2033 611 -2033 0 3
rlabel polysilicon 618 -2027 618 -2027 0 1
rlabel polysilicon 618 -2033 618 -2033 0 3
rlabel polysilicon 625 -2027 625 -2027 0 1
rlabel polysilicon 625 -2033 625 -2033 0 3
rlabel polysilicon 632 -2027 632 -2027 0 1
rlabel polysilicon 635 -2027 635 -2027 0 2
rlabel polysilicon 632 -2033 632 -2033 0 3
rlabel polysilicon 635 -2033 635 -2033 0 4
rlabel polysilicon 642 -2027 642 -2027 0 2
rlabel polysilicon 639 -2033 639 -2033 0 3
rlabel polysilicon 642 -2033 642 -2033 0 4
rlabel polysilicon 646 -2027 646 -2027 0 1
rlabel polysilicon 649 -2027 649 -2027 0 2
rlabel polysilicon 653 -2027 653 -2027 0 1
rlabel polysilicon 653 -2033 653 -2033 0 3
rlabel polysilicon 660 -2027 660 -2027 0 1
rlabel polysilicon 660 -2033 660 -2033 0 3
rlabel polysilicon 670 -2033 670 -2033 0 4
rlabel polysilicon 695 -2027 695 -2027 0 1
rlabel polysilicon 695 -2033 695 -2033 0 3
rlabel polysilicon 16 -2092 16 -2092 0 1
rlabel polysilicon 16 -2098 16 -2098 0 3
rlabel polysilicon 23 -2098 23 -2098 0 3
rlabel polysilicon 33 -2092 33 -2092 0 2
rlabel polysilicon 37 -2092 37 -2092 0 1
rlabel polysilicon 37 -2098 37 -2098 0 3
rlabel polysilicon 44 -2092 44 -2092 0 1
rlabel polysilicon 44 -2098 44 -2098 0 3
rlabel polysilicon 51 -2092 51 -2092 0 1
rlabel polysilicon 51 -2098 51 -2098 0 3
rlabel polysilicon 58 -2092 58 -2092 0 1
rlabel polysilicon 58 -2098 58 -2098 0 3
rlabel polysilicon 65 -2092 65 -2092 0 1
rlabel polysilicon 65 -2098 65 -2098 0 3
rlabel polysilicon 75 -2092 75 -2092 0 2
rlabel polysilicon 72 -2098 72 -2098 0 3
rlabel polysilicon 75 -2098 75 -2098 0 4
rlabel polysilicon 79 -2092 79 -2092 0 1
rlabel polysilicon 79 -2098 79 -2098 0 3
rlabel polysilicon 86 -2092 86 -2092 0 1
rlabel polysilicon 86 -2098 86 -2098 0 3
rlabel polysilicon 96 -2092 96 -2092 0 2
rlabel polysilicon 100 -2092 100 -2092 0 1
rlabel polysilicon 100 -2098 100 -2098 0 3
rlabel polysilicon 107 -2092 107 -2092 0 1
rlabel polysilicon 107 -2098 107 -2098 0 3
rlabel polysilicon 114 -2092 114 -2092 0 1
rlabel polysilicon 117 -2092 117 -2092 0 2
rlabel polysilicon 117 -2098 117 -2098 0 4
rlabel polysilicon 121 -2092 121 -2092 0 1
rlabel polysilicon 121 -2098 121 -2098 0 3
rlabel polysilicon 128 -2092 128 -2092 0 1
rlabel polysilicon 128 -2098 128 -2098 0 3
rlabel polysilicon 135 -2092 135 -2092 0 1
rlabel polysilicon 135 -2098 135 -2098 0 3
rlabel polysilicon 142 -2092 142 -2092 0 1
rlabel polysilicon 142 -2098 142 -2098 0 3
rlabel polysilicon 149 -2092 149 -2092 0 1
rlabel polysilicon 149 -2098 149 -2098 0 3
rlabel polysilicon 156 -2092 156 -2092 0 1
rlabel polysilicon 159 -2092 159 -2092 0 2
rlabel polysilicon 163 -2092 163 -2092 0 1
rlabel polysilicon 163 -2098 163 -2098 0 3
rlabel polysilicon 170 -2092 170 -2092 0 1
rlabel polysilicon 170 -2098 170 -2098 0 3
rlabel polysilicon 177 -2092 177 -2092 0 1
rlabel polysilicon 177 -2098 177 -2098 0 3
rlabel polysilicon 184 -2098 184 -2098 0 3
rlabel polysilicon 187 -2098 187 -2098 0 4
rlabel polysilicon 191 -2092 191 -2092 0 1
rlabel polysilicon 194 -2092 194 -2092 0 2
rlabel polysilicon 198 -2092 198 -2092 0 1
rlabel polysilicon 198 -2098 198 -2098 0 3
rlabel polysilicon 205 -2098 205 -2098 0 3
rlabel polysilicon 208 -2098 208 -2098 0 4
rlabel polysilicon 212 -2092 212 -2092 0 1
rlabel polysilicon 212 -2098 212 -2098 0 3
rlabel polysilicon 219 -2092 219 -2092 0 1
rlabel polysilicon 222 -2092 222 -2092 0 2
rlabel polysilicon 226 -2092 226 -2092 0 1
rlabel polysilicon 226 -2098 226 -2098 0 3
rlabel polysilicon 236 -2092 236 -2092 0 2
rlabel polysilicon 233 -2098 233 -2098 0 3
rlabel polysilicon 240 -2092 240 -2092 0 1
rlabel polysilicon 240 -2098 240 -2098 0 3
rlabel polysilicon 247 -2092 247 -2092 0 1
rlabel polysilicon 247 -2098 247 -2098 0 3
rlabel polysilicon 254 -2092 254 -2092 0 1
rlabel polysilicon 254 -2098 254 -2098 0 3
rlabel polysilicon 261 -2092 261 -2092 0 1
rlabel polysilicon 261 -2098 261 -2098 0 3
rlabel polysilicon 268 -2092 268 -2092 0 1
rlabel polysilicon 268 -2098 268 -2098 0 3
rlabel polysilicon 275 -2092 275 -2092 0 1
rlabel polysilicon 275 -2098 275 -2098 0 3
rlabel polysilicon 282 -2092 282 -2092 0 1
rlabel polysilicon 282 -2098 282 -2098 0 3
rlabel polysilicon 289 -2092 289 -2092 0 1
rlabel polysilicon 289 -2098 289 -2098 0 3
rlabel polysilicon 296 -2092 296 -2092 0 1
rlabel polysilicon 296 -2098 296 -2098 0 3
rlabel polysilicon 303 -2092 303 -2092 0 1
rlabel polysilicon 306 -2092 306 -2092 0 2
rlabel polysilicon 306 -2098 306 -2098 0 4
rlabel polysilicon 313 -2092 313 -2092 0 2
rlabel polysilicon 310 -2098 310 -2098 0 3
rlabel polysilicon 317 -2092 317 -2092 0 1
rlabel polysilicon 320 -2092 320 -2092 0 2
rlabel polysilicon 317 -2098 317 -2098 0 3
rlabel polysilicon 320 -2098 320 -2098 0 4
rlabel polysilicon 324 -2092 324 -2092 0 1
rlabel polysilicon 327 -2092 327 -2092 0 2
rlabel polysilicon 331 -2092 331 -2092 0 1
rlabel polysilicon 331 -2098 331 -2098 0 3
rlabel polysilicon 338 -2092 338 -2092 0 1
rlabel polysilicon 338 -2098 338 -2098 0 3
rlabel polysilicon 345 -2092 345 -2092 0 1
rlabel polysilicon 345 -2098 345 -2098 0 3
rlabel polysilicon 352 -2092 352 -2092 0 1
rlabel polysilicon 359 -2092 359 -2092 0 1
rlabel polysilicon 359 -2098 359 -2098 0 3
rlabel polysilicon 366 -2092 366 -2092 0 1
rlabel polysilicon 369 -2092 369 -2092 0 2
rlabel polysilicon 369 -2098 369 -2098 0 4
rlabel polysilicon 373 -2092 373 -2092 0 1
rlabel polysilicon 373 -2098 373 -2098 0 3
rlabel polysilicon 380 -2092 380 -2092 0 1
rlabel polysilicon 383 -2092 383 -2092 0 2
rlabel polysilicon 383 -2098 383 -2098 0 4
rlabel polysilicon 387 -2092 387 -2092 0 1
rlabel polysilicon 387 -2098 387 -2098 0 3
rlabel polysilicon 394 -2092 394 -2092 0 1
rlabel polysilicon 394 -2098 394 -2098 0 3
rlabel polysilicon 401 -2092 401 -2092 0 1
rlabel polysilicon 404 -2092 404 -2092 0 2
rlabel polysilicon 408 -2092 408 -2092 0 1
rlabel polysilicon 415 -2092 415 -2092 0 1
rlabel polysilicon 418 -2092 418 -2092 0 2
rlabel polysilicon 425 -2092 425 -2092 0 2
rlabel polysilicon 422 -2098 422 -2098 0 3
rlabel polysilicon 429 -2092 429 -2092 0 1
rlabel polysilicon 429 -2098 429 -2098 0 3
rlabel polysilicon 436 -2092 436 -2092 0 1
rlabel polysilicon 436 -2098 436 -2098 0 3
rlabel polysilicon 443 -2092 443 -2092 0 1
rlabel polysilicon 443 -2098 443 -2098 0 3
rlabel polysilicon 450 -2092 450 -2092 0 1
rlabel polysilicon 450 -2098 450 -2098 0 3
rlabel polysilicon 457 -2092 457 -2092 0 1
rlabel polysilicon 457 -2098 457 -2098 0 3
rlabel polysilicon 464 -2092 464 -2092 0 1
rlabel polysilicon 464 -2098 464 -2098 0 3
rlabel polysilicon 471 -2092 471 -2092 0 1
rlabel polysilicon 471 -2098 471 -2098 0 3
rlabel polysilicon 478 -2092 478 -2092 0 1
rlabel polysilicon 481 -2092 481 -2092 0 2
rlabel polysilicon 485 -2092 485 -2092 0 1
rlabel polysilicon 485 -2098 485 -2098 0 3
rlabel polysilicon 492 -2092 492 -2092 0 1
rlabel polysilicon 492 -2098 492 -2098 0 3
rlabel polysilicon 499 -2092 499 -2092 0 1
rlabel polysilicon 502 -2098 502 -2098 0 4
rlabel polysilicon 506 -2092 506 -2092 0 1
rlabel polysilicon 506 -2098 506 -2098 0 3
rlabel polysilicon 513 -2092 513 -2092 0 1
rlabel polysilicon 513 -2098 513 -2098 0 3
rlabel polysilicon 520 -2092 520 -2092 0 1
rlabel polysilicon 520 -2098 520 -2098 0 3
rlabel polysilicon 527 -2092 527 -2092 0 1
rlabel polysilicon 527 -2098 527 -2098 0 3
rlabel polysilicon 534 -2092 534 -2092 0 1
rlabel polysilicon 534 -2098 534 -2098 0 3
rlabel polysilicon 541 -2092 541 -2092 0 1
rlabel polysilicon 541 -2098 541 -2098 0 3
rlabel polysilicon 548 -2092 548 -2092 0 1
rlabel polysilicon 548 -2098 548 -2098 0 3
rlabel polysilicon 555 -2092 555 -2092 0 1
rlabel polysilicon 558 -2098 558 -2098 0 4
rlabel polysilicon 562 -2092 562 -2092 0 1
rlabel polysilicon 562 -2098 562 -2098 0 3
rlabel polysilicon 569 -2092 569 -2092 0 1
rlabel polysilicon 569 -2098 569 -2098 0 3
rlabel polysilicon 576 -2092 576 -2092 0 1
rlabel polysilicon 576 -2098 576 -2098 0 3
rlabel polysilicon 583 -2092 583 -2092 0 1
rlabel polysilicon 583 -2098 583 -2098 0 3
rlabel polysilicon 590 -2092 590 -2092 0 1
rlabel polysilicon 590 -2098 590 -2098 0 3
rlabel polysilicon 604 -2092 604 -2092 0 1
rlabel polysilicon 604 -2098 604 -2098 0 3
rlabel polysilicon 611 -2092 611 -2092 0 1
rlabel polysilicon 611 -2098 611 -2098 0 3
rlabel polysilicon 618 -2098 618 -2098 0 3
rlabel polysilicon 621 -2098 621 -2098 0 4
rlabel polysilicon 642 -2092 642 -2092 0 2
rlabel polysilicon 642 -2098 642 -2098 0 4
rlabel polysilicon 646 -2092 646 -2092 0 1
rlabel polysilicon 646 -2098 646 -2098 0 3
rlabel polysilicon 674 -2092 674 -2092 0 1
rlabel polysilicon 674 -2098 674 -2098 0 3
rlabel polysilicon 688 -2092 688 -2092 0 1
rlabel polysilicon 688 -2098 688 -2098 0 3
rlabel polysilicon 26 -2149 26 -2149 0 2
rlabel polysilicon 33 -2149 33 -2149 0 2
rlabel polysilicon 37 -2149 37 -2149 0 1
rlabel polysilicon 37 -2155 37 -2155 0 3
rlabel polysilicon 44 -2149 44 -2149 0 1
rlabel polysilicon 44 -2155 44 -2155 0 3
rlabel polysilicon 51 -2149 51 -2149 0 1
rlabel polysilicon 51 -2155 51 -2155 0 3
rlabel polysilicon 58 -2149 58 -2149 0 1
rlabel polysilicon 58 -2155 58 -2155 0 3
rlabel polysilicon 65 -2149 65 -2149 0 1
rlabel polysilicon 65 -2155 65 -2155 0 3
rlabel polysilicon 72 -2155 72 -2155 0 3
rlabel polysilicon 79 -2149 79 -2149 0 1
rlabel polysilicon 86 -2149 86 -2149 0 1
rlabel polysilicon 86 -2155 86 -2155 0 3
rlabel polysilicon 93 -2155 93 -2155 0 3
rlabel polysilicon 96 -2155 96 -2155 0 4
rlabel polysilicon 100 -2149 100 -2149 0 1
rlabel polysilicon 100 -2155 100 -2155 0 3
rlabel polysilicon 107 -2149 107 -2149 0 1
rlabel polysilicon 107 -2155 107 -2155 0 3
rlabel polysilicon 117 -2149 117 -2149 0 2
rlabel polysilicon 121 -2155 121 -2155 0 3
rlabel polysilicon 128 -2155 128 -2155 0 3
rlabel polysilicon 131 -2155 131 -2155 0 4
rlabel polysilicon 135 -2149 135 -2149 0 1
rlabel polysilicon 135 -2155 135 -2155 0 3
rlabel polysilicon 142 -2149 142 -2149 0 1
rlabel polysilicon 142 -2155 142 -2155 0 3
rlabel polysilicon 152 -2149 152 -2149 0 2
rlabel polysilicon 156 -2149 156 -2149 0 1
rlabel polysilicon 156 -2155 156 -2155 0 3
rlabel polysilicon 163 -2149 163 -2149 0 1
rlabel polysilicon 163 -2155 163 -2155 0 3
rlabel polysilicon 170 -2149 170 -2149 0 1
rlabel polysilicon 170 -2155 170 -2155 0 3
rlabel polysilicon 177 -2149 177 -2149 0 1
rlabel polysilicon 177 -2155 177 -2155 0 3
rlabel polysilicon 180 -2155 180 -2155 0 4
rlabel polysilicon 184 -2155 184 -2155 0 3
rlabel polysilicon 187 -2155 187 -2155 0 4
rlabel polysilicon 191 -2149 191 -2149 0 1
rlabel polysilicon 191 -2155 191 -2155 0 3
rlabel polysilicon 198 -2149 198 -2149 0 1
rlabel polysilicon 198 -2155 198 -2155 0 3
rlabel polysilicon 205 -2149 205 -2149 0 1
rlabel polysilicon 205 -2155 205 -2155 0 3
rlabel polysilicon 215 -2149 215 -2149 0 2
rlabel polysilicon 212 -2155 212 -2155 0 3
rlabel polysilicon 222 -2149 222 -2149 0 2
rlabel polysilicon 219 -2155 219 -2155 0 3
rlabel polysilicon 226 -2149 226 -2149 0 1
rlabel polysilicon 226 -2155 226 -2155 0 3
rlabel polysilicon 233 -2149 233 -2149 0 1
rlabel polysilicon 233 -2155 233 -2155 0 3
rlabel polysilicon 240 -2149 240 -2149 0 1
rlabel polysilicon 240 -2155 240 -2155 0 3
rlabel polysilicon 247 -2149 247 -2149 0 1
rlabel polysilicon 247 -2155 247 -2155 0 3
rlabel polysilicon 254 -2149 254 -2149 0 1
rlabel polysilicon 261 -2149 261 -2149 0 1
rlabel polysilicon 264 -2149 264 -2149 0 2
rlabel polysilicon 268 -2149 268 -2149 0 1
rlabel polysilicon 268 -2155 268 -2155 0 3
rlabel polysilicon 275 -2149 275 -2149 0 1
rlabel polysilicon 275 -2155 275 -2155 0 3
rlabel polysilicon 282 -2155 282 -2155 0 3
rlabel polysilicon 289 -2149 289 -2149 0 1
rlabel polysilicon 292 -2149 292 -2149 0 2
rlabel polysilicon 292 -2155 292 -2155 0 4
rlabel polysilicon 296 -2149 296 -2149 0 1
rlabel polysilicon 296 -2155 296 -2155 0 3
rlabel polysilicon 303 -2149 303 -2149 0 1
rlabel polysilicon 306 -2149 306 -2149 0 2
rlabel polysilicon 303 -2155 303 -2155 0 3
rlabel polysilicon 310 -2149 310 -2149 0 1
rlabel polysilicon 310 -2155 310 -2155 0 3
rlabel polysilicon 317 -2155 317 -2155 0 3
rlabel polysilicon 324 -2149 324 -2149 0 1
rlabel polysilicon 324 -2155 324 -2155 0 3
rlabel polysilicon 334 -2149 334 -2149 0 2
rlabel polysilicon 334 -2155 334 -2155 0 4
rlabel polysilicon 338 -2149 338 -2149 0 1
rlabel polysilicon 338 -2155 338 -2155 0 3
rlabel polysilicon 345 -2149 345 -2149 0 1
rlabel polysilicon 345 -2155 345 -2155 0 3
rlabel polysilicon 352 -2149 352 -2149 0 1
rlabel polysilicon 352 -2155 352 -2155 0 3
rlabel polysilicon 359 -2155 359 -2155 0 3
rlabel polysilicon 362 -2155 362 -2155 0 4
rlabel polysilicon 366 -2149 366 -2149 0 1
rlabel polysilicon 366 -2155 366 -2155 0 3
rlabel polysilicon 373 -2149 373 -2149 0 1
rlabel polysilicon 380 -2149 380 -2149 0 1
rlabel polysilicon 380 -2155 380 -2155 0 3
rlabel polysilicon 387 -2149 387 -2149 0 1
rlabel polysilicon 387 -2155 387 -2155 0 3
rlabel polysilicon 394 -2149 394 -2149 0 1
rlabel polysilicon 394 -2155 394 -2155 0 3
rlabel polysilicon 401 -2149 401 -2149 0 1
rlabel polysilicon 401 -2155 401 -2155 0 3
rlabel polysilicon 408 -2149 408 -2149 0 1
rlabel polysilicon 408 -2155 408 -2155 0 3
rlabel polysilicon 415 -2155 415 -2155 0 3
rlabel polysilicon 422 -2149 422 -2149 0 1
rlabel polysilicon 422 -2155 422 -2155 0 3
rlabel polysilicon 429 -2149 429 -2149 0 1
rlabel polysilicon 429 -2155 429 -2155 0 3
rlabel polysilicon 436 -2149 436 -2149 0 1
rlabel polysilicon 436 -2155 436 -2155 0 3
rlabel polysilicon 443 -2149 443 -2149 0 1
rlabel polysilicon 443 -2155 443 -2155 0 3
rlabel polysilicon 450 -2149 450 -2149 0 1
rlabel polysilicon 450 -2155 450 -2155 0 3
rlabel polysilicon 457 -2149 457 -2149 0 1
rlabel polysilicon 457 -2155 457 -2155 0 3
rlabel polysilicon 467 -2155 467 -2155 0 4
rlabel polysilicon 471 -2149 471 -2149 0 1
rlabel polysilicon 471 -2155 471 -2155 0 3
rlabel polysilicon 478 -2149 478 -2149 0 1
rlabel polysilicon 478 -2155 478 -2155 0 3
rlabel polysilicon 485 -2149 485 -2149 0 1
rlabel polysilicon 485 -2155 485 -2155 0 3
rlabel polysilicon 492 -2149 492 -2149 0 1
rlabel polysilicon 492 -2155 492 -2155 0 3
rlabel polysilicon 499 -2155 499 -2155 0 3
rlabel polysilicon 509 -2149 509 -2149 0 2
rlabel polysilicon 509 -2155 509 -2155 0 4
rlabel polysilicon 513 -2149 513 -2149 0 1
rlabel polysilicon 513 -2155 513 -2155 0 3
rlabel polysilicon 523 -2149 523 -2149 0 2
rlabel polysilicon 530 -2149 530 -2149 0 2
rlabel polysilicon 534 -2149 534 -2149 0 1
rlabel polysilicon 534 -2155 534 -2155 0 3
rlabel polysilicon 541 -2149 541 -2149 0 1
rlabel polysilicon 541 -2155 541 -2155 0 3
rlabel polysilicon 548 -2149 548 -2149 0 1
rlabel polysilicon 548 -2155 548 -2155 0 3
rlabel polysilicon 555 -2149 555 -2149 0 1
rlabel polysilicon 555 -2155 555 -2155 0 3
rlabel polysilicon 562 -2149 562 -2149 0 1
rlabel polysilicon 562 -2155 562 -2155 0 3
rlabel polysilicon 569 -2149 569 -2149 0 1
rlabel polysilicon 569 -2155 569 -2155 0 3
rlabel polysilicon 590 -2149 590 -2149 0 1
rlabel polysilicon 590 -2155 590 -2155 0 3
rlabel polysilicon 597 -2149 597 -2149 0 1
rlabel polysilicon 597 -2155 597 -2155 0 3
rlabel polysilicon 611 -2149 611 -2149 0 1
rlabel polysilicon 611 -2155 611 -2155 0 3
rlabel polysilicon 9 -2196 9 -2196 0 1
rlabel polysilicon 9 -2202 9 -2202 0 3
rlabel polysilicon 19 -2196 19 -2196 0 2
rlabel polysilicon 23 -2202 23 -2202 0 3
rlabel polysilicon 40 -2196 40 -2196 0 2
rlabel polysilicon 44 -2202 44 -2202 0 3
rlabel polysilicon 51 -2196 51 -2196 0 1
rlabel polysilicon 51 -2202 51 -2202 0 3
rlabel polysilicon 58 -2196 58 -2196 0 1
rlabel polysilicon 58 -2202 58 -2202 0 3
rlabel polysilicon 65 -2196 65 -2196 0 1
rlabel polysilicon 65 -2202 65 -2202 0 3
rlabel polysilicon 72 -2196 72 -2196 0 1
rlabel polysilicon 72 -2202 72 -2202 0 3
rlabel polysilicon 79 -2196 79 -2196 0 1
rlabel polysilicon 79 -2202 79 -2202 0 3
rlabel polysilicon 86 -2196 86 -2196 0 1
rlabel polysilicon 86 -2202 86 -2202 0 3
rlabel polysilicon 93 -2196 93 -2196 0 1
rlabel polysilicon 93 -2202 93 -2202 0 3
rlabel polysilicon 100 -2196 100 -2196 0 1
rlabel polysilicon 100 -2202 100 -2202 0 3
rlabel polysilicon 107 -2196 107 -2196 0 1
rlabel polysilicon 107 -2202 107 -2202 0 3
rlabel polysilicon 114 -2202 114 -2202 0 3
rlabel polysilicon 121 -2196 121 -2196 0 1
rlabel polysilicon 121 -2202 121 -2202 0 3
rlabel polysilicon 128 -2196 128 -2196 0 1
rlabel polysilicon 131 -2196 131 -2196 0 2
rlabel polysilicon 128 -2202 128 -2202 0 3
rlabel polysilicon 135 -2196 135 -2196 0 1
rlabel polysilicon 138 -2196 138 -2196 0 2
rlabel polysilicon 145 -2202 145 -2202 0 4
rlabel polysilicon 149 -2196 149 -2196 0 1
rlabel polysilicon 149 -2202 149 -2202 0 3
rlabel polysilicon 156 -2196 156 -2196 0 1
rlabel polysilicon 156 -2202 156 -2202 0 3
rlabel polysilicon 163 -2196 163 -2196 0 1
rlabel polysilicon 163 -2202 163 -2202 0 3
rlabel polysilicon 170 -2196 170 -2196 0 1
rlabel polysilicon 170 -2202 170 -2202 0 3
rlabel polysilicon 177 -2196 177 -2196 0 1
rlabel polysilicon 177 -2202 177 -2202 0 3
rlabel polysilicon 187 -2196 187 -2196 0 2
rlabel polysilicon 191 -2196 191 -2196 0 1
rlabel polysilicon 191 -2202 191 -2202 0 3
rlabel polysilicon 198 -2196 198 -2196 0 1
rlabel polysilicon 201 -2202 201 -2202 0 4
rlabel polysilicon 208 -2196 208 -2196 0 2
rlabel polysilicon 205 -2202 205 -2202 0 3
rlabel polysilicon 212 -2196 212 -2196 0 1
rlabel polysilicon 215 -2196 215 -2196 0 2
rlabel polysilicon 219 -2196 219 -2196 0 1
rlabel polysilicon 219 -2202 219 -2202 0 3
rlabel polysilicon 226 -2196 226 -2196 0 1
rlabel polysilicon 226 -2202 226 -2202 0 3
rlabel polysilicon 233 -2196 233 -2196 0 1
rlabel polysilicon 247 -2196 247 -2196 0 1
rlabel polysilicon 247 -2202 247 -2202 0 3
rlabel polysilicon 257 -2196 257 -2196 0 2
rlabel polysilicon 254 -2202 254 -2202 0 3
rlabel polysilicon 261 -2196 261 -2196 0 1
rlabel polysilicon 261 -2202 261 -2202 0 3
rlabel polysilicon 268 -2196 268 -2196 0 1
rlabel polysilicon 268 -2202 268 -2202 0 3
rlabel polysilicon 278 -2196 278 -2196 0 2
rlabel polysilicon 285 -2196 285 -2196 0 2
rlabel polysilicon 289 -2196 289 -2196 0 1
rlabel polysilicon 289 -2202 289 -2202 0 3
rlabel polysilicon 296 -2196 296 -2196 0 1
rlabel polysilicon 299 -2202 299 -2202 0 4
rlabel polysilicon 303 -2196 303 -2196 0 1
rlabel polysilicon 303 -2202 303 -2202 0 3
rlabel polysilicon 317 -2196 317 -2196 0 1
rlabel polysilicon 317 -2202 317 -2202 0 3
rlabel polysilicon 324 -2196 324 -2196 0 1
rlabel polysilicon 324 -2202 324 -2202 0 3
rlabel polysilicon 331 -2196 331 -2196 0 1
rlabel polysilicon 331 -2202 331 -2202 0 3
rlabel polysilicon 345 -2196 345 -2196 0 1
rlabel polysilicon 348 -2196 348 -2196 0 2
rlabel polysilicon 345 -2202 345 -2202 0 3
rlabel polysilicon 352 -2196 352 -2196 0 1
rlabel polysilicon 352 -2202 352 -2202 0 3
rlabel polysilicon 359 -2202 359 -2202 0 3
rlabel polysilicon 362 -2202 362 -2202 0 4
rlabel polysilicon 366 -2202 366 -2202 0 3
rlabel polysilicon 373 -2196 373 -2196 0 1
rlabel polysilicon 380 -2196 380 -2196 0 1
rlabel polysilicon 380 -2202 380 -2202 0 3
rlabel polysilicon 387 -2196 387 -2196 0 1
rlabel polysilicon 387 -2202 387 -2202 0 3
rlabel polysilicon 394 -2196 394 -2196 0 1
rlabel polysilicon 394 -2202 394 -2202 0 3
rlabel polysilicon 401 -2196 401 -2196 0 1
rlabel polysilicon 401 -2202 401 -2202 0 3
rlabel polysilicon 408 -2196 408 -2196 0 1
rlabel polysilicon 408 -2202 408 -2202 0 3
rlabel polysilicon 415 -2196 415 -2196 0 1
rlabel polysilicon 418 -2202 418 -2202 0 4
rlabel polysilicon 425 -2196 425 -2196 0 2
rlabel polysilicon 422 -2202 422 -2202 0 3
rlabel polysilicon 429 -2196 429 -2196 0 1
rlabel polysilicon 429 -2202 429 -2202 0 3
rlabel polysilicon 436 -2196 436 -2196 0 1
rlabel polysilicon 436 -2202 436 -2202 0 3
rlabel polysilicon 443 -2196 443 -2196 0 1
rlabel polysilicon 443 -2202 443 -2202 0 3
rlabel polysilicon 453 -2196 453 -2196 0 2
rlabel polysilicon 457 -2196 457 -2196 0 1
rlabel polysilicon 457 -2202 457 -2202 0 3
rlabel polysilicon 464 -2196 464 -2196 0 1
rlabel polysilicon 464 -2202 464 -2202 0 3
rlabel polysilicon 481 -2196 481 -2196 0 2
rlabel polysilicon 492 -2196 492 -2196 0 1
rlabel polysilicon 492 -2202 492 -2202 0 3
rlabel polysilicon 499 -2196 499 -2196 0 1
rlabel polysilicon 520 -2196 520 -2196 0 1
rlabel polysilicon 520 -2202 520 -2202 0 3
rlabel polysilicon 534 -2196 534 -2196 0 1
rlabel polysilicon 534 -2202 534 -2202 0 3
rlabel polysilicon 548 -2202 548 -2202 0 3
rlabel polysilicon 555 -2196 555 -2196 0 1
rlabel polysilicon 555 -2202 555 -2202 0 3
rlabel polysilicon 600 -2196 600 -2196 0 2
rlabel polysilicon 600 -2202 600 -2202 0 4
rlabel polysilicon 604 -2196 604 -2196 0 1
rlabel polysilicon 604 -2202 604 -2202 0 3
rlabel polysilicon 611 -2196 611 -2196 0 1
rlabel polysilicon 611 -2202 611 -2202 0 3
rlabel polysilicon 16 -2225 16 -2225 0 1
rlabel polysilicon 26 -2225 26 -2225 0 2
rlabel polysilicon 44 -2225 44 -2225 0 1
rlabel polysilicon 51 -2225 51 -2225 0 1
rlabel polysilicon 58 -2225 58 -2225 0 1
rlabel polysilicon 58 -2231 58 -2231 0 3
rlabel polysilicon 75 -2231 75 -2231 0 4
rlabel polysilicon 82 -2225 82 -2225 0 2
rlabel polysilicon 93 -2231 93 -2231 0 3
rlabel polysilicon 103 -2225 103 -2225 0 2
rlabel polysilicon 107 -2225 107 -2225 0 1
rlabel polysilicon 107 -2231 107 -2231 0 3
rlabel polysilicon 114 -2225 114 -2225 0 1
rlabel polysilicon 114 -2231 114 -2231 0 3
rlabel polysilicon 131 -2231 131 -2231 0 4
rlabel polysilicon 149 -2225 149 -2225 0 1
rlabel polysilicon 149 -2231 149 -2231 0 3
rlabel polysilicon 163 -2231 163 -2231 0 3
rlabel polysilicon 173 -2231 173 -2231 0 4
rlabel polysilicon 177 -2225 177 -2225 0 1
rlabel polysilicon 187 -2225 187 -2225 0 2
rlabel polysilicon 191 -2225 191 -2225 0 1
rlabel polysilicon 201 -2231 201 -2231 0 4
rlabel polysilicon 205 -2225 205 -2225 0 1
rlabel polysilicon 208 -2225 208 -2225 0 2
rlabel polysilicon 212 -2225 212 -2225 0 1
rlabel polysilicon 219 -2231 219 -2231 0 3
rlabel polysilicon 226 -2225 226 -2225 0 1
rlabel polysilicon 226 -2231 226 -2231 0 3
rlabel polysilicon 240 -2225 240 -2225 0 1
rlabel polysilicon 240 -2231 240 -2231 0 3
rlabel polysilicon 247 -2225 247 -2225 0 1
rlabel polysilicon 247 -2231 247 -2231 0 3
rlabel polysilicon 254 -2225 254 -2225 0 1
rlabel polysilicon 254 -2231 254 -2231 0 3
rlabel polysilicon 268 -2225 268 -2225 0 1
rlabel polysilicon 268 -2231 268 -2231 0 3
rlabel polysilicon 275 -2225 275 -2225 0 1
rlabel polysilicon 275 -2231 275 -2231 0 3
rlabel polysilicon 282 -2225 282 -2225 0 1
rlabel polysilicon 282 -2231 282 -2231 0 3
rlabel polysilicon 289 -2225 289 -2225 0 1
rlabel polysilicon 289 -2231 289 -2231 0 3
rlabel polysilicon 303 -2231 303 -2231 0 3
rlabel polysilicon 310 -2231 310 -2231 0 3
rlabel polysilicon 313 -2231 313 -2231 0 4
rlabel polysilicon 327 -2225 327 -2225 0 2
rlabel polysilicon 327 -2231 327 -2231 0 4
rlabel polysilicon 331 -2225 331 -2225 0 1
rlabel polysilicon 331 -2231 331 -2231 0 3
rlabel polysilicon 341 -2225 341 -2225 0 2
rlabel polysilicon 348 -2225 348 -2225 0 2
rlabel polysilicon 355 -2231 355 -2231 0 4
rlabel polysilicon 373 -2225 373 -2225 0 1
rlabel polysilicon 373 -2231 373 -2231 0 3
rlabel polysilicon 383 -2231 383 -2231 0 4
rlabel polysilicon 390 -2231 390 -2231 0 4
rlabel polysilicon 408 -2225 408 -2225 0 1
rlabel polysilicon 408 -2231 408 -2231 0 3
rlabel polysilicon 429 -2231 429 -2231 0 3
rlabel polysilicon 450 -2225 450 -2225 0 1
rlabel polysilicon 450 -2231 450 -2231 0 3
rlabel polysilicon 474 -2231 474 -2231 0 4
rlabel polysilicon 485 -2231 485 -2231 0 3
rlabel polysilicon 506 -2225 506 -2225 0 1
rlabel polysilicon 506 -2231 506 -2231 0 3
rlabel polysilicon 534 -2225 534 -2225 0 1
rlabel polysilicon 537 -2225 537 -2225 0 2
rlabel polysilicon 611 -2225 611 -2225 0 1
rlabel metal2 131 1 131 1 0 net=3179
rlabel metal2 163 1 163 1 0 net=1303
rlabel metal2 191 1 191 1 0 net=5287
rlabel metal2 261 1 261 1 0 net=1883
rlabel metal2 177 -1 177 -1 0 net=4069
rlabel metal2 215 -1 215 -1 0 net=2799
rlabel metal2 268 -1 268 -1 0 net=3757
rlabel metal2 226 -3 226 -3 0 net=2525
rlabel metal2 26 -14 26 -14 0 net=652
rlabel metal2 26 -14 26 -14 0 net=652
rlabel metal2 86 -14 86 -14 0 net=1305
rlabel metal2 170 -14 170 -14 0 net=2793
rlabel metal2 240 -14 240 -14 0 net=1885
rlabel metal2 268 -14 268 -14 0 net=3759
rlabel metal2 369 -14 369 -14 0 net=4853
rlabel metal2 93 -16 93 -16 0 net=4153
rlabel metal2 107 -16 107 -16 0 net=896
rlabel metal2 142 -16 142 -16 0 net=2526
rlabel metal2 247 -16 247 -16 0 net=2801
rlabel metal2 327 -16 327 -16 0 net=4679
rlabel metal2 376 -16 376 -16 0 net=4267
rlabel metal2 110 -18 110 -18 0 net=2265
rlabel metal2 257 -18 257 -18 0 net=4463
rlabel metal2 138 -20 138 -20 0 net=2079
rlabel metal2 149 -20 149 -20 0 net=2093
rlabel metal2 170 -20 170 -20 0 net=4071
rlabel metal2 180 -20 180 -20 0 net=1031
rlabel metal2 243 -20 243 -20 0 net=1323
rlabel metal2 275 -20 275 -20 0 net=3405
rlabel metal2 156 -22 156 -22 0 net=3180
rlabel metal2 184 -22 184 -22 0 net=4979
rlabel metal2 215 -22 215 -22 0 net=3525
rlabel metal2 117 -24 117 -24 0 net=1001
rlabel metal2 191 -24 191 -24 0 net=5289
rlabel metal2 128 -26 128 -26 0 net=1359
rlabel metal2 198 -26 198 -26 0 net=3783
rlabel metal2 198 -28 198 -28 0 net=1437
rlabel metal2 222 -28 222 -28 0 net=3705
rlabel metal2 282 -28 282 -28 0 net=3831
rlabel metal2 205 -30 205 -30 0 net=2937
rlabel metal2 282 -30 282 -30 0 net=3557
rlabel metal2 65 -41 65 -41 0 net=4155
rlabel metal2 100 -41 100 -41 0 net=4980
rlabel metal2 212 -41 212 -41 0 net=3832
rlabel metal2 72 -43 72 -43 0 net=414
rlabel metal2 149 -43 149 -43 0 net=2094
rlabel metal2 184 -43 184 -43 0 net=1439
rlabel metal2 226 -43 226 -43 0 net=4237
rlabel metal2 75 -45 75 -45 0 net=3611
rlabel metal2 156 -45 156 -45 0 net=1002
rlabel metal2 229 -45 229 -45 0 net=3706
rlabel metal2 275 -45 275 -45 0 net=3407
rlabel metal2 282 -45 282 -45 0 net=4793
rlabel metal2 79 -47 79 -47 0 net=1409
rlabel metal2 233 -47 233 -47 0 net=1032
rlabel metal2 324 -47 324 -47 0 net=4464
rlabel metal2 86 -49 86 -49 0 net=1306
rlabel metal2 233 -49 233 -49 0 net=1887
rlabel metal2 261 -49 261 -49 0 net=2939
rlabel metal2 275 -49 275 -49 0 net=3558
rlabel metal2 44 -51 44 -51 0 net=4401
rlabel metal2 114 -51 114 -51 0 net=904
rlabel metal2 163 -51 163 -51 0 net=1003
rlabel metal2 240 -51 240 -51 0 net=1325
rlabel metal2 107 -53 107 -53 0 net=1077
rlabel metal2 117 -53 117 -53 0 net=735
rlabel metal2 191 -53 191 -53 0 net=1361
rlabel metal2 282 -53 282 -53 0 net=4268
rlabel metal2 121 -55 121 -55 0 net=816
rlabel metal2 205 -55 205 -55 0 net=4269
rlabel metal2 121 -57 121 -57 0 net=515
rlabel metal2 170 -57 170 -57 0 net=4073
rlabel metal2 131 -59 131 -59 0 net=4577
rlabel metal2 135 -61 135 -61 0 net=2081
rlabel metal2 170 -61 170 -61 0 net=4854
rlabel metal2 285 -63 285 -63 0 net=3760
rlabel metal2 289 -65 289 -65 0 net=2803
rlabel metal2 331 -65 331 -65 0 net=4681
rlabel metal2 219 -67 219 -67 0 net=2795
rlabel metal2 296 -67 296 -67 0 net=3527
rlabel metal2 338 -67 338 -67 0 net=3589
rlabel metal2 219 -69 219 -69 0 net=4371
rlabel metal2 254 -71 254 -71 0 net=2267
rlabel metal2 303 -71 303 -71 0 net=3785
rlabel metal2 303 -71 303 -71 0 net=3785
rlabel metal2 338 -71 338 -71 0 net=3915
rlabel metal2 51 -73 51 -73 0 net=1581
rlabel metal2 257 -73 257 -73 0 net=3643
rlabel metal2 352 -73 352 -73 0 net=5291
rlabel metal2 44 -84 44 -84 0 net=4402
rlabel metal2 121 -84 121 -84 0 net=2083
rlabel metal2 159 -84 159 -84 0 net=987
rlabel metal2 194 -84 194 -84 0 net=1803
rlabel metal2 250 -84 250 -84 0 net=4682
rlabel metal2 51 -86 51 -86 0 net=1582
rlabel metal2 163 -86 163 -86 0 net=1005
rlabel metal2 201 -86 201 -86 0 net=1362
rlabel metal2 254 -86 254 -86 0 net=3786
rlabel metal2 331 -86 331 -86 0 net=3644
rlabel metal2 394 -86 394 -86 0 net=5293
rlabel metal2 58 -88 58 -88 0 net=1835
rlabel metal2 205 -88 205 -88 0 net=1327
rlabel metal2 257 -88 257 -88 0 net=4238
rlabel metal2 401 -88 401 -88 0 net=4707
rlabel metal2 65 -90 65 -90 0 net=4156
rlabel metal2 128 -90 128 -90 0 net=1983
rlabel metal2 65 -92 65 -92 0 net=1410
rlabel metal2 86 -92 86 -92 0 net=1079
rlabel metal2 131 -92 131 -92 0 net=2796
rlabel metal2 317 -92 317 -92 0 net=3409
rlabel metal2 352 -92 352 -92 0 net=4794
rlabel metal2 93 -94 93 -94 0 net=1821
rlabel metal2 142 -94 142 -94 0 net=176
rlabel metal2 212 -94 212 -94 0 net=2940
rlabel metal2 271 -94 271 -94 0 net=4578
rlabel metal2 408 -94 408 -94 0 net=4087
rlabel metal2 107 -96 107 -96 0 net=2485
rlabel metal2 275 -96 275 -96 0 net=2837
rlabel metal2 289 -96 289 -96 0 net=4075
rlabel metal2 366 -96 366 -96 0 net=4373
rlabel metal2 96 -98 96 -98 0 net=3545
rlabel metal2 149 -100 149 -100 0 net=3613
rlabel metal2 149 -102 149 -102 0 net=1441
rlabel metal2 212 -102 212 -102 0 net=409
rlabel metal2 222 -102 222 -102 0 net=4495
rlabel metal2 177 -104 177 -104 0 net=2167
rlabel metal2 278 -104 278 -104 0 net=4270
rlabel metal2 184 -106 184 -106 0 net=2191
rlabel metal2 215 -106 215 -106 0 net=3528
rlabel metal2 338 -106 338 -106 0 net=3917
rlabel metal2 79 -108 79 -108 0 net=2061
rlabel metal2 233 -108 233 -108 0 net=1889
rlabel metal2 271 -108 271 -108 0 net=1949
rlabel metal2 345 -108 345 -108 0 net=3591
rlabel metal2 198 -110 198 -110 0 net=2989
rlabel metal2 240 -112 240 -112 0 net=4511
rlabel metal2 278 -114 278 -114 0 net=2931
rlabel metal2 310 -114 310 -114 0 net=2805
rlabel metal2 296 -116 296 -116 0 net=2269
rlabel metal2 296 -118 296 -118 0 net=4117
rlabel metal2 37 -129 37 -129 0 net=1443
rlabel metal2 156 -129 156 -129 0 net=1339
rlabel metal2 215 -129 215 -129 0 net=4512
rlabel metal2 436 -129 436 -129 0 net=4497
rlabel metal2 44 -131 44 -131 0 net=1823
rlabel metal2 110 -131 110 -131 0 net=1733
rlabel metal2 128 -131 128 -131 0 net=1329
rlabel metal2 219 -131 219 -131 0 net=1217
rlabel metal2 226 -131 226 -131 0 net=1804
rlabel metal2 254 -131 254 -131 0 net=1891
rlabel metal2 275 -131 275 -131 0 net=4669
rlabel metal2 51 -133 51 -133 0 net=3123
rlabel metal2 170 -133 170 -133 0 net=1007
rlabel metal2 58 -135 58 -135 0 net=1836
rlabel metal2 145 -135 145 -135 0 net=4419
rlabel metal2 233 -135 233 -135 0 net=307
rlabel metal2 247 -135 247 -135 0 net=1950
rlabel metal2 359 -135 359 -135 0 net=3547
rlabel metal2 380 -135 380 -135 0 net=4795
rlabel metal2 58 -137 58 -137 0 net=4965
rlabel metal2 170 -137 170 -137 0 net=2193
rlabel metal2 236 -137 236 -137 0 net=4374
rlabel metal2 72 -139 72 -139 0 net=2085
rlabel metal2 131 -139 131 -139 0 net=4496
rlabel metal2 79 -141 79 -141 0 net=2062
rlabel metal2 177 -141 177 -141 0 net=2169
rlabel metal2 254 -141 254 -141 0 net=4721
rlabel metal2 79 -143 79 -143 0 net=4121
rlabel metal2 184 -143 184 -143 0 net=1867
rlabel metal2 261 -143 261 -143 0 net=1497
rlabel metal2 289 -143 289 -143 0 net=4077
rlabel metal2 387 -143 387 -143 0 net=3919
rlabel metal2 89 -145 89 -145 0 net=225
rlabel metal2 103 -145 103 -145 0 net=239
rlabel metal2 191 -145 191 -145 0 net=2807
rlabel metal2 352 -145 352 -145 0 net=3593
rlabel metal2 401 -145 401 -145 0 net=4709
rlabel metal2 100 -147 100 -147 0 net=2487
rlabel metal2 117 -147 117 -147 0 net=3399
rlabel metal2 345 -147 345 -147 0 net=2991
rlabel metal2 415 -147 415 -147 0 net=5295
rlabel metal2 138 -149 138 -149 0 net=747
rlabel metal2 208 -149 208 -149 0 net=4239
rlabel metal2 86 -151 86 -151 0 net=1080
rlabel metal2 282 -151 282 -151 0 net=2839
rlabel metal2 296 -153 296 -153 0 net=4118
rlabel metal2 317 -153 317 -153 0 net=2271
rlabel metal2 296 -155 296 -155 0 net=3095
rlabel metal2 303 -157 303 -157 0 net=2933
rlabel metal2 306 -159 306 -159 0 net=4617
rlabel metal2 310 -161 310 -161 0 net=4088
rlabel metal2 317 -163 317 -163 0 net=5053
rlabel metal2 320 -165 320 -165 0 net=1984
rlabel metal2 373 -167 373 -167 0 net=3615
rlabel metal2 331 -169 331 -169 0 net=3411
rlabel metal2 331 -171 331 -171 0 net=615
rlabel metal2 16 -182 16 -182 0 net=4387
rlabel metal2 100 -182 100 -182 0 net=2488
rlabel metal2 100 -182 100 -182 0 net=2488
rlabel metal2 114 -182 114 -182 0 net=1734
rlabel metal2 191 -182 191 -182 0 net=2808
rlabel metal2 292 -182 292 -182 0 net=3412
rlabel metal2 380 -182 380 -182 0 net=4078
rlabel metal2 583 -182 583 -182 0 net=5427
rlabel metal2 30 -184 30 -184 0 net=1065
rlabel metal2 226 -184 226 -184 0 net=4421
rlabel metal2 534 -184 534 -184 0 net=5103
rlabel metal2 37 -186 37 -186 0 net=1444
rlabel metal2 212 -186 212 -186 0 net=169
rlabel metal2 212 -186 212 -186 0 net=169
rlabel metal2 254 -186 254 -186 0 net=363
rlabel metal2 380 -186 380 -186 0 net=3391
rlabel metal2 37 -188 37 -188 0 net=4122
rlabel metal2 86 -188 86 -188 0 net=1527
rlabel metal2 114 -188 114 -188 0 net=2969
rlabel metal2 387 -188 387 -188 0 net=3096
rlabel metal2 44 -190 44 -190 0 net=1824
rlabel metal2 191 -190 191 -190 0 net=1485
rlabel metal2 257 -190 257 -190 0 net=1892
rlabel metal2 275 -190 275 -190 0 net=2841
rlabel metal2 366 -190 366 -190 0 net=3549
rlabel metal2 464 -190 464 -190 0 net=4723
rlabel metal2 51 -192 51 -192 0 net=3124
rlabel metal2 296 -192 296 -192 0 net=3400
rlabel metal2 450 -192 450 -192 0 net=4671
rlabel metal2 471 -192 471 -192 0 net=4797
rlabel metal2 58 -194 58 -194 0 net=4967
rlabel metal2 58 -196 58 -196 0 net=1115
rlabel metal2 121 -196 121 -196 0 net=1868
rlabel metal2 261 -196 261 -196 0 net=1499
rlabel metal2 306 -196 306 -196 0 net=3920
rlabel metal2 65 -198 65 -198 0 net=664
rlabel metal2 72 -198 72 -198 0 net=2086
rlabel metal2 156 -198 156 -198 0 net=1341
rlabel metal2 278 -198 278 -198 0 net=1008
rlabel metal2 443 -198 443 -198 0 net=4619
rlabel metal2 457 -198 457 -198 0 net=4711
rlabel metal2 79 -200 79 -200 0 net=4253
rlabel metal2 436 -200 436 -200 0 net=4499
rlabel metal2 89 -202 89 -202 0 net=5296
rlabel metal2 103 -204 103 -204 0 net=4299
rlabel metal2 121 -206 121 -206 0 net=3961
rlabel metal2 408 -206 408 -206 0 net=5055
rlabel metal2 124 -208 124 -208 0 net=876
rlabel metal2 243 -208 243 -208 0 net=1239
rlabel metal2 282 -208 282 -208 0 net=4049
rlabel metal2 128 -210 128 -210 0 net=1331
rlabel metal2 187 -210 187 -210 0 net=3879
rlabel metal2 408 -210 408 -210 0 net=4021
rlabel metal2 82 -212 82 -212 0 net=2691
rlabel metal2 135 -212 135 -212 0 net=152
rlabel metal2 317 -212 317 -212 0 net=2273
rlabel metal2 135 -214 135 -214 0 net=2029
rlabel metal2 170 -214 170 -214 0 net=2195
rlabel metal2 324 -214 324 -214 0 net=4815
rlabel metal2 142 -216 142 -216 0 net=1375
rlabel metal2 233 -216 233 -216 0 net=2935
rlabel metal2 401 -216 401 -216 0 net=4241
rlabel metal2 96 -218 96 -218 0 net=4645
rlabel metal2 142 -220 142 -220 0 net=2475
rlabel metal2 331 -220 331 -220 0 net=4885
rlabel metal2 170 -222 170 -222 0 net=2007
rlabel metal2 198 -222 198 -222 0 net=2170
rlabel metal2 310 -222 310 -222 0 net=3351
rlabel metal2 345 -222 345 -222 0 net=3617
rlabel metal2 156 -224 156 -224 0 net=1119
rlabel metal2 198 -224 198 -224 0 net=2993
rlabel metal2 359 -224 359 -224 0 net=3595
rlabel metal2 205 -226 205 -226 0 net=1219
rlabel metal2 359 -226 359 -226 0 net=4683
rlabel metal2 149 -228 149 -228 0 net=463
rlabel metal2 16 -239 16 -239 0 net=4388
rlabel metal2 180 -239 180 -239 0 net=2196
rlabel metal2 285 -239 285 -239 0 net=4242
rlabel metal2 499 -239 499 -239 0 net=4725
rlabel metal2 586 -239 586 -239 0 net=5327
rlabel metal2 639 -239 639 -239 0 net=5429
rlabel metal2 30 -241 30 -241 0 net=1066
rlabel metal2 184 -241 184 -241 0 net=1333
rlabel metal2 184 -241 184 -241 0 net=1333
rlabel metal2 205 -241 205 -241 0 net=1220
rlabel metal2 240 -241 240 -241 0 net=5059
rlabel metal2 653 -241 653 -241 0 net=5331
rlabel metal2 653 -241 653 -241 0 net=5331
rlabel metal2 30 -243 30 -243 0 net=2995
rlabel metal2 205 -243 205 -243 0 net=1507
rlabel metal2 243 -243 243 -243 0 net=2842
rlabel metal2 278 -243 278 -243 0 net=3997
rlabel metal2 506 -243 506 -243 0 net=4799
rlabel metal2 44 -245 44 -245 0 net=1943
rlabel metal2 82 -245 82 -245 0 net=4422
rlabel metal2 481 -245 481 -245 0 net=4823
rlabel metal2 51 -247 51 -247 0 net=4968
rlabel metal2 534 -247 534 -247 0 net=5104
rlabel metal2 58 -249 58 -249 0 net=1117
rlabel metal2 103 -249 103 -249 0 net=3618
rlabel metal2 352 -249 352 -249 0 net=4886
rlabel metal2 513 -249 513 -249 0 net=4817
rlabel metal2 72 -251 72 -251 0 net=2031
rlabel metal2 156 -251 156 -251 0 net=2483
rlabel metal2 362 -251 362 -251 0 net=4646
rlabel metal2 408 -251 408 -251 0 net=4023
rlabel metal2 555 -251 555 -251 0 net=4929
rlabel metal2 86 -253 86 -253 0 net=2365
rlabel metal2 198 -253 198 -253 0 net=2491
rlabel metal2 366 -253 366 -253 0 net=3881
rlabel metal2 558 -253 558 -253 0 net=5243
rlabel metal2 93 -255 93 -255 0 net=1427
rlabel metal2 124 -255 124 -255 0 net=2709
rlabel metal2 156 -255 156 -255 0 net=1121
rlabel metal2 212 -255 212 -255 0 net=1376
rlabel metal2 247 -255 247 -255 0 net=5165
rlabel metal2 422 -255 422 -255 0 net=4255
rlabel metal2 100 -257 100 -257 0 net=3847
rlabel metal2 226 -257 226 -257 0 net=3447
rlabel metal2 268 -257 268 -257 0 net=1240
rlabel metal2 285 -257 285 -257 0 net=5395
rlabel metal2 254 -259 254 -259 0 net=3681
rlabel metal2 429 -259 429 -259 0 net=4301
rlabel metal2 268 -261 268 -261 0 net=2543
rlabel metal2 331 -261 331 -261 0 net=3353
rlabel metal2 233 -263 233 -263 0 net=2936
rlabel metal2 338 -263 338 -263 0 net=4217
rlabel metal2 289 -265 289 -265 0 net=1500
rlabel metal2 303 -265 303 -265 0 net=2477
rlabel metal2 380 -265 380 -265 0 net=3392
rlabel metal2 443 -265 443 -265 0 net=4501
rlabel metal2 114 -267 114 -267 0 net=2971
rlabel metal2 310 -267 310 -267 0 net=3009
rlabel metal2 415 -267 415 -267 0 net=4051
rlabel metal2 457 -267 457 -267 0 net=5057
rlabel metal2 114 -269 114 -269 0 net=1343
rlabel metal2 282 -269 282 -269 0 net=3509
rlabel metal2 457 -269 457 -269 0 net=4673
rlabel metal2 471 -269 471 -269 0 net=4713
rlabel metal2 128 -271 128 -271 0 net=2693
rlabel metal2 387 -271 387 -271 0 net=3551
rlabel metal2 107 -273 107 -273 0 net=1529
rlabel metal2 152 -273 152 -273 0 net=2095
rlabel metal2 299 -273 299 -273 0 net=3087
rlabel metal2 107 -275 107 -275 0 net=1487
rlabel metal2 222 -275 222 -275 0 net=3749
rlabel metal2 152 -277 152 -277 0 net=257
rlabel metal2 170 -277 170 -277 0 net=2009
rlabel metal2 313 -277 313 -277 0 net=979
rlabel metal2 40 -279 40 -279 0 net=2671
rlabel metal2 317 -279 317 -279 0 net=2275
rlabel metal2 366 -279 366 -279 0 net=2623
rlabel metal2 394 -279 394 -279 0 net=3597
rlabel metal2 215 -281 215 -281 0 net=2955
rlabel metal2 450 -281 450 -281 0 net=4621
rlabel metal2 215 -283 215 -283 0 net=1503
rlabel metal2 373 -283 373 -283 0 net=3963
rlabel metal2 163 -285 163 -285 0 net=1629
rlabel metal2 436 -285 436 -285 0 net=4685
rlabel metal2 9 -296 9 -296 0 net=2707
rlabel metal2 320 -296 320 -296 0 net=4302
rlabel metal2 653 -296 653 -296 0 net=5332
rlabel metal2 660 -296 660 -296 0 net=5431
rlabel metal2 30 -298 30 -298 0 net=2996
rlabel metal2 191 -298 191 -298 0 net=2694
rlabel metal2 387 -298 387 -298 0 net=4714
rlabel metal2 653 -298 653 -298 0 net=4455
rlabel metal2 30 -300 30 -300 0 net=2689
rlabel metal2 247 -300 247 -300 0 net=2484
rlabel metal2 359 -300 359 -300 0 net=5058
rlabel metal2 44 -302 44 -302 0 net=1944
rlabel metal2 247 -302 247 -302 0 net=1735
rlabel metal2 310 -302 310 -302 0 net=4024
rlabel metal2 534 -302 534 -302 0 net=4801
rlabel metal2 569 -302 569 -302 0 net=5061
rlabel metal2 611 -302 611 -302 0 net=5397
rlabel metal2 51 -304 51 -304 0 net=2745
rlabel metal2 215 -304 215 -304 0 net=3882
rlabel metal2 506 -304 506 -304 0 net=4219
rlabel metal2 562 -304 562 -304 0 net=4931
rlabel metal2 604 -304 604 -304 0 net=5245
rlabel metal2 58 -306 58 -306 0 net=1118
rlabel metal2 156 -306 156 -306 0 net=1122
rlabel metal2 191 -306 191 -306 0 net=3448
rlabel metal2 254 -306 254 -306 0 net=3354
rlabel metal2 597 -306 597 -306 0 net=5329
rlabel metal2 65 -308 65 -308 0 net=2544
rlabel metal2 289 -308 289 -308 0 net=2973
rlabel metal2 79 -310 79 -310 0 net=2956
rlabel metal2 401 -310 401 -310 0 net=3011
rlabel metal2 429 -310 429 -310 0 net=4053
rlabel metal2 79 -312 79 -312 0 net=2711
rlabel metal2 170 -312 170 -312 0 net=2673
rlabel metal2 289 -312 289 -312 0 net=1863
rlabel metal2 401 -312 401 -312 0 net=3683
rlabel metal2 432 -312 432 -312 0 net=4726
rlabel metal2 23 -314 23 -314 0 net=4969
rlabel metal2 205 -314 205 -314 0 net=1504
rlabel metal2 240 -314 240 -314 0 net=1509
rlabel metal2 257 -314 257 -314 0 net=2010
rlabel metal2 310 -314 310 -314 0 net=2625
rlabel metal2 373 -314 373 -314 0 net=1630
rlabel metal2 408 -314 408 -314 0 net=5167
rlabel metal2 86 -316 86 -316 0 net=2366
rlabel metal2 313 -316 313 -316 0 net=4256
rlabel metal2 86 -318 86 -318 0 net=1831
rlabel metal2 317 -318 317 -318 0 net=2479
rlabel metal2 352 -318 352 -318 0 net=3552
rlabel metal2 26 -320 26 -320 0 net=3311
rlabel metal2 373 -320 373 -320 0 net=3965
rlabel metal2 478 -320 478 -320 0 net=3999
rlabel metal2 527 -320 527 -320 0 net=4825
rlabel metal2 93 -322 93 -322 0 net=1429
rlabel metal2 331 -322 331 -322 0 net=5149
rlabel metal2 93 -324 93 -324 0 net=1805
rlabel metal2 261 -324 261 -324 0 net=2097
rlabel metal2 338 -324 338 -324 0 net=3598
rlabel metal2 100 -326 100 -326 0 net=3848
rlabel metal2 324 -326 324 -326 0 net=2277
rlabel metal2 341 -326 341 -326 0 net=2833
rlabel metal2 408 -326 408 -326 0 net=4623
rlabel metal2 548 -326 548 -326 0 net=4839
rlabel metal2 100 -328 100 -328 0 net=2089
rlabel metal2 415 -328 415 -328 0 net=3089
rlabel metal2 436 -328 436 -328 0 net=5183
rlabel metal2 110 -330 110 -330 0 net=731
rlabel metal2 222 -330 222 -330 0 net=2917
rlabel metal2 457 -330 457 -330 0 net=4675
rlabel metal2 492 -330 492 -330 0 net=4503
rlabel metal2 541 -330 541 -330 0 net=4819
rlabel metal2 72 -332 72 -332 0 net=2032
rlabel metal2 222 -332 222 -332 0 net=266
rlabel metal2 450 -332 450 -332 0 net=4687
rlabel metal2 72 -334 72 -334 0 net=2493
rlabel metal2 362 -334 362 -334 0 net=760
rlabel metal2 457 -334 457 -334 0 net=3751
rlabel metal2 107 -336 107 -336 0 net=1489
rlabel metal2 299 -336 299 -336 0 net=3909
rlabel metal2 107 -338 107 -338 0 net=3439
rlabel metal2 114 -340 114 -340 0 net=1344
rlabel metal2 299 -340 299 -340 0 net=3510
rlabel metal2 114 -342 114 -342 0 net=2423
rlabel metal2 443 -342 443 -342 0 net=3467
rlabel metal2 121 -344 121 -344 0 net=233
rlabel metal2 166 -344 166 -344 0 net=5201
rlabel metal2 128 -346 128 -346 0 net=1531
rlabel metal2 135 -348 135 -348 0 net=1355
rlabel metal2 58 -350 58 -350 0 net=2283
rlabel metal2 142 -352 142 -352 0 net=1335
rlabel metal2 128 -354 128 -354 0 net=1903
rlabel metal2 9 -365 9 -365 0 net=2708
rlabel metal2 128 -365 128 -365 0 net=1904
rlabel metal2 324 -365 324 -365 0 net=5063
rlabel metal2 653 -365 653 -365 0 net=64
rlabel metal2 674 -365 674 -365 0 net=5433
rlabel metal2 16 -367 16 -367 0 net=1337
rlabel metal2 170 -367 170 -367 0 net=3440
rlabel metal2 453 -367 453 -367 0 net=5062
rlabel metal2 583 -367 583 -367 0 net=5203
rlabel metal2 660 -367 660 -367 0 net=4456
rlabel metal2 23 -369 23 -369 0 net=4970
rlabel metal2 128 -369 128 -369 0 net=1405
rlabel metal2 219 -369 219 -369 0 net=3927
rlabel metal2 520 -369 520 -369 0 net=4689
rlabel metal2 30 -371 30 -371 0 net=2690
rlabel metal2 341 -371 341 -371 0 net=3684
rlabel metal2 408 -371 408 -371 0 net=4625
rlabel metal2 583 -371 583 -371 0 net=5399
rlabel metal2 44 -373 44 -373 0 net=3731
rlabel metal2 212 -373 212 -373 0 net=2747
rlabel metal2 429 -373 429 -373 0 net=4889
rlabel metal2 51 -375 51 -375 0 net=3623
rlabel metal2 229 -375 229 -375 0 net=4971
rlabel metal2 58 -377 58 -377 0 net=2284
rlabel metal2 359 -377 359 -377 0 net=4504
rlabel metal2 506 -377 506 -377 0 net=4221
rlabel metal2 548 -377 548 -377 0 net=4841
rlabel metal2 33 -379 33 -379 0 net=4517
rlabel metal2 555 -379 555 -379 0 net=5151
rlabel metal2 72 -381 72 -381 0 net=2494
rlabel metal2 177 -381 177 -381 0 net=272
rlabel metal2 254 -381 254 -381 0 net=1511
rlabel metal2 366 -381 366 -381 0 net=3752
rlabel metal2 464 -381 464 -381 0 net=3911
rlabel metal2 562 -381 562 -381 0 net=4933
rlabel metal2 72 -383 72 -383 0 net=1833
rlabel metal2 100 -383 100 -383 0 net=1557
rlabel metal2 275 -383 275 -383 0 net=3966
rlabel metal2 383 -383 383 -383 0 net=5168
rlabel metal2 604 -383 604 -383 0 net=5247
rlabel metal2 65 -385 65 -385 0 net=1713
rlabel metal2 275 -385 275 -385 0 net=2425
rlabel metal2 345 -385 345 -385 0 net=3313
rlabel metal2 471 -385 471 -385 0 net=4677
rlabel metal2 79 -387 79 -387 0 net=2712
rlabel metal2 240 -387 240 -387 0 net=1533
rlabel metal2 338 -387 338 -387 0 net=2279
rlabel metal2 352 -387 352 -387 0 net=3443
rlabel metal2 478 -387 478 -387 0 net=4001
rlabel metal2 527 -387 527 -387 0 net=4827
rlabel metal2 86 -389 86 -389 0 net=1231
rlabel metal2 282 -389 282 -389 0 net=2027
rlabel metal2 383 -389 383 -389 0 net=4325
rlabel metal2 93 -391 93 -391 0 net=1806
rlabel metal2 261 -391 261 -391 0 net=2918
rlabel metal2 289 -391 289 -391 0 net=1865
rlabel metal2 387 -391 387 -391 0 net=4611
rlabel metal2 481 -391 481 -391 0 net=5184
rlabel metal2 93 -393 93 -393 0 net=1419
rlabel metal2 198 -393 198 -393 0 net=1491
rlabel metal2 331 -393 331 -393 0 net=2099
rlabel metal2 355 -393 355 -393 0 net=4693
rlabel metal2 107 -395 107 -395 0 net=943
rlabel metal2 233 -395 233 -395 0 net=1431
rlabel metal2 310 -395 310 -395 0 net=2627
rlabel metal2 362 -395 362 -395 0 net=3341
rlabel metal2 107 -397 107 -397 0 net=2347
rlabel metal2 317 -397 317 -397 0 net=2480
rlabel metal2 390 -397 390 -397 0 net=5330
rlabel metal2 114 -399 114 -399 0 net=4563
rlabel metal2 121 -401 121 -401 0 net=1129
rlabel metal2 401 -401 401 -401 0 net=3013
rlabel metal2 422 -401 422 -401 0 net=3091
rlabel metal2 436 -401 436 -401 0 net=3469
rlabel metal2 534 -401 534 -401 0 net=4803
rlabel metal2 135 -403 135 -403 0 net=1356
rlabel metal2 268 -403 268 -403 0 net=2675
rlabel metal2 135 -405 135 -405 0 net=1221
rlabel metal2 170 -405 170 -405 0 net=168
rlabel metal2 317 -405 317 -405 0 net=2974
rlabel metal2 138 -407 138 -407 0 net=264
rlabel metal2 387 -407 387 -407 0 net=4457
rlabel metal2 142 -409 142 -409 0 net=1191
rlabel metal2 226 -409 226 -409 0 net=2091
rlabel metal2 394 -409 394 -409 0 net=2835
rlabel metal2 485 -409 485 -409 0 net=4055
rlabel metal2 117 -411 117 -411 0 net=3825
rlabel metal2 149 -413 149 -413 0 net=496
rlabel metal2 247 -413 247 -413 0 net=1737
rlabel metal2 149 -415 149 -415 0 net=1657
rlabel metal2 247 -415 247 -415 0 net=3337
rlabel metal2 184 -417 184 -417 0 net=1445
rlabel metal2 191 -419 191 -419 0 net=4820
rlabel metal2 474 -421 474 -421 0 net=4479
rlabel metal2 16 -432 16 -432 0 net=1338
rlabel metal2 257 -432 257 -432 0 net=2028
rlabel metal2 380 -432 380 -432 0 net=4056
rlabel metal2 541 -432 541 -432 0 net=4481
rlabel metal2 583 -432 583 -432 0 net=5401
rlabel metal2 33 -434 33 -434 0 net=1192
rlabel metal2 149 -434 149 -434 0 net=1658
rlabel metal2 201 -434 201 -434 0 net=3342
rlabel metal2 646 -434 646 -434 0 net=5153
rlabel metal2 681 -434 681 -434 0 net=5435
rlabel metal2 681 -434 681 -434 0 net=5435
rlabel metal2 40 -436 40 -436 0 net=738
rlabel metal2 219 -436 219 -436 0 net=4518
rlabel metal2 653 -436 653 -436 0 net=5205
rlabel metal2 44 -438 44 -438 0 net=3733
rlabel metal2 527 -438 527 -438 0 net=4327
rlabel metal2 639 -438 639 -438 0 net=5065
rlabel metal2 44 -440 44 -440 0 net=1223
rlabel metal2 205 -440 205 -440 0 net=3314
rlabel metal2 471 -440 471 -440 0 net=4934
rlabel metal2 632 -440 632 -440 0 net=4973
rlabel metal2 51 -442 51 -442 0 net=3624
rlabel metal2 390 -442 390 -442 0 net=4678
rlabel metal2 611 -442 611 -442 0 net=4843
rlabel metal2 58 -444 58 -444 0 net=1513
rlabel metal2 320 -444 320 -444 0 net=3092
rlabel metal2 450 -444 450 -444 0 net=4613
rlabel metal2 618 -444 618 -444 0 net=4891
rlabel metal2 65 -446 65 -446 0 net=1715
rlabel metal2 222 -446 222 -446 0 net=4103
rlabel metal2 65 -448 65 -448 0 net=2017
rlabel metal2 352 -448 352 -448 0 net=2101
rlabel metal2 390 -448 390 -448 0 net=4690
rlabel metal2 72 -450 72 -450 0 net=1834
rlabel metal2 177 -450 177 -450 0 net=5093
rlabel metal2 72 -452 72 -452 0 net=2033
rlabel metal2 229 -452 229 -452 0 net=1492
rlabel metal2 257 -452 257 -452 0 net=2919
rlabel metal2 478 -452 478 -452 0 net=5013
rlabel metal2 79 -454 79 -454 0 net=1131
rlabel metal2 128 -454 128 -454 0 net=1407
rlabel metal2 135 -454 135 -454 0 net=2285
rlabel metal2 264 -454 264 -454 0 net=2836
rlabel metal2 425 -454 425 -454 0 net=4694
rlabel metal2 82 -456 82 -456 0 net=1133
rlabel metal2 156 -456 156 -456 0 net=1535
rlabel metal2 331 -456 331 -456 0 net=2629
rlabel metal2 439 -456 439 -456 0 net=3807
rlabel metal2 485 -456 485 -456 0 net=3827
rlabel metal2 534 -456 534 -456 0 net=4459
rlabel metal2 93 -458 93 -458 0 net=1421
rlabel metal2 177 -458 177 -458 0 net=2891
rlabel metal2 345 -458 345 -458 0 net=2281
rlabel metal2 401 -458 401 -458 0 net=3015
rlabel metal2 492 -458 492 -458 0 net=3913
rlabel metal2 541 -458 541 -458 0 net=4805
rlabel metal2 100 -460 100 -460 0 net=1559
rlabel metal2 338 -460 338 -460 0 net=2749
rlabel metal2 443 -460 443 -460 0 net=3339
rlabel metal2 499 -460 499 -460 0 net=3929
rlabel metal2 100 -462 100 -462 0 net=4029
rlabel metal2 215 -462 215 -462 0 net=2503
rlabel metal2 436 -462 436 -462 0 net=3471
rlabel metal2 520 -462 520 -462 0 net=4223
rlabel metal2 107 -464 107 -464 0 net=2348
rlabel metal2 275 -464 275 -464 0 net=2427
rlabel metal2 61 -466 61 -466 0 net=326
rlabel metal2 310 -466 310 -466 0 net=2489
rlabel metal2 450 -466 450 -466 0 net=5161
rlabel metal2 110 -468 110 -468 0 net=2773
rlabel metal2 457 -468 457 -468 0 net=3445
rlabel metal2 114 -470 114 -470 0 net=4626
rlabel metal2 114 -472 114 -472 0 net=1011
rlabel metal2 117 -474 117 -474 0 net=1866
rlabel metal2 128 -476 128 -476 0 net=1433
rlabel metal2 327 -476 327 -476 0 net=2179
rlabel metal2 184 -478 184 -478 0 net=1447
rlabel metal2 355 -478 355 -478 0 net=4123
rlabel metal2 86 -480 86 -480 0 net=1233
rlabel metal2 191 -480 191 -480 0 net=2137
rlabel metal2 359 -480 359 -480 0 net=4002
rlabel metal2 544 -480 544 -480 0 net=1
rlabel metal2 86 -482 86 -482 0 net=1269
rlabel metal2 194 -482 194 -482 0 net=3647
rlabel metal2 215 -484 215 -484 0 net=2676
rlabel metal2 226 -486 226 -486 0 net=2905
rlabel metal2 226 -488 226 -488 0 net=2092
rlabel metal2 359 -488 359 -488 0 net=4828
rlabel metal2 229 -490 229 -490 0 net=256
rlabel metal2 268 -490 268 -490 0 net=2451
rlabel metal2 422 -490 422 -490 0 net=4025
rlabel metal2 555 -490 555 -490 0 net=4565
rlabel metal2 37 -492 37 -492 0 net=1075
rlabel metal2 233 -494 233 -494 0 net=248
rlabel metal2 233 -496 233 -496 0 net=1049
rlabel metal2 240 -498 240 -498 0 net=1738
rlabel metal2 247 -500 247 -500 0 net=2547
rlabel metal2 387 -500 387 -500 0 net=3017
rlabel metal2 261 -502 261 -502 0 net=1181
rlabel metal2 317 -504 317 -504 0 net=5248
rlabel metal2 282 -506 282 -506 0 net=5087
rlabel metal2 282 -508 282 -508 0 net=5333
rlabel metal2 16 -519 16 -519 0 net=882
rlabel metal2 348 -519 348 -519 0 net=4614
rlabel metal2 23 -521 23 -521 0 net=3473
rlabel metal2 558 -521 558 -521 0 net=5154
rlabel metal2 26 -523 26 -523 0 net=1448
rlabel metal2 324 -523 324 -523 0 net=3016
rlabel metal2 502 -523 502 -523 0 net=5413
rlabel metal2 30 -525 30 -525 0 net=491
rlabel metal2 460 -525 460 -525 0 net=3930
rlabel metal2 30 -527 30 -527 0 net=2921
rlabel metal2 611 -527 611 -527 0 net=5335
rlabel metal2 37 -529 37 -529 0 net=3645
rlabel metal2 310 -529 310 -529 0 net=2383
rlabel metal2 464 -529 464 -529 0 net=3735
rlabel metal2 618 -529 618 -529 0 net=4975
rlabel metal2 44 -531 44 -531 0 net=1224
rlabel metal2 296 -531 296 -531 0 net=2630
rlabel metal2 513 -531 513 -531 0 net=5095
rlabel metal2 44 -533 44 -533 0 net=4031
rlabel metal2 107 -533 107 -533 0 net=4104
rlabel metal2 576 -533 576 -533 0 net=4225
rlabel metal2 58 -535 58 -535 0 net=1514
rlabel metal2 282 -535 282 -535 0 net=1408
rlabel metal2 327 -535 327 -535 0 net=3340
rlabel metal2 562 -535 562 -535 0 net=4329
rlabel metal2 639 -535 639 -535 0 net=5089
rlabel metal2 51 -537 51 -537 0 net=5325
rlabel metal2 58 -539 58 -539 0 net=2181
rlabel metal2 387 -539 387 -539 0 net=530
rlabel metal2 65 -541 65 -541 0 net=2019
rlabel metal2 352 -541 352 -541 0 net=3463
rlabel metal2 401 -541 401 -541 0 net=2428
rlabel metal2 65 -543 65 -543 0 net=1681
rlabel metal2 306 -543 306 -543 0 net=4585
rlabel metal2 68 -545 68 -545 0 net=4573
rlabel metal2 72 -547 72 -547 0 net=2034
rlabel metal2 128 -547 128 -547 0 net=1434
rlabel metal2 355 -547 355 -547 0 net=5066
rlabel metal2 54 -549 54 -549 0 net=984
rlabel metal2 79 -549 79 -549 0 net=1132
rlabel metal2 240 -549 240 -549 0 net=2429
rlabel metal2 254 -549 254 -549 0 net=2504
rlabel metal2 425 -549 425 -549 0 net=3151
rlabel metal2 520 -549 520 -549 0 net=4461
rlabel metal2 79 -551 79 -551 0 net=3165
rlabel metal2 131 -551 131 -551 0 net=2665
rlabel metal2 404 -551 404 -551 0 net=5206
rlabel metal2 86 -553 86 -553 0 net=1235
rlabel metal2 194 -553 194 -553 0 net=1076
rlabel metal2 93 -555 93 -555 0 net=1271
rlabel metal2 93 -555 93 -555 0 net=1271
rlabel metal2 114 -555 114 -555 0 net=1013
rlabel metal2 233 -555 233 -555 0 net=1051
rlabel metal2 285 -555 285 -555 0 net=3828
rlabel metal2 541 -555 541 -555 0 net=4807
rlabel metal2 107 -557 107 -557 0 net=4061
rlabel metal2 541 -557 541 -557 0 net=4483
rlabel metal2 114 -559 114 -559 0 net=4124
rlabel metal2 135 -561 135 -561 0 net=2287
rlabel metal2 366 -561 366 -561 0 net=2103
rlabel metal2 366 -561 366 -561 0 net=2103
rlabel metal2 387 -561 387 -561 0 net=2461
rlabel metal2 478 -561 478 -561 0 net=3809
rlabel metal2 135 -563 135 -563 0 net=3446
rlabel metal2 569 -563 569 -563 0 net=4845
rlabel metal2 145 -565 145 -565 0 net=3914
rlabel metal2 625 -565 625 -565 0 net=5015
rlabel metal2 170 -567 170 -567 0 net=1751
rlabel metal2 201 -567 201 -567 0 net=2750
rlabel metal2 408 -567 408 -567 0 net=2490
rlabel metal2 478 -567 478 -567 0 net=3649
rlabel metal2 534 -567 534 -567 0 net=4893
rlabel metal2 177 -569 177 -569 0 net=2892
rlabel metal2 205 -569 205 -569 0 net=1717
rlabel metal2 289 -569 289 -569 0 net=3327
rlabel metal2 320 -569 320 -569 0 net=3797
rlabel metal2 506 -569 506 -569 0 net=4567
rlabel metal2 163 -571 163 -571 0 net=1423
rlabel metal2 184 -571 184 -571 0 net=3241
rlabel metal2 394 -571 394 -571 0 net=3018
rlabel metal2 411 -571 411 -571 0 net=5277
rlabel metal2 159 -573 159 -573 0 net=1721
rlabel metal2 205 -573 205 -573 0 net=1311
rlabel metal2 215 -573 215 -573 0 net=5045
rlabel metal2 215 -575 215 -575 0 net=2906
rlabel metal2 492 -575 492 -575 0 net=4855
rlabel metal2 219 -577 219 -577 0 net=1560
rlabel metal2 422 -577 422 -577 0 net=3025
rlabel metal2 457 -577 457 -577 0 net=5162
rlabel metal2 233 -579 233 -579 0 net=1059
rlabel metal2 548 -579 548 -579 0 net=4027
rlabel metal2 681 -579 681 -579 0 net=5437
rlabel metal2 121 -581 121 -581 0 net=4347
rlabel metal2 121 -583 121 -583 0 net=2775
rlabel metal2 173 -583 173 -583 0 net=5423
rlabel metal2 142 -585 142 -585 0 net=1537
rlabel metal2 240 -585 240 -585 0 net=1183
rlabel metal2 275 -585 275 -585 0 net=2051
rlabel metal2 243 -587 243 -587 0 net=3693
rlabel metal2 247 -589 247 -589 0 net=2549
rlabel metal2 149 -591 149 -591 0 net=1135
rlabel metal2 275 -591 275 -591 0 net=2774
rlabel metal2 149 -593 149 -593 0 net=2139
rlabel metal2 317 -593 317 -593 0 net=2282
rlabel metal2 443 -593 443 -593 0 net=5402
rlabel metal2 303 -595 303 -595 0 net=2453
rlabel metal2 23 -606 23 -606 0 net=3474
rlabel metal2 411 -606 411 -606 0 net=4586
rlabel metal2 611 -606 611 -606 0 net=5337
rlabel metal2 30 -608 30 -608 0 net=2923
rlabel metal2 709 -608 709 -608 0 net=5439
rlabel metal2 37 -610 37 -610 0 net=3646
rlabel metal2 93 -610 93 -610 0 net=1272
rlabel metal2 107 -610 107 -610 0 net=4330
rlabel metal2 625 -610 625 -610 0 net=5017
rlabel metal2 625 -610 625 -610 0 net=5017
rlabel metal2 632 -610 632 -610 0 net=5047
rlabel metal2 37 -612 37 -612 0 net=3243
rlabel metal2 187 -612 187 -612 0 net=430
rlabel metal2 219 -612 219 -612 0 net=5326
rlabel metal2 674 -612 674 -612 0 net=5415
rlabel metal2 44 -614 44 -614 0 net=4032
rlabel metal2 93 -614 93 -614 0 net=2455
rlabel metal2 415 -614 415 -614 0 net=4063
rlabel metal2 541 -614 541 -614 0 net=4485
rlabel metal2 44 -616 44 -616 0 net=2203
rlabel metal2 222 -616 222 -616 0 net=1175
rlabel metal2 51 -618 51 -618 0 net=3465
rlabel metal2 355 -618 355 -618 0 net=5343
rlabel metal2 58 -620 58 -620 0 net=2183
rlabel metal2 100 -620 100 -620 0 net=588
rlabel metal2 212 -620 212 -620 0 net=1095
rlabel metal2 226 -620 226 -620 0 net=1015
rlabel metal2 226 -620 226 -620 0 net=1015
rlabel metal2 233 -620 233 -620 0 net=1061
rlabel metal2 348 -620 348 -620 0 net=3739
rlabel metal2 569 -620 569 -620 0 net=4847
rlabel metal2 681 -620 681 -620 0 net=5425
rlabel metal2 23 -622 23 -622 0 net=428
rlabel metal2 75 -622 75 -622 0 net=1941
rlabel metal2 254 -622 254 -622 0 net=1053
rlabel metal2 254 -622 254 -622 0 net=1053
rlabel metal2 275 -622 275 -622 0 net=2462
rlabel metal2 418 -622 418 -622 0 net=4568
rlabel metal2 513 -622 513 -622 0 net=5097
rlabel metal2 79 -624 79 -624 0 net=3167
rlabel metal2 107 -624 107 -624 0 net=1539
rlabel metal2 170 -624 170 -624 0 net=1753
rlabel metal2 282 -624 282 -624 0 net=3665
rlabel metal2 555 -624 555 -624 0 net=5029
rlabel metal2 79 -626 79 -626 0 net=1313
rlabel metal2 303 -626 303 -626 0 net=2052
rlabel metal2 366 -626 366 -626 0 net=2105
rlabel metal2 366 -626 366 -626 0 net=2105
rlabel metal2 380 -626 380 -626 0 net=2667
rlabel metal2 422 -626 422 -626 0 net=3027
rlabel metal2 450 -626 450 -626 0 net=3799
rlabel metal2 583 -626 583 -626 0 net=5209
rlabel metal2 639 -626 639 -626 0 net=5091
rlabel metal2 114 -628 114 -628 0 net=2431
rlabel metal2 296 -628 296 -628 0 net=1683
rlabel metal2 425 -628 425 -628 0 net=5278
rlabel metal2 117 -630 117 -630 0 net=1136
rlabel metal2 261 -630 261 -630 0 net=4667
rlabel metal2 439 -630 439 -630 0 net=4894
rlabel metal2 590 -630 590 -630 0 net=4809
rlabel metal2 54 -632 54 -632 0 net=555
rlabel metal2 453 -632 453 -632 0 net=4691
rlabel metal2 121 -634 121 -634 0 net=2777
rlabel metal2 457 -634 457 -634 0 net=4395
rlabel metal2 618 -634 618 -634 0 net=4977
rlabel metal2 124 -636 124 -636 0 net=4887
rlabel metal2 128 -638 128 -638 0 net=2288
rlabel metal2 457 -638 457 -638 0 net=4462
rlabel metal2 135 -640 135 -640 0 net=3497
rlabel metal2 142 -642 142 -642 0 net=614
rlabel metal2 464 -642 464 -642 0 net=3737
rlabel metal2 163 -644 163 -644 0 net=1723
rlabel metal2 198 -644 198 -644 0 net=4091
rlabel metal2 149 -646 149 -646 0 net=2141
rlabel metal2 247 -646 247 -646 0 net=1719
rlabel metal2 296 -646 296 -646 0 net=2681
rlabel metal2 429 -646 429 -646 0 net=3152
rlabel metal2 471 -646 471 -646 0 net=3685
rlabel metal2 19 -648 19 -648 0 net=1571
rlabel metal2 303 -648 303 -648 0 net=1369
rlabel metal2 478 -648 478 -648 0 net=3651
rlabel metal2 86 -650 86 -650 0 net=1237
rlabel metal2 310 -650 310 -650 0 net=2385
rlabel metal2 478 -650 478 -650 0 net=4226
rlabel metal2 86 -652 86 -652 0 net=2577
rlabel metal2 317 -652 317 -652 0 net=5307
rlabel metal2 177 -654 177 -654 0 net=1425
rlabel metal2 320 -654 320 -654 0 net=4574
rlabel metal2 604 -654 604 -654 0 net=4857
rlabel metal2 177 -656 177 -656 0 net=1185
rlabel metal2 359 -656 359 -656 0 net=1781
rlabel metal2 485 -656 485 -656 0 net=3695
rlabel metal2 548 -656 548 -656 0 net=4349
rlabel metal2 159 -658 159 -658 0 net=1225
rlabel metal2 373 -658 373 -658 0 net=3971
rlabel metal2 194 -660 194 -660 0 net=969
rlabel metal2 324 -660 324 -660 0 net=2021
rlabel metal2 394 -660 394 -660 0 net=2551
rlabel metal2 467 -660 467 -660 0 net=2785
rlabel metal2 492 -660 492 -660 0 net=4028
rlabel metal2 201 -662 201 -662 0 net=3707
rlabel metal2 205 -664 205 -664 0 net=1147
rlabel metal2 460 -664 460 -664 0 net=4695
rlabel metal2 324 -666 324 -666 0 net=4429
rlabel metal2 499 -668 499 -668 0 net=3810
rlabel metal2 135 -670 135 -670 0 net=4127
rlabel metal2 289 -672 289 -672 0 net=3329
rlabel metal2 289 -674 289 -674 0 net=1273
rlabel metal2 30 -685 30 -685 0 net=587
rlabel metal2 467 -685 467 -685 0 net=5426
rlabel metal2 765 -685 765 -685 0 net=5441
rlabel metal2 37 -687 37 -687 0 net=3245
rlabel metal2 338 -687 338 -687 0 net=1063
rlabel metal2 338 -687 338 -687 0 net=1063
rlabel metal2 345 -687 345 -687 0 net=4692
rlabel metal2 730 -687 730 -687 0 net=5309
rlabel metal2 37 -689 37 -689 0 net=1541
rlabel metal2 114 -689 114 -689 0 net=2433
rlabel metal2 443 -689 443 -689 0 net=3029
rlabel metal2 485 -689 485 -689 0 net=2787
rlabel metal2 506 -689 506 -689 0 net=5273
rlabel metal2 772 -689 772 -689 0 net=5049
rlabel metal2 44 -691 44 -691 0 net=2204
rlabel metal2 362 -691 362 -691 0 net=2106
rlabel metal2 380 -691 380 -691 0 net=2669
rlabel metal2 495 -691 495 -691 0 net=5299
rlabel metal2 44 -693 44 -693 0 net=2457
rlabel metal2 107 -693 107 -693 0 net=1371
rlabel metal2 320 -693 320 -693 0 net=3738
rlabel metal2 586 -693 586 -693 0 net=5416
rlabel metal2 51 -695 51 -695 0 net=3466
rlabel metal2 450 -695 450 -695 0 net=4093
rlabel metal2 604 -695 604 -695 0 net=4351
rlabel metal2 744 -695 744 -695 0 net=5345
rlabel metal2 54 -697 54 -697 0 net=476
rlabel metal2 359 -697 359 -697 0 net=1783
rlabel metal2 383 -697 383 -697 0 net=2924
rlabel metal2 58 -699 58 -699 0 net=1317
rlabel metal2 65 -699 65 -699 0 net=2184
rlabel metal2 345 -699 345 -699 0 net=777
rlabel metal2 397 -699 397 -699 0 net=4978
rlabel metal2 65 -701 65 -701 0 net=3331
rlabel metal2 506 -701 506 -701 0 net=3499
rlabel metal2 520 -701 520 -701 0 net=3653
rlabel metal2 520 -701 520 -701 0 net=3653
rlabel metal2 527 -701 527 -701 0 net=3667
rlabel metal2 527 -701 527 -701 0 net=3667
rlabel metal2 541 -701 541 -701 0 net=3697
rlabel metal2 541 -701 541 -701 0 net=3697
rlabel metal2 548 -701 548 -701 0 net=3709
rlabel metal2 548 -701 548 -701 0 net=3709
rlabel metal2 555 -701 555 -701 0 net=3741
rlabel metal2 597 -701 597 -701 0 net=4129
rlabel metal2 632 -701 632 -701 0 net=5211
rlabel metal2 72 -703 72 -703 0 net=5113
rlabel metal2 72 -705 72 -705 0 net=4191
rlabel metal2 124 -705 124 -705 0 net=1274
rlabel metal2 296 -705 296 -705 0 net=2683
rlabel metal2 478 -705 478 -705 0 net=4319
rlabel metal2 646 -705 646 -705 0 net=4697
rlabel metal2 86 -707 86 -707 0 net=2578
rlabel metal2 212 -707 212 -707 0 net=1097
rlabel metal2 212 -707 212 -707 0 net=1097
rlabel metal2 222 -707 222 -707 0 net=1426
rlabel metal2 320 -707 320 -707 0 net=533
rlabel metal2 89 -709 89 -709 0 net=13
rlabel metal2 415 -709 415 -709 0 net=4065
rlabel metal2 625 -709 625 -709 0 net=5019
rlabel metal2 653 -709 653 -709 0 net=4811
rlabel metal2 128 -711 128 -711 0 net=4668
rlabel metal2 268 -711 268 -711 0 net=1238
rlabel metal2 289 -711 289 -711 0 net=492
rlabel metal2 562 -711 562 -711 0 net=3801
rlabel metal2 611 -711 611 -711 0 net=4397
rlabel metal2 79 -713 79 -713 0 net=1315
rlabel metal2 282 -713 282 -713 0 net=5189
rlabel metal2 79 -715 79 -715 0 net=1176
rlabel metal2 131 -717 131 -717 0 net=2778
rlabel metal2 397 -717 397 -717 0 net=4486
rlabel metal2 695 -717 695 -717 0 net=5031
rlabel metal2 16 -719 16 -719 0 net=4717
rlabel metal2 135 -721 135 -721 0 net=4019
rlabel metal2 618 -721 618 -721 0 net=4431
rlabel metal2 135 -723 135 -723 0 net=1149
rlabel metal2 233 -723 233 -723 0 net=1942
rlabel metal2 401 -723 401 -723 0 net=5338
rlabel metal2 114 -725 114 -725 0 net=2125
rlabel metal2 408 -725 408 -725 0 net=2387
rlabel metal2 429 -725 429 -725 0 net=2553
rlabel metal2 621 -725 621 -725 0 net=4737
rlabel metal2 121 -727 121 -727 0 net=1971
rlabel metal2 247 -727 247 -727 0 net=1720
rlabel metal2 348 -727 348 -727 0 net=480
rlabel metal2 499 -727 499 -727 0 net=3687
rlabel metal2 142 -729 142 -729 0 net=4888
rlabel metal2 124 -731 124 -731 0 net=1395
rlabel metal2 145 -731 145 -731 0 net=67
rlabel metal2 163 -731 163 -731 0 net=2143
rlabel metal2 429 -731 429 -731 0 net=4848
rlabel metal2 86 -733 86 -733 0 net=4251
rlabel metal2 156 -735 156 -735 0 net=5098
rlabel metal2 156 -737 156 -737 0 net=1493
rlabel metal2 247 -737 247 -737 0 net=1779
rlabel metal2 348 -737 348 -737 0 net=4385
rlabel metal2 163 -739 163 -739 0 net=1647
rlabel metal2 373 -739 373 -739 0 net=2023
rlabel metal2 394 -739 394 -739 0 net=4829
rlabel metal2 184 -741 184 -741 0 net=5105
rlabel metal2 170 -743 170 -743 0 net=1725
rlabel metal2 191 -743 191 -743 0 net=1755
rlabel metal2 254 -743 254 -743 0 net=1054
rlabel metal2 373 -743 373 -743 0 net=1797
rlabel metal2 149 -745 149 -745 0 net=1573
rlabel metal2 436 -745 436 -745 0 net=4579
rlabel metal2 149 -747 149 -747 0 net=5092
rlabel metal2 170 -749 170 -749 0 net=1017
rlabel metal2 254 -749 254 -749 0 net=1505
rlabel metal2 453 -749 453 -749 0 net=3561
rlabel metal2 576 -749 576 -749 0 net=3973
rlabel metal2 177 -751 177 -751 0 net=1187
rlabel metal2 201 -751 201 -751 0 net=4171
rlabel metal2 96 -753 96 -753 0 net=2107
rlabel metal2 201 -753 201 -753 0 net=1321
rlabel metal2 446 -753 446 -753 0 net=4005
rlabel metal2 226 -755 226 -755 0 net=1227
rlabel metal2 261 -755 261 -755 0 net=1685
rlabel metal2 481 -755 481 -755 0 net=4858
rlabel metal2 100 -757 100 -757 0 net=3169
rlabel metal2 439 -757 439 -757 0 net=4505
rlabel metal2 30 -759 30 -759 0 net=2505
rlabel metal2 240 -759 240 -759 0 net=2527
rlabel metal2 439 -759 439 -759 0 net=54
rlabel metal2 19 -770 19 -770 0 net=260
rlabel metal2 30 -770 30 -770 0 net=2065
rlabel metal2 408 -770 408 -770 0 net=2145
rlabel metal2 488 -770 488 -770 0 net=5271
rlabel metal2 849 -770 849 -770 0 net=5051
rlabel metal2 23 -772 23 -772 0 net=1687
rlabel metal2 159 -772 159 -772 0 net=1574
rlabel metal2 289 -772 289 -772 0 net=1322
rlabel metal2 310 -772 310 -772 0 net=3562
rlabel metal2 534 -772 534 -772 0 net=3974
rlabel metal2 751 -772 751 -772 0 net=5191
rlabel metal2 37 -774 37 -774 0 net=1542
rlabel metal2 177 -774 177 -774 0 net=2109
rlabel metal2 201 -774 201 -774 0 net=1686
rlabel metal2 268 -774 268 -774 0 net=1316
rlabel metal2 292 -774 292 -774 0 net=2670
rlabel metal2 460 -774 460 -774 0 net=3802
rlabel metal2 621 -774 621 -774 0 net=5300
rlabel metal2 779 -774 779 -774 0 net=5311
rlabel metal2 37 -776 37 -776 0 net=910
rlabel metal2 446 -776 446 -776 0 net=4812
rlabel metal2 758 -776 758 -776 0 net=5213
rlabel metal2 40 -778 40 -778 0 net=3081
rlabel metal2 296 -778 296 -778 0 net=3991
rlabel metal2 646 -778 646 -778 0 net=5021
rlabel metal2 793 -778 793 -778 0 net=5443
rlabel metal2 54 -780 54 -780 0 net=3332
rlabel metal2 86 -780 86 -780 0 net=124
rlabel metal2 222 -780 222 -780 0 net=4252
rlabel metal2 667 -780 667 -780 0 net=4507
rlabel metal2 765 -780 765 -780 0 net=5275
rlabel metal2 44 -782 44 -782 0 net=2459
rlabel metal2 226 -782 226 -782 0 net=1229
rlabel metal2 317 -782 317 -782 0 net=2159
rlabel metal2 352 -782 352 -782 0 net=4859
rlabel metal2 44 -784 44 -784 0 net=1495
rlabel metal2 166 -784 166 -784 0 net=4157
rlabel metal2 674 -784 674 -784 0 net=4581
rlabel metal2 58 -786 58 -786 0 net=1318
rlabel metal2 100 -786 100 -786 0 net=2507
rlabel metal2 320 -786 320 -786 0 net=2554
rlabel metal2 688 -786 688 -786 0 net=4719
rlabel metal2 65 -788 65 -788 0 net=2685
rlabel metal2 467 -788 467 -788 0 net=5106
rlabel metal2 72 -790 72 -790 0 net=4193
rlabel metal2 681 -790 681 -790 0 net=4699
rlabel metal2 79 -792 79 -792 0 net=3939
rlabel metal2 639 -792 639 -792 0 net=4353
rlabel metal2 695 -792 695 -792 0 net=4739
rlabel metal2 79 -794 79 -794 0 net=1373
rlabel metal2 114 -794 114 -794 0 net=1151
rlabel metal2 149 -794 149 -794 0 net=3115
rlabel metal2 327 -794 327 -794 0 net=889
rlabel metal2 411 -794 411 -794 0 net=4386
rlabel metal2 86 -796 86 -796 0 net=4627
rlabel metal2 89 -798 89 -798 0 net=298
rlabel metal2 89 -798 89 -798 0 net=298
rlabel metal2 93 -798 93 -798 0 net=1501
rlabel metal2 397 -798 397 -798 0 net=5346
rlabel metal2 117 -800 117 -800 0 net=4020
rlabel metal2 604 -800 604 -800 0 net=4131
rlabel metal2 653 -800 653 -800 0 net=4399
rlabel metal2 702 -800 702 -800 0 net=5033
rlabel metal2 121 -802 121 -802 0 net=2126
rlabel metal2 408 -802 408 -802 0 net=3943
rlabel metal2 611 -802 611 -802 0 net=4173
rlabel metal2 723 -802 723 -802 0 net=5115
rlabel metal2 72 -804 72 -804 0 net=1309
rlabel metal2 135 -804 135 -804 0 net=1189
rlabel metal2 198 -804 198 -804 0 net=96
rlabel metal2 436 -804 436 -804 0 net=2849
rlabel metal2 152 -806 152 -806 0 net=1817
rlabel metal2 338 -806 338 -806 0 net=1064
rlabel metal2 446 -806 446 -806 0 net=4997
rlabel metal2 58 -808 58 -808 0 net=2049
rlabel metal2 352 -808 352 -808 0 net=1799
rlabel metal2 429 -808 429 -808 0 net=4185
rlabel metal2 674 -808 674 -808 0 net=5363
rlabel metal2 156 -810 156 -810 0 net=1879
rlabel metal2 212 -810 212 -810 0 net=1099
rlabel metal2 212 -810 212 -810 0 net=1099
rlabel metal2 226 -810 226 -810 0 net=1123
rlabel metal2 401 -810 401 -810 0 net=2357
rlabel metal2 464 -810 464 -810 0 net=3773
rlabel metal2 625 -810 625 -810 0 net=4433
rlabel metal2 177 -812 177 -812 0 net=1727
rlabel metal2 233 -812 233 -812 0 net=1973
rlabel metal2 513 -812 513 -812 0 net=5463
rlabel metal2 170 -814 170 -814 0 net=1019
rlabel metal2 240 -814 240 -814 0 net=2529
rlabel metal2 247 -814 247 -814 0 net=1780
rlabel metal2 254 -814 254 -814 0 net=1506
rlabel metal2 520 -814 520 -814 0 net=3655
rlabel metal2 537 -814 537 -814 0 net=3933
rlabel metal2 142 -816 142 -816 0 net=1397
rlabel metal2 184 -816 184 -816 0 net=1757
rlabel metal2 240 -816 240 -816 0 net=2025
rlabel metal2 548 -816 548 -816 0 net=3711
rlabel metal2 569 -816 569 -816 0 net=4831
rlabel metal2 142 -818 142 -818 0 net=4066
rlabel metal2 163 -820 163 -820 0 net=1649
rlabel metal2 268 -820 268 -820 0 net=2879
rlabel metal2 499 -820 499 -820 0 net=3689
rlabel metal2 555 -820 555 -820 0 net=3743
rlabel metal2 576 -820 576 -820 0 net=4007
rlabel metal2 128 -822 128 -822 0 net=3753
rlabel metal2 128 -824 128 -824 0 net=2435
rlabel metal2 471 -824 471 -824 0 net=3031
rlabel metal2 541 -824 541 -824 0 net=3699
rlabel metal2 163 -826 163 -826 0 net=3246
rlabel metal2 331 -826 331 -826 0 net=3171
rlabel metal2 527 -826 527 -826 0 net=3669
rlabel metal2 107 -828 107 -828 0 net=1475
rlabel metal2 331 -828 331 -828 0 net=5077
rlabel metal2 243 -830 243 -830 0 net=1
rlabel metal2 471 -830 471 -830 0 net=2789
rlabel metal2 506 -830 506 -830 0 net=3501
rlabel metal2 299 -832 299 -832 0 net=2261
rlabel metal2 506 -832 506 -832 0 net=5193
rlabel metal2 306 -834 306 -834 0 net=4569
rlabel metal2 100 -836 100 -836 0 net=232
rlabel metal2 355 -836 355 -836 0 net=2388
rlabel metal2 359 -838 359 -838 0 net=3947
rlabel metal2 198 -840 198 -840 0 net=1673
rlabel metal2 366 -840 366 -840 0 net=1785
rlabel metal2 366 -842 366 -842 0 net=4321
rlabel metal2 383 -844 383 -844 0 net=2975
rlabel metal2 450 -846 450 -846 0 net=4095
rlabel metal2 450 -848 450 -848 0 net=4477
rlabel metal2 9 -859 9 -859 0 net=5265
rlabel metal2 674 -859 674 -859 0 net=5444
rlabel metal2 16 -861 16 -861 0 net=1881
rlabel metal2 201 -861 201 -861 0 net=720
rlabel metal2 282 -861 282 -861 0 net=1230
rlabel metal2 338 -861 338 -861 0 net=4322
rlabel metal2 404 -861 404 -861 0 net=3712
rlabel metal2 576 -861 576 -861 0 net=3755
rlabel metal2 576 -861 576 -861 0 net=3755
rlabel metal2 660 -861 660 -861 0 net=4187
rlabel metal2 831 -861 831 -861 0 net=5052
rlabel metal2 30 -863 30 -863 0 net=2066
rlabel metal2 240 -863 240 -863 0 net=2026
rlabel metal2 317 -863 317 -863 0 net=1819
rlabel metal2 411 -863 411 -863 0 net=2850
rlabel metal2 44 -865 44 -865 0 net=1496
rlabel metal2 163 -865 163 -865 0 net=5235
rlabel metal2 44 -867 44 -867 0 net=1801
rlabel metal2 359 -867 359 -867 0 net=3656
rlabel metal2 562 -867 562 -867 0 net=3949
rlabel metal2 653 -867 653 -867 0 net=4175
rlabel metal2 58 -869 58 -869 0 net=2050
rlabel metal2 261 -869 261 -869 0 net=2115
rlabel metal2 429 -869 429 -869 0 net=5192
rlabel metal2 72 -871 72 -871 0 net=4132
rlabel metal2 653 -871 653 -871 0 net=4629
rlabel metal2 744 -871 744 -871 0 net=5365
rlabel metal2 72 -873 72 -873 0 net=1477
rlabel metal2 121 -873 121 -873 0 net=1310
rlabel metal2 135 -873 135 -873 0 net=1190
rlabel metal2 268 -873 268 -873 0 net=2881
rlabel metal2 327 -873 327 -873 0 net=4720
rlabel metal2 23 -875 23 -875 0 net=1689
rlabel metal2 142 -875 142 -875 0 net=3116
rlabel metal2 317 -875 317 -875 0 net=2301
rlabel metal2 387 -875 387 -875 0 net=2531
rlabel metal2 443 -875 443 -875 0 net=5272
rlabel metal2 23 -877 23 -877 0 net=3173
rlabel metal2 590 -877 590 -877 0 net=4571
rlabel metal2 75 -879 75 -879 0 net=1974
rlabel metal2 387 -879 387 -879 0 net=2263
rlabel metal2 453 -879 453 -879 0 net=3502
rlabel metal2 597 -879 597 -879 0 net=3941
rlabel metal2 730 -879 730 -879 0 net=4833
rlabel metal2 79 -881 79 -881 0 net=1374
rlabel metal2 310 -881 310 -881 0 net=2509
rlabel metal2 457 -881 457 -881 0 net=3033
rlabel metal2 506 -881 506 -881 0 net=4508
rlabel metal2 744 -881 744 -881 0 net=4861
rlabel metal2 79 -883 79 -883 0 net=3449
rlabel metal2 611 -883 611 -883 0 net=4009
rlabel metal2 702 -883 702 -883 0 net=5035
rlabel metal2 765 -883 765 -883 0 net=5079
rlabel metal2 82 -885 82 -885 0 net=2146
rlabel metal2 506 -885 506 -885 0 net=4400
rlabel metal2 709 -885 709 -885 0 net=4701
rlabel metal2 800 -885 800 -885 0 net=5215
rlabel metal2 86 -887 86 -887 0 net=1152
rlabel metal2 142 -887 142 -887 0 net=2495
rlabel metal2 166 -887 166 -887 0 net=1728
rlabel metal2 184 -887 184 -887 0 net=1759
rlabel metal2 345 -887 345 -887 0 net=2161
rlabel metal2 439 -887 439 -887 0 net=3145
rlabel metal2 534 -887 534 -887 0 net=3529
rlabel metal2 30 -889 30 -889 0 net=1679
rlabel metal2 362 -889 362 -889 0 net=2593
rlabel metal2 460 -889 460 -889 0 net=5276
rlabel metal2 51 -891 51 -891 0 net=1839
rlabel metal2 177 -891 177 -891 0 net=1125
rlabel metal2 233 -891 233 -891 0 net=1021
rlabel metal2 464 -891 464 -891 0 net=3857
rlabel metal2 625 -891 625 -891 0 net=4435
rlabel metal2 737 -891 737 -891 0 net=4741
rlabel metal2 842 -891 842 -891 0 net=5465
rlabel metal2 40 -893 40 -893 0 net=4513
rlabel metal2 254 -893 254 -893 0 net=1651
rlabel metal2 467 -893 467 -893 0 net=3744
rlabel metal2 583 -893 583 -893 0 net=3775
rlabel metal2 751 -893 751 -893 0 net=4999
rlabel metal2 51 -895 51 -895 0 net=1786
rlabel metal2 478 -895 478 -895 0 net=4478
rlabel metal2 555 -895 555 -895 0 net=3701
rlabel metal2 681 -895 681 -895 0 net=4355
rlabel metal2 695 -895 695 -895 0 net=5023
rlabel metal2 86 -897 86 -897 0 net=3495
rlabel metal2 170 -897 170 -897 0 net=1399
rlabel metal2 254 -897 254 -897 0 net=1281
rlabel metal2 471 -897 471 -897 0 net=2790
rlabel metal2 541 -897 541 -897 0 net=3671
rlabel metal2 667 -897 667 -897 0 net=4195
rlabel metal2 716 -897 716 -897 0 net=3935
rlabel metal2 93 -899 93 -899 0 net=1502
rlabel metal2 156 -899 156 -899 0 net=1965
rlabel metal2 446 -899 446 -899 0 net=4183
rlabel metal2 716 -899 716 -899 0 net=5117
rlabel metal2 772 -899 772 -899 0 net=5195
rlabel metal2 93 -901 93 -901 0 net=2359
rlabel metal2 471 -901 471 -901 0 net=2977
rlabel metal2 646 -901 646 -901 0 net=4159
rlabel metal2 821 -901 821 -901 0 net=5313
rlabel metal2 54 -903 54 -903 0 net=3247
rlabel metal2 632 -903 632 -903 0 net=4097
rlabel metal2 835 -903 835 -903 0 net=5409
rlabel metal2 100 -905 100 -905 0 net=4582
rlabel metal2 65 -907 65 -907 0 net=2687
rlabel metal2 103 -907 103 -907 0 net=600
rlabel metal2 401 -907 401 -907 0 net=4467
rlabel metal2 618 -907 618 -907 0 net=3993
rlabel metal2 107 -909 107 -909 0 net=3147
rlabel metal2 191 -909 191 -909 0 net=1675
rlabel metal2 205 -909 205 -909 0 net=2111
rlabel metal2 485 -909 485 -909 0 net=3129
rlabel metal2 604 -909 604 -909 0 net=3945
rlabel metal2 58 -911 58 -911 0 net=2679
rlabel metal2 212 -911 212 -911 0 net=1101
rlabel metal2 261 -911 261 -911 0 net=1345
rlabel metal2 548 -911 548 -911 0 net=3691
rlabel metal2 128 -913 128 -913 0 net=2436
rlabel metal2 128 -915 128 -915 0 net=1261
rlabel metal2 215 -915 215 -915 0 net=3371
rlabel metal2 170 -917 170 -917 0 net=1363
rlabel metal2 219 -917 219 -917 0 net=2460
rlabel metal2 380 -917 380 -917 0 net=2171
rlabel metal2 219 -919 219 -919 0 net=2821
rlabel metal2 275 -921 275 -921 0 net=3083
rlabel metal2 303 -923 303 -923 0 net=5249
rlabel metal2 19 -925 19 -925 0 net=3839
rlabel metal2 331 -925 331 -925 0 net=2397
rlabel metal2 2 -936 2 -936 0 net=4515
rlabel metal2 247 -936 247 -936 0 net=1346
rlabel metal2 275 -936 275 -936 0 net=2113
rlabel metal2 390 -936 390 -936 0 net=4160
rlabel metal2 779 -936 779 -936 0 net=3937
rlabel metal2 9 -938 9 -938 0 net=5266
rlabel metal2 100 -938 100 -938 0 net=2688
rlabel metal2 348 -938 348 -938 0 net=4572
rlabel metal2 814 -938 814 -938 0 net=5367
rlabel metal2 9 -940 9 -940 0 net=1263
rlabel metal2 149 -940 149 -940 0 net=1365
rlabel metal2 173 -940 173 -940 0 net=2264
rlabel metal2 394 -940 394 -940 0 net=2594
rlabel metal2 450 -940 450 -940 0 net=5417
rlabel metal2 16 -942 16 -942 0 net=1882
rlabel metal2 352 -942 352 -942 0 net=3146
rlabel metal2 509 -942 509 -942 0 net=4742
rlabel metal2 786 -942 786 -942 0 net=5143
rlabel metal2 842 -942 842 -942 0 net=5467
rlabel metal2 842 -942 842 -942 0 net=5467
rlabel metal2 30 -944 30 -944 0 net=1680
rlabel metal2 331 -944 331 -944 0 net=2399
rlabel metal2 397 -944 397 -944 0 net=4188
rlabel metal2 716 -944 716 -944 0 net=5119
rlabel metal2 814 -944 814 -944 0 net=5411
rlabel metal2 37 -946 37 -946 0 net=2571
rlabel metal2 128 -946 128 -946 0 net=730
rlabel metal2 247 -946 247 -946 0 net=1205
rlabel metal2 331 -946 331 -946 0 net=3776
rlabel metal2 737 -946 737 -946 0 net=4863
rlabel metal2 40 -948 40 -948 0 net=1478
rlabel metal2 79 -948 79 -948 0 net=2173
rlabel metal2 401 -948 401 -948 0 net=4184
rlabel metal2 744 -948 744 -948 0 net=5001
rlabel metal2 44 -950 44 -950 0 net=1802
rlabel metal2 404 -950 404 -950 0 net=1820
rlabel metal2 429 -950 429 -950 0 net=2532
rlabel metal2 513 -950 513 -950 0 net=4176
rlabel metal2 751 -950 751 -950 0 net=5251
rlabel metal2 51 -952 51 -952 0 net=2361
rlabel metal2 117 -952 117 -952 0 net=3756
rlabel metal2 590 -952 590 -952 0 net=5314
rlabel metal2 58 -954 58 -954 0 net=2680
rlabel metal2 408 -954 408 -954 0 net=3692
rlabel metal2 646 -954 646 -954 0 net=4099
rlabel metal2 793 -954 793 -954 0 net=5237
rlabel metal2 58 -956 58 -956 0 net=2925
rlabel metal2 121 -956 121 -956 0 net=10
rlabel metal2 201 -956 201 -956 0 net=2621
rlabel metal2 303 -956 303 -956 0 net=3841
rlabel metal2 646 -956 646 -956 0 net=4357
rlabel metal2 44 -958 44 -958 0 net=2441
rlabel metal2 152 -958 152 -958 0 net=5267
rlabel metal2 61 -960 61 -960 0 net=880
rlabel metal2 429 -960 429 -960 0 net=5261
rlabel metal2 65 -962 65 -962 0 net=3496
rlabel metal2 163 -962 163 -962 0 net=3131
rlabel metal2 516 -962 516 -962 0 net=5155
rlabel metal2 65 -964 65 -964 0 net=2163
rlabel metal2 436 -964 436 -964 0 net=3994
rlabel metal2 653 -964 653 -964 0 net=4631
rlabel metal2 72 -966 72 -966 0 net=1967
rlabel metal2 177 -966 177 -966 0 net=1127
rlabel metal2 373 -966 373 -966 0 net=3335
rlabel metal2 443 -966 443 -966 0 net=5255
rlabel metal2 86 -968 86 -968 0 net=2303
rlabel metal2 443 -968 443 -968 0 net=3035
rlabel metal2 464 -968 464 -968 0 net=2979
rlabel metal2 474 -968 474 -968 0 net=4905
rlabel metal2 135 -970 135 -970 0 net=1691
rlabel metal2 177 -970 177 -970 0 net=1401
rlabel metal2 254 -970 254 -970 0 net=1283
rlabel metal2 317 -970 317 -970 0 net=2713
rlabel metal2 446 -970 446 -970 0 net=4731
rlabel metal2 135 -972 135 -972 0 net=1193
rlabel metal2 205 -972 205 -972 0 net=1643
rlabel metal2 170 -974 170 -974 0 net=3423
rlabel metal2 254 -974 254 -974 0 net=3967
rlabel metal2 457 -974 457 -974 0 net=3249
rlabel metal2 520 -974 520 -974 0 net=3373
rlabel metal2 520 -974 520 -974 0 net=3373
rlabel metal2 527 -974 527 -974 0 net=3451
rlabel metal2 527 -974 527 -974 0 net=3451
rlabel metal2 534 -974 534 -974 0 net=3531
rlabel metal2 534 -974 534 -974 0 net=3531
rlabel metal2 541 -974 541 -974 0 net=3946
rlabel metal2 653 -974 653 -974 0 net=4197
rlabel metal2 688 -974 688 -974 0 net=5025
rlabel metal2 191 -976 191 -976 0 net=1677
rlabel metal2 261 -976 261 -976 0 net=1023
rlabel metal2 278 -976 278 -976 0 net=2510
rlabel metal2 450 -976 450 -976 0 net=3085
rlabel metal2 481 -976 481 -976 0 net=3581
rlabel metal2 548 -976 548 -976 0 net=5216
rlabel metal2 208 -978 208 -978 0 net=3942
rlabel metal2 695 -978 695 -978 0 net=4835
rlabel metal2 772 -978 772 -978 0 net=5197
rlabel metal2 212 -980 212 -980 0 net=1739
rlabel metal2 478 -980 478 -980 0 net=4303
rlabel metal2 765 -980 765 -980 0 net=5081
rlabel metal2 215 -982 215 -982 0 net=1760
rlabel metal2 338 -982 338 -982 0 net=3605
rlabel metal2 562 -982 562 -982 0 net=3951
rlabel metal2 639 -982 639 -982 0 net=4703
rlabel metal2 758 -982 758 -982 0 net=5037
rlabel metal2 184 -984 184 -984 0 net=4751
rlabel metal2 758 -984 758 -984 0 net=5297
rlabel metal2 142 -986 142 -986 0 net=2497
rlabel metal2 219 -986 219 -986 0 net=1102
rlabel metal2 268 -986 268 -986 0 net=2147
rlabel metal2 376 -986 376 -986 0 net=4527
rlabel metal2 114 -988 114 -988 0 net=1841
rlabel metal2 240 -988 240 -988 0 net=2823
rlabel metal2 485 -988 485 -988 0 net=3703
rlabel metal2 576 -988 576 -988 0 net=3859
rlabel metal2 114 -990 114 -990 0 net=4403
rlabel metal2 289 -992 289 -992 0 net=1653
rlabel metal2 289 -994 289 -994 0 net=2883
rlabel metal2 345 -994 345 -994 0 net=2117
rlabel metal2 404 -994 404 -994 0 net=2869
rlabel metal2 555 -994 555 -994 0 net=3673
rlabel metal2 583 -994 583 -994 0 net=4469
rlabel metal2 23 -996 23 -996 0 net=3174
rlabel metal2 555 -996 555 -996 0 net=4436
rlabel metal2 23 -998 23 -998 0 net=3149
rlabel metal2 299 -998 299 -998 0 net=3811
rlabel metal2 558 -998 558 -998 0 net=3291
rlabel metal2 597 -998 597 -998 0 net=3713
rlabel metal2 107 -1000 107 -1000 0 net=2229
rlabel metal2 324 -1000 324 -1000 0 net=1869
rlabel metal2 611 -1000 611 -1000 0 net=4011
rlabel metal2 425 -1002 425 -1002 0 net=4067
rlabel metal2 506 -1004 506 -1004 0 net=3887
rlabel metal2 2 -1015 2 -1015 0 net=4516
rlabel metal2 422 -1015 422 -1015 0 net=3583
rlabel metal2 551 -1015 551 -1015 0 net=4906
rlabel metal2 786 -1015 786 -1015 0 net=5145
rlabel metal2 863 -1015 863 -1015 0 net=5419
rlabel metal2 9 -1017 9 -1017 0 net=1264
rlabel metal2 212 -1017 212 -1017 0 net=1741
rlabel metal2 341 -1017 341 -1017 0 net=3812
rlabel metal2 502 -1017 502 -1017 0 net=5468
rlabel metal2 849 -1017 849 -1017 0 net=5369
rlabel metal2 16 -1019 16 -1019 0 net=1645
rlabel metal2 212 -1019 212 -1019 0 net=1167
rlabel metal2 404 -1019 404 -1019 0 net=3704
rlabel metal2 492 -1019 492 -1019 0 net=5451
rlabel metal2 898 -1019 898 -1019 0 net=3938
rlabel metal2 19 -1021 19 -1021 0 net=4821
rlabel metal2 793 -1021 793 -1021 0 net=5157
rlabel metal2 793 -1021 793 -1021 0 net=5157
rlabel metal2 800 -1021 800 -1021 0 net=5199
rlabel metal2 23 -1023 23 -1023 0 net=3150
rlabel metal2 30 -1023 30 -1023 0 net=2573
rlabel metal2 205 -1023 205 -1023 0 net=1025
rlabel metal2 303 -1023 303 -1023 0 net=1128
rlabel metal2 478 -1023 478 -1023 0 net=4704
rlabel metal2 642 -1023 642 -1023 0 net=5123
rlabel metal2 23 -1025 23 -1025 0 net=1693
rlabel metal2 166 -1025 166 -1025 0 net=1678
rlabel metal2 261 -1025 261 -1025 0 net=1469
rlabel metal2 590 -1025 590 -1025 0 net=3843
rlabel metal2 33 -1027 33 -1027 0 net=4752
rlabel metal2 772 -1027 772 -1027 0 net=5083
rlabel metal2 807 -1027 807 -1027 0 net=5239
rlabel metal2 37 -1029 37 -1029 0 net=2572
rlabel metal2 219 -1029 219 -1029 0 net=2622
rlabel metal2 303 -1029 303 -1029 0 net=1871
rlabel metal2 331 -1029 331 -1029 0 net=4528
rlabel metal2 772 -1029 772 -1029 0 net=4913
rlabel metal2 37 -1031 37 -1031 0 net=2305
rlabel metal2 93 -1031 93 -1031 0 net=2927
rlabel metal2 439 -1031 439 -1031 0 net=2639
rlabel metal2 506 -1031 506 -1031 0 net=4068
rlabel metal2 618 -1031 618 -1031 0 net=3953
rlabel metal2 618 -1031 618 -1031 0 net=3953
rlabel metal2 660 -1031 660 -1031 0 net=4305
rlabel metal2 779 -1031 779 -1031 0 net=5121
rlabel metal2 54 -1033 54 -1033 0 net=1663
rlabel metal2 107 -1033 107 -1033 0 net=2231
rlabel metal2 415 -1033 415 -1033 0 net=2871
rlabel metal2 513 -1033 513 -1033 0 net=5252
rlabel metal2 821 -1033 821 -1033 0 net=5257
rlabel metal2 58 -1035 58 -1035 0 net=1853
rlabel metal2 163 -1035 163 -1035 0 net=3133
rlabel metal2 516 -1035 516 -1035 0 net=3714
rlabel metal2 604 -1035 604 -1035 0 net=3889
rlabel metal2 681 -1035 681 -1035 0 net=4471
rlabel metal2 828 -1035 828 -1035 0 net=5263
rlabel metal2 65 -1037 65 -1037 0 net=2165
rlabel metal2 432 -1037 432 -1037 0 net=3036
rlabel metal2 446 -1037 446 -1037 0 net=4951
rlabel metal2 835 -1037 835 -1037 0 net=5269
rlabel metal2 65 -1039 65 -1039 0 net=3968
rlabel metal2 278 -1039 278 -1039 0 net=1457
rlabel metal2 289 -1039 289 -1039 0 net=2885
rlabel metal2 527 -1039 527 -1039 0 net=3453
rlabel metal2 604 -1039 604 -1039 0 net=5002
rlabel metal2 72 -1041 72 -1041 0 net=1968
rlabel metal2 121 -1041 121 -1041 0 net=1843
rlabel metal2 163 -1041 163 -1041 0 net=5412
rlabel metal2 72 -1043 72 -1043 0 net=1367
rlabel metal2 152 -1043 152 -1043 0 net=4491
rlabel metal2 79 -1045 79 -1045 0 net=2175
rlabel metal2 317 -1045 317 -1045 0 net=2715
rlabel metal2 453 -1045 453 -1045 0 net=612
rlabel metal2 576 -1045 576 -1045 0 net=3861
rlabel metal2 674 -1045 674 -1045 0 net=4405
rlabel metal2 79 -1047 79 -1047 0 net=2114
rlabel metal2 296 -1047 296 -1047 0 net=1285
rlabel metal2 352 -1047 352 -1047 0 net=2149
rlabel metal2 499 -1047 499 -1047 0 net=5067
rlabel metal2 103 -1049 103 -1049 0 net=1893
rlabel metal2 128 -1049 128 -1049 0 net=4100
rlabel metal2 688 -1049 688 -1049 0 net=5027
rlabel metal2 107 -1051 107 -1051 0 net=1137
rlabel metal2 128 -1051 128 -1051 0 net=2131
rlabel metal2 352 -1051 352 -1051 0 net=3393
rlabel metal2 614 -1051 614 -1051 0 net=1
rlabel metal2 695 -1051 695 -1051 0 net=4837
rlabel metal2 135 -1053 135 -1053 0 net=1195
rlabel metal2 170 -1053 170 -1053 0 net=3287
rlabel metal2 275 -1053 275 -1053 0 net=3086
rlabel metal2 464 -1053 464 -1053 0 net=2981
rlabel metal2 520 -1053 520 -1053 0 net=3375
rlabel metal2 702 -1053 702 -1053 0 net=4633
rlabel metal2 702 -1053 702 -1053 0 net=4633
rlabel metal2 716 -1053 716 -1053 0 net=4733
rlabel metal2 177 -1055 177 -1055 0 net=1403
rlabel metal2 243 -1055 243 -1055 0 net=1463
rlabel metal2 317 -1055 317 -1055 0 net=2511
rlabel metal2 527 -1055 527 -1055 0 net=3921
rlabel metal2 737 -1055 737 -1055 0 net=4865
rlabel metal2 100 -1057 100 -1057 0 net=1037
rlabel metal2 184 -1057 184 -1057 0 net=2499
rlabel metal2 268 -1057 268 -1057 0 net=1975
rlabel metal2 359 -1057 359 -1057 0 net=2401
rlabel metal2 380 -1057 380 -1057 0 net=3336
rlabel metal2 429 -1057 429 -1057 0 net=3023
rlabel metal2 534 -1057 534 -1057 0 net=3533
rlabel metal2 191 -1059 191 -1059 0 net=1515
rlabel metal2 226 -1059 226 -1059 0 net=3425
rlabel metal2 565 -1059 565 -1059 0 net=5279
rlabel metal2 44 -1061 44 -1061 0 net=2442
rlabel metal2 226 -1061 226 -1061 0 net=2825
rlabel metal2 247 -1061 247 -1061 0 net=1207
rlabel metal2 345 -1061 345 -1061 0 net=2119
rlabel metal2 387 -1061 387 -1061 0 net=1654
rlabel metal2 646 -1061 646 -1061 0 net=4359
rlabel metal2 44 -1063 44 -1063 0 net=2363
rlabel metal2 201 -1063 201 -1063 0 net=3213
rlabel metal2 345 -1063 345 -1063 0 net=5298
rlabel metal2 359 -1065 359 -1065 0 net=1913
rlabel metal2 548 -1065 548 -1065 0 net=3607
rlabel metal2 653 -1065 653 -1065 0 net=4199
rlabel metal2 758 -1065 758 -1065 0 net=5039
rlabel metal2 184 -1067 184 -1067 0 net=3153
rlabel metal2 562 -1067 562 -1067 0 net=3675
rlabel metal2 366 -1069 366 -1069 0 net=3535
rlabel metal2 625 -1069 625 -1069 0 net=4013
rlabel metal2 366 -1071 366 -1071 0 net=1931
rlabel metal2 534 -1071 534 -1071 0 net=4537
rlabel metal2 376 -1073 376 -1073 0 net=3745
rlabel metal2 390 -1075 390 -1075 0 net=2581
rlabel metal2 562 -1075 562 -1075 0 net=4423
rlabel metal2 429 -1077 429 -1077 0 net=3251
rlabel metal2 569 -1077 569 -1077 0 net=3293
rlabel metal2 607 -1077 607 -1077 0 net=4113
rlabel metal2 194 -1079 194 -1079 0 net=3435
rlabel metal2 450 -1081 450 -1081 0 net=3503
rlabel metal2 9 -1092 9 -1092 0 net=4822
rlabel metal2 807 -1092 807 -1092 0 net=4953
rlabel metal2 807 -1092 807 -1092 0 net=4953
rlabel metal2 884 -1092 884 -1092 0 net=5453
rlabel metal2 982 -1092 982 -1092 0 net=2185
rlabel metal2 9 -1094 9 -1094 0 net=3289
rlabel metal2 198 -1094 198 -1094 0 net=2826
rlabel metal2 240 -1094 240 -1094 0 net=1459
rlabel metal2 317 -1094 317 -1094 0 net=2513
rlabel metal2 446 -1094 446 -1094 0 net=3844
rlabel metal2 898 -1094 898 -1094 0 net=5264
rlabel metal2 16 -1096 16 -1096 0 net=1646
rlabel metal2 642 -1096 642 -1096 0 net=5122
rlabel metal2 856 -1096 856 -1096 0 net=5147
rlabel metal2 912 -1096 912 -1096 0 net=5371
rlabel metal2 16 -1098 16 -1098 0 net=2575
rlabel metal2 44 -1098 44 -1098 0 net=2364
rlabel metal2 103 -1098 103 -1098 0 net=4200
rlabel metal2 828 -1098 828 -1098 0 net=5069
rlabel metal2 940 -1098 940 -1098 0 net=5259
rlabel metal2 940 -1098 940 -1098 0 net=5259
rlabel metal2 30 -1100 30 -1100 0 net=2307
rlabel metal2 44 -1100 44 -1100 0 net=1027
rlabel metal2 226 -1100 226 -1100 0 net=2177
rlabel metal2 345 -1100 345 -1100 0 net=1933
rlabel metal2 387 -1100 387 -1100 0 net=2233
rlabel metal2 436 -1100 436 -1100 0 net=2929
rlabel metal2 450 -1100 450 -1100 0 net=629
rlabel metal2 667 -1100 667 -1100 0 net=5281
rlabel metal2 37 -1102 37 -1102 0 net=1977
rlabel metal2 275 -1102 275 -1102 0 net=3787
rlabel metal2 348 -1102 348 -1102 0 net=2166
rlabel metal2 436 -1102 436 -1102 0 net=2241
rlabel metal2 506 -1102 506 -1102 0 net=2887
rlabel metal2 544 -1102 544 -1102 0 net=5028
rlabel metal2 842 -1102 842 -1102 0 net=5125
rlabel metal2 51 -1104 51 -1104 0 net=1665
rlabel metal2 93 -1104 93 -1104 0 net=5229
rlabel metal2 58 -1106 58 -1106 0 net=1855
rlabel metal2 72 -1106 72 -1106 0 net=1368
rlabel metal2 156 -1106 156 -1106 0 net=1039
rlabel metal2 198 -1106 198 -1106 0 net=2913
rlabel metal2 558 -1106 558 -1106 0 net=4838
rlabel metal2 58 -1108 58 -1108 0 net=2501
rlabel metal2 268 -1108 268 -1108 0 net=1209
rlabel metal2 303 -1108 303 -1108 0 net=1873
rlabel metal2 355 -1108 355 -1108 0 net=3534
rlabel metal2 702 -1108 702 -1108 0 net=4635
rlabel metal2 863 -1108 863 -1108 0 net=4655
rlabel metal2 72 -1110 72 -1110 0 net=712
rlabel metal2 205 -1110 205 -1110 0 net=2077
rlabel metal2 366 -1110 366 -1110 0 net=3609
rlabel metal2 684 -1110 684 -1110 0 net=5200
rlabel metal2 82 -1112 82 -1112 0 net=247
rlabel metal2 247 -1112 247 -1112 0 net=1465
rlabel metal2 303 -1112 303 -1112 0 net=1287
rlabel metal2 355 -1112 355 -1112 0 net=2415
rlabel metal2 520 -1112 520 -1112 0 net=3024
rlabel metal2 607 -1112 607 -1112 0 net=3517
rlabel metal2 702 -1112 702 -1112 0 net=3717
rlabel metal2 751 -1112 751 -1112 0 net=4539
rlabel metal2 849 -1112 849 -1112 0 net=4559
rlabel metal2 86 -1114 86 -1114 0 net=1139
rlabel metal2 128 -1114 128 -1114 0 net=2133
rlabel metal2 331 -1114 331 -1114 0 net=3215
rlabel metal2 758 -1114 758 -1114 0 net=5041
rlabel metal2 103 -1116 103 -1116 0 net=1577
rlabel metal2 278 -1116 278 -1116 0 net=3957
rlabel metal2 800 -1116 800 -1116 0 net=5085
rlabel metal2 107 -1118 107 -1118 0 net=1895
rlabel metal2 128 -1118 128 -1118 0 net=1197
rlabel metal2 152 -1118 152 -1118 0 net=349
rlabel metal2 527 -1118 527 -1118 0 net=4360
rlabel metal2 114 -1120 114 -1120 0 net=2121
rlabel metal2 390 -1120 390 -1120 0 net=5420
rlabel metal2 135 -1122 135 -1122 0 net=4263
rlabel metal2 870 -1122 870 -1122 0 net=5241
rlabel metal2 135 -1124 135 -1124 0 net=2753
rlabel metal2 530 -1124 530 -1124 0 net=5270
rlabel metal2 138 -1126 138 -1126 0 net=1404
rlabel metal2 250 -1126 250 -1126 0 net=3661
rlabel metal2 772 -1126 772 -1126 0 net=4915
rlabel metal2 23 -1128 23 -1128 0 net=1695
rlabel metal2 282 -1128 282 -1128 0 net=2759
rlabel metal2 562 -1128 562 -1128 0 net=4492
rlabel metal2 93 -1130 93 -1130 0 net=4105
rlabel metal2 793 -1130 793 -1130 0 net=5159
rlabel metal2 142 -1132 142 -1132 0 net=3253
rlabel metal2 453 -1132 453 -1132 0 net=3504
rlabel metal2 709 -1132 709 -1132 0 net=4425
rlabel metal2 163 -1134 163 -1134 0 net=1471
rlabel metal2 289 -1134 289 -1134 0 net=1915
rlabel metal2 380 -1134 380 -1134 0 net=2151
rlabel metal2 422 -1134 422 -1134 0 net=3585
rlabel metal2 166 -1136 166 -1136 0 net=4943
rlabel metal2 177 -1138 177 -1138 0 net=1517
rlabel metal2 261 -1138 261 -1138 0 net=2873
rlabel metal2 562 -1138 562 -1138 0 net=2997
rlabel metal2 184 -1140 184 -1140 0 net=3155
rlabel metal2 464 -1140 464 -1140 0 net=4866
rlabel metal2 170 -1142 170 -1142 0 net=1043
rlabel metal2 191 -1142 191 -1142 0 net=1169
rlabel metal2 324 -1142 324 -1142 0 net=1543
rlabel metal2 485 -1142 485 -1142 0 net=2611
rlabel metal2 569 -1142 569 -1142 0 net=4331
rlabel metal2 331 -1144 331 -1144 0 net=3455
rlabel metal2 618 -1144 618 -1144 0 net=3955
rlabel metal2 338 -1146 338 -1146 0 net=1742
rlabel metal2 513 -1146 513 -1146 0 net=3135
rlabel metal2 572 -1146 572 -1146 0 net=4014
rlabel metal2 222 -1148 222 -1148 0 net=3969
rlabel metal2 222 -1150 222 -1150 0 net=3381
rlabel metal2 401 -1150 401 -1150 0 net=2717
rlabel metal2 576 -1150 576 -1150 0 net=3377
rlabel metal2 646 -1150 646 -1150 0 net=3677
rlabel metal2 730 -1150 730 -1150 0 net=4473
rlabel metal2 338 -1152 338 -1152 0 net=2403
rlabel metal2 583 -1152 583 -1152 0 net=3395
rlabel metal2 646 -1152 646 -1152 0 net=3923
rlabel metal2 359 -1154 359 -1154 0 net=4734
rlabel metal2 373 -1156 373 -1156 0 net=1389
rlabel metal2 548 -1156 548 -1156 0 net=2855
rlabel metal2 744 -1156 744 -1156 0 net=4407
rlabel metal2 79 -1158 79 -1158 0 net=4437
rlabel metal2 79 -1160 79 -1160 0 net=1845
rlabel metal2 425 -1160 425 -1160 0 net=3553
rlabel metal2 618 -1160 618 -1160 0 net=4306
rlabel metal2 625 -1162 625 -1162 0 net=4115
rlabel metal2 611 -1164 611 -1164 0 net=3537
rlabel metal2 653 -1164 653 -1164 0 net=3747
rlabel metal2 597 -1166 597 -1166 0 net=3295
rlabel metal2 656 -1166 656 -1166 0 net=5357
rlabel metal2 499 -1168 499 -1168 0 net=2983
rlabel metal2 660 -1168 660 -1168 0 net=3863
rlabel metal2 478 -1170 478 -1170 0 net=2641
rlabel metal2 541 -1170 541 -1170 0 net=3427
rlabel metal2 674 -1170 674 -1170 0 net=3891
rlabel metal2 401 -1172 401 -1172 0 net=1449
rlabel metal2 541 -1172 541 -1172 0 net=3097
rlabel metal2 457 -1174 457 -1174 0 net=3437
rlabel metal2 457 -1176 457 -1176 0 net=2583
rlabel metal2 212 -1178 212 -1178 0 net=2601
rlabel metal2 5 -1189 5 -1189 0 net=263
rlabel metal2 222 -1189 222 -1189 0 net=3438
rlabel metal2 719 -1189 719 -1189 0 net=5086
rlabel metal2 940 -1189 940 -1189 0 net=5260
rlabel metal2 975 -1189 975 -1189 0 net=5455
rlabel metal2 985 -1189 985 -1189 0 net=4615
rlabel metal2 9 -1191 9 -1191 0 net=3290
rlabel metal2 215 -1191 215 -1191 0 net=3748
rlabel metal2 737 -1191 737 -1191 0 net=3893
rlabel metal2 751 -1191 751 -1191 0 net=3959
rlabel metal2 989 -1191 989 -1191 0 net=2187
rlabel metal2 16 -1193 16 -1193 0 net=2576
rlabel metal2 247 -1193 247 -1193 0 net=1467
rlabel metal2 247 -1193 247 -1193 0 net=1467
rlabel metal2 254 -1193 254 -1193 0 net=1578
rlabel metal2 341 -1193 341 -1193 0 net=408
rlabel metal2 625 -1193 625 -1193 0 net=3539
rlabel metal2 723 -1193 723 -1193 0 net=4439
rlabel metal2 800 -1193 800 -1193 0 net=4333
rlabel metal2 968 -1193 968 -1193 0 net=2481
rlabel metal2 16 -1195 16 -1195 0 net=1519
rlabel metal2 201 -1195 201 -1195 0 net=3970
rlabel metal2 800 -1195 800 -1195 0 net=5071
rlabel metal2 912 -1195 912 -1195 0 net=5231
rlabel metal2 26 -1197 26 -1197 0 net=466
rlabel metal2 26 -1197 26 -1197 0 net=466
rlabel metal2 44 -1197 44 -1197 0 net=1028
rlabel metal2 352 -1197 352 -1197 0 net=2613
rlabel metal2 506 -1197 506 -1197 0 net=5148
rlabel metal2 58 -1199 58 -1199 0 net=2502
rlabel metal2 254 -1199 254 -1199 0 net=2907
rlabel metal2 373 -1199 373 -1199 0 net=1391
rlabel metal2 429 -1199 429 -1199 0 net=3157
rlabel metal2 814 -1199 814 -1199 0 net=4427
rlabel metal2 58 -1201 58 -1201 0 net=2205
rlabel metal2 464 -1201 464 -1201 0 net=4116
rlabel metal2 814 -1201 814 -1201 0 net=5359
rlabel metal2 72 -1203 72 -1203 0 net=2437
rlabel metal2 268 -1203 268 -1203 0 net=1211
rlabel metal2 355 -1203 355 -1203 0 net=3610
rlabel metal2 411 -1203 411 -1203 0 net=3586
rlabel metal2 737 -1203 737 -1203 0 net=4637
rlabel metal2 65 -1205 65 -1205 0 net=1857
rlabel metal2 411 -1205 411 -1205 0 net=3401
rlabel metal2 842 -1205 842 -1205 0 net=4541
rlabel metal2 65 -1207 65 -1207 0 net=2643
rlabel metal2 534 -1207 534 -1207 0 net=2889
rlabel metal2 786 -1207 786 -1207 0 net=4265
rlabel metal2 849 -1207 849 -1207 0 net=4561
rlabel metal2 86 -1209 86 -1209 0 net=1140
rlabel metal2 135 -1209 135 -1209 0 net=2178
rlabel metal2 268 -1209 268 -1209 0 net=1289
rlabel metal2 310 -1209 310 -1209 0 net=1875
rlabel metal2 429 -1209 429 -1209 0 net=2999
rlabel metal2 579 -1209 579 -1209 0 net=4101
rlabel metal2 79 -1211 79 -1211 0 net=1847
rlabel metal2 142 -1211 142 -1211 0 net=3254
rlabel metal2 359 -1211 359 -1211 0 net=4954
rlabel metal2 30 -1213 30 -1213 0 net=2309
rlabel metal2 149 -1213 149 -1213 0 net=3456
rlabel metal2 446 -1213 446 -1213 0 net=3678
rlabel metal2 772 -1213 772 -1213 0 net=4107
rlabel metal2 30 -1215 30 -1215 0 net=1265
rlabel metal2 450 -1215 450 -1215 0 net=2984
rlabel metal2 604 -1215 604 -1215 0 net=3217
rlabel metal2 779 -1215 779 -1215 0 net=4409
rlabel metal2 12 -1217 12 -1217 0 net=511
rlabel metal2 436 -1217 436 -1217 0 net=2243
rlabel metal2 453 -1217 453 -1217 0 net=3956
rlabel metal2 79 -1219 79 -1219 0 net=1545
rlabel metal2 464 -1219 464 -1219 0 net=5282
rlabel metal2 86 -1221 86 -1221 0 net=2367
rlabel metal2 163 -1221 163 -1221 0 net=1473
rlabel metal2 226 -1221 226 -1221 0 net=1009
rlabel metal2 520 -1221 520 -1221 0 net=2755
rlabel metal2 583 -1221 583 -1221 0 net=3555
rlabel metal2 93 -1223 93 -1223 0 net=2078
rlabel metal2 233 -1223 233 -1223 0 net=1697
rlabel metal2 467 -1223 467 -1223 0 net=784
rlabel metal2 656 -1223 656 -1223 0 net=5160
rlabel metal2 37 -1225 37 -1225 0 net=1979
rlabel metal2 233 -1225 233 -1225 0 net=1451
rlabel metal2 474 -1225 474 -1225 0 net=2765
rlabel metal2 527 -1225 527 -1225 0 net=2761
rlabel metal2 541 -1225 541 -1225 0 net=697
rlabel metal2 93 -1227 93 -1227 0 net=3378
rlabel metal2 635 -1227 635 -1227 0 net=4145
rlabel metal2 877 -1227 877 -1227 0 net=4945
rlabel metal2 96 -1229 96 -1229 0 net=1583
rlabel metal2 170 -1229 170 -1229 0 net=3019
rlabel metal2 275 -1229 275 -1229 0 net=3789
rlabel metal2 758 -1229 758 -1229 0 net=4917
rlabel metal2 877 -1229 877 -1229 0 net=5373
rlabel metal2 96 -1231 96 -1231 0 net=3233
rlabel metal2 401 -1231 401 -1231 0 net=2197
rlabel metal2 471 -1231 471 -1231 0 net=2603
rlabel metal2 544 -1231 544 -1231 0 net=4525
rlabel metal2 100 -1233 100 -1233 0 net=1041
rlabel metal2 285 -1233 285 -1233 0 net=2930
rlabel metal2 555 -1233 555 -1233 0 net=2915
rlabel metal2 639 -1233 639 -1233 0 net=3397
rlabel metal2 863 -1233 863 -1233 0 net=4657
rlabel metal2 103 -1235 103 -1235 0 net=3662
rlabel metal2 107 -1237 107 -1237 0 net=1897
rlabel metal2 128 -1237 128 -1237 0 net=1199
rlabel metal2 296 -1237 296 -1237 0 net=2135
rlabel metal2 457 -1237 457 -1237 0 net=2585
rlabel metal2 583 -1237 583 -1237 0 net=3099
rlabel metal2 597 -1237 597 -1237 0 net=3301
rlabel metal2 44 -1239 44 -1239 0 net=2063
rlabel metal2 149 -1239 149 -1239 0 net=1045
rlabel metal2 296 -1239 296 -1239 0 net=1935
rlabel metal2 394 -1239 394 -1239 0 net=3383
rlabel metal2 646 -1239 646 -1239 0 net=3925
rlabel metal2 110 -1241 110 -1241 0 net=1170
rlabel metal2 303 -1241 303 -1241 0 net=25
rlabel metal2 457 -1241 457 -1241 0 net=3864
rlabel metal2 114 -1243 114 -1243 0 net=2123
rlabel metal2 604 -1243 604 -1243 0 net=3883
rlabel metal2 51 -1245 51 -1245 0 net=1667
rlabel metal2 184 -1245 184 -1245 0 net=1787
rlabel metal2 338 -1245 338 -1245 0 net=2405
rlabel metal2 471 -1245 471 -1245 0 net=546
rlabel metal2 51 -1247 51 -1247 0 net=2875
rlabel metal2 345 -1247 345 -1247 0 net=2153
rlabel metal2 478 -1247 478 -1247 0 net=4901
rlabel metal2 191 -1249 191 -1249 0 net=2001
rlabel metal2 261 -1249 261 -1249 0 net=1917
rlabel metal2 380 -1249 380 -1249 0 net=4389
rlabel metal2 607 -1249 607 -1249 0 net=5042
rlabel metal2 891 -1249 891 -1249 0 net=5127
rlabel metal2 212 -1251 212 -1251 0 net=3441
rlabel metal2 835 -1251 835 -1251 0 net=4475
rlabel metal2 289 -1253 289 -1253 0 net=2235
rlabel metal2 443 -1253 443 -1253 0 net=2515
rlabel metal2 492 -1253 492 -1253 0 net=3987
rlabel metal2 310 -1255 310 -1255 0 net=4375
rlabel metal2 387 -1257 387 -1257 0 net=2417
rlabel metal2 443 -1257 443 -1257 0 net=3175
rlabel metal2 513 -1257 513 -1257 0 net=2719
rlabel metal2 600 -1257 600 -1257 0 net=4227
rlabel metal2 282 -1259 282 -1259 0 net=1357
rlabel metal2 513 -1259 513 -1259 0 net=2857
rlabel metal2 611 -1259 611 -1259 0 net=3297
rlabel metal2 611 -1259 611 -1259 0 net=3297
rlabel metal2 646 -1259 646 -1259 0 net=2783
rlabel metal2 240 -1261 240 -1261 0 net=1461
rlabel metal2 548 -1261 548 -1261 0 net=3137
rlabel metal2 656 -1261 656 -1261 0 net=5242
rlabel metal2 40 -1263 40 -1263 0 net=2035
rlabel metal2 569 -1263 569 -1263 0 net=4705
rlabel metal2 660 -1265 660 -1265 0 net=3429
rlabel metal2 660 -1267 660 -1267 0 net=3719
rlabel metal2 124 -1269 124 -1269 0 net=3521
rlabel metal2 667 -1271 667 -1271 0 net=3519
rlabel metal2 670 -1273 670 -1273 0 net=5003
rlabel metal2 9 -1284 9 -1284 0 net=1266
rlabel metal2 37 -1284 37 -1284 0 net=1047
rlabel metal2 170 -1284 170 -1284 0 net=1743
rlabel metal2 222 -1284 222 -1284 0 net=2236
rlabel metal2 310 -1284 310 -1284 0 net=2124
rlabel metal2 579 -1284 579 -1284 0 net=3556
rlabel metal2 943 -1284 943 -1284 0 net=4616
rlabel metal2 30 -1286 30 -1286 0 net=2890
rlabel metal2 723 -1286 723 -1286 0 net=4441
rlabel metal2 723 -1286 723 -1286 0 net=4441
rlabel metal2 772 -1286 772 -1286 0 net=3895
rlabel metal2 772 -1286 772 -1286 0 net=3895
rlabel metal2 971 -1286 971 -1286 0 net=2482
rlabel metal2 44 -1288 44 -1288 0 net=2064
rlabel metal2 226 -1288 226 -1288 0 net=1010
rlabel metal2 509 -1288 509 -1288 0 net=3302
rlabel metal2 940 -1288 940 -1288 0 net=3005
rlabel metal2 44 -1290 44 -1290 0 net=2369
rlabel metal2 89 -1290 89 -1290 0 net=820
rlabel metal2 457 -1290 457 -1290 0 net=2605
rlabel metal2 569 -1290 569 -1290 0 net=3960
rlabel metal2 51 -1292 51 -1292 0 net=2876
rlabel metal2 408 -1292 408 -1292 0 net=2136
rlabel metal2 446 -1292 446 -1292 0 net=1267
rlabel metal2 499 -1292 499 -1292 0 net=3398
rlabel metal2 954 -1292 954 -1292 0 net=2189
rlabel metal2 51 -1294 51 -1294 0 net=3197
rlabel metal2 124 -1294 124 -1294 0 net=405
rlabel metal2 240 -1294 240 -1294 0 net=2037
rlabel metal2 310 -1294 310 -1294 0 net=1213
rlabel metal2 352 -1294 352 -1294 0 net=2615
rlabel metal2 569 -1294 569 -1294 0 net=3101
rlabel metal2 597 -1294 597 -1294 0 net=3299
rlabel metal2 618 -1294 618 -1294 0 net=4706
rlabel metal2 58 -1296 58 -1296 0 net=2206
rlabel metal2 184 -1296 184 -1296 0 net=3430
rlabel metal2 919 -1296 919 -1296 0 net=4102
rlabel metal2 61 -1298 61 -1298 0 net=1659
rlabel metal2 135 -1298 135 -1298 0 net=1849
rlabel metal2 198 -1298 198 -1298 0 net=1474
rlabel metal2 229 -1298 229 -1298 0 net=5175
rlabel metal2 65 -1300 65 -1300 0 net=2645
rlabel metal2 387 -1300 387 -1300 0 net=2419
rlabel metal2 411 -1300 411 -1300 0 net=4526
rlabel metal2 65 -1302 65 -1302 0 net=359
rlabel metal2 387 -1302 387 -1302 0 net=2721
rlabel metal2 576 -1302 576 -1302 0 net=4562
rlabel metal2 72 -1304 72 -1304 0 net=2438
rlabel metal2 149 -1304 149 -1304 0 net=1919
rlabel metal2 282 -1304 282 -1304 0 net=1462
rlabel metal2 415 -1304 415 -1304 0 net=1358
rlabel metal2 467 -1304 467 -1304 0 net=868
rlabel metal2 502 -1304 502 -1304 0 net=3059
rlabel metal2 632 -1304 632 -1304 0 net=3721
rlabel metal2 667 -1304 667 -1304 0 net=4476
rlabel metal2 898 -1304 898 -1304 0 net=5457
rlabel metal2 16 -1306 16 -1306 0 net=1521
rlabel metal2 296 -1306 296 -1306 0 net=1937
rlabel metal2 366 -1306 366 -1306 0 net=1858
rlabel metal2 471 -1306 471 -1306 0 net=3926
rlabel metal2 16 -1308 16 -1308 0 net=1793
rlabel metal2 114 -1308 114 -1308 0 net=1669
rlabel metal2 163 -1308 163 -1308 0 net=1585
rlabel metal2 303 -1308 303 -1308 0 net=3479
rlabel metal2 474 -1308 474 -1308 0 net=2784
rlabel metal2 653 -1308 653 -1308 0 net=5381
rlabel metal2 72 -1310 72 -1310 0 net=3442
rlabel metal2 793 -1310 793 -1310 0 net=4411
rlabel metal2 12 -1312 12 -1312 0 net=4211
rlabel metal2 93 -1314 93 -1314 0 net=1251
rlabel metal2 548 -1314 548 -1314 0 net=3139
rlabel metal2 646 -1314 646 -1314 0 net=3541
rlabel metal2 114 -1316 114 -1316 0 net=1899
rlabel metal2 128 -1316 128 -1316 0 net=2909
rlabel metal2 317 -1316 317 -1316 0 net=1699
rlabel metal2 331 -1316 331 -1316 0 net=3235
rlabel metal2 653 -1316 653 -1316 0 net=3523
rlabel metal2 709 -1316 709 -1316 0 net=4377
rlabel metal2 121 -1318 121 -1318 0 net=2916
rlabel metal2 656 -1318 656 -1318 0 net=4428
rlabel metal2 156 -1320 156 -1320 0 net=1201
rlabel metal2 177 -1320 177 -1320 0 net=3021
rlabel metal2 415 -1320 415 -1320 0 net=2211
rlabel metal2 142 -1322 142 -1322 0 net=2311
rlabel metal2 191 -1322 191 -1322 0 net=2003
rlabel metal2 208 -1322 208 -1322 0 net=2647
rlabel metal2 534 -1322 534 -1322 0 net=2763
rlabel metal2 590 -1322 590 -1322 0 net=4391
rlabel metal2 667 -1322 667 -1322 0 net=4147
rlabel metal2 835 -1322 835 -1322 0 net=4947
rlabel metal2 100 -1324 100 -1324 0 net=1042
rlabel metal2 212 -1324 212 -1324 0 net=2439
rlabel metal2 313 -1324 313 -1324 0 net=5403
rlabel metal2 625 -1324 625 -1324 0 net=3403
rlabel metal2 688 -1324 688 -1324 0 net=3989
rlabel metal2 100 -1326 100 -1326 0 net=3093
rlabel metal2 233 -1326 233 -1326 0 net=1452
rlabel metal2 429 -1326 429 -1326 0 net=3001
rlabel metal2 674 -1326 674 -1326 0 net=3219
rlabel metal2 142 -1328 142 -1328 0 net=2587
rlabel metal2 562 -1328 562 -1328 0 net=2757
rlabel metal2 702 -1328 702 -1328 0 net=4109
rlabel metal2 233 -1330 233 -1330 0 net=2199
rlabel metal2 432 -1330 432 -1330 0 net=3158
rlabel metal2 240 -1332 240 -1332 0 net=1393
rlabel metal2 436 -1332 436 -1332 0 net=2245
rlabel metal2 460 -1332 460 -1332 0 net=4989
rlabel metal2 247 -1334 247 -1334 0 net=1468
rlabel metal2 394 -1334 394 -1334 0 net=2407
rlabel metal2 443 -1334 443 -1334 0 net=4923
rlabel metal2 205 -1336 205 -1336 0 net=1981
rlabel metal2 254 -1336 254 -1336 0 net=2155
rlabel metal2 366 -1336 366 -1336 0 net=2053
rlabel metal2 443 -1336 443 -1336 0 net=2517
rlabel metal2 481 -1336 481 -1336 0 net=3520
rlabel metal2 303 -1338 303 -1338 0 net=2011
rlabel metal2 450 -1338 450 -1338 0 net=2766
rlabel metal2 527 -1338 527 -1338 0 net=3415
rlabel metal2 716 -1338 716 -1338 0 net=3885
rlabel metal2 765 -1338 765 -1338 0 net=4335
rlabel metal2 877 -1338 877 -1338 0 net=5375
rlabel metal2 338 -1340 338 -1340 0 net=2381
rlabel metal2 478 -1340 478 -1340 0 net=2779
rlabel metal2 639 -1340 639 -1340 0 net=3385
rlabel metal2 814 -1340 814 -1340 0 net=5361
rlabel metal2 338 -1342 338 -1342 0 net=1877
rlabel metal2 383 -1342 383 -1342 0 net=4753
rlabel metal2 814 -1342 814 -1342 0 net=4543
rlabel metal2 268 -1344 268 -1344 0 net=1290
rlabel metal2 485 -1344 485 -1344 0 net=3177
rlabel metal2 737 -1344 737 -1344 0 net=4639
rlabel metal2 800 -1344 800 -1344 0 net=5073
rlabel metal2 268 -1346 268 -1346 0 net=1789
rlabel metal2 513 -1346 513 -1346 0 net=2859
rlabel metal2 639 -1346 639 -1346 0 net=3791
rlabel metal2 758 -1346 758 -1346 0 net=4919
rlabel metal2 828 -1346 828 -1346 0 net=4903
rlabel metal2 79 -1348 79 -1348 0 net=1547
rlabel metal2 485 -1348 485 -1348 0 net=4519
rlabel metal2 758 -1348 758 -1348 0 net=5233
rlabel metal2 79 -1350 79 -1350 0 net=2559
rlabel metal2 695 -1350 695 -1350 0 net=4079
rlabel metal2 513 -1352 513 -1352 0 net=4266
rlabel metal2 520 -1354 520 -1354 0 net=2741
rlabel metal2 737 -1354 737 -1354 0 net=4229
rlabel metal2 842 -1354 842 -1354 0 net=5005
rlabel metal2 821 -1356 821 -1356 0 net=4659
rlabel metal2 870 -1358 870 -1358 0 net=5129
rlabel metal2 2 -1369 2 -1369 0 net=2371
rlabel metal2 58 -1369 58 -1369 0 net=2561
rlabel metal2 86 -1369 86 -1369 0 net=1671
rlabel metal2 156 -1369 156 -1369 0 net=2646
rlabel metal2 376 -1369 376 -1369 0 net=3896
rlabel metal2 856 -1369 856 -1369 0 net=5075
rlabel metal2 908 -1369 908 -1369 0 net=2190
rlabel metal2 971 -1369 971 -1369 0 net=3006
rlabel metal2 9 -1371 9 -1371 0 net=3022
rlabel metal2 394 -1371 394 -1371 0 net=3178
rlabel metal2 712 -1371 712 -1371 0 net=3886
rlabel metal2 765 -1371 765 -1371 0 net=4337
rlabel metal2 947 -1371 947 -1371 0 net=2851
rlabel metal2 9 -1373 9 -1373 0 net=4212
rlabel metal2 765 -1373 765 -1373 0 net=5459
rlabel metal2 912 -1373 912 -1373 0 net=3221
rlabel metal2 37 -1375 37 -1375 0 net=1048
rlabel metal2 240 -1375 240 -1375 0 net=1394
rlabel metal2 397 -1375 397 -1375 0 net=2420
rlabel metal2 450 -1375 450 -1375 0 net=962
rlabel metal2 467 -1375 467 -1375 0 net=5234
rlabel metal2 856 -1375 856 -1375 0 net=5131
rlabel metal2 891 -1375 891 -1375 0 net=5383
rlabel metal2 37 -1377 37 -1377 0 net=3559
rlabel metal2 198 -1377 198 -1377 0 net=2005
rlabel metal2 198 -1377 198 -1377 0 net=2005
rlabel metal2 205 -1377 205 -1377 0 net=1878
rlabel metal2 348 -1377 348 -1377 0 net=4279
rlabel metal2 744 -1377 744 -1377 0 net=4521
rlabel metal2 800 -1377 800 -1377 0 net=4921
rlabel metal2 51 -1379 51 -1379 0 net=3199
rlabel metal2 401 -1379 401 -1379 0 net=2382
rlabel metal2 478 -1379 478 -1379 0 net=3524
rlabel metal2 681 -1379 681 -1379 0 net=4081
rlabel metal2 702 -1379 702 -1379 0 net=4111
rlabel metal2 800 -1379 800 -1379 0 net=4661
rlabel metal2 849 -1379 849 -1379 0 net=4991
rlabel metal2 51 -1381 51 -1381 0 net=1791
rlabel metal2 275 -1381 275 -1381 0 net=1549
rlabel metal2 275 -1381 275 -1381 0 net=1549
rlabel metal2 296 -1381 296 -1381 0 net=2440
rlabel metal2 401 -1381 401 -1381 0 net=2861
rlabel metal2 576 -1381 576 -1381 0 net=3300
rlabel metal2 604 -1381 604 -1381 0 net=4904
rlabel metal2 842 -1381 842 -1381 0 net=5007
rlabel metal2 863 -1381 863 -1381 0 net=5177
rlabel metal2 65 -1383 65 -1383 0 net=157
rlabel metal2 191 -1383 191 -1383 0 net=4317
rlabel metal2 807 -1383 807 -1383 0 net=4925
rlabel metal2 863 -1383 863 -1383 0 net=4899
rlabel metal2 33 -1385 33 -1385 0 net=3635
rlabel metal2 72 -1385 72 -1385 0 net=915
rlabel metal2 555 -1385 555 -1385 0 net=3003
rlabel metal2 702 -1385 702 -1385 0 net=4231
rlabel metal2 72 -1387 72 -1387 0 net=2607
rlabel metal2 464 -1387 464 -1387 0 net=3975
rlabel metal2 590 -1387 590 -1387 0 net=5405
rlabel metal2 79 -1389 79 -1389 0 net=2473
rlabel metal2 338 -1389 338 -1389 0 net=1268
rlabel metal2 516 -1389 516 -1389 0 net=3990
rlabel metal2 723 -1389 723 -1389 0 net=4443
rlabel metal2 89 -1391 89 -1391 0 net=3060
rlabel metal2 593 -1391 593 -1391 0 net=5362
rlabel metal2 93 -1393 93 -1393 0 net=1253
rlabel metal2 226 -1393 226 -1393 0 net=1985
rlabel metal2 569 -1393 569 -1393 0 net=3103
rlabel metal2 604 -1393 604 -1393 0 net=4849
rlabel metal2 877 -1393 877 -1393 0 net=5377
rlabel metal2 93 -1395 93 -1395 0 net=1901
rlabel metal2 124 -1395 124 -1395 0 net=3386
rlabel metal2 835 -1395 835 -1395 0 net=4949
rlabel metal2 100 -1397 100 -1397 0 net=3094
rlabel metal2 667 -1397 667 -1397 0 net=4149
rlabel metal2 709 -1397 709 -1397 0 net=4379
rlabel metal2 751 -1397 751 -1397 0 net=4413
rlabel metal2 835 -1397 835 -1397 0 net=4867
rlabel metal2 23 -1399 23 -1399 0 net=1613
rlabel metal2 128 -1399 128 -1399 0 net=2911
rlabel metal2 310 -1399 310 -1399 0 net=1214
rlabel metal2 453 -1399 453 -1399 0 net=4189
rlabel metal2 779 -1399 779 -1399 0 net=4755
rlabel metal2 943 -1399 943 -1399 0 net=4647
rlabel metal2 23 -1401 23 -1401 0 net=2157
rlabel metal2 261 -1401 261 -1401 0 net=1522
rlabel metal2 373 -1401 373 -1401 0 net=3833
rlabel metal2 121 -1403 121 -1403 0 net=3181
rlabel metal2 478 -1403 478 -1403 0 net=2617
rlabel metal2 527 -1403 527 -1403 0 net=4640
rlabel metal2 121 -1405 121 -1405 0 net=295
rlabel metal2 233 -1405 233 -1405 0 net=2201
rlabel metal2 471 -1405 471 -1405 0 net=3481
rlabel metal2 530 -1405 530 -1405 0 net=2758
rlabel metal2 786 -1405 786 -1405 0 net=4545
rlabel metal2 135 -1407 135 -1407 0 net=2039
rlabel metal2 310 -1407 310 -1407 0 net=1701
rlabel metal2 331 -1407 331 -1407 0 net=3007
rlabel metal2 646 -1407 646 -1407 0 net=3543
rlabel metal2 149 -1409 149 -1409 0 net=1921
rlabel metal2 289 -1409 289 -1409 0 net=2055
rlabel metal2 390 -1409 390 -1409 0 net=1067
rlabel metal2 481 -1409 481 -1409 0 net=4599
rlabel metal2 107 -1411 107 -1411 0 net=1661
rlabel metal2 159 -1411 159 -1411 0 net=3037
rlabel metal2 247 -1411 247 -1411 0 net=1982
rlabel metal2 366 -1411 366 -1411 0 net=2723
rlabel metal2 485 -1411 485 -1411 0 net=2764
rlabel metal2 632 -1411 632 -1411 0 net=3723
rlabel metal2 660 -1411 660 -1411 0 net=4393
rlabel metal2 30 -1413 30 -1413 0 net=4003
rlabel metal2 166 -1413 166 -1413 0 net=1945
rlabel metal2 219 -1413 219 -1413 0 net=2443
rlabel metal2 233 -1413 233 -1413 0 net=1033
rlabel metal2 537 -1413 537 -1413 0 net=3404
rlabel metal2 632 -1413 632 -1413 0 net=4583
rlabel metal2 107 -1415 107 -1415 0 net=1453
rlabel metal2 170 -1415 170 -1415 0 net=1745
rlabel metal2 317 -1415 317 -1415 0 net=1141
rlabel metal2 492 -1415 492 -1415 0 net=2649
rlabel metal2 513 -1415 513 -1415 0 net=2743
rlabel metal2 534 -1415 534 -1415 0 net=2781
rlabel metal2 639 -1415 639 -1415 0 net=3793
rlabel metal2 16 -1417 16 -1417 0 net=1794
rlabel metal2 541 -1417 541 -1417 0 net=3417
rlabel metal2 16 -1419 16 -1419 0 net=2013
rlabel metal2 464 -1419 464 -1419 0 net=2751
rlabel metal2 541 -1419 541 -1419 0 net=3141
rlabel metal2 163 -1421 163 -1421 0 net=1203
rlabel metal2 177 -1421 177 -1421 0 net=2313
rlabel metal2 254 -1421 254 -1421 0 net=1939
rlabel metal2 488 -1421 488 -1421 0 net=3619
rlabel metal2 128 -1423 128 -1423 0 net=1085
rlabel metal2 184 -1423 184 -1423 0 net=1851
rlabel metal2 499 -1423 499 -1423 0 net=3237
rlabel metal2 212 -1425 212 -1425 0 net=2903
rlabel metal2 509 -1425 509 -1425 0 net=3255
rlabel metal2 282 -1427 282 -1427 0 net=1587
rlabel metal2 579 -1427 579 -1427 0 net=3571
rlabel metal2 282 -1429 282 -1429 0 net=2213
rlabel metal2 579 -1429 579 -1429 0 net=5315
rlabel metal2 415 -1431 415 -1431 0 net=2409
rlabel metal2 422 -1433 422 -1433 0 net=2247
rlabel metal2 436 -1435 436 -1435 0 net=2519
rlabel metal2 142 -1437 142 -1437 0 net=2589
rlabel metal2 9 -1448 9 -1448 0 net=2015
rlabel metal2 23 -1448 23 -1448 0 net=2158
rlabel metal2 432 -1448 432 -1448 0 net=2752
rlabel metal2 548 -1448 548 -1448 0 net=4922
rlabel metal2 940 -1448 940 -1448 0 net=3223
rlabel metal2 16 -1450 16 -1450 0 net=1987
rlabel metal2 282 -1450 282 -1450 0 net=2215
rlabel metal2 457 -1450 457 -1450 0 net=3239
rlabel metal2 502 -1450 502 -1450 0 net=4112
rlabel metal2 800 -1450 800 -1450 0 net=4663
rlabel metal2 800 -1450 800 -1450 0 net=4663
rlabel metal2 856 -1450 856 -1450 0 net=5133
rlabel metal2 856 -1450 856 -1450 0 net=5133
rlabel metal2 961 -1450 961 -1450 0 net=4648
rlabel metal2 23 -1452 23 -1452 0 net=3560
rlabel metal2 44 -1452 44 -1452 0 net=1455
rlabel metal2 114 -1452 114 -1452 0 net=1245
rlabel metal2 285 -1452 285 -1452 0 net=2744
rlabel metal2 555 -1452 555 -1452 0 net=4950
rlabel metal2 982 -1452 982 -1452 0 net=3875
rlabel metal2 51 -1454 51 -1454 0 net=1792
rlabel metal2 373 -1454 373 -1454 0 net=2411
rlabel metal2 432 -1454 432 -1454 0 net=924
rlabel metal2 506 -1454 506 -1454 0 net=4900
rlabel metal2 51 -1456 51 -1456 0 net=2631
rlabel metal2 558 -1456 558 -1456 0 net=4338
rlabel metal2 79 -1458 79 -1458 0 net=2474
rlabel metal2 604 -1458 604 -1458 0 net=4394
rlabel metal2 79 -1460 79 -1460 0 net=2941
rlabel metal2 303 -1460 303 -1460 0 net=2904
rlabel metal2 397 -1460 397 -1460 0 net=4873
rlabel metal2 93 -1462 93 -1462 0 net=1902
rlabel metal2 142 -1462 142 -1462 0 net=1852
rlabel metal2 338 -1462 338 -1462 0 net=1809
rlabel metal2 460 -1462 460 -1462 0 net=4600
rlabel metal2 93 -1464 93 -1464 0 net=1143
rlabel metal2 345 -1464 345 -1464 0 net=3183
rlabel metal2 576 -1464 576 -1464 0 net=3257
rlabel metal2 632 -1464 632 -1464 0 net=5076
rlabel metal2 100 -1466 100 -1466 0 net=1615
rlabel metal2 352 -1466 352 -1466 0 net=2724
rlabel metal2 376 -1466 376 -1466 0 net=3200
rlabel metal2 415 -1466 415 -1466 0 net=2249
rlabel metal2 467 -1466 467 -1466 0 net=4993
rlabel metal2 887 -1466 887 -1466 0 net=5393
rlabel metal2 905 -1466 905 -1466 0 net=5385
rlabel metal2 100 -1468 100 -1468 0 net=1829
rlabel metal2 422 -1468 422 -1468 0 net=2619
rlabel metal2 485 -1468 485 -1468 0 net=418
rlabel metal2 611 -1468 611 -1468 0 net=3795
rlabel metal2 688 -1468 688 -1468 0 net=4151
rlabel metal2 712 -1468 712 -1468 0 net=4584
rlabel metal2 912 -1468 912 -1468 0 net=5179
rlabel metal2 65 -1470 65 -1470 0 net=3637
rlabel metal2 688 -1470 688 -1470 0 net=4757
rlabel metal2 65 -1472 65 -1472 0 net=2609
rlabel metal2 117 -1472 117 -1472 0 net=1662
rlabel metal2 156 -1472 156 -1472 0 net=4190
rlabel metal2 793 -1472 793 -1472 0 net=4927
rlabel metal2 86 -1474 86 -1474 0 net=1672
rlabel metal2 159 -1474 159 -1474 0 net=2782
rlabel metal2 632 -1474 632 -1474 0 net=2207
rlabel metal2 653 -1474 653 -1474 0 net=4992
rlabel metal2 86 -1476 86 -1476 0 net=2963
rlabel metal2 198 -1476 198 -1476 0 net=2006
rlabel metal2 198 -1476 198 -1476 0 net=2006
rlabel metal2 201 -1476 201 -1476 0 net=1746
rlabel metal2 310 -1476 310 -1476 0 net=1703
rlabel metal2 310 -1476 310 -1476 0 net=1703
rlabel metal2 352 -1476 352 -1476 0 net=1907
rlabel metal2 467 -1476 467 -1476 0 net=3004
rlabel metal2 730 -1476 730 -1476 0 net=4445
rlabel metal2 821 -1476 821 -1476 0 net=5317
rlabel metal2 107 -1478 107 -1478 0 net=1029
rlabel metal2 471 -1478 471 -1478 0 net=1068
rlabel metal2 590 -1478 590 -1478 0 net=4083
rlabel metal2 695 -1478 695 -1478 0 net=4381
rlabel metal2 737 -1478 737 -1478 0 net=3829
rlabel metal2 58 -1480 58 -1480 0 net=2563
rlabel metal2 478 -1480 478 -1480 0 net=4318
rlabel metal2 842 -1480 842 -1480 0 net=5407
rlabel metal2 58 -1482 58 -1482 0 net=1035
rlabel metal2 240 -1482 240 -1482 0 net=3039
rlabel metal2 355 -1482 355 -1482 0 net=59
rlabel metal2 485 -1482 485 -1482 0 net=3143
rlabel metal2 597 -1482 597 -1482 0 net=3419
rlabel metal2 625 -1482 625 -1482 0 net=3931
rlabel metal2 681 -1482 681 -1482 0 net=4233
rlabel metal2 723 -1482 723 -1482 0 net=4415
rlabel metal2 765 -1482 765 -1482 0 net=5461
rlabel metal2 919 -1482 919 -1482 0 net=2853
rlabel metal2 121 -1484 121 -1484 0 net=1619
rlabel metal2 324 -1484 324 -1484 0 net=2985
rlabel metal2 597 -1484 597 -1484 0 net=3621
rlabel metal2 653 -1484 653 -1484 0 net=4281
rlabel metal2 744 -1484 744 -1484 0 net=4523
rlabel metal2 933 -1484 933 -1484 0 net=5207
rlabel metal2 128 -1486 128 -1486 0 net=1385
rlabel metal2 509 -1486 509 -1486 0 net=3544
rlabel metal2 702 -1486 702 -1486 0 net=4869
rlabel metal2 135 -1488 135 -1488 0 net=2041
rlabel metal2 443 -1488 443 -1488 0 net=2591
rlabel metal2 751 -1488 751 -1488 0 net=4547
rlabel metal2 835 -1488 835 -1488 0 net=5009
rlabel metal2 40 -1490 40 -1490 0 net=5099
rlabel metal2 142 -1492 142 -1492 0 net=1605
rlabel metal2 184 -1492 184 -1492 0 net=1957
rlabel metal2 366 -1492 366 -1492 0 net=2202
rlabel metal2 443 -1492 443 -1492 0 net=3315
rlabel metal2 537 -1492 537 -1492 0 net=4909
rlabel metal2 149 -1494 149 -1494 0 net=1940
rlabel metal2 261 -1494 261 -1494 0 net=1923
rlabel metal2 369 -1494 369 -1494 0 net=4557
rlabel metal2 786 -1494 786 -1494 0 net=4851
rlabel metal2 163 -1496 163 -1496 0 net=1204
rlabel metal2 173 -1496 173 -1496 0 net=1588
rlabel metal2 492 -1496 492 -1496 0 net=2651
rlabel metal2 537 -1496 537 -1496 0 net=4877
rlabel metal2 30 -1498 30 -1498 0 net=4004
rlabel metal2 184 -1498 184 -1498 0 net=3511
rlabel metal2 492 -1498 492 -1498 0 net=3483
rlabel metal2 618 -1498 618 -1498 0 net=3573
rlabel metal2 667 -1498 667 -1498 0 net=3835
rlabel metal2 807 -1498 807 -1498 0 net=5379
rlabel metal2 30 -1500 30 -1500 0 net=2057
rlabel metal2 359 -1500 359 -1500 0 net=3567
rlabel metal2 646 -1500 646 -1500 0 net=3725
rlabel metal2 152 -1502 152 -1502 0 net=3629
rlabel metal2 187 -1504 187 -1504 0 net=2314
rlabel metal2 261 -1504 261 -1504 0 net=1413
rlabel metal2 187 -1506 187 -1506 0 net=3008
rlabel metal2 191 -1508 191 -1508 0 net=1947
rlabel metal2 289 -1508 289 -1508 0 net=2579
rlabel metal2 562 -1508 562 -1508 0 net=3977
rlabel metal2 191 -1510 191 -1510 0 net=131
rlabel metal2 401 -1510 401 -1510 0 net=2863
rlabel metal2 562 -1510 562 -1510 0 net=3105
rlabel metal2 205 -1512 205 -1512 0 net=1255
rlabel metal2 401 -1512 401 -1512 0 net=2521
rlabel metal2 583 -1512 583 -1512 0 net=3207
rlabel metal2 166 -1514 166 -1514 0 net=2463
rlabel metal2 177 -1516 177 -1516 0 net=1087
rlabel metal2 219 -1516 219 -1516 0 net=2445
rlabel metal2 233 -1516 233 -1516 0 net=2331
rlabel metal2 177 -1518 177 -1518 0 net=1349
rlabel metal2 219 -1520 219 -1520 0 net=2912
rlabel metal2 240 -1522 240 -1522 0 net=1593
rlabel metal2 275 -1524 275 -1524 0 net=1551
rlabel metal2 2 -1526 2 -1526 0 net=2373
rlabel metal2 23 -1537 23 -1537 0 net=1319
rlabel metal2 44 -1537 44 -1537 0 net=1456
rlabel metal2 166 -1537 166 -1537 0 net=2580
rlabel metal2 306 -1537 306 -1537 0 net=2412
rlabel metal2 415 -1537 415 -1537 0 net=2251
rlabel metal2 415 -1537 415 -1537 0 net=2251
rlabel metal2 432 -1537 432 -1537 0 net=3144
rlabel metal2 509 -1537 509 -1537 0 net=5408
rlabel metal2 849 -1537 849 -1537 0 net=5101
rlabel metal2 947 -1537 947 -1537 0 net=4773
rlabel metal2 982 -1537 982 -1537 0 net=3877
rlabel metal2 30 -1539 30 -1539 0 net=2058
rlabel metal2 345 -1539 345 -1539 0 net=3040
rlabel metal2 373 -1539 373 -1539 0 net=2523
rlabel metal2 436 -1539 436 -1539 0 net=2464
rlabel metal2 884 -1539 884 -1539 0 net=3224
rlabel metal2 954 -1539 954 -1539 0 net=5208
rlabel metal2 16 -1541 16 -1541 0 net=1989
rlabel metal2 37 -1541 37 -1541 0 net=2374
rlabel metal2 282 -1541 282 -1541 0 net=3051
rlabel metal2 352 -1541 352 -1541 0 net=1909
rlabel metal2 478 -1541 478 -1541 0 net=4084
rlabel metal2 604 -1541 604 -1541 0 net=3421
rlabel metal2 898 -1541 898 -1541 0 net=5394
rlabel metal2 940 -1541 940 -1541 0 net=5391
rlabel metal2 16 -1543 16 -1543 0 net=4161
rlabel metal2 352 -1543 352 -1543 0 net=2043
rlabel metal2 401 -1543 401 -1543 0 net=3631
rlabel metal2 705 -1543 705 -1543 0 net=5462
rlabel metal2 800 -1543 800 -1543 0 net=4664
rlabel metal2 898 -1543 898 -1543 0 net=5181
rlabel metal2 37 -1545 37 -1545 0 net=1379
rlabel metal2 100 -1545 100 -1545 0 net=1830
rlabel metal2 142 -1545 142 -1545 0 net=1607
rlabel metal2 142 -1545 142 -1545 0 net=1607
rlabel metal2 149 -1545 149 -1545 0 net=3240
rlabel metal2 478 -1545 478 -1545 0 net=3484
rlabel metal2 520 -1545 520 -1545 0 net=3317
rlabel metal2 534 -1545 534 -1545 0 net=4446
rlabel metal2 733 -1545 733 -1545 0 net=5380
rlabel metal2 814 -1545 814 -1545 0 net=4879
rlabel metal2 44 -1547 44 -1547 0 net=1387
rlabel metal2 135 -1547 135 -1547 0 net=721
rlabel metal2 436 -1547 436 -1547 0 net=2595
rlabel metal2 485 -1547 485 -1547 0 net=2865
rlabel metal2 586 -1547 586 -1547 0 net=2592
rlabel metal2 723 -1547 723 -1547 0 net=4417
rlabel metal2 723 -1547 723 -1547 0 net=4417
rlabel metal2 814 -1547 814 -1547 0 net=5387
rlabel metal2 9 -1549 9 -1549 0 net=2016
rlabel metal2 492 -1549 492 -1549 0 net=2208
rlabel metal2 646 -1549 646 -1549 0 net=4383
rlabel metal2 716 -1549 716 -1549 0 net=4549
rlabel metal2 65 -1551 65 -1551 0 net=2610
rlabel metal2 446 -1551 446 -1551 0 net=4152
rlabel metal2 751 -1551 751 -1551 0 net=5319
rlabel metal2 65 -1553 65 -1553 0 net=3599
rlabel metal2 194 -1553 194 -1553 0 net=3622
rlabel metal2 604 -1553 604 -1553 0 net=4283
rlabel metal2 709 -1553 709 -1553 0 net=4995
rlabel metal2 86 -1555 86 -1555 0 net=2965
rlabel metal2 408 -1555 408 -1555 0 net=2565
rlabel metal2 520 -1555 520 -1555 0 net=3259
rlabel metal2 590 -1555 590 -1555 0 net=4759
rlabel metal2 86 -1557 86 -1557 0 net=3579
rlabel metal2 114 -1557 114 -1557 0 net=1246
rlabel metal2 555 -1557 555 -1557 0 net=4743
rlabel metal2 618 -1557 618 -1557 0 net=3569
rlabel metal2 93 -1559 93 -1559 0 net=1144
rlabel metal2 450 -1559 450 -1559 0 net=3830
rlabel metal2 100 -1561 100 -1561 0 net=4487
rlabel metal2 341 -1561 341 -1561 0 net=5219
rlabel metal2 107 -1563 107 -1563 0 net=1030
rlabel metal2 369 -1563 369 -1563 0 net=3485
rlabel metal2 453 -1563 453 -1563 0 net=4524
rlabel metal2 58 -1565 58 -1565 0 net=1036
rlabel metal2 457 -1565 457 -1565 0 net=2653
rlabel metal2 530 -1565 530 -1565 0 net=4177
rlabel metal2 632 -1565 632 -1565 0 net=3639
rlabel metal2 688 -1565 688 -1565 0 net=4871
rlabel metal2 744 -1565 744 -1565 0 net=5011
rlabel metal2 58 -1567 58 -1567 0 net=4957
rlabel metal2 702 -1567 702 -1567 0 net=2854
rlabel metal2 128 -1569 128 -1569 0 net=1959
rlabel metal2 411 -1569 411 -1569 0 net=4465
rlabel metal2 660 -1569 660 -1569 0 net=4235
rlabel metal2 880 -1569 880 -1569 0 net=4985
rlabel metal2 135 -1571 135 -1571 0 net=1089
rlabel metal2 212 -1571 212 -1571 0 net=1257
rlabel metal2 261 -1571 261 -1571 0 net=1415
rlabel metal2 282 -1571 282 -1571 0 net=1925
rlabel metal2 331 -1571 331 -1571 0 net=4935
rlabel metal2 513 -1571 513 -1571 0 net=3185
rlabel metal2 75 -1573 75 -1573 0 net=1381
rlabel metal2 289 -1573 289 -1573 0 net=4033
rlabel metal2 534 -1573 534 -1573 0 net=4489
rlabel metal2 149 -1575 149 -1575 0 net=2657
rlabel metal2 429 -1575 429 -1575 0 net=3229
rlabel metal2 548 -1575 548 -1575 0 net=3107
rlabel metal2 156 -1577 156 -1577 0 net=1948
rlabel metal2 303 -1577 303 -1577 0 net=1617
rlabel metal2 324 -1577 324 -1577 0 net=2987
rlabel metal2 562 -1577 562 -1577 0 net=4558
rlabel metal2 156 -1579 156 -1579 0 net=4928
rlabel metal2 159 -1581 159 -1581 0 net=3061
rlabel metal2 317 -1581 317 -1581 0 net=2217
rlabel metal2 429 -1581 429 -1581 0 net=3679
rlabel metal2 765 -1581 765 -1581 0 net=4911
rlabel metal2 72 -1583 72 -1583 0 net=3457
rlabel metal2 793 -1583 793 -1583 0 net=5135
rlabel metal2 72 -1585 72 -1585 0 net=1595
rlabel metal2 247 -1585 247 -1585 0 net=1553
rlabel metal2 362 -1585 362 -1585 0 net=5339
rlabel metal2 177 -1587 177 -1587 0 net=3796
rlabel metal2 177 -1589 177 -1589 0 net=3837
rlabel metal2 198 -1591 198 -1591 0 net=1351
rlabel metal2 296 -1591 296 -1591 0 net=1811
rlabel metal2 362 -1591 362 -1591 0 net=2620
rlabel metal2 569 -1591 569 -1591 0 net=3979
rlabel metal2 674 -1591 674 -1591 0 net=4875
rlabel metal2 173 -1593 173 -1593 0 net=2819
rlabel metal2 338 -1593 338 -1593 0 net=3932
rlabel metal2 201 -1595 201 -1595 0 net=3117
rlabel metal2 240 -1595 240 -1595 0 net=3075
rlabel metal2 569 -1595 569 -1595 0 net=3575
rlabel metal2 215 -1597 215 -1597 0 net=2446
rlabel metal2 639 -1597 639 -1597 0 net=3727
rlabel metal2 226 -1599 226 -1599 0 net=1705
rlabel metal2 506 -1599 506 -1599 0 net=4339
rlabel metal2 667 -1599 667 -1599 0 net=5253
rlabel metal2 233 -1601 233 -1601 0 net=2333
rlabel metal2 506 -1601 506 -1601 0 net=3209
rlabel metal2 51 -1603 51 -1603 0 net=2633
rlabel metal2 523 -1603 523 -1603 0 net=1
rlabel metal2 51 -1605 51 -1605 0 net=2943
rlabel metal2 537 -1605 537 -1605 0 net=4852
rlabel metal2 26 -1607 26 -1607 0 net=5169
rlabel metal2 79 -1609 79 -1609 0 net=1621
rlabel metal2 121 -1611 121 -1611 0 net=5043
rlabel metal2 9 -1622 9 -1622 0 net=1320
rlabel metal2 30 -1622 30 -1622 0 net=1991
rlabel metal2 124 -1622 124 -1622 0 net=4490
rlabel metal2 695 -1622 695 -1622 0 net=4958
rlabel metal2 943 -1622 943 -1622 0 net=3333
rlabel metal2 971 -1622 971 -1622 0 net=5392
rlabel metal2 9 -1624 9 -1624 0 net=3077
rlabel metal2 247 -1624 247 -1624 0 net=1555
rlabel metal2 289 -1624 289 -1624 0 net=3053
rlabel metal2 390 -1624 390 -1624 0 net=4575
rlabel metal2 793 -1624 793 -1624 0 net=5136
rlabel metal2 877 -1624 877 -1624 0 net=5182
rlabel metal2 912 -1624 912 -1624 0 net=4987
rlabel metal2 975 -1624 975 -1624 0 net=3878
rlabel metal2 16 -1626 16 -1626 0 net=4162
rlabel metal2 240 -1626 240 -1626 0 net=1813
rlabel metal2 299 -1626 299 -1626 0 net=4466
rlabel metal2 660 -1626 660 -1626 0 net=4236
rlabel metal2 712 -1626 712 -1626 0 net=4912
rlabel metal2 835 -1626 835 -1626 0 net=5341
rlabel metal2 894 -1626 894 -1626 0 net=5102
rlabel metal2 16 -1628 16 -1628 0 net=847
rlabel metal2 93 -1628 93 -1628 0 net=4340
rlabel metal2 639 -1628 639 -1628 0 net=3729
rlabel metal2 926 -1628 926 -1628 0 net=4775
rlabel metal2 23 -1630 23 -1630 0 net=2395
rlabel metal2 100 -1630 100 -1630 0 net=4488
rlabel metal2 247 -1630 247 -1630 0 net=2335
rlabel metal2 341 -1630 341 -1630 0 net=47
rlabel metal2 723 -1630 723 -1630 0 net=4418
rlabel metal2 842 -1630 842 -1630 0 net=4880
rlabel metal2 30 -1632 30 -1632 0 net=1955
rlabel metal2 303 -1632 303 -1632 0 net=1618
rlabel metal2 341 -1632 341 -1632 0 net=3640
rlabel metal2 660 -1632 660 -1632 0 net=5012
rlabel metal2 828 -1632 828 -1632 0 net=5221
rlabel metal2 37 -1634 37 -1634 0 net=1380
rlabel metal2 93 -1634 93 -1634 0 net=1575
rlabel metal2 163 -1634 163 -1634 0 net=3849
rlabel metal2 667 -1634 667 -1634 0 net=5321
rlabel metal2 37 -1636 37 -1636 0 net=4085
rlabel metal2 439 -1636 439 -1636 0 net=3779
rlabel metal2 716 -1636 716 -1636 0 net=4551
rlabel metal2 44 -1638 44 -1638 0 net=1388
rlabel metal2 331 -1638 331 -1638 0 net=4937
rlabel metal2 44 -1640 44 -1640 0 net=2945
rlabel metal2 58 -1640 58 -1640 0 net=3580
rlabel metal2 107 -1640 107 -1640 0 net=1707
rlabel metal2 303 -1640 303 -1640 0 net=1291
rlabel metal2 404 -1640 404 -1640 0 net=4895
rlabel metal2 51 -1642 51 -1642 0 net=1259
rlabel metal2 226 -1642 226 -1642 0 net=1655
rlabel metal2 348 -1642 348 -1642 0 net=2524
rlabel metal2 383 -1642 383 -1642 0 net=4181
rlabel metal2 86 -1644 86 -1644 0 net=2087
rlabel metal2 110 -1644 110 -1644 0 net=2988
rlabel metal2 359 -1644 359 -1644 0 net=2967
rlabel metal2 387 -1644 387 -1644 0 net=3680
rlabel metal2 450 -1644 450 -1644 0 net=4529
rlabel metal2 128 -1646 128 -1646 0 net=1961
rlabel metal2 282 -1646 282 -1646 0 net=1927
rlabel metal2 352 -1646 352 -1646 0 net=2045
rlabel metal2 429 -1646 429 -1646 0 net=2655
rlabel metal2 464 -1646 464 -1646 0 net=1910
rlabel metal2 65 -1648 65 -1648 0 net=3601
rlabel metal2 401 -1648 401 -1648 0 net=3633
rlabel metal2 464 -1648 464 -1648 0 net=4133
rlabel metal2 65 -1650 65 -1650 0 net=1623
rlabel metal2 128 -1650 128 -1650 0 net=3657
rlabel metal2 282 -1650 282 -1650 0 net=2567
rlabel metal2 450 -1650 450 -1650 0 net=5107
rlabel metal2 135 -1652 135 -1652 0 net=1090
rlabel metal2 317 -1652 317 -1652 0 net=2219
rlabel metal2 401 -1652 401 -1652 0 net=4813
rlabel metal2 135 -1654 135 -1654 0 net=2659
rlabel metal2 163 -1654 163 -1654 0 net=1591
rlabel metal2 219 -1654 219 -1654 0 net=3119
rlabel metal2 331 -1654 331 -1654 0 net=4125
rlabel metal2 72 -1656 72 -1656 0 net=1597
rlabel metal2 408 -1656 408 -1656 0 net=2253
rlabel metal2 453 -1656 453 -1656 0 net=4996
rlabel metal2 145 -1658 145 -1658 0 net=2421
rlabel metal2 471 -1658 471 -1658 0 net=4035
rlabel metal2 149 -1660 149 -1660 0 net=5044
rlabel metal2 166 -1662 166 -1662 0 net=2820
rlabel metal2 471 -1662 471 -1662 0 net=3187
rlabel metal2 527 -1662 527 -1662 0 net=4876
rlabel metal2 170 -1664 170 -1664 0 net=3838
rlabel metal2 198 -1664 198 -1664 0 net=1353
rlabel metal2 478 -1664 478 -1664 0 net=2827
rlabel metal2 495 -1664 495 -1664 0 net=4872
rlabel metal2 173 -1666 173 -1666 0 net=2325
rlabel metal2 254 -1666 254 -1666 0 net=3063
rlabel metal2 527 -1666 527 -1666 0 net=3109
rlabel metal2 555 -1666 555 -1666 0 net=4179
rlabel metal2 173 -1668 173 -1668 0 net=2067
rlabel metal2 198 -1668 198 -1668 0 net=2843
rlabel metal2 254 -1668 254 -1668 0 net=1383
rlabel metal2 268 -1668 268 -1668 0 net=1347
rlabel metal2 488 -1668 488 -1668 0 net=3570
rlabel metal2 79 -1670 79 -1670 0 net=1729
rlabel metal2 261 -1670 261 -1670 0 net=1417
rlabel metal2 492 -1670 492 -1670 0 net=3231
rlabel metal2 506 -1670 506 -1670 0 net=3211
rlabel metal2 555 -1670 555 -1670 0 net=3319
rlabel metal2 586 -1670 586 -1670 0 net=4307
rlabel metal2 233 -1672 233 -1672 0 net=2635
rlabel metal2 499 -1672 499 -1672 0 net=3261
rlabel metal2 534 -1672 534 -1672 0 net=5254
rlabel metal2 156 -1674 156 -1674 0 net=2809
rlabel metal2 537 -1674 537 -1674 0 net=5185
rlabel metal2 142 -1676 142 -1676 0 net=1609
rlabel metal2 509 -1676 509 -1676 0 net=3422
rlabel metal2 142 -1678 142 -1678 0 net=3355
rlabel metal2 590 -1678 590 -1678 0 net=4761
rlabel metal2 786 -1678 786 -1678 0 net=5171
rlabel metal2 814 -1678 814 -1678 0 net=5389
rlabel metal2 485 -1680 485 -1680 0 net=2867
rlabel metal2 541 -1682 541 -1682 0 net=3515
rlabel metal2 520 -1684 520 -1684 0 net=3343
rlabel metal2 544 -1684 544 -1684 0 net=4384
rlabel metal2 562 -1686 562 -1686 0 net=4284
rlabel metal2 611 -1686 611 -1686 0 net=3981
rlabel metal2 152 -1688 152 -1688 0 net=3505
rlabel metal2 443 -1690 443 -1690 0 net=3487
rlabel metal2 436 -1692 436 -1692 0 net=2597
rlabel metal2 481 -1692 481 -1692 0 net=4777
rlabel metal2 565 -1692 565 -1692 0 net=4981
rlabel metal2 380 -1694 380 -1694 0 net=2071
rlabel metal2 569 -1694 569 -1694 0 net=3577
rlabel metal2 569 -1696 569 -1696 0 net=4213
rlabel metal2 583 -1698 583 -1698 0 net=3897
rlabel metal2 572 -1700 572 -1700 0 net=5301
rlabel metal2 590 -1700 590 -1700 0 net=3387
rlabel metal2 597 -1702 597 -1702 0 net=4745
rlabel metal2 394 -1704 394 -1704 0 net=3459
rlabel metal2 16 -1715 16 -1715 0 net=593
rlabel metal2 72 -1715 72 -1715 0 net=1093
rlabel metal2 79 -1715 79 -1715 0 net=1730
rlabel metal2 506 -1715 506 -1715 0 net=3212
rlabel metal2 572 -1715 572 -1715 0 net=3730
rlabel metal2 905 -1715 905 -1715 0 net=4988
rlabel metal2 926 -1715 926 -1715 0 net=4776
rlabel metal2 961 -1715 961 -1715 0 net=3334
rlabel metal2 16 -1717 16 -1717 0 net=2221
rlabel metal2 355 -1717 355 -1717 0 net=4814
rlabel metal2 37 -1719 37 -1719 0 net=4086
rlabel metal2 397 -1719 397 -1719 0 net=2656
rlabel metal2 436 -1719 436 -1719 0 net=4215
rlabel metal2 709 -1719 709 -1719 0 net=4763
rlabel metal2 37 -1721 37 -1721 0 net=121
rlabel metal2 523 -1721 523 -1721 0 net=4126
rlabel metal2 51 -1723 51 -1723 0 net=1260
rlabel metal2 376 -1723 376 -1723 0 net=4182
rlabel metal2 58 -1725 58 -1725 0 net=1625
rlabel metal2 93 -1725 93 -1725 0 net=1576
rlabel metal2 439 -1725 439 -1725 0 net=2868
rlabel metal2 9 -1727 9 -1727 0 net=3079
rlabel metal2 103 -1727 103 -1727 0 net=3634
rlabel metal2 467 -1727 467 -1727 0 net=3516
rlabel metal2 9 -1729 9 -1729 0 net=144
rlabel metal2 387 -1729 387 -1729 0 net=2255
rlabel metal2 450 -1729 450 -1729 0 net=3578
rlabel metal2 86 -1731 86 -1731 0 net=2088
rlabel metal2 117 -1731 117 -1731 0 net=2810
rlabel metal2 548 -1731 548 -1731 0 net=3321
rlabel metal2 642 -1731 642 -1731 0 net=5390
rlabel metal2 23 -1733 23 -1733 0 net=2396
rlabel metal2 121 -1733 121 -1733 0 net=1993
rlabel metal2 159 -1733 159 -1733 0 net=4576
rlabel metal2 23 -1735 23 -1735 0 net=3269
rlabel metal2 191 -1735 191 -1735 0 net=1599
rlabel metal2 222 -1735 222 -1735 0 net=563
rlabel metal2 450 -1735 450 -1735 0 net=2829
rlabel metal2 485 -1735 485 -1735 0 net=3232
rlabel metal2 534 -1735 534 -1735 0 net=3389
rlabel metal2 667 -1735 667 -1735 0 net=5323
rlabel metal2 82 -1737 82 -1737 0 net=361
rlabel metal2 124 -1737 124 -1737 0 net=3641
rlabel metal2 702 -1737 702 -1737 0 net=4897
rlabel metal2 128 -1739 128 -1739 0 net=3659
rlabel metal2 730 -1739 730 -1739 0 net=5173
rlabel metal2 142 -1741 142 -1741 0 net=1479
rlabel metal2 737 -1741 737 -1741 0 net=5187
rlabel metal2 163 -1743 163 -1743 0 net=1592
rlabel metal2 173 -1743 173 -1743 0 net=1418
rlabel metal2 268 -1743 268 -1743 0 net=1348
rlabel metal2 471 -1743 471 -1743 0 net=3189
rlabel metal2 488 -1743 488 -1743 0 net=4601
rlabel metal2 166 -1745 166 -1745 0 net=2422
rlabel metal2 474 -1745 474 -1745 0 net=4180
rlabel metal2 170 -1747 170 -1747 0 net=4769
rlabel metal2 422 -1747 422 -1747 0 net=1969
rlabel metal2 191 -1749 191 -1749 0 net=2337
rlabel metal2 261 -1749 261 -1749 0 net=1293
rlabel metal2 310 -1749 310 -1749 0 net=1556
rlabel metal2 478 -1749 478 -1749 0 net=3111
rlabel metal2 555 -1749 555 -1749 0 net=3507
rlabel metal2 660 -1749 660 -1749 0 net=4531
rlabel metal2 107 -1751 107 -1751 0 net=1709
rlabel metal2 324 -1751 324 -1751 0 net=1929
rlabel metal2 527 -1751 527 -1751 0 net=3357
rlabel metal2 716 -1751 716 -1751 0 net=5223
rlabel metal2 107 -1753 107 -1753 0 net=2661
rlabel metal2 156 -1753 156 -1753 0 net=1611
rlabel metal2 271 -1753 271 -1753 0 net=5342
rlabel metal2 30 -1755 30 -1755 0 net=1956
rlabel metal2 219 -1755 219 -1755 0 net=2327
rlabel metal2 324 -1755 324 -1755 0 net=2725
rlabel metal2 576 -1755 576 -1755 0 net=3851
rlabel metal2 723 -1755 723 -1755 0 net=5109
rlabel metal2 30 -1757 30 -1757 0 net=2569
rlabel metal2 219 -1757 219 -1757 0 net=2957
rlabel metal2 625 -1757 625 -1757 0 net=4309
rlabel metal2 226 -1759 226 -1759 0 net=1656
rlabel metal2 695 -1759 695 -1759 0 net=4553
rlabel metal2 114 -1761 114 -1761 0 net=1815
rlabel metal2 233 -1761 233 -1761 0 net=1354
rlabel metal2 541 -1761 541 -1761 0 net=3461
rlabel metal2 639 -1761 639 -1761 0 net=4983
rlabel metal2 198 -1763 198 -1763 0 net=2845
rlabel metal2 236 -1763 236 -1763 0 net=4041
rlabel metal2 198 -1765 198 -1765 0 net=2533
rlabel metal2 338 -1765 338 -1765 0 net=2047
rlabel metal2 415 -1765 415 -1765 0 net=3345
rlabel metal2 597 -1765 597 -1765 0 net=3899
rlabel metal2 240 -1767 240 -1767 0 net=1814
rlabel metal2 443 -1767 443 -1767 0 net=2599
rlabel metal2 44 -1769 44 -1769 0 net=2947
rlabel metal2 44 -1771 44 -1771 0 net=3263
rlabel metal2 240 -1773 240 -1773 0 net=1215
rlabel metal2 499 -1773 499 -1773 0 net=4036
rlabel metal2 254 -1775 254 -1775 0 net=1384
rlabel metal2 653 -1775 653 -1775 0 net=4747
rlabel metal2 184 -1777 184 -1777 0 net=2069
rlabel metal2 275 -1777 275 -1777 0 net=2637
rlabel metal2 184 -1779 184 -1779 0 net=2968
rlabel metal2 583 -1779 583 -1779 0 net=5303
rlabel metal2 212 -1781 212 -1781 0 net=1963
rlabel metal2 282 -1781 282 -1781 0 net=2568
rlabel metal2 583 -1781 583 -1781 0 net=3781
rlabel metal2 93 -1783 93 -1783 0 net=1109
rlabel metal2 282 -1783 282 -1783 0 net=1153
rlabel metal2 464 -1783 464 -1783 0 net=3065
rlabel metal2 618 -1783 618 -1783 0 net=4135
rlabel metal2 289 -1785 289 -1785 0 net=3055
rlabel metal2 562 -1785 562 -1785 0 net=4779
rlabel metal2 180 -1787 180 -1787 0 net=1145
rlabel metal2 296 -1787 296 -1787 0 net=33
rlabel metal2 352 -1787 352 -1787 0 net=3603
rlabel metal2 296 -1789 296 -1789 0 net=2073
rlabel metal2 401 -1789 401 -1789 0 net=4341
rlabel metal2 299 -1791 299 -1791 0 net=115
rlabel metal2 317 -1793 317 -1793 0 net=3121
rlabel metal2 359 -1793 359 -1793 0 net=3489
rlabel metal2 604 -1795 604 -1795 0 net=3983
rlabel metal2 632 -1797 632 -1797 0 net=4939
rlabel metal2 352 -1799 352 -1799 0 net=4285
rlabel metal2 9 -1810 9 -1810 0 net=2570
rlabel metal2 33 -1810 33 -1810 0 net=1905
rlabel metal2 40 -1810 40 -1810 0 net=122
rlabel metal2 89 -1810 89 -1810 0 net=1970
rlabel metal2 457 -1810 457 -1810 0 net=3057
rlabel metal2 457 -1810 457 -1810 0 net=3057
rlabel metal2 471 -1810 471 -1810 0 net=3113
rlabel metal2 492 -1810 492 -1810 0 net=5324
rlabel metal2 23 -1812 23 -1812 0 net=3271
rlabel metal2 93 -1812 93 -1812 0 net=1111
rlabel metal2 219 -1812 219 -1812 0 net=1964
rlabel metal2 306 -1812 306 -1812 0 net=2048
rlabel metal2 345 -1812 345 -1812 0 net=1930
rlabel metal2 366 -1812 366 -1812 0 net=2677
rlabel metal2 380 -1812 380 -1812 0 net=3508
rlabel metal2 579 -1812 579 -1812 0 net=5188
rlabel metal2 744 -1812 744 -1812 0 net=4984
rlabel metal2 744 -1812 744 -1812 0 net=4984
rlabel metal2 44 -1814 44 -1814 0 net=3265
rlabel metal2 492 -1814 492 -1814 0 net=3277
rlabel metal2 506 -1814 506 -1814 0 net=3984
rlabel metal2 667 -1814 667 -1814 0 net=4603
rlabel metal2 667 -1814 667 -1814 0 net=4603
rlabel metal2 674 -1814 674 -1814 0 net=4941
rlabel metal2 723 -1814 723 -1814 0 net=5111
rlabel metal2 723 -1814 723 -1814 0 net=5111
rlabel metal2 737 -1814 737 -1814 0 net=5305
rlabel metal2 51 -1816 51 -1816 0 net=2663
rlabel metal2 121 -1816 121 -1816 0 net=3122
rlabel metal2 348 -1816 348 -1816 0 net=2638
rlabel metal2 58 -1818 58 -1818 0 net=1627
rlabel metal2 58 -1818 58 -1818 0 net=1627
rlabel metal2 65 -1818 65 -1818 0 net=3080
rlabel metal2 219 -1818 219 -1818 0 net=1155
rlabel metal2 331 -1818 331 -1818 0 net=3067
rlabel metal2 495 -1818 495 -1818 0 net=4163
rlabel metal2 65 -1820 65 -1820 0 net=2847
rlabel metal2 240 -1820 240 -1820 0 net=1216
rlabel metal2 513 -1820 513 -1820 0 net=3359
rlabel metal2 604 -1820 604 -1820 0 net=4043
rlabel metal2 653 -1820 653 -1820 0 net=4749
rlabel metal2 72 -1822 72 -1822 0 net=1094
rlabel metal2 240 -1822 240 -1822 0 net=2075
rlabel metal2 352 -1822 352 -1822 0 net=2811
rlabel metal2 464 -1822 464 -1822 0 net=3390
rlabel metal2 611 -1822 611 -1822 0 net=4137
rlabel metal2 674 -1822 674 -1822 0 net=4781
rlabel metal2 72 -1824 72 -1824 0 net=1481
rlabel metal2 149 -1824 149 -1824 0 net=1995
rlabel metal2 184 -1824 184 -1824 0 net=2339
rlabel metal2 201 -1824 201 -1824 0 net=21
rlabel metal2 415 -1824 415 -1824 0 net=3347
rlabel metal2 516 -1824 516 -1824 0 net=5174
rlabel metal2 47 -1826 47 -1826 0 net=2791
rlabel metal2 453 -1826 453 -1826 0 net=3761
rlabel metal2 618 -1826 618 -1826 0 net=4287
rlabel metal2 681 -1826 681 -1826 0 net=4765
rlabel metal2 79 -1828 79 -1828 0 net=2465
rlabel metal2 121 -1828 121 -1828 0 net=1241
rlabel metal2 268 -1828 268 -1828 0 net=3660
rlabel metal2 695 -1828 695 -1828 0 net=4555
rlabel metal2 93 -1830 93 -1830 0 net=2315
rlabel metal2 509 -1830 509 -1830 0 net=4587
rlabel metal2 695 -1830 695 -1830 0 net=5225
rlabel metal2 103 -1832 103 -1832 0 net=1146
rlabel metal2 296 -1832 296 -1832 0 net=1711
rlabel metal2 338 -1832 338 -1832 0 net=5217
rlabel metal2 107 -1834 107 -1834 0 net=2535
rlabel metal2 275 -1834 275 -1834 0 net=2949
rlabel metal2 520 -1834 520 -1834 0 net=3323
rlabel metal2 590 -1834 590 -1834 0 net=4311
rlabel metal2 100 -1836 100 -1836 0 net=3125
rlabel metal2 282 -1836 282 -1836 0 net=3191
rlabel metal2 625 -1836 625 -1836 0 net=4533
rlabel metal2 124 -1838 124 -1838 0 net=3431
rlabel metal2 642 -1838 642 -1838 0 net=3865
rlabel metal2 128 -1840 128 -1840 0 net=1612
rlabel metal2 352 -1840 352 -1840 0 net=4089
rlabel metal2 135 -1842 135 -1842 0 net=4216
rlabel metal2 443 -1842 443 -1842 0 net=3462
rlabel metal2 142 -1844 142 -1844 0 net=2070
rlabel metal2 355 -1844 355 -1844 0 net=3642
rlabel metal2 156 -1846 156 -1846 0 net=1601
rlabel metal2 247 -1846 247 -1846 0 net=1295
rlabel metal2 310 -1846 310 -1846 0 net=2329
rlabel metal2 16 -1848 16 -1848 0 net=2223
rlabel metal2 254 -1848 254 -1848 0 net=1767
rlabel metal2 369 -1848 369 -1848 0 net=3900
rlabel metal2 16 -1850 16 -1850 0 net=2289
rlabel metal2 310 -1850 310 -1850 0 net=2727
rlabel metal2 359 -1850 359 -1850 0 net=3491
rlabel metal2 387 -1850 387 -1850 0 net=2257
rlabel metal2 450 -1850 450 -1850 0 net=2831
rlabel metal2 163 -1852 163 -1852 0 net=3604
rlabel metal2 12 -1854 12 -1854 0 net=3803
rlabel metal2 131 -1856 131 -1856 0 net=921
rlabel metal2 166 -1856 166 -1856 0 net=3715
rlabel metal2 170 -1858 170 -1858 0 net=1377
rlabel metal2 261 -1858 261 -1858 0 net=4343
rlabel metal2 485 -1858 485 -1858 0 net=3159
rlabel metal2 135 -1860 135 -1860 0 net=1275
rlabel metal2 173 -1860 173 -1860 0 net=3815
rlabel metal2 187 -1862 187 -1862 0 net=1816
rlabel metal2 268 -1862 268 -1862 0 net=1055
rlabel metal2 114 -1864 114 -1864 0 net=1171
rlabel metal2 324 -1864 324 -1864 0 net=3767
rlabel metal2 373 -1866 373 -1866 0 net=4898
rlabel metal2 303 -1868 303 -1868 0 net=214
rlabel metal2 387 -1868 387 -1868 0 net=3782
rlabel metal2 390 -1870 390 -1870 0 net=2600
rlabel metal2 180 -1872 180 -1872 0 net=4271
rlabel metal2 408 -1874 408 -1874 0 net=4771
rlabel metal2 408 -1876 408 -1876 0 net=2959
rlabel metal2 576 -1876 576 -1876 0 net=3853
rlabel metal2 317 -1878 317 -1878 0 net=4015
rlabel metal2 138 -1880 138 -1880 0 net=3771
rlabel metal2 2 -1891 2 -1891 0 net=1483
rlabel metal2 107 -1891 107 -1891 0 net=2536
rlabel metal2 177 -1891 177 -1891 0 net=1997
rlabel metal2 194 -1891 194 -1891 0 net=2792
rlabel metal2 432 -1891 432 -1891 0 net=5306
rlabel metal2 5 -1893 5 -1893 0 net=9
rlabel metal2 201 -1893 201 -1893 0 net=630
rlabel metal2 376 -1893 376 -1893 0 net=4272
rlabel metal2 709 -1893 709 -1893 0 net=4556
rlabel metal2 9 -1895 9 -1895 0 net=2695
rlabel metal2 397 -1895 397 -1895 0 net=3716
rlabel metal2 583 -1895 583 -1895 0 net=3855
rlabel metal2 583 -1895 583 -1895 0 net=3855
rlabel metal2 604 -1895 604 -1895 0 net=4045
rlabel metal2 604 -1895 604 -1895 0 net=4045
rlabel metal2 611 -1895 611 -1895 0 net=4139
rlabel metal2 611 -1895 611 -1895 0 net=4139
rlabel metal2 12 -1897 12 -1897 0 net=933
rlabel metal2 177 -1897 177 -1897 0 net=1435
rlabel metal2 240 -1897 240 -1897 0 net=2076
rlabel metal2 338 -1897 338 -1897 0 net=3763
rlabel metal2 541 -1897 541 -1897 0 net=3769
rlabel metal2 23 -1899 23 -1899 0 net=1378
rlabel metal2 292 -1899 292 -1899 0 net=2330
rlabel metal2 23 -1901 23 -1901 0 net=2349
rlabel metal2 471 -1901 471 -1901 0 net=3114
rlabel metal2 562 -1901 562 -1901 0 net=3805
rlabel metal2 33 -1903 33 -1903 0 net=1906
rlabel metal2 44 -1903 44 -1903 0 net=1057
rlabel metal2 296 -1903 296 -1903 0 net=1712
rlabel metal2 317 -1903 317 -1903 0 net=3772
rlabel metal2 436 -1903 436 -1903 0 net=2832
rlabel metal2 26 -1905 26 -1905 0 net=786
rlabel metal2 296 -1905 296 -1905 0 net=1603
rlabel metal2 345 -1905 345 -1905 0 net=4772
rlabel metal2 51 -1907 51 -1907 0 net=2664
rlabel metal2 156 -1907 156 -1907 0 net=1602
rlabel metal2 324 -1907 324 -1907 0 net=3349
rlabel metal2 520 -1907 520 -1907 0 net=3325
rlabel metal2 541 -1907 541 -1907 0 net=4313
rlabel metal2 597 -1907 597 -1907 0 net=4589
rlabel metal2 674 -1907 674 -1907 0 net=4783
rlabel metal2 51 -1909 51 -1909 0 net=1628
rlabel metal2 61 -1909 61 -1909 0 net=2466
rlabel metal2 117 -1909 117 -1909 0 net=549
rlabel metal2 184 -1909 184 -1909 0 net=2340
rlabel metal2 254 -1909 254 -1909 0 net=1769
rlabel metal2 359 -1909 359 -1909 0 net=3777
rlabel metal2 590 -1909 590 -1909 0 net=3867
rlabel metal2 667 -1909 667 -1909 0 net=4605
rlabel metal2 65 -1911 65 -1911 0 net=2848
rlabel metal2 184 -1911 184 -1911 0 net=1157
rlabel metal2 303 -1911 303 -1911 0 net=1635
rlabel metal2 471 -1911 471 -1911 0 net=3587
rlabel metal2 502 -1911 502 -1911 0 net=5112
rlabel metal2 65 -1913 65 -1913 0 net=3193
rlabel metal2 331 -1913 331 -1913 0 net=3069
rlabel metal2 362 -1913 362 -1913 0 net=2678
rlabel metal2 380 -1913 380 -1913 0 net=3493
rlabel metal2 625 -1913 625 -1913 0 net=4535
rlabel metal2 16 -1915 16 -1915 0 net=2291
rlabel metal2 366 -1915 366 -1915 0 net=4447
rlabel metal2 72 -1917 72 -1917 0 net=573
rlabel metal2 618 -1917 618 -1917 0 net=4289
rlabel metal2 639 -1917 639 -1917 0 net=5347
rlabel metal2 79 -1919 79 -1919 0 net=3413
rlabel metal2 506 -1919 506 -1919 0 net=3433
rlabel metal2 618 -1919 618 -1919 0 net=4165
rlabel metal2 19 -1921 19 -1921 0 net=3563
rlabel metal2 114 -1923 114 -1923 0 net=1173
rlabel metal2 261 -1923 261 -1923 0 net=4345
rlabel metal2 380 -1923 380 -1923 0 net=2259
rlabel metal2 401 -1923 401 -1923 0 net=3817
rlabel metal2 100 -1925 100 -1925 0 net=3127
rlabel metal2 355 -1925 355 -1925 0 net=209
rlabel metal2 401 -1925 401 -1925 0 net=2813
rlabel metal2 429 -1925 429 -1925 0 net=4017
rlabel metal2 100 -1927 100 -1927 0 net=3663
rlabel metal2 121 -1929 121 -1929 0 net=1243
rlabel metal2 121 -1929 121 -1929 0 net=1243
rlabel metal2 128 -1929 128 -1929 0 net=2729
rlabel metal2 429 -1929 429 -1929 0 net=838
rlabel metal2 131 -1931 131 -1931 0 net=4090
rlabel metal2 145 -1933 145 -1933 0 net=2377
rlabel metal2 436 -1933 436 -1933 0 net=3161
rlabel metal2 205 -1935 205 -1935 0 net=2225
rlabel metal2 310 -1935 310 -1935 0 net=3058
rlabel metal2 485 -1935 485 -1935 0 net=3361
rlabel metal2 149 -1937 149 -1937 0 net=1761
rlabel metal2 208 -1937 208 -1937 0 net=5218
rlabel metal2 142 -1939 142 -1939 0 net=5445
rlabel metal2 86 -1941 86 -1941 0 net=3273
rlabel metal2 212 -1941 212 -1941 0 net=1113
rlabel metal2 271 -1941 271 -1941 0 net=4451
rlabel metal2 86 -1943 86 -1943 0 net=1277
rlabel metal2 163 -1943 163 -1943 0 net=1103
rlabel metal2 219 -1943 219 -1943 0 net=1837
rlabel metal2 352 -1943 352 -1943 0 net=3475
rlabel metal2 135 -1945 135 -1945 0 net=2961
rlabel metal2 439 -1945 439 -1945 0 net=4955
rlabel metal2 275 -1947 275 -1947 0 net=2951
rlabel metal2 443 -1947 443 -1947 0 net=3279
rlabel metal2 247 -1949 247 -1949 0 net=1297
rlabel metal2 422 -1949 422 -1949 0 net=3379
rlabel metal2 93 -1951 93 -1951 0 net=2317
rlabel metal2 450 -1951 450 -1951 0 net=4750
rlabel metal2 37 -1953 37 -1953 0 net=4735
rlabel metal2 93 -1955 93 -1955 0 net=2389
rlabel metal2 450 -1955 450 -1955 0 net=3267
rlabel metal2 478 -1957 478 -1957 0 net=4942
rlabel metal2 695 -1959 695 -1959 0 net=5227
rlabel metal2 681 -1961 681 -1961 0 net=4767
rlabel metal2 54 -1963 54 -1963 0 net=4649
rlabel metal2 16 -1974 16 -1974 0 net=3275
rlabel metal2 156 -1974 156 -1974 0 net=3128
rlabel metal2 285 -1974 285 -1974 0 net=3664
rlabel metal2 635 -1974 635 -1974 0 net=5228
rlabel metal2 19 -1976 19 -1976 0 net=4346
rlabel metal2 366 -1976 366 -1976 0 net=3868
rlabel metal2 642 -1976 642 -1976 0 net=4768
rlabel metal2 23 -1978 23 -1978 0 net=2351
rlabel metal2 240 -1978 240 -1978 0 net=1114
rlabel metal2 324 -1978 324 -1978 0 net=3350
rlabel metal2 450 -1978 450 -1978 0 net=3268
rlabel metal2 534 -1978 534 -1978 0 net=3326
rlabel metal2 551 -1978 551 -1978 0 net=4536
rlabel metal2 695 -1978 695 -1978 0 net=5349
rlabel metal2 23 -1980 23 -1980 0 net=596
rlabel metal2 37 -1980 37 -1980 0 net=1579
rlabel metal2 100 -1980 100 -1980 0 net=3070
rlabel metal2 366 -1980 366 -1980 0 net=3047
rlabel metal2 562 -1980 562 -1980 0 net=3778
rlabel metal2 30 -1982 30 -1982 0 net=2375
rlabel metal2 110 -1982 110 -1982 0 net=710
rlabel metal2 163 -1982 163 -1982 0 net=1105
rlabel metal2 331 -1982 331 -1982 0 net=3813
rlabel metal2 404 -1982 404 -1982 0 net=3588
rlabel metal2 478 -1982 478 -1982 0 net=3901
rlabel metal2 44 -1984 44 -1984 0 net=1058
rlabel metal2 443 -1984 443 -1984 0 net=3281
rlabel metal2 457 -1984 457 -1984 0 net=3856
rlabel metal2 618 -1984 618 -1984 0 net=4167
rlabel metal2 44 -1986 44 -1986 0 net=1279
rlabel metal2 93 -1986 93 -1986 0 net=2391
rlabel metal2 170 -1986 170 -1986 0 net=1604
rlabel metal2 303 -1986 303 -1986 0 net=1637
rlabel metal2 369 -1986 369 -1986 0 net=4018
rlabel metal2 51 -1988 51 -1988 0 net=4736
rlabel metal2 58 -1990 58 -1990 0 net=2059
rlabel metal2 107 -1990 107 -1990 0 net=2962
rlabel metal2 142 -1990 142 -1990 0 net=3625
rlabel metal2 219 -1990 219 -1990 0 net=3041
rlabel metal2 387 -1990 387 -1990 0 net=3806
rlabel metal2 583 -1990 583 -1990 0 net=4449
rlabel metal2 65 -1992 65 -1992 0 net=3195
rlabel metal2 100 -1992 100 -1992 0 net=4956
rlabel metal2 2 -1994 2 -1994 0 net=1484
rlabel metal2 68 -1994 68 -1994 0 net=4201
rlabel metal2 177 -1994 177 -1994 0 net=482
rlabel metal2 215 -1994 215 -1994 0 net=217
rlabel metal2 72 -1996 72 -1996 0 net=1301
rlabel metal2 117 -1996 117 -1996 0 net=3414
rlabel metal2 534 -1996 534 -1996 0 net=4651
rlabel metal2 117 -1998 117 -1998 0 net=4273
rlabel metal2 149 -1998 149 -1998 0 net=1763
rlabel metal2 177 -1998 177 -1998 0 net=1159
rlabel metal2 191 -1998 191 -1998 0 net=1999
rlabel metal2 254 -1998 254 -1998 0 net=1174
rlabel metal2 289 -1998 289 -1998 0 net=2227
rlabel metal2 387 -1998 387 -1998 0 net=2953
rlabel metal2 415 -1998 415 -1998 0 net=5141
rlabel metal2 604 -1998 604 -1998 0 net=4047
rlabel metal2 9 -2000 9 -2000 0 net=2697
rlabel metal2 184 -2000 184 -2000 0 net=3770
rlabel metal2 562 -2000 562 -2000 0 net=4591
rlabel metal2 604 -2000 604 -2000 0 net=4607
rlabel metal2 9 -2002 9 -2002 0 net=4961
rlabel metal2 219 -2002 219 -2002 0 net=1838
rlabel metal2 247 -2002 247 -2002 0 net=2319
rlabel metal2 289 -2002 289 -2002 0 net=3765
rlabel metal2 380 -2002 380 -2002 0 net=2260
rlabel metal2 418 -2002 418 -2002 0 net=3434
rlabel metal2 569 -2002 569 -2002 0 net=4453
rlabel metal2 54 -2004 54 -2004 0 net=4257
rlabel metal2 394 -2004 394 -2004 0 net=2815
rlabel metal2 408 -2004 408 -2004 0 net=3163
rlabel metal2 443 -2004 443 -2004 0 net=3477
rlabel metal2 597 -2004 597 -2004 0 net=5447
rlabel metal2 54 -2006 54 -2006 0 net=4963
rlabel metal2 506 -2006 506 -2006 0 net=3819
rlabel metal2 642 -2006 642 -2006 0 net=346
rlabel metal2 121 -2008 121 -2008 0 net=1244
rlabel metal2 226 -2008 226 -2008 0 net=1436
rlabel metal2 261 -2008 261 -2008 0 net=1299
rlabel metal2 422 -2008 422 -2008 0 net=2893
rlabel metal2 513 -2008 513 -2008 0 net=4315
rlabel metal2 576 -2008 576 -2008 0 net=4291
rlabel metal2 128 -2010 128 -2010 0 net=2731
rlabel metal2 457 -2010 457 -2010 0 net=3363
rlabel metal2 541 -2010 541 -2010 0 net=4141
rlabel metal2 625 -2010 625 -2010 0 net=5449
rlabel metal2 121 -2012 121 -2012 0 net=2467
rlabel metal2 131 -2012 131 -2012 0 net=182
rlabel metal2 464 -2012 464 -2012 0 net=3494
rlabel metal2 611 -2012 611 -2012 0 net=4785
rlabel metal2 226 -2014 226 -2014 0 net=2379
rlabel metal2 474 -2014 474 -2014 0 net=4641
rlabel metal2 233 -2016 233 -2016 0 net=1561
rlabel metal2 373 -2016 373 -2016 0 net=2767
rlabel metal2 492 -2016 492 -2016 0 net=3380
rlabel metal2 275 -2018 275 -2018 0 net=1771
rlabel metal2 429 -2018 429 -2018 0 net=3565
rlabel metal2 282 -2020 282 -2020 0 net=2293
rlabel metal2 348 -2020 348 -2020 0 net=4653
rlabel metal2 282 -2022 282 -2022 0 net=4323
rlabel metal2 303 -2024 303 -2024 0 net=2877
rlabel metal2 436 -2024 436 -2024 0 net=4361
rlabel metal2 9 -2035 9 -2035 0 net=4962
rlabel metal2 212 -2035 212 -2035 0 net=3566
rlabel metal2 436 -2035 436 -2035 0 net=5450
rlabel metal2 632 -2035 632 -2035 0 net=410
rlabel metal2 646 -2035 646 -2035 0 net=4169
rlabel metal2 688 -2035 688 -2035 0 net=5351
rlabel metal2 16 -2037 16 -2037 0 net=3276
rlabel metal2 114 -2037 114 -2037 0 net=3766
rlabel metal2 296 -2037 296 -2037 0 net=3043
rlabel metal2 296 -2037 296 -2037 0 net=3043
rlabel metal2 303 -2037 303 -2037 0 net=2228
rlabel metal2 380 -2037 380 -2037 0 net=3478
rlabel metal2 474 -2037 474 -2037 0 net=4316
rlabel metal2 520 -2037 520 -2037 0 net=4143
rlabel metal2 548 -2037 548 -2037 0 net=4450
rlabel metal2 16 -2039 16 -2039 0 net=4509
rlabel metal2 177 -2039 177 -2039 0 net=1161
rlabel metal2 177 -2039 177 -2039 0 net=1161
rlabel metal2 191 -2039 191 -2039 0 net=2954
rlabel metal2 415 -2039 415 -2039 0 net=4652
rlabel metal2 541 -2039 541 -2039 0 net=4593
rlabel metal2 30 -2041 30 -2041 0 net=2376
rlabel metal2 121 -2041 121 -2041 0 net=2469
rlabel metal2 121 -2041 121 -2041 0 net=2469
rlabel metal2 128 -2041 128 -2041 0 net=4275
rlabel metal2 191 -2041 191 -2041 0 net=2000
rlabel metal2 257 -2041 257 -2041 0 net=1300
rlabel metal2 289 -2041 289 -2041 0 net=1069
rlabel metal2 481 -2041 481 -2041 0 net=4454
rlabel metal2 37 -2043 37 -2043 0 net=1580
rlabel metal2 303 -2043 303 -2043 0 net=3201
rlabel metal2 443 -2043 443 -2043 0 net=3283
rlabel metal2 471 -2043 471 -2043 0 net=3821
rlabel metal2 548 -2043 548 -2043 0 net=4293
rlabel metal2 33 -2045 33 -2045 0 net=1731
rlabel metal2 44 -2045 44 -2045 0 net=1280
rlabel metal2 100 -2045 100 -2045 0 net=1177
rlabel metal2 117 -2045 117 -2045 0 net=475
rlabel metal2 198 -2045 198 -2045 0 net=589
rlabel metal2 425 -2045 425 -2045 0 net=5448
rlabel metal2 44 -2047 44 -2047 0 net=3627
rlabel metal2 194 -2047 194 -2047 0 net=2341
rlabel metal2 205 -2047 205 -2047 0 net=2353
rlabel metal2 313 -2047 313 -2047 0 net=5353
rlabel metal2 51 -2049 51 -2049 0 net=1302
rlabel metal2 79 -2049 79 -2049 0 net=3196
rlabel metal2 429 -2049 429 -2049 0 net=3903
rlabel metal2 485 -2049 485 -2049 0 net=4243
rlabel metal2 51 -2051 51 -2051 0 net=4037
rlabel metal2 212 -2051 212 -2051 0 net=1639
rlabel metal2 320 -2051 320 -2051 0 net=4643
rlabel metal2 555 -2051 555 -2051 0 net=4642
rlabel metal2 65 -2053 65 -2053 0 net=4964
rlabel metal2 555 -2053 555 -2053 0 net=4048
rlabel metal2 642 -2053 642 -2053 0 net=473
rlabel metal2 65 -2055 65 -2055 0 net=1765
rlabel metal2 215 -2055 215 -2055 0 net=91
rlabel metal2 75 -2057 75 -2057 0 net=1747
rlabel metal2 86 -2057 86 -2057 0 net=3071
rlabel metal2 170 -2057 170 -2057 0 net=1773
rlabel metal2 327 -2057 327 -2057 0 net=2878
rlabel metal2 359 -2057 359 -2057 0 net=2733
rlabel metal2 418 -2057 418 -2057 0 net=5163
rlabel metal2 107 -2059 107 -2059 0 net=2393
rlabel metal2 219 -2059 219 -2059 0 net=4654
rlabel metal2 562 -2059 562 -2059 0 net=4787
rlabel metal2 58 -2061 58 -2061 0 net=2060
rlabel metal2 222 -2061 222 -2061 0 net=2380
rlabel metal2 236 -2061 236 -2061 0 net=4907
rlabel metal2 604 -2061 604 -2061 0 net=4609
rlabel metal2 58 -2063 58 -2063 0 net=998
rlabel metal2 149 -2063 149 -2063 0 net=2699
rlabel metal2 383 -2063 383 -2063 0 net=3164
rlabel metal2 450 -2063 450 -2063 0 net=3365
rlabel metal2 492 -2063 492 -2063 0 net=4363
rlabel metal2 149 -2065 149 -2065 0 net=1563
rlabel metal2 240 -2065 240 -2065 0 net=1107
rlabel metal2 331 -2065 331 -2065 0 net=3814
rlabel metal2 408 -2065 408 -2065 0 net=4715
rlabel metal2 135 -2067 135 -2067 0 net=3869
rlabel metal2 338 -2067 338 -2067 0 net=4259
rlabel metal2 499 -2067 499 -2067 0 net=719
rlabel metal2 156 -2069 156 -2069 0 net=4203
rlabel metal2 142 -2071 142 -2071 0 net=1247
rlabel metal2 159 -2071 159 -2071 0 net=3305
rlabel metal2 222 -2071 222 -2071 0 net=1411
rlabel metal2 254 -2071 254 -2071 0 net=2769
rlabel metal2 394 -2071 394 -2071 0 net=2817
rlabel metal2 226 -2073 226 -2073 0 net=2537
rlabel metal2 373 -2073 373 -2073 0 net=2555
rlabel metal2 268 -2075 268 -2075 0 net=2321
rlabel metal2 345 -2075 345 -2075 0 net=1951
rlabel metal2 394 -2075 394 -2075 0 net=2895
rlabel metal2 268 -2077 268 -2077 0 net=3049
rlabel metal2 401 -2077 401 -2077 0 net=4324
rlabel metal2 275 -2079 275 -2079 0 net=1567
rlabel metal2 317 -2081 317 -2081 0 net=2295
rlabel metal2 352 -2081 352 -2081 0 net=4057
rlabel metal2 317 -2083 317 -2083 0 net=4881
rlabel metal2 366 -2085 366 -2085 0 net=5142
rlabel metal2 282 -2087 282 -2087 0 net=911
rlabel metal2 282 -2089 282 -2089 0 net=1631
rlabel metal2 23 -2100 23 -2100 0 net=299
rlabel metal2 65 -2100 65 -2100 0 net=1766
rlabel metal2 324 -2100 324 -2100 0 net=1953
rlabel metal2 366 -2100 366 -2100 0 net=3995
rlabel metal2 429 -2100 429 -2100 0 net=3905
rlabel metal2 429 -2100 429 -2100 0 net=3905
rlabel metal2 509 -2100 509 -2100 0 net=4144
rlabel metal2 523 -2100 523 -2100 0 net=4908
rlabel metal2 590 -2100 590 -2100 0 net=1307
rlabel metal2 611 -2100 611 -2100 0 net=4610
rlabel metal2 642 -2100 642 -2100 0 net=4170
rlabel metal2 674 -2100 674 -2100 0 net=5352
rlabel metal2 26 -2102 26 -2102 0 net=474
rlabel metal2 100 -2102 100 -2102 0 net=1179
rlabel metal2 100 -2102 100 -2102 0 net=1179
rlabel metal2 107 -2102 107 -2102 0 net=2394
rlabel metal2 310 -2102 310 -2102 0 net=2323
rlabel metal2 345 -2102 345 -2102 0 net=3303
rlabel metal2 394 -2102 394 -2102 0 net=2897
rlabel metal2 530 -2102 530 -2102 0 net=5164
rlabel metal2 611 -2102 611 -2102 0 net=5137
rlabel metal2 33 -2104 33 -2104 0 net=1732
rlabel metal2 44 -2104 44 -2104 0 net=3628
rlabel metal2 331 -2104 331 -2104 0 net=2297
rlabel metal2 37 -2106 37 -2106 0 net=4277
rlabel metal2 135 -2106 135 -2106 0 net=3871
rlabel metal2 156 -2106 156 -2106 0 net=1163
rlabel metal2 187 -2106 187 -2106 0 net=799
rlabel metal2 338 -2106 338 -2106 0 net=3985
rlabel metal2 387 -2106 387 -2106 0 net=2735
rlabel metal2 534 -2106 534 -2106 0 net=4883
rlabel metal2 562 -2106 562 -2106 0 net=4789
rlabel metal2 44 -2108 44 -2108 0 net=1091
rlabel metal2 208 -2108 208 -2108 0 net=3050
rlabel metal2 282 -2108 282 -2108 0 net=1633
rlabel metal2 359 -2108 359 -2108 0 net=2701
rlabel metal2 464 -2108 464 -2108 0 net=4059
rlabel metal2 541 -2108 541 -2108 0 net=4595
rlabel metal2 541 -2108 541 -2108 0 net=4595
rlabel metal2 51 -2110 51 -2110 0 net=4038
rlabel metal2 163 -2110 163 -2110 0 net=3306
rlabel metal2 215 -2110 215 -2110 0 net=4716
rlabel metal2 51 -2112 51 -2112 0 net=2343
rlabel metal2 205 -2112 205 -2112 0 net=1641
rlabel metal2 222 -2112 222 -2112 0 net=740
rlabel metal2 58 -2114 58 -2114 0 net=3073
rlabel metal2 107 -2114 107 -2114 0 net=2471
rlabel metal2 135 -2114 135 -2114 0 net=1249
rlabel metal2 149 -2114 149 -2114 0 net=1565
rlabel metal2 170 -2114 170 -2114 0 net=1775
rlabel metal2 198 -2114 198 -2114 0 net=1071
rlabel metal2 296 -2114 296 -2114 0 net=3045
rlabel metal2 296 -2114 296 -2114 0 net=3045
rlabel metal2 303 -2114 303 -2114 0 net=2545
rlabel metal2 65 -2116 65 -2116 0 net=1749
rlabel metal2 86 -2116 86 -2116 0 net=2539
rlabel metal2 233 -2116 233 -2116 0 net=1108
rlabel metal2 247 -2116 247 -2116 0 net=1412
rlabel metal2 16 -2118 16 -2118 0 net=4510
rlabel metal2 170 -2118 170 -2118 0 net=2237
rlabel metal2 268 -2118 268 -2118 0 net=2447
rlabel metal2 369 -2118 369 -2118 0 net=2818
rlabel metal2 72 -2120 72 -2120 0 net=758
rlabel metal2 177 -2120 177 -2120 0 net=4665
rlabel metal2 117 -2122 117 -2122 0 net=967
rlabel metal2 233 -2124 233 -2124 0 net=1569
rlabel metal2 240 -2126 240 -2126 0 net=4119
rlabel metal2 247 -2128 247 -2128 0 net=3285
rlabel metal2 254 -2130 254 -2130 0 net=2770
rlabel metal2 443 -2130 443 -2130 0 net=3367
rlabel metal2 226 -2132 226 -2132 0 net=4205
rlabel metal2 261 -2132 261 -2132 0 net=2355
rlabel metal2 450 -2132 450 -2132 0 net=3823
rlabel metal2 261 -2134 261 -2134 0 net=4644
rlabel metal2 422 -2136 422 -2136 0 net=4039
rlabel metal2 513 -2136 513 -2136 0 net=4295
rlabel metal2 422 -2138 422 -2138 0 net=3203
rlabel metal2 492 -2138 492 -2138 0 net=4261
rlabel metal2 373 -2140 373 -2140 0 net=2557
rlabel metal2 492 -2140 492 -2140 0 net=4365
rlabel metal2 373 -2142 373 -2142 0 net=4204
rlabel metal2 457 -2144 457 -2144 0 net=4245
rlabel metal2 485 -2146 485 -2146 0 net=5355
rlabel metal2 9 -2157 9 -2157 0 net=4493
rlabel metal2 37 -2157 37 -2157 0 net=4278
rlabel metal2 240 -2157 240 -2157 0 net=4120
rlabel metal2 285 -2157 285 -2157 0 net=3046
rlabel metal2 317 -2157 317 -2157 0 net=3996
rlabel metal2 415 -2157 415 -2157 0 net=4262
rlabel metal2 590 -2157 590 -2157 0 net=4791
rlabel metal2 611 -2157 611 -2157 0 net=5139
rlabel metal2 611 -2157 611 -2157 0 net=5139
rlabel metal2 44 -2159 44 -2159 0 net=1092
rlabel metal2 208 -2159 208 -2159 0 net=1859
rlabel metal2 292 -2159 292 -2159 0 net=2324
rlabel metal2 317 -2159 317 -2159 0 net=2703
rlabel metal2 408 -2159 408 -2159 0 net=3369
rlabel metal2 450 -2159 450 -2159 0 net=3824
rlabel metal2 499 -2159 499 -2159 0 net=4884
rlabel metal2 597 -2159 597 -2159 0 net=1308
rlabel metal2 51 -2161 51 -2161 0 net=2345
rlabel metal2 275 -2161 275 -2161 0 net=2356
rlabel metal2 324 -2161 324 -2161 0 net=1954
rlabel metal2 352 -2161 352 -2161 0 net=1634
rlabel metal2 362 -2161 362 -2161 0 net=5356
rlabel metal2 541 -2161 541 -2161 0 net=4597
rlabel metal2 51 -2163 51 -2163 0 net=2797
rlabel metal2 163 -2163 163 -2163 0 net=1566
rlabel metal2 247 -2163 247 -2163 0 net=3286
rlabel metal2 387 -2163 387 -2163 0 net=3205
rlabel metal2 425 -2163 425 -2163 0 net=4666
rlabel metal2 58 -2165 58 -2165 0 net=3074
rlabel metal2 107 -2165 107 -2165 0 net=2472
rlabel metal2 131 -2165 131 -2165 0 net=1250
rlabel metal2 163 -2165 163 -2165 0 net=1523
rlabel metal2 268 -2165 268 -2165 0 net=2449
rlabel metal2 324 -2165 324 -2165 0 net=3304
rlabel metal2 352 -2165 352 -2165 0 net=2299
rlabel metal2 58 -2167 58 -2167 0 net=3845
rlabel metal2 278 -2167 278 -2167 0 net=412
rlabel metal2 366 -2167 366 -2167 0 net=2546
rlabel metal2 65 -2169 65 -2169 0 net=1750
rlabel metal2 79 -2169 79 -2169 0 net=1165
rlabel metal2 177 -2169 177 -2169 0 net=1911
rlabel metal2 345 -2169 345 -2169 0 net=4060
rlabel metal2 40 -2171 40 -2171 0 net=5283
rlabel metal2 86 -2171 86 -2171 0 net=2541
rlabel metal2 296 -2171 296 -2171 0 net=5421
rlabel metal2 513 -2171 513 -2171 0 net=4297
rlabel metal2 65 -2173 65 -2173 0 net=1807
rlabel metal2 331 -2173 331 -2173 0 net=2737
rlabel metal2 415 -2173 415 -2173 0 net=2771
rlabel metal2 86 -2175 86 -2175 0 net=3873
rlabel metal2 156 -2175 156 -2175 0 net=2239
rlabel metal2 219 -2175 219 -2175 0 net=2413
rlabel metal2 394 -2175 394 -2175 0 net=3307
rlabel metal2 93 -2177 93 -2177 0 net=1180
rlabel metal2 107 -2177 107 -2177 0 net=2209
rlabel metal2 135 -2177 135 -2177 0 net=709
rlabel metal2 429 -2177 429 -2177 0 net=3907
rlabel metal2 453 -2177 453 -2177 0 net=4040
rlabel metal2 93 -2179 93 -2179 0 net=1825
rlabel metal2 205 -2179 205 -2179 0 net=1642
rlabel metal2 429 -2179 429 -2179 0 net=4367
rlabel metal2 100 -2181 100 -2181 0 net=1073
rlabel metal2 380 -2181 380 -2181 0 net=3986
rlabel metal2 121 -2183 121 -2183 0 net=1570
rlabel metal2 380 -2183 380 -2183 0 net=2899
rlabel metal2 436 -2183 436 -2183 0 net=2558
rlabel metal2 121 -2185 121 -2185 0 net=1795
rlabel metal2 170 -2185 170 -2185 0 net=1081
rlabel metal2 436 -2185 436 -2185 0 net=4247
rlabel metal2 198 -2187 198 -2187 0 net=3225
rlabel metal2 457 -2187 457 -2187 0 net=4727
rlabel metal2 226 -2189 226 -2189 0 net=4207
rlabel metal2 191 -2191 191 -2191 0 net=1777
rlabel metal2 187 -2193 187 -2193 0 net=2127
rlabel metal2 9 -2204 9 -2204 0 net=4494
rlabel metal2 23 -2204 23 -2204 0 net=279
rlabel metal2 44 -2204 44 -2204 0 net=465
rlabel metal2 44 -2204 44 -2204 0 net=465
rlabel metal2 51 -2204 51 -2204 0 net=2798
rlabel metal2 107 -2204 107 -2204 0 net=2210
rlabel metal2 240 -2204 240 -2204 0 net=2901
rlabel metal2 408 -2204 408 -2204 0 net=3370
rlabel metal2 429 -2204 429 -2204 0 net=4369
rlabel metal2 457 -2204 457 -2204 0 net=4729
rlabel metal2 534 -2204 534 -2204 0 net=4298
rlabel metal2 600 -2204 600 -2204 0 net=4792
rlabel metal2 611 -2204 611 -2204 0 net=5140
rlabel metal2 611 -2204 611 -2204 0 net=5140
rlabel metal2 51 -2206 51 -2206 0 net=689
rlabel metal2 86 -2206 86 -2206 0 net=3874
rlabel metal2 254 -2206 254 -2206 0 net=5422
rlabel metal2 537 -2206 537 -2206 0 net=4598
rlabel metal2 58 -2208 58 -2208 0 net=3846
rlabel metal2 149 -2208 149 -2208 0 net=2240
rlabel metal2 177 -2208 177 -2208 0 net=1912
rlabel metal2 254 -2208 254 -2208 0 net=1861
rlabel metal2 299 -2208 299 -2208 0 net=133
rlabel metal2 366 -2208 366 -2208 0 net=3206
rlabel metal2 394 -2208 394 -2208 0 net=3309
rlabel metal2 422 -2208 422 -2208 0 net=234
rlabel metal2 58 -2210 58 -2210 0 net=1827
rlabel metal2 100 -2210 100 -2210 0 net=1074
rlabel metal2 247 -2210 247 -2210 0 net=3227
rlabel metal2 303 -2210 303 -2210 0 net=2450
rlabel metal2 359 -2210 359 -2210 0 net=2772
rlabel metal2 65 -2212 65 -2212 0 net=1808
rlabel metal2 149 -2212 149 -2212 0 net=1525
rlabel metal2 177 -2212 177 -2212 0 net=2346
rlabel metal2 268 -2212 268 -2212 0 net=2542
rlabel metal2 373 -2212 373 -2212 0 net=4249
rlabel metal2 443 -2212 443 -2212 0 net=3908
rlabel metal2 79 -2214 79 -2214 0 net=1166
rlabel metal2 247 -2214 247 -2214 0 net=2705
rlabel metal2 324 -2214 324 -2214 0 net=2300
rlabel metal2 107 -2216 107 -2216 0 net=1083
rlabel metal2 187 -2216 187 -2216 0 net=2414
rlabel metal2 268 -2216 268 -2216 0 net=4959
rlabel metal2 114 -2218 114 -2218 0 net=1796
rlabel metal2 191 -2218 191 -2218 0 net=2129
rlabel metal2 72 -2220 72 -2220 0 net=5285
rlabel metal2 191 -2220 191 -2220 0 net=1778
rlabel metal2 275 -2220 275 -2220 0 net=2739
rlabel metal2 226 -2222 226 -2222 0 net=1589
rlabel metal2 331 -2222 331 -2222 0 net=4209
rlabel metal2 58 -2233 58 -2233 0 net=1828
rlabel metal2 107 -2233 107 -2233 0 net=1084
rlabel metal2 201 -2233 201 -2233 0 net=4960
rlabel metal2 275 -2233 275 -2233 0 net=2740
rlabel metal2 331 -2233 331 -2233 0 net=4210
rlabel metal2 408 -2233 408 -2233 0 net=3310
rlabel metal2 450 -2233 450 -2233 0 net=4370
rlabel metal2 485 -2233 485 -2233 0 net=4730
rlabel metal2 75 -2235 75 -2235 0 net=5286
rlabel metal2 131 -2235 131 -2235 0 net=1590
rlabel metal2 240 -2235 240 -2235 0 net=2902
rlabel metal2 149 -2237 149 -2237 0 net=1526
rlabel metal2 219 -2237 219 -2237 0 net=2130
rlabel metal2 289 -2237 289 -2237 0 net=3228
rlabel metal2 310 -2237 310 -2237 0 net=4250
rlabel metal2 247 -2239 247 -2239 0 net=2706
rlabel metal2 254 -2241 254 -2241 0 net=1862
<< end >>
