magic
tech scmos
timestamp 1555017187 
<< pdiffusion >>
rect 1 -12 7 -6
rect 8 -12 14 -6
rect 15 -12 21 -6
rect 22 -12 28 -6
rect 113 -12 119 -6
rect 120 -12 123 -6
rect 127 -12 133 -6
rect 134 -12 137 -6
rect 141 -12 147 -6
rect 148 -12 154 -6
rect 155 -12 158 -6
rect 162 -12 168 -6
rect 169 -12 175 -6
rect 176 -12 179 -6
rect 183 -12 189 -6
rect 190 -12 193 -6
rect 197 -12 203 -6
rect 204 -12 210 -6
rect 211 -12 217 -6
rect 232 -12 238 -6
rect 246 -12 249 -6
rect 295 -12 298 -6
rect 309 -12 315 -6
rect 316 -12 319 -6
rect 330 -12 333 -6
rect 337 -12 343 -6
rect 344 -12 350 -6
rect 351 -12 354 -6
rect 372 -12 378 -6
rect 421 -12 427 -6
rect 1 -31 7 -25
rect 8 -31 14 -25
rect 64 -31 70 -25
rect 71 -31 74 -25
rect 78 -31 81 -25
rect 85 -31 91 -25
rect 92 -31 98 -25
rect 99 -31 102 -25
rect 106 -31 109 -25
rect 113 -31 119 -25
rect 120 -31 126 -25
rect 127 -31 133 -25
rect 134 -31 137 -25
rect 141 -31 144 -25
rect 148 -31 151 -25
rect 155 -31 161 -25
rect 162 -31 168 -25
rect 169 -31 172 -25
rect 176 -31 179 -25
rect 183 -31 186 -25
rect 190 -31 193 -25
rect 197 -31 203 -25
rect 204 -31 210 -25
rect 211 -31 214 -25
rect 218 -31 224 -25
rect 225 -31 231 -25
rect 232 -31 235 -25
rect 239 -31 242 -25
rect 246 -31 252 -25
rect 253 -31 256 -25
rect 260 -31 266 -25
rect 281 -31 284 -25
rect 295 -31 298 -25
rect 302 -31 305 -25
rect 309 -31 315 -25
rect 323 -31 329 -25
rect 330 -31 333 -25
rect 344 -31 347 -25
rect 351 -31 354 -25
rect 393 -31 396 -25
rect 400 -31 406 -25
rect 428 -31 431 -25
rect 435 -31 438 -25
rect 484 -31 490 -25
rect 554 -31 557 -25
rect 1 -60 7 -54
rect 8 -60 14 -54
rect 15 -60 21 -54
rect 22 -60 28 -54
rect 50 -60 53 -54
rect 57 -60 63 -54
rect 64 -60 67 -54
rect 71 -60 74 -54
rect 78 -60 84 -54
rect 85 -60 88 -54
rect 92 -60 95 -54
rect 99 -60 105 -54
rect 106 -60 109 -54
rect 113 -60 116 -54
rect 120 -60 123 -54
rect 127 -60 133 -54
rect 134 -60 137 -54
rect 141 -60 144 -54
rect 148 -60 151 -54
rect 155 -60 161 -54
rect 162 -60 165 -54
rect 169 -60 172 -54
rect 176 -60 179 -54
rect 183 -60 186 -54
rect 190 -60 196 -54
rect 197 -60 200 -54
rect 204 -60 207 -54
rect 211 -60 217 -54
rect 218 -60 221 -54
rect 225 -60 231 -54
rect 232 -60 235 -54
rect 239 -60 245 -54
rect 246 -60 249 -54
rect 253 -60 256 -54
rect 260 -60 263 -54
rect 267 -60 270 -54
rect 274 -60 277 -54
rect 281 -60 287 -54
rect 288 -60 291 -54
rect 295 -60 298 -54
rect 302 -60 308 -54
rect 309 -60 315 -54
rect 316 -60 322 -54
rect 323 -60 326 -54
rect 330 -60 333 -54
rect 337 -60 340 -54
rect 344 -60 347 -54
rect 351 -60 354 -54
rect 358 -60 361 -54
rect 365 -60 368 -54
rect 372 -60 375 -54
rect 379 -60 385 -54
rect 386 -60 389 -54
rect 393 -60 396 -54
rect 400 -60 406 -54
rect 414 -60 417 -54
rect 442 -60 445 -54
rect 449 -60 452 -54
rect 456 -60 462 -54
rect 575 -60 578 -54
rect 29 -99 32 -93
rect 36 -99 39 -93
rect 43 -99 46 -93
rect 50 -99 53 -93
rect 57 -99 60 -93
rect 64 -99 70 -93
rect 71 -99 74 -93
rect 78 -99 84 -93
rect 85 -99 88 -93
rect 92 -99 98 -93
rect 99 -99 102 -93
rect 106 -99 109 -93
rect 113 -99 116 -93
rect 120 -99 126 -93
rect 127 -99 133 -93
rect 134 -99 137 -93
rect 141 -99 144 -93
rect 148 -99 154 -93
rect 155 -99 161 -93
rect 162 -99 165 -93
rect 169 -99 172 -93
rect 176 -99 179 -93
rect 183 -99 186 -93
rect 190 -99 193 -93
rect 197 -99 200 -93
rect 204 -99 207 -93
rect 211 -99 214 -93
rect 218 -99 221 -93
rect 225 -99 228 -93
rect 232 -99 235 -93
rect 239 -99 245 -93
rect 246 -99 249 -93
rect 253 -99 259 -93
rect 260 -99 263 -93
rect 267 -99 270 -93
rect 274 -99 277 -93
rect 281 -99 287 -93
rect 288 -99 291 -93
rect 295 -99 298 -93
rect 302 -99 305 -93
rect 309 -99 315 -93
rect 316 -99 322 -93
rect 323 -99 326 -93
rect 330 -99 333 -93
rect 337 -99 340 -93
rect 344 -99 347 -93
rect 351 -99 357 -93
rect 358 -99 361 -93
rect 365 -99 371 -93
rect 372 -99 378 -93
rect 379 -99 382 -93
rect 386 -99 389 -93
rect 393 -99 396 -93
rect 400 -99 403 -93
rect 407 -99 410 -93
rect 414 -99 417 -93
rect 421 -99 427 -93
rect 428 -99 431 -93
rect 435 -99 438 -93
rect 442 -99 448 -93
rect 449 -99 452 -93
rect 456 -99 462 -93
rect 463 -99 466 -93
rect 470 -99 473 -93
rect 477 -99 480 -93
rect 491 -99 494 -93
rect 519 -99 525 -93
rect 526 -99 532 -93
rect 575 -99 578 -93
rect 589 -99 592 -93
rect 1 -150 7 -144
rect 8 -150 11 -144
rect 15 -150 18 -144
rect 22 -150 28 -144
rect 29 -150 32 -144
rect 36 -150 39 -144
rect 43 -150 46 -144
rect 50 -150 53 -144
rect 57 -150 60 -144
rect 64 -150 67 -144
rect 71 -150 77 -144
rect 78 -150 84 -144
rect 85 -150 91 -144
rect 92 -150 98 -144
rect 99 -150 102 -144
rect 106 -150 109 -144
rect 113 -150 116 -144
rect 120 -150 123 -144
rect 127 -150 130 -144
rect 134 -150 137 -144
rect 141 -150 144 -144
rect 148 -150 151 -144
rect 155 -150 158 -144
rect 162 -150 168 -144
rect 169 -150 175 -144
rect 176 -150 179 -144
rect 183 -150 186 -144
rect 190 -150 193 -144
rect 197 -150 200 -144
rect 204 -150 207 -144
rect 211 -150 214 -144
rect 218 -150 224 -144
rect 225 -150 228 -144
rect 232 -150 235 -144
rect 239 -150 242 -144
rect 246 -150 249 -144
rect 253 -150 259 -144
rect 260 -150 266 -144
rect 267 -150 270 -144
rect 274 -150 280 -144
rect 281 -150 284 -144
rect 288 -150 294 -144
rect 295 -150 298 -144
rect 302 -150 305 -144
rect 309 -150 315 -144
rect 316 -150 322 -144
rect 323 -150 326 -144
rect 330 -150 333 -144
rect 337 -150 340 -144
rect 344 -150 347 -144
rect 351 -150 354 -144
rect 358 -150 361 -144
rect 365 -150 368 -144
rect 372 -150 375 -144
rect 379 -150 382 -144
rect 386 -150 389 -144
rect 393 -150 396 -144
rect 400 -150 403 -144
rect 407 -150 410 -144
rect 414 -150 420 -144
rect 421 -150 424 -144
rect 428 -150 431 -144
rect 435 -150 438 -144
rect 442 -150 445 -144
rect 449 -150 452 -144
rect 456 -150 459 -144
rect 463 -150 466 -144
rect 470 -150 476 -144
rect 477 -150 480 -144
rect 484 -150 487 -144
rect 491 -150 494 -144
rect 498 -150 504 -144
rect 505 -150 508 -144
rect 512 -150 515 -144
rect 519 -150 522 -144
rect 526 -150 529 -144
rect 533 -150 536 -144
rect 540 -150 543 -144
rect 547 -150 550 -144
rect 554 -150 557 -144
rect 561 -150 564 -144
rect 568 -150 571 -144
rect 575 -150 578 -144
rect 582 -150 588 -144
rect 589 -150 592 -144
rect 596 -150 599 -144
rect 603 -150 606 -144
rect 610 -150 613 -144
rect 617 -150 620 -144
rect 624 -150 630 -144
rect 1 -211 7 -205
rect 8 -211 14 -205
rect 15 -211 18 -205
rect 22 -211 25 -205
rect 29 -211 32 -205
rect 36 -211 39 -205
rect 43 -211 46 -205
rect 50 -211 53 -205
rect 57 -211 60 -205
rect 64 -211 67 -205
rect 71 -211 77 -205
rect 78 -211 81 -205
rect 85 -211 88 -205
rect 92 -211 98 -205
rect 99 -211 105 -205
rect 106 -211 109 -205
rect 113 -211 116 -205
rect 120 -211 123 -205
rect 127 -211 130 -205
rect 134 -211 140 -205
rect 141 -211 144 -205
rect 148 -211 151 -205
rect 155 -211 158 -205
rect 162 -211 165 -205
rect 169 -211 172 -205
rect 176 -211 182 -205
rect 183 -211 186 -205
rect 190 -211 193 -205
rect 197 -211 200 -205
rect 204 -211 210 -205
rect 211 -211 217 -205
rect 218 -211 221 -205
rect 225 -211 228 -205
rect 232 -211 235 -205
rect 239 -211 242 -205
rect 246 -211 249 -205
rect 253 -211 256 -205
rect 260 -211 263 -205
rect 267 -211 270 -205
rect 274 -211 280 -205
rect 281 -211 284 -205
rect 288 -211 291 -205
rect 295 -211 301 -205
rect 302 -211 308 -205
rect 309 -211 312 -205
rect 316 -211 322 -205
rect 323 -211 329 -205
rect 330 -211 336 -205
rect 337 -211 343 -205
rect 344 -211 347 -205
rect 351 -211 354 -205
rect 358 -211 361 -205
rect 365 -211 371 -205
rect 372 -211 375 -205
rect 379 -211 382 -205
rect 386 -211 392 -205
rect 393 -211 396 -205
rect 400 -211 403 -205
rect 407 -211 410 -205
rect 414 -211 417 -205
rect 421 -211 424 -205
rect 428 -211 431 -205
rect 435 -211 438 -205
rect 442 -211 448 -205
rect 449 -211 452 -205
rect 456 -211 459 -205
rect 463 -211 466 -205
rect 470 -211 473 -205
rect 477 -211 480 -205
rect 484 -211 490 -205
rect 491 -211 494 -205
rect 498 -211 501 -205
rect 505 -211 508 -205
rect 512 -211 515 -205
rect 519 -211 522 -205
rect 526 -211 529 -205
rect 533 -211 536 -205
rect 540 -211 543 -205
rect 547 -211 550 -205
rect 554 -211 557 -205
rect 561 -211 564 -205
rect 568 -211 571 -205
rect 575 -211 578 -205
rect 582 -211 585 -205
rect 589 -211 592 -205
rect 596 -211 599 -205
rect 603 -211 606 -205
rect 610 -211 613 -205
rect 617 -211 620 -205
rect 624 -211 627 -205
rect 631 -211 634 -205
rect 638 -211 641 -205
rect 645 -211 648 -205
rect 652 -211 655 -205
rect 659 -211 662 -205
rect 666 -211 669 -205
rect 673 -211 676 -205
rect 1 -276 4 -270
rect 8 -276 14 -270
rect 15 -276 18 -270
rect 22 -276 25 -270
rect 29 -276 35 -270
rect 36 -276 39 -270
rect 43 -276 46 -270
rect 50 -276 56 -270
rect 57 -276 60 -270
rect 64 -276 67 -270
rect 71 -276 74 -270
rect 78 -276 84 -270
rect 85 -276 88 -270
rect 92 -276 95 -270
rect 99 -276 105 -270
rect 106 -276 112 -270
rect 113 -276 119 -270
rect 120 -276 123 -270
rect 127 -276 130 -270
rect 134 -276 137 -270
rect 141 -276 144 -270
rect 148 -276 154 -270
rect 155 -276 158 -270
rect 162 -276 165 -270
rect 169 -276 172 -270
rect 176 -276 179 -270
rect 183 -276 186 -270
rect 190 -276 193 -270
rect 197 -276 200 -270
rect 204 -276 207 -270
rect 211 -276 214 -270
rect 218 -276 221 -270
rect 225 -276 228 -270
rect 232 -276 235 -270
rect 239 -276 245 -270
rect 246 -276 252 -270
rect 253 -276 256 -270
rect 260 -276 266 -270
rect 267 -276 270 -270
rect 274 -276 280 -270
rect 281 -276 284 -270
rect 288 -276 294 -270
rect 295 -276 301 -270
rect 302 -276 305 -270
rect 309 -276 315 -270
rect 316 -276 319 -270
rect 323 -276 326 -270
rect 330 -276 333 -270
rect 337 -276 340 -270
rect 344 -276 347 -270
rect 351 -276 354 -270
rect 358 -276 361 -270
rect 365 -276 371 -270
rect 372 -276 375 -270
rect 379 -276 385 -270
rect 386 -276 389 -270
rect 393 -276 396 -270
rect 400 -276 403 -270
rect 407 -276 410 -270
rect 414 -276 417 -270
rect 421 -276 424 -270
rect 428 -276 431 -270
rect 435 -276 438 -270
rect 442 -276 445 -270
rect 449 -276 452 -270
rect 456 -276 459 -270
rect 463 -276 469 -270
rect 470 -276 473 -270
rect 477 -276 480 -270
rect 484 -276 487 -270
rect 491 -276 494 -270
rect 498 -276 501 -270
rect 505 -276 508 -270
rect 512 -276 515 -270
rect 519 -276 522 -270
rect 526 -276 529 -270
rect 533 -276 536 -270
rect 540 -276 543 -270
rect 547 -276 550 -270
rect 554 -276 557 -270
rect 561 -276 564 -270
rect 568 -276 571 -270
rect 575 -276 578 -270
rect 582 -276 585 -270
rect 589 -276 592 -270
rect 596 -276 599 -270
rect 603 -276 606 -270
rect 610 -276 613 -270
rect 617 -276 620 -270
rect 624 -276 627 -270
rect 631 -276 634 -270
rect 638 -276 641 -270
rect 645 -276 648 -270
rect 652 -276 655 -270
rect 659 -276 662 -270
rect 666 -276 669 -270
rect 673 -276 676 -270
rect 680 -276 683 -270
rect 687 -276 690 -270
rect 694 -276 697 -270
rect 701 -276 704 -270
rect 708 -276 714 -270
rect 715 -276 718 -270
rect 722 -276 725 -270
rect 729 -276 735 -270
rect 1 -343 7 -337
rect 8 -343 14 -337
rect 15 -343 18 -337
rect 22 -343 28 -337
rect 29 -343 32 -337
rect 36 -343 39 -337
rect 43 -343 49 -337
rect 50 -343 56 -337
rect 57 -343 63 -337
rect 64 -343 67 -337
rect 71 -343 74 -337
rect 78 -343 81 -337
rect 85 -343 88 -337
rect 92 -343 95 -337
rect 99 -343 102 -337
rect 106 -343 112 -337
rect 113 -343 116 -337
rect 120 -343 123 -337
rect 127 -343 130 -337
rect 134 -343 137 -337
rect 141 -343 144 -337
rect 148 -343 151 -337
rect 155 -343 158 -337
rect 162 -343 168 -337
rect 169 -343 172 -337
rect 176 -343 179 -337
rect 183 -343 189 -337
rect 190 -343 193 -337
rect 197 -343 200 -337
rect 204 -343 207 -337
rect 211 -343 214 -337
rect 218 -343 221 -337
rect 225 -343 231 -337
rect 232 -343 235 -337
rect 239 -343 242 -337
rect 246 -343 249 -337
rect 253 -343 259 -337
rect 260 -343 263 -337
rect 267 -343 270 -337
rect 274 -343 280 -337
rect 281 -343 287 -337
rect 288 -343 291 -337
rect 295 -343 301 -337
rect 302 -343 305 -337
rect 309 -343 312 -337
rect 316 -343 319 -337
rect 323 -343 329 -337
rect 330 -343 333 -337
rect 337 -343 340 -337
rect 344 -343 350 -337
rect 351 -343 354 -337
rect 358 -343 364 -337
rect 365 -343 371 -337
rect 372 -343 375 -337
rect 379 -343 382 -337
rect 386 -343 389 -337
rect 393 -343 396 -337
rect 400 -343 406 -337
rect 407 -343 410 -337
rect 414 -343 417 -337
rect 421 -343 424 -337
rect 428 -343 434 -337
rect 435 -343 438 -337
rect 442 -343 445 -337
rect 449 -343 452 -337
rect 456 -343 459 -337
rect 463 -343 466 -337
rect 470 -343 473 -337
rect 477 -343 480 -337
rect 484 -343 487 -337
rect 491 -343 494 -337
rect 498 -343 501 -337
rect 505 -343 508 -337
rect 512 -343 515 -337
rect 519 -343 522 -337
rect 526 -343 529 -337
rect 533 -343 536 -337
rect 540 -343 543 -337
rect 547 -343 550 -337
rect 554 -343 557 -337
rect 561 -343 564 -337
rect 568 -343 571 -337
rect 575 -343 578 -337
rect 582 -343 585 -337
rect 589 -343 592 -337
rect 596 -343 599 -337
rect 603 -343 606 -337
rect 610 -343 613 -337
rect 617 -343 620 -337
rect 624 -343 627 -337
rect 631 -343 634 -337
rect 638 -343 641 -337
rect 645 -343 648 -337
rect 652 -343 655 -337
rect 659 -343 662 -337
rect 666 -343 669 -337
rect 673 -343 676 -337
rect 680 -343 683 -337
rect 687 -343 690 -337
rect 694 -343 697 -337
rect 701 -343 704 -337
rect 708 -343 711 -337
rect 715 -343 718 -337
rect 722 -343 725 -337
rect 729 -343 732 -337
rect 736 -343 739 -337
rect 1 -422 7 -416
rect 8 -422 14 -416
rect 15 -422 18 -416
rect 22 -422 25 -416
rect 29 -422 32 -416
rect 36 -422 39 -416
rect 43 -422 46 -416
rect 50 -422 53 -416
rect 57 -422 63 -416
rect 64 -422 67 -416
rect 71 -422 74 -416
rect 78 -422 81 -416
rect 85 -422 88 -416
rect 92 -422 95 -416
rect 99 -422 102 -416
rect 106 -422 112 -416
rect 113 -422 116 -416
rect 120 -422 126 -416
rect 127 -422 130 -416
rect 134 -422 137 -416
rect 141 -422 144 -416
rect 148 -422 151 -416
rect 155 -422 158 -416
rect 162 -422 165 -416
rect 169 -422 172 -416
rect 176 -422 179 -416
rect 183 -422 186 -416
rect 190 -422 193 -416
rect 197 -422 200 -416
rect 204 -422 207 -416
rect 211 -422 214 -416
rect 218 -422 224 -416
rect 225 -422 228 -416
rect 232 -422 235 -416
rect 239 -422 242 -416
rect 246 -422 249 -416
rect 253 -422 256 -416
rect 260 -422 263 -416
rect 267 -422 270 -416
rect 274 -422 277 -416
rect 281 -422 284 -416
rect 288 -422 294 -416
rect 295 -422 298 -416
rect 302 -422 305 -416
rect 309 -422 312 -416
rect 316 -422 319 -416
rect 323 -422 326 -416
rect 330 -422 336 -416
rect 337 -422 343 -416
rect 344 -422 350 -416
rect 351 -422 354 -416
rect 358 -422 361 -416
rect 365 -422 368 -416
rect 372 -422 378 -416
rect 379 -422 385 -416
rect 386 -422 389 -416
rect 393 -422 399 -416
rect 400 -422 406 -416
rect 407 -422 410 -416
rect 414 -422 420 -416
rect 421 -422 424 -416
rect 428 -422 434 -416
rect 435 -422 438 -416
rect 442 -422 445 -416
rect 449 -422 452 -416
rect 456 -422 459 -416
rect 463 -422 466 -416
rect 470 -422 476 -416
rect 477 -422 480 -416
rect 484 -422 487 -416
rect 491 -422 494 -416
rect 498 -422 501 -416
rect 505 -422 511 -416
rect 512 -422 515 -416
rect 519 -422 525 -416
rect 526 -422 529 -416
rect 533 -422 536 -416
rect 540 -422 543 -416
rect 547 -422 550 -416
rect 554 -422 560 -416
rect 561 -422 564 -416
rect 568 -422 571 -416
rect 575 -422 578 -416
rect 582 -422 585 -416
rect 589 -422 592 -416
rect 596 -422 599 -416
rect 603 -422 606 -416
rect 610 -422 613 -416
rect 617 -422 620 -416
rect 624 -422 627 -416
rect 631 -422 634 -416
rect 638 -422 641 -416
rect 645 -422 648 -416
rect 652 -422 655 -416
rect 659 -422 662 -416
rect 666 -422 669 -416
rect 673 -422 676 -416
rect 680 -422 683 -416
rect 687 -422 690 -416
rect 694 -422 697 -416
rect 701 -422 704 -416
rect 708 -422 711 -416
rect 715 -422 718 -416
rect 722 -422 725 -416
rect 729 -422 732 -416
rect 736 -422 739 -416
rect 743 -422 746 -416
rect 750 -422 753 -416
rect 757 -422 760 -416
rect 764 -422 767 -416
rect 771 -422 774 -416
rect 778 -422 781 -416
rect 785 -422 788 -416
rect 792 -422 795 -416
rect 799 -422 802 -416
rect 806 -422 809 -416
rect 813 -422 816 -416
rect 1 -515 7 -509
rect 8 -515 11 -509
rect 15 -515 18 -509
rect 22 -515 25 -509
rect 29 -515 32 -509
rect 36 -515 39 -509
rect 43 -515 49 -509
rect 50 -515 53 -509
rect 57 -515 63 -509
rect 64 -515 67 -509
rect 71 -515 74 -509
rect 78 -515 81 -509
rect 85 -515 88 -509
rect 92 -515 95 -509
rect 99 -515 105 -509
rect 106 -515 109 -509
rect 113 -515 116 -509
rect 120 -515 123 -509
rect 127 -515 130 -509
rect 134 -515 140 -509
rect 141 -515 144 -509
rect 148 -515 151 -509
rect 155 -515 158 -509
rect 162 -515 165 -509
rect 169 -515 172 -509
rect 176 -515 179 -509
rect 183 -515 186 -509
rect 190 -515 193 -509
rect 197 -515 200 -509
rect 204 -515 207 -509
rect 211 -515 214 -509
rect 218 -515 224 -509
rect 225 -515 231 -509
rect 232 -515 235 -509
rect 239 -515 242 -509
rect 246 -515 249 -509
rect 253 -515 256 -509
rect 260 -515 266 -509
rect 267 -515 270 -509
rect 274 -515 277 -509
rect 281 -515 284 -509
rect 288 -515 291 -509
rect 295 -515 298 -509
rect 302 -515 308 -509
rect 309 -515 315 -509
rect 316 -515 319 -509
rect 323 -515 326 -509
rect 330 -515 333 -509
rect 337 -515 340 -509
rect 344 -515 347 -509
rect 351 -515 357 -509
rect 358 -515 361 -509
rect 365 -515 371 -509
rect 372 -515 375 -509
rect 379 -515 385 -509
rect 386 -515 392 -509
rect 393 -515 396 -509
rect 400 -515 406 -509
rect 407 -515 413 -509
rect 414 -515 417 -509
rect 421 -515 424 -509
rect 428 -515 434 -509
rect 435 -515 438 -509
rect 442 -515 445 -509
rect 449 -515 452 -509
rect 456 -515 459 -509
rect 463 -515 466 -509
rect 470 -515 476 -509
rect 477 -515 480 -509
rect 484 -515 487 -509
rect 491 -515 497 -509
rect 498 -515 501 -509
rect 505 -515 508 -509
rect 512 -515 515 -509
rect 519 -515 522 -509
rect 526 -515 529 -509
rect 533 -515 536 -509
rect 540 -515 543 -509
rect 547 -515 550 -509
rect 554 -515 560 -509
rect 561 -515 564 -509
rect 568 -515 571 -509
rect 575 -515 578 -509
rect 582 -515 585 -509
rect 589 -515 592 -509
rect 596 -515 599 -509
rect 603 -515 606 -509
rect 610 -515 613 -509
rect 617 -515 620 -509
rect 624 -515 627 -509
rect 631 -515 634 -509
rect 638 -515 641 -509
rect 645 -515 648 -509
rect 652 -515 655 -509
rect 659 -515 662 -509
rect 666 -515 669 -509
rect 673 -515 676 -509
rect 680 -515 683 -509
rect 687 -515 690 -509
rect 694 -515 697 -509
rect 701 -515 704 -509
rect 708 -515 711 -509
rect 715 -515 718 -509
rect 722 -515 725 -509
rect 729 -515 732 -509
rect 736 -515 739 -509
rect 743 -515 746 -509
rect 750 -515 753 -509
rect 757 -515 760 -509
rect 764 -515 767 -509
rect 771 -515 774 -509
rect 778 -515 781 -509
rect 785 -515 788 -509
rect 792 -515 795 -509
rect 799 -515 802 -509
rect 1 -584 7 -578
rect 8 -584 11 -578
rect 15 -584 18 -578
rect 22 -584 28 -578
rect 29 -584 32 -578
rect 36 -584 39 -578
rect 43 -584 46 -578
rect 50 -584 56 -578
rect 57 -584 60 -578
rect 64 -584 67 -578
rect 71 -584 74 -578
rect 78 -584 81 -578
rect 85 -584 88 -578
rect 92 -584 95 -578
rect 99 -584 102 -578
rect 106 -584 112 -578
rect 113 -584 116 -578
rect 120 -584 126 -578
rect 127 -584 133 -578
rect 134 -584 140 -578
rect 141 -584 144 -578
rect 148 -584 151 -578
rect 155 -584 158 -578
rect 162 -584 165 -578
rect 169 -584 172 -578
rect 176 -584 179 -578
rect 183 -584 186 -578
rect 190 -584 193 -578
rect 197 -584 200 -578
rect 204 -584 207 -578
rect 211 -584 214 -578
rect 218 -584 221 -578
rect 225 -584 228 -578
rect 232 -584 235 -578
rect 239 -584 242 -578
rect 246 -584 249 -578
rect 253 -584 259 -578
rect 260 -584 263 -578
rect 267 -584 270 -578
rect 274 -584 277 -578
rect 281 -584 284 -578
rect 288 -584 291 -578
rect 295 -584 301 -578
rect 302 -584 305 -578
rect 309 -584 315 -578
rect 316 -584 322 -578
rect 323 -584 326 -578
rect 330 -584 336 -578
rect 337 -584 340 -578
rect 344 -584 347 -578
rect 351 -584 354 -578
rect 358 -584 361 -578
rect 365 -584 368 -578
rect 372 -584 375 -578
rect 379 -584 385 -578
rect 386 -584 389 -578
rect 393 -584 396 -578
rect 400 -584 403 -578
rect 407 -584 410 -578
rect 414 -584 420 -578
rect 421 -584 424 -578
rect 428 -584 431 -578
rect 435 -584 438 -578
rect 442 -584 445 -578
rect 449 -584 452 -578
rect 456 -584 462 -578
rect 463 -584 469 -578
rect 470 -584 473 -578
rect 477 -584 480 -578
rect 484 -584 490 -578
rect 491 -584 494 -578
rect 498 -584 501 -578
rect 505 -584 511 -578
rect 512 -584 518 -578
rect 519 -584 522 -578
rect 526 -584 529 -578
rect 533 -584 536 -578
rect 540 -584 543 -578
rect 547 -584 553 -578
rect 554 -584 557 -578
rect 561 -584 564 -578
rect 568 -584 571 -578
rect 575 -584 578 -578
rect 582 -584 585 -578
rect 589 -584 592 -578
rect 596 -584 599 -578
rect 603 -584 606 -578
rect 610 -584 613 -578
rect 617 -584 620 -578
rect 624 -584 627 -578
rect 631 -584 634 -578
rect 638 -584 641 -578
rect 645 -584 648 -578
rect 652 -584 655 -578
rect 659 -584 662 -578
rect 666 -584 669 -578
rect 673 -584 676 -578
rect 680 -584 683 -578
rect 687 -584 690 -578
rect 694 -584 697 -578
rect 701 -584 704 -578
rect 708 -584 711 -578
rect 715 -584 718 -578
rect 722 -584 725 -578
rect 729 -584 732 -578
rect 736 -584 739 -578
rect 743 -584 746 -578
rect 750 -584 753 -578
rect 757 -584 760 -578
rect 764 -584 767 -578
rect 771 -584 774 -578
rect 778 -584 781 -578
rect 785 -584 788 -578
rect 792 -584 795 -578
rect 799 -584 802 -578
rect 806 -584 809 -578
rect 813 -584 816 -578
rect 820 -584 823 -578
rect 1 -673 4 -667
rect 8 -673 11 -667
rect 15 -673 18 -667
rect 22 -673 25 -667
rect 29 -673 32 -667
rect 36 -673 39 -667
rect 43 -673 46 -667
rect 50 -673 56 -667
rect 57 -673 63 -667
rect 64 -673 70 -667
rect 71 -673 74 -667
rect 78 -673 81 -667
rect 85 -673 88 -667
rect 92 -673 95 -667
rect 99 -673 102 -667
rect 106 -673 112 -667
rect 113 -673 119 -667
rect 120 -673 123 -667
rect 127 -673 130 -667
rect 134 -673 137 -667
rect 141 -673 147 -667
rect 148 -673 151 -667
rect 155 -673 158 -667
rect 162 -673 165 -667
rect 169 -673 172 -667
rect 176 -673 179 -667
rect 183 -673 186 -667
rect 190 -673 193 -667
rect 197 -673 200 -667
rect 204 -673 207 -667
rect 211 -673 217 -667
rect 218 -673 221 -667
rect 225 -673 231 -667
rect 232 -673 235 -667
rect 239 -673 242 -667
rect 246 -673 249 -667
rect 253 -673 256 -667
rect 260 -673 263 -667
rect 267 -673 273 -667
rect 274 -673 277 -667
rect 281 -673 284 -667
rect 288 -673 294 -667
rect 295 -673 301 -667
rect 302 -673 305 -667
rect 309 -673 312 -667
rect 316 -673 319 -667
rect 323 -673 326 -667
rect 330 -673 333 -667
rect 337 -673 340 -667
rect 344 -673 350 -667
rect 351 -673 354 -667
rect 358 -673 361 -667
rect 365 -673 371 -667
rect 372 -673 375 -667
rect 379 -673 385 -667
rect 386 -673 389 -667
rect 393 -673 396 -667
rect 400 -673 403 -667
rect 407 -673 410 -667
rect 414 -673 420 -667
rect 421 -673 424 -667
rect 428 -673 431 -667
rect 435 -673 438 -667
rect 442 -673 445 -667
rect 449 -673 455 -667
rect 456 -673 462 -667
rect 463 -673 466 -667
rect 470 -673 473 -667
rect 477 -673 480 -667
rect 484 -673 487 -667
rect 491 -673 494 -667
rect 498 -673 501 -667
rect 505 -673 508 -667
rect 512 -673 515 -667
rect 519 -673 522 -667
rect 526 -673 529 -667
rect 533 -673 536 -667
rect 540 -673 546 -667
rect 547 -673 550 -667
rect 554 -673 557 -667
rect 561 -673 564 -667
rect 568 -673 571 -667
rect 575 -673 578 -667
rect 582 -673 585 -667
rect 589 -673 592 -667
rect 596 -673 599 -667
rect 603 -673 606 -667
rect 610 -673 613 -667
rect 617 -673 620 -667
rect 624 -673 627 -667
rect 631 -673 634 -667
rect 638 -673 641 -667
rect 645 -673 648 -667
rect 652 -673 655 -667
rect 659 -673 662 -667
rect 666 -673 669 -667
rect 673 -673 676 -667
rect 680 -673 683 -667
rect 687 -673 690 -667
rect 694 -673 697 -667
rect 701 -673 704 -667
rect 708 -673 711 -667
rect 715 -673 718 -667
rect 722 -673 725 -667
rect 729 -673 732 -667
rect 736 -673 739 -667
rect 743 -673 746 -667
rect 750 -673 753 -667
rect 757 -673 760 -667
rect 764 -673 767 -667
rect 771 -673 774 -667
rect 778 -673 781 -667
rect 785 -673 791 -667
rect 792 -673 798 -667
rect 8 -740 14 -734
rect 15 -740 21 -734
rect 22 -740 25 -734
rect 29 -740 32 -734
rect 36 -740 39 -734
rect 43 -740 46 -734
rect 50 -740 53 -734
rect 57 -740 60 -734
rect 64 -740 70 -734
rect 71 -740 74 -734
rect 78 -740 81 -734
rect 85 -740 91 -734
rect 92 -740 95 -734
rect 99 -740 102 -734
rect 106 -740 109 -734
rect 113 -740 116 -734
rect 120 -740 123 -734
rect 127 -740 133 -734
rect 134 -740 137 -734
rect 141 -740 144 -734
rect 148 -740 151 -734
rect 155 -740 158 -734
rect 162 -740 168 -734
rect 169 -740 172 -734
rect 176 -740 179 -734
rect 183 -740 186 -734
rect 190 -740 193 -734
rect 197 -740 200 -734
rect 204 -740 207 -734
rect 211 -740 214 -734
rect 218 -740 221 -734
rect 225 -740 231 -734
rect 232 -740 235 -734
rect 239 -740 242 -734
rect 246 -740 249 -734
rect 253 -740 256 -734
rect 260 -740 263 -734
rect 267 -740 273 -734
rect 274 -740 277 -734
rect 281 -740 284 -734
rect 288 -740 291 -734
rect 295 -740 298 -734
rect 302 -740 305 -734
rect 309 -740 312 -734
rect 316 -740 322 -734
rect 323 -740 326 -734
rect 330 -740 333 -734
rect 337 -740 340 -734
rect 344 -740 350 -734
rect 351 -740 354 -734
rect 358 -740 361 -734
rect 365 -740 368 -734
rect 372 -740 375 -734
rect 379 -740 385 -734
rect 386 -740 389 -734
rect 393 -740 399 -734
rect 400 -740 403 -734
rect 407 -740 410 -734
rect 414 -740 417 -734
rect 421 -740 427 -734
rect 428 -740 431 -734
rect 435 -740 438 -734
rect 442 -740 448 -734
rect 449 -740 452 -734
rect 456 -740 459 -734
rect 463 -740 466 -734
rect 470 -740 473 -734
rect 477 -740 480 -734
rect 484 -740 487 -734
rect 491 -740 494 -734
rect 498 -740 501 -734
rect 505 -740 508 -734
rect 512 -740 515 -734
rect 519 -740 525 -734
rect 526 -740 532 -734
rect 533 -740 536 -734
rect 540 -740 543 -734
rect 547 -740 553 -734
rect 554 -740 557 -734
rect 561 -740 564 -734
rect 568 -740 574 -734
rect 575 -740 578 -734
rect 582 -740 585 -734
rect 589 -740 592 -734
rect 596 -740 599 -734
rect 603 -740 606 -734
rect 610 -740 613 -734
rect 617 -740 620 -734
rect 624 -740 627 -734
rect 631 -740 634 -734
rect 638 -740 641 -734
rect 645 -740 648 -734
rect 652 -740 655 -734
rect 659 -740 662 -734
rect 666 -740 669 -734
rect 673 -740 676 -734
rect 680 -740 683 -734
rect 687 -740 690 -734
rect 694 -740 697 -734
rect 701 -740 704 -734
rect 708 -740 711 -734
rect 715 -740 718 -734
rect 722 -740 725 -734
rect 729 -740 732 -734
rect 736 -740 739 -734
rect 743 -740 746 -734
rect 750 -740 753 -734
rect 757 -740 760 -734
rect 764 -740 767 -734
rect 771 -740 774 -734
rect 778 -740 784 -734
rect 785 -740 788 -734
rect 792 -740 798 -734
rect 799 -740 802 -734
rect 806 -740 809 -734
rect 1 -811 7 -805
rect 8 -811 11 -805
rect 15 -811 18 -805
rect 22 -811 25 -805
rect 29 -811 32 -805
rect 36 -811 42 -805
rect 43 -811 46 -805
rect 50 -811 53 -805
rect 57 -811 60 -805
rect 64 -811 67 -805
rect 71 -811 77 -805
rect 78 -811 81 -805
rect 85 -811 88 -805
rect 92 -811 95 -805
rect 99 -811 102 -805
rect 106 -811 109 -805
rect 113 -811 116 -805
rect 120 -811 123 -805
rect 127 -811 133 -805
rect 134 -811 137 -805
rect 141 -811 144 -805
rect 148 -811 151 -805
rect 155 -811 161 -805
rect 162 -811 165 -805
rect 169 -811 172 -805
rect 176 -811 179 -805
rect 183 -811 186 -805
rect 190 -811 193 -805
rect 197 -811 200 -805
rect 204 -811 207 -805
rect 211 -811 217 -805
rect 218 -811 221 -805
rect 225 -811 228 -805
rect 232 -811 235 -805
rect 239 -811 242 -805
rect 246 -811 252 -805
rect 253 -811 259 -805
rect 260 -811 263 -805
rect 267 -811 270 -805
rect 274 -811 277 -805
rect 281 -811 287 -805
rect 288 -811 291 -805
rect 295 -811 298 -805
rect 302 -811 305 -805
rect 309 -811 315 -805
rect 316 -811 319 -805
rect 323 -811 326 -805
rect 330 -811 333 -805
rect 337 -811 340 -805
rect 344 -811 347 -805
rect 351 -811 354 -805
rect 358 -811 364 -805
rect 365 -811 368 -805
rect 372 -811 378 -805
rect 379 -811 382 -805
rect 386 -811 389 -805
rect 393 -811 399 -805
rect 400 -811 406 -805
rect 407 -811 413 -805
rect 414 -811 417 -805
rect 421 -811 424 -805
rect 428 -811 431 -805
rect 435 -811 438 -805
rect 442 -811 445 -805
rect 449 -811 452 -805
rect 456 -811 459 -805
rect 463 -811 466 -805
rect 470 -811 473 -805
rect 477 -811 483 -805
rect 484 -811 487 -805
rect 491 -811 494 -805
rect 498 -811 501 -805
rect 505 -811 508 -805
rect 512 -811 515 -805
rect 519 -811 522 -805
rect 526 -811 529 -805
rect 533 -811 536 -805
rect 540 -811 543 -805
rect 547 -811 553 -805
rect 554 -811 557 -805
rect 561 -811 564 -805
rect 568 -811 571 -805
rect 575 -811 578 -805
rect 582 -811 585 -805
rect 589 -811 592 -805
rect 596 -811 602 -805
rect 603 -811 606 -805
rect 610 -811 613 -805
rect 617 -811 623 -805
rect 624 -811 627 -805
rect 631 -811 634 -805
rect 638 -811 641 -805
rect 645 -811 648 -805
rect 652 -811 655 -805
rect 659 -811 662 -805
rect 666 -811 669 -805
rect 673 -811 676 -805
rect 680 -811 683 -805
rect 687 -811 690 -805
rect 694 -811 697 -805
rect 701 -811 704 -805
rect 708 -811 711 -805
rect 715 -811 718 -805
rect 722 -811 725 -805
rect 729 -811 732 -805
rect 736 -811 739 -805
rect 743 -811 746 -805
rect 750 -811 753 -805
rect 757 -811 760 -805
rect 764 -811 767 -805
rect 771 -811 777 -805
rect 778 -811 781 -805
rect 785 -811 788 -805
rect 1 -866 7 -860
rect 8 -866 11 -860
rect 15 -866 21 -860
rect 22 -866 25 -860
rect 29 -866 32 -860
rect 36 -866 42 -860
rect 43 -866 46 -860
rect 50 -866 56 -860
rect 57 -866 60 -860
rect 64 -866 67 -860
rect 71 -866 74 -860
rect 78 -866 81 -860
rect 85 -866 88 -860
rect 92 -866 95 -860
rect 99 -866 102 -860
rect 106 -866 112 -860
rect 113 -866 119 -860
rect 120 -866 123 -860
rect 127 -866 130 -860
rect 134 -866 140 -860
rect 141 -866 144 -860
rect 148 -866 151 -860
rect 155 -866 158 -860
rect 162 -866 165 -860
rect 169 -866 175 -860
rect 176 -866 179 -860
rect 183 -866 186 -860
rect 190 -866 193 -860
rect 197 -866 200 -860
rect 204 -866 207 -860
rect 211 -866 214 -860
rect 218 -866 221 -860
rect 225 -866 228 -860
rect 232 -866 235 -860
rect 239 -866 242 -860
rect 246 -866 249 -860
rect 253 -866 256 -860
rect 260 -866 266 -860
rect 267 -866 273 -860
rect 274 -866 277 -860
rect 281 -866 284 -860
rect 288 -866 291 -860
rect 295 -866 298 -860
rect 302 -866 305 -860
rect 309 -866 312 -860
rect 316 -866 319 -860
rect 323 -866 326 -860
rect 330 -866 333 -860
rect 337 -866 340 -860
rect 344 -866 350 -860
rect 351 -866 354 -860
rect 358 -866 361 -860
rect 365 -866 371 -860
rect 372 -866 375 -860
rect 379 -866 385 -860
rect 386 -866 392 -860
rect 393 -866 396 -860
rect 400 -866 403 -860
rect 407 -866 410 -860
rect 414 -866 417 -860
rect 421 -866 424 -860
rect 428 -866 431 -860
rect 435 -866 438 -860
rect 442 -866 445 -860
rect 449 -866 452 -860
rect 456 -866 459 -860
rect 463 -866 466 -860
rect 470 -866 473 -860
rect 477 -866 480 -860
rect 484 -866 487 -860
rect 491 -866 494 -860
rect 498 -866 504 -860
rect 505 -866 508 -860
rect 512 -866 515 -860
rect 519 -866 522 -860
rect 526 -866 529 -860
rect 533 -866 536 -860
rect 540 -866 546 -860
rect 547 -866 550 -860
rect 554 -866 557 -860
rect 561 -866 564 -860
rect 568 -866 571 -860
rect 575 -866 578 -860
rect 582 -866 585 -860
rect 589 -866 592 -860
rect 596 -866 599 -860
rect 603 -866 609 -860
rect 610 -866 613 -860
rect 617 -866 620 -860
rect 624 -866 627 -860
rect 631 -866 634 -860
rect 638 -866 641 -860
rect 645 -866 648 -860
rect 652 -866 655 -860
rect 659 -866 662 -860
rect 666 -866 669 -860
rect 680 -866 686 -860
rect 687 -866 690 -860
rect 694 -866 697 -860
rect 701 -866 704 -860
rect 722 -866 728 -860
rect 729 -866 735 -860
rect 736 -866 739 -860
rect 743 -866 746 -860
rect 750 -866 753 -860
rect 757 -866 760 -860
rect 1 -919 7 -913
rect 43 -919 46 -913
rect 50 -919 53 -913
rect 57 -919 60 -913
rect 64 -919 67 -913
rect 71 -919 77 -913
rect 78 -919 81 -913
rect 85 -919 88 -913
rect 92 -919 95 -913
rect 99 -919 102 -913
rect 106 -919 109 -913
rect 113 -919 116 -913
rect 120 -919 126 -913
rect 127 -919 130 -913
rect 134 -919 137 -913
rect 141 -919 144 -913
rect 148 -919 151 -913
rect 155 -919 161 -913
rect 162 -919 165 -913
rect 169 -919 172 -913
rect 176 -919 182 -913
rect 183 -919 186 -913
rect 190 -919 193 -913
rect 197 -919 203 -913
rect 204 -919 210 -913
rect 211 -919 214 -913
rect 218 -919 221 -913
rect 225 -919 228 -913
rect 232 -919 235 -913
rect 239 -919 242 -913
rect 246 -919 249 -913
rect 253 -919 259 -913
rect 260 -919 263 -913
rect 267 -919 273 -913
rect 274 -919 277 -913
rect 281 -919 284 -913
rect 288 -919 291 -913
rect 295 -919 301 -913
rect 302 -919 305 -913
rect 309 -919 312 -913
rect 316 -919 319 -913
rect 323 -919 329 -913
rect 330 -919 333 -913
rect 337 -919 340 -913
rect 344 -919 347 -913
rect 351 -919 354 -913
rect 358 -919 361 -913
rect 365 -919 371 -913
rect 372 -919 378 -913
rect 379 -919 382 -913
rect 386 -919 389 -913
rect 393 -919 399 -913
rect 400 -919 403 -913
rect 407 -919 410 -913
rect 414 -919 417 -913
rect 421 -919 424 -913
rect 428 -919 431 -913
rect 435 -919 438 -913
rect 442 -919 445 -913
rect 449 -919 452 -913
rect 456 -919 459 -913
rect 463 -919 469 -913
rect 470 -919 473 -913
rect 477 -919 480 -913
rect 484 -919 487 -913
rect 491 -919 494 -913
rect 498 -919 501 -913
rect 505 -919 508 -913
rect 512 -919 515 -913
rect 519 -919 525 -913
rect 526 -919 529 -913
rect 533 -919 536 -913
rect 540 -919 543 -913
rect 547 -919 550 -913
rect 554 -919 557 -913
rect 561 -919 564 -913
rect 568 -919 571 -913
rect 575 -919 578 -913
rect 582 -919 585 -913
rect 589 -919 592 -913
rect 596 -919 599 -913
rect 603 -919 606 -913
rect 610 -919 613 -913
rect 617 -919 620 -913
rect 624 -919 627 -913
rect 631 -919 634 -913
rect 638 -919 644 -913
rect 645 -919 648 -913
rect 652 -919 658 -913
rect 659 -919 665 -913
rect 666 -919 669 -913
rect 673 -919 676 -913
rect 680 -919 683 -913
rect 715 -919 718 -913
rect 743 -919 749 -913
rect 1 -978 7 -972
rect 8 -978 14 -972
rect 15 -978 21 -972
rect 64 -978 67 -972
rect 71 -978 74 -972
rect 78 -978 81 -972
rect 85 -978 88 -972
rect 92 -978 98 -972
rect 99 -978 105 -972
rect 106 -978 112 -972
rect 113 -978 119 -972
rect 120 -978 123 -972
rect 127 -978 130 -972
rect 134 -978 137 -972
rect 141 -978 144 -972
rect 148 -978 151 -972
rect 155 -978 158 -972
rect 162 -978 165 -972
rect 169 -978 172 -972
rect 176 -978 179 -972
rect 183 -978 186 -972
rect 190 -978 193 -972
rect 197 -978 203 -972
rect 204 -978 207 -972
rect 211 -978 214 -972
rect 218 -978 221 -972
rect 225 -978 231 -972
rect 232 -978 235 -972
rect 239 -978 242 -972
rect 246 -978 249 -972
rect 253 -978 256 -972
rect 260 -978 263 -972
rect 267 -978 270 -972
rect 274 -978 277 -972
rect 281 -978 284 -972
rect 288 -978 291 -972
rect 295 -978 298 -972
rect 302 -978 305 -972
rect 309 -978 315 -972
rect 316 -978 322 -972
rect 323 -978 326 -972
rect 330 -978 333 -972
rect 337 -978 340 -972
rect 344 -978 347 -972
rect 351 -978 354 -972
rect 358 -978 361 -972
rect 365 -978 371 -972
rect 372 -978 378 -972
rect 379 -978 382 -972
rect 386 -978 392 -972
rect 393 -978 396 -972
rect 400 -978 403 -972
rect 407 -978 410 -972
rect 414 -978 420 -972
rect 421 -978 427 -972
rect 428 -978 431 -972
rect 435 -978 438 -972
rect 442 -978 445 -972
rect 449 -978 455 -972
rect 456 -978 459 -972
rect 463 -978 466 -972
rect 470 -978 473 -972
rect 477 -978 480 -972
rect 484 -978 487 -972
rect 491 -978 494 -972
rect 498 -978 501 -972
rect 505 -978 508 -972
rect 512 -978 515 -972
rect 519 -978 525 -972
rect 526 -978 529 -972
rect 533 -978 536 -972
rect 540 -978 546 -972
rect 547 -978 550 -972
rect 554 -978 557 -972
rect 561 -978 564 -972
rect 568 -978 571 -972
rect 575 -978 578 -972
rect 582 -978 585 -972
rect 589 -978 592 -972
rect 596 -978 599 -972
rect 603 -978 606 -972
rect 610 -978 613 -972
rect 617 -978 620 -972
rect 624 -978 630 -972
rect 659 -978 662 -972
rect 673 -978 676 -972
rect 1 -1017 7 -1011
rect 8 -1017 14 -1011
rect 99 -1017 102 -1011
rect 141 -1017 144 -1011
rect 148 -1017 151 -1011
rect 155 -1017 158 -1011
rect 162 -1017 165 -1011
rect 169 -1017 172 -1011
rect 176 -1017 179 -1011
rect 183 -1017 186 -1011
rect 190 -1017 193 -1011
rect 197 -1017 200 -1011
rect 204 -1017 207 -1011
rect 211 -1017 217 -1011
rect 218 -1017 221 -1011
rect 225 -1017 228 -1011
rect 232 -1017 235 -1011
rect 239 -1017 242 -1011
rect 246 -1017 252 -1011
rect 253 -1017 256 -1011
rect 260 -1017 266 -1011
rect 267 -1017 270 -1011
rect 274 -1017 277 -1011
rect 281 -1017 284 -1011
rect 288 -1017 291 -1011
rect 295 -1017 301 -1011
rect 302 -1017 305 -1011
rect 309 -1017 312 -1011
rect 316 -1017 322 -1011
rect 323 -1017 326 -1011
rect 330 -1017 336 -1011
rect 337 -1017 340 -1011
rect 344 -1017 350 -1011
rect 351 -1017 354 -1011
rect 358 -1017 364 -1011
rect 365 -1017 371 -1011
rect 372 -1017 375 -1011
rect 379 -1017 382 -1011
rect 386 -1017 389 -1011
rect 393 -1017 396 -1011
rect 400 -1017 403 -1011
rect 407 -1017 410 -1011
rect 414 -1017 417 -1011
rect 421 -1017 424 -1011
rect 428 -1017 434 -1011
rect 435 -1017 441 -1011
rect 442 -1017 448 -1011
rect 449 -1017 452 -1011
rect 456 -1017 462 -1011
rect 463 -1017 466 -1011
rect 491 -1017 494 -1011
rect 498 -1017 501 -1011
rect 505 -1017 508 -1011
rect 526 -1017 532 -1011
rect 540 -1017 546 -1011
rect 547 -1017 550 -1011
rect 568 -1017 571 -1011
rect 575 -1017 578 -1011
rect 582 -1017 585 -1011
rect 589 -1017 592 -1011
rect 603 -1017 609 -1011
rect 610 -1017 613 -1011
rect 645 -1017 651 -1011
rect 666 -1017 672 -1011
rect 1 -1046 7 -1040
rect 8 -1046 14 -1040
rect 99 -1046 102 -1040
rect 113 -1046 116 -1040
rect 120 -1046 126 -1040
rect 127 -1046 130 -1040
rect 134 -1046 137 -1040
rect 141 -1046 144 -1040
rect 148 -1046 151 -1040
rect 155 -1046 158 -1040
rect 162 -1046 165 -1040
rect 169 -1046 175 -1040
rect 176 -1046 182 -1040
rect 183 -1046 189 -1040
rect 190 -1046 193 -1040
rect 197 -1046 200 -1040
rect 204 -1046 207 -1040
rect 211 -1046 217 -1040
rect 218 -1046 221 -1040
rect 225 -1046 231 -1040
rect 232 -1046 235 -1040
rect 239 -1046 245 -1040
rect 246 -1046 249 -1040
rect 253 -1046 256 -1040
rect 260 -1046 266 -1040
rect 267 -1046 270 -1040
rect 274 -1046 280 -1040
rect 281 -1046 287 -1040
rect 288 -1046 291 -1040
rect 295 -1046 298 -1040
rect 302 -1046 308 -1040
rect 309 -1046 312 -1040
rect 316 -1046 319 -1040
rect 365 -1046 368 -1040
rect 372 -1046 378 -1040
rect 379 -1046 385 -1040
rect 386 -1046 389 -1040
rect 393 -1046 396 -1040
rect 400 -1046 406 -1040
rect 407 -1046 410 -1040
rect 414 -1046 420 -1040
rect 421 -1046 424 -1040
rect 428 -1046 431 -1040
rect 435 -1046 438 -1040
rect 442 -1046 445 -1040
rect 456 -1046 459 -1040
rect 470 -1046 476 -1040
rect 477 -1046 480 -1040
rect 484 -1046 487 -1040
rect 540 -1046 546 -1040
rect 547 -1046 550 -1040
rect 561 -1046 564 -1040
rect 568 -1046 571 -1040
rect 575 -1046 581 -1040
rect 582 -1046 585 -1040
rect 589 -1046 592 -1040
rect 1 -1067 7 -1061
rect 8 -1067 14 -1061
rect 99 -1067 105 -1061
rect 106 -1067 109 -1061
rect 134 -1067 140 -1061
rect 141 -1067 147 -1061
rect 148 -1067 151 -1061
rect 155 -1067 161 -1061
rect 162 -1067 165 -1061
rect 169 -1067 175 -1061
rect 190 -1067 196 -1061
rect 197 -1067 200 -1061
rect 204 -1067 210 -1061
rect 211 -1067 217 -1061
rect 218 -1067 224 -1061
rect 225 -1067 228 -1061
rect 232 -1067 235 -1061
rect 281 -1067 287 -1061
rect 295 -1067 301 -1061
rect 379 -1067 382 -1061
rect 393 -1067 399 -1061
rect 407 -1067 413 -1061
rect 428 -1067 431 -1061
rect 435 -1067 441 -1061
rect 442 -1067 448 -1061
rect 449 -1067 455 -1061
rect 456 -1067 459 -1061
rect 561 -1067 567 -1061
rect 575 -1067 581 -1061
rect 582 -1067 585 -1061
<< polysilicon >>
rect 114 -7 115 -5
rect 121 -7 122 -5
rect 121 -13 122 -11
rect 128 -7 129 -5
rect 131 -7 132 -5
rect 135 -7 136 -5
rect 135 -13 136 -11
rect 142 -7 143 -5
rect 149 -7 150 -5
rect 156 -7 157 -5
rect 156 -13 157 -11
rect 163 -7 164 -5
rect 166 -7 167 -5
rect 173 -13 174 -11
rect 177 -7 178 -5
rect 177 -13 178 -11
rect 184 -13 185 -11
rect 187 -13 188 -11
rect 191 -7 192 -5
rect 191 -13 192 -11
rect 198 -7 199 -5
rect 201 -13 202 -11
rect 208 -7 209 -5
rect 215 -13 216 -11
rect 236 -7 237 -5
rect 236 -13 237 -11
rect 247 -7 248 -5
rect 247 -13 248 -11
rect 296 -7 297 -5
rect 296 -13 297 -11
rect 313 -7 314 -5
rect 313 -13 314 -11
rect 317 -7 318 -5
rect 317 -13 318 -11
rect 331 -7 332 -5
rect 331 -13 332 -11
rect 338 -7 339 -5
rect 348 -7 349 -5
rect 352 -7 353 -5
rect 352 -13 353 -11
rect 373 -7 374 -5
rect 373 -13 374 -11
rect 422 -13 423 -11
rect 65 -32 66 -30
rect 72 -26 73 -24
rect 72 -32 73 -30
rect 79 -26 80 -24
rect 79 -32 80 -30
rect 89 -26 90 -24
rect 96 -26 97 -24
rect 96 -32 97 -30
rect 100 -26 101 -24
rect 100 -32 101 -30
rect 107 -26 108 -24
rect 107 -32 108 -30
rect 117 -26 118 -24
rect 117 -32 118 -30
rect 121 -32 122 -30
rect 128 -26 129 -24
rect 131 -26 132 -24
rect 135 -26 136 -24
rect 135 -32 136 -30
rect 142 -26 143 -24
rect 142 -32 143 -30
rect 149 -26 150 -24
rect 149 -32 150 -30
rect 156 -26 157 -24
rect 159 -26 160 -24
rect 159 -32 160 -30
rect 166 -32 167 -30
rect 170 -26 171 -24
rect 170 -32 171 -30
rect 177 -26 178 -24
rect 177 -32 178 -30
rect 184 -26 185 -24
rect 184 -32 185 -30
rect 191 -26 192 -24
rect 191 -32 192 -30
rect 198 -26 199 -24
rect 205 -32 206 -30
rect 212 -26 213 -24
rect 212 -32 213 -30
rect 219 -26 220 -24
rect 222 -32 223 -30
rect 229 -26 230 -24
rect 226 -32 227 -30
rect 233 -26 234 -24
rect 233 -32 234 -30
rect 240 -26 241 -24
rect 240 -32 241 -30
rect 250 -32 251 -30
rect 254 -26 255 -24
rect 254 -32 255 -30
rect 261 -32 262 -30
rect 264 -32 265 -30
rect 282 -26 283 -24
rect 282 -32 283 -30
rect 296 -26 297 -24
rect 296 -32 297 -30
rect 303 -26 304 -24
rect 303 -32 304 -30
rect 313 -32 314 -30
rect 327 -32 328 -30
rect 331 -26 332 -24
rect 331 -32 332 -30
rect 345 -26 346 -24
rect 345 -32 346 -30
rect 352 -26 353 -24
rect 352 -32 353 -30
rect 394 -26 395 -24
rect 394 -32 395 -30
rect 404 -26 405 -24
rect 429 -26 430 -24
rect 429 -32 430 -30
rect 436 -26 437 -24
rect 436 -32 437 -30
rect 485 -26 486 -24
rect 488 -32 489 -30
rect 555 -26 556 -24
rect 555 -32 556 -30
rect 51 -55 52 -53
rect 51 -61 52 -59
rect 58 -55 59 -53
rect 65 -55 66 -53
rect 65 -61 66 -59
rect 72 -55 73 -53
rect 72 -61 73 -59
rect 82 -61 83 -59
rect 86 -55 87 -53
rect 86 -61 87 -59
rect 93 -55 94 -53
rect 93 -61 94 -59
rect 100 -55 101 -53
rect 100 -61 101 -59
rect 107 -55 108 -53
rect 107 -61 108 -59
rect 114 -55 115 -53
rect 114 -61 115 -59
rect 121 -55 122 -53
rect 121 -61 122 -59
rect 128 -61 129 -59
rect 131 -61 132 -59
rect 135 -55 136 -53
rect 135 -61 136 -59
rect 142 -55 143 -53
rect 142 -61 143 -59
rect 149 -55 150 -53
rect 149 -61 150 -59
rect 156 -55 157 -53
rect 159 -55 160 -53
rect 163 -55 164 -53
rect 163 -61 164 -59
rect 170 -55 171 -53
rect 170 -61 171 -59
rect 177 -55 178 -53
rect 177 -61 178 -59
rect 184 -55 185 -53
rect 184 -61 185 -59
rect 194 -55 195 -53
rect 191 -61 192 -59
rect 198 -55 199 -53
rect 198 -61 199 -59
rect 205 -55 206 -53
rect 205 -61 206 -59
rect 215 -55 216 -53
rect 215 -61 216 -59
rect 219 -55 220 -53
rect 219 -61 220 -59
rect 226 -55 227 -53
rect 229 -61 230 -59
rect 233 -55 234 -53
rect 233 -61 234 -59
rect 240 -61 241 -59
rect 243 -61 244 -59
rect 247 -55 248 -53
rect 247 -61 248 -59
rect 254 -55 255 -53
rect 254 -61 255 -59
rect 261 -55 262 -53
rect 261 -61 262 -59
rect 268 -55 269 -53
rect 268 -61 269 -59
rect 275 -55 276 -53
rect 275 -61 276 -59
rect 285 -55 286 -53
rect 285 -61 286 -59
rect 289 -55 290 -53
rect 289 -61 290 -59
rect 296 -55 297 -53
rect 296 -61 297 -59
rect 303 -55 304 -53
rect 313 -61 314 -59
rect 317 -55 318 -53
rect 324 -55 325 -53
rect 324 -61 325 -59
rect 331 -55 332 -53
rect 331 -61 332 -59
rect 338 -55 339 -53
rect 338 -61 339 -59
rect 345 -55 346 -53
rect 345 -61 346 -59
rect 352 -55 353 -53
rect 352 -61 353 -59
rect 359 -55 360 -53
rect 359 -61 360 -59
rect 366 -55 367 -53
rect 366 -61 367 -59
rect 373 -55 374 -53
rect 373 -61 374 -59
rect 380 -55 381 -53
rect 387 -55 388 -53
rect 387 -61 388 -59
rect 394 -55 395 -53
rect 394 -61 395 -59
rect 404 -55 405 -53
rect 401 -61 402 -59
rect 415 -55 416 -53
rect 415 -61 416 -59
rect 443 -55 444 -53
rect 443 -61 444 -59
rect 450 -55 451 -53
rect 450 -61 451 -59
rect 457 -61 458 -59
rect 576 -55 577 -53
rect 576 -61 577 -59
rect 30 -94 31 -92
rect 30 -100 31 -98
rect 37 -94 38 -92
rect 37 -100 38 -98
rect 44 -94 45 -92
rect 44 -100 45 -98
rect 51 -94 52 -92
rect 51 -100 52 -98
rect 58 -94 59 -92
rect 58 -100 59 -98
rect 65 -94 66 -92
rect 68 -100 69 -98
rect 72 -94 73 -92
rect 72 -100 73 -98
rect 79 -94 80 -92
rect 79 -100 80 -98
rect 86 -94 87 -92
rect 86 -100 87 -98
rect 96 -94 97 -92
rect 96 -100 97 -98
rect 100 -94 101 -92
rect 100 -100 101 -98
rect 107 -94 108 -92
rect 107 -100 108 -98
rect 114 -94 115 -92
rect 114 -100 115 -98
rect 121 -100 122 -98
rect 124 -100 125 -98
rect 128 -94 129 -92
rect 131 -94 132 -92
rect 135 -94 136 -92
rect 135 -100 136 -98
rect 142 -94 143 -92
rect 142 -100 143 -98
rect 152 -94 153 -92
rect 149 -100 150 -98
rect 156 -94 157 -92
rect 156 -100 157 -98
rect 159 -100 160 -98
rect 163 -94 164 -92
rect 163 -100 164 -98
rect 170 -94 171 -92
rect 170 -100 171 -98
rect 177 -94 178 -92
rect 177 -100 178 -98
rect 184 -94 185 -92
rect 184 -100 185 -98
rect 191 -94 192 -92
rect 191 -100 192 -98
rect 198 -94 199 -92
rect 198 -100 199 -98
rect 205 -94 206 -92
rect 205 -100 206 -98
rect 212 -94 213 -92
rect 212 -100 213 -98
rect 219 -94 220 -92
rect 219 -100 220 -98
rect 226 -94 227 -92
rect 226 -100 227 -98
rect 233 -94 234 -92
rect 233 -100 234 -98
rect 240 -94 241 -92
rect 240 -100 241 -98
rect 243 -100 244 -98
rect 247 -94 248 -92
rect 247 -100 248 -98
rect 257 -100 258 -98
rect 261 -94 262 -92
rect 261 -100 262 -98
rect 268 -94 269 -92
rect 268 -100 269 -98
rect 275 -94 276 -92
rect 275 -100 276 -98
rect 282 -100 283 -98
rect 289 -94 290 -92
rect 289 -100 290 -98
rect 296 -94 297 -92
rect 296 -100 297 -98
rect 303 -94 304 -92
rect 303 -100 304 -98
rect 313 -94 314 -92
rect 313 -100 314 -98
rect 320 -100 321 -98
rect 324 -94 325 -92
rect 324 -100 325 -98
rect 331 -94 332 -92
rect 331 -100 332 -98
rect 338 -94 339 -92
rect 338 -100 339 -98
rect 345 -94 346 -92
rect 345 -100 346 -98
rect 355 -100 356 -98
rect 359 -94 360 -92
rect 359 -100 360 -98
rect 369 -94 370 -92
rect 366 -100 367 -98
rect 373 -94 374 -92
rect 373 -100 374 -98
rect 380 -94 381 -92
rect 380 -100 381 -98
rect 387 -94 388 -92
rect 387 -100 388 -98
rect 394 -94 395 -92
rect 394 -100 395 -98
rect 401 -94 402 -92
rect 401 -100 402 -98
rect 408 -94 409 -92
rect 408 -100 409 -98
rect 415 -94 416 -92
rect 415 -100 416 -98
rect 425 -94 426 -92
rect 429 -94 430 -92
rect 429 -100 430 -98
rect 436 -94 437 -92
rect 436 -100 437 -98
rect 443 -100 444 -98
rect 446 -100 447 -98
rect 450 -94 451 -92
rect 450 -100 451 -98
rect 457 -94 458 -92
rect 460 -100 461 -98
rect 464 -94 465 -92
rect 464 -100 465 -98
rect 471 -94 472 -92
rect 471 -100 472 -98
rect 478 -94 479 -92
rect 478 -100 479 -98
rect 492 -94 493 -92
rect 492 -100 493 -98
rect 523 -100 524 -98
rect 527 -94 528 -92
rect 530 -94 531 -92
rect 576 -94 577 -92
rect 576 -100 577 -98
rect 590 -94 591 -92
rect 590 -100 591 -98
rect 9 -145 10 -143
rect 9 -151 10 -149
rect 16 -145 17 -143
rect 16 -151 17 -149
rect 26 -145 27 -143
rect 30 -145 31 -143
rect 30 -151 31 -149
rect 37 -145 38 -143
rect 37 -151 38 -149
rect 44 -145 45 -143
rect 44 -151 45 -149
rect 51 -145 52 -143
rect 51 -151 52 -149
rect 58 -145 59 -143
rect 58 -151 59 -149
rect 65 -145 66 -143
rect 65 -151 66 -149
rect 72 -145 73 -143
rect 75 -145 76 -143
rect 72 -151 73 -149
rect 79 -151 80 -149
rect 82 -151 83 -149
rect 86 -145 87 -143
rect 86 -151 87 -149
rect 93 -145 94 -143
rect 96 -151 97 -149
rect 100 -145 101 -143
rect 100 -151 101 -149
rect 107 -145 108 -143
rect 107 -151 108 -149
rect 114 -145 115 -143
rect 114 -151 115 -149
rect 121 -145 122 -143
rect 121 -151 122 -149
rect 128 -145 129 -143
rect 128 -151 129 -149
rect 135 -145 136 -143
rect 135 -151 136 -149
rect 142 -145 143 -143
rect 142 -151 143 -149
rect 149 -145 150 -143
rect 149 -151 150 -149
rect 156 -145 157 -143
rect 156 -151 157 -149
rect 166 -145 167 -143
rect 170 -145 171 -143
rect 173 -145 174 -143
rect 170 -151 171 -149
rect 173 -151 174 -149
rect 177 -145 178 -143
rect 177 -151 178 -149
rect 184 -145 185 -143
rect 184 -151 185 -149
rect 191 -145 192 -143
rect 191 -151 192 -149
rect 198 -145 199 -143
rect 198 -151 199 -149
rect 205 -145 206 -143
rect 205 -151 206 -149
rect 212 -145 213 -143
rect 212 -151 213 -149
rect 219 -145 220 -143
rect 222 -145 223 -143
rect 219 -151 220 -149
rect 222 -151 223 -149
rect 226 -145 227 -143
rect 226 -151 227 -149
rect 233 -145 234 -143
rect 233 -151 234 -149
rect 240 -145 241 -143
rect 240 -151 241 -149
rect 247 -145 248 -143
rect 247 -151 248 -149
rect 257 -145 258 -143
rect 257 -151 258 -149
rect 261 -145 262 -143
rect 261 -151 262 -149
rect 268 -145 269 -143
rect 268 -151 269 -149
rect 275 -145 276 -143
rect 278 -151 279 -149
rect 282 -145 283 -143
rect 282 -151 283 -149
rect 289 -145 290 -143
rect 292 -151 293 -149
rect 296 -145 297 -143
rect 296 -151 297 -149
rect 303 -145 304 -143
rect 303 -151 304 -149
rect 310 -145 311 -143
rect 313 -145 314 -143
rect 313 -151 314 -149
rect 320 -145 321 -143
rect 317 -151 318 -149
rect 320 -151 321 -149
rect 324 -145 325 -143
rect 324 -151 325 -149
rect 331 -145 332 -143
rect 331 -151 332 -149
rect 338 -145 339 -143
rect 338 -151 339 -149
rect 345 -145 346 -143
rect 345 -151 346 -149
rect 352 -145 353 -143
rect 352 -151 353 -149
rect 359 -145 360 -143
rect 359 -151 360 -149
rect 366 -145 367 -143
rect 366 -151 367 -149
rect 373 -145 374 -143
rect 373 -151 374 -149
rect 380 -145 381 -143
rect 380 -151 381 -149
rect 387 -145 388 -143
rect 387 -151 388 -149
rect 394 -145 395 -143
rect 394 -151 395 -149
rect 401 -145 402 -143
rect 401 -151 402 -149
rect 408 -145 409 -143
rect 408 -151 409 -149
rect 415 -145 416 -143
rect 415 -151 416 -149
rect 418 -151 419 -149
rect 422 -145 423 -143
rect 422 -151 423 -149
rect 429 -145 430 -143
rect 429 -151 430 -149
rect 436 -145 437 -143
rect 436 -151 437 -149
rect 443 -145 444 -143
rect 443 -151 444 -149
rect 450 -145 451 -143
rect 450 -151 451 -149
rect 457 -145 458 -143
rect 457 -151 458 -149
rect 464 -145 465 -143
rect 464 -151 465 -149
rect 474 -145 475 -143
rect 471 -151 472 -149
rect 478 -145 479 -143
rect 478 -151 479 -149
rect 485 -145 486 -143
rect 485 -151 486 -149
rect 492 -145 493 -143
rect 492 -151 493 -149
rect 499 -145 500 -143
rect 506 -145 507 -143
rect 506 -151 507 -149
rect 513 -145 514 -143
rect 513 -151 514 -149
rect 520 -145 521 -143
rect 520 -151 521 -149
rect 527 -145 528 -143
rect 527 -151 528 -149
rect 534 -145 535 -143
rect 534 -151 535 -149
rect 541 -145 542 -143
rect 541 -151 542 -149
rect 548 -145 549 -143
rect 548 -151 549 -149
rect 555 -145 556 -143
rect 555 -151 556 -149
rect 562 -145 563 -143
rect 562 -151 563 -149
rect 569 -145 570 -143
rect 569 -151 570 -149
rect 576 -145 577 -143
rect 576 -151 577 -149
rect 586 -145 587 -143
rect 583 -151 584 -149
rect 586 -151 587 -149
rect 590 -145 591 -143
rect 590 -151 591 -149
rect 597 -145 598 -143
rect 597 -151 598 -149
rect 604 -145 605 -143
rect 604 -151 605 -149
rect 611 -145 612 -143
rect 611 -151 612 -149
rect 618 -145 619 -143
rect 618 -151 619 -149
rect 625 -151 626 -149
rect 628 -151 629 -149
rect 16 -206 17 -204
rect 16 -212 17 -210
rect 23 -206 24 -204
rect 23 -212 24 -210
rect 30 -206 31 -204
rect 30 -212 31 -210
rect 37 -206 38 -204
rect 37 -212 38 -210
rect 44 -206 45 -204
rect 44 -212 45 -210
rect 51 -206 52 -204
rect 51 -212 52 -210
rect 58 -206 59 -204
rect 58 -212 59 -210
rect 65 -206 66 -204
rect 65 -212 66 -210
rect 75 -212 76 -210
rect 79 -206 80 -204
rect 79 -212 80 -210
rect 86 -206 87 -204
rect 86 -212 87 -210
rect 93 -206 94 -204
rect 96 -206 97 -204
rect 96 -212 97 -210
rect 100 -206 101 -204
rect 107 -206 108 -204
rect 107 -212 108 -210
rect 114 -206 115 -204
rect 114 -212 115 -210
rect 121 -206 122 -204
rect 121 -212 122 -210
rect 128 -206 129 -204
rect 128 -212 129 -210
rect 135 -206 136 -204
rect 138 -206 139 -204
rect 135 -212 136 -210
rect 142 -206 143 -204
rect 142 -212 143 -210
rect 149 -206 150 -204
rect 149 -212 150 -210
rect 156 -206 157 -204
rect 156 -212 157 -210
rect 163 -206 164 -204
rect 163 -212 164 -210
rect 170 -206 171 -204
rect 170 -212 171 -210
rect 177 -206 178 -204
rect 180 -206 181 -204
rect 177 -212 178 -210
rect 180 -212 181 -210
rect 184 -206 185 -204
rect 184 -212 185 -210
rect 191 -206 192 -204
rect 191 -212 192 -210
rect 198 -206 199 -204
rect 198 -212 199 -210
rect 208 -206 209 -204
rect 212 -206 213 -204
rect 215 -206 216 -204
rect 219 -206 220 -204
rect 219 -212 220 -210
rect 226 -206 227 -204
rect 226 -212 227 -210
rect 233 -206 234 -204
rect 233 -212 234 -210
rect 240 -206 241 -204
rect 240 -212 241 -210
rect 247 -206 248 -204
rect 247 -212 248 -210
rect 254 -206 255 -204
rect 254 -212 255 -210
rect 261 -206 262 -204
rect 261 -212 262 -210
rect 268 -206 269 -204
rect 268 -212 269 -210
rect 278 -206 279 -204
rect 275 -212 276 -210
rect 278 -212 279 -210
rect 282 -206 283 -204
rect 282 -212 283 -210
rect 289 -206 290 -204
rect 289 -212 290 -210
rect 296 -206 297 -204
rect 299 -206 300 -204
rect 299 -212 300 -210
rect 306 -206 307 -204
rect 310 -206 311 -204
rect 310 -212 311 -210
rect 317 -206 318 -204
rect 317 -212 318 -210
rect 327 -212 328 -210
rect 331 -206 332 -204
rect 334 -206 335 -204
rect 331 -212 332 -210
rect 341 -206 342 -204
rect 341 -212 342 -210
rect 345 -206 346 -204
rect 345 -212 346 -210
rect 352 -206 353 -204
rect 352 -212 353 -210
rect 359 -206 360 -204
rect 359 -212 360 -210
rect 369 -206 370 -204
rect 366 -212 367 -210
rect 369 -212 370 -210
rect 373 -206 374 -204
rect 373 -212 374 -210
rect 380 -206 381 -204
rect 380 -212 381 -210
rect 387 -206 388 -204
rect 390 -206 391 -204
rect 387 -212 388 -210
rect 394 -206 395 -204
rect 394 -212 395 -210
rect 401 -206 402 -204
rect 401 -212 402 -210
rect 408 -206 409 -204
rect 408 -212 409 -210
rect 415 -206 416 -204
rect 415 -212 416 -210
rect 422 -206 423 -204
rect 422 -212 423 -210
rect 429 -206 430 -204
rect 429 -212 430 -210
rect 436 -206 437 -204
rect 436 -212 437 -210
rect 443 -212 444 -210
rect 446 -212 447 -210
rect 450 -206 451 -204
rect 450 -212 451 -210
rect 457 -206 458 -204
rect 457 -212 458 -210
rect 464 -206 465 -204
rect 464 -212 465 -210
rect 471 -206 472 -204
rect 471 -212 472 -210
rect 478 -206 479 -204
rect 478 -212 479 -210
rect 488 -206 489 -204
rect 488 -212 489 -210
rect 492 -206 493 -204
rect 492 -212 493 -210
rect 499 -206 500 -204
rect 499 -212 500 -210
rect 506 -206 507 -204
rect 506 -212 507 -210
rect 513 -206 514 -204
rect 513 -212 514 -210
rect 520 -206 521 -204
rect 520 -212 521 -210
rect 527 -206 528 -204
rect 527 -212 528 -210
rect 534 -206 535 -204
rect 534 -212 535 -210
rect 541 -206 542 -204
rect 541 -212 542 -210
rect 548 -206 549 -204
rect 548 -212 549 -210
rect 555 -206 556 -204
rect 555 -212 556 -210
rect 562 -206 563 -204
rect 562 -212 563 -210
rect 569 -206 570 -204
rect 569 -212 570 -210
rect 576 -206 577 -204
rect 576 -212 577 -210
rect 583 -206 584 -204
rect 583 -212 584 -210
rect 590 -206 591 -204
rect 590 -212 591 -210
rect 597 -206 598 -204
rect 597 -212 598 -210
rect 604 -206 605 -204
rect 604 -212 605 -210
rect 611 -206 612 -204
rect 611 -212 612 -210
rect 618 -206 619 -204
rect 618 -212 619 -210
rect 625 -206 626 -204
rect 625 -212 626 -210
rect 632 -206 633 -204
rect 632 -212 633 -210
rect 639 -206 640 -204
rect 639 -212 640 -210
rect 646 -206 647 -204
rect 646 -212 647 -210
rect 653 -206 654 -204
rect 653 -212 654 -210
rect 660 -206 661 -204
rect 660 -212 661 -210
rect 667 -206 668 -204
rect 667 -212 668 -210
rect 674 -206 675 -204
rect 674 -212 675 -210
rect 2 -271 3 -269
rect 2 -277 3 -275
rect 9 -271 10 -269
rect 16 -271 17 -269
rect 16 -277 17 -275
rect 23 -271 24 -269
rect 23 -277 24 -275
rect 30 -271 31 -269
rect 33 -271 34 -269
rect 33 -277 34 -275
rect 37 -271 38 -269
rect 37 -277 38 -275
rect 44 -271 45 -269
rect 44 -277 45 -275
rect 51 -271 52 -269
rect 54 -271 55 -269
rect 51 -277 52 -275
rect 54 -277 55 -275
rect 58 -271 59 -269
rect 58 -277 59 -275
rect 65 -271 66 -269
rect 65 -277 66 -275
rect 72 -271 73 -269
rect 72 -277 73 -275
rect 79 -271 80 -269
rect 82 -271 83 -269
rect 82 -277 83 -275
rect 86 -271 87 -269
rect 86 -277 87 -275
rect 93 -271 94 -269
rect 93 -277 94 -275
rect 100 -271 101 -269
rect 103 -271 104 -269
rect 107 -271 108 -269
rect 107 -277 108 -275
rect 110 -277 111 -275
rect 117 -271 118 -269
rect 114 -277 115 -275
rect 121 -271 122 -269
rect 121 -277 122 -275
rect 128 -271 129 -269
rect 128 -277 129 -275
rect 135 -271 136 -269
rect 135 -277 136 -275
rect 142 -271 143 -269
rect 142 -277 143 -275
rect 152 -271 153 -269
rect 156 -271 157 -269
rect 156 -277 157 -275
rect 163 -271 164 -269
rect 163 -277 164 -275
rect 170 -271 171 -269
rect 170 -277 171 -275
rect 177 -271 178 -269
rect 177 -277 178 -275
rect 184 -271 185 -269
rect 184 -277 185 -275
rect 191 -271 192 -269
rect 191 -277 192 -275
rect 198 -271 199 -269
rect 198 -277 199 -275
rect 205 -271 206 -269
rect 205 -277 206 -275
rect 212 -271 213 -269
rect 212 -277 213 -275
rect 219 -271 220 -269
rect 219 -277 220 -275
rect 226 -271 227 -269
rect 226 -277 227 -275
rect 233 -271 234 -269
rect 233 -277 234 -275
rect 243 -271 244 -269
rect 240 -277 241 -275
rect 247 -271 248 -269
rect 250 -271 251 -269
rect 247 -277 248 -275
rect 250 -277 251 -275
rect 254 -271 255 -269
rect 254 -277 255 -275
rect 264 -271 265 -269
rect 261 -277 262 -275
rect 264 -277 265 -275
rect 268 -271 269 -269
rect 268 -277 269 -275
rect 278 -271 279 -269
rect 275 -277 276 -275
rect 278 -277 279 -275
rect 282 -271 283 -269
rect 282 -277 283 -275
rect 289 -271 290 -269
rect 292 -271 293 -269
rect 292 -277 293 -275
rect 296 -271 297 -269
rect 299 -271 300 -269
rect 296 -277 297 -275
rect 299 -277 300 -275
rect 303 -271 304 -269
rect 303 -277 304 -275
rect 310 -271 311 -269
rect 313 -271 314 -269
rect 310 -277 311 -275
rect 313 -277 314 -275
rect 317 -271 318 -269
rect 317 -277 318 -275
rect 324 -271 325 -269
rect 324 -277 325 -275
rect 331 -271 332 -269
rect 331 -277 332 -275
rect 338 -271 339 -269
rect 338 -277 339 -275
rect 345 -271 346 -269
rect 345 -277 346 -275
rect 352 -271 353 -269
rect 352 -277 353 -275
rect 359 -271 360 -269
rect 359 -277 360 -275
rect 369 -271 370 -269
rect 369 -277 370 -275
rect 373 -271 374 -269
rect 373 -277 374 -275
rect 380 -271 381 -269
rect 383 -271 384 -269
rect 380 -277 381 -275
rect 383 -277 384 -275
rect 387 -271 388 -269
rect 387 -277 388 -275
rect 394 -271 395 -269
rect 394 -277 395 -275
rect 401 -271 402 -269
rect 401 -277 402 -275
rect 408 -271 409 -269
rect 408 -277 409 -275
rect 415 -271 416 -269
rect 415 -277 416 -275
rect 422 -271 423 -269
rect 422 -277 423 -275
rect 429 -271 430 -269
rect 429 -277 430 -275
rect 436 -271 437 -269
rect 436 -277 437 -275
rect 443 -271 444 -269
rect 443 -277 444 -275
rect 450 -271 451 -269
rect 450 -277 451 -275
rect 457 -271 458 -269
rect 457 -277 458 -275
rect 467 -277 468 -275
rect 471 -271 472 -269
rect 471 -277 472 -275
rect 478 -271 479 -269
rect 478 -277 479 -275
rect 485 -271 486 -269
rect 485 -277 486 -275
rect 492 -271 493 -269
rect 492 -277 493 -275
rect 499 -271 500 -269
rect 499 -277 500 -275
rect 506 -271 507 -269
rect 506 -277 507 -275
rect 513 -271 514 -269
rect 513 -277 514 -275
rect 520 -271 521 -269
rect 520 -277 521 -275
rect 527 -271 528 -269
rect 527 -277 528 -275
rect 534 -271 535 -269
rect 534 -277 535 -275
rect 541 -271 542 -269
rect 541 -277 542 -275
rect 548 -271 549 -269
rect 548 -277 549 -275
rect 555 -271 556 -269
rect 555 -277 556 -275
rect 562 -271 563 -269
rect 562 -277 563 -275
rect 569 -271 570 -269
rect 569 -277 570 -275
rect 576 -271 577 -269
rect 576 -277 577 -275
rect 583 -271 584 -269
rect 583 -277 584 -275
rect 590 -271 591 -269
rect 590 -277 591 -275
rect 597 -271 598 -269
rect 597 -277 598 -275
rect 604 -271 605 -269
rect 604 -277 605 -275
rect 611 -271 612 -269
rect 611 -277 612 -275
rect 618 -271 619 -269
rect 618 -277 619 -275
rect 625 -271 626 -269
rect 625 -277 626 -275
rect 632 -271 633 -269
rect 632 -277 633 -275
rect 639 -271 640 -269
rect 639 -277 640 -275
rect 646 -271 647 -269
rect 646 -277 647 -275
rect 653 -271 654 -269
rect 653 -277 654 -275
rect 660 -271 661 -269
rect 660 -277 661 -275
rect 667 -271 668 -269
rect 667 -277 668 -275
rect 674 -271 675 -269
rect 674 -277 675 -275
rect 681 -271 682 -269
rect 681 -277 682 -275
rect 688 -271 689 -269
rect 688 -277 689 -275
rect 695 -271 696 -269
rect 695 -277 696 -275
rect 702 -271 703 -269
rect 702 -277 703 -275
rect 712 -271 713 -269
rect 709 -277 710 -275
rect 716 -271 717 -269
rect 716 -277 717 -275
rect 723 -271 724 -269
rect 723 -277 724 -275
rect 730 -271 731 -269
rect 16 -338 17 -336
rect 16 -344 17 -342
rect 26 -338 27 -336
rect 26 -344 27 -342
rect 30 -338 31 -336
rect 30 -344 31 -342
rect 37 -338 38 -336
rect 37 -344 38 -342
rect 44 -338 45 -336
rect 47 -338 48 -336
rect 47 -344 48 -342
rect 51 -338 52 -336
rect 54 -338 55 -336
rect 54 -344 55 -342
rect 58 -338 59 -336
rect 58 -344 59 -342
rect 61 -344 62 -342
rect 65 -338 66 -336
rect 65 -344 66 -342
rect 72 -338 73 -336
rect 72 -344 73 -342
rect 79 -338 80 -336
rect 79 -344 80 -342
rect 86 -338 87 -336
rect 86 -344 87 -342
rect 93 -338 94 -336
rect 93 -344 94 -342
rect 100 -338 101 -336
rect 100 -344 101 -342
rect 110 -338 111 -336
rect 110 -344 111 -342
rect 114 -338 115 -336
rect 114 -344 115 -342
rect 121 -338 122 -336
rect 121 -344 122 -342
rect 128 -338 129 -336
rect 128 -344 129 -342
rect 135 -338 136 -336
rect 135 -344 136 -342
rect 142 -338 143 -336
rect 142 -344 143 -342
rect 149 -338 150 -336
rect 149 -344 150 -342
rect 156 -338 157 -336
rect 156 -344 157 -342
rect 163 -344 164 -342
rect 170 -338 171 -336
rect 170 -344 171 -342
rect 177 -338 178 -336
rect 177 -344 178 -342
rect 184 -338 185 -336
rect 187 -338 188 -336
rect 187 -344 188 -342
rect 191 -338 192 -336
rect 191 -344 192 -342
rect 198 -338 199 -336
rect 198 -344 199 -342
rect 205 -338 206 -336
rect 205 -344 206 -342
rect 212 -338 213 -336
rect 212 -344 213 -342
rect 219 -338 220 -336
rect 219 -344 220 -342
rect 226 -338 227 -336
rect 226 -344 227 -342
rect 229 -344 230 -342
rect 233 -338 234 -336
rect 233 -344 234 -342
rect 240 -338 241 -336
rect 240 -344 241 -342
rect 247 -338 248 -336
rect 247 -344 248 -342
rect 257 -338 258 -336
rect 254 -344 255 -342
rect 261 -338 262 -336
rect 261 -344 262 -342
rect 268 -338 269 -336
rect 268 -344 269 -342
rect 275 -338 276 -336
rect 278 -338 279 -336
rect 278 -344 279 -342
rect 282 -338 283 -336
rect 282 -344 283 -342
rect 285 -344 286 -342
rect 289 -338 290 -336
rect 289 -344 290 -342
rect 299 -338 300 -336
rect 296 -344 297 -342
rect 299 -344 300 -342
rect 303 -338 304 -336
rect 303 -344 304 -342
rect 310 -338 311 -336
rect 310 -344 311 -342
rect 317 -338 318 -336
rect 317 -344 318 -342
rect 324 -338 325 -336
rect 327 -338 328 -336
rect 331 -338 332 -336
rect 331 -344 332 -342
rect 338 -338 339 -336
rect 338 -344 339 -342
rect 345 -338 346 -336
rect 348 -338 349 -336
rect 345 -344 346 -342
rect 348 -344 349 -342
rect 352 -338 353 -336
rect 352 -344 353 -342
rect 362 -338 363 -336
rect 366 -344 367 -342
rect 369 -344 370 -342
rect 373 -338 374 -336
rect 373 -344 374 -342
rect 380 -338 381 -336
rect 380 -344 381 -342
rect 387 -338 388 -336
rect 387 -344 388 -342
rect 394 -338 395 -336
rect 394 -344 395 -342
rect 401 -338 402 -336
rect 401 -344 402 -342
rect 408 -338 409 -336
rect 408 -344 409 -342
rect 415 -338 416 -336
rect 415 -344 416 -342
rect 422 -338 423 -336
rect 422 -344 423 -342
rect 429 -338 430 -336
rect 432 -338 433 -336
rect 429 -344 430 -342
rect 436 -338 437 -336
rect 436 -344 437 -342
rect 443 -338 444 -336
rect 443 -344 444 -342
rect 450 -338 451 -336
rect 450 -344 451 -342
rect 457 -338 458 -336
rect 457 -344 458 -342
rect 464 -338 465 -336
rect 464 -344 465 -342
rect 471 -338 472 -336
rect 471 -344 472 -342
rect 478 -338 479 -336
rect 478 -344 479 -342
rect 485 -338 486 -336
rect 485 -344 486 -342
rect 492 -338 493 -336
rect 492 -344 493 -342
rect 499 -338 500 -336
rect 499 -344 500 -342
rect 506 -338 507 -336
rect 506 -344 507 -342
rect 513 -338 514 -336
rect 513 -344 514 -342
rect 520 -338 521 -336
rect 520 -344 521 -342
rect 527 -338 528 -336
rect 527 -344 528 -342
rect 534 -338 535 -336
rect 534 -344 535 -342
rect 541 -338 542 -336
rect 541 -344 542 -342
rect 548 -338 549 -336
rect 548 -344 549 -342
rect 555 -338 556 -336
rect 555 -344 556 -342
rect 562 -338 563 -336
rect 562 -344 563 -342
rect 569 -338 570 -336
rect 569 -344 570 -342
rect 576 -338 577 -336
rect 576 -344 577 -342
rect 583 -338 584 -336
rect 583 -344 584 -342
rect 590 -338 591 -336
rect 590 -344 591 -342
rect 597 -338 598 -336
rect 597 -344 598 -342
rect 604 -338 605 -336
rect 604 -344 605 -342
rect 611 -338 612 -336
rect 611 -344 612 -342
rect 618 -338 619 -336
rect 618 -344 619 -342
rect 625 -338 626 -336
rect 625 -344 626 -342
rect 632 -338 633 -336
rect 632 -344 633 -342
rect 639 -338 640 -336
rect 639 -344 640 -342
rect 646 -338 647 -336
rect 646 -344 647 -342
rect 653 -338 654 -336
rect 653 -344 654 -342
rect 660 -338 661 -336
rect 660 -344 661 -342
rect 667 -338 668 -336
rect 667 -344 668 -342
rect 674 -338 675 -336
rect 674 -344 675 -342
rect 681 -338 682 -336
rect 681 -344 682 -342
rect 688 -338 689 -336
rect 688 -344 689 -342
rect 695 -338 696 -336
rect 695 -344 696 -342
rect 702 -338 703 -336
rect 702 -344 703 -342
rect 709 -338 710 -336
rect 709 -344 710 -342
rect 716 -338 717 -336
rect 716 -344 717 -342
rect 723 -338 724 -336
rect 723 -344 724 -342
rect 730 -338 731 -336
rect 730 -344 731 -342
rect 737 -338 738 -336
rect 737 -344 738 -342
rect 2 -417 3 -415
rect 5 -417 6 -415
rect 9 -423 10 -421
rect 16 -417 17 -415
rect 16 -423 17 -421
rect 23 -417 24 -415
rect 23 -423 24 -421
rect 30 -417 31 -415
rect 30 -423 31 -421
rect 37 -417 38 -415
rect 37 -423 38 -421
rect 44 -417 45 -415
rect 44 -423 45 -421
rect 51 -417 52 -415
rect 51 -423 52 -421
rect 58 -423 59 -421
rect 65 -417 66 -415
rect 65 -423 66 -421
rect 72 -417 73 -415
rect 72 -423 73 -421
rect 79 -417 80 -415
rect 79 -423 80 -421
rect 86 -417 87 -415
rect 86 -423 87 -421
rect 93 -417 94 -415
rect 93 -423 94 -421
rect 100 -417 101 -415
rect 100 -423 101 -421
rect 107 -417 108 -415
rect 110 -417 111 -415
rect 107 -423 108 -421
rect 110 -423 111 -421
rect 114 -417 115 -415
rect 114 -423 115 -421
rect 124 -417 125 -415
rect 124 -423 125 -421
rect 128 -417 129 -415
rect 128 -423 129 -421
rect 135 -417 136 -415
rect 135 -423 136 -421
rect 142 -417 143 -415
rect 142 -423 143 -421
rect 149 -417 150 -415
rect 149 -423 150 -421
rect 156 -417 157 -415
rect 156 -423 157 -421
rect 163 -417 164 -415
rect 163 -423 164 -421
rect 170 -417 171 -415
rect 170 -423 171 -421
rect 177 -417 178 -415
rect 177 -423 178 -421
rect 184 -417 185 -415
rect 184 -423 185 -421
rect 191 -417 192 -415
rect 191 -423 192 -421
rect 198 -417 199 -415
rect 198 -423 199 -421
rect 205 -417 206 -415
rect 205 -423 206 -421
rect 212 -417 213 -415
rect 212 -423 213 -421
rect 219 -417 220 -415
rect 222 -417 223 -415
rect 219 -423 220 -421
rect 222 -423 223 -421
rect 226 -417 227 -415
rect 226 -423 227 -421
rect 233 -417 234 -415
rect 233 -423 234 -421
rect 240 -417 241 -415
rect 240 -423 241 -421
rect 247 -417 248 -415
rect 247 -423 248 -421
rect 254 -417 255 -415
rect 254 -423 255 -421
rect 261 -417 262 -415
rect 261 -423 262 -421
rect 268 -417 269 -415
rect 268 -423 269 -421
rect 275 -417 276 -415
rect 275 -423 276 -421
rect 282 -417 283 -415
rect 282 -423 283 -421
rect 289 -417 290 -415
rect 292 -417 293 -415
rect 296 -417 297 -415
rect 296 -423 297 -421
rect 303 -417 304 -415
rect 303 -423 304 -421
rect 310 -417 311 -415
rect 310 -423 311 -421
rect 317 -417 318 -415
rect 317 -423 318 -421
rect 324 -417 325 -415
rect 324 -423 325 -421
rect 331 -417 332 -415
rect 334 -417 335 -415
rect 331 -423 332 -421
rect 334 -423 335 -421
rect 338 -417 339 -415
rect 341 -417 342 -415
rect 338 -423 339 -421
rect 345 -417 346 -415
rect 348 -417 349 -415
rect 345 -423 346 -421
rect 348 -423 349 -421
rect 352 -417 353 -415
rect 352 -423 353 -421
rect 359 -417 360 -415
rect 359 -423 360 -421
rect 366 -417 367 -415
rect 366 -423 367 -421
rect 373 -417 374 -415
rect 376 -417 377 -415
rect 380 -417 381 -415
rect 383 -417 384 -415
rect 380 -423 381 -421
rect 383 -423 384 -421
rect 387 -417 388 -415
rect 387 -423 388 -421
rect 394 -417 395 -415
rect 397 -417 398 -415
rect 394 -423 395 -421
rect 401 -417 402 -415
rect 404 -417 405 -415
rect 404 -423 405 -421
rect 408 -417 409 -415
rect 408 -423 409 -421
rect 415 -417 416 -415
rect 418 -417 419 -415
rect 415 -423 416 -421
rect 418 -423 419 -421
rect 422 -417 423 -415
rect 422 -423 423 -421
rect 432 -417 433 -415
rect 432 -423 433 -421
rect 436 -417 437 -415
rect 436 -423 437 -421
rect 443 -417 444 -415
rect 443 -423 444 -421
rect 450 -417 451 -415
rect 450 -423 451 -421
rect 457 -417 458 -415
rect 457 -423 458 -421
rect 464 -417 465 -415
rect 464 -423 465 -421
rect 474 -417 475 -415
rect 471 -423 472 -421
rect 474 -423 475 -421
rect 478 -417 479 -415
rect 478 -423 479 -421
rect 485 -417 486 -415
rect 485 -423 486 -421
rect 492 -417 493 -415
rect 492 -423 493 -421
rect 499 -417 500 -415
rect 499 -423 500 -421
rect 506 -423 507 -421
rect 513 -417 514 -415
rect 513 -423 514 -421
rect 523 -417 524 -415
rect 520 -423 521 -421
rect 523 -423 524 -421
rect 527 -417 528 -415
rect 527 -423 528 -421
rect 534 -417 535 -415
rect 534 -423 535 -421
rect 541 -417 542 -415
rect 541 -423 542 -421
rect 548 -417 549 -415
rect 548 -423 549 -421
rect 558 -417 559 -415
rect 555 -423 556 -421
rect 562 -417 563 -415
rect 562 -423 563 -421
rect 569 -417 570 -415
rect 569 -423 570 -421
rect 576 -417 577 -415
rect 576 -423 577 -421
rect 583 -417 584 -415
rect 590 -417 591 -415
rect 590 -423 591 -421
rect 597 -417 598 -415
rect 597 -423 598 -421
rect 604 -417 605 -415
rect 604 -423 605 -421
rect 611 -417 612 -415
rect 611 -423 612 -421
rect 618 -417 619 -415
rect 618 -423 619 -421
rect 625 -417 626 -415
rect 625 -423 626 -421
rect 632 -417 633 -415
rect 632 -423 633 -421
rect 639 -417 640 -415
rect 639 -423 640 -421
rect 646 -417 647 -415
rect 646 -423 647 -421
rect 653 -417 654 -415
rect 653 -423 654 -421
rect 660 -417 661 -415
rect 660 -423 661 -421
rect 667 -417 668 -415
rect 667 -423 668 -421
rect 674 -417 675 -415
rect 674 -423 675 -421
rect 681 -417 682 -415
rect 681 -423 682 -421
rect 688 -417 689 -415
rect 688 -423 689 -421
rect 695 -417 696 -415
rect 695 -423 696 -421
rect 702 -417 703 -415
rect 702 -423 703 -421
rect 705 -423 706 -421
rect 709 -417 710 -415
rect 709 -423 710 -421
rect 716 -417 717 -415
rect 716 -423 717 -421
rect 723 -417 724 -415
rect 723 -423 724 -421
rect 730 -417 731 -415
rect 730 -423 731 -421
rect 737 -417 738 -415
rect 737 -423 738 -421
rect 744 -417 745 -415
rect 744 -423 745 -421
rect 751 -417 752 -415
rect 751 -423 752 -421
rect 758 -417 759 -415
rect 758 -423 759 -421
rect 765 -417 766 -415
rect 765 -423 766 -421
rect 772 -417 773 -415
rect 772 -423 773 -421
rect 779 -417 780 -415
rect 779 -423 780 -421
rect 786 -417 787 -415
rect 786 -423 787 -421
rect 793 -417 794 -415
rect 793 -423 794 -421
rect 800 -417 801 -415
rect 800 -423 801 -421
rect 807 -417 808 -415
rect 807 -423 808 -421
rect 814 -417 815 -415
rect 814 -423 815 -421
rect 9 -510 10 -508
rect 9 -516 10 -514
rect 16 -510 17 -508
rect 16 -516 17 -514
rect 23 -510 24 -508
rect 23 -516 24 -514
rect 30 -510 31 -508
rect 30 -516 31 -514
rect 37 -510 38 -508
rect 37 -516 38 -514
rect 44 -510 45 -508
rect 47 -510 48 -508
rect 47 -516 48 -514
rect 51 -510 52 -508
rect 51 -516 52 -514
rect 58 -510 59 -508
rect 61 -510 62 -508
rect 61 -516 62 -514
rect 65 -510 66 -508
rect 65 -516 66 -514
rect 72 -510 73 -508
rect 72 -516 73 -514
rect 79 -510 80 -508
rect 79 -516 80 -514
rect 86 -510 87 -508
rect 86 -516 87 -514
rect 93 -510 94 -508
rect 93 -516 94 -514
rect 100 -510 101 -508
rect 100 -516 101 -514
rect 103 -516 104 -514
rect 107 -510 108 -508
rect 107 -516 108 -514
rect 114 -510 115 -508
rect 114 -516 115 -514
rect 121 -510 122 -508
rect 121 -516 122 -514
rect 128 -510 129 -508
rect 128 -516 129 -514
rect 138 -510 139 -508
rect 135 -516 136 -514
rect 142 -510 143 -508
rect 142 -516 143 -514
rect 149 -510 150 -508
rect 149 -516 150 -514
rect 156 -510 157 -508
rect 156 -516 157 -514
rect 163 -510 164 -508
rect 163 -516 164 -514
rect 170 -510 171 -508
rect 170 -516 171 -514
rect 177 -510 178 -508
rect 177 -516 178 -514
rect 184 -510 185 -508
rect 184 -516 185 -514
rect 191 -510 192 -508
rect 191 -516 192 -514
rect 198 -510 199 -508
rect 198 -516 199 -514
rect 205 -510 206 -508
rect 205 -516 206 -514
rect 212 -510 213 -508
rect 212 -516 213 -514
rect 222 -510 223 -508
rect 219 -516 220 -514
rect 222 -516 223 -514
rect 226 -516 227 -514
rect 233 -510 234 -508
rect 233 -516 234 -514
rect 240 -510 241 -508
rect 240 -516 241 -514
rect 247 -510 248 -508
rect 247 -516 248 -514
rect 254 -510 255 -508
rect 254 -516 255 -514
rect 264 -510 265 -508
rect 261 -516 262 -514
rect 264 -516 265 -514
rect 268 -510 269 -508
rect 268 -516 269 -514
rect 275 -510 276 -508
rect 275 -516 276 -514
rect 282 -510 283 -508
rect 282 -516 283 -514
rect 289 -510 290 -508
rect 289 -516 290 -514
rect 296 -510 297 -508
rect 296 -516 297 -514
rect 303 -510 304 -508
rect 306 -516 307 -514
rect 310 -510 311 -508
rect 310 -516 311 -514
rect 313 -516 314 -514
rect 317 -510 318 -508
rect 317 -516 318 -514
rect 324 -510 325 -508
rect 324 -516 325 -514
rect 331 -510 332 -508
rect 331 -516 332 -514
rect 338 -510 339 -508
rect 338 -516 339 -514
rect 345 -510 346 -508
rect 345 -516 346 -514
rect 355 -510 356 -508
rect 359 -510 360 -508
rect 359 -516 360 -514
rect 366 -510 367 -508
rect 366 -516 367 -514
rect 369 -516 370 -514
rect 373 -510 374 -508
rect 373 -516 374 -514
rect 380 -510 381 -508
rect 383 -510 384 -508
rect 383 -516 384 -514
rect 387 -516 388 -514
rect 390 -516 391 -514
rect 394 -510 395 -508
rect 394 -516 395 -514
rect 401 -510 402 -508
rect 404 -510 405 -508
rect 401 -516 402 -514
rect 411 -516 412 -514
rect 415 -510 416 -508
rect 415 -516 416 -514
rect 422 -510 423 -508
rect 422 -516 423 -514
rect 429 -516 430 -514
rect 432 -516 433 -514
rect 436 -510 437 -508
rect 436 -516 437 -514
rect 443 -510 444 -508
rect 443 -516 444 -514
rect 450 -510 451 -508
rect 450 -516 451 -514
rect 457 -510 458 -508
rect 457 -516 458 -514
rect 464 -510 465 -508
rect 464 -516 465 -514
rect 474 -510 475 -508
rect 474 -516 475 -514
rect 478 -510 479 -508
rect 478 -516 479 -514
rect 485 -510 486 -508
rect 485 -516 486 -514
rect 492 -510 493 -508
rect 492 -516 493 -514
rect 495 -516 496 -514
rect 499 -510 500 -508
rect 499 -516 500 -514
rect 506 -510 507 -508
rect 506 -516 507 -514
rect 513 -510 514 -508
rect 513 -516 514 -514
rect 520 -510 521 -508
rect 520 -516 521 -514
rect 527 -510 528 -508
rect 527 -516 528 -514
rect 534 -510 535 -508
rect 534 -516 535 -514
rect 541 -510 542 -508
rect 541 -516 542 -514
rect 548 -510 549 -508
rect 548 -516 549 -514
rect 558 -510 559 -508
rect 558 -516 559 -514
rect 562 -510 563 -508
rect 562 -516 563 -514
rect 569 -510 570 -508
rect 569 -516 570 -514
rect 576 -510 577 -508
rect 576 -516 577 -514
rect 583 -516 584 -514
rect 590 -510 591 -508
rect 590 -516 591 -514
rect 597 -510 598 -508
rect 597 -516 598 -514
rect 604 -510 605 -508
rect 604 -516 605 -514
rect 611 -510 612 -508
rect 611 -516 612 -514
rect 618 -510 619 -508
rect 618 -516 619 -514
rect 625 -510 626 -508
rect 625 -516 626 -514
rect 632 -510 633 -508
rect 632 -516 633 -514
rect 639 -510 640 -508
rect 639 -516 640 -514
rect 646 -510 647 -508
rect 646 -516 647 -514
rect 653 -510 654 -508
rect 653 -516 654 -514
rect 660 -510 661 -508
rect 660 -516 661 -514
rect 667 -510 668 -508
rect 667 -516 668 -514
rect 674 -510 675 -508
rect 674 -516 675 -514
rect 681 -510 682 -508
rect 681 -516 682 -514
rect 688 -510 689 -508
rect 688 -516 689 -514
rect 695 -510 696 -508
rect 695 -516 696 -514
rect 702 -510 703 -508
rect 705 -510 706 -508
rect 702 -516 703 -514
rect 709 -510 710 -508
rect 709 -516 710 -514
rect 716 -510 717 -508
rect 716 -516 717 -514
rect 723 -510 724 -508
rect 723 -516 724 -514
rect 730 -510 731 -508
rect 730 -516 731 -514
rect 737 -510 738 -508
rect 737 -516 738 -514
rect 744 -510 745 -508
rect 744 -516 745 -514
rect 751 -510 752 -508
rect 751 -516 752 -514
rect 758 -510 759 -508
rect 758 -516 759 -514
rect 765 -510 766 -508
rect 765 -516 766 -514
rect 772 -510 773 -508
rect 772 -516 773 -514
rect 779 -510 780 -508
rect 779 -516 780 -514
rect 786 -510 787 -508
rect 786 -516 787 -514
rect 793 -510 794 -508
rect 793 -516 794 -514
rect 800 -510 801 -508
rect 800 -516 801 -514
rect 9 -579 10 -577
rect 9 -585 10 -583
rect 16 -579 17 -577
rect 16 -585 17 -583
rect 23 -579 24 -577
rect 23 -585 24 -583
rect 26 -585 27 -583
rect 30 -579 31 -577
rect 30 -585 31 -583
rect 37 -579 38 -577
rect 37 -585 38 -583
rect 44 -579 45 -577
rect 44 -585 45 -583
rect 54 -579 55 -577
rect 58 -579 59 -577
rect 58 -585 59 -583
rect 65 -579 66 -577
rect 65 -585 66 -583
rect 72 -579 73 -577
rect 72 -585 73 -583
rect 79 -579 80 -577
rect 79 -585 80 -583
rect 86 -579 87 -577
rect 86 -585 87 -583
rect 93 -579 94 -577
rect 93 -585 94 -583
rect 100 -579 101 -577
rect 100 -585 101 -583
rect 110 -579 111 -577
rect 107 -585 108 -583
rect 110 -585 111 -583
rect 114 -579 115 -577
rect 114 -585 115 -583
rect 121 -585 122 -583
rect 124 -585 125 -583
rect 128 -579 129 -577
rect 131 -579 132 -577
rect 135 -579 136 -577
rect 135 -585 136 -583
rect 138 -585 139 -583
rect 142 -579 143 -577
rect 142 -585 143 -583
rect 149 -579 150 -577
rect 149 -585 150 -583
rect 156 -579 157 -577
rect 156 -585 157 -583
rect 163 -579 164 -577
rect 163 -585 164 -583
rect 170 -579 171 -577
rect 170 -585 171 -583
rect 177 -579 178 -577
rect 177 -585 178 -583
rect 184 -579 185 -577
rect 184 -585 185 -583
rect 191 -579 192 -577
rect 191 -585 192 -583
rect 198 -579 199 -577
rect 198 -585 199 -583
rect 205 -579 206 -577
rect 205 -585 206 -583
rect 212 -579 213 -577
rect 212 -585 213 -583
rect 219 -579 220 -577
rect 219 -585 220 -583
rect 226 -579 227 -577
rect 226 -585 227 -583
rect 233 -579 234 -577
rect 233 -585 234 -583
rect 240 -579 241 -577
rect 240 -585 241 -583
rect 247 -579 248 -577
rect 247 -585 248 -583
rect 254 -579 255 -577
rect 257 -579 258 -577
rect 254 -585 255 -583
rect 257 -585 258 -583
rect 261 -579 262 -577
rect 261 -585 262 -583
rect 268 -579 269 -577
rect 268 -585 269 -583
rect 275 -579 276 -577
rect 275 -585 276 -583
rect 282 -579 283 -577
rect 282 -585 283 -583
rect 289 -579 290 -577
rect 289 -585 290 -583
rect 296 -585 297 -583
rect 303 -579 304 -577
rect 303 -585 304 -583
rect 313 -579 314 -577
rect 310 -585 311 -583
rect 313 -585 314 -583
rect 317 -579 318 -577
rect 317 -585 318 -583
rect 320 -585 321 -583
rect 324 -579 325 -577
rect 324 -585 325 -583
rect 331 -579 332 -577
rect 334 -579 335 -577
rect 331 -585 332 -583
rect 334 -585 335 -583
rect 338 -579 339 -577
rect 338 -585 339 -583
rect 345 -579 346 -577
rect 345 -585 346 -583
rect 352 -579 353 -577
rect 352 -585 353 -583
rect 359 -579 360 -577
rect 359 -585 360 -583
rect 366 -579 367 -577
rect 366 -585 367 -583
rect 373 -579 374 -577
rect 373 -585 374 -583
rect 380 -579 381 -577
rect 383 -579 384 -577
rect 380 -585 381 -583
rect 383 -585 384 -583
rect 387 -579 388 -577
rect 387 -585 388 -583
rect 394 -579 395 -577
rect 394 -585 395 -583
rect 401 -579 402 -577
rect 401 -585 402 -583
rect 408 -579 409 -577
rect 408 -585 409 -583
rect 415 -579 416 -577
rect 418 -579 419 -577
rect 415 -585 416 -583
rect 422 -579 423 -577
rect 422 -585 423 -583
rect 429 -579 430 -577
rect 429 -585 430 -583
rect 436 -579 437 -577
rect 436 -585 437 -583
rect 443 -579 444 -577
rect 443 -585 444 -583
rect 450 -579 451 -577
rect 450 -585 451 -583
rect 457 -579 458 -577
rect 460 -585 461 -583
rect 464 -579 465 -577
rect 467 -579 468 -577
rect 464 -585 465 -583
rect 467 -585 468 -583
rect 471 -579 472 -577
rect 471 -585 472 -583
rect 478 -579 479 -577
rect 478 -585 479 -583
rect 485 -579 486 -577
rect 488 -579 489 -577
rect 485 -585 486 -583
rect 492 -579 493 -577
rect 492 -585 493 -583
rect 499 -579 500 -577
rect 499 -585 500 -583
rect 506 -579 507 -577
rect 506 -585 507 -583
rect 509 -585 510 -583
rect 513 -585 514 -583
rect 516 -585 517 -583
rect 520 -579 521 -577
rect 520 -585 521 -583
rect 527 -579 528 -577
rect 527 -585 528 -583
rect 534 -579 535 -577
rect 534 -585 535 -583
rect 541 -579 542 -577
rect 541 -585 542 -583
rect 551 -579 552 -577
rect 548 -585 549 -583
rect 555 -579 556 -577
rect 555 -585 556 -583
rect 562 -579 563 -577
rect 562 -585 563 -583
rect 569 -579 570 -577
rect 569 -585 570 -583
rect 576 -579 577 -577
rect 576 -585 577 -583
rect 583 -579 584 -577
rect 583 -585 584 -583
rect 590 -579 591 -577
rect 590 -585 591 -583
rect 597 -579 598 -577
rect 597 -585 598 -583
rect 604 -579 605 -577
rect 604 -585 605 -583
rect 611 -579 612 -577
rect 611 -585 612 -583
rect 618 -579 619 -577
rect 618 -585 619 -583
rect 625 -579 626 -577
rect 625 -585 626 -583
rect 632 -579 633 -577
rect 632 -585 633 -583
rect 639 -579 640 -577
rect 639 -585 640 -583
rect 646 -579 647 -577
rect 646 -585 647 -583
rect 653 -579 654 -577
rect 653 -585 654 -583
rect 660 -579 661 -577
rect 660 -585 661 -583
rect 667 -579 668 -577
rect 667 -585 668 -583
rect 674 -579 675 -577
rect 674 -585 675 -583
rect 681 -579 682 -577
rect 681 -585 682 -583
rect 688 -579 689 -577
rect 688 -585 689 -583
rect 695 -579 696 -577
rect 695 -585 696 -583
rect 702 -579 703 -577
rect 702 -585 703 -583
rect 709 -579 710 -577
rect 709 -585 710 -583
rect 716 -579 717 -577
rect 716 -585 717 -583
rect 723 -579 724 -577
rect 723 -585 724 -583
rect 730 -579 731 -577
rect 730 -585 731 -583
rect 737 -579 738 -577
rect 737 -585 738 -583
rect 744 -579 745 -577
rect 744 -585 745 -583
rect 751 -579 752 -577
rect 751 -585 752 -583
rect 758 -579 759 -577
rect 758 -585 759 -583
rect 765 -579 766 -577
rect 765 -585 766 -583
rect 772 -579 773 -577
rect 772 -585 773 -583
rect 779 -579 780 -577
rect 779 -585 780 -583
rect 786 -579 787 -577
rect 786 -585 787 -583
rect 793 -579 794 -577
rect 793 -585 794 -583
rect 800 -579 801 -577
rect 800 -585 801 -583
rect 807 -579 808 -577
rect 807 -585 808 -583
rect 814 -579 815 -577
rect 814 -585 815 -583
rect 821 -579 822 -577
rect 821 -585 822 -583
rect 2 -668 3 -666
rect 2 -674 3 -672
rect 9 -668 10 -666
rect 9 -674 10 -672
rect 16 -668 17 -666
rect 16 -674 17 -672
rect 23 -668 24 -666
rect 23 -674 24 -672
rect 30 -668 31 -666
rect 30 -674 31 -672
rect 37 -668 38 -666
rect 37 -674 38 -672
rect 44 -668 45 -666
rect 44 -674 45 -672
rect 51 -668 52 -666
rect 54 -668 55 -666
rect 51 -674 52 -672
rect 58 -668 59 -666
rect 61 -668 62 -666
rect 61 -674 62 -672
rect 68 -668 69 -666
rect 65 -674 66 -672
rect 68 -674 69 -672
rect 72 -668 73 -666
rect 72 -674 73 -672
rect 79 -668 80 -666
rect 79 -674 80 -672
rect 86 -668 87 -666
rect 86 -674 87 -672
rect 93 -668 94 -666
rect 93 -674 94 -672
rect 100 -668 101 -666
rect 100 -674 101 -672
rect 107 -668 108 -666
rect 110 -668 111 -666
rect 107 -674 108 -672
rect 114 -668 115 -666
rect 114 -674 115 -672
rect 121 -668 122 -666
rect 121 -674 122 -672
rect 128 -668 129 -666
rect 128 -674 129 -672
rect 135 -668 136 -666
rect 135 -674 136 -672
rect 142 -668 143 -666
rect 142 -674 143 -672
rect 149 -668 150 -666
rect 149 -674 150 -672
rect 156 -668 157 -666
rect 156 -674 157 -672
rect 163 -668 164 -666
rect 163 -674 164 -672
rect 170 -668 171 -666
rect 170 -674 171 -672
rect 177 -668 178 -666
rect 177 -674 178 -672
rect 184 -668 185 -666
rect 184 -674 185 -672
rect 191 -668 192 -666
rect 191 -674 192 -672
rect 198 -668 199 -666
rect 198 -674 199 -672
rect 205 -668 206 -666
rect 205 -674 206 -672
rect 212 -668 213 -666
rect 215 -668 216 -666
rect 212 -674 213 -672
rect 219 -668 220 -666
rect 219 -674 220 -672
rect 226 -668 227 -666
rect 229 -668 230 -666
rect 229 -674 230 -672
rect 233 -668 234 -666
rect 233 -674 234 -672
rect 240 -668 241 -666
rect 240 -674 241 -672
rect 247 -668 248 -666
rect 247 -674 248 -672
rect 254 -668 255 -666
rect 254 -674 255 -672
rect 261 -668 262 -666
rect 261 -674 262 -672
rect 268 -668 269 -666
rect 271 -668 272 -666
rect 268 -674 269 -672
rect 271 -674 272 -672
rect 275 -668 276 -666
rect 275 -674 276 -672
rect 282 -668 283 -666
rect 282 -674 283 -672
rect 289 -668 290 -666
rect 292 -668 293 -666
rect 296 -668 297 -666
rect 299 -668 300 -666
rect 296 -674 297 -672
rect 303 -668 304 -666
rect 303 -674 304 -672
rect 310 -668 311 -666
rect 310 -674 311 -672
rect 317 -668 318 -666
rect 317 -674 318 -672
rect 324 -668 325 -666
rect 324 -674 325 -672
rect 331 -668 332 -666
rect 331 -674 332 -672
rect 338 -668 339 -666
rect 338 -674 339 -672
rect 345 -668 346 -666
rect 348 -668 349 -666
rect 348 -674 349 -672
rect 352 -668 353 -666
rect 352 -674 353 -672
rect 359 -668 360 -666
rect 359 -674 360 -672
rect 366 -668 367 -666
rect 369 -668 370 -666
rect 369 -674 370 -672
rect 373 -668 374 -666
rect 373 -674 374 -672
rect 383 -668 384 -666
rect 380 -674 381 -672
rect 387 -668 388 -666
rect 387 -674 388 -672
rect 394 -668 395 -666
rect 394 -674 395 -672
rect 401 -668 402 -666
rect 401 -674 402 -672
rect 408 -668 409 -666
rect 408 -674 409 -672
rect 415 -668 416 -666
rect 415 -674 416 -672
rect 418 -674 419 -672
rect 422 -668 423 -666
rect 422 -674 423 -672
rect 429 -668 430 -666
rect 429 -674 430 -672
rect 436 -668 437 -666
rect 436 -674 437 -672
rect 443 -668 444 -666
rect 443 -674 444 -672
rect 450 -668 451 -666
rect 453 -668 454 -666
rect 453 -674 454 -672
rect 457 -668 458 -666
rect 460 -668 461 -666
rect 460 -674 461 -672
rect 464 -668 465 -666
rect 464 -674 465 -672
rect 471 -668 472 -666
rect 471 -674 472 -672
rect 478 -668 479 -666
rect 478 -674 479 -672
rect 485 -668 486 -666
rect 485 -674 486 -672
rect 492 -668 493 -666
rect 492 -674 493 -672
rect 499 -668 500 -666
rect 499 -674 500 -672
rect 506 -668 507 -666
rect 506 -674 507 -672
rect 513 -668 514 -666
rect 513 -674 514 -672
rect 520 -668 521 -666
rect 520 -674 521 -672
rect 527 -668 528 -666
rect 527 -674 528 -672
rect 534 -668 535 -666
rect 534 -674 535 -672
rect 544 -674 545 -672
rect 548 -668 549 -666
rect 548 -674 549 -672
rect 555 -668 556 -666
rect 555 -674 556 -672
rect 562 -668 563 -666
rect 562 -674 563 -672
rect 569 -668 570 -666
rect 569 -674 570 -672
rect 576 -668 577 -666
rect 576 -674 577 -672
rect 583 -668 584 -666
rect 583 -674 584 -672
rect 590 -668 591 -666
rect 590 -674 591 -672
rect 597 -668 598 -666
rect 597 -674 598 -672
rect 604 -668 605 -666
rect 604 -674 605 -672
rect 611 -668 612 -666
rect 611 -674 612 -672
rect 618 -668 619 -666
rect 618 -674 619 -672
rect 625 -668 626 -666
rect 625 -674 626 -672
rect 632 -668 633 -666
rect 632 -674 633 -672
rect 639 -668 640 -666
rect 639 -674 640 -672
rect 646 -668 647 -666
rect 646 -674 647 -672
rect 653 -668 654 -666
rect 653 -674 654 -672
rect 660 -668 661 -666
rect 660 -674 661 -672
rect 667 -668 668 -666
rect 667 -674 668 -672
rect 674 -668 675 -666
rect 674 -674 675 -672
rect 681 -668 682 -666
rect 681 -674 682 -672
rect 688 -668 689 -666
rect 688 -674 689 -672
rect 695 -668 696 -666
rect 695 -674 696 -672
rect 702 -668 703 -666
rect 702 -674 703 -672
rect 709 -668 710 -666
rect 709 -674 710 -672
rect 716 -668 717 -666
rect 716 -674 717 -672
rect 723 -668 724 -666
rect 723 -674 724 -672
rect 730 -668 731 -666
rect 730 -674 731 -672
rect 737 -668 738 -666
rect 737 -674 738 -672
rect 744 -668 745 -666
rect 744 -674 745 -672
rect 751 -668 752 -666
rect 751 -674 752 -672
rect 758 -668 759 -666
rect 758 -674 759 -672
rect 765 -668 766 -666
rect 765 -674 766 -672
rect 772 -668 773 -666
rect 772 -674 773 -672
rect 779 -668 780 -666
rect 779 -674 780 -672
rect 786 -668 787 -666
rect 793 -668 794 -666
rect 12 -735 13 -733
rect 16 -735 17 -733
rect 19 -741 20 -739
rect 23 -735 24 -733
rect 23 -741 24 -739
rect 30 -735 31 -733
rect 30 -741 31 -739
rect 37 -735 38 -733
rect 37 -741 38 -739
rect 44 -735 45 -733
rect 44 -741 45 -739
rect 51 -735 52 -733
rect 51 -741 52 -739
rect 58 -735 59 -733
rect 58 -741 59 -739
rect 65 -735 66 -733
rect 68 -735 69 -733
rect 68 -741 69 -739
rect 72 -735 73 -733
rect 72 -741 73 -739
rect 79 -735 80 -733
rect 79 -741 80 -739
rect 89 -735 90 -733
rect 86 -741 87 -739
rect 89 -741 90 -739
rect 93 -735 94 -733
rect 93 -741 94 -739
rect 100 -735 101 -733
rect 100 -741 101 -739
rect 107 -735 108 -733
rect 107 -741 108 -739
rect 114 -735 115 -733
rect 114 -741 115 -739
rect 121 -735 122 -733
rect 121 -741 122 -739
rect 128 -735 129 -733
rect 131 -735 132 -733
rect 135 -735 136 -733
rect 135 -741 136 -739
rect 142 -735 143 -733
rect 142 -741 143 -739
rect 149 -735 150 -733
rect 149 -741 150 -739
rect 156 -735 157 -733
rect 156 -741 157 -739
rect 163 -735 164 -733
rect 166 -735 167 -733
rect 166 -741 167 -739
rect 170 -735 171 -733
rect 170 -741 171 -739
rect 177 -735 178 -733
rect 177 -741 178 -739
rect 184 -735 185 -733
rect 184 -741 185 -739
rect 191 -735 192 -733
rect 191 -741 192 -739
rect 198 -735 199 -733
rect 198 -741 199 -739
rect 205 -735 206 -733
rect 205 -741 206 -739
rect 212 -735 213 -733
rect 212 -741 213 -739
rect 219 -735 220 -733
rect 219 -741 220 -739
rect 226 -735 227 -733
rect 229 -735 230 -733
rect 229 -741 230 -739
rect 233 -735 234 -733
rect 233 -741 234 -739
rect 240 -735 241 -733
rect 247 -735 248 -733
rect 247 -741 248 -739
rect 254 -735 255 -733
rect 254 -741 255 -739
rect 261 -735 262 -733
rect 261 -741 262 -739
rect 268 -735 269 -733
rect 271 -735 272 -733
rect 268 -741 269 -739
rect 275 -735 276 -733
rect 275 -741 276 -739
rect 282 -735 283 -733
rect 282 -741 283 -739
rect 289 -735 290 -733
rect 289 -741 290 -739
rect 296 -735 297 -733
rect 296 -741 297 -739
rect 303 -735 304 -733
rect 303 -741 304 -739
rect 310 -735 311 -733
rect 310 -741 311 -739
rect 317 -735 318 -733
rect 320 -735 321 -733
rect 317 -741 318 -739
rect 320 -741 321 -739
rect 324 -735 325 -733
rect 324 -741 325 -739
rect 331 -735 332 -733
rect 331 -741 332 -739
rect 338 -735 339 -733
rect 338 -741 339 -739
rect 345 -735 346 -733
rect 345 -741 346 -739
rect 348 -741 349 -739
rect 352 -735 353 -733
rect 352 -741 353 -739
rect 359 -735 360 -733
rect 359 -741 360 -739
rect 366 -735 367 -733
rect 366 -741 367 -739
rect 373 -735 374 -733
rect 373 -741 374 -739
rect 380 -735 381 -733
rect 380 -741 381 -739
rect 383 -741 384 -739
rect 387 -735 388 -733
rect 387 -741 388 -739
rect 394 -735 395 -733
rect 397 -741 398 -739
rect 401 -735 402 -733
rect 401 -741 402 -739
rect 408 -735 409 -733
rect 408 -741 409 -739
rect 415 -735 416 -733
rect 415 -741 416 -739
rect 422 -735 423 -733
rect 425 -735 426 -733
rect 422 -741 423 -739
rect 425 -741 426 -739
rect 429 -735 430 -733
rect 429 -741 430 -739
rect 436 -735 437 -733
rect 436 -741 437 -739
rect 443 -735 444 -733
rect 446 -735 447 -733
rect 443 -741 444 -739
rect 446 -741 447 -739
rect 450 -735 451 -733
rect 450 -741 451 -739
rect 453 -741 454 -739
rect 457 -735 458 -733
rect 457 -741 458 -739
rect 464 -735 465 -733
rect 464 -741 465 -739
rect 471 -735 472 -733
rect 471 -741 472 -739
rect 478 -735 479 -733
rect 478 -741 479 -739
rect 485 -735 486 -733
rect 485 -741 486 -739
rect 492 -735 493 -733
rect 492 -741 493 -739
rect 499 -735 500 -733
rect 499 -741 500 -739
rect 506 -735 507 -733
rect 506 -741 507 -739
rect 513 -735 514 -733
rect 513 -741 514 -739
rect 523 -735 524 -733
rect 527 -735 528 -733
rect 530 -735 531 -733
rect 527 -741 528 -739
rect 530 -741 531 -739
rect 534 -735 535 -733
rect 534 -741 535 -739
rect 541 -735 542 -733
rect 541 -741 542 -739
rect 551 -735 552 -733
rect 548 -741 549 -739
rect 555 -735 556 -733
rect 555 -741 556 -739
rect 562 -735 563 -733
rect 562 -741 563 -739
rect 569 -741 570 -739
rect 572 -741 573 -739
rect 576 -735 577 -733
rect 576 -741 577 -739
rect 583 -735 584 -733
rect 583 -741 584 -739
rect 590 -735 591 -733
rect 590 -741 591 -739
rect 597 -735 598 -733
rect 597 -741 598 -739
rect 604 -735 605 -733
rect 604 -741 605 -739
rect 611 -735 612 -733
rect 611 -741 612 -739
rect 618 -735 619 -733
rect 618 -741 619 -739
rect 625 -735 626 -733
rect 625 -741 626 -739
rect 632 -735 633 -733
rect 632 -741 633 -739
rect 639 -735 640 -733
rect 639 -741 640 -739
rect 646 -735 647 -733
rect 646 -741 647 -739
rect 653 -735 654 -733
rect 653 -741 654 -739
rect 660 -735 661 -733
rect 660 -741 661 -739
rect 667 -735 668 -733
rect 667 -741 668 -739
rect 674 -735 675 -733
rect 674 -741 675 -739
rect 681 -735 682 -733
rect 681 -741 682 -739
rect 688 -735 689 -733
rect 688 -741 689 -739
rect 695 -735 696 -733
rect 695 -741 696 -739
rect 702 -735 703 -733
rect 702 -741 703 -739
rect 709 -735 710 -733
rect 709 -741 710 -739
rect 716 -735 717 -733
rect 716 -741 717 -739
rect 723 -735 724 -733
rect 723 -741 724 -739
rect 730 -735 731 -733
rect 730 -741 731 -739
rect 737 -735 738 -733
rect 737 -741 738 -739
rect 744 -735 745 -733
rect 744 -741 745 -739
rect 751 -735 752 -733
rect 751 -741 752 -739
rect 758 -735 759 -733
rect 758 -741 759 -739
rect 765 -735 766 -733
rect 765 -741 766 -739
rect 772 -735 773 -733
rect 772 -741 773 -739
rect 779 -735 780 -733
rect 782 -735 783 -733
rect 782 -741 783 -739
rect 786 -735 787 -733
rect 786 -741 787 -739
rect 793 -735 794 -733
rect 793 -741 794 -739
rect 800 -735 801 -733
rect 800 -741 801 -739
rect 807 -735 808 -733
rect 807 -741 808 -739
rect 2 -806 3 -804
rect 9 -806 10 -804
rect 9 -812 10 -810
rect 16 -806 17 -804
rect 16 -812 17 -810
rect 23 -806 24 -804
rect 23 -812 24 -810
rect 30 -806 31 -804
rect 30 -812 31 -810
rect 37 -806 38 -804
rect 40 -806 41 -804
rect 40 -812 41 -810
rect 44 -806 45 -804
rect 44 -812 45 -810
rect 51 -806 52 -804
rect 51 -812 52 -810
rect 58 -806 59 -804
rect 58 -812 59 -810
rect 65 -806 66 -804
rect 65 -812 66 -810
rect 72 -806 73 -804
rect 75 -806 76 -804
rect 72 -812 73 -810
rect 75 -812 76 -810
rect 79 -806 80 -804
rect 79 -812 80 -810
rect 86 -806 87 -804
rect 86 -812 87 -810
rect 93 -806 94 -804
rect 93 -812 94 -810
rect 100 -806 101 -804
rect 100 -812 101 -810
rect 107 -806 108 -804
rect 107 -812 108 -810
rect 114 -806 115 -804
rect 114 -812 115 -810
rect 121 -806 122 -804
rect 121 -812 122 -810
rect 128 -806 129 -804
rect 128 -812 129 -810
rect 131 -812 132 -810
rect 135 -806 136 -804
rect 135 -812 136 -810
rect 142 -806 143 -804
rect 142 -812 143 -810
rect 149 -806 150 -804
rect 149 -812 150 -810
rect 159 -806 160 -804
rect 156 -812 157 -810
rect 159 -812 160 -810
rect 163 -806 164 -804
rect 163 -812 164 -810
rect 170 -806 171 -804
rect 170 -812 171 -810
rect 177 -806 178 -804
rect 177 -812 178 -810
rect 184 -806 185 -804
rect 184 -812 185 -810
rect 191 -806 192 -804
rect 191 -812 192 -810
rect 198 -806 199 -804
rect 198 -812 199 -810
rect 205 -806 206 -804
rect 205 -812 206 -810
rect 212 -806 213 -804
rect 215 -806 216 -804
rect 219 -806 220 -804
rect 219 -812 220 -810
rect 226 -806 227 -804
rect 226 -812 227 -810
rect 233 -806 234 -804
rect 233 -812 234 -810
rect 240 -812 241 -810
rect 247 -806 248 -804
rect 247 -812 248 -810
rect 250 -812 251 -810
rect 254 -806 255 -804
rect 257 -812 258 -810
rect 261 -806 262 -804
rect 261 -812 262 -810
rect 268 -806 269 -804
rect 268 -812 269 -810
rect 275 -806 276 -804
rect 275 -812 276 -810
rect 282 -806 283 -804
rect 285 -806 286 -804
rect 282 -812 283 -810
rect 289 -806 290 -804
rect 289 -812 290 -810
rect 296 -806 297 -804
rect 296 -812 297 -810
rect 303 -806 304 -804
rect 303 -812 304 -810
rect 310 -806 311 -804
rect 317 -806 318 -804
rect 317 -812 318 -810
rect 324 -806 325 -804
rect 324 -812 325 -810
rect 331 -806 332 -804
rect 331 -812 332 -810
rect 338 -806 339 -804
rect 338 -812 339 -810
rect 345 -806 346 -804
rect 345 -812 346 -810
rect 352 -806 353 -804
rect 352 -812 353 -810
rect 359 -806 360 -804
rect 362 -806 363 -804
rect 366 -806 367 -804
rect 366 -812 367 -810
rect 373 -806 374 -804
rect 376 -806 377 -804
rect 373 -812 374 -810
rect 376 -812 377 -810
rect 380 -806 381 -804
rect 380 -812 381 -810
rect 387 -806 388 -804
rect 387 -812 388 -810
rect 397 -812 398 -810
rect 401 -806 402 -804
rect 404 -806 405 -804
rect 404 -812 405 -810
rect 411 -806 412 -804
rect 411 -812 412 -810
rect 415 -806 416 -804
rect 415 -812 416 -810
rect 422 -806 423 -804
rect 422 -812 423 -810
rect 429 -806 430 -804
rect 429 -812 430 -810
rect 436 -806 437 -804
rect 436 -812 437 -810
rect 443 -806 444 -804
rect 443 -812 444 -810
rect 450 -806 451 -804
rect 453 -806 454 -804
rect 450 -812 451 -810
rect 457 -806 458 -804
rect 457 -812 458 -810
rect 464 -806 465 -804
rect 464 -812 465 -810
rect 471 -806 472 -804
rect 471 -812 472 -810
rect 478 -806 479 -804
rect 481 -806 482 -804
rect 481 -812 482 -810
rect 485 -806 486 -804
rect 485 -812 486 -810
rect 492 -806 493 -804
rect 492 -812 493 -810
rect 499 -806 500 -804
rect 499 -812 500 -810
rect 506 -806 507 -804
rect 506 -812 507 -810
rect 513 -806 514 -804
rect 513 -812 514 -810
rect 520 -806 521 -804
rect 520 -812 521 -810
rect 527 -806 528 -804
rect 527 -812 528 -810
rect 534 -806 535 -804
rect 534 -812 535 -810
rect 541 -806 542 -804
rect 541 -812 542 -810
rect 548 -806 549 -804
rect 551 -806 552 -804
rect 548 -812 549 -810
rect 555 -806 556 -804
rect 555 -812 556 -810
rect 562 -806 563 -804
rect 562 -812 563 -810
rect 569 -806 570 -804
rect 569 -812 570 -810
rect 576 -806 577 -804
rect 576 -812 577 -810
rect 583 -806 584 -804
rect 583 -812 584 -810
rect 590 -806 591 -804
rect 590 -812 591 -810
rect 597 -806 598 -804
rect 600 -806 601 -804
rect 597 -812 598 -810
rect 604 -806 605 -804
rect 604 -812 605 -810
rect 611 -806 612 -804
rect 611 -812 612 -810
rect 618 -806 619 -804
rect 618 -812 619 -810
rect 625 -806 626 -804
rect 625 -812 626 -810
rect 632 -806 633 -804
rect 632 -812 633 -810
rect 639 -806 640 -804
rect 639 -812 640 -810
rect 646 -806 647 -804
rect 646 -812 647 -810
rect 653 -806 654 -804
rect 653 -812 654 -810
rect 660 -806 661 -804
rect 660 -812 661 -810
rect 667 -806 668 -804
rect 667 -812 668 -810
rect 674 -806 675 -804
rect 674 -812 675 -810
rect 681 -806 682 -804
rect 681 -812 682 -810
rect 688 -806 689 -804
rect 688 -812 689 -810
rect 695 -806 696 -804
rect 695 -812 696 -810
rect 702 -806 703 -804
rect 702 -812 703 -810
rect 709 -806 710 -804
rect 709 -812 710 -810
rect 716 -806 717 -804
rect 716 -812 717 -810
rect 723 -806 724 -804
rect 723 -812 724 -810
rect 730 -806 731 -804
rect 730 -812 731 -810
rect 737 -806 738 -804
rect 737 -812 738 -810
rect 744 -806 745 -804
rect 744 -812 745 -810
rect 751 -806 752 -804
rect 751 -812 752 -810
rect 758 -806 759 -804
rect 758 -812 759 -810
rect 765 -806 766 -804
rect 765 -812 766 -810
rect 772 -806 773 -804
rect 779 -806 780 -804
rect 779 -812 780 -810
rect 786 -806 787 -804
rect 786 -812 787 -810
rect 9 -861 10 -859
rect 9 -867 10 -865
rect 19 -867 20 -865
rect 23 -861 24 -859
rect 23 -867 24 -865
rect 30 -861 31 -859
rect 30 -867 31 -865
rect 40 -867 41 -865
rect 44 -861 45 -859
rect 44 -867 45 -865
rect 51 -861 52 -859
rect 54 -867 55 -865
rect 58 -861 59 -859
rect 58 -867 59 -865
rect 65 -861 66 -859
rect 65 -867 66 -865
rect 72 -861 73 -859
rect 72 -867 73 -865
rect 79 -861 80 -859
rect 79 -867 80 -865
rect 86 -861 87 -859
rect 86 -867 87 -865
rect 93 -861 94 -859
rect 93 -867 94 -865
rect 100 -861 101 -859
rect 100 -867 101 -865
rect 107 -861 108 -859
rect 110 -861 111 -859
rect 107 -867 108 -865
rect 110 -867 111 -865
rect 114 -861 115 -859
rect 117 -861 118 -859
rect 117 -867 118 -865
rect 121 -861 122 -859
rect 121 -867 122 -865
rect 128 -861 129 -859
rect 128 -867 129 -865
rect 138 -861 139 -859
rect 135 -867 136 -865
rect 138 -867 139 -865
rect 142 -861 143 -859
rect 142 -867 143 -865
rect 149 -861 150 -859
rect 149 -867 150 -865
rect 156 -861 157 -859
rect 156 -867 157 -865
rect 163 -861 164 -859
rect 163 -867 164 -865
rect 173 -861 174 -859
rect 170 -867 171 -865
rect 173 -867 174 -865
rect 177 -861 178 -859
rect 177 -867 178 -865
rect 184 -861 185 -859
rect 184 -867 185 -865
rect 191 -861 192 -859
rect 191 -867 192 -865
rect 198 -861 199 -859
rect 198 -867 199 -865
rect 205 -861 206 -859
rect 205 -867 206 -865
rect 212 -861 213 -859
rect 212 -867 213 -865
rect 219 -861 220 -859
rect 219 -867 220 -865
rect 226 -861 227 -859
rect 226 -867 227 -865
rect 233 -861 234 -859
rect 233 -867 234 -865
rect 240 -861 241 -859
rect 240 -867 241 -865
rect 247 -861 248 -859
rect 247 -867 248 -865
rect 254 -861 255 -859
rect 254 -867 255 -865
rect 261 -861 262 -859
rect 264 -861 265 -859
rect 268 -861 269 -859
rect 271 -861 272 -859
rect 271 -867 272 -865
rect 275 -861 276 -859
rect 275 -867 276 -865
rect 282 -861 283 -859
rect 282 -867 283 -865
rect 289 -861 290 -859
rect 289 -867 290 -865
rect 296 -861 297 -859
rect 296 -867 297 -865
rect 303 -861 304 -859
rect 303 -867 304 -865
rect 310 -861 311 -859
rect 310 -867 311 -865
rect 317 -861 318 -859
rect 317 -867 318 -865
rect 324 -861 325 -859
rect 324 -867 325 -865
rect 331 -861 332 -859
rect 331 -867 332 -865
rect 338 -861 339 -859
rect 338 -867 339 -865
rect 345 -861 346 -859
rect 348 -861 349 -859
rect 348 -867 349 -865
rect 352 -861 353 -859
rect 352 -867 353 -865
rect 359 -861 360 -859
rect 359 -867 360 -865
rect 366 -861 367 -859
rect 366 -867 367 -865
rect 369 -867 370 -865
rect 373 -861 374 -859
rect 373 -867 374 -865
rect 380 -861 381 -859
rect 383 -867 384 -865
rect 387 -861 388 -859
rect 390 -861 391 -859
rect 390 -867 391 -865
rect 394 -861 395 -859
rect 394 -867 395 -865
rect 401 -861 402 -859
rect 401 -867 402 -865
rect 408 -861 409 -859
rect 408 -867 409 -865
rect 415 -861 416 -859
rect 415 -867 416 -865
rect 422 -861 423 -859
rect 422 -867 423 -865
rect 429 -861 430 -859
rect 429 -867 430 -865
rect 436 -861 437 -859
rect 436 -867 437 -865
rect 443 -861 444 -859
rect 443 -867 444 -865
rect 450 -861 451 -859
rect 450 -867 451 -865
rect 457 -861 458 -859
rect 457 -867 458 -865
rect 464 -861 465 -859
rect 464 -867 465 -865
rect 471 -861 472 -859
rect 471 -867 472 -865
rect 478 -861 479 -859
rect 478 -867 479 -865
rect 485 -861 486 -859
rect 485 -867 486 -865
rect 492 -861 493 -859
rect 492 -867 493 -865
rect 502 -861 503 -859
rect 502 -867 503 -865
rect 506 -861 507 -859
rect 506 -867 507 -865
rect 513 -861 514 -859
rect 513 -867 514 -865
rect 520 -861 521 -859
rect 520 -867 521 -865
rect 527 -861 528 -859
rect 527 -867 528 -865
rect 534 -861 535 -859
rect 534 -867 535 -865
rect 544 -861 545 -859
rect 541 -867 542 -865
rect 544 -867 545 -865
rect 548 -861 549 -859
rect 548 -867 549 -865
rect 555 -861 556 -859
rect 555 -867 556 -865
rect 562 -861 563 -859
rect 562 -867 563 -865
rect 569 -861 570 -859
rect 569 -867 570 -865
rect 576 -861 577 -859
rect 576 -867 577 -865
rect 583 -861 584 -859
rect 583 -867 584 -865
rect 590 -861 591 -859
rect 590 -867 591 -865
rect 597 -861 598 -859
rect 597 -867 598 -865
rect 607 -861 608 -859
rect 604 -867 605 -865
rect 611 -861 612 -859
rect 611 -867 612 -865
rect 618 -861 619 -859
rect 618 -867 619 -865
rect 625 -861 626 -859
rect 625 -867 626 -865
rect 632 -861 633 -859
rect 632 -867 633 -865
rect 639 -861 640 -859
rect 639 -867 640 -865
rect 646 -861 647 -859
rect 646 -867 647 -865
rect 653 -861 654 -859
rect 653 -867 654 -865
rect 660 -861 661 -859
rect 660 -867 661 -865
rect 667 -861 668 -859
rect 667 -867 668 -865
rect 681 -867 682 -865
rect 684 -867 685 -865
rect 688 -861 689 -859
rect 688 -867 689 -865
rect 695 -861 696 -859
rect 695 -867 696 -865
rect 702 -861 703 -859
rect 702 -867 703 -865
rect 726 -861 727 -859
rect 726 -867 727 -865
rect 730 -867 731 -865
rect 733 -867 734 -865
rect 737 -861 738 -859
rect 737 -867 738 -865
rect 744 -861 745 -859
rect 744 -867 745 -865
rect 751 -861 752 -859
rect 751 -867 752 -865
rect 758 -861 759 -859
rect 758 -867 759 -865
rect 44 -914 45 -912
rect 44 -920 45 -918
rect 51 -914 52 -912
rect 51 -920 52 -918
rect 58 -914 59 -912
rect 58 -920 59 -918
rect 65 -914 66 -912
rect 65 -920 66 -918
rect 72 -914 73 -912
rect 79 -914 80 -912
rect 79 -920 80 -918
rect 86 -914 87 -912
rect 86 -920 87 -918
rect 93 -914 94 -912
rect 93 -920 94 -918
rect 100 -914 101 -912
rect 100 -920 101 -918
rect 107 -914 108 -912
rect 107 -920 108 -918
rect 114 -914 115 -912
rect 114 -920 115 -918
rect 124 -914 125 -912
rect 121 -920 122 -918
rect 128 -914 129 -912
rect 128 -920 129 -918
rect 135 -914 136 -912
rect 135 -920 136 -918
rect 142 -914 143 -912
rect 142 -920 143 -918
rect 149 -914 150 -912
rect 149 -920 150 -918
rect 156 -914 157 -912
rect 156 -920 157 -918
rect 159 -920 160 -918
rect 163 -914 164 -912
rect 163 -920 164 -918
rect 170 -914 171 -912
rect 170 -920 171 -918
rect 177 -914 178 -912
rect 180 -914 181 -912
rect 184 -914 185 -912
rect 184 -920 185 -918
rect 191 -914 192 -912
rect 191 -920 192 -918
rect 198 -914 199 -912
rect 198 -920 199 -918
rect 205 -914 206 -912
rect 208 -914 209 -912
rect 205 -920 206 -918
rect 212 -914 213 -912
rect 212 -920 213 -918
rect 219 -914 220 -912
rect 219 -920 220 -918
rect 226 -914 227 -912
rect 226 -920 227 -918
rect 233 -914 234 -912
rect 233 -920 234 -918
rect 240 -914 241 -912
rect 240 -920 241 -918
rect 247 -914 248 -912
rect 247 -920 248 -918
rect 257 -914 258 -912
rect 254 -920 255 -918
rect 257 -920 258 -918
rect 261 -914 262 -912
rect 261 -920 262 -918
rect 271 -914 272 -912
rect 268 -920 269 -918
rect 275 -914 276 -912
rect 275 -920 276 -918
rect 282 -914 283 -912
rect 282 -920 283 -918
rect 289 -914 290 -912
rect 289 -920 290 -918
rect 296 -914 297 -912
rect 299 -914 300 -912
rect 299 -920 300 -918
rect 303 -914 304 -912
rect 303 -920 304 -918
rect 310 -914 311 -912
rect 310 -920 311 -918
rect 317 -914 318 -912
rect 317 -920 318 -918
rect 324 -920 325 -918
rect 331 -914 332 -912
rect 331 -920 332 -918
rect 338 -914 339 -912
rect 338 -920 339 -918
rect 345 -914 346 -912
rect 345 -920 346 -918
rect 352 -914 353 -912
rect 352 -920 353 -918
rect 359 -914 360 -912
rect 359 -920 360 -918
rect 366 -920 367 -918
rect 369 -920 370 -918
rect 373 -914 374 -912
rect 376 -914 377 -912
rect 380 -914 381 -912
rect 380 -920 381 -918
rect 387 -914 388 -912
rect 387 -920 388 -918
rect 394 -914 395 -912
rect 397 -914 398 -912
rect 401 -914 402 -912
rect 401 -920 402 -918
rect 408 -914 409 -912
rect 408 -920 409 -918
rect 415 -914 416 -912
rect 415 -920 416 -918
rect 422 -914 423 -912
rect 422 -920 423 -918
rect 429 -914 430 -912
rect 429 -920 430 -918
rect 436 -914 437 -912
rect 436 -920 437 -918
rect 443 -914 444 -912
rect 443 -920 444 -918
rect 450 -914 451 -912
rect 450 -920 451 -918
rect 457 -914 458 -912
rect 457 -920 458 -918
rect 467 -914 468 -912
rect 464 -920 465 -918
rect 471 -914 472 -912
rect 471 -920 472 -918
rect 478 -914 479 -912
rect 478 -920 479 -918
rect 485 -914 486 -912
rect 485 -920 486 -918
rect 492 -914 493 -912
rect 492 -920 493 -918
rect 499 -914 500 -912
rect 499 -920 500 -918
rect 506 -914 507 -912
rect 506 -920 507 -918
rect 513 -914 514 -912
rect 513 -920 514 -918
rect 523 -914 524 -912
rect 520 -920 521 -918
rect 527 -914 528 -912
rect 527 -920 528 -918
rect 534 -914 535 -912
rect 534 -920 535 -918
rect 541 -914 542 -912
rect 541 -920 542 -918
rect 548 -914 549 -912
rect 548 -920 549 -918
rect 555 -914 556 -912
rect 555 -920 556 -918
rect 562 -914 563 -912
rect 562 -920 563 -918
rect 569 -914 570 -912
rect 569 -920 570 -918
rect 576 -914 577 -912
rect 576 -920 577 -918
rect 583 -914 584 -912
rect 583 -920 584 -918
rect 590 -914 591 -912
rect 590 -920 591 -918
rect 597 -914 598 -912
rect 597 -920 598 -918
rect 604 -914 605 -912
rect 604 -920 605 -918
rect 611 -914 612 -912
rect 611 -920 612 -918
rect 618 -914 619 -912
rect 618 -920 619 -918
rect 625 -914 626 -912
rect 625 -920 626 -918
rect 632 -914 633 -912
rect 632 -920 633 -918
rect 642 -914 643 -912
rect 639 -920 640 -918
rect 642 -920 643 -918
rect 646 -914 647 -912
rect 646 -920 647 -918
rect 653 -920 654 -918
rect 660 -914 661 -912
rect 663 -914 664 -912
rect 667 -914 668 -912
rect 667 -920 668 -918
rect 674 -914 675 -912
rect 674 -920 675 -918
rect 681 -914 682 -912
rect 681 -920 682 -918
rect 716 -914 717 -912
rect 716 -920 717 -918
rect 747 -914 748 -912
rect 744 -920 745 -918
rect 65 -973 66 -971
rect 65 -979 66 -977
rect 72 -973 73 -971
rect 72 -979 73 -977
rect 79 -973 80 -971
rect 79 -979 80 -977
rect 86 -973 87 -971
rect 86 -979 87 -977
rect 93 -979 94 -977
rect 96 -979 97 -977
rect 103 -973 104 -971
rect 100 -979 101 -977
rect 107 -973 108 -971
rect 107 -979 108 -977
rect 117 -979 118 -977
rect 121 -973 122 -971
rect 121 -979 122 -977
rect 128 -973 129 -971
rect 128 -979 129 -977
rect 135 -973 136 -971
rect 135 -979 136 -977
rect 142 -973 143 -971
rect 142 -979 143 -977
rect 149 -973 150 -971
rect 149 -979 150 -977
rect 156 -973 157 -971
rect 156 -979 157 -977
rect 163 -973 164 -971
rect 163 -979 164 -977
rect 170 -973 171 -971
rect 170 -979 171 -977
rect 177 -973 178 -971
rect 177 -979 178 -977
rect 184 -973 185 -971
rect 184 -979 185 -977
rect 191 -973 192 -971
rect 191 -979 192 -977
rect 198 -973 199 -971
rect 201 -979 202 -977
rect 205 -973 206 -971
rect 205 -979 206 -977
rect 212 -973 213 -971
rect 212 -979 213 -977
rect 219 -973 220 -971
rect 219 -979 220 -977
rect 226 -973 227 -971
rect 226 -979 227 -977
rect 229 -979 230 -977
rect 233 -973 234 -971
rect 233 -979 234 -977
rect 240 -973 241 -971
rect 240 -979 241 -977
rect 247 -973 248 -971
rect 247 -979 248 -977
rect 254 -973 255 -971
rect 254 -979 255 -977
rect 261 -973 262 -971
rect 261 -979 262 -977
rect 268 -973 269 -971
rect 268 -979 269 -977
rect 275 -973 276 -971
rect 275 -979 276 -977
rect 282 -973 283 -971
rect 282 -979 283 -977
rect 289 -973 290 -971
rect 289 -979 290 -977
rect 296 -973 297 -971
rect 296 -979 297 -977
rect 303 -973 304 -971
rect 303 -979 304 -977
rect 313 -973 314 -971
rect 313 -979 314 -977
rect 317 -973 318 -971
rect 320 -973 321 -971
rect 324 -973 325 -971
rect 324 -979 325 -977
rect 331 -973 332 -971
rect 331 -979 332 -977
rect 338 -973 339 -971
rect 338 -979 339 -977
rect 345 -973 346 -971
rect 345 -979 346 -977
rect 352 -973 353 -971
rect 352 -979 353 -977
rect 359 -973 360 -971
rect 359 -979 360 -977
rect 366 -973 367 -971
rect 366 -979 367 -977
rect 369 -979 370 -977
rect 373 -973 374 -971
rect 373 -979 374 -977
rect 380 -973 381 -971
rect 380 -979 381 -977
rect 390 -979 391 -977
rect 394 -973 395 -971
rect 394 -979 395 -977
rect 401 -973 402 -971
rect 401 -979 402 -977
rect 408 -973 409 -971
rect 408 -979 409 -977
rect 415 -979 416 -977
rect 418 -979 419 -977
rect 425 -973 426 -971
rect 422 -979 423 -977
rect 425 -979 426 -977
rect 429 -973 430 -971
rect 429 -979 430 -977
rect 436 -973 437 -971
rect 436 -979 437 -977
rect 443 -973 444 -971
rect 443 -979 444 -977
rect 453 -973 454 -971
rect 450 -979 451 -977
rect 453 -979 454 -977
rect 457 -973 458 -971
rect 457 -979 458 -977
rect 464 -973 465 -971
rect 464 -979 465 -977
rect 471 -973 472 -971
rect 471 -979 472 -977
rect 478 -973 479 -971
rect 478 -979 479 -977
rect 485 -973 486 -971
rect 485 -979 486 -977
rect 492 -973 493 -971
rect 492 -979 493 -977
rect 499 -973 500 -971
rect 499 -979 500 -977
rect 506 -973 507 -971
rect 506 -979 507 -977
rect 513 -973 514 -971
rect 513 -979 514 -977
rect 523 -979 524 -977
rect 527 -973 528 -971
rect 527 -979 528 -977
rect 534 -973 535 -971
rect 534 -979 535 -977
rect 541 -973 542 -971
rect 544 -973 545 -971
rect 548 -973 549 -971
rect 548 -979 549 -977
rect 555 -973 556 -971
rect 555 -979 556 -977
rect 562 -973 563 -971
rect 562 -979 563 -977
rect 569 -973 570 -971
rect 569 -979 570 -977
rect 576 -973 577 -971
rect 576 -979 577 -977
rect 583 -973 584 -971
rect 583 -979 584 -977
rect 590 -973 591 -971
rect 590 -979 591 -977
rect 597 -973 598 -971
rect 597 -979 598 -977
rect 604 -973 605 -971
rect 604 -979 605 -977
rect 611 -973 612 -971
rect 611 -979 612 -977
rect 618 -973 619 -971
rect 618 -979 619 -977
rect 625 -973 626 -971
rect 628 -973 629 -971
rect 660 -973 661 -971
rect 660 -979 661 -977
rect 674 -973 675 -971
rect 674 -979 675 -977
rect 100 -1012 101 -1010
rect 100 -1018 101 -1016
rect 142 -1012 143 -1010
rect 142 -1018 143 -1016
rect 149 -1012 150 -1010
rect 149 -1018 150 -1016
rect 156 -1012 157 -1010
rect 156 -1018 157 -1016
rect 163 -1012 164 -1010
rect 163 -1018 164 -1016
rect 170 -1012 171 -1010
rect 170 -1018 171 -1016
rect 177 -1012 178 -1010
rect 177 -1018 178 -1016
rect 184 -1012 185 -1010
rect 184 -1018 185 -1016
rect 191 -1012 192 -1010
rect 191 -1018 192 -1016
rect 198 -1012 199 -1010
rect 198 -1018 199 -1016
rect 205 -1012 206 -1010
rect 205 -1018 206 -1016
rect 215 -1018 216 -1016
rect 219 -1012 220 -1010
rect 219 -1018 220 -1016
rect 226 -1012 227 -1010
rect 226 -1018 227 -1016
rect 233 -1012 234 -1010
rect 233 -1018 234 -1016
rect 240 -1012 241 -1010
rect 240 -1018 241 -1016
rect 247 -1012 248 -1010
rect 250 -1012 251 -1010
rect 247 -1018 248 -1016
rect 254 -1012 255 -1010
rect 254 -1018 255 -1016
rect 264 -1012 265 -1010
rect 261 -1018 262 -1016
rect 264 -1018 265 -1016
rect 268 -1012 269 -1010
rect 268 -1018 269 -1016
rect 275 -1012 276 -1010
rect 275 -1018 276 -1016
rect 282 -1012 283 -1010
rect 282 -1018 283 -1016
rect 289 -1012 290 -1010
rect 289 -1018 290 -1016
rect 299 -1018 300 -1016
rect 303 -1012 304 -1010
rect 303 -1018 304 -1016
rect 310 -1012 311 -1010
rect 310 -1018 311 -1016
rect 317 -1012 318 -1010
rect 317 -1018 318 -1016
rect 324 -1012 325 -1010
rect 324 -1018 325 -1016
rect 331 -1012 332 -1010
rect 338 -1012 339 -1010
rect 338 -1018 339 -1016
rect 345 -1012 346 -1010
rect 348 -1018 349 -1016
rect 352 -1012 353 -1010
rect 352 -1018 353 -1016
rect 359 -1012 360 -1010
rect 362 -1012 363 -1010
rect 359 -1018 360 -1016
rect 369 -1012 370 -1010
rect 366 -1018 367 -1016
rect 373 -1012 374 -1010
rect 373 -1018 374 -1016
rect 380 -1012 381 -1010
rect 380 -1018 381 -1016
rect 387 -1012 388 -1010
rect 387 -1018 388 -1016
rect 394 -1012 395 -1010
rect 394 -1018 395 -1016
rect 401 -1012 402 -1010
rect 401 -1018 402 -1016
rect 408 -1012 409 -1010
rect 408 -1018 409 -1016
rect 415 -1012 416 -1010
rect 415 -1018 416 -1016
rect 422 -1012 423 -1010
rect 422 -1018 423 -1016
rect 429 -1012 430 -1010
rect 436 -1012 437 -1010
rect 439 -1012 440 -1010
rect 439 -1018 440 -1016
rect 446 -1012 447 -1010
rect 443 -1018 444 -1016
rect 450 -1012 451 -1010
rect 450 -1018 451 -1016
rect 457 -1012 458 -1010
rect 460 -1018 461 -1016
rect 464 -1012 465 -1010
rect 464 -1018 465 -1016
rect 492 -1012 493 -1010
rect 492 -1018 493 -1016
rect 499 -1012 500 -1010
rect 499 -1018 500 -1016
rect 506 -1012 507 -1010
rect 506 -1018 507 -1016
rect 527 -1012 528 -1010
rect 527 -1018 528 -1016
rect 544 -1012 545 -1010
rect 548 -1012 549 -1010
rect 548 -1018 549 -1016
rect 569 -1012 570 -1010
rect 569 -1018 570 -1016
rect 576 -1012 577 -1010
rect 576 -1018 577 -1016
rect 583 -1012 584 -1010
rect 583 -1018 584 -1016
rect 590 -1012 591 -1010
rect 590 -1018 591 -1016
rect 607 -1012 608 -1010
rect 604 -1018 605 -1016
rect 611 -1012 612 -1010
rect 611 -1018 612 -1016
rect 646 -1012 647 -1010
rect 649 -1012 650 -1010
rect 670 -1012 671 -1010
rect 100 -1041 101 -1039
rect 100 -1047 101 -1045
rect 114 -1041 115 -1039
rect 114 -1047 115 -1045
rect 124 -1041 125 -1039
rect 128 -1041 129 -1039
rect 128 -1047 129 -1045
rect 135 -1041 136 -1039
rect 135 -1047 136 -1045
rect 142 -1041 143 -1039
rect 142 -1047 143 -1045
rect 149 -1041 150 -1039
rect 149 -1047 150 -1045
rect 156 -1041 157 -1039
rect 156 -1047 157 -1045
rect 163 -1041 164 -1039
rect 163 -1047 164 -1045
rect 170 -1041 171 -1039
rect 173 -1041 174 -1039
rect 173 -1047 174 -1045
rect 177 -1041 178 -1039
rect 180 -1047 181 -1045
rect 184 -1047 185 -1045
rect 191 -1041 192 -1039
rect 191 -1047 192 -1045
rect 198 -1041 199 -1039
rect 198 -1047 199 -1045
rect 205 -1041 206 -1039
rect 205 -1047 206 -1045
rect 215 -1041 216 -1039
rect 212 -1047 213 -1045
rect 219 -1041 220 -1039
rect 219 -1047 220 -1045
rect 229 -1041 230 -1039
rect 233 -1041 234 -1039
rect 233 -1047 234 -1045
rect 243 -1041 244 -1039
rect 247 -1041 248 -1039
rect 247 -1047 248 -1045
rect 254 -1041 255 -1039
rect 254 -1047 255 -1045
rect 264 -1041 265 -1039
rect 268 -1041 269 -1039
rect 268 -1047 269 -1045
rect 275 -1047 276 -1045
rect 278 -1047 279 -1045
rect 285 -1047 286 -1045
rect 289 -1041 290 -1039
rect 289 -1047 290 -1045
rect 296 -1041 297 -1039
rect 296 -1047 297 -1045
rect 306 -1041 307 -1039
rect 303 -1047 304 -1045
rect 310 -1041 311 -1039
rect 310 -1047 311 -1045
rect 317 -1041 318 -1039
rect 317 -1047 318 -1045
rect 366 -1041 367 -1039
rect 366 -1047 367 -1045
rect 373 -1041 374 -1039
rect 376 -1047 377 -1045
rect 383 -1047 384 -1045
rect 387 -1041 388 -1039
rect 387 -1047 388 -1045
rect 394 -1041 395 -1039
rect 394 -1047 395 -1045
rect 404 -1047 405 -1045
rect 408 -1041 409 -1039
rect 408 -1047 409 -1045
rect 418 -1041 419 -1039
rect 415 -1047 416 -1045
rect 422 -1041 423 -1039
rect 422 -1047 423 -1045
rect 429 -1041 430 -1039
rect 429 -1047 430 -1045
rect 436 -1041 437 -1039
rect 436 -1047 437 -1045
rect 443 -1041 444 -1039
rect 443 -1047 444 -1045
rect 457 -1041 458 -1039
rect 457 -1047 458 -1045
rect 474 -1041 475 -1039
rect 471 -1047 472 -1045
rect 478 -1041 479 -1039
rect 478 -1047 479 -1045
rect 485 -1041 486 -1039
rect 485 -1047 486 -1045
rect 541 -1047 542 -1045
rect 548 -1041 549 -1039
rect 548 -1047 549 -1045
rect 562 -1041 563 -1039
rect 562 -1047 563 -1045
rect 569 -1041 570 -1039
rect 569 -1047 570 -1045
rect 579 -1047 580 -1045
rect 583 -1041 584 -1039
rect 583 -1047 584 -1045
rect 590 -1041 591 -1039
rect 590 -1047 591 -1045
rect 100 -1068 101 -1066
rect 107 -1062 108 -1060
rect 107 -1068 108 -1066
rect 135 -1062 136 -1060
rect 142 -1062 143 -1060
rect 149 -1062 150 -1060
rect 149 -1068 150 -1066
rect 159 -1068 160 -1066
rect 163 -1062 164 -1060
rect 163 -1068 164 -1066
rect 170 -1068 171 -1066
rect 194 -1062 195 -1060
rect 198 -1062 199 -1060
rect 198 -1068 199 -1066
rect 205 -1068 206 -1066
rect 215 -1068 216 -1066
rect 219 -1068 220 -1066
rect 226 -1062 227 -1060
rect 226 -1068 227 -1066
rect 233 -1062 234 -1060
rect 233 -1068 234 -1066
rect 282 -1062 283 -1060
rect 296 -1062 297 -1060
rect 299 -1062 300 -1060
rect 380 -1062 381 -1060
rect 380 -1068 381 -1066
rect 394 -1068 395 -1066
rect 411 -1062 412 -1060
rect 429 -1062 430 -1060
rect 429 -1068 430 -1066
rect 439 -1068 440 -1066
rect 443 -1062 444 -1060
rect 446 -1068 447 -1066
rect 453 -1062 454 -1060
rect 457 -1062 458 -1060
rect 457 -1068 458 -1066
rect 562 -1062 563 -1060
rect 579 -1062 580 -1060
rect 576 -1068 577 -1066
rect 583 -1062 584 -1060
rect 583 -1068 584 -1066
<< metal1 >>
rect 114 0 122 1
rect 128 0 150 1
rect 156 0 167 1
rect 177 0 199 1
rect 236 0 248 1
rect 296 0 314 1
rect 317 0 374 1
rect 131 -2 164 -1
rect 191 -2 209 -1
rect 331 -2 339 -1
rect 348 -2 353 -1
rect 135 -4 143 -3
rect 72 -15 90 -14
rect 100 -15 129 -14
rect 131 -15 150 -14
rect 156 -15 185 -14
rect 187 -15 237 -14
rect 247 -15 255 -14
rect 296 -15 304 -14
rect 331 -15 346 -14
rect 373 -15 437 -14
rect 485 -15 556 -14
rect 79 -17 97 -16
rect 107 -17 136 -16
rect 142 -17 192 -16
rect 201 -17 213 -16
rect 215 -17 234 -16
rect 296 -17 318 -16
rect 394 -17 405 -16
rect 422 -17 430 -16
rect 117 -19 122 -18
rect 135 -19 160 -18
rect 170 -19 178 -18
rect 184 -19 199 -18
rect 219 -19 283 -18
rect 313 -19 332 -18
rect 156 -21 192 -20
rect 229 -21 241 -20
rect 173 -23 178 -22
rect 51 -34 59 -33
rect 65 -34 69 -33
rect 79 -34 94 -33
rect 96 -34 115 -33
rect 149 -34 164 -33
rect 166 -34 171 -33
rect 191 -34 227 -33
rect 233 -34 269 -33
rect 275 -34 318 -33
rect 345 -34 367 -33
rect 387 -34 395 -33
rect 415 -34 489 -33
rect 555 -34 577 -33
rect 65 -36 73 -35
rect 86 -36 101 -35
rect 107 -36 171 -35
rect 212 -36 220 -35
rect 233 -36 251 -35
rect 254 -36 265 -35
rect 285 -36 339 -35
rect 352 -36 374 -35
rect 380 -36 395 -35
rect 429 -36 444 -35
rect 68 -38 73 -37
rect 100 -38 118 -37
rect 149 -38 206 -37
rect 240 -38 248 -37
rect 289 -38 314 -37
rect 327 -38 346 -37
rect 359 -38 405 -37
rect 436 -38 451 -37
rect 107 -40 223 -39
rect 303 -40 325 -39
rect 331 -40 353 -39
rect 156 -42 199 -41
rect 254 -42 304 -41
rect 159 -44 178 -43
rect 194 -44 206 -43
rect 282 -44 332 -43
rect 121 -46 160 -45
rect 177 -46 227 -45
rect 121 -48 136 -47
rect 135 -50 143 -49
rect 142 -52 216 -51
rect 30 -63 153 -62
rect 156 -63 171 -62
rect 191 -63 269 -62
rect 366 -63 409 -62
rect 425 -63 465 -62
rect 471 -63 528 -62
rect 530 -63 591 -62
rect 37 -65 52 -64
rect 58 -65 83 -64
rect 93 -65 227 -64
rect 233 -65 269 -64
rect 373 -65 430 -64
rect 443 -65 493 -64
rect 44 -67 136 -66
rect 142 -67 213 -66
rect 240 -67 248 -66
rect 261 -67 286 -66
rect 303 -67 374 -66
rect 380 -67 388 -66
rect 401 -67 479 -66
rect 51 -69 122 -68
rect 131 -69 171 -68
rect 205 -69 234 -68
rect 240 -69 255 -68
rect 261 -69 290 -68
rect 387 -69 395 -68
rect 401 -69 416 -68
rect 65 -71 97 -70
rect 100 -71 178 -70
rect 289 -71 360 -70
rect 72 -73 80 -72
rect 86 -73 101 -72
rect 128 -73 178 -72
rect 324 -73 416 -72
rect 65 -75 87 -74
rect 128 -75 248 -74
rect 313 -75 325 -74
rect 331 -75 395 -74
rect 72 -77 216 -76
rect 296 -77 332 -76
rect 345 -77 360 -76
rect 131 -79 136 -78
rect 142 -79 185 -78
rect 219 -79 297 -78
rect 313 -79 437 -78
rect 149 -81 192 -80
rect 219 -81 244 -80
rect 345 -81 370 -80
rect 163 -83 206 -82
rect 163 -85 230 -84
rect 184 -87 276 -86
rect 275 -89 339 -88
rect 338 -91 353 -90
rect 9 -102 38 -101
rect 51 -102 122 -101
rect 128 -102 258 -101
rect 282 -102 528 -101
rect 555 -102 577 -101
rect 590 -102 619 -101
rect 16 -104 59 -103
rect 65 -104 101 -103
rect 121 -104 157 -103
rect 170 -104 314 -103
rect 331 -104 458 -103
rect 460 -104 591 -103
rect 26 -106 69 -105
rect 75 -106 157 -105
rect 173 -106 192 -105
rect 240 -106 563 -105
rect 30 -108 94 -107
rect 100 -108 108 -107
rect 149 -108 241 -107
rect 243 -108 269 -107
rect 282 -108 290 -107
rect 313 -108 360 -107
rect 366 -108 570 -107
rect 37 -110 80 -109
rect 86 -110 150 -109
rect 191 -110 199 -109
rect 226 -110 269 -109
rect 275 -110 290 -109
rect 338 -110 360 -109
rect 366 -110 451 -109
rect 478 -110 577 -109
rect 30 -112 276 -111
rect 345 -112 353 -111
rect 355 -112 605 -111
rect 51 -114 97 -113
rect 107 -114 115 -113
rect 142 -114 339 -113
rect 345 -114 402 -113
rect 415 -114 535 -113
rect 58 -116 87 -115
rect 114 -116 125 -115
rect 142 -116 164 -115
rect 198 -116 213 -115
rect 226 -116 447 -115
rect 492 -116 612 -115
rect 205 -118 213 -117
rect 233 -118 402 -117
rect 415 -118 493 -117
rect 499 -118 507 -117
rect 520 -118 524 -117
rect 135 -120 234 -119
rect 247 -120 549 -119
rect 44 -122 136 -121
rect 205 -122 220 -121
rect 247 -122 304 -121
rect 373 -122 514 -121
rect 44 -124 73 -123
rect 184 -124 304 -123
rect 320 -124 374 -123
rect 387 -124 451 -123
rect 72 -126 332 -125
rect 394 -126 598 -125
rect 159 -128 185 -127
rect 219 -128 223 -127
rect 261 -128 321 -127
rect 324 -128 388 -127
rect 422 -128 465 -127
rect 170 -130 262 -129
rect 296 -130 395 -129
rect 408 -130 465 -129
rect 177 -132 297 -131
rect 310 -132 325 -131
rect 408 -132 472 -131
rect 166 -134 178 -133
rect 429 -134 479 -133
rect 429 -136 475 -135
rect 436 -138 486 -137
rect 380 -140 437 -139
rect 443 -140 542 -139
rect 257 -142 381 -141
rect 443 -142 587 -141
rect 23 -153 192 -152
rect 205 -153 258 -152
rect 261 -153 570 -152
rect 611 -153 661 -152
rect 51 -155 181 -154
rect 184 -155 419 -154
rect 464 -155 640 -154
rect 51 -157 129 -156
rect 142 -157 185 -156
rect 191 -157 293 -156
rect 306 -157 598 -156
rect 618 -157 626 -156
rect 628 -157 647 -156
rect 65 -159 94 -158
rect 100 -159 129 -158
rect 135 -159 143 -158
rect 156 -159 164 -158
rect 173 -159 199 -158
rect 212 -159 311 -158
rect 313 -159 591 -158
rect 604 -159 626 -158
rect 58 -161 66 -160
rect 72 -161 139 -160
rect 198 -161 248 -160
rect 254 -161 297 -160
rect 334 -161 668 -160
rect 16 -163 59 -162
rect 79 -163 157 -162
rect 212 -163 262 -162
rect 278 -163 535 -162
rect 541 -163 570 -162
rect 576 -163 591 -162
rect 16 -165 45 -164
rect 79 -165 108 -164
rect 135 -165 300 -164
rect 387 -165 675 -164
rect 44 -167 283 -166
rect 289 -167 325 -166
rect 387 -167 619 -166
rect 82 -169 97 -168
rect 100 -169 402 -168
rect 436 -169 465 -168
rect 471 -169 598 -168
rect 86 -171 150 -170
rect 215 -171 395 -170
rect 457 -171 535 -170
rect 562 -171 605 -170
rect 86 -173 115 -172
rect 149 -173 528 -172
rect 555 -173 563 -172
rect 107 -175 122 -174
rect 219 -175 339 -174
rect 341 -175 472 -174
rect 485 -175 633 -174
rect 30 -177 220 -176
rect 247 -177 587 -176
rect 30 -179 241 -178
rect 268 -179 395 -178
rect 422 -179 458 -178
rect 492 -179 612 -178
rect 37 -181 122 -180
rect 222 -181 423 -180
rect 499 -181 514 -180
rect 520 -181 542 -180
rect 37 -183 97 -182
rect 114 -183 227 -182
rect 240 -183 279 -182
rect 282 -183 370 -182
rect 390 -183 654 -182
rect 177 -185 227 -184
rect 296 -185 381 -184
rect 488 -185 514 -184
rect 520 -185 584 -184
rect 177 -187 209 -186
rect 317 -187 556 -186
rect 268 -189 318 -188
rect 320 -189 437 -188
rect 506 -189 528 -188
rect 548 -189 584 -188
rect 359 -191 493 -190
rect 331 -193 360 -192
rect 366 -193 402 -192
rect 415 -193 549 -192
rect 331 -195 577 -194
rect 345 -197 416 -196
rect 478 -197 507 -196
rect 170 -199 346 -198
rect 373 -199 381 -198
rect 408 -199 479 -198
rect 9 -201 171 -200
rect 352 -201 374 -200
rect 408 -201 430 -200
rect 303 -203 353 -202
rect 429 -203 444 -202
rect 23 -214 213 -213
rect 275 -214 535 -213
rect 548 -214 689 -213
rect 23 -216 97 -215
rect 100 -216 108 -215
rect 152 -216 244 -215
rect 292 -216 535 -215
rect 548 -216 598 -215
rect 653 -216 696 -215
rect 44 -218 94 -217
rect 103 -218 234 -217
rect 296 -218 430 -217
rect 446 -218 598 -217
rect 660 -218 717 -217
rect 44 -220 55 -219
rect 65 -220 76 -219
rect 86 -220 136 -219
rect 156 -220 279 -219
rect 303 -220 353 -219
rect 369 -220 619 -219
rect 51 -222 73 -221
rect 86 -222 279 -221
rect 313 -222 570 -221
rect 583 -222 619 -221
rect 51 -224 150 -223
rect 170 -224 325 -223
rect 331 -224 640 -223
rect 37 -226 332 -225
rect 338 -226 360 -225
rect 369 -226 570 -225
rect 590 -226 654 -225
rect 9 -228 38 -227
rect 65 -228 83 -227
rect 128 -228 157 -227
rect 177 -228 311 -227
rect 341 -228 493 -227
rect 499 -228 591 -227
rect 611 -228 661 -227
rect 16 -230 178 -229
rect 191 -230 206 -229
rect 233 -230 241 -229
rect 254 -230 353 -229
rect 387 -230 633 -229
rect 16 -232 118 -231
rect 128 -232 185 -231
rect 191 -232 227 -231
rect 254 -232 269 -231
rect 299 -232 640 -231
rect 30 -234 311 -233
rect 345 -234 360 -233
rect 422 -234 724 -233
rect 33 -236 227 -235
rect 247 -236 346 -235
rect 408 -236 423 -235
rect 457 -236 486 -235
rect 488 -236 605 -235
rect 79 -238 171 -237
rect 198 -238 202 -237
rect 247 -238 682 -237
rect 2 -240 80 -239
rect 107 -240 388 -239
rect 464 -240 493 -239
rect 513 -240 703 -239
rect 121 -242 185 -241
rect 198 -242 290 -241
rect 299 -242 430 -241
rect 471 -242 500 -241
rect 513 -242 675 -241
rect 121 -244 265 -243
rect 268 -244 283 -243
rect 327 -244 458 -243
rect 471 -244 479 -243
rect 527 -244 584 -243
rect 135 -246 181 -245
rect 201 -246 290 -245
rect 366 -246 528 -245
rect 555 -246 605 -245
rect 250 -248 556 -247
rect 562 -248 633 -247
rect 261 -250 283 -249
rect 380 -250 409 -249
rect 436 -250 479 -249
rect 506 -250 563 -249
rect 576 -250 612 -249
rect 380 -252 647 -251
rect 383 -254 675 -253
rect 394 -256 437 -255
rect 506 -256 668 -255
rect 394 -258 402 -257
rect 541 -258 577 -257
rect 625 -258 668 -257
rect 373 -260 402 -259
rect 415 -260 542 -259
rect 646 -260 713 -259
rect 30 -262 374 -261
rect 443 -262 626 -261
rect 317 -264 416 -263
rect 443 -264 451 -263
rect 114 -266 318 -265
rect 450 -266 521 -265
rect 520 -268 731 -267
rect 23 -279 55 -278
rect 58 -279 111 -278
rect 128 -279 279 -278
rect 289 -279 353 -278
rect 362 -279 542 -278
rect 569 -279 731 -278
rect 26 -281 227 -280
rect 240 -281 528 -280
rect 534 -281 570 -280
rect 716 -281 738 -280
rect 2 -283 227 -282
rect 247 -283 304 -282
rect 310 -283 339 -282
rect 345 -283 353 -282
rect 380 -283 640 -282
rect 30 -285 73 -284
rect 82 -285 668 -284
rect 16 -287 73 -286
rect 86 -287 304 -286
rect 310 -287 314 -286
rect 338 -287 416 -286
rect 422 -287 465 -286
rect 467 -287 549 -286
rect 639 -287 654 -286
rect 667 -287 682 -286
rect 16 -289 206 -288
rect 212 -289 251 -288
rect 292 -289 717 -288
rect 33 -291 535 -290
rect 541 -291 591 -290
rect 653 -291 675 -290
rect 37 -293 80 -292
rect 100 -293 171 -292
rect 198 -293 349 -292
rect 380 -293 402 -292
rect 422 -293 507 -292
rect 548 -293 563 -292
rect 590 -293 612 -292
rect 44 -295 528 -294
rect 555 -295 682 -294
rect 47 -297 437 -296
rect 499 -297 507 -296
rect 555 -297 598 -296
rect 51 -299 87 -298
rect 107 -299 206 -298
rect 212 -299 384 -298
rect 394 -299 416 -298
rect 432 -299 521 -298
rect 562 -299 584 -298
rect 597 -299 626 -298
rect 54 -301 115 -300
rect 121 -301 129 -300
rect 135 -301 150 -300
rect 156 -301 241 -300
rect 257 -301 612 -300
rect 625 -301 633 -300
rect 58 -303 297 -302
rect 345 -303 703 -302
rect 65 -305 188 -304
rect 191 -305 199 -304
rect 219 -305 248 -304
rect 261 -305 675 -304
rect 65 -307 269 -306
rect 299 -307 703 -306
rect 93 -309 269 -308
rect 299 -309 514 -308
rect 583 -309 619 -308
rect 632 -309 647 -308
rect 110 -311 115 -310
rect 121 -311 370 -310
rect 394 -311 409 -310
rect 436 -311 710 -310
rect 135 -313 185 -312
rect 191 -313 283 -312
rect 401 -313 724 -312
rect 37 -315 185 -314
rect 275 -315 619 -314
rect 646 -315 661 -314
rect 695 -315 724 -314
rect 44 -317 696 -316
rect 93 -319 283 -318
rect 443 -319 500 -318
rect 660 -319 689 -318
rect 142 -321 171 -320
rect 177 -321 262 -320
rect 275 -321 409 -320
rect 457 -321 521 -320
rect 142 -323 265 -322
rect 324 -323 458 -322
rect 471 -323 514 -322
rect 156 -325 234 -324
rect 324 -325 388 -324
rect 450 -325 472 -324
rect 51 -327 234 -326
rect 278 -327 388 -326
rect 429 -327 451 -326
rect 163 -329 220 -328
rect 327 -329 689 -328
rect 177 -331 255 -330
rect 331 -331 444 -330
rect 317 -333 332 -332
rect 429 -333 710 -332
rect 317 -335 360 -334
rect 5 -346 360 -345
rect 369 -346 479 -345
rect 555 -346 759 -345
rect 23 -348 367 -347
rect 376 -348 801 -347
rect 26 -350 451 -349
rect 474 -350 766 -349
rect 30 -352 185 -351
rect 187 -352 248 -351
rect 268 -352 279 -351
rect 282 -352 570 -351
rect 667 -352 745 -351
rect 30 -354 157 -353
rect 219 -354 255 -353
rect 268 -354 458 -353
rect 513 -354 570 -353
rect 583 -354 668 -353
rect 674 -354 752 -353
rect 2 -356 584 -355
rect 688 -356 773 -355
rect 44 -358 398 -357
rect 408 -358 458 -357
rect 464 -358 514 -357
rect 527 -358 675 -357
rect 695 -358 780 -357
rect 47 -360 297 -359
rect 324 -360 346 -359
rect 352 -360 367 -359
rect 408 -360 416 -359
rect 432 -360 724 -359
rect 730 -360 808 -359
rect 51 -362 192 -361
rect 219 -362 444 -361
rect 485 -362 528 -361
rect 558 -362 815 -361
rect 54 -364 405 -363
rect 415 -364 738 -363
rect 61 -366 230 -365
rect 233 -366 419 -365
rect 422 -366 444 -365
rect 471 -366 486 -365
rect 618 -366 689 -365
rect 709 -366 787 -365
rect 72 -368 234 -367
rect 247 -368 339 -367
rect 345 -368 703 -367
rect 716 -368 794 -367
rect 72 -370 87 -369
rect 93 -370 276 -369
rect 282 -370 332 -369
rect 338 -370 451 -369
rect 625 -370 696 -369
rect 37 -372 332 -371
rect 348 -372 724 -371
rect 79 -374 192 -373
rect 226 -374 353 -373
rect 387 -374 423 -373
rect 429 -374 619 -373
rect 639 -374 703 -373
rect 79 -376 178 -375
rect 226 -376 318 -375
rect 348 -376 738 -375
rect 86 -378 136 -377
rect 285 -378 524 -377
rect 541 -378 640 -377
rect 646 -378 710 -377
rect 93 -380 342 -379
rect 436 -380 479 -379
rect 492 -380 542 -379
rect 576 -380 626 -379
rect 646 -380 661 -379
rect 681 -380 731 -379
rect 100 -382 136 -381
rect 289 -382 388 -381
rect 394 -382 437 -381
rect 492 -382 500 -381
rect 520 -382 577 -381
rect 590 -382 661 -381
rect 100 -384 206 -383
rect 292 -384 465 -383
rect 590 -384 598 -383
rect 611 -384 682 -383
rect 107 -386 633 -385
rect 653 -386 717 -385
rect 110 -388 255 -387
rect 296 -388 304 -387
rect 310 -388 318 -387
rect 534 -388 598 -387
rect 604 -388 612 -387
rect 110 -390 500 -389
rect 548 -390 654 -389
rect 121 -392 206 -391
rect 222 -392 311 -391
rect 383 -392 605 -391
rect 124 -394 157 -393
rect 163 -394 290 -393
rect 299 -394 633 -393
rect 114 -396 164 -395
rect 303 -396 335 -395
rect 401 -396 535 -395
rect 37 -398 402 -397
rect 506 -398 549 -397
rect 114 -400 241 -399
rect 128 -402 178 -401
rect 240 -402 381 -401
rect 128 -404 143 -403
rect 212 -404 381 -403
rect 16 -406 213 -405
rect 16 -408 199 -407
rect 142 -410 171 -409
rect 198 -410 395 -409
rect 65 -412 171 -411
rect 58 -414 66 -413
rect 9 -425 52 -424
rect 58 -425 69 -424
rect 72 -425 139 -424
rect 170 -425 220 -424
rect 264 -425 752 -424
rect 9 -427 45 -426
rect 47 -427 668 -426
rect 702 -427 706 -426
rect 51 -429 101 -428
rect 107 -429 675 -428
rect 702 -429 745 -428
rect 58 -431 759 -430
rect 61 -433 269 -432
rect 275 -433 374 -432
rect 380 -433 661 -432
rect 730 -433 745 -432
rect 72 -435 199 -434
rect 205 -435 290 -434
rect 334 -435 598 -434
rect 611 -435 675 -434
rect 716 -435 731 -434
rect 79 -437 276 -436
rect 338 -437 654 -436
rect 79 -439 297 -438
rect 348 -439 724 -438
rect 86 -441 122 -440
rect 163 -441 206 -440
rect 233 -441 339 -440
rect 366 -441 384 -440
rect 394 -441 640 -440
rect 646 -441 759 -440
rect 44 -443 234 -442
rect 254 -443 297 -442
rect 387 -443 395 -442
rect 401 -443 633 -442
rect 709 -443 724 -442
rect 86 -445 360 -444
rect 404 -445 794 -444
rect 93 -447 164 -446
rect 170 -447 223 -446
rect 226 -447 367 -446
rect 443 -447 612 -446
rect 618 -447 640 -446
rect 695 -447 710 -446
rect 793 -447 808 -446
rect 93 -449 346 -448
rect 352 -449 360 -448
rect 474 -449 773 -448
rect 100 -451 405 -450
rect 474 -451 661 -450
rect 681 -451 696 -450
rect 772 -451 787 -450
rect 107 -453 129 -452
rect 198 -453 318 -452
rect 324 -453 346 -452
rect 355 -453 619 -452
rect 625 -453 647 -452
rect 786 -453 801 -452
rect 30 -455 129 -454
rect 191 -455 325 -454
rect 506 -455 598 -454
rect 604 -455 633 -454
rect 800 -455 815 -454
rect 30 -457 433 -456
rect 520 -457 738 -456
rect 37 -459 507 -458
rect 523 -459 766 -458
rect 37 -461 150 -460
rect 212 -461 255 -460
rect 261 -461 269 -460
rect 303 -461 318 -460
rect 418 -461 521 -460
rect 541 -461 545 -460
rect 558 -461 752 -460
rect 765 -461 780 -460
rect 110 -463 192 -462
rect 222 -463 780 -462
rect 135 -465 213 -464
rect 247 -465 444 -464
rect 541 -465 584 -464
rect 590 -465 682 -464
rect 688 -465 738 -464
rect 149 -467 384 -466
rect 562 -467 654 -466
rect 705 -467 717 -466
rect 247 -469 283 -468
rect 303 -469 465 -468
rect 492 -469 563 -468
rect 569 -469 591 -468
rect 282 -471 311 -470
rect 380 -471 689 -470
rect 16 -473 311 -472
rect 422 -473 465 -472
rect 492 -473 668 -472
rect 16 -475 125 -474
rect 422 -475 479 -474
rect 548 -475 570 -474
rect 576 -475 605 -474
rect 415 -477 479 -476
rect 527 -477 549 -476
rect 555 -477 577 -476
rect 408 -479 416 -478
rect 485 -479 528 -478
rect 485 -481 535 -480
rect 457 -483 535 -482
rect 457 -485 514 -484
rect 499 -487 514 -486
rect 331 -489 500 -488
rect 156 -491 332 -490
rect 156 -493 185 -492
rect 142 -495 185 -494
rect 142 -497 178 -496
rect 23 -499 178 -498
rect 23 -501 241 -500
rect 65 -503 241 -502
rect 65 -505 115 -504
rect 114 -507 472 -506
rect 9 -518 104 -517
rect 163 -518 433 -517
rect 467 -518 773 -517
rect 793 -518 808 -517
rect 9 -520 101 -519
rect 163 -520 178 -519
rect 184 -520 220 -519
rect 222 -520 535 -519
rect 555 -520 577 -519
rect 583 -520 822 -519
rect 16 -522 265 -521
rect 313 -522 360 -521
rect 380 -522 559 -521
rect 618 -522 622 -521
rect 779 -522 794 -521
rect 800 -522 815 -521
rect 16 -524 451 -523
rect 471 -524 493 -523
rect 495 -524 703 -523
rect 758 -524 780 -523
rect 786 -524 801 -523
rect 44 -526 111 -525
rect 135 -526 451 -525
rect 457 -526 493 -525
rect 520 -526 535 -525
rect 541 -526 584 -525
rect 618 -526 654 -525
rect 744 -526 759 -525
rect 765 -526 787 -525
rect 47 -528 332 -527
rect 383 -528 549 -527
rect 621 -528 654 -527
rect 54 -530 192 -529
rect 226 -530 276 -529
rect 303 -530 314 -529
rect 317 -530 332 -529
rect 383 -530 563 -529
rect 625 -530 745 -529
rect 58 -532 94 -531
rect 131 -532 192 -531
rect 212 -532 227 -531
rect 233 -532 360 -531
rect 387 -532 773 -531
rect 61 -534 101 -533
rect 121 -534 234 -533
rect 240 -534 388 -533
rect 390 -534 514 -533
rect 520 -534 528 -533
rect 541 -534 591 -533
rect 625 -534 640 -533
rect 79 -536 220 -535
rect 240 -536 374 -535
rect 394 -536 409 -535
rect 429 -536 731 -535
rect 79 -538 206 -537
rect 257 -538 283 -537
rect 310 -538 766 -537
rect 51 -540 206 -539
rect 275 -540 307 -539
rect 345 -540 374 -539
rect 401 -540 577 -539
rect 639 -540 661 -539
rect 30 -542 346 -541
rect 401 -542 416 -541
rect 422 -542 430 -541
rect 457 -542 717 -541
rect 30 -544 199 -543
rect 282 -544 507 -543
rect 562 -544 598 -543
rect 86 -546 353 -545
rect 369 -546 717 -545
rect 86 -548 262 -547
rect 317 -548 661 -547
rect 93 -550 171 -549
rect 177 -550 269 -549
rect 415 -550 612 -549
rect 114 -552 395 -551
rect 422 -552 437 -551
rect 474 -552 570 -551
rect 597 -552 633 -551
rect 23 -554 115 -553
rect 135 -554 269 -553
rect 436 -554 465 -553
rect 478 -554 552 -553
rect 569 -554 605 -553
rect 611 -554 724 -553
rect 23 -556 325 -555
rect 411 -556 724 -555
rect 149 -558 262 -557
rect 324 -558 339 -557
rect 443 -558 479 -557
rect 485 -558 528 -557
rect 604 -558 675 -557
rect 72 -560 444 -559
rect 488 -560 703 -559
rect 142 -562 150 -561
rect 156 -562 213 -561
rect 296 -562 339 -561
rect 499 -562 731 -561
rect 37 -564 157 -563
rect 170 -564 290 -563
rect 464 -564 500 -563
rect 506 -564 591 -563
rect 632 -564 647 -563
rect 674 -564 752 -563
rect 37 -566 108 -565
rect 198 -566 367 -565
rect 646 -566 668 -565
rect 737 -566 752 -565
rect 65 -568 143 -567
rect 289 -568 486 -567
rect 667 -568 689 -567
rect 65 -570 248 -569
rect 418 -570 738 -569
rect 128 -572 367 -571
rect 688 -572 696 -571
rect 72 -574 129 -573
rect 247 -574 255 -573
rect 334 -574 696 -573
rect 184 -576 255 -575
rect 2 -587 73 -586
rect 107 -587 157 -586
rect 163 -587 370 -586
rect 457 -587 556 -586
rect 9 -589 293 -588
rect 296 -589 395 -588
rect 464 -589 510 -588
rect 513 -589 633 -588
rect 9 -591 332 -590
rect 334 -591 731 -590
rect 54 -593 346 -592
rect 467 -593 577 -592
rect 730 -593 808 -592
rect 68 -595 283 -594
rect 299 -595 367 -594
rect 485 -595 682 -594
rect 72 -597 101 -596
rect 107 -597 745 -596
rect 100 -599 461 -598
rect 506 -599 654 -598
rect 110 -601 185 -600
rect 205 -601 258 -600
rect 271 -601 395 -600
rect 460 -601 682 -600
rect 110 -603 241 -602
rect 254 -603 633 -602
rect 653 -603 738 -602
rect 121 -605 409 -604
rect 506 -605 542 -604
rect 576 -605 612 -604
rect 737 -605 794 -604
rect 121 -607 178 -606
rect 184 -607 479 -606
rect 513 -607 563 -606
rect 611 -607 689 -606
rect 26 -609 689 -608
rect 124 -611 773 -610
rect 128 -613 171 -612
rect 177 -613 290 -612
rect 303 -613 318 -612
rect 320 -613 409 -612
rect 478 -613 493 -612
rect 534 -613 556 -612
rect 562 -613 619 -612
rect 772 -613 801 -612
rect 138 -615 143 -614
rect 149 -615 318 -614
rect 331 -615 374 -614
rect 492 -615 528 -614
rect 534 -615 591 -614
rect 618 -615 703 -614
rect 37 -617 143 -616
rect 156 -617 297 -616
rect 303 -617 360 -616
rect 366 -617 815 -616
rect 30 -619 38 -618
rect 61 -619 150 -618
rect 163 -619 227 -618
rect 240 -619 248 -618
rect 282 -619 325 -618
rect 359 -619 423 -618
rect 527 -619 584 -618
rect 590 -619 661 -618
rect 702 -619 752 -618
rect 170 -621 230 -620
rect 289 -621 486 -620
rect 583 -621 605 -620
rect 751 -621 787 -620
rect 191 -623 255 -622
rect 310 -623 626 -622
rect 191 -625 346 -624
rect 348 -625 661 -624
rect 205 -627 234 -626
rect 275 -627 311 -626
rect 324 -627 353 -626
rect 373 -627 444 -626
rect 453 -627 787 -626
rect 198 -629 234 -628
rect 268 -629 276 -628
rect 338 -629 353 -628
rect 422 -629 430 -628
rect 443 -629 517 -628
rect 548 -629 605 -628
rect 625 -629 710 -628
rect 65 -631 199 -630
rect 212 -631 269 -630
rect 338 -631 388 -630
rect 548 -631 598 -630
rect 709 -631 780 -630
rect 30 -633 213 -632
rect 215 -633 724 -632
rect 758 -633 780 -632
rect 219 -635 248 -634
rect 380 -635 724 -634
rect 758 -635 794 -634
rect 51 -637 220 -636
rect 226 -637 262 -636
rect 383 -637 430 -636
rect 597 -637 668 -636
rect 44 -639 262 -638
rect 383 -639 465 -638
rect 646 -639 668 -638
rect 44 -641 314 -640
rect 387 -641 402 -640
rect 646 -641 696 -640
rect 16 -643 402 -642
rect 499 -643 696 -642
rect 16 -645 59 -644
rect 499 -645 640 -644
rect 58 -647 136 -646
rect 639 -647 717 -646
rect 79 -649 136 -648
rect 674 -649 717 -648
rect 79 -651 115 -650
rect 674 -651 766 -650
rect 23 -653 115 -652
rect 415 -653 766 -652
rect 23 -655 451 -654
rect 415 -657 745 -656
rect 450 -659 472 -658
rect 471 -661 521 -660
rect 520 -663 570 -662
rect 569 -665 822 -664
rect 2 -676 90 -675
rect 142 -676 419 -675
rect 425 -676 507 -675
rect 520 -676 524 -675
rect 551 -676 661 -675
rect 779 -676 787 -675
rect 16 -678 69 -677
rect 142 -678 164 -677
rect 184 -678 349 -677
rect 415 -678 437 -677
rect 446 -678 528 -677
rect 660 -678 675 -677
rect 779 -678 808 -677
rect 16 -680 94 -679
rect 107 -680 437 -679
rect 450 -680 486 -679
rect 499 -680 503 -679
rect 527 -680 710 -679
rect 51 -682 87 -681
rect 107 -682 269 -681
rect 271 -682 668 -681
rect 37 -684 52 -683
rect 58 -684 122 -683
rect 149 -684 185 -683
rect 212 -684 318 -683
rect 415 -684 430 -683
rect 453 -684 654 -683
rect 9 -686 318 -685
rect 457 -686 465 -685
rect 471 -686 801 -685
rect 37 -688 80 -687
rect 93 -688 272 -687
rect 296 -688 773 -687
rect 61 -690 171 -689
rect 198 -690 297 -689
rect 310 -690 430 -689
rect 443 -690 472 -689
rect 485 -690 493 -689
rect 499 -690 514 -689
rect 604 -690 668 -689
rect 772 -690 794 -689
rect 12 -692 311 -691
rect 443 -692 738 -691
rect 68 -694 80 -693
rect 114 -694 122 -693
rect 135 -694 150 -693
rect 170 -694 262 -693
rect 268 -694 367 -693
rect 460 -694 738 -693
rect 72 -696 164 -695
rect 198 -696 241 -695
rect 261 -696 304 -695
rect 464 -696 535 -695
rect 583 -696 605 -695
rect 646 -696 675 -695
rect 23 -698 73 -697
rect 114 -698 129 -697
rect 135 -698 230 -697
rect 233 -698 290 -697
rect 303 -698 370 -697
rect 492 -698 570 -697
rect 583 -698 612 -697
rect 646 -698 703 -697
rect 23 -700 192 -699
rect 212 -700 255 -699
rect 513 -700 556 -699
rect 590 -700 612 -699
rect 618 -700 703 -699
rect 44 -702 129 -701
rect 191 -702 206 -701
rect 226 -702 710 -701
rect 44 -704 66 -703
rect 205 -704 220 -703
rect 229 -704 381 -703
rect 534 -704 783 -703
rect 30 -706 66 -705
rect 219 -706 409 -705
rect 544 -706 591 -705
rect 618 -706 689 -705
rect 30 -708 325 -707
rect 345 -708 409 -707
rect 555 -708 563 -707
rect 597 -708 689 -707
rect 233 -710 248 -709
rect 254 -710 339 -709
rect 380 -710 696 -709
rect 240 -712 276 -711
rect 324 -712 360 -711
rect 502 -712 563 -711
rect 597 -712 633 -711
rect 653 -712 682 -711
rect 695 -712 717 -711
rect 166 -714 360 -713
rect 478 -714 717 -713
rect 247 -716 332 -715
rect 338 -716 353 -715
rect 478 -716 549 -715
rect 576 -716 633 -715
rect 681 -716 724 -715
rect 275 -718 283 -717
rect 331 -718 388 -717
rect 530 -718 577 -717
rect 723 -718 745 -717
rect 282 -720 395 -719
rect 744 -720 759 -719
rect 320 -722 388 -721
rect 394 -722 507 -721
rect 730 -722 759 -721
rect 131 -724 731 -723
rect 352 -726 374 -725
rect 373 -728 402 -727
rect 401 -730 423 -729
rect 422 -732 542 -731
rect 2 -743 227 -742
rect 268 -743 276 -742
rect 289 -743 349 -742
rect 397 -743 465 -742
rect 481 -743 570 -742
rect 572 -743 738 -742
rect 782 -743 787 -742
rect 793 -743 808 -742
rect 9 -745 129 -744
rect 166 -745 220 -744
rect 268 -745 388 -744
rect 422 -745 703 -744
rect 737 -745 745 -744
rect 16 -747 59 -746
rect 65 -747 73 -746
rect 79 -747 318 -746
rect 345 -747 689 -746
rect 702 -747 724 -746
rect 744 -747 752 -746
rect 30 -749 230 -748
rect 275 -749 297 -748
rect 310 -749 346 -748
rect 366 -749 465 -748
rect 506 -749 570 -748
rect 576 -749 787 -748
rect 19 -751 367 -750
rect 376 -751 507 -750
rect 520 -751 556 -750
rect 600 -751 661 -750
rect 751 -751 759 -750
rect 30 -753 45 -752
rect 58 -753 122 -752
rect 184 -753 216 -752
rect 233 -753 297 -752
rect 310 -753 353 -752
rect 380 -753 689 -752
rect 758 -753 773 -752
rect 40 -755 164 -754
rect 184 -755 213 -754
rect 282 -755 388 -754
rect 408 -755 423 -754
rect 446 -755 724 -754
rect 772 -755 780 -754
rect 44 -757 412 -756
rect 450 -757 454 -756
rect 530 -757 640 -756
rect 72 -759 178 -758
rect 198 -759 202 -758
rect 205 -759 220 -758
rect 247 -759 283 -758
rect 289 -759 374 -758
rect 450 -759 493 -758
rect 541 -759 577 -758
rect 618 -759 661 -758
rect 75 -761 206 -760
rect 233 -761 248 -760
rect 320 -761 619 -760
rect 632 -761 640 -760
rect 79 -763 304 -762
rect 331 -763 353 -762
rect 359 -763 381 -762
rect 485 -763 493 -762
rect 534 -763 542 -762
rect 548 -763 605 -762
rect 86 -765 384 -764
rect 471 -765 535 -764
rect 551 -765 668 -764
rect 86 -767 101 -766
rect 107 -767 122 -766
rect 177 -767 262 -766
rect 303 -767 339 -766
rect 359 -767 458 -766
rect 471 -767 479 -766
rect 555 -767 591 -766
rect 597 -767 633 -766
rect 667 -767 696 -766
rect 89 -769 682 -768
rect 695 -769 710 -768
rect 93 -771 318 -770
rect 324 -771 339 -770
rect 362 -771 591 -770
rect 646 -771 682 -770
rect 23 -773 94 -772
rect 100 -773 150 -772
rect 170 -773 262 -772
rect 373 -773 717 -772
rect 23 -775 136 -774
rect 149 -775 192 -774
rect 198 -775 241 -774
rect 254 -775 325 -774
rect 404 -775 598 -774
rect 646 -775 675 -774
rect 716 -775 731 -774
rect 51 -777 171 -776
rect 191 -777 444 -776
rect 453 -777 486 -776
rect 548 -777 731 -776
rect 51 -779 426 -778
rect 443 -779 528 -778
rect 583 -779 605 -778
rect 107 -781 115 -780
rect 135 -781 143 -780
rect 159 -781 528 -780
rect 37 -783 115 -782
rect 142 -783 157 -782
rect 212 -783 332 -782
rect 457 -783 801 -782
rect 37 -785 612 -784
rect 254 -787 675 -786
rect 285 -789 612 -788
rect 478 -791 710 -790
rect 499 -793 584 -792
rect 436 -795 500 -794
rect 429 -797 437 -796
rect 415 -799 430 -798
rect 401 -801 416 -800
rect 68 -803 402 -802
rect 23 -814 157 -813
rect 170 -814 251 -813
rect 254 -814 276 -813
rect 282 -814 297 -813
rect 310 -814 381 -813
rect 394 -814 430 -813
rect 478 -814 528 -813
rect 544 -814 682 -813
rect 9 -816 24 -815
rect 30 -816 41 -815
rect 65 -816 132 -815
rect 156 -816 234 -815
rect 240 -816 258 -815
rect 271 -816 444 -815
rect 481 -816 563 -815
rect 597 -816 745 -815
rect 9 -818 129 -817
rect 177 -818 213 -817
rect 219 -818 223 -817
rect 226 -818 377 -817
rect 397 -818 486 -817
rect 513 -818 528 -817
rect 548 -818 647 -817
rect 744 -818 787 -817
rect 16 -820 66 -819
rect 72 -820 87 -819
rect 93 -820 227 -819
rect 240 -820 423 -819
rect 429 -820 458 -819
rect 485 -820 570 -819
rect 618 -820 766 -819
rect 86 -822 115 -821
rect 117 -822 160 -821
rect 184 -822 234 -821
rect 275 -822 332 -821
rect 345 -822 402 -821
rect 408 -822 503 -821
rect 513 -822 521 -821
rect 548 -822 605 -821
rect 618 -822 703 -821
rect 75 -824 115 -823
rect 121 -824 129 -823
rect 135 -824 178 -823
rect 184 -824 206 -823
rect 219 -824 304 -823
rect 331 -824 339 -823
rect 345 -824 591 -823
rect 646 -824 717 -823
rect 93 -826 108 -825
rect 110 -826 192 -825
rect 205 -826 269 -825
rect 282 -826 437 -825
rect 443 -826 507 -825
rect 562 -826 612 -825
rect 702 -826 752 -825
rect 72 -828 108 -827
rect 121 -828 150 -827
rect 191 -828 325 -827
rect 338 -828 388 -827
rect 404 -828 507 -827
rect 569 -828 633 -827
rect 751 -828 759 -827
rect 79 -830 269 -829
rect 296 -830 318 -829
rect 348 -830 689 -829
rect 758 -830 780 -829
rect 51 -832 80 -831
rect 100 -832 150 -831
rect 163 -832 318 -831
rect 359 -832 391 -831
rect 411 -832 584 -831
rect 590 -832 640 -831
rect 688 -832 727 -831
rect 30 -834 52 -833
rect 142 -834 164 -833
rect 222 -834 304 -833
rect 366 -834 521 -833
rect 583 -834 654 -833
rect 44 -836 101 -835
rect 247 -836 388 -835
rect 422 -836 493 -835
rect 611 -836 675 -835
rect 44 -838 139 -837
rect 198 -838 248 -837
rect 324 -838 367 -837
rect 373 -838 598 -837
rect 632 -838 661 -837
rect 58 -840 143 -839
rect 198 -840 290 -839
rect 373 -840 465 -839
rect 492 -840 608 -839
rect 639 -840 668 -839
rect 58 -842 174 -841
rect 264 -842 465 -841
rect 653 -842 696 -841
rect 289 -844 353 -843
rect 380 -844 661 -843
rect 667 -844 724 -843
rect 352 -846 416 -845
rect 436 -846 472 -845
rect 695 -846 731 -845
rect 415 -848 542 -847
rect 457 -850 535 -849
rect 471 -852 500 -851
rect 534 -852 556 -851
rect 555 -854 577 -853
rect 576 -856 626 -855
rect 625 -858 710 -857
rect 9 -869 398 -868
rect 471 -869 524 -868
rect 544 -869 584 -868
rect 604 -869 731 -868
rect 733 -869 738 -868
rect 747 -869 752 -868
rect 19 -871 24 -870
rect 51 -871 94 -870
rect 114 -871 118 -870
rect 124 -871 479 -870
rect 499 -871 535 -870
rect 583 -871 598 -870
rect 604 -871 640 -870
rect 663 -871 689 -870
rect 726 -871 759 -870
rect 54 -873 108 -872
rect 135 -873 178 -872
rect 180 -873 276 -872
rect 282 -873 384 -872
rect 387 -873 423 -872
rect 502 -873 633 -872
rect 674 -873 703 -872
rect 30 -875 283 -874
rect 317 -875 381 -874
rect 390 -875 451 -874
rect 520 -875 598 -874
rect 632 -875 647 -874
rect 681 -875 745 -874
rect 58 -877 178 -876
rect 212 -877 300 -876
rect 317 -877 339 -876
rect 345 -877 542 -876
rect 642 -877 647 -876
rect 681 -877 696 -876
rect 58 -879 87 -878
rect 93 -879 111 -878
rect 121 -879 136 -878
rect 142 -879 146 -878
rect 149 -879 171 -878
rect 257 -879 304 -878
rect 352 -879 370 -878
rect 401 -879 423 -878
rect 450 -879 528 -878
rect 534 -879 577 -878
rect 684 -879 717 -878
rect 65 -881 349 -880
rect 352 -881 395 -880
rect 401 -881 444 -880
rect 527 -881 570 -880
rect 576 -881 619 -880
rect 65 -883 220 -882
rect 261 -883 374 -882
rect 394 -883 654 -882
rect 79 -885 150 -884
rect 170 -885 311 -884
rect 366 -885 444 -884
rect 492 -885 570 -884
rect 618 -885 668 -884
rect 79 -887 241 -886
rect 271 -887 297 -886
rect 303 -887 332 -886
rect 373 -887 479 -886
rect 541 -887 563 -886
rect 86 -889 139 -888
rect 142 -889 192 -888
rect 198 -889 241 -888
rect 271 -889 377 -888
rect 464 -889 493 -888
rect 555 -889 668 -888
rect 100 -891 213 -890
rect 219 -891 255 -890
rect 275 -891 325 -890
rect 331 -891 437 -890
rect 562 -891 591 -890
rect 72 -893 101 -892
rect 107 -893 129 -892
rect 145 -893 192 -892
rect 198 -893 234 -892
rect 289 -893 339 -892
rect 415 -893 437 -892
rect 590 -893 612 -892
rect 72 -895 227 -894
rect 289 -895 409 -894
rect 415 -895 468 -894
rect 611 -895 626 -894
rect 40 -897 227 -896
rect 310 -897 360 -896
rect 408 -897 430 -896
rect 625 -897 661 -896
rect 128 -899 157 -898
rect 173 -899 556 -898
rect 156 -901 360 -900
rect 429 -901 458 -900
rect 506 -901 661 -900
rect 184 -903 234 -902
rect 457 -903 486 -902
rect 506 -903 549 -902
rect 184 -905 248 -904
rect 296 -905 549 -904
rect 44 -907 248 -906
rect 485 -907 514 -906
rect 44 -909 206 -908
rect 208 -909 514 -908
rect 205 -911 472 -910
rect 44 -922 454 -921
rect 464 -922 493 -921
rect 520 -922 577 -921
rect 646 -922 654 -921
rect 660 -922 675 -921
rect 716 -922 745 -921
rect 51 -924 122 -923
rect 170 -924 178 -923
rect 191 -924 206 -923
rect 219 -924 269 -923
rect 282 -924 314 -923
rect 320 -924 423 -923
rect 464 -924 556 -923
rect 674 -924 682 -923
rect 72 -926 94 -925
rect 103 -926 122 -925
rect 142 -926 220 -925
rect 226 -926 426 -925
rect 492 -926 570 -925
rect 107 -928 157 -927
rect 159 -928 171 -927
rect 184 -928 206 -927
rect 240 -928 325 -927
rect 394 -928 430 -927
rect 499 -928 577 -927
rect 86 -930 108 -929
rect 128 -930 143 -929
rect 184 -930 234 -929
rect 240 -930 353 -929
rect 499 -930 619 -929
rect 58 -932 87 -931
rect 100 -932 129 -931
rect 191 -932 367 -931
rect 527 -932 570 -931
rect 618 -932 640 -931
rect 114 -934 234 -933
rect 254 -934 430 -933
rect 450 -934 528 -933
rect 541 -934 643 -933
rect 198 -936 542 -935
rect 555 -936 612 -935
rect 149 -938 199 -937
rect 254 -938 437 -937
rect 534 -938 612 -937
rect 149 -940 227 -939
rect 268 -940 318 -939
rect 324 -940 472 -939
rect 156 -942 318 -941
rect 352 -942 416 -941
rect 436 -942 458 -941
rect 471 -942 486 -941
rect 275 -944 283 -943
rect 289 -944 300 -943
rect 310 -944 545 -943
rect 79 -946 290 -945
rect 296 -946 339 -945
rect 366 -946 633 -945
rect 79 -948 304 -947
rect 338 -948 360 -947
rect 408 -948 535 -947
rect 275 -950 346 -949
rect 359 -950 381 -949
rect 408 -950 444 -949
rect 457 -950 584 -949
rect 247 -952 346 -951
rect 380 -952 388 -951
rect 443 -952 514 -951
rect 583 -952 598 -951
rect 212 -954 248 -953
rect 303 -954 370 -953
rect 478 -954 486 -953
rect 513 -954 563 -953
rect 65 -956 213 -955
rect 331 -956 598 -955
rect 65 -958 258 -957
rect 261 -958 332 -957
rect 478 -958 549 -957
rect 261 -960 402 -959
rect 506 -960 563 -959
rect 373 -962 402 -961
rect 506 -962 629 -961
rect 548 -964 591 -963
rect 590 -966 626 -965
rect 604 -968 626 -967
rect 604 -970 668 -969
rect 65 -981 230 -980
rect 254 -981 419 -980
rect 422 -981 493 -980
rect 523 -981 528 -980
rect 544 -981 570 -980
rect 576 -981 580 -980
rect 607 -981 612 -980
rect 649 -981 661 -980
rect 670 -981 675 -980
rect 72 -983 97 -982
rect 100 -983 251 -982
rect 254 -983 363 -982
rect 373 -983 444 -982
rect 453 -983 500 -982
rect 527 -983 535 -982
rect 555 -983 570 -982
rect 576 -983 591 -982
rect 611 -983 619 -982
rect 79 -985 199 -984
rect 212 -985 370 -984
rect 380 -985 447 -984
rect 471 -985 500 -984
rect 579 -985 591 -984
rect 93 -987 101 -986
rect 107 -987 129 -986
rect 170 -987 202 -986
rect 264 -987 325 -986
rect 352 -987 391 -986
rect 394 -987 423 -986
rect 425 -987 437 -986
rect 439 -987 507 -986
rect 86 -989 171 -988
rect 191 -989 227 -988
rect 240 -989 353 -988
rect 369 -989 598 -988
rect 117 -991 122 -990
rect 177 -991 241 -990
rect 268 -991 374 -990
rect 380 -991 451 -990
rect 492 -991 514 -990
rect 163 -993 178 -992
rect 184 -993 269 -992
rect 296 -993 395 -992
rect 429 -993 647 -992
rect 156 -995 164 -994
rect 184 -995 206 -994
rect 226 -995 290 -994
rect 303 -995 437 -994
rect 450 -995 479 -994
rect 506 -995 584 -994
rect 142 -997 157 -996
rect 191 -997 283 -996
rect 310 -997 346 -996
rect 429 -997 486 -996
rect 562 -997 584 -996
rect 135 -999 143 -998
rect 205 -999 276 -998
rect 282 -999 367 -998
rect 233 -1001 276 -1000
rect 317 -1001 458 -1000
rect 219 -1003 234 -1002
rect 261 -1003 290 -1002
rect 324 -1003 339 -1002
rect 345 -1003 409 -1002
rect 457 -1003 605 -1002
rect 219 -1005 248 -1004
rect 338 -1005 360 -1004
rect 408 -1005 416 -1004
rect 247 -1007 304 -1006
rect 313 -1007 416 -1006
rect 359 -1009 388 -1008
rect 114 -1020 174 -1019
rect 198 -1020 349 -1019
rect 352 -1020 461 -1019
rect 478 -1020 507 -1019
rect 562 -1020 577 -1019
rect 604 -1020 612 -1019
rect 128 -1022 164 -1021
rect 198 -1022 220 -1021
rect 229 -1022 248 -1021
rect 268 -1022 367 -1021
rect 373 -1022 430 -1021
rect 436 -1022 451 -1021
rect 457 -1022 465 -1021
rect 485 -1022 493 -1021
rect 499 -1022 528 -1021
rect 135 -1024 150 -1023
rect 163 -1024 178 -1023
rect 191 -1024 248 -1023
rect 275 -1024 318 -1023
rect 366 -1024 381 -1023
rect 394 -1024 475 -1023
rect 149 -1026 157 -1025
rect 177 -1026 220 -1025
rect 226 -1026 269 -1025
rect 289 -1026 360 -1025
rect 373 -1026 416 -1025
rect 418 -1026 423 -1025
rect 142 -1028 157 -1027
rect 184 -1028 192 -1027
rect 205 -1028 307 -1027
rect 317 -1028 339 -1027
rect 394 -1028 402 -1027
rect 422 -1028 444 -1027
rect 124 -1030 143 -1029
rect 170 -1030 206 -1029
rect 215 -1030 234 -1029
rect 240 -1030 244 -1029
rect 254 -1030 290 -1029
rect 296 -1030 311 -1029
rect 439 -1030 444 -1029
rect 170 -1032 283 -1031
rect 299 -1032 304 -1031
rect 310 -1032 325 -1031
rect 215 -1034 255 -1033
rect 233 -1036 265 -1035
rect 261 -1038 265 -1037
rect 100 -1049 108 -1048
rect 128 -1049 195 -1048
rect 198 -1049 213 -1048
rect 219 -1049 227 -1048
rect 247 -1049 304 -1048
rect 366 -1049 381 -1048
rect 383 -1049 388 -1048
rect 394 -1049 405 -1048
rect 408 -1049 412 -1048
rect 415 -1049 430 -1048
rect 443 -1049 454 -1048
rect 471 -1049 486 -1048
rect 541 -1049 549 -1048
rect 579 -1049 584 -1048
rect 142 -1051 174 -1050
rect 180 -1051 234 -1050
rect 254 -1051 276 -1050
rect 278 -1051 297 -1050
rect 299 -1051 311 -1050
rect 376 -1051 423 -1050
rect 429 -1051 437 -1050
rect 443 -1051 479 -1050
rect 569 -1051 584 -1050
rect 142 -1053 157 -1052
rect 163 -1053 185 -1052
rect 191 -1053 199 -1052
rect 205 -1053 234 -1052
rect 268 -1053 283 -1052
rect 285 -1053 318 -1052
rect 579 -1053 591 -1052
rect 149 -1055 164 -1054
rect 289 -1055 297 -1054
rect 135 -1057 150 -1056
rect 114 -1059 136 -1058
rect 100 -1070 108 -1069
rect 149 -1070 160 -1069
rect 163 -1070 171 -1069
rect 198 -1070 206 -1069
rect 215 -1070 234 -1069
rect 380 -1070 395 -1069
rect 429 -1070 440 -1069
rect 446 -1070 458 -1069
rect 576 -1070 584 -1069
rect 219 -1072 227 -1071
<< m2contact >>
rect 114 0 115 1
rect 121 0 122 1
rect 128 0 129 1
rect 149 0 150 1
rect 156 0 157 1
rect 166 0 167 1
rect 177 0 178 1
rect 198 0 199 1
rect 236 0 237 1
rect 247 0 248 1
rect 296 0 297 1
rect 313 0 314 1
rect 317 0 318 1
rect 373 0 374 1
rect 131 -2 132 -1
rect 163 -2 164 -1
rect 191 -2 192 -1
rect 208 -2 209 -1
rect 331 -2 332 -1
rect 338 -2 339 -1
rect 348 -2 349 -1
rect 352 -2 353 -1
rect 135 -4 136 -3
rect 142 -4 143 -3
rect 72 -15 73 -14
rect 89 -15 90 -14
rect 100 -15 101 -14
rect 128 -15 129 -14
rect 131 -15 132 -14
rect 149 -15 150 -14
rect 156 -15 157 -14
rect 184 -15 185 -14
rect 187 -15 188 -14
rect 236 -15 237 -14
rect 247 -15 248 -14
rect 254 -15 255 -14
rect 296 -15 297 -14
rect 303 -15 304 -14
rect 331 -15 332 -14
rect 345 -15 346 -14
rect 373 -15 374 -14
rect 436 -15 437 -14
rect 485 -15 486 -14
rect 555 -15 556 -14
rect 79 -17 80 -16
rect 96 -17 97 -16
rect 107 -17 108 -16
rect 135 -17 136 -16
rect 142 -17 143 -16
rect 191 -17 192 -16
rect 201 -17 202 -16
rect 212 -17 213 -16
rect 215 -17 216 -16
rect 233 -17 234 -16
rect 296 -17 297 -16
rect 317 -17 318 -16
rect 394 -17 395 -16
rect 404 -17 405 -16
rect 422 -17 423 -16
rect 429 -17 430 -16
rect 117 -19 118 -18
rect 121 -19 122 -18
rect 135 -19 136 -18
rect 159 -19 160 -18
rect 170 -19 171 -18
rect 177 -19 178 -18
rect 184 -19 185 -18
rect 198 -19 199 -18
rect 219 -19 220 -18
rect 282 -19 283 -18
rect 313 -19 314 -18
rect 331 -19 332 -18
rect 156 -21 157 -20
rect 191 -21 192 -20
rect 229 -21 230 -20
rect 240 -21 241 -20
rect 173 -23 174 -22
rect 177 -23 178 -22
rect 51 -34 52 -33
rect 58 -34 59 -33
rect 65 -34 66 -33
rect 68 -34 69 -33
rect 79 -34 80 -33
rect 93 -34 94 -33
rect 96 -34 97 -33
rect 114 -34 115 -33
rect 149 -34 150 -33
rect 163 -34 164 -33
rect 166 -34 167 -33
rect 170 -34 171 -33
rect 191 -34 192 -33
rect 226 -34 227 -33
rect 233 -34 234 -33
rect 268 -34 269 -33
rect 275 -34 276 -33
rect 317 -34 318 -33
rect 345 -34 346 -33
rect 366 -34 367 -33
rect 387 -34 388 -33
rect 394 -34 395 -33
rect 415 -34 416 -33
rect 488 -34 489 -33
rect 555 -34 556 -33
rect 576 -34 577 -33
rect 65 -36 66 -35
rect 72 -36 73 -35
rect 86 -36 87 -35
rect 100 -36 101 -35
rect 107 -36 108 -35
rect 170 -36 171 -35
rect 212 -36 213 -35
rect 219 -36 220 -35
rect 233 -36 234 -35
rect 250 -36 251 -35
rect 254 -36 255 -35
rect 264 -36 265 -35
rect 285 -36 286 -35
rect 338 -36 339 -35
rect 352 -36 353 -35
rect 373 -36 374 -35
rect 380 -36 381 -35
rect 394 -36 395 -35
rect 429 -36 430 -35
rect 443 -36 444 -35
rect 68 -38 69 -37
rect 72 -38 73 -37
rect 100 -38 101 -37
rect 117 -38 118 -37
rect 149 -38 150 -37
rect 205 -38 206 -37
rect 240 -38 241 -37
rect 247 -38 248 -37
rect 289 -38 290 -37
rect 313 -38 314 -37
rect 327 -38 328 -37
rect 345 -38 346 -37
rect 359 -38 360 -37
rect 404 -38 405 -37
rect 436 -38 437 -37
rect 450 -38 451 -37
rect 107 -40 108 -39
rect 222 -40 223 -39
rect 303 -40 304 -39
rect 324 -40 325 -39
rect 331 -40 332 -39
rect 352 -40 353 -39
rect 156 -42 157 -41
rect 198 -42 199 -41
rect 254 -42 255 -41
rect 303 -42 304 -41
rect 159 -44 160 -43
rect 177 -44 178 -43
rect 194 -44 195 -43
rect 205 -44 206 -43
rect 282 -44 283 -43
rect 331 -44 332 -43
rect 121 -46 122 -45
rect 159 -46 160 -45
rect 177 -46 178 -45
rect 226 -46 227 -45
rect 121 -48 122 -47
rect 135 -48 136 -47
rect 135 -50 136 -49
rect 142 -50 143 -49
rect 142 -52 143 -51
rect 215 -52 216 -51
rect 30 -63 31 -62
rect 152 -63 153 -62
rect 156 -63 157 -62
rect 170 -63 171 -62
rect 191 -63 192 -62
rect 268 -63 269 -62
rect 366 -63 367 -62
rect 408 -63 409 -62
rect 425 -63 426 -62
rect 464 -63 465 -62
rect 471 -63 472 -62
rect 527 -63 528 -62
rect 530 -63 531 -62
rect 590 -63 591 -62
rect 37 -65 38 -64
rect 51 -65 52 -64
rect 58 -65 59 -64
rect 82 -65 83 -64
rect 93 -65 94 -64
rect 226 -65 227 -64
rect 233 -65 234 -64
rect 268 -65 269 -64
rect 373 -65 374 -64
rect 429 -65 430 -64
rect 443 -65 444 -64
rect 492 -65 493 -64
rect 44 -67 45 -66
rect 135 -67 136 -66
rect 142 -67 143 -66
rect 212 -67 213 -66
rect 240 -67 241 -66
rect 247 -67 248 -66
rect 261 -67 262 -66
rect 285 -67 286 -66
rect 303 -67 304 -66
rect 373 -67 374 -66
rect 380 -67 381 -66
rect 387 -67 388 -66
rect 401 -67 402 -66
rect 478 -67 479 -66
rect 51 -69 52 -68
rect 121 -69 122 -68
rect 131 -69 132 -68
rect 170 -69 171 -68
rect 205 -69 206 -68
rect 233 -69 234 -68
rect 240 -69 241 -68
rect 254 -69 255 -68
rect 261 -69 262 -68
rect 289 -69 290 -68
rect 387 -69 388 -68
rect 394 -69 395 -68
rect 401 -69 402 -68
rect 415 -69 416 -68
rect 65 -71 66 -70
rect 96 -71 97 -70
rect 100 -71 101 -70
rect 177 -71 178 -70
rect 289 -71 290 -70
rect 359 -71 360 -70
rect 72 -73 73 -72
rect 79 -73 80 -72
rect 86 -73 87 -72
rect 100 -73 101 -72
rect 128 -73 129 -72
rect 177 -73 178 -72
rect 324 -73 325 -72
rect 415 -73 416 -72
rect 65 -75 66 -74
rect 86 -75 87 -74
rect 128 -75 129 -74
rect 247 -75 248 -74
rect 313 -75 314 -74
rect 324 -75 325 -74
rect 331 -75 332 -74
rect 394 -75 395 -74
rect 72 -77 73 -76
rect 215 -77 216 -76
rect 296 -77 297 -76
rect 331 -77 332 -76
rect 345 -77 346 -76
rect 359 -77 360 -76
rect 131 -79 132 -78
rect 135 -79 136 -78
rect 142 -79 143 -78
rect 184 -79 185 -78
rect 219 -79 220 -78
rect 296 -79 297 -78
rect 313 -79 314 -78
rect 436 -79 437 -78
rect 149 -81 150 -80
rect 191 -81 192 -80
rect 219 -81 220 -80
rect 243 -81 244 -80
rect 345 -81 346 -80
rect 369 -81 370 -80
rect 163 -83 164 -82
rect 205 -83 206 -82
rect 163 -85 164 -84
rect 229 -85 230 -84
rect 184 -87 185 -86
rect 275 -87 276 -86
rect 275 -89 276 -88
rect 338 -89 339 -88
rect 338 -91 339 -90
rect 352 -91 353 -90
rect 9 -102 10 -101
rect 37 -102 38 -101
rect 51 -102 52 -101
rect 121 -102 122 -101
rect 128 -102 129 -101
rect 257 -102 258 -101
rect 282 -102 283 -101
rect 527 -102 528 -101
rect 555 -102 556 -101
rect 576 -102 577 -101
rect 590 -102 591 -101
rect 618 -102 619 -101
rect 16 -104 17 -103
rect 58 -104 59 -103
rect 65 -104 66 -103
rect 100 -104 101 -103
rect 121 -104 122 -103
rect 156 -104 157 -103
rect 170 -104 171 -103
rect 313 -104 314 -103
rect 331 -104 332 -103
rect 457 -104 458 -103
rect 460 -104 461 -103
rect 590 -104 591 -103
rect 26 -106 27 -105
rect 68 -106 69 -105
rect 75 -106 76 -105
rect 156 -106 157 -105
rect 173 -106 174 -105
rect 191 -106 192 -105
rect 240 -106 241 -105
rect 562 -106 563 -105
rect 30 -108 31 -107
rect 93 -108 94 -107
rect 100 -108 101 -107
rect 107 -108 108 -107
rect 149 -108 150 -107
rect 240 -108 241 -107
rect 243 -108 244 -107
rect 268 -108 269 -107
rect 282 -108 283 -107
rect 289 -108 290 -107
rect 313 -108 314 -107
rect 359 -108 360 -107
rect 366 -108 367 -107
rect 569 -108 570 -107
rect 37 -110 38 -109
rect 79 -110 80 -109
rect 86 -110 87 -109
rect 149 -110 150 -109
rect 191 -110 192 -109
rect 198 -110 199 -109
rect 226 -110 227 -109
rect 268 -110 269 -109
rect 275 -110 276 -109
rect 289 -110 290 -109
rect 338 -110 339 -109
rect 359 -110 360 -109
rect 366 -110 367 -109
rect 450 -110 451 -109
rect 478 -110 479 -109
rect 576 -110 577 -109
rect 30 -112 31 -111
rect 275 -112 276 -111
rect 345 -112 346 -111
rect 352 -112 353 -111
rect 355 -112 356 -111
rect 604 -112 605 -111
rect 51 -114 52 -113
rect 96 -114 97 -113
rect 107 -114 108 -113
rect 114 -114 115 -113
rect 142 -114 143 -113
rect 338 -114 339 -113
rect 345 -114 346 -113
rect 401 -114 402 -113
rect 415 -114 416 -113
rect 534 -114 535 -113
rect 58 -116 59 -115
rect 86 -116 87 -115
rect 114 -116 115 -115
rect 124 -116 125 -115
rect 142 -116 143 -115
rect 163 -116 164 -115
rect 198 -116 199 -115
rect 212 -116 213 -115
rect 226 -116 227 -115
rect 446 -116 447 -115
rect 492 -116 493 -115
rect 611 -116 612 -115
rect 205 -118 206 -117
rect 212 -118 213 -117
rect 233 -118 234 -117
rect 401 -118 402 -117
rect 415 -118 416 -117
rect 492 -118 493 -117
rect 499 -118 500 -117
rect 506 -118 507 -117
rect 520 -118 521 -117
rect 523 -118 524 -117
rect 135 -120 136 -119
rect 233 -120 234 -119
rect 247 -120 248 -119
rect 548 -120 549 -119
rect 44 -122 45 -121
rect 135 -122 136 -121
rect 205 -122 206 -121
rect 219 -122 220 -121
rect 247 -122 248 -121
rect 303 -122 304 -121
rect 373 -122 374 -121
rect 513 -122 514 -121
rect 44 -124 45 -123
rect 72 -124 73 -123
rect 184 -124 185 -123
rect 303 -124 304 -123
rect 320 -124 321 -123
rect 373 -124 374 -123
rect 387 -124 388 -123
rect 450 -124 451 -123
rect 72 -126 73 -125
rect 331 -126 332 -125
rect 394 -126 395 -125
rect 597 -126 598 -125
rect 159 -128 160 -127
rect 184 -128 185 -127
rect 219 -128 220 -127
rect 222 -128 223 -127
rect 261 -128 262 -127
rect 320 -128 321 -127
rect 324 -128 325 -127
rect 387 -128 388 -127
rect 422 -128 423 -127
rect 464 -128 465 -127
rect 170 -130 171 -129
rect 261 -130 262 -129
rect 296 -130 297 -129
rect 394 -130 395 -129
rect 408 -130 409 -129
rect 464 -130 465 -129
rect 177 -132 178 -131
rect 296 -132 297 -131
rect 310 -132 311 -131
rect 324 -132 325 -131
rect 408 -132 409 -131
rect 471 -132 472 -131
rect 166 -134 167 -133
rect 177 -134 178 -133
rect 429 -134 430 -133
rect 478 -134 479 -133
rect 429 -136 430 -135
rect 474 -136 475 -135
rect 436 -138 437 -137
rect 485 -138 486 -137
rect 380 -140 381 -139
rect 436 -140 437 -139
rect 443 -140 444 -139
rect 541 -140 542 -139
rect 257 -142 258 -141
rect 380 -142 381 -141
rect 443 -142 444 -141
rect 586 -142 587 -141
rect 23 -153 24 -152
rect 191 -153 192 -152
rect 205 -153 206 -152
rect 257 -153 258 -152
rect 261 -153 262 -152
rect 569 -153 570 -152
rect 611 -153 612 -152
rect 660 -153 661 -152
rect 51 -155 52 -154
rect 180 -155 181 -154
rect 184 -155 185 -154
rect 418 -155 419 -154
rect 464 -155 465 -154
rect 639 -155 640 -154
rect 51 -157 52 -156
rect 128 -157 129 -156
rect 142 -157 143 -156
rect 184 -157 185 -156
rect 191 -157 192 -156
rect 292 -157 293 -156
rect 306 -157 307 -156
rect 597 -157 598 -156
rect 618 -157 619 -156
rect 625 -157 626 -156
rect 628 -157 629 -156
rect 646 -157 647 -156
rect 65 -159 66 -158
rect 93 -159 94 -158
rect 100 -159 101 -158
rect 128 -159 129 -158
rect 135 -159 136 -158
rect 142 -159 143 -158
rect 156 -159 157 -158
rect 163 -159 164 -158
rect 173 -159 174 -158
rect 198 -159 199 -158
rect 212 -159 213 -158
rect 310 -159 311 -158
rect 313 -159 314 -158
rect 590 -159 591 -158
rect 604 -159 605 -158
rect 625 -159 626 -158
rect 58 -161 59 -160
rect 65 -161 66 -160
rect 72 -161 73 -160
rect 138 -161 139 -160
rect 198 -161 199 -160
rect 247 -161 248 -160
rect 254 -161 255 -160
rect 296 -161 297 -160
rect 334 -161 335 -160
rect 667 -161 668 -160
rect 16 -163 17 -162
rect 58 -163 59 -162
rect 79 -163 80 -162
rect 156 -163 157 -162
rect 212 -163 213 -162
rect 261 -163 262 -162
rect 278 -163 279 -162
rect 534 -163 535 -162
rect 541 -163 542 -162
rect 569 -163 570 -162
rect 576 -163 577 -162
rect 590 -163 591 -162
rect 16 -165 17 -164
rect 44 -165 45 -164
rect 79 -165 80 -164
rect 107 -165 108 -164
rect 135 -165 136 -164
rect 299 -165 300 -164
rect 387 -165 388 -164
rect 674 -165 675 -164
rect 44 -167 45 -166
rect 282 -167 283 -166
rect 289 -167 290 -166
rect 324 -167 325 -166
rect 387 -167 388 -166
rect 618 -167 619 -166
rect 82 -169 83 -168
rect 96 -169 97 -168
rect 100 -169 101 -168
rect 401 -169 402 -168
rect 436 -169 437 -168
rect 464 -169 465 -168
rect 471 -169 472 -168
rect 597 -169 598 -168
rect 86 -171 87 -170
rect 149 -171 150 -170
rect 215 -171 216 -170
rect 394 -171 395 -170
rect 457 -171 458 -170
rect 534 -171 535 -170
rect 562 -171 563 -170
rect 604 -171 605 -170
rect 86 -173 87 -172
rect 114 -173 115 -172
rect 149 -173 150 -172
rect 527 -173 528 -172
rect 555 -173 556 -172
rect 562 -173 563 -172
rect 107 -175 108 -174
rect 121 -175 122 -174
rect 219 -175 220 -174
rect 338 -175 339 -174
rect 341 -175 342 -174
rect 471 -175 472 -174
rect 485 -175 486 -174
rect 632 -175 633 -174
rect 30 -177 31 -176
rect 219 -177 220 -176
rect 247 -177 248 -176
rect 586 -177 587 -176
rect 30 -179 31 -178
rect 240 -179 241 -178
rect 268 -179 269 -178
rect 394 -179 395 -178
rect 422 -179 423 -178
rect 457 -179 458 -178
rect 492 -179 493 -178
rect 611 -179 612 -178
rect 37 -181 38 -180
rect 121 -181 122 -180
rect 222 -181 223 -180
rect 422 -181 423 -180
rect 499 -181 500 -180
rect 513 -181 514 -180
rect 520 -181 521 -180
rect 541 -181 542 -180
rect 37 -183 38 -182
rect 96 -183 97 -182
rect 114 -183 115 -182
rect 226 -183 227 -182
rect 240 -183 241 -182
rect 278 -183 279 -182
rect 282 -183 283 -182
rect 369 -183 370 -182
rect 390 -183 391 -182
rect 653 -183 654 -182
rect 177 -185 178 -184
rect 226 -185 227 -184
rect 296 -185 297 -184
rect 380 -185 381 -184
rect 488 -185 489 -184
rect 513 -185 514 -184
rect 520 -185 521 -184
rect 583 -185 584 -184
rect 177 -187 178 -186
rect 208 -187 209 -186
rect 317 -187 318 -186
rect 555 -187 556 -186
rect 268 -189 269 -188
rect 317 -189 318 -188
rect 320 -189 321 -188
rect 436 -189 437 -188
rect 506 -189 507 -188
rect 527 -189 528 -188
rect 548 -189 549 -188
rect 583 -189 584 -188
rect 359 -191 360 -190
rect 492 -191 493 -190
rect 331 -193 332 -192
rect 359 -193 360 -192
rect 366 -193 367 -192
rect 401 -193 402 -192
rect 415 -193 416 -192
rect 548 -193 549 -192
rect 331 -195 332 -194
rect 576 -195 577 -194
rect 345 -197 346 -196
rect 415 -197 416 -196
rect 478 -197 479 -196
rect 506 -197 507 -196
rect 170 -199 171 -198
rect 345 -199 346 -198
rect 373 -199 374 -198
rect 380 -199 381 -198
rect 408 -199 409 -198
rect 478 -199 479 -198
rect 9 -201 10 -200
rect 170 -201 171 -200
rect 352 -201 353 -200
rect 373 -201 374 -200
rect 408 -201 409 -200
rect 429 -201 430 -200
rect 303 -203 304 -202
rect 352 -203 353 -202
rect 429 -203 430 -202
rect 443 -203 444 -202
rect 23 -214 24 -213
rect 212 -214 213 -213
rect 275 -214 276 -213
rect 534 -214 535 -213
rect 548 -214 549 -213
rect 688 -214 689 -213
rect 23 -216 24 -215
rect 96 -216 97 -215
rect 100 -216 101 -215
rect 107 -216 108 -215
rect 152 -216 153 -215
rect 243 -216 244 -215
rect 292 -216 293 -215
rect 534 -216 535 -215
rect 548 -216 549 -215
rect 597 -216 598 -215
rect 653 -216 654 -215
rect 695 -216 696 -215
rect 44 -218 45 -217
rect 93 -218 94 -217
rect 103 -218 104 -217
rect 233 -218 234 -217
rect 296 -218 297 -217
rect 429 -218 430 -217
rect 446 -218 447 -217
rect 597 -218 598 -217
rect 660 -218 661 -217
rect 716 -218 717 -217
rect 44 -220 45 -219
rect 54 -220 55 -219
rect 65 -220 66 -219
rect 75 -220 76 -219
rect 86 -220 87 -219
rect 135 -220 136 -219
rect 156 -220 157 -219
rect 278 -220 279 -219
rect 303 -220 304 -219
rect 352 -220 353 -219
rect 369 -220 370 -219
rect 618 -220 619 -219
rect 51 -222 52 -221
rect 72 -222 73 -221
rect 86 -222 87 -221
rect 278 -222 279 -221
rect 313 -222 314 -221
rect 569 -222 570 -221
rect 583 -222 584 -221
rect 618 -222 619 -221
rect 51 -224 52 -223
rect 149 -224 150 -223
rect 170 -224 171 -223
rect 324 -224 325 -223
rect 331 -224 332 -223
rect 639 -224 640 -223
rect 37 -226 38 -225
rect 331 -226 332 -225
rect 338 -226 339 -225
rect 359 -226 360 -225
rect 369 -226 370 -225
rect 569 -226 570 -225
rect 590 -226 591 -225
rect 653 -226 654 -225
rect 9 -228 10 -227
rect 37 -228 38 -227
rect 65 -228 66 -227
rect 82 -228 83 -227
rect 128 -228 129 -227
rect 156 -228 157 -227
rect 177 -228 178 -227
rect 310 -228 311 -227
rect 341 -228 342 -227
rect 492 -228 493 -227
rect 499 -228 500 -227
rect 590 -228 591 -227
rect 611 -228 612 -227
rect 660 -228 661 -227
rect 16 -230 17 -229
rect 177 -230 178 -229
rect 191 -230 192 -229
rect 205 -230 206 -229
rect 233 -230 234 -229
rect 240 -230 241 -229
rect 254 -230 255 -229
rect 352 -230 353 -229
rect 387 -230 388 -229
rect 632 -230 633 -229
rect 16 -232 17 -231
rect 117 -232 118 -231
rect 128 -232 129 -231
rect 184 -232 185 -231
rect 191 -232 192 -231
rect 226 -232 227 -231
rect 254 -232 255 -231
rect 268 -232 269 -231
rect 299 -232 300 -231
rect 639 -232 640 -231
rect 30 -234 31 -233
rect 310 -234 311 -233
rect 345 -234 346 -233
rect 359 -234 360 -233
rect 422 -234 423 -233
rect 723 -234 724 -233
rect 33 -236 34 -235
rect 226 -236 227 -235
rect 247 -236 248 -235
rect 345 -236 346 -235
rect 408 -236 409 -235
rect 422 -236 423 -235
rect 457 -236 458 -235
rect 485 -236 486 -235
rect 488 -236 489 -235
rect 604 -236 605 -235
rect 79 -238 80 -237
rect 170 -238 171 -237
rect 198 -238 199 -237
rect 201 -238 202 -237
rect 247 -238 248 -237
rect 681 -238 682 -237
rect 2 -240 3 -239
rect 79 -240 80 -239
rect 107 -240 108 -239
rect 387 -240 388 -239
rect 464 -240 465 -239
rect 492 -240 493 -239
rect 513 -240 514 -239
rect 702 -240 703 -239
rect 121 -242 122 -241
rect 184 -242 185 -241
rect 198 -242 199 -241
rect 289 -242 290 -241
rect 299 -242 300 -241
rect 429 -242 430 -241
rect 471 -242 472 -241
rect 499 -242 500 -241
rect 513 -242 514 -241
rect 674 -242 675 -241
rect 121 -244 122 -243
rect 264 -244 265 -243
rect 268 -244 269 -243
rect 282 -244 283 -243
rect 327 -244 328 -243
rect 457 -244 458 -243
rect 471 -244 472 -243
rect 478 -244 479 -243
rect 527 -244 528 -243
rect 583 -244 584 -243
rect 135 -246 136 -245
rect 180 -246 181 -245
rect 201 -246 202 -245
rect 289 -246 290 -245
rect 366 -246 367 -245
rect 527 -246 528 -245
rect 555 -246 556 -245
rect 604 -246 605 -245
rect 250 -248 251 -247
rect 555 -248 556 -247
rect 562 -248 563 -247
rect 632 -248 633 -247
rect 261 -250 262 -249
rect 282 -250 283 -249
rect 380 -250 381 -249
rect 408 -250 409 -249
rect 436 -250 437 -249
rect 478 -250 479 -249
rect 506 -250 507 -249
rect 562 -250 563 -249
rect 576 -250 577 -249
rect 611 -250 612 -249
rect 380 -252 381 -251
rect 646 -252 647 -251
rect 383 -254 384 -253
rect 674 -254 675 -253
rect 394 -256 395 -255
rect 436 -256 437 -255
rect 506 -256 507 -255
rect 667 -256 668 -255
rect 394 -258 395 -257
rect 401 -258 402 -257
rect 541 -258 542 -257
rect 576 -258 577 -257
rect 625 -258 626 -257
rect 667 -258 668 -257
rect 373 -260 374 -259
rect 401 -260 402 -259
rect 415 -260 416 -259
rect 541 -260 542 -259
rect 646 -260 647 -259
rect 712 -260 713 -259
rect 30 -262 31 -261
rect 373 -262 374 -261
rect 443 -262 444 -261
rect 625 -262 626 -261
rect 317 -264 318 -263
rect 415 -264 416 -263
rect 443 -264 444 -263
rect 450 -264 451 -263
rect 114 -266 115 -265
rect 317 -266 318 -265
rect 450 -266 451 -265
rect 520 -266 521 -265
rect 520 -268 521 -267
rect 730 -268 731 -267
rect 23 -279 24 -278
rect 54 -279 55 -278
rect 58 -279 59 -278
rect 110 -279 111 -278
rect 128 -279 129 -278
rect 278 -279 279 -278
rect 289 -279 290 -278
rect 352 -279 353 -278
rect 362 -279 363 -278
rect 541 -279 542 -278
rect 569 -279 570 -278
rect 730 -279 731 -278
rect 26 -281 27 -280
rect 226 -281 227 -280
rect 240 -281 241 -280
rect 527 -281 528 -280
rect 534 -281 535 -280
rect 569 -281 570 -280
rect 716 -281 717 -280
rect 737 -281 738 -280
rect 2 -283 3 -282
rect 226 -283 227 -282
rect 247 -283 248 -282
rect 303 -283 304 -282
rect 310 -283 311 -282
rect 338 -283 339 -282
rect 345 -283 346 -282
rect 352 -283 353 -282
rect 380 -283 381 -282
rect 639 -283 640 -282
rect 30 -285 31 -284
rect 72 -285 73 -284
rect 82 -285 83 -284
rect 667 -285 668 -284
rect 16 -287 17 -286
rect 72 -287 73 -286
rect 86 -287 87 -286
rect 303 -287 304 -286
rect 310 -287 311 -286
rect 313 -287 314 -286
rect 338 -287 339 -286
rect 415 -287 416 -286
rect 422 -287 423 -286
rect 464 -287 465 -286
rect 467 -287 468 -286
rect 548 -287 549 -286
rect 639 -287 640 -286
rect 653 -287 654 -286
rect 667 -287 668 -286
rect 681 -287 682 -286
rect 16 -289 17 -288
rect 205 -289 206 -288
rect 212 -289 213 -288
rect 250 -289 251 -288
rect 292 -289 293 -288
rect 716 -289 717 -288
rect 33 -291 34 -290
rect 534 -291 535 -290
rect 541 -291 542 -290
rect 590 -291 591 -290
rect 653 -291 654 -290
rect 674 -291 675 -290
rect 37 -293 38 -292
rect 79 -293 80 -292
rect 100 -293 101 -292
rect 170 -293 171 -292
rect 198 -293 199 -292
rect 348 -293 349 -292
rect 380 -293 381 -292
rect 401 -293 402 -292
rect 422 -293 423 -292
rect 506 -293 507 -292
rect 548 -293 549 -292
rect 562 -293 563 -292
rect 590 -293 591 -292
rect 611 -293 612 -292
rect 44 -295 45 -294
rect 527 -295 528 -294
rect 555 -295 556 -294
rect 681 -295 682 -294
rect 47 -297 48 -296
rect 436 -297 437 -296
rect 499 -297 500 -296
rect 506 -297 507 -296
rect 555 -297 556 -296
rect 597 -297 598 -296
rect 51 -299 52 -298
rect 86 -299 87 -298
rect 107 -299 108 -298
rect 205 -299 206 -298
rect 212 -299 213 -298
rect 383 -299 384 -298
rect 394 -299 395 -298
rect 415 -299 416 -298
rect 432 -299 433 -298
rect 520 -299 521 -298
rect 562 -299 563 -298
rect 583 -299 584 -298
rect 597 -299 598 -298
rect 625 -299 626 -298
rect 54 -301 55 -300
rect 114 -301 115 -300
rect 121 -301 122 -300
rect 128 -301 129 -300
rect 135 -301 136 -300
rect 149 -301 150 -300
rect 156 -301 157 -300
rect 240 -301 241 -300
rect 257 -301 258 -300
rect 611 -301 612 -300
rect 625 -301 626 -300
rect 632 -301 633 -300
rect 58 -303 59 -302
rect 296 -303 297 -302
rect 345 -303 346 -302
rect 702 -303 703 -302
rect 65 -305 66 -304
rect 187 -305 188 -304
rect 191 -305 192 -304
rect 198 -305 199 -304
rect 219 -305 220 -304
rect 247 -305 248 -304
rect 261 -305 262 -304
rect 674 -305 675 -304
rect 65 -307 66 -306
rect 268 -307 269 -306
rect 299 -307 300 -306
rect 702 -307 703 -306
rect 93 -309 94 -308
rect 268 -309 269 -308
rect 299 -309 300 -308
rect 513 -309 514 -308
rect 583 -309 584 -308
rect 618 -309 619 -308
rect 632 -309 633 -308
rect 646 -309 647 -308
rect 110 -311 111 -310
rect 114 -311 115 -310
rect 121 -311 122 -310
rect 369 -311 370 -310
rect 394 -311 395 -310
rect 408 -311 409 -310
rect 436 -311 437 -310
rect 709 -311 710 -310
rect 135 -313 136 -312
rect 184 -313 185 -312
rect 191 -313 192 -312
rect 282 -313 283 -312
rect 401 -313 402 -312
rect 723 -313 724 -312
rect 37 -315 38 -314
rect 184 -315 185 -314
rect 275 -315 276 -314
rect 618 -315 619 -314
rect 646 -315 647 -314
rect 660 -315 661 -314
rect 695 -315 696 -314
rect 723 -315 724 -314
rect 44 -317 45 -316
rect 695 -317 696 -316
rect 93 -319 94 -318
rect 282 -319 283 -318
rect 443 -319 444 -318
rect 499 -319 500 -318
rect 660 -319 661 -318
rect 688 -319 689 -318
rect 142 -321 143 -320
rect 170 -321 171 -320
rect 177 -321 178 -320
rect 261 -321 262 -320
rect 275 -321 276 -320
rect 408 -321 409 -320
rect 457 -321 458 -320
rect 520 -321 521 -320
rect 142 -323 143 -322
rect 264 -323 265 -322
rect 324 -323 325 -322
rect 457 -323 458 -322
rect 471 -323 472 -322
rect 513 -323 514 -322
rect 156 -325 157 -324
rect 233 -325 234 -324
rect 324 -325 325 -324
rect 387 -325 388 -324
rect 450 -325 451 -324
rect 471 -325 472 -324
rect 51 -327 52 -326
rect 233 -327 234 -326
rect 278 -327 279 -326
rect 387 -327 388 -326
rect 429 -327 430 -326
rect 450 -327 451 -326
rect 163 -329 164 -328
rect 219 -329 220 -328
rect 327 -329 328 -328
rect 688 -329 689 -328
rect 177 -331 178 -330
rect 254 -331 255 -330
rect 331 -331 332 -330
rect 443 -331 444 -330
rect 317 -333 318 -332
rect 331 -333 332 -332
rect 429 -333 430 -332
rect 709 -333 710 -332
rect 317 -335 318 -334
rect 359 -335 360 -334
rect 5 -346 6 -345
rect 359 -346 360 -345
rect 369 -346 370 -345
rect 478 -346 479 -345
rect 555 -346 556 -345
rect 758 -346 759 -345
rect 23 -348 24 -347
rect 366 -348 367 -347
rect 376 -348 377 -347
rect 800 -348 801 -347
rect 26 -350 27 -349
rect 450 -350 451 -349
rect 474 -350 475 -349
rect 765 -350 766 -349
rect 30 -352 31 -351
rect 184 -352 185 -351
rect 187 -352 188 -351
rect 247 -352 248 -351
rect 268 -352 269 -351
rect 278 -352 279 -351
rect 282 -352 283 -351
rect 569 -352 570 -351
rect 667 -352 668 -351
rect 744 -352 745 -351
rect 30 -354 31 -353
rect 156 -354 157 -353
rect 219 -354 220 -353
rect 254 -354 255 -353
rect 268 -354 269 -353
rect 457 -354 458 -353
rect 513 -354 514 -353
rect 569 -354 570 -353
rect 583 -354 584 -353
rect 667 -354 668 -353
rect 674 -354 675 -353
rect 751 -354 752 -353
rect 2 -356 3 -355
rect 583 -356 584 -355
rect 688 -356 689 -355
rect 772 -356 773 -355
rect 44 -358 45 -357
rect 397 -358 398 -357
rect 408 -358 409 -357
rect 457 -358 458 -357
rect 464 -358 465 -357
rect 513 -358 514 -357
rect 527 -358 528 -357
rect 674 -358 675 -357
rect 695 -358 696 -357
rect 779 -358 780 -357
rect 47 -360 48 -359
rect 296 -360 297 -359
rect 324 -360 325 -359
rect 345 -360 346 -359
rect 352 -360 353 -359
rect 366 -360 367 -359
rect 408 -360 409 -359
rect 415 -360 416 -359
rect 432 -360 433 -359
rect 723 -360 724 -359
rect 730 -360 731 -359
rect 807 -360 808 -359
rect 51 -362 52 -361
rect 191 -362 192 -361
rect 219 -362 220 -361
rect 443 -362 444 -361
rect 485 -362 486 -361
rect 527 -362 528 -361
rect 558 -362 559 -361
rect 814 -362 815 -361
rect 54 -364 55 -363
rect 404 -364 405 -363
rect 415 -364 416 -363
rect 737 -364 738 -363
rect 61 -366 62 -365
rect 229 -366 230 -365
rect 233 -366 234 -365
rect 418 -366 419 -365
rect 422 -366 423 -365
rect 443 -366 444 -365
rect 471 -366 472 -365
rect 485 -366 486 -365
rect 618 -366 619 -365
rect 688 -366 689 -365
rect 709 -366 710 -365
rect 786 -366 787 -365
rect 72 -368 73 -367
rect 233 -368 234 -367
rect 247 -368 248 -367
rect 338 -368 339 -367
rect 345 -368 346 -367
rect 702 -368 703 -367
rect 716 -368 717 -367
rect 793 -368 794 -367
rect 72 -370 73 -369
rect 86 -370 87 -369
rect 93 -370 94 -369
rect 275 -370 276 -369
rect 282 -370 283 -369
rect 331 -370 332 -369
rect 338 -370 339 -369
rect 450 -370 451 -369
rect 625 -370 626 -369
rect 695 -370 696 -369
rect 37 -372 38 -371
rect 331 -372 332 -371
rect 348 -372 349 -371
rect 723 -372 724 -371
rect 79 -374 80 -373
rect 191 -374 192 -373
rect 226 -374 227 -373
rect 352 -374 353 -373
rect 387 -374 388 -373
rect 422 -374 423 -373
rect 429 -374 430 -373
rect 618 -374 619 -373
rect 639 -374 640 -373
rect 702 -374 703 -373
rect 79 -376 80 -375
rect 177 -376 178 -375
rect 226 -376 227 -375
rect 317 -376 318 -375
rect 348 -376 349 -375
rect 737 -376 738 -375
rect 86 -378 87 -377
rect 135 -378 136 -377
rect 285 -378 286 -377
rect 523 -378 524 -377
rect 541 -378 542 -377
rect 639 -378 640 -377
rect 646 -378 647 -377
rect 709 -378 710 -377
rect 93 -380 94 -379
rect 341 -380 342 -379
rect 436 -380 437 -379
rect 478 -380 479 -379
rect 492 -380 493 -379
rect 541 -380 542 -379
rect 576 -380 577 -379
rect 625 -380 626 -379
rect 646 -380 647 -379
rect 660 -380 661 -379
rect 681 -380 682 -379
rect 730 -380 731 -379
rect 100 -382 101 -381
rect 135 -382 136 -381
rect 289 -382 290 -381
rect 387 -382 388 -381
rect 394 -382 395 -381
rect 436 -382 437 -381
rect 492 -382 493 -381
rect 499 -382 500 -381
rect 520 -382 521 -381
rect 576 -382 577 -381
rect 590 -382 591 -381
rect 660 -382 661 -381
rect 100 -384 101 -383
rect 205 -384 206 -383
rect 292 -384 293 -383
rect 464 -384 465 -383
rect 590 -384 591 -383
rect 597 -384 598 -383
rect 611 -384 612 -383
rect 681 -384 682 -383
rect 107 -386 108 -385
rect 632 -386 633 -385
rect 653 -386 654 -385
rect 716 -386 717 -385
rect 110 -388 111 -387
rect 254 -388 255 -387
rect 296 -388 297 -387
rect 303 -388 304 -387
rect 310 -388 311 -387
rect 317 -388 318 -387
rect 534 -388 535 -387
rect 597 -388 598 -387
rect 604 -388 605 -387
rect 611 -388 612 -387
rect 110 -390 111 -389
rect 499 -390 500 -389
rect 548 -390 549 -389
rect 653 -390 654 -389
rect 121 -392 122 -391
rect 205 -392 206 -391
rect 222 -392 223 -391
rect 310 -392 311 -391
rect 383 -392 384 -391
rect 604 -392 605 -391
rect 124 -394 125 -393
rect 156 -394 157 -393
rect 163 -394 164 -393
rect 289 -394 290 -393
rect 299 -394 300 -393
rect 632 -394 633 -393
rect 114 -396 115 -395
rect 163 -396 164 -395
rect 303 -396 304 -395
rect 334 -396 335 -395
rect 401 -396 402 -395
rect 534 -396 535 -395
rect 37 -398 38 -397
rect 401 -398 402 -397
rect 506 -398 507 -397
rect 548 -398 549 -397
rect 114 -400 115 -399
rect 240 -400 241 -399
rect 128 -402 129 -401
rect 177 -402 178 -401
rect 240 -402 241 -401
rect 380 -402 381 -401
rect 128 -404 129 -403
rect 142 -404 143 -403
rect 212 -404 213 -403
rect 380 -404 381 -403
rect 16 -406 17 -405
rect 212 -406 213 -405
rect 16 -408 17 -407
rect 198 -408 199 -407
rect 142 -410 143 -409
rect 170 -410 171 -409
rect 198 -410 199 -409
rect 394 -410 395 -409
rect 65 -412 66 -411
rect 170 -412 171 -411
rect 58 -414 59 -413
rect 65 -414 66 -413
rect 9 -425 10 -424
rect 51 -425 52 -424
rect 58 -425 59 -424
rect 68 -425 69 -424
rect 72 -425 73 -424
rect 138 -425 139 -424
rect 170 -425 171 -424
rect 219 -425 220 -424
rect 264 -425 265 -424
rect 751 -425 752 -424
rect 9 -427 10 -426
rect 44 -427 45 -426
rect 47 -427 48 -426
rect 667 -427 668 -426
rect 702 -427 703 -426
rect 705 -427 706 -426
rect 51 -429 52 -428
rect 100 -429 101 -428
rect 107 -429 108 -428
rect 674 -429 675 -428
rect 702 -429 703 -428
rect 744 -429 745 -428
rect 58 -431 59 -430
rect 758 -431 759 -430
rect 61 -433 62 -432
rect 268 -433 269 -432
rect 275 -433 276 -432
rect 373 -433 374 -432
rect 380 -433 381 -432
rect 660 -433 661 -432
rect 730 -433 731 -432
rect 744 -433 745 -432
rect 72 -435 73 -434
rect 198 -435 199 -434
rect 205 -435 206 -434
rect 289 -435 290 -434
rect 334 -435 335 -434
rect 597 -435 598 -434
rect 611 -435 612 -434
rect 674 -435 675 -434
rect 716 -435 717 -434
rect 730 -435 731 -434
rect 79 -437 80 -436
rect 275 -437 276 -436
rect 338 -437 339 -436
rect 653 -437 654 -436
rect 79 -439 80 -438
rect 296 -439 297 -438
rect 348 -439 349 -438
rect 723 -439 724 -438
rect 86 -441 87 -440
rect 121 -441 122 -440
rect 163 -441 164 -440
rect 205 -441 206 -440
rect 233 -441 234 -440
rect 338 -441 339 -440
rect 366 -441 367 -440
rect 383 -441 384 -440
rect 394 -441 395 -440
rect 639 -441 640 -440
rect 646 -441 647 -440
rect 758 -441 759 -440
rect 44 -443 45 -442
rect 233 -443 234 -442
rect 254 -443 255 -442
rect 296 -443 297 -442
rect 387 -443 388 -442
rect 394 -443 395 -442
rect 401 -443 402 -442
rect 632 -443 633 -442
rect 709 -443 710 -442
rect 723 -443 724 -442
rect 86 -445 87 -444
rect 359 -445 360 -444
rect 404 -445 405 -444
rect 793 -445 794 -444
rect 93 -447 94 -446
rect 163 -447 164 -446
rect 170 -447 171 -446
rect 222 -447 223 -446
rect 226 -447 227 -446
rect 366 -447 367 -446
rect 443 -447 444 -446
rect 611 -447 612 -446
rect 618 -447 619 -446
rect 639 -447 640 -446
rect 695 -447 696 -446
rect 709 -447 710 -446
rect 793 -447 794 -446
rect 807 -447 808 -446
rect 93 -449 94 -448
rect 345 -449 346 -448
rect 352 -449 353 -448
rect 359 -449 360 -448
rect 474 -449 475 -448
rect 772 -449 773 -448
rect 100 -451 101 -450
rect 404 -451 405 -450
rect 474 -451 475 -450
rect 660 -451 661 -450
rect 681 -451 682 -450
rect 695 -451 696 -450
rect 772 -451 773 -450
rect 786 -451 787 -450
rect 107 -453 108 -452
rect 128 -453 129 -452
rect 198 -453 199 -452
rect 317 -453 318 -452
rect 324 -453 325 -452
rect 345 -453 346 -452
rect 355 -453 356 -452
rect 618 -453 619 -452
rect 625 -453 626 -452
rect 646 -453 647 -452
rect 786 -453 787 -452
rect 800 -453 801 -452
rect 30 -455 31 -454
rect 128 -455 129 -454
rect 191 -455 192 -454
rect 324 -455 325 -454
rect 506 -455 507 -454
rect 597 -455 598 -454
rect 604 -455 605 -454
rect 632 -455 633 -454
rect 800 -455 801 -454
rect 814 -455 815 -454
rect 30 -457 31 -456
rect 432 -457 433 -456
rect 520 -457 521 -456
rect 737 -457 738 -456
rect 37 -459 38 -458
rect 506 -459 507 -458
rect 523 -459 524 -458
rect 765 -459 766 -458
rect 37 -461 38 -460
rect 149 -461 150 -460
rect 212 -461 213 -460
rect 254 -461 255 -460
rect 261 -461 262 -460
rect 268 -461 269 -460
rect 303 -461 304 -460
rect 317 -461 318 -460
rect 418 -461 419 -460
rect 520 -461 521 -460
rect 541 -461 542 -460
rect 544 -461 545 -460
rect 558 -461 559 -460
rect 751 -461 752 -460
rect 765 -461 766 -460
rect 779 -461 780 -460
rect 110 -463 111 -462
rect 191 -463 192 -462
rect 222 -463 223 -462
rect 779 -463 780 -462
rect 135 -465 136 -464
rect 212 -465 213 -464
rect 247 -465 248 -464
rect 443 -465 444 -464
rect 541 -465 542 -464
rect 583 -465 584 -464
rect 590 -465 591 -464
rect 681 -465 682 -464
rect 688 -465 689 -464
rect 737 -465 738 -464
rect 149 -467 150 -466
rect 383 -467 384 -466
rect 562 -467 563 -466
rect 653 -467 654 -466
rect 705 -467 706 -466
rect 716 -467 717 -466
rect 247 -469 248 -468
rect 282 -469 283 -468
rect 303 -469 304 -468
rect 464 -469 465 -468
rect 492 -469 493 -468
rect 562 -469 563 -468
rect 569 -469 570 -468
rect 590 -469 591 -468
rect 282 -471 283 -470
rect 310 -471 311 -470
rect 380 -471 381 -470
rect 688 -471 689 -470
rect 16 -473 17 -472
rect 310 -473 311 -472
rect 422 -473 423 -472
rect 464 -473 465 -472
rect 492 -473 493 -472
rect 667 -473 668 -472
rect 16 -475 17 -474
rect 124 -475 125 -474
rect 422 -475 423 -474
rect 478 -475 479 -474
rect 548 -475 549 -474
rect 569 -475 570 -474
rect 576 -475 577 -474
rect 604 -475 605 -474
rect 415 -477 416 -476
rect 478 -477 479 -476
rect 527 -477 528 -476
rect 548 -477 549 -476
rect 555 -477 556 -476
rect 576 -477 577 -476
rect 408 -479 409 -478
rect 415 -479 416 -478
rect 485 -479 486 -478
rect 527 -479 528 -478
rect 485 -481 486 -480
rect 534 -481 535 -480
rect 457 -483 458 -482
rect 534 -483 535 -482
rect 457 -485 458 -484
rect 513 -485 514 -484
rect 499 -487 500 -486
rect 513 -487 514 -486
rect 331 -489 332 -488
rect 499 -489 500 -488
rect 156 -491 157 -490
rect 331 -491 332 -490
rect 156 -493 157 -492
rect 184 -493 185 -492
rect 142 -495 143 -494
rect 184 -495 185 -494
rect 142 -497 143 -496
rect 177 -497 178 -496
rect 23 -499 24 -498
rect 177 -499 178 -498
rect 23 -501 24 -500
rect 240 -501 241 -500
rect 65 -503 66 -502
rect 240 -503 241 -502
rect 65 -505 66 -504
rect 114 -505 115 -504
rect 114 -507 115 -506
rect 471 -507 472 -506
rect 9 -518 10 -517
rect 103 -518 104 -517
rect 163 -518 164 -517
rect 432 -518 433 -517
rect 467 -518 468 -517
rect 772 -518 773 -517
rect 793 -518 794 -517
rect 807 -518 808 -517
rect 9 -520 10 -519
rect 100 -520 101 -519
rect 163 -520 164 -519
rect 177 -520 178 -519
rect 184 -520 185 -519
rect 219 -520 220 -519
rect 222 -520 223 -519
rect 534 -520 535 -519
rect 555 -520 556 -519
rect 576 -520 577 -519
rect 583 -520 584 -519
rect 821 -520 822 -519
rect 16 -522 17 -521
rect 264 -522 265 -521
rect 313 -522 314 -521
rect 359 -522 360 -521
rect 380 -522 381 -521
rect 558 -522 559 -521
rect 618 -522 619 -521
rect 621 -522 622 -521
rect 779 -522 780 -521
rect 793 -522 794 -521
rect 800 -522 801 -521
rect 814 -522 815 -521
rect 16 -524 17 -523
rect 450 -524 451 -523
rect 471 -524 472 -523
rect 492 -524 493 -523
rect 495 -524 496 -523
rect 702 -524 703 -523
rect 758 -524 759 -523
rect 779 -524 780 -523
rect 786 -524 787 -523
rect 800 -524 801 -523
rect 44 -526 45 -525
rect 110 -526 111 -525
rect 135 -526 136 -525
rect 450 -526 451 -525
rect 457 -526 458 -525
rect 492 -526 493 -525
rect 520 -526 521 -525
rect 534 -526 535 -525
rect 541 -526 542 -525
rect 583 -526 584 -525
rect 618 -526 619 -525
rect 653 -526 654 -525
rect 744 -526 745 -525
rect 758 -526 759 -525
rect 765 -526 766 -525
rect 786 -526 787 -525
rect 47 -528 48 -527
rect 331 -528 332 -527
rect 383 -528 384 -527
rect 548 -528 549 -527
rect 621 -528 622 -527
rect 653 -528 654 -527
rect 54 -530 55 -529
rect 191 -530 192 -529
rect 226 -530 227 -529
rect 275 -530 276 -529
rect 303 -530 304 -529
rect 313 -530 314 -529
rect 317 -530 318 -529
rect 331 -530 332 -529
rect 383 -530 384 -529
rect 562 -530 563 -529
rect 625 -530 626 -529
rect 744 -530 745 -529
rect 58 -532 59 -531
rect 93 -532 94 -531
rect 131 -532 132 -531
rect 191 -532 192 -531
rect 212 -532 213 -531
rect 226 -532 227 -531
rect 233 -532 234 -531
rect 359 -532 360 -531
rect 387 -532 388 -531
rect 772 -532 773 -531
rect 61 -534 62 -533
rect 100 -534 101 -533
rect 121 -534 122 -533
rect 233 -534 234 -533
rect 240 -534 241 -533
rect 387 -534 388 -533
rect 390 -534 391 -533
rect 513 -534 514 -533
rect 520 -534 521 -533
rect 527 -534 528 -533
rect 541 -534 542 -533
rect 590 -534 591 -533
rect 625 -534 626 -533
rect 639 -534 640 -533
rect 79 -536 80 -535
rect 219 -536 220 -535
rect 240 -536 241 -535
rect 373 -536 374 -535
rect 394 -536 395 -535
rect 408 -536 409 -535
rect 429 -536 430 -535
rect 730 -536 731 -535
rect 79 -538 80 -537
rect 205 -538 206 -537
rect 257 -538 258 -537
rect 282 -538 283 -537
rect 310 -538 311 -537
rect 765 -538 766 -537
rect 51 -540 52 -539
rect 205 -540 206 -539
rect 275 -540 276 -539
rect 306 -540 307 -539
rect 345 -540 346 -539
rect 373 -540 374 -539
rect 401 -540 402 -539
rect 576 -540 577 -539
rect 639 -540 640 -539
rect 660 -540 661 -539
rect 30 -542 31 -541
rect 345 -542 346 -541
rect 401 -542 402 -541
rect 415 -542 416 -541
rect 422 -542 423 -541
rect 429 -542 430 -541
rect 457 -542 458 -541
rect 716 -542 717 -541
rect 30 -544 31 -543
rect 198 -544 199 -543
rect 282 -544 283 -543
rect 506 -544 507 -543
rect 562 -544 563 -543
rect 597 -544 598 -543
rect 86 -546 87 -545
rect 352 -546 353 -545
rect 369 -546 370 -545
rect 716 -546 717 -545
rect 86 -548 87 -547
rect 261 -548 262 -547
rect 317 -548 318 -547
rect 660 -548 661 -547
rect 93 -550 94 -549
rect 170 -550 171 -549
rect 177 -550 178 -549
rect 268 -550 269 -549
rect 415 -550 416 -549
rect 611 -550 612 -549
rect 114 -552 115 -551
rect 394 -552 395 -551
rect 422 -552 423 -551
rect 436 -552 437 -551
rect 474 -552 475 -551
rect 569 -552 570 -551
rect 597 -552 598 -551
rect 632 -552 633 -551
rect 23 -554 24 -553
rect 114 -554 115 -553
rect 135 -554 136 -553
rect 268 -554 269 -553
rect 436 -554 437 -553
rect 464 -554 465 -553
rect 478 -554 479 -553
rect 551 -554 552 -553
rect 569 -554 570 -553
rect 604 -554 605 -553
rect 611 -554 612 -553
rect 723 -554 724 -553
rect 23 -556 24 -555
rect 324 -556 325 -555
rect 411 -556 412 -555
rect 723 -556 724 -555
rect 149 -558 150 -557
rect 261 -558 262 -557
rect 324 -558 325 -557
rect 338 -558 339 -557
rect 443 -558 444 -557
rect 478 -558 479 -557
rect 485 -558 486 -557
rect 527 -558 528 -557
rect 604 -558 605 -557
rect 674 -558 675 -557
rect 72 -560 73 -559
rect 443 -560 444 -559
rect 488 -560 489 -559
rect 702 -560 703 -559
rect 142 -562 143 -561
rect 149 -562 150 -561
rect 156 -562 157 -561
rect 212 -562 213 -561
rect 296 -562 297 -561
rect 338 -562 339 -561
rect 499 -562 500 -561
rect 730 -562 731 -561
rect 37 -564 38 -563
rect 156 -564 157 -563
rect 170 -564 171 -563
rect 289 -564 290 -563
rect 464 -564 465 -563
rect 499 -564 500 -563
rect 506 -564 507 -563
rect 590 -564 591 -563
rect 632 -564 633 -563
rect 646 -564 647 -563
rect 674 -564 675 -563
rect 751 -564 752 -563
rect 37 -566 38 -565
rect 107 -566 108 -565
rect 198 -566 199 -565
rect 366 -566 367 -565
rect 646 -566 647 -565
rect 667 -566 668 -565
rect 737 -566 738 -565
rect 751 -566 752 -565
rect 65 -568 66 -567
rect 142 -568 143 -567
rect 289 -568 290 -567
rect 485 -568 486 -567
rect 667 -568 668 -567
rect 688 -568 689 -567
rect 65 -570 66 -569
rect 247 -570 248 -569
rect 418 -570 419 -569
rect 737 -570 738 -569
rect 128 -572 129 -571
rect 366 -572 367 -571
rect 688 -572 689 -571
rect 695 -572 696 -571
rect 72 -574 73 -573
rect 128 -574 129 -573
rect 247 -574 248 -573
rect 254 -574 255 -573
rect 334 -574 335 -573
rect 695 -574 696 -573
rect 184 -576 185 -575
rect 254 -576 255 -575
rect 2 -587 3 -586
rect 72 -587 73 -586
rect 107 -587 108 -586
rect 156 -587 157 -586
rect 163 -587 164 -586
rect 369 -587 370 -586
rect 457 -587 458 -586
rect 555 -587 556 -586
rect 9 -589 10 -588
rect 292 -589 293 -588
rect 296 -589 297 -588
rect 394 -589 395 -588
rect 464 -589 465 -588
rect 509 -589 510 -588
rect 513 -589 514 -588
rect 632 -589 633 -588
rect 9 -591 10 -590
rect 331 -591 332 -590
rect 334 -591 335 -590
rect 730 -591 731 -590
rect 54 -593 55 -592
rect 345 -593 346 -592
rect 467 -593 468 -592
rect 576 -593 577 -592
rect 730 -593 731 -592
rect 807 -593 808 -592
rect 68 -595 69 -594
rect 282 -595 283 -594
rect 299 -595 300 -594
rect 366 -595 367 -594
rect 485 -595 486 -594
rect 681 -595 682 -594
rect 72 -597 73 -596
rect 100 -597 101 -596
rect 107 -597 108 -596
rect 744 -597 745 -596
rect 100 -599 101 -598
rect 460 -599 461 -598
rect 506 -599 507 -598
rect 653 -599 654 -598
rect 110 -601 111 -600
rect 184 -601 185 -600
rect 205 -601 206 -600
rect 257 -601 258 -600
rect 271 -601 272 -600
rect 394 -601 395 -600
rect 460 -601 461 -600
rect 681 -601 682 -600
rect 110 -603 111 -602
rect 240 -603 241 -602
rect 254 -603 255 -602
rect 632 -603 633 -602
rect 653 -603 654 -602
rect 737 -603 738 -602
rect 121 -605 122 -604
rect 408 -605 409 -604
rect 506 -605 507 -604
rect 541 -605 542 -604
rect 576 -605 577 -604
rect 611 -605 612 -604
rect 737 -605 738 -604
rect 793 -605 794 -604
rect 121 -607 122 -606
rect 177 -607 178 -606
rect 184 -607 185 -606
rect 478 -607 479 -606
rect 513 -607 514 -606
rect 562 -607 563 -606
rect 611 -607 612 -606
rect 688 -607 689 -606
rect 26 -609 27 -608
rect 688 -609 689 -608
rect 124 -611 125 -610
rect 772 -611 773 -610
rect 128 -613 129 -612
rect 170 -613 171 -612
rect 177 -613 178 -612
rect 289 -613 290 -612
rect 303 -613 304 -612
rect 317 -613 318 -612
rect 320 -613 321 -612
rect 408 -613 409 -612
rect 478 -613 479 -612
rect 492 -613 493 -612
rect 534 -613 535 -612
rect 555 -613 556 -612
rect 562 -613 563 -612
rect 618 -613 619 -612
rect 772 -613 773 -612
rect 800 -613 801 -612
rect 138 -615 139 -614
rect 142 -615 143 -614
rect 149 -615 150 -614
rect 317 -615 318 -614
rect 331 -615 332 -614
rect 373 -615 374 -614
rect 492 -615 493 -614
rect 527 -615 528 -614
rect 534 -615 535 -614
rect 590 -615 591 -614
rect 618 -615 619 -614
rect 702 -615 703 -614
rect 37 -617 38 -616
rect 142 -617 143 -616
rect 156 -617 157 -616
rect 296 -617 297 -616
rect 303 -617 304 -616
rect 359 -617 360 -616
rect 366 -617 367 -616
rect 814 -617 815 -616
rect 30 -619 31 -618
rect 37 -619 38 -618
rect 61 -619 62 -618
rect 149 -619 150 -618
rect 163 -619 164 -618
rect 226 -619 227 -618
rect 240 -619 241 -618
rect 247 -619 248 -618
rect 282 -619 283 -618
rect 324 -619 325 -618
rect 359 -619 360 -618
rect 422 -619 423 -618
rect 527 -619 528 -618
rect 583 -619 584 -618
rect 590 -619 591 -618
rect 660 -619 661 -618
rect 702 -619 703 -618
rect 751 -619 752 -618
rect 170 -621 171 -620
rect 229 -621 230 -620
rect 289 -621 290 -620
rect 485 -621 486 -620
rect 583 -621 584 -620
rect 604 -621 605 -620
rect 751 -621 752 -620
rect 786 -621 787 -620
rect 191 -623 192 -622
rect 254 -623 255 -622
rect 310 -623 311 -622
rect 625 -623 626 -622
rect 191 -625 192 -624
rect 345 -625 346 -624
rect 348 -625 349 -624
rect 660 -625 661 -624
rect 205 -627 206 -626
rect 233 -627 234 -626
rect 275 -627 276 -626
rect 310 -627 311 -626
rect 324 -627 325 -626
rect 352 -627 353 -626
rect 373 -627 374 -626
rect 443 -627 444 -626
rect 453 -627 454 -626
rect 786 -627 787 -626
rect 198 -629 199 -628
rect 233 -629 234 -628
rect 268 -629 269 -628
rect 275 -629 276 -628
rect 338 -629 339 -628
rect 352 -629 353 -628
rect 422 -629 423 -628
rect 429 -629 430 -628
rect 443 -629 444 -628
rect 516 -629 517 -628
rect 548 -629 549 -628
rect 604 -629 605 -628
rect 625 -629 626 -628
rect 709 -629 710 -628
rect 65 -631 66 -630
rect 198 -631 199 -630
rect 212 -631 213 -630
rect 268 -631 269 -630
rect 338 -631 339 -630
rect 387 -631 388 -630
rect 548 -631 549 -630
rect 597 -631 598 -630
rect 709 -631 710 -630
rect 779 -631 780 -630
rect 30 -633 31 -632
rect 212 -633 213 -632
rect 215 -633 216 -632
rect 723 -633 724 -632
rect 758 -633 759 -632
rect 779 -633 780 -632
rect 219 -635 220 -634
rect 247 -635 248 -634
rect 380 -635 381 -634
rect 723 -635 724 -634
rect 758 -635 759 -634
rect 793 -635 794 -634
rect 51 -637 52 -636
rect 219 -637 220 -636
rect 226 -637 227 -636
rect 261 -637 262 -636
rect 383 -637 384 -636
rect 429 -637 430 -636
rect 597 -637 598 -636
rect 667 -637 668 -636
rect 44 -639 45 -638
rect 261 -639 262 -638
rect 383 -639 384 -638
rect 464 -639 465 -638
rect 646 -639 647 -638
rect 667 -639 668 -638
rect 44 -641 45 -640
rect 313 -641 314 -640
rect 387 -641 388 -640
rect 401 -641 402 -640
rect 646 -641 647 -640
rect 695 -641 696 -640
rect 16 -643 17 -642
rect 401 -643 402 -642
rect 499 -643 500 -642
rect 695 -643 696 -642
rect 16 -645 17 -644
rect 58 -645 59 -644
rect 499 -645 500 -644
rect 639 -645 640 -644
rect 58 -647 59 -646
rect 135 -647 136 -646
rect 639 -647 640 -646
rect 716 -647 717 -646
rect 79 -649 80 -648
rect 135 -649 136 -648
rect 674 -649 675 -648
rect 716 -649 717 -648
rect 79 -651 80 -650
rect 114 -651 115 -650
rect 674 -651 675 -650
rect 765 -651 766 -650
rect 23 -653 24 -652
rect 114 -653 115 -652
rect 415 -653 416 -652
rect 765 -653 766 -652
rect 23 -655 24 -654
rect 450 -655 451 -654
rect 415 -657 416 -656
rect 744 -657 745 -656
rect 450 -659 451 -658
rect 471 -659 472 -658
rect 471 -661 472 -660
rect 520 -661 521 -660
rect 520 -663 521 -662
rect 569 -663 570 -662
rect 569 -665 570 -664
rect 821 -665 822 -664
rect 2 -676 3 -675
rect 89 -676 90 -675
rect 142 -676 143 -675
rect 418 -676 419 -675
rect 425 -676 426 -675
rect 506 -676 507 -675
rect 520 -676 521 -675
rect 523 -676 524 -675
rect 551 -676 552 -675
rect 660 -676 661 -675
rect 779 -676 780 -675
rect 786 -676 787 -675
rect 16 -678 17 -677
rect 68 -678 69 -677
rect 142 -678 143 -677
rect 163 -678 164 -677
rect 184 -678 185 -677
rect 348 -678 349 -677
rect 415 -678 416 -677
rect 436 -678 437 -677
rect 446 -678 447 -677
rect 527 -678 528 -677
rect 660 -678 661 -677
rect 674 -678 675 -677
rect 779 -678 780 -677
rect 807 -678 808 -677
rect 16 -680 17 -679
rect 93 -680 94 -679
rect 107 -680 108 -679
rect 436 -680 437 -679
rect 450 -680 451 -679
rect 485 -680 486 -679
rect 499 -680 500 -679
rect 502 -680 503 -679
rect 527 -680 528 -679
rect 709 -680 710 -679
rect 51 -682 52 -681
rect 86 -682 87 -681
rect 107 -682 108 -681
rect 268 -682 269 -681
rect 271 -682 272 -681
rect 667 -682 668 -681
rect 37 -684 38 -683
rect 51 -684 52 -683
rect 58 -684 59 -683
rect 121 -684 122 -683
rect 149 -684 150 -683
rect 184 -684 185 -683
rect 212 -684 213 -683
rect 317 -684 318 -683
rect 415 -684 416 -683
rect 429 -684 430 -683
rect 453 -684 454 -683
rect 653 -684 654 -683
rect 9 -686 10 -685
rect 317 -686 318 -685
rect 457 -686 458 -685
rect 464 -686 465 -685
rect 471 -686 472 -685
rect 800 -686 801 -685
rect 37 -688 38 -687
rect 79 -688 80 -687
rect 93 -688 94 -687
rect 271 -688 272 -687
rect 296 -688 297 -687
rect 772 -688 773 -687
rect 61 -690 62 -689
rect 170 -690 171 -689
rect 198 -690 199 -689
rect 296 -690 297 -689
rect 310 -690 311 -689
rect 429 -690 430 -689
rect 443 -690 444 -689
rect 471 -690 472 -689
rect 485 -690 486 -689
rect 492 -690 493 -689
rect 499 -690 500 -689
rect 513 -690 514 -689
rect 604 -690 605 -689
rect 667 -690 668 -689
rect 772 -690 773 -689
rect 793 -690 794 -689
rect 12 -692 13 -691
rect 310 -692 311 -691
rect 443 -692 444 -691
rect 737 -692 738 -691
rect 68 -694 69 -693
rect 79 -694 80 -693
rect 114 -694 115 -693
rect 121 -694 122 -693
rect 135 -694 136 -693
rect 149 -694 150 -693
rect 170 -694 171 -693
rect 261 -694 262 -693
rect 268 -694 269 -693
rect 366 -694 367 -693
rect 460 -694 461 -693
rect 737 -694 738 -693
rect 72 -696 73 -695
rect 163 -696 164 -695
rect 198 -696 199 -695
rect 240 -696 241 -695
rect 261 -696 262 -695
rect 303 -696 304 -695
rect 464 -696 465 -695
rect 534 -696 535 -695
rect 583 -696 584 -695
rect 604 -696 605 -695
rect 646 -696 647 -695
rect 674 -696 675 -695
rect 23 -698 24 -697
rect 72 -698 73 -697
rect 114 -698 115 -697
rect 128 -698 129 -697
rect 135 -698 136 -697
rect 229 -698 230 -697
rect 233 -698 234 -697
rect 289 -698 290 -697
rect 303 -698 304 -697
rect 369 -698 370 -697
rect 492 -698 493 -697
rect 569 -698 570 -697
rect 583 -698 584 -697
rect 611 -698 612 -697
rect 646 -698 647 -697
rect 702 -698 703 -697
rect 23 -700 24 -699
rect 191 -700 192 -699
rect 212 -700 213 -699
rect 254 -700 255 -699
rect 513 -700 514 -699
rect 555 -700 556 -699
rect 590 -700 591 -699
rect 611 -700 612 -699
rect 618 -700 619 -699
rect 702 -700 703 -699
rect 44 -702 45 -701
rect 128 -702 129 -701
rect 191 -702 192 -701
rect 205 -702 206 -701
rect 226 -702 227 -701
rect 709 -702 710 -701
rect 44 -704 45 -703
rect 65 -704 66 -703
rect 205 -704 206 -703
rect 219 -704 220 -703
rect 229 -704 230 -703
rect 380 -704 381 -703
rect 534 -704 535 -703
rect 782 -704 783 -703
rect 30 -706 31 -705
rect 65 -706 66 -705
rect 219 -706 220 -705
rect 408 -706 409 -705
rect 544 -706 545 -705
rect 590 -706 591 -705
rect 618 -706 619 -705
rect 688 -706 689 -705
rect 30 -708 31 -707
rect 324 -708 325 -707
rect 345 -708 346 -707
rect 408 -708 409 -707
rect 555 -708 556 -707
rect 562 -708 563 -707
rect 597 -708 598 -707
rect 688 -708 689 -707
rect 233 -710 234 -709
rect 247 -710 248 -709
rect 254 -710 255 -709
rect 338 -710 339 -709
rect 380 -710 381 -709
rect 695 -710 696 -709
rect 240 -712 241 -711
rect 275 -712 276 -711
rect 324 -712 325 -711
rect 359 -712 360 -711
rect 502 -712 503 -711
rect 562 -712 563 -711
rect 597 -712 598 -711
rect 632 -712 633 -711
rect 653 -712 654 -711
rect 681 -712 682 -711
rect 695 -712 696 -711
rect 716 -712 717 -711
rect 166 -714 167 -713
rect 359 -714 360 -713
rect 478 -714 479 -713
rect 716 -714 717 -713
rect 247 -716 248 -715
rect 331 -716 332 -715
rect 338 -716 339 -715
rect 352 -716 353 -715
rect 478 -716 479 -715
rect 548 -716 549 -715
rect 576 -716 577 -715
rect 632 -716 633 -715
rect 681 -716 682 -715
rect 723 -716 724 -715
rect 275 -718 276 -717
rect 282 -718 283 -717
rect 331 -718 332 -717
rect 387 -718 388 -717
rect 530 -718 531 -717
rect 576 -718 577 -717
rect 723 -718 724 -717
rect 744 -718 745 -717
rect 282 -720 283 -719
rect 394 -720 395 -719
rect 744 -720 745 -719
rect 758 -720 759 -719
rect 320 -722 321 -721
rect 387 -722 388 -721
rect 394 -722 395 -721
rect 506 -722 507 -721
rect 730 -722 731 -721
rect 758 -722 759 -721
rect 131 -724 132 -723
rect 730 -724 731 -723
rect 352 -726 353 -725
rect 373 -726 374 -725
rect 373 -728 374 -727
rect 401 -728 402 -727
rect 401 -730 402 -729
rect 422 -730 423 -729
rect 422 -732 423 -731
rect 541 -732 542 -731
rect 2 -743 3 -742
rect 226 -743 227 -742
rect 268 -743 269 -742
rect 275 -743 276 -742
rect 289 -743 290 -742
rect 348 -743 349 -742
rect 397 -743 398 -742
rect 464 -743 465 -742
rect 481 -743 482 -742
rect 569 -743 570 -742
rect 572 -743 573 -742
rect 737 -743 738 -742
rect 782 -743 783 -742
rect 786 -743 787 -742
rect 793 -743 794 -742
rect 807 -743 808 -742
rect 9 -745 10 -744
rect 128 -745 129 -744
rect 166 -745 167 -744
rect 219 -745 220 -744
rect 268 -745 269 -744
rect 387 -745 388 -744
rect 422 -745 423 -744
rect 702 -745 703 -744
rect 737 -745 738 -744
rect 744 -745 745 -744
rect 16 -747 17 -746
rect 58 -747 59 -746
rect 65 -747 66 -746
rect 72 -747 73 -746
rect 79 -747 80 -746
rect 317 -747 318 -746
rect 345 -747 346 -746
rect 688 -747 689 -746
rect 702 -747 703 -746
rect 723 -747 724 -746
rect 744 -747 745 -746
rect 751 -747 752 -746
rect 30 -749 31 -748
rect 229 -749 230 -748
rect 275 -749 276 -748
rect 296 -749 297 -748
rect 310 -749 311 -748
rect 345 -749 346 -748
rect 366 -749 367 -748
rect 464 -749 465 -748
rect 506 -749 507 -748
rect 569 -749 570 -748
rect 576 -749 577 -748
rect 786 -749 787 -748
rect 19 -751 20 -750
rect 366 -751 367 -750
rect 376 -751 377 -750
rect 506 -751 507 -750
rect 520 -751 521 -750
rect 555 -751 556 -750
rect 600 -751 601 -750
rect 660 -751 661 -750
rect 751 -751 752 -750
rect 758 -751 759 -750
rect 30 -753 31 -752
rect 44 -753 45 -752
rect 58 -753 59 -752
rect 121 -753 122 -752
rect 184 -753 185 -752
rect 215 -753 216 -752
rect 233 -753 234 -752
rect 296 -753 297 -752
rect 310 -753 311 -752
rect 352 -753 353 -752
rect 380 -753 381 -752
rect 688 -753 689 -752
rect 758 -753 759 -752
rect 772 -753 773 -752
rect 40 -755 41 -754
rect 163 -755 164 -754
rect 184 -755 185 -754
rect 212 -755 213 -754
rect 282 -755 283 -754
rect 387 -755 388 -754
rect 408 -755 409 -754
rect 422 -755 423 -754
rect 446 -755 447 -754
rect 723 -755 724 -754
rect 772 -755 773 -754
rect 779 -755 780 -754
rect 44 -757 45 -756
rect 411 -757 412 -756
rect 450 -757 451 -756
rect 453 -757 454 -756
rect 530 -757 531 -756
rect 639 -757 640 -756
rect 72 -759 73 -758
rect 177 -759 178 -758
rect 198 -759 199 -758
rect 201 -759 202 -758
rect 205 -759 206 -758
rect 219 -759 220 -758
rect 247 -759 248 -758
rect 282 -759 283 -758
rect 289 -759 290 -758
rect 373 -759 374 -758
rect 450 -759 451 -758
rect 492 -759 493 -758
rect 541 -759 542 -758
rect 576 -759 577 -758
rect 618 -759 619 -758
rect 660 -759 661 -758
rect 75 -761 76 -760
rect 205 -761 206 -760
rect 233 -761 234 -760
rect 247 -761 248 -760
rect 320 -761 321 -760
rect 618 -761 619 -760
rect 632 -761 633 -760
rect 639 -761 640 -760
rect 79 -763 80 -762
rect 303 -763 304 -762
rect 331 -763 332 -762
rect 352 -763 353 -762
rect 359 -763 360 -762
rect 380 -763 381 -762
rect 485 -763 486 -762
rect 492 -763 493 -762
rect 534 -763 535 -762
rect 541 -763 542 -762
rect 548 -763 549 -762
rect 604 -763 605 -762
rect 86 -765 87 -764
rect 383 -765 384 -764
rect 471 -765 472 -764
rect 534 -765 535 -764
rect 551 -765 552 -764
rect 667 -765 668 -764
rect 86 -767 87 -766
rect 100 -767 101 -766
rect 107 -767 108 -766
rect 121 -767 122 -766
rect 177 -767 178 -766
rect 261 -767 262 -766
rect 303 -767 304 -766
rect 338 -767 339 -766
rect 359 -767 360 -766
rect 457 -767 458 -766
rect 471 -767 472 -766
rect 478 -767 479 -766
rect 555 -767 556 -766
rect 590 -767 591 -766
rect 597 -767 598 -766
rect 632 -767 633 -766
rect 667 -767 668 -766
rect 695 -767 696 -766
rect 89 -769 90 -768
rect 681 -769 682 -768
rect 695 -769 696 -768
rect 709 -769 710 -768
rect 93 -771 94 -770
rect 317 -771 318 -770
rect 324 -771 325 -770
rect 338 -771 339 -770
rect 362 -771 363 -770
rect 590 -771 591 -770
rect 646 -771 647 -770
rect 681 -771 682 -770
rect 23 -773 24 -772
rect 93 -773 94 -772
rect 100 -773 101 -772
rect 149 -773 150 -772
rect 170 -773 171 -772
rect 261 -773 262 -772
rect 373 -773 374 -772
rect 716 -773 717 -772
rect 23 -775 24 -774
rect 135 -775 136 -774
rect 149 -775 150 -774
rect 191 -775 192 -774
rect 198 -775 199 -774
rect 240 -775 241 -774
rect 254 -775 255 -774
rect 324 -775 325 -774
rect 404 -775 405 -774
rect 597 -775 598 -774
rect 646 -775 647 -774
rect 674 -775 675 -774
rect 716 -775 717 -774
rect 730 -775 731 -774
rect 51 -777 52 -776
rect 170 -777 171 -776
rect 191 -777 192 -776
rect 443 -777 444 -776
rect 453 -777 454 -776
rect 485 -777 486 -776
rect 548 -777 549 -776
rect 730 -777 731 -776
rect 51 -779 52 -778
rect 425 -779 426 -778
rect 443 -779 444 -778
rect 527 -779 528 -778
rect 583 -779 584 -778
rect 604 -779 605 -778
rect 107 -781 108 -780
rect 114 -781 115 -780
rect 135 -781 136 -780
rect 142 -781 143 -780
rect 159 -781 160 -780
rect 527 -781 528 -780
rect 37 -783 38 -782
rect 114 -783 115 -782
rect 142 -783 143 -782
rect 156 -783 157 -782
rect 212 -783 213 -782
rect 331 -783 332 -782
rect 457 -783 458 -782
rect 800 -783 801 -782
rect 37 -785 38 -784
rect 611 -785 612 -784
rect 254 -787 255 -786
rect 674 -787 675 -786
rect 285 -789 286 -788
rect 611 -789 612 -788
rect 478 -791 479 -790
rect 709 -791 710 -790
rect 499 -793 500 -792
rect 583 -793 584 -792
rect 436 -795 437 -794
rect 499 -795 500 -794
rect 429 -797 430 -796
rect 436 -797 437 -796
rect 415 -799 416 -798
rect 429 -799 430 -798
rect 401 -801 402 -800
rect 415 -801 416 -800
rect 68 -803 69 -802
rect 401 -803 402 -802
rect 23 -814 24 -813
rect 156 -814 157 -813
rect 170 -814 171 -813
rect 250 -814 251 -813
rect 254 -814 255 -813
rect 275 -814 276 -813
rect 282 -814 283 -813
rect 296 -814 297 -813
rect 310 -814 311 -813
rect 380 -814 381 -813
rect 394 -814 395 -813
rect 429 -814 430 -813
rect 478 -814 479 -813
rect 527 -814 528 -813
rect 544 -814 545 -813
rect 681 -814 682 -813
rect 9 -816 10 -815
rect 23 -816 24 -815
rect 30 -816 31 -815
rect 40 -816 41 -815
rect 65 -816 66 -815
rect 131 -816 132 -815
rect 156 -816 157 -815
rect 233 -816 234 -815
rect 240 -816 241 -815
rect 257 -816 258 -815
rect 271 -816 272 -815
rect 443 -816 444 -815
rect 481 -816 482 -815
rect 562 -816 563 -815
rect 597 -816 598 -815
rect 744 -816 745 -815
rect 9 -818 10 -817
rect 128 -818 129 -817
rect 177 -818 178 -817
rect 212 -818 213 -817
rect 219 -818 220 -817
rect 222 -818 223 -817
rect 226 -818 227 -817
rect 376 -818 377 -817
rect 397 -818 398 -817
rect 485 -818 486 -817
rect 513 -818 514 -817
rect 527 -818 528 -817
rect 548 -818 549 -817
rect 646 -818 647 -817
rect 744 -818 745 -817
rect 786 -818 787 -817
rect 16 -820 17 -819
rect 65 -820 66 -819
rect 72 -820 73 -819
rect 86 -820 87 -819
rect 93 -820 94 -819
rect 226 -820 227 -819
rect 240 -820 241 -819
rect 422 -820 423 -819
rect 429 -820 430 -819
rect 457 -820 458 -819
rect 485 -820 486 -819
rect 569 -820 570 -819
rect 618 -820 619 -819
rect 765 -820 766 -819
rect 86 -822 87 -821
rect 114 -822 115 -821
rect 117 -822 118 -821
rect 159 -822 160 -821
rect 184 -822 185 -821
rect 233 -822 234 -821
rect 275 -822 276 -821
rect 331 -822 332 -821
rect 345 -822 346 -821
rect 401 -822 402 -821
rect 408 -822 409 -821
rect 502 -822 503 -821
rect 513 -822 514 -821
rect 520 -822 521 -821
rect 548 -822 549 -821
rect 604 -822 605 -821
rect 618 -822 619 -821
rect 702 -822 703 -821
rect 75 -824 76 -823
rect 114 -824 115 -823
rect 121 -824 122 -823
rect 128 -824 129 -823
rect 135 -824 136 -823
rect 177 -824 178 -823
rect 184 -824 185 -823
rect 205 -824 206 -823
rect 219 -824 220 -823
rect 303 -824 304 -823
rect 331 -824 332 -823
rect 338 -824 339 -823
rect 345 -824 346 -823
rect 590 -824 591 -823
rect 646 -824 647 -823
rect 716 -824 717 -823
rect 93 -826 94 -825
rect 107 -826 108 -825
rect 110 -826 111 -825
rect 191 -826 192 -825
rect 205 -826 206 -825
rect 268 -826 269 -825
rect 282 -826 283 -825
rect 436 -826 437 -825
rect 443 -826 444 -825
rect 506 -826 507 -825
rect 562 -826 563 -825
rect 611 -826 612 -825
rect 702 -826 703 -825
rect 751 -826 752 -825
rect 72 -828 73 -827
rect 107 -828 108 -827
rect 121 -828 122 -827
rect 149 -828 150 -827
rect 191 -828 192 -827
rect 324 -828 325 -827
rect 338 -828 339 -827
rect 387 -828 388 -827
rect 404 -828 405 -827
rect 506 -828 507 -827
rect 569 -828 570 -827
rect 632 -828 633 -827
rect 751 -828 752 -827
rect 758 -828 759 -827
rect 79 -830 80 -829
rect 268 -830 269 -829
rect 296 -830 297 -829
rect 317 -830 318 -829
rect 348 -830 349 -829
rect 688 -830 689 -829
rect 758 -830 759 -829
rect 779 -830 780 -829
rect 51 -832 52 -831
rect 79 -832 80 -831
rect 100 -832 101 -831
rect 149 -832 150 -831
rect 163 -832 164 -831
rect 317 -832 318 -831
rect 359 -832 360 -831
rect 390 -832 391 -831
rect 411 -832 412 -831
rect 583 -832 584 -831
rect 590 -832 591 -831
rect 639 -832 640 -831
rect 688 -832 689 -831
rect 726 -832 727 -831
rect 30 -834 31 -833
rect 51 -834 52 -833
rect 142 -834 143 -833
rect 163 -834 164 -833
rect 222 -834 223 -833
rect 303 -834 304 -833
rect 366 -834 367 -833
rect 520 -834 521 -833
rect 583 -834 584 -833
rect 653 -834 654 -833
rect 44 -836 45 -835
rect 100 -836 101 -835
rect 247 -836 248 -835
rect 387 -836 388 -835
rect 422 -836 423 -835
rect 492 -836 493 -835
rect 611 -836 612 -835
rect 674 -836 675 -835
rect 44 -838 45 -837
rect 138 -838 139 -837
rect 198 -838 199 -837
rect 247 -838 248 -837
rect 324 -838 325 -837
rect 366 -838 367 -837
rect 373 -838 374 -837
rect 597 -838 598 -837
rect 632 -838 633 -837
rect 660 -838 661 -837
rect 58 -840 59 -839
rect 142 -840 143 -839
rect 198 -840 199 -839
rect 289 -840 290 -839
rect 373 -840 374 -839
rect 464 -840 465 -839
rect 492 -840 493 -839
rect 607 -840 608 -839
rect 639 -840 640 -839
rect 667 -840 668 -839
rect 58 -842 59 -841
rect 173 -842 174 -841
rect 264 -842 265 -841
rect 464 -842 465 -841
rect 653 -842 654 -841
rect 695 -842 696 -841
rect 289 -844 290 -843
rect 352 -844 353 -843
rect 380 -844 381 -843
rect 660 -844 661 -843
rect 667 -844 668 -843
rect 723 -844 724 -843
rect 352 -846 353 -845
rect 415 -846 416 -845
rect 436 -846 437 -845
rect 471 -846 472 -845
rect 695 -846 696 -845
rect 730 -846 731 -845
rect 415 -848 416 -847
rect 541 -848 542 -847
rect 457 -850 458 -849
rect 534 -850 535 -849
rect 471 -852 472 -851
rect 499 -852 500 -851
rect 534 -852 535 -851
rect 555 -852 556 -851
rect 555 -854 556 -853
rect 576 -854 577 -853
rect 576 -856 577 -855
rect 625 -856 626 -855
rect 625 -858 626 -857
rect 709 -858 710 -857
rect 9 -869 10 -868
rect 397 -869 398 -868
rect 471 -869 472 -868
rect 523 -869 524 -868
rect 544 -869 545 -868
rect 583 -869 584 -868
rect 604 -869 605 -868
rect 730 -869 731 -868
rect 733 -869 734 -868
rect 737 -869 738 -868
rect 747 -869 748 -868
rect 751 -869 752 -868
rect 19 -871 20 -870
rect 23 -871 24 -870
rect 51 -871 52 -870
rect 93 -871 94 -870
rect 114 -871 115 -870
rect 117 -871 118 -870
rect 124 -871 125 -870
rect 478 -871 479 -870
rect 499 -871 500 -870
rect 534 -871 535 -870
rect 583 -871 584 -870
rect 597 -871 598 -870
rect 604 -871 605 -870
rect 639 -871 640 -870
rect 663 -871 664 -870
rect 688 -871 689 -870
rect 726 -871 727 -870
rect 758 -871 759 -870
rect 54 -873 55 -872
rect 107 -873 108 -872
rect 135 -873 136 -872
rect 177 -873 178 -872
rect 180 -873 181 -872
rect 275 -873 276 -872
rect 282 -873 283 -872
rect 383 -873 384 -872
rect 387 -873 388 -872
rect 422 -873 423 -872
rect 502 -873 503 -872
rect 632 -873 633 -872
rect 674 -873 675 -872
rect 702 -873 703 -872
rect 30 -875 31 -874
rect 282 -875 283 -874
rect 317 -875 318 -874
rect 380 -875 381 -874
rect 390 -875 391 -874
rect 450 -875 451 -874
rect 520 -875 521 -874
rect 597 -875 598 -874
rect 632 -875 633 -874
rect 646 -875 647 -874
rect 681 -875 682 -874
rect 744 -875 745 -874
rect 58 -877 59 -876
rect 177 -877 178 -876
rect 212 -877 213 -876
rect 299 -877 300 -876
rect 317 -877 318 -876
rect 338 -877 339 -876
rect 345 -877 346 -876
rect 541 -877 542 -876
rect 642 -877 643 -876
rect 646 -877 647 -876
rect 681 -877 682 -876
rect 695 -877 696 -876
rect 58 -879 59 -878
rect 86 -879 87 -878
rect 93 -879 94 -878
rect 110 -879 111 -878
rect 121 -879 122 -878
rect 135 -879 136 -878
rect 142 -879 143 -878
rect 145 -879 146 -878
rect 149 -879 150 -878
rect 170 -879 171 -878
rect 257 -879 258 -878
rect 303 -879 304 -878
rect 352 -879 353 -878
rect 369 -879 370 -878
rect 401 -879 402 -878
rect 422 -879 423 -878
rect 450 -879 451 -878
rect 527 -879 528 -878
rect 534 -879 535 -878
rect 576 -879 577 -878
rect 684 -879 685 -878
rect 716 -879 717 -878
rect 65 -881 66 -880
rect 348 -881 349 -880
rect 352 -881 353 -880
rect 394 -881 395 -880
rect 401 -881 402 -880
rect 443 -881 444 -880
rect 527 -881 528 -880
rect 569 -881 570 -880
rect 576 -881 577 -880
rect 618 -881 619 -880
rect 65 -883 66 -882
rect 219 -883 220 -882
rect 261 -883 262 -882
rect 373 -883 374 -882
rect 394 -883 395 -882
rect 653 -883 654 -882
rect 79 -885 80 -884
rect 149 -885 150 -884
rect 170 -885 171 -884
rect 310 -885 311 -884
rect 366 -885 367 -884
rect 443 -885 444 -884
rect 492 -885 493 -884
rect 569 -885 570 -884
rect 618 -885 619 -884
rect 667 -885 668 -884
rect 79 -887 80 -886
rect 240 -887 241 -886
rect 271 -887 272 -886
rect 296 -887 297 -886
rect 303 -887 304 -886
rect 331 -887 332 -886
rect 373 -887 374 -886
rect 478 -887 479 -886
rect 541 -887 542 -886
rect 562 -887 563 -886
rect 86 -889 87 -888
rect 138 -889 139 -888
rect 142 -889 143 -888
rect 191 -889 192 -888
rect 198 -889 199 -888
rect 240 -889 241 -888
rect 271 -889 272 -888
rect 376 -889 377 -888
rect 464 -889 465 -888
rect 492 -889 493 -888
rect 555 -889 556 -888
rect 667 -889 668 -888
rect 100 -891 101 -890
rect 212 -891 213 -890
rect 219 -891 220 -890
rect 254 -891 255 -890
rect 275 -891 276 -890
rect 324 -891 325 -890
rect 331 -891 332 -890
rect 436 -891 437 -890
rect 562 -891 563 -890
rect 590 -891 591 -890
rect 72 -893 73 -892
rect 100 -893 101 -892
rect 107 -893 108 -892
rect 128 -893 129 -892
rect 145 -893 146 -892
rect 191 -893 192 -892
rect 198 -893 199 -892
rect 233 -893 234 -892
rect 289 -893 290 -892
rect 338 -893 339 -892
rect 415 -893 416 -892
rect 436 -893 437 -892
rect 590 -893 591 -892
rect 611 -893 612 -892
rect 72 -895 73 -894
rect 226 -895 227 -894
rect 289 -895 290 -894
rect 408 -895 409 -894
rect 415 -895 416 -894
rect 467 -895 468 -894
rect 611 -895 612 -894
rect 625 -895 626 -894
rect 40 -897 41 -896
rect 226 -897 227 -896
rect 310 -897 311 -896
rect 359 -897 360 -896
rect 408 -897 409 -896
rect 429 -897 430 -896
rect 625 -897 626 -896
rect 660 -897 661 -896
rect 128 -899 129 -898
rect 156 -899 157 -898
rect 173 -899 174 -898
rect 555 -899 556 -898
rect 156 -901 157 -900
rect 359 -901 360 -900
rect 429 -901 430 -900
rect 457 -901 458 -900
rect 506 -901 507 -900
rect 660 -901 661 -900
rect 184 -903 185 -902
rect 233 -903 234 -902
rect 457 -903 458 -902
rect 485 -903 486 -902
rect 506 -903 507 -902
rect 548 -903 549 -902
rect 184 -905 185 -904
rect 247 -905 248 -904
rect 296 -905 297 -904
rect 548 -905 549 -904
rect 44 -907 45 -906
rect 247 -907 248 -906
rect 485 -907 486 -906
rect 513 -907 514 -906
rect 44 -909 45 -908
rect 205 -909 206 -908
rect 208 -909 209 -908
rect 513 -909 514 -908
rect 205 -911 206 -910
rect 471 -911 472 -910
rect 44 -922 45 -921
rect 453 -922 454 -921
rect 464 -922 465 -921
rect 492 -922 493 -921
rect 520 -922 521 -921
rect 576 -922 577 -921
rect 646 -922 647 -921
rect 653 -922 654 -921
rect 660 -922 661 -921
rect 674 -922 675 -921
rect 716 -922 717 -921
rect 744 -922 745 -921
rect 51 -924 52 -923
rect 121 -924 122 -923
rect 170 -924 171 -923
rect 177 -924 178 -923
rect 191 -924 192 -923
rect 205 -924 206 -923
rect 219 -924 220 -923
rect 268 -924 269 -923
rect 282 -924 283 -923
rect 313 -924 314 -923
rect 320 -924 321 -923
rect 422 -924 423 -923
rect 464 -924 465 -923
rect 555 -924 556 -923
rect 674 -924 675 -923
rect 681 -924 682 -923
rect 72 -926 73 -925
rect 93 -926 94 -925
rect 103 -926 104 -925
rect 121 -926 122 -925
rect 142 -926 143 -925
rect 219 -926 220 -925
rect 226 -926 227 -925
rect 425 -926 426 -925
rect 492 -926 493 -925
rect 569 -926 570 -925
rect 107 -928 108 -927
rect 156 -928 157 -927
rect 159 -928 160 -927
rect 170 -928 171 -927
rect 184 -928 185 -927
rect 205 -928 206 -927
rect 240 -928 241 -927
rect 324 -928 325 -927
rect 394 -928 395 -927
rect 429 -928 430 -927
rect 499 -928 500 -927
rect 576 -928 577 -927
rect 86 -930 87 -929
rect 107 -930 108 -929
rect 128 -930 129 -929
rect 142 -930 143 -929
rect 184 -930 185 -929
rect 233 -930 234 -929
rect 240 -930 241 -929
rect 352 -930 353 -929
rect 499 -930 500 -929
rect 618 -930 619 -929
rect 58 -932 59 -931
rect 86 -932 87 -931
rect 100 -932 101 -931
rect 128 -932 129 -931
rect 191 -932 192 -931
rect 366 -932 367 -931
rect 527 -932 528 -931
rect 569 -932 570 -931
rect 618 -932 619 -931
rect 639 -932 640 -931
rect 114 -934 115 -933
rect 233 -934 234 -933
rect 254 -934 255 -933
rect 429 -934 430 -933
rect 450 -934 451 -933
rect 527 -934 528 -933
rect 541 -934 542 -933
rect 642 -934 643 -933
rect 198 -936 199 -935
rect 541 -936 542 -935
rect 555 -936 556 -935
rect 611 -936 612 -935
rect 149 -938 150 -937
rect 198 -938 199 -937
rect 254 -938 255 -937
rect 436 -938 437 -937
rect 534 -938 535 -937
rect 611 -938 612 -937
rect 149 -940 150 -939
rect 226 -940 227 -939
rect 268 -940 269 -939
rect 317 -940 318 -939
rect 324 -940 325 -939
rect 471 -940 472 -939
rect 156 -942 157 -941
rect 317 -942 318 -941
rect 352 -942 353 -941
rect 415 -942 416 -941
rect 436 -942 437 -941
rect 457 -942 458 -941
rect 471 -942 472 -941
rect 485 -942 486 -941
rect 275 -944 276 -943
rect 282 -944 283 -943
rect 289 -944 290 -943
rect 299 -944 300 -943
rect 310 -944 311 -943
rect 544 -944 545 -943
rect 79 -946 80 -945
rect 289 -946 290 -945
rect 296 -946 297 -945
rect 338 -946 339 -945
rect 366 -946 367 -945
rect 632 -946 633 -945
rect 79 -948 80 -947
rect 303 -948 304 -947
rect 338 -948 339 -947
rect 359 -948 360 -947
rect 408 -948 409 -947
rect 534 -948 535 -947
rect 275 -950 276 -949
rect 345 -950 346 -949
rect 359 -950 360 -949
rect 380 -950 381 -949
rect 408 -950 409 -949
rect 443 -950 444 -949
rect 457 -950 458 -949
rect 583 -950 584 -949
rect 247 -952 248 -951
rect 345 -952 346 -951
rect 380 -952 381 -951
rect 387 -952 388 -951
rect 443 -952 444 -951
rect 513 -952 514 -951
rect 583 -952 584 -951
rect 597 -952 598 -951
rect 212 -954 213 -953
rect 247 -954 248 -953
rect 303 -954 304 -953
rect 369 -954 370 -953
rect 478 -954 479 -953
rect 485 -954 486 -953
rect 513 -954 514 -953
rect 562 -954 563 -953
rect 65 -956 66 -955
rect 212 -956 213 -955
rect 331 -956 332 -955
rect 597 -956 598 -955
rect 65 -958 66 -957
rect 257 -958 258 -957
rect 261 -958 262 -957
rect 331 -958 332 -957
rect 478 -958 479 -957
rect 548 -958 549 -957
rect 261 -960 262 -959
rect 401 -960 402 -959
rect 506 -960 507 -959
rect 562 -960 563 -959
rect 373 -962 374 -961
rect 401 -962 402 -961
rect 506 -962 507 -961
rect 628 -962 629 -961
rect 548 -964 549 -963
rect 590 -964 591 -963
rect 590 -966 591 -965
rect 625 -966 626 -965
rect 604 -968 605 -967
rect 625 -968 626 -967
rect 604 -970 605 -969
rect 667 -970 668 -969
rect 65 -981 66 -980
rect 229 -981 230 -980
rect 254 -981 255 -980
rect 418 -981 419 -980
rect 422 -981 423 -980
rect 492 -981 493 -980
rect 523 -981 524 -980
rect 527 -981 528 -980
rect 544 -981 545 -980
rect 569 -981 570 -980
rect 576 -981 577 -980
rect 579 -981 580 -980
rect 607 -981 608 -980
rect 611 -981 612 -980
rect 649 -981 650 -980
rect 660 -981 661 -980
rect 670 -981 671 -980
rect 674 -981 675 -980
rect 72 -983 73 -982
rect 96 -983 97 -982
rect 100 -983 101 -982
rect 250 -983 251 -982
rect 254 -983 255 -982
rect 362 -983 363 -982
rect 373 -983 374 -982
rect 443 -983 444 -982
rect 453 -983 454 -982
rect 499 -983 500 -982
rect 527 -983 528 -982
rect 534 -983 535 -982
rect 555 -983 556 -982
rect 569 -983 570 -982
rect 576 -983 577 -982
rect 590 -983 591 -982
rect 611 -983 612 -982
rect 618 -983 619 -982
rect 79 -985 80 -984
rect 198 -985 199 -984
rect 212 -985 213 -984
rect 369 -985 370 -984
rect 380 -985 381 -984
rect 446 -985 447 -984
rect 471 -985 472 -984
rect 499 -985 500 -984
rect 579 -985 580 -984
rect 590 -985 591 -984
rect 93 -987 94 -986
rect 100 -987 101 -986
rect 107 -987 108 -986
rect 128 -987 129 -986
rect 170 -987 171 -986
rect 201 -987 202 -986
rect 264 -987 265 -986
rect 324 -987 325 -986
rect 352 -987 353 -986
rect 390 -987 391 -986
rect 394 -987 395 -986
rect 422 -987 423 -986
rect 425 -987 426 -986
rect 436 -987 437 -986
rect 439 -987 440 -986
rect 506 -987 507 -986
rect 86 -989 87 -988
rect 170 -989 171 -988
rect 191 -989 192 -988
rect 226 -989 227 -988
rect 240 -989 241 -988
rect 352 -989 353 -988
rect 369 -989 370 -988
rect 597 -989 598 -988
rect 117 -991 118 -990
rect 121 -991 122 -990
rect 177 -991 178 -990
rect 240 -991 241 -990
rect 268 -991 269 -990
rect 373 -991 374 -990
rect 380 -991 381 -990
rect 450 -991 451 -990
rect 492 -991 493 -990
rect 513 -991 514 -990
rect 163 -993 164 -992
rect 177 -993 178 -992
rect 184 -993 185 -992
rect 268 -993 269 -992
rect 296 -993 297 -992
rect 394 -993 395 -992
rect 429 -993 430 -992
rect 646 -993 647 -992
rect 156 -995 157 -994
rect 163 -995 164 -994
rect 184 -995 185 -994
rect 205 -995 206 -994
rect 226 -995 227 -994
rect 289 -995 290 -994
rect 303 -995 304 -994
rect 436 -995 437 -994
rect 450 -995 451 -994
rect 478 -995 479 -994
rect 506 -995 507 -994
rect 583 -995 584 -994
rect 142 -997 143 -996
rect 156 -997 157 -996
rect 191 -997 192 -996
rect 282 -997 283 -996
rect 310 -997 311 -996
rect 345 -997 346 -996
rect 429 -997 430 -996
rect 485 -997 486 -996
rect 562 -997 563 -996
rect 583 -997 584 -996
rect 135 -999 136 -998
rect 142 -999 143 -998
rect 205 -999 206 -998
rect 275 -999 276 -998
rect 282 -999 283 -998
rect 366 -999 367 -998
rect 233 -1001 234 -1000
rect 275 -1001 276 -1000
rect 317 -1001 318 -1000
rect 457 -1001 458 -1000
rect 219 -1003 220 -1002
rect 233 -1003 234 -1002
rect 261 -1003 262 -1002
rect 289 -1003 290 -1002
rect 324 -1003 325 -1002
rect 338 -1003 339 -1002
rect 345 -1003 346 -1002
rect 408 -1003 409 -1002
rect 457 -1003 458 -1002
rect 604 -1003 605 -1002
rect 219 -1005 220 -1004
rect 247 -1005 248 -1004
rect 338 -1005 339 -1004
rect 359 -1005 360 -1004
rect 408 -1005 409 -1004
rect 415 -1005 416 -1004
rect 247 -1007 248 -1006
rect 303 -1007 304 -1006
rect 313 -1007 314 -1006
rect 415 -1007 416 -1006
rect 359 -1009 360 -1008
rect 387 -1009 388 -1008
rect 114 -1020 115 -1019
rect 173 -1020 174 -1019
rect 198 -1020 199 -1019
rect 348 -1020 349 -1019
rect 352 -1020 353 -1019
rect 460 -1020 461 -1019
rect 478 -1020 479 -1019
rect 506 -1020 507 -1019
rect 562 -1020 563 -1019
rect 576 -1020 577 -1019
rect 604 -1020 605 -1019
rect 611 -1020 612 -1019
rect 128 -1022 129 -1021
rect 163 -1022 164 -1021
rect 198 -1022 199 -1021
rect 219 -1022 220 -1021
rect 229 -1022 230 -1021
rect 247 -1022 248 -1021
rect 268 -1022 269 -1021
rect 366 -1022 367 -1021
rect 373 -1022 374 -1021
rect 429 -1022 430 -1021
rect 436 -1022 437 -1021
rect 450 -1022 451 -1021
rect 457 -1022 458 -1021
rect 464 -1022 465 -1021
rect 485 -1022 486 -1021
rect 492 -1022 493 -1021
rect 499 -1022 500 -1021
rect 527 -1022 528 -1021
rect 135 -1024 136 -1023
rect 149 -1024 150 -1023
rect 163 -1024 164 -1023
rect 177 -1024 178 -1023
rect 191 -1024 192 -1023
rect 247 -1024 248 -1023
rect 275 -1024 276 -1023
rect 317 -1024 318 -1023
rect 366 -1024 367 -1023
rect 380 -1024 381 -1023
rect 394 -1024 395 -1023
rect 474 -1024 475 -1023
rect 149 -1026 150 -1025
rect 156 -1026 157 -1025
rect 177 -1026 178 -1025
rect 219 -1026 220 -1025
rect 226 -1026 227 -1025
rect 268 -1026 269 -1025
rect 289 -1026 290 -1025
rect 359 -1026 360 -1025
rect 373 -1026 374 -1025
rect 415 -1026 416 -1025
rect 418 -1026 419 -1025
rect 422 -1026 423 -1025
rect 142 -1028 143 -1027
rect 156 -1028 157 -1027
rect 184 -1028 185 -1027
rect 191 -1028 192 -1027
rect 205 -1028 206 -1027
rect 306 -1028 307 -1027
rect 317 -1028 318 -1027
rect 338 -1028 339 -1027
rect 394 -1028 395 -1027
rect 401 -1028 402 -1027
rect 422 -1028 423 -1027
rect 443 -1028 444 -1027
rect 124 -1030 125 -1029
rect 142 -1030 143 -1029
rect 170 -1030 171 -1029
rect 205 -1030 206 -1029
rect 215 -1030 216 -1029
rect 233 -1030 234 -1029
rect 240 -1030 241 -1029
rect 243 -1030 244 -1029
rect 254 -1030 255 -1029
rect 289 -1030 290 -1029
rect 296 -1030 297 -1029
rect 310 -1030 311 -1029
rect 439 -1030 440 -1029
rect 443 -1030 444 -1029
rect 170 -1032 171 -1031
rect 282 -1032 283 -1031
rect 299 -1032 300 -1031
rect 303 -1032 304 -1031
rect 310 -1032 311 -1031
rect 324 -1032 325 -1031
rect 215 -1034 216 -1033
rect 254 -1034 255 -1033
rect 233 -1036 234 -1035
rect 264 -1036 265 -1035
rect 261 -1038 262 -1037
rect 264 -1038 265 -1037
rect 100 -1049 101 -1048
rect 107 -1049 108 -1048
rect 128 -1049 129 -1048
rect 194 -1049 195 -1048
rect 198 -1049 199 -1048
rect 212 -1049 213 -1048
rect 219 -1049 220 -1048
rect 226 -1049 227 -1048
rect 247 -1049 248 -1048
rect 303 -1049 304 -1048
rect 366 -1049 367 -1048
rect 380 -1049 381 -1048
rect 383 -1049 384 -1048
rect 387 -1049 388 -1048
rect 394 -1049 395 -1048
rect 404 -1049 405 -1048
rect 408 -1049 409 -1048
rect 411 -1049 412 -1048
rect 415 -1049 416 -1048
rect 429 -1049 430 -1048
rect 443 -1049 444 -1048
rect 453 -1049 454 -1048
rect 471 -1049 472 -1048
rect 485 -1049 486 -1048
rect 541 -1049 542 -1048
rect 548 -1049 549 -1048
rect 579 -1049 580 -1048
rect 583 -1049 584 -1048
rect 142 -1051 143 -1050
rect 173 -1051 174 -1050
rect 180 -1051 181 -1050
rect 233 -1051 234 -1050
rect 254 -1051 255 -1050
rect 275 -1051 276 -1050
rect 278 -1051 279 -1050
rect 296 -1051 297 -1050
rect 299 -1051 300 -1050
rect 310 -1051 311 -1050
rect 376 -1051 377 -1050
rect 422 -1051 423 -1050
rect 429 -1051 430 -1050
rect 436 -1051 437 -1050
rect 443 -1051 444 -1050
rect 478 -1051 479 -1050
rect 569 -1051 570 -1050
rect 583 -1051 584 -1050
rect 142 -1053 143 -1052
rect 156 -1053 157 -1052
rect 163 -1053 164 -1052
rect 184 -1053 185 -1052
rect 191 -1053 192 -1052
rect 198 -1053 199 -1052
rect 205 -1053 206 -1052
rect 233 -1053 234 -1052
rect 268 -1053 269 -1052
rect 282 -1053 283 -1052
rect 285 -1053 286 -1052
rect 317 -1053 318 -1052
rect 579 -1053 580 -1052
rect 590 -1053 591 -1052
rect 149 -1055 150 -1054
rect 163 -1055 164 -1054
rect 289 -1055 290 -1054
rect 296 -1055 297 -1054
rect 135 -1057 136 -1056
rect 149 -1057 150 -1056
rect 114 -1059 115 -1058
rect 135 -1059 136 -1058
rect 100 -1070 101 -1069
rect 107 -1070 108 -1069
rect 149 -1070 150 -1069
rect 159 -1070 160 -1069
rect 163 -1070 164 -1069
rect 170 -1070 171 -1069
rect 198 -1070 199 -1069
rect 205 -1070 206 -1069
rect 215 -1070 216 -1069
rect 233 -1070 234 -1069
rect 380 -1070 381 -1069
rect 394 -1070 395 -1069
rect 429 -1070 430 -1069
rect 439 -1070 440 -1069
rect 446 -1070 447 -1069
rect 457 -1070 458 -1069
rect 576 -1070 577 -1069
rect 583 -1070 584 -1069
rect 219 -1072 220 -1071
rect 226 -1072 227 -1071
<< metal2 >>
rect 114 -5 115 1
rect 121 -5 122 1
rect 128 -5 129 1
rect 149 -5 150 1
rect 156 -5 157 1
rect 166 -5 167 1
rect 177 -5 178 1
rect 198 -5 199 1
rect 236 -5 237 1
rect 247 -5 248 1
rect 296 -5 297 1
rect 313 -5 314 1
rect 317 -5 318 1
rect 373 -5 374 1
rect 131 -5 132 -1
rect 163 -5 164 -1
rect 191 -5 192 -1
rect 208 -5 209 -1
rect 331 -5 332 -1
rect 338 -5 339 -1
rect 348 -5 349 -1
rect 352 -5 353 -1
rect 135 -5 136 -3
rect 142 -5 143 -3
rect 72 -24 73 -14
rect 89 -24 90 -14
rect 100 -24 101 -14
rect 128 -24 129 -14
rect 131 -24 132 -14
rect 149 -24 150 -14
rect 156 -15 157 -13
rect 184 -15 185 -13
rect 187 -15 188 -13
rect 236 -15 237 -13
rect 247 -15 248 -13
rect 254 -24 255 -14
rect 296 -15 297 -13
rect 303 -24 304 -14
rect 331 -15 332 -13
rect 345 -24 346 -14
rect 352 -15 353 -13
rect 352 -24 353 -14
rect 352 -15 353 -13
rect 352 -24 353 -14
rect 373 -15 374 -13
rect 436 -24 437 -14
rect 485 -24 486 -14
rect 555 -24 556 -14
rect 79 -24 80 -16
rect 96 -24 97 -16
rect 107 -24 108 -16
rect 135 -17 136 -13
rect 142 -24 143 -16
rect 191 -17 192 -13
rect 201 -17 202 -13
rect 212 -24 213 -16
rect 215 -17 216 -13
rect 233 -24 234 -16
rect 296 -24 297 -16
rect 317 -17 318 -13
rect 394 -24 395 -16
rect 404 -24 405 -16
rect 422 -17 423 -13
rect 429 -24 430 -16
rect 117 -24 118 -18
rect 121 -19 122 -13
rect 135 -24 136 -18
rect 159 -24 160 -18
rect 170 -24 171 -18
rect 177 -19 178 -13
rect 184 -24 185 -18
rect 198 -24 199 -18
rect 219 -24 220 -18
rect 282 -24 283 -18
rect 313 -19 314 -13
rect 331 -24 332 -18
rect 156 -24 157 -20
rect 191 -24 192 -20
rect 229 -24 230 -20
rect 240 -24 241 -20
rect 173 -23 174 -13
rect 177 -24 178 -22
rect 51 -53 52 -33
rect 58 -53 59 -33
rect 65 -34 66 -32
rect 68 -38 69 -33
rect 79 -34 80 -32
rect 93 -53 94 -33
rect 96 -34 97 -32
rect 114 -53 115 -33
rect 149 -34 150 -32
rect 163 -53 164 -33
rect 166 -34 167 -32
rect 170 -34 171 -32
rect 184 -34 185 -32
rect 184 -53 185 -33
rect 184 -34 185 -32
rect 184 -53 185 -33
rect 191 -34 192 -32
rect 226 -34 227 -32
rect 233 -34 234 -32
rect 268 -53 269 -33
rect 275 -53 276 -33
rect 317 -53 318 -33
rect 345 -34 346 -32
rect 366 -53 367 -33
rect 387 -53 388 -33
rect 394 -34 395 -32
rect 415 -53 416 -33
rect 488 -34 489 -32
rect 555 -34 556 -32
rect 576 -53 577 -33
rect 65 -53 66 -35
rect 72 -36 73 -32
rect 86 -53 87 -35
rect 100 -36 101 -32
rect 107 -36 108 -32
rect 170 -53 171 -35
rect 212 -36 213 -32
rect 219 -53 220 -35
rect 233 -53 234 -35
rect 250 -36 251 -32
rect 254 -36 255 -32
rect 264 -36 265 -32
rect 285 -53 286 -35
rect 338 -53 339 -35
rect 352 -36 353 -32
rect 373 -53 374 -35
rect 380 -53 381 -35
rect 394 -53 395 -35
rect 429 -36 430 -32
rect 443 -53 444 -35
rect 72 -53 73 -37
rect 100 -53 101 -37
rect 117 -38 118 -32
rect 149 -53 150 -37
rect 205 -38 206 -32
rect 240 -38 241 -32
rect 247 -53 248 -37
rect 261 -38 262 -32
rect 261 -53 262 -37
rect 261 -38 262 -32
rect 261 -53 262 -37
rect 289 -53 290 -37
rect 313 -38 314 -32
rect 327 -38 328 -32
rect 345 -53 346 -37
rect 359 -53 360 -37
rect 404 -53 405 -37
rect 436 -38 437 -32
rect 450 -53 451 -37
rect 107 -53 108 -39
rect 222 -40 223 -32
rect 296 -40 297 -32
rect 296 -53 297 -39
rect 296 -40 297 -32
rect 296 -53 297 -39
rect 303 -40 304 -32
rect 324 -53 325 -39
rect 331 -40 332 -32
rect 352 -53 353 -39
rect 156 -53 157 -41
rect 198 -53 199 -41
rect 254 -53 255 -41
rect 303 -53 304 -41
rect 159 -44 160 -32
rect 177 -44 178 -32
rect 194 -53 195 -43
rect 205 -53 206 -43
rect 282 -44 283 -32
rect 331 -53 332 -43
rect 121 -46 122 -32
rect 159 -53 160 -45
rect 177 -53 178 -45
rect 226 -53 227 -45
rect 121 -53 122 -47
rect 135 -48 136 -32
rect 135 -53 136 -49
rect 142 -50 143 -32
rect 142 -53 143 -51
rect 215 -53 216 -51
rect 30 -92 31 -62
rect 152 -92 153 -62
rect 156 -92 157 -62
rect 170 -63 171 -61
rect 191 -63 192 -61
rect 268 -63 269 -61
rect 366 -63 367 -61
rect 408 -92 409 -62
rect 425 -92 426 -62
rect 464 -92 465 -62
rect 471 -92 472 -62
rect 527 -92 528 -62
rect 530 -92 531 -62
rect 590 -92 591 -62
rect 37 -92 38 -64
rect 51 -65 52 -61
rect 58 -92 59 -64
rect 82 -65 83 -61
rect 93 -65 94 -61
rect 226 -92 227 -64
rect 233 -65 234 -61
rect 268 -92 269 -64
rect 373 -65 374 -61
rect 429 -92 430 -64
rect 443 -65 444 -61
rect 492 -92 493 -64
rect 576 -65 577 -61
rect 576 -92 577 -64
rect 576 -65 577 -61
rect 576 -92 577 -64
rect 44 -92 45 -66
rect 135 -67 136 -61
rect 142 -67 143 -61
rect 212 -92 213 -66
rect 240 -67 241 -61
rect 247 -67 248 -61
rect 261 -67 262 -61
rect 285 -67 286 -61
rect 303 -92 304 -66
rect 373 -92 374 -66
rect 380 -92 381 -66
rect 387 -67 388 -61
rect 401 -67 402 -61
rect 478 -92 479 -66
rect 51 -92 52 -68
rect 121 -69 122 -61
rect 131 -69 132 -61
rect 170 -92 171 -68
rect 198 -69 199 -61
rect 198 -92 199 -68
rect 198 -69 199 -61
rect 198 -92 199 -68
rect 205 -69 206 -61
rect 233 -92 234 -68
rect 240 -92 241 -68
rect 254 -69 255 -61
rect 261 -92 262 -68
rect 289 -69 290 -61
rect 387 -92 388 -68
rect 394 -69 395 -61
rect 401 -92 402 -68
rect 415 -69 416 -61
rect 450 -69 451 -61
rect 450 -92 451 -68
rect 450 -69 451 -61
rect 450 -92 451 -68
rect 457 -69 458 -61
rect 457 -92 458 -68
rect 457 -69 458 -61
rect 457 -92 458 -68
rect 65 -71 66 -61
rect 96 -92 97 -70
rect 100 -71 101 -61
rect 177 -71 178 -61
rect 289 -92 290 -70
rect 359 -71 360 -61
rect 72 -73 73 -61
rect 79 -92 80 -72
rect 86 -73 87 -61
rect 100 -92 101 -72
rect 107 -73 108 -61
rect 107 -92 108 -72
rect 107 -73 108 -61
rect 107 -92 108 -72
rect 114 -73 115 -61
rect 114 -92 115 -72
rect 114 -73 115 -61
rect 114 -92 115 -72
rect 128 -73 129 -61
rect 177 -92 178 -72
rect 324 -73 325 -61
rect 415 -92 416 -72
rect 65 -92 66 -74
rect 86 -92 87 -74
rect 128 -92 129 -74
rect 247 -92 248 -74
rect 313 -75 314 -61
rect 324 -92 325 -74
rect 331 -75 332 -61
rect 394 -92 395 -74
rect 72 -92 73 -76
rect 215 -77 216 -61
rect 296 -77 297 -61
rect 331 -92 332 -76
rect 345 -77 346 -61
rect 359 -92 360 -76
rect 131 -92 132 -78
rect 135 -92 136 -78
rect 142 -92 143 -78
rect 184 -79 185 -61
rect 219 -79 220 -61
rect 296 -92 297 -78
rect 313 -92 314 -78
rect 436 -92 437 -78
rect 149 -81 150 -61
rect 191 -92 192 -80
rect 219 -92 220 -80
rect 243 -81 244 -61
rect 345 -92 346 -80
rect 369 -92 370 -80
rect 163 -83 164 -61
rect 205 -92 206 -82
rect 163 -92 164 -84
rect 229 -85 230 -61
rect 184 -92 185 -86
rect 275 -87 276 -61
rect 275 -92 276 -88
rect 338 -89 339 -61
rect 338 -92 339 -90
rect 352 -91 353 -61
rect 9 -143 10 -101
rect 37 -102 38 -100
rect 51 -102 52 -100
rect 121 -102 122 -100
rect 128 -143 129 -101
rect 257 -102 258 -100
rect 282 -102 283 -100
rect 527 -143 528 -101
rect 555 -143 556 -101
rect 576 -102 577 -100
rect 590 -102 591 -100
rect 618 -143 619 -101
rect 16 -143 17 -103
rect 58 -104 59 -100
rect 65 -143 66 -103
rect 100 -104 101 -100
rect 121 -143 122 -103
rect 156 -104 157 -100
rect 170 -104 171 -100
rect 313 -104 314 -100
rect 331 -104 332 -100
rect 457 -143 458 -103
rect 460 -104 461 -100
rect 590 -143 591 -103
rect 26 -143 27 -105
rect 68 -106 69 -100
rect 75 -143 76 -105
rect 156 -143 157 -105
rect 173 -143 174 -105
rect 191 -106 192 -100
rect 240 -106 241 -100
rect 562 -143 563 -105
rect 30 -108 31 -100
rect 93 -143 94 -107
rect 100 -143 101 -107
rect 107 -108 108 -100
rect 149 -108 150 -100
rect 240 -143 241 -107
rect 243 -108 244 -100
rect 268 -108 269 -100
rect 282 -143 283 -107
rect 289 -108 290 -100
rect 313 -143 314 -107
rect 359 -108 360 -100
rect 366 -108 367 -100
rect 569 -143 570 -107
rect 37 -143 38 -109
rect 79 -110 80 -100
rect 86 -110 87 -100
rect 149 -143 150 -109
rect 191 -143 192 -109
rect 198 -110 199 -100
rect 226 -110 227 -100
rect 268 -143 269 -109
rect 275 -110 276 -100
rect 289 -143 290 -109
rect 338 -110 339 -100
rect 359 -143 360 -109
rect 366 -143 367 -109
rect 450 -110 451 -100
rect 478 -110 479 -100
rect 576 -143 577 -109
rect 30 -143 31 -111
rect 275 -143 276 -111
rect 345 -112 346 -100
rect 352 -143 353 -111
rect 355 -112 356 -100
rect 604 -143 605 -111
rect 51 -143 52 -113
rect 96 -114 97 -100
rect 107 -143 108 -113
rect 114 -114 115 -100
rect 142 -114 143 -100
rect 338 -143 339 -113
rect 345 -143 346 -113
rect 401 -114 402 -100
rect 415 -114 416 -100
rect 534 -143 535 -113
rect 58 -143 59 -115
rect 86 -143 87 -115
rect 114 -143 115 -115
rect 124 -116 125 -100
rect 142 -143 143 -115
rect 163 -116 164 -100
rect 198 -143 199 -115
rect 212 -116 213 -100
rect 226 -143 227 -115
rect 446 -116 447 -100
rect 492 -116 493 -100
rect 611 -143 612 -115
rect 205 -118 206 -100
rect 212 -143 213 -117
rect 233 -118 234 -100
rect 401 -143 402 -117
rect 415 -143 416 -117
rect 492 -143 493 -117
rect 499 -143 500 -117
rect 506 -143 507 -117
rect 520 -143 521 -117
rect 523 -118 524 -100
rect 135 -120 136 -100
rect 233 -143 234 -119
rect 247 -120 248 -100
rect 548 -143 549 -119
rect 44 -122 45 -100
rect 135 -143 136 -121
rect 205 -143 206 -121
rect 219 -122 220 -100
rect 247 -143 248 -121
rect 303 -122 304 -100
rect 373 -122 374 -100
rect 513 -143 514 -121
rect 44 -143 45 -123
rect 72 -124 73 -100
rect 184 -124 185 -100
rect 303 -143 304 -123
rect 320 -124 321 -100
rect 373 -143 374 -123
rect 387 -124 388 -100
rect 450 -143 451 -123
rect 72 -143 73 -125
rect 331 -143 332 -125
rect 394 -126 395 -100
rect 597 -143 598 -125
rect 159 -128 160 -100
rect 184 -143 185 -127
rect 219 -143 220 -127
rect 222 -143 223 -127
rect 261 -128 262 -100
rect 320 -143 321 -127
rect 324 -128 325 -100
rect 387 -143 388 -127
rect 422 -143 423 -127
rect 464 -128 465 -100
rect 170 -143 171 -129
rect 261 -143 262 -129
rect 296 -130 297 -100
rect 394 -143 395 -129
rect 408 -130 409 -100
rect 464 -143 465 -129
rect 177 -132 178 -100
rect 296 -143 297 -131
rect 310 -143 311 -131
rect 324 -143 325 -131
rect 408 -143 409 -131
rect 471 -132 472 -100
rect 166 -143 167 -133
rect 177 -143 178 -133
rect 429 -134 430 -100
rect 478 -143 479 -133
rect 429 -143 430 -135
rect 474 -143 475 -135
rect 436 -138 437 -100
rect 485 -143 486 -137
rect 380 -140 381 -100
rect 436 -143 437 -139
rect 443 -140 444 -100
rect 541 -143 542 -139
rect 257 -143 258 -141
rect 380 -143 381 -141
rect 443 -143 444 -141
rect 586 -143 587 -141
rect 23 -204 24 -152
rect 191 -153 192 -151
rect 205 -153 206 -151
rect 257 -153 258 -151
rect 261 -153 262 -151
rect 569 -153 570 -151
rect 611 -153 612 -151
rect 660 -204 661 -152
rect 51 -155 52 -151
rect 180 -204 181 -154
rect 184 -155 185 -151
rect 418 -155 419 -151
rect 450 -155 451 -151
rect 450 -204 451 -154
rect 450 -155 451 -151
rect 450 -204 451 -154
rect 464 -155 465 -151
rect 639 -204 640 -154
rect 51 -204 52 -156
rect 128 -157 129 -151
rect 142 -157 143 -151
rect 184 -204 185 -156
rect 191 -204 192 -156
rect 292 -157 293 -151
rect 306 -204 307 -156
rect 597 -157 598 -151
rect 618 -157 619 -151
rect 625 -157 626 -151
rect 628 -157 629 -151
rect 646 -204 647 -156
rect 65 -159 66 -151
rect 93 -204 94 -158
rect 100 -159 101 -151
rect 128 -204 129 -158
rect 135 -159 136 -151
rect 142 -204 143 -158
rect 156 -159 157 -151
rect 163 -204 164 -158
rect 173 -159 174 -151
rect 198 -159 199 -151
rect 212 -159 213 -151
rect 310 -204 311 -158
rect 313 -159 314 -151
rect 590 -159 591 -151
rect 604 -159 605 -151
rect 625 -204 626 -158
rect 58 -161 59 -151
rect 65 -204 66 -160
rect 72 -161 73 -151
rect 138 -204 139 -160
rect 198 -204 199 -160
rect 247 -161 248 -151
rect 254 -204 255 -160
rect 296 -161 297 -151
rect 334 -204 335 -160
rect 667 -204 668 -160
rect 16 -163 17 -151
rect 58 -204 59 -162
rect 79 -163 80 -151
rect 156 -204 157 -162
rect 212 -204 213 -162
rect 261 -204 262 -162
rect 278 -163 279 -151
rect 534 -163 535 -151
rect 541 -163 542 -151
rect 569 -204 570 -162
rect 576 -163 577 -151
rect 590 -204 591 -162
rect 16 -204 17 -164
rect 44 -165 45 -151
rect 79 -204 80 -164
rect 107 -165 108 -151
rect 135 -204 136 -164
rect 299 -204 300 -164
rect 387 -165 388 -151
rect 674 -204 675 -164
rect 44 -204 45 -166
rect 282 -167 283 -151
rect 289 -204 290 -166
rect 324 -167 325 -151
rect 387 -204 388 -166
rect 618 -204 619 -166
rect 82 -169 83 -151
rect 96 -169 97 -151
rect 100 -204 101 -168
rect 401 -169 402 -151
rect 436 -169 437 -151
rect 464 -204 465 -168
rect 471 -169 472 -151
rect 597 -204 598 -168
rect 86 -171 87 -151
rect 149 -171 150 -151
rect 215 -204 216 -170
rect 394 -171 395 -151
rect 457 -171 458 -151
rect 534 -204 535 -170
rect 562 -171 563 -151
rect 604 -204 605 -170
rect 86 -204 87 -172
rect 114 -173 115 -151
rect 149 -204 150 -172
rect 527 -173 528 -151
rect 555 -173 556 -151
rect 562 -204 563 -172
rect 107 -204 108 -174
rect 121 -175 122 -151
rect 219 -175 220 -151
rect 338 -175 339 -151
rect 341 -204 342 -174
rect 471 -204 472 -174
rect 485 -175 486 -151
rect 632 -204 633 -174
rect 30 -177 31 -151
rect 219 -204 220 -176
rect 233 -177 234 -151
rect 233 -204 234 -176
rect 233 -177 234 -151
rect 233 -204 234 -176
rect 247 -204 248 -176
rect 586 -177 587 -151
rect 30 -204 31 -178
rect 240 -179 241 -151
rect 268 -179 269 -151
rect 394 -204 395 -178
rect 422 -179 423 -151
rect 457 -204 458 -178
rect 492 -179 493 -151
rect 611 -204 612 -178
rect 37 -181 38 -151
rect 121 -204 122 -180
rect 222 -181 223 -151
rect 422 -204 423 -180
rect 499 -204 500 -180
rect 513 -181 514 -151
rect 520 -181 521 -151
rect 541 -204 542 -180
rect 37 -204 38 -182
rect 96 -204 97 -182
rect 114 -204 115 -182
rect 226 -183 227 -151
rect 240 -204 241 -182
rect 278 -204 279 -182
rect 282 -204 283 -182
rect 369 -204 370 -182
rect 390 -204 391 -182
rect 653 -204 654 -182
rect 177 -185 178 -151
rect 226 -204 227 -184
rect 296 -204 297 -184
rect 380 -185 381 -151
rect 488 -204 489 -184
rect 513 -204 514 -184
rect 520 -204 521 -184
rect 583 -185 584 -151
rect 177 -204 178 -186
rect 208 -204 209 -186
rect 317 -187 318 -151
rect 555 -204 556 -186
rect 268 -204 269 -188
rect 317 -204 318 -188
rect 320 -189 321 -151
rect 436 -204 437 -188
rect 506 -189 507 -151
rect 527 -204 528 -188
rect 548 -189 549 -151
rect 583 -204 584 -188
rect 359 -191 360 -151
rect 492 -204 493 -190
rect 331 -193 332 -151
rect 359 -204 360 -192
rect 366 -193 367 -151
rect 401 -204 402 -192
rect 415 -193 416 -151
rect 548 -204 549 -192
rect 331 -204 332 -194
rect 576 -204 577 -194
rect 345 -197 346 -151
rect 415 -204 416 -196
rect 478 -197 479 -151
rect 506 -204 507 -196
rect 170 -199 171 -151
rect 345 -204 346 -198
rect 373 -199 374 -151
rect 380 -204 381 -198
rect 408 -199 409 -151
rect 478 -204 479 -198
rect 9 -201 10 -151
rect 170 -204 171 -200
rect 352 -201 353 -151
rect 373 -204 374 -200
rect 408 -204 409 -200
rect 429 -201 430 -151
rect 303 -203 304 -151
rect 352 -204 353 -202
rect 429 -204 430 -202
rect 443 -203 444 -151
rect 23 -214 24 -212
rect 212 -269 213 -213
rect 219 -214 220 -212
rect 219 -269 220 -213
rect 219 -214 220 -212
rect 219 -269 220 -213
rect 275 -214 276 -212
rect 534 -214 535 -212
rect 548 -214 549 -212
rect 688 -269 689 -213
rect 23 -269 24 -215
rect 96 -216 97 -212
rect 100 -269 101 -215
rect 107 -216 108 -212
rect 142 -216 143 -212
rect 142 -269 143 -215
rect 142 -216 143 -212
rect 142 -269 143 -215
rect 152 -269 153 -215
rect 243 -269 244 -215
rect 292 -269 293 -215
rect 534 -269 535 -215
rect 548 -269 549 -215
rect 597 -216 598 -212
rect 653 -216 654 -212
rect 695 -269 696 -215
rect 44 -218 45 -212
rect 93 -269 94 -217
rect 103 -269 104 -217
rect 233 -218 234 -212
rect 296 -269 297 -217
rect 429 -218 430 -212
rect 446 -218 447 -212
rect 597 -269 598 -217
rect 660 -218 661 -212
rect 716 -269 717 -217
rect 44 -269 45 -219
rect 54 -269 55 -219
rect 58 -220 59 -212
rect 58 -269 59 -219
rect 58 -220 59 -212
rect 58 -269 59 -219
rect 65 -220 66 -212
rect 75 -220 76 -212
rect 86 -220 87 -212
rect 135 -220 136 -212
rect 156 -220 157 -212
rect 278 -220 279 -212
rect 303 -269 304 -219
rect 352 -220 353 -212
rect 369 -220 370 -212
rect 618 -220 619 -212
rect 51 -222 52 -212
rect 72 -269 73 -221
rect 86 -269 87 -221
rect 278 -269 279 -221
rect 313 -269 314 -221
rect 569 -222 570 -212
rect 583 -222 584 -212
rect 618 -269 619 -221
rect 51 -269 52 -223
rect 149 -224 150 -212
rect 163 -224 164 -212
rect 163 -269 164 -223
rect 163 -224 164 -212
rect 163 -269 164 -223
rect 170 -224 171 -212
rect 324 -269 325 -223
rect 331 -224 332 -212
rect 639 -224 640 -212
rect 37 -226 38 -212
rect 331 -269 332 -225
rect 338 -269 339 -225
rect 359 -226 360 -212
rect 369 -269 370 -225
rect 569 -269 570 -225
rect 590 -226 591 -212
rect 653 -269 654 -225
rect 9 -269 10 -227
rect 37 -269 38 -227
rect 65 -269 66 -227
rect 82 -269 83 -227
rect 128 -228 129 -212
rect 156 -269 157 -227
rect 177 -228 178 -212
rect 310 -228 311 -212
rect 341 -228 342 -212
rect 492 -228 493 -212
rect 499 -228 500 -212
rect 590 -269 591 -227
rect 611 -228 612 -212
rect 660 -269 661 -227
rect 16 -230 17 -212
rect 177 -269 178 -229
rect 191 -230 192 -212
rect 205 -269 206 -229
rect 233 -269 234 -229
rect 240 -230 241 -212
rect 254 -230 255 -212
rect 352 -269 353 -229
rect 387 -230 388 -212
rect 632 -230 633 -212
rect 16 -269 17 -231
rect 117 -269 118 -231
rect 128 -269 129 -231
rect 184 -232 185 -212
rect 191 -269 192 -231
rect 226 -232 227 -212
rect 254 -269 255 -231
rect 268 -232 269 -212
rect 299 -232 300 -212
rect 639 -269 640 -231
rect 30 -234 31 -212
rect 310 -269 311 -233
rect 345 -234 346 -212
rect 359 -269 360 -233
rect 422 -234 423 -212
rect 723 -269 724 -233
rect 33 -269 34 -235
rect 226 -269 227 -235
rect 247 -236 248 -212
rect 345 -269 346 -235
rect 408 -236 409 -212
rect 422 -269 423 -235
rect 457 -236 458 -212
rect 485 -269 486 -235
rect 488 -236 489 -212
rect 604 -236 605 -212
rect 79 -238 80 -212
rect 170 -269 171 -237
rect 198 -238 199 -212
rect 201 -246 202 -237
rect 247 -269 248 -237
rect 681 -269 682 -237
rect 2 -269 3 -239
rect 79 -269 80 -239
rect 107 -269 108 -239
rect 387 -269 388 -239
rect 464 -240 465 -212
rect 492 -269 493 -239
rect 513 -240 514 -212
rect 702 -269 703 -239
rect 121 -242 122 -212
rect 184 -269 185 -241
rect 198 -269 199 -241
rect 289 -242 290 -212
rect 299 -269 300 -241
rect 429 -269 430 -241
rect 471 -242 472 -212
rect 499 -269 500 -241
rect 513 -269 514 -241
rect 674 -242 675 -212
rect 121 -269 122 -243
rect 264 -269 265 -243
rect 268 -269 269 -243
rect 282 -244 283 -212
rect 327 -244 328 -212
rect 457 -269 458 -243
rect 471 -269 472 -243
rect 478 -244 479 -212
rect 527 -244 528 -212
rect 583 -269 584 -243
rect 135 -269 136 -245
rect 180 -246 181 -212
rect 289 -269 290 -245
rect 366 -246 367 -212
rect 527 -269 528 -245
rect 555 -246 556 -212
rect 604 -269 605 -245
rect 250 -269 251 -247
rect 555 -269 556 -247
rect 562 -248 563 -212
rect 632 -269 633 -247
rect 261 -250 262 -212
rect 282 -269 283 -249
rect 380 -250 381 -212
rect 408 -269 409 -249
rect 436 -250 437 -212
rect 478 -269 479 -249
rect 506 -250 507 -212
rect 562 -269 563 -249
rect 576 -250 577 -212
rect 611 -269 612 -249
rect 380 -269 381 -251
rect 646 -252 647 -212
rect 383 -269 384 -253
rect 674 -269 675 -253
rect 394 -256 395 -212
rect 436 -269 437 -255
rect 506 -269 507 -255
rect 667 -256 668 -212
rect 394 -269 395 -257
rect 401 -258 402 -212
rect 541 -258 542 -212
rect 576 -269 577 -257
rect 625 -258 626 -212
rect 667 -269 668 -257
rect 373 -260 374 -212
rect 401 -269 402 -259
rect 415 -260 416 -212
rect 541 -269 542 -259
rect 646 -269 647 -259
rect 712 -269 713 -259
rect 30 -269 31 -261
rect 373 -269 374 -261
rect 443 -262 444 -212
rect 625 -269 626 -261
rect 317 -264 318 -212
rect 415 -269 416 -263
rect 443 -269 444 -263
rect 450 -264 451 -212
rect 114 -266 115 -212
rect 317 -269 318 -265
rect 450 -269 451 -265
rect 520 -266 521 -212
rect 520 -269 521 -267
rect 730 -269 731 -267
rect 23 -279 24 -277
rect 54 -279 55 -277
rect 58 -279 59 -277
rect 110 -279 111 -277
rect 128 -279 129 -277
rect 278 -279 279 -277
rect 289 -336 290 -278
rect 352 -279 353 -277
rect 362 -336 363 -278
rect 541 -279 542 -277
rect 569 -279 570 -277
rect 730 -336 731 -278
rect 26 -336 27 -280
rect 226 -281 227 -277
rect 240 -281 241 -277
rect 527 -281 528 -277
rect 534 -281 535 -277
rect 569 -336 570 -280
rect 576 -281 577 -277
rect 576 -336 577 -280
rect 576 -281 577 -277
rect 576 -336 577 -280
rect 604 -281 605 -277
rect 604 -336 605 -280
rect 604 -281 605 -277
rect 604 -336 605 -280
rect 716 -281 717 -277
rect 737 -336 738 -280
rect 2 -283 3 -277
rect 226 -336 227 -282
rect 247 -283 248 -277
rect 303 -283 304 -277
rect 310 -283 311 -277
rect 338 -283 339 -277
rect 345 -283 346 -277
rect 352 -336 353 -282
rect 373 -283 374 -277
rect 373 -336 374 -282
rect 373 -283 374 -277
rect 373 -336 374 -282
rect 380 -283 381 -277
rect 639 -283 640 -277
rect 30 -336 31 -284
rect 72 -285 73 -277
rect 82 -285 83 -277
rect 667 -285 668 -277
rect 16 -287 17 -277
rect 72 -336 73 -286
rect 86 -287 87 -277
rect 303 -336 304 -286
rect 310 -336 311 -286
rect 313 -287 314 -277
rect 338 -336 339 -286
rect 415 -287 416 -277
rect 422 -287 423 -277
rect 464 -336 465 -286
rect 467 -287 468 -277
rect 548 -287 549 -277
rect 639 -336 640 -286
rect 653 -287 654 -277
rect 667 -336 668 -286
rect 681 -287 682 -277
rect 16 -336 17 -288
rect 205 -289 206 -277
rect 212 -289 213 -277
rect 250 -289 251 -277
rect 292 -289 293 -277
rect 716 -336 717 -288
rect 33 -291 34 -277
rect 534 -336 535 -290
rect 541 -336 542 -290
rect 590 -291 591 -277
rect 653 -336 654 -290
rect 674 -291 675 -277
rect 37 -293 38 -277
rect 79 -336 80 -292
rect 100 -336 101 -292
rect 170 -293 171 -277
rect 198 -293 199 -277
rect 348 -336 349 -292
rect 380 -336 381 -292
rect 401 -293 402 -277
rect 422 -336 423 -292
rect 506 -293 507 -277
rect 548 -336 549 -292
rect 562 -293 563 -277
rect 590 -336 591 -292
rect 611 -293 612 -277
rect 44 -295 45 -277
rect 527 -336 528 -294
rect 555 -295 556 -277
rect 681 -336 682 -294
rect 47 -336 48 -296
rect 436 -297 437 -277
rect 478 -297 479 -277
rect 478 -336 479 -296
rect 478 -297 479 -277
rect 478 -336 479 -296
rect 485 -297 486 -277
rect 485 -336 486 -296
rect 485 -297 486 -277
rect 485 -336 486 -296
rect 492 -297 493 -277
rect 492 -336 493 -296
rect 492 -297 493 -277
rect 492 -336 493 -296
rect 499 -297 500 -277
rect 506 -336 507 -296
rect 555 -336 556 -296
rect 597 -297 598 -277
rect 51 -299 52 -277
rect 86 -336 87 -298
rect 107 -299 108 -277
rect 205 -336 206 -298
rect 212 -336 213 -298
rect 383 -299 384 -277
rect 394 -299 395 -277
rect 415 -336 416 -298
rect 432 -336 433 -298
rect 520 -299 521 -277
rect 562 -336 563 -298
rect 583 -299 584 -277
rect 597 -336 598 -298
rect 625 -299 626 -277
rect 54 -336 55 -300
rect 114 -301 115 -277
rect 121 -301 122 -277
rect 128 -336 129 -300
rect 135 -301 136 -277
rect 149 -336 150 -300
rect 156 -301 157 -277
rect 240 -336 241 -300
rect 257 -336 258 -300
rect 611 -336 612 -300
rect 625 -336 626 -300
rect 632 -301 633 -277
rect 58 -336 59 -302
rect 296 -303 297 -277
rect 345 -336 346 -302
rect 702 -303 703 -277
rect 65 -305 66 -277
rect 187 -336 188 -304
rect 191 -305 192 -277
rect 198 -336 199 -304
rect 219 -305 220 -277
rect 247 -336 248 -304
rect 261 -305 262 -277
rect 674 -336 675 -304
rect 65 -336 66 -306
rect 268 -307 269 -277
rect 299 -307 300 -277
rect 702 -336 703 -306
rect 93 -309 94 -277
rect 268 -336 269 -308
rect 299 -336 300 -308
rect 513 -309 514 -277
rect 583 -336 584 -308
rect 618 -309 619 -277
rect 632 -336 633 -308
rect 646 -309 647 -277
rect 110 -336 111 -310
rect 114 -336 115 -310
rect 121 -336 122 -310
rect 369 -311 370 -277
rect 394 -336 395 -310
rect 408 -311 409 -277
rect 436 -336 437 -310
rect 709 -311 710 -277
rect 135 -336 136 -312
rect 184 -313 185 -277
rect 191 -336 192 -312
rect 282 -313 283 -277
rect 401 -336 402 -312
rect 723 -313 724 -277
rect 37 -336 38 -314
rect 184 -336 185 -314
rect 275 -315 276 -277
rect 618 -336 619 -314
rect 646 -336 647 -314
rect 660 -315 661 -277
rect 695 -315 696 -277
rect 723 -336 724 -314
rect 44 -336 45 -316
rect 695 -336 696 -316
rect 93 -336 94 -318
rect 282 -336 283 -318
rect 443 -319 444 -277
rect 499 -336 500 -318
rect 660 -336 661 -318
rect 688 -319 689 -277
rect 142 -321 143 -277
rect 170 -336 171 -320
rect 177 -321 178 -277
rect 261 -336 262 -320
rect 275 -336 276 -320
rect 408 -336 409 -320
rect 457 -321 458 -277
rect 520 -336 521 -320
rect 142 -336 143 -322
rect 264 -323 265 -277
rect 324 -323 325 -277
rect 457 -336 458 -322
rect 471 -323 472 -277
rect 513 -336 514 -322
rect 156 -336 157 -324
rect 233 -325 234 -277
rect 324 -336 325 -324
rect 387 -325 388 -277
rect 450 -325 451 -277
rect 471 -336 472 -324
rect 51 -336 52 -326
rect 233 -336 234 -326
rect 278 -336 279 -326
rect 387 -336 388 -326
rect 429 -327 430 -277
rect 450 -336 451 -326
rect 163 -329 164 -277
rect 219 -336 220 -328
rect 327 -336 328 -328
rect 688 -336 689 -328
rect 177 -336 178 -330
rect 254 -331 255 -277
rect 331 -331 332 -277
rect 443 -336 444 -330
rect 317 -333 318 -277
rect 331 -336 332 -332
rect 429 -336 430 -332
rect 709 -336 710 -332
rect 317 -336 318 -334
rect 359 -335 360 -277
rect 5 -415 6 -345
rect 359 -415 360 -345
rect 369 -346 370 -344
rect 478 -346 479 -344
rect 555 -346 556 -344
rect 758 -415 759 -345
rect 23 -415 24 -347
rect 366 -348 367 -344
rect 373 -348 374 -344
rect 373 -415 374 -347
rect 373 -348 374 -344
rect 373 -415 374 -347
rect 376 -415 377 -347
rect 800 -415 801 -347
rect 26 -350 27 -344
rect 450 -350 451 -344
rect 474 -415 475 -349
rect 765 -415 766 -349
rect 30 -352 31 -344
rect 184 -415 185 -351
rect 187 -352 188 -344
rect 247 -352 248 -344
rect 261 -352 262 -344
rect 261 -415 262 -351
rect 261 -352 262 -344
rect 261 -415 262 -351
rect 268 -352 269 -344
rect 278 -352 279 -344
rect 282 -352 283 -344
rect 569 -352 570 -344
rect 667 -352 668 -344
rect 744 -415 745 -351
rect 30 -415 31 -353
rect 156 -354 157 -344
rect 219 -354 220 -344
rect 254 -354 255 -344
rect 268 -415 269 -353
rect 457 -354 458 -344
rect 513 -354 514 -344
rect 569 -415 570 -353
rect 583 -354 584 -344
rect 667 -415 668 -353
rect 674 -354 675 -344
rect 751 -415 752 -353
rect 2 -415 3 -355
rect 583 -415 584 -355
rect 688 -356 689 -344
rect 772 -415 773 -355
rect 44 -415 45 -357
rect 397 -415 398 -357
rect 408 -358 409 -344
rect 457 -415 458 -357
rect 464 -358 465 -344
rect 513 -415 514 -357
rect 527 -358 528 -344
rect 674 -415 675 -357
rect 695 -358 696 -344
rect 779 -415 780 -357
rect 47 -360 48 -344
rect 296 -360 297 -344
rect 324 -415 325 -359
rect 345 -360 346 -344
rect 352 -360 353 -344
rect 366 -415 367 -359
rect 408 -415 409 -359
rect 415 -360 416 -344
rect 432 -415 433 -359
rect 723 -360 724 -344
rect 730 -360 731 -344
rect 807 -415 808 -359
rect 51 -415 52 -361
rect 191 -362 192 -344
rect 219 -415 220 -361
rect 443 -362 444 -344
rect 485 -362 486 -344
rect 527 -415 528 -361
rect 558 -415 559 -361
rect 814 -415 815 -361
rect 54 -364 55 -344
rect 404 -415 405 -363
rect 415 -415 416 -363
rect 737 -364 738 -344
rect 61 -366 62 -344
rect 229 -366 230 -344
rect 233 -366 234 -344
rect 418 -415 419 -365
rect 422 -366 423 -344
rect 443 -415 444 -365
rect 471 -366 472 -344
rect 485 -415 486 -365
rect 562 -366 563 -344
rect 562 -415 563 -365
rect 562 -366 563 -344
rect 562 -415 563 -365
rect 618 -366 619 -344
rect 688 -415 689 -365
rect 709 -366 710 -344
rect 786 -415 787 -365
rect 72 -368 73 -344
rect 233 -415 234 -367
rect 247 -415 248 -367
rect 338 -368 339 -344
rect 345 -415 346 -367
rect 702 -368 703 -344
rect 716 -368 717 -344
rect 793 -415 794 -367
rect 72 -415 73 -369
rect 86 -370 87 -344
rect 93 -370 94 -344
rect 275 -415 276 -369
rect 282 -415 283 -369
rect 331 -370 332 -344
rect 338 -415 339 -369
rect 450 -415 451 -369
rect 625 -370 626 -344
rect 695 -415 696 -369
rect 37 -372 38 -344
rect 331 -415 332 -371
rect 348 -372 349 -344
rect 723 -415 724 -371
rect 79 -374 80 -344
rect 191 -415 192 -373
rect 226 -374 227 -344
rect 352 -415 353 -373
rect 387 -374 388 -344
rect 422 -415 423 -373
rect 429 -374 430 -344
rect 618 -415 619 -373
rect 639 -374 640 -344
rect 702 -415 703 -373
rect 79 -415 80 -375
rect 177 -376 178 -344
rect 226 -415 227 -375
rect 317 -376 318 -344
rect 348 -415 349 -375
rect 737 -415 738 -375
rect 86 -415 87 -377
rect 135 -378 136 -344
rect 149 -378 150 -344
rect 149 -415 150 -377
rect 149 -378 150 -344
rect 149 -415 150 -377
rect 285 -378 286 -344
rect 523 -415 524 -377
rect 541 -378 542 -344
rect 639 -415 640 -377
rect 646 -378 647 -344
rect 709 -415 710 -377
rect 93 -415 94 -379
rect 341 -415 342 -379
rect 436 -380 437 -344
rect 478 -415 479 -379
rect 492 -380 493 -344
rect 541 -415 542 -379
rect 576 -380 577 -344
rect 625 -415 626 -379
rect 646 -415 647 -379
rect 660 -380 661 -344
rect 681 -380 682 -344
rect 730 -415 731 -379
rect 100 -382 101 -344
rect 135 -415 136 -381
rect 289 -382 290 -344
rect 387 -415 388 -381
rect 394 -382 395 -344
rect 436 -415 437 -381
rect 492 -415 493 -381
rect 499 -382 500 -344
rect 520 -382 521 -344
rect 576 -415 577 -381
rect 590 -382 591 -344
rect 660 -415 661 -381
rect 100 -415 101 -383
rect 205 -384 206 -344
rect 292 -415 293 -383
rect 464 -415 465 -383
rect 590 -415 591 -383
rect 597 -384 598 -344
rect 611 -384 612 -344
rect 681 -415 682 -383
rect 107 -415 108 -385
rect 632 -386 633 -344
rect 653 -386 654 -344
rect 716 -415 717 -385
rect 110 -388 111 -344
rect 254 -415 255 -387
rect 296 -415 297 -387
rect 303 -388 304 -344
rect 310 -388 311 -344
rect 317 -415 318 -387
rect 534 -388 535 -344
rect 597 -415 598 -387
rect 604 -388 605 -344
rect 611 -415 612 -387
rect 110 -415 111 -389
rect 499 -415 500 -389
rect 548 -390 549 -344
rect 653 -415 654 -389
rect 121 -392 122 -344
rect 205 -415 206 -391
rect 222 -415 223 -391
rect 310 -415 311 -391
rect 383 -415 384 -391
rect 604 -415 605 -391
rect 124 -415 125 -393
rect 156 -415 157 -393
rect 163 -394 164 -344
rect 289 -415 290 -393
rect 299 -394 300 -344
rect 632 -415 633 -393
rect 114 -396 115 -344
rect 163 -415 164 -395
rect 303 -415 304 -395
rect 334 -415 335 -395
rect 401 -396 402 -344
rect 534 -415 535 -395
rect 37 -415 38 -397
rect 401 -415 402 -397
rect 506 -398 507 -344
rect 548 -415 549 -397
rect 114 -415 115 -399
rect 240 -400 241 -344
rect 128 -402 129 -344
rect 177 -415 178 -401
rect 240 -415 241 -401
rect 380 -402 381 -344
rect 128 -415 129 -403
rect 142 -404 143 -344
rect 212 -404 213 -344
rect 380 -415 381 -403
rect 16 -406 17 -344
rect 212 -415 213 -405
rect 16 -415 17 -407
rect 198 -408 199 -344
rect 142 -415 143 -409
rect 170 -410 171 -344
rect 198 -415 199 -409
rect 394 -415 395 -409
rect 65 -412 66 -344
rect 170 -415 171 -411
rect 58 -414 59 -344
rect 65 -415 66 -413
rect 9 -425 10 -423
rect 51 -425 52 -423
rect 58 -425 59 -423
rect 68 -467 69 -424
rect 72 -425 73 -423
rect 138 -508 139 -424
rect 170 -425 171 -423
rect 219 -425 220 -423
rect 264 -508 265 -424
rect 751 -425 752 -423
rect 9 -508 10 -426
rect 44 -427 45 -423
rect 47 -508 48 -426
rect 667 -427 668 -423
rect 702 -427 703 -423
rect 705 -427 706 -423
rect 51 -508 52 -428
rect 100 -429 101 -423
rect 107 -429 108 -423
rect 674 -429 675 -423
rect 702 -508 703 -428
rect 744 -429 745 -423
rect 58 -508 59 -430
rect 758 -431 759 -423
rect 61 -508 62 -432
rect 268 -433 269 -423
rect 275 -433 276 -423
rect 373 -508 374 -432
rect 380 -433 381 -423
rect 660 -433 661 -423
rect 730 -433 731 -423
rect 744 -508 745 -432
rect 72 -508 73 -434
rect 198 -435 199 -423
rect 205 -435 206 -423
rect 289 -508 290 -434
rect 334 -435 335 -423
rect 597 -435 598 -423
rect 611 -435 612 -423
rect 674 -508 675 -434
rect 716 -435 717 -423
rect 730 -508 731 -434
rect 79 -437 80 -423
rect 275 -508 276 -436
rect 338 -437 339 -423
rect 653 -437 654 -423
rect 79 -508 80 -438
rect 296 -439 297 -423
rect 348 -439 349 -423
rect 723 -439 724 -423
rect 86 -441 87 -423
rect 121 -508 122 -440
rect 163 -441 164 -423
rect 205 -508 206 -440
rect 233 -441 234 -423
rect 338 -508 339 -440
rect 366 -441 367 -423
rect 383 -441 384 -423
rect 394 -441 395 -423
rect 639 -441 640 -423
rect 646 -441 647 -423
rect 758 -508 759 -440
rect 44 -508 45 -442
rect 233 -508 234 -442
rect 254 -443 255 -423
rect 296 -508 297 -442
rect 387 -443 388 -423
rect 394 -508 395 -442
rect 401 -508 402 -442
rect 632 -443 633 -423
rect 709 -443 710 -423
rect 723 -508 724 -442
rect 86 -508 87 -444
rect 359 -445 360 -423
rect 404 -445 405 -423
rect 793 -445 794 -423
rect 93 -447 94 -423
rect 163 -508 164 -446
rect 170 -508 171 -446
rect 222 -447 223 -423
rect 226 -447 227 -423
rect 366 -508 367 -446
rect 436 -447 437 -423
rect 436 -508 437 -446
rect 436 -447 437 -423
rect 436 -508 437 -446
rect 443 -447 444 -423
rect 611 -508 612 -446
rect 618 -447 619 -423
rect 639 -508 640 -446
rect 695 -447 696 -423
rect 709 -508 710 -446
rect 793 -508 794 -446
rect 807 -447 808 -423
rect 93 -508 94 -448
rect 345 -449 346 -423
rect 352 -449 353 -423
rect 359 -508 360 -448
rect 450 -449 451 -423
rect 450 -508 451 -448
rect 450 -449 451 -423
rect 450 -508 451 -448
rect 474 -449 475 -423
rect 772 -449 773 -423
rect 100 -508 101 -450
rect 404 -508 405 -450
rect 474 -508 475 -450
rect 660 -508 661 -450
rect 681 -451 682 -423
rect 695 -508 696 -450
rect 772 -508 773 -450
rect 786 -451 787 -423
rect 107 -508 108 -452
rect 128 -453 129 -423
rect 198 -508 199 -452
rect 317 -453 318 -423
rect 324 -453 325 -423
rect 345 -508 346 -452
rect 355 -508 356 -452
rect 618 -508 619 -452
rect 625 -453 626 -423
rect 646 -508 647 -452
rect 786 -508 787 -452
rect 800 -453 801 -423
rect 30 -455 31 -423
rect 128 -508 129 -454
rect 191 -455 192 -423
rect 324 -508 325 -454
rect 506 -455 507 -423
rect 597 -508 598 -454
rect 604 -455 605 -423
rect 632 -508 633 -454
rect 800 -508 801 -454
rect 814 -455 815 -423
rect 30 -508 31 -456
rect 432 -457 433 -423
rect 520 -457 521 -423
rect 737 -457 738 -423
rect 37 -459 38 -423
rect 506 -508 507 -458
rect 523 -459 524 -423
rect 765 -459 766 -423
rect 37 -508 38 -460
rect 149 -461 150 -423
rect 212 -461 213 -423
rect 254 -508 255 -460
rect 261 -461 262 -423
rect 268 -508 269 -460
rect 303 -461 304 -423
rect 317 -508 318 -460
rect 418 -461 419 -423
rect 520 -508 521 -460
rect 541 -461 542 -423
rect 544 -467 545 -460
rect 558 -508 559 -460
rect 751 -508 752 -460
rect 765 -508 766 -460
rect 779 -461 780 -423
rect 110 -463 111 -423
rect 191 -508 192 -462
rect 222 -508 223 -462
rect 779 -508 780 -462
rect 135 -465 136 -423
rect 212 -508 213 -464
rect 247 -465 248 -423
rect 443 -508 444 -464
rect 541 -508 542 -464
rect 590 -465 591 -423
rect 681 -508 682 -464
rect 688 -465 689 -423
rect 737 -508 738 -464
rect 149 -508 150 -466
rect 383 -508 384 -466
rect 562 -467 563 -423
rect 653 -508 654 -466
rect 705 -508 706 -466
rect 716 -508 717 -466
rect 247 -508 248 -468
rect 282 -469 283 -423
rect 303 -508 304 -468
rect 464 -469 465 -423
rect 492 -469 493 -423
rect 562 -508 563 -468
rect 569 -469 570 -423
rect 590 -508 591 -468
rect 282 -508 283 -470
rect 310 -471 311 -423
rect 380 -508 381 -470
rect 688 -508 689 -470
rect 16 -473 17 -423
rect 310 -508 311 -472
rect 422 -473 423 -423
rect 464 -508 465 -472
rect 492 -508 493 -472
rect 667 -508 668 -472
rect 16 -508 17 -474
rect 124 -475 125 -423
rect 422 -508 423 -474
rect 478 -475 479 -423
rect 548 -475 549 -423
rect 569 -508 570 -474
rect 576 -475 577 -423
rect 604 -508 605 -474
rect 415 -477 416 -423
rect 478 -508 479 -476
rect 527 -477 528 -423
rect 548 -508 549 -476
rect 555 -477 556 -423
rect 576 -508 577 -476
rect 408 -479 409 -423
rect 415 -508 416 -478
rect 485 -479 486 -423
rect 527 -508 528 -478
rect 485 -508 486 -480
rect 534 -481 535 -423
rect 457 -483 458 -423
rect 534 -508 535 -482
rect 457 -508 458 -484
rect 513 -485 514 -423
rect 499 -487 500 -423
rect 513 -508 514 -486
rect 331 -489 332 -423
rect 499 -508 500 -488
rect 156 -491 157 -423
rect 331 -508 332 -490
rect 156 -508 157 -492
rect 184 -493 185 -423
rect 142 -495 143 -423
rect 184 -508 185 -494
rect 142 -508 143 -496
rect 177 -497 178 -423
rect 23 -499 24 -423
rect 177 -508 178 -498
rect 23 -508 24 -500
rect 240 -501 241 -423
rect 65 -503 66 -423
rect 240 -508 241 -502
rect 65 -508 66 -504
rect 114 -505 115 -423
rect 114 -508 115 -506
rect 471 -507 472 -423
rect 9 -518 10 -516
rect 103 -518 104 -516
rect 163 -518 164 -516
rect 432 -518 433 -516
rect 467 -577 468 -517
rect 772 -518 773 -516
rect 793 -518 794 -516
rect 807 -577 808 -517
rect 9 -577 10 -519
rect 100 -520 101 -516
rect 163 -577 164 -519
rect 177 -520 178 -516
rect 184 -520 185 -516
rect 219 -520 220 -516
rect 222 -520 223 -516
rect 534 -520 535 -516
rect 555 -577 556 -519
rect 576 -520 577 -516
rect 583 -520 584 -516
rect 821 -577 822 -519
rect 16 -522 17 -516
rect 264 -522 265 -516
rect 313 -522 314 -516
rect 359 -522 360 -516
rect 380 -577 381 -521
rect 558 -522 559 -516
rect 618 -522 619 -516
rect 621 -528 622 -521
rect 681 -522 682 -516
rect 681 -577 682 -521
rect 681 -522 682 -516
rect 681 -577 682 -521
rect 709 -522 710 -516
rect 709 -577 710 -521
rect 709 -522 710 -516
rect 709 -577 710 -521
rect 779 -522 780 -516
rect 793 -577 794 -521
rect 800 -522 801 -516
rect 814 -577 815 -521
rect 16 -577 17 -523
rect 450 -524 451 -516
rect 471 -577 472 -523
rect 492 -524 493 -516
rect 495 -524 496 -516
rect 702 -524 703 -516
rect 758 -524 759 -516
rect 779 -577 780 -523
rect 786 -524 787 -516
rect 800 -577 801 -523
rect 44 -577 45 -525
rect 110 -577 111 -525
rect 135 -526 136 -516
rect 450 -577 451 -525
rect 457 -526 458 -516
rect 492 -577 493 -525
rect 520 -526 521 -516
rect 534 -577 535 -525
rect 541 -526 542 -516
rect 583 -577 584 -525
rect 618 -577 619 -525
rect 653 -526 654 -516
rect 744 -526 745 -516
rect 758 -577 759 -525
rect 765 -526 766 -516
rect 786 -577 787 -525
rect 47 -528 48 -516
rect 331 -528 332 -516
rect 383 -528 384 -516
rect 548 -528 549 -516
rect 653 -577 654 -527
rect 54 -577 55 -529
rect 191 -530 192 -516
rect 226 -530 227 -516
rect 275 -530 276 -516
rect 303 -577 304 -529
rect 313 -577 314 -529
rect 317 -530 318 -516
rect 331 -577 332 -529
rect 383 -577 384 -529
rect 562 -530 563 -516
rect 625 -530 626 -516
rect 744 -577 745 -529
rect 58 -577 59 -531
rect 93 -532 94 -516
rect 131 -577 132 -531
rect 191 -577 192 -531
rect 212 -532 213 -516
rect 226 -577 227 -531
rect 233 -532 234 -516
rect 359 -577 360 -531
rect 387 -532 388 -516
rect 772 -577 773 -531
rect 61 -534 62 -516
rect 100 -577 101 -533
rect 121 -534 122 -516
rect 233 -577 234 -533
rect 240 -534 241 -516
rect 387 -577 388 -533
rect 390 -534 391 -516
rect 513 -534 514 -516
rect 520 -577 521 -533
rect 527 -534 528 -516
rect 541 -577 542 -533
rect 590 -534 591 -516
rect 625 -577 626 -533
rect 639 -534 640 -516
rect 79 -536 80 -516
rect 219 -577 220 -535
rect 240 -577 241 -535
rect 373 -536 374 -516
rect 394 -536 395 -516
rect 408 -577 409 -535
rect 429 -536 430 -516
rect 730 -536 731 -516
rect 79 -577 80 -537
rect 205 -538 206 -516
rect 257 -577 258 -537
rect 282 -538 283 -516
rect 310 -538 311 -516
rect 765 -577 766 -537
rect 51 -540 52 -516
rect 205 -577 206 -539
rect 275 -577 276 -539
rect 306 -540 307 -516
rect 345 -540 346 -516
rect 373 -577 374 -539
rect 401 -540 402 -516
rect 576 -577 577 -539
rect 639 -577 640 -539
rect 660 -540 661 -516
rect 30 -542 31 -516
rect 345 -577 346 -541
rect 401 -577 402 -541
rect 415 -542 416 -516
rect 422 -542 423 -516
rect 429 -577 430 -541
rect 457 -577 458 -541
rect 716 -542 717 -516
rect 30 -577 31 -543
rect 198 -544 199 -516
rect 282 -577 283 -543
rect 506 -544 507 -516
rect 562 -577 563 -543
rect 597 -544 598 -516
rect 86 -546 87 -516
rect 352 -577 353 -545
rect 369 -546 370 -516
rect 716 -577 717 -545
rect 86 -577 87 -547
rect 261 -548 262 -516
rect 317 -577 318 -547
rect 660 -577 661 -547
rect 93 -577 94 -549
rect 170 -550 171 -516
rect 177 -577 178 -549
rect 268 -550 269 -516
rect 415 -577 416 -549
rect 611 -550 612 -516
rect 114 -552 115 -516
rect 394 -577 395 -551
rect 422 -577 423 -551
rect 436 -552 437 -516
rect 474 -552 475 -516
rect 569 -552 570 -516
rect 597 -577 598 -551
rect 632 -552 633 -516
rect 23 -554 24 -516
rect 114 -577 115 -553
rect 135 -577 136 -553
rect 268 -577 269 -553
rect 436 -577 437 -553
rect 464 -554 465 -516
rect 478 -554 479 -516
rect 551 -577 552 -553
rect 569 -577 570 -553
rect 604 -554 605 -516
rect 611 -577 612 -553
rect 723 -554 724 -516
rect 23 -577 24 -555
rect 324 -556 325 -516
rect 411 -556 412 -516
rect 723 -577 724 -555
rect 149 -558 150 -516
rect 261 -577 262 -557
rect 324 -577 325 -557
rect 338 -558 339 -516
rect 443 -558 444 -516
rect 478 -577 479 -557
rect 485 -558 486 -516
rect 527 -577 528 -557
rect 604 -577 605 -557
rect 674 -558 675 -516
rect 72 -560 73 -516
rect 443 -577 444 -559
rect 488 -577 489 -559
rect 702 -577 703 -559
rect 142 -562 143 -516
rect 149 -577 150 -561
rect 156 -562 157 -516
rect 212 -577 213 -561
rect 296 -562 297 -516
rect 338 -577 339 -561
rect 499 -562 500 -516
rect 730 -577 731 -561
rect 37 -564 38 -516
rect 156 -577 157 -563
rect 170 -577 171 -563
rect 289 -564 290 -516
rect 464 -577 465 -563
rect 499 -577 500 -563
rect 506 -577 507 -563
rect 590 -577 591 -563
rect 632 -577 633 -563
rect 646 -564 647 -516
rect 674 -577 675 -563
rect 751 -564 752 -516
rect 37 -577 38 -565
rect 107 -566 108 -516
rect 198 -577 199 -565
rect 366 -566 367 -516
rect 646 -577 647 -565
rect 667 -566 668 -516
rect 737 -566 738 -516
rect 751 -577 752 -565
rect 65 -568 66 -516
rect 142 -577 143 -567
rect 289 -577 290 -567
rect 485 -577 486 -567
rect 667 -577 668 -567
rect 688 -568 689 -516
rect 65 -577 66 -569
rect 247 -570 248 -516
rect 418 -577 419 -569
rect 737 -577 738 -569
rect 128 -572 129 -516
rect 366 -577 367 -571
rect 688 -577 689 -571
rect 695 -572 696 -516
rect 72 -577 73 -573
rect 128 -577 129 -573
rect 247 -577 248 -573
rect 254 -574 255 -516
rect 334 -577 335 -573
rect 695 -577 696 -573
rect 184 -577 185 -575
rect 254 -577 255 -575
rect 2 -666 3 -586
rect 72 -587 73 -585
rect 86 -587 87 -585
rect 86 -666 87 -586
rect 86 -587 87 -585
rect 86 -666 87 -586
rect 93 -587 94 -585
rect 93 -666 94 -586
rect 93 -587 94 -585
rect 93 -666 94 -586
rect 107 -587 108 -585
rect 156 -587 157 -585
rect 163 -587 164 -585
rect 369 -666 370 -586
rect 436 -587 437 -585
rect 436 -666 437 -586
rect 436 -587 437 -585
rect 436 -666 437 -586
rect 457 -666 458 -586
rect 555 -587 556 -585
rect 9 -589 10 -585
rect 292 -666 293 -588
rect 296 -589 297 -585
rect 394 -589 395 -585
rect 464 -589 465 -585
rect 509 -589 510 -585
rect 513 -589 514 -585
rect 632 -589 633 -585
rect 9 -666 10 -590
rect 331 -591 332 -585
rect 334 -591 335 -585
rect 730 -591 731 -585
rect 54 -666 55 -592
rect 345 -593 346 -585
rect 467 -593 468 -585
rect 576 -593 577 -585
rect 730 -666 731 -592
rect 807 -593 808 -585
rect 68 -666 69 -594
rect 282 -595 283 -585
rect 299 -666 300 -594
rect 366 -595 367 -585
rect 485 -595 486 -585
rect 681 -595 682 -585
rect 72 -666 73 -596
rect 100 -597 101 -585
rect 107 -666 108 -596
rect 744 -597 745 -585
rect 100 -666 101 -598
rect 460 -599 461 -585
rect 506 -599 507 -585
rect 653 -599 654 -585
rect 110 -601 111 -585
rect 184 -601 185 -585
rect 205 -601 206 -585
rect 257 -601 258 -585
rect 271 -666 272 -600
rect 394 -666 395 -600
rect 460 -666 461 -600
rect 681 -666 682 -600
rect 110 -666 111 -602
rect 240 -603 241 -585
rect 254 -603 255 -585
rect 632 -666 633 -602
rect 653 -666 654 -602
rect 737 -603 738 -585
rect 121 -605 122 -585
rect 408 -605 409 -585
rect 506 -666 507 -604
rect 541 -605 542 -585
rect 576 -666 577 -604
rect 611 -605 612 -585
rect 737 -666 738 -604
rect 793 -605 794 -585
rect 121 -666 122 -606
rect 177 -607 178 -585
rect 184 -666 185 -606
rect 478 -607 479 -585
rect 513 -666 514 -606
rect 562 -607 563 -585
rect 611 -666 612 -606
rect 688 -607 689 -585
rect 26 -609 27 -585
rect 688 -666 689 -608
rect 124 -611 125 -585
rect 772 -611 773 -585
rect 128 -666 129 -612
rect 170 -613 171 -585
rect 177 -666 178 -612
rect 289 -613 290 -585
rect 303 -613 304 -585
rect 317 -613 318 -585
rect 320 -613 321 -585
rect 408 -666 409 -612
rect 478 -666 479 -612
rect 492 -613 493 -585
rect 534 -613 535 -585
rect 555 -666 556 -612
rect 562 -666 563 -612
rect 618 -613 619 -585
rect 772 -666 773 -612
rect 800 -613 801 -585
rect 138 -615 139 -585
rect 142 -615 143 -585
rect 149 -615 150 -585
rect 317 -666 318 -614
rect 331 -666 332 -614
rect 373 -615 374 -585
rect 492 -666 493 -614
rect 527 -615 528 -585
rect 534 -666 535 -614
rect 590 -615 591 -585
rect 618 -666 619 -614
rect 702 -615 703 -585
rect 37 -617 38 -585
rect 142 -666 143 -616
rect 156 -666 157 -616
rect 296 -666 297 -616
rect 303 -666 304 -616
rect 359 -617 360 -585
rect 366 -666 367 -616
rect 814 -617 815 -585
rect 30 -619 31 -585
rect 37 -666 38 -618
rect 61 -666 62 -618
rect 149 -666 150 -618
rect 163 -666 164 -618
rect 226 -619 227 -585
rect 240 -666 241 -618
rect 247 -619 248 -585
rect 282 -666 283 -618
rect 324 -619 325 -585
rect 359 -666 360 -618
rect 422 -619 423 -585
rect 527 -666 528 -618
rect 583 -619 584 -585
rect 590 -666 591 -618
rect 660 -619 661 -585
rect 702 -666 703 -618
rect 751 -619 752 -585
rect 170 -666 171 -620
rect 229 -666 230 -620
rect 289 -666 290 -620
rect 485 -666 486 -620
rect 583 -666 584 -620
rect 604 -621 605 -585
rect 751 -666 752 -620
rect 786 -621 787 -585
rect 191 -623 192 -585
rect 254 -666 255 -622
rect 310 -623 311 -585
rect 625 -623 626 -585
rect 191 -666 192 -624
rect 345 -666 346 -624
rect 348 -666 349 -624
rect 660 -666 661 -624
rect 205 -666 206 -626
rect 233 -627 234 -585
rect 275 -627 276 -585
rect 310 -666 311 -626
rect 324 -666 325 -626
rect 352 -627 353 -585
rect 373 -666 374 -626
rect 443 -627 444 -585
rect 453 -666 454 -626
rect 786 -666 787 -626
rect 198 -629 199 -585
rect 233 -666 234 -628
rect 268 -629 269 -585
rect 275 -666 276 -628
rect 338 -629 339 -585
rect 352 -666 353 -628
rect 422 -666 423 -628
rect 429 -629 430 -585
rect 443 -666 444 -628
rect 516 -629 517 -585
rect 548 -629 549 -585
rect 604 -666 605 -628
rect 625 -666 626 -628
rect 709 -629 710 -585
rect 65 -631 66 -585
rect 198 -666 199 -630
rect 212 -631 213 -585
rect 268 -666 269 -630
rect 338 -666 339 -630
rect 387 -631 388 -585
rect 548 -666 549 -630
rect 597 -631 598 -585
rect 709 -666 710 -630
rect 779 -631 780 -585
rect 30 -666 31 -632
rect 212 -666 213 -632
rect 215 -666 216 -632
rect 723 -633 724 -585
rect 758 -633 759 -585
rect 779 -666 780 -632
rect 219 -635 220 -585
rect 247 -666 248 -634
rect 380 -635 381 -585
rect 723 -666 724 -634
rect 758 -666 759 -634
rect 793 -666 794 -634
rect 51 -666 52 -636
rect 219 -666 220 -636
rect 226 -666 227 -636
rect 261 -637 262 -585
rect 383 -637 384 -585
rect 429 -666 430 -636
rect 597 -666 598 -636
rect 667 -637 668 -585
rect 44 -639 45 -585
rect 261 -666 262 -638
rect 383 -666 384 -638
rect 464 -666 465 -638
rect 646 -639 647 -585
rect 667 -666 668 -638
rect 44 -666 45 -640
rect 313 -641 314 -585
rect 387 -666 388 -640
rect 401 -641 402 -585
rect 646 -666 647 -640
rect 695 -641 696 -585
rect 16 -643 17 -585
rect 401 -666 402 -642
rect 499 -643 500 -585
rect 695 -666 696 -642
rect 16 -666 17 -644
rect 58 -645 59 -585
rect 499 -666 500 -644
rect 639 -645 640 -585
rect 58 -666 59 -646
rect 135 -647 136 -585
rect 639 -666 640 -646
rect 716 -647 717 -585
rect 79 -649 80 -585
rect 135 -666 136 -648
rect 674 -649 675 -585
rect 716 -666 717 -648
rect 79 -666 80 -650
rect 114 -651 115 -585
rect 674 -666 675 -650
rect 765 -651 766 -585
rect 23 -653 24 -585
rect 114 -666 115 -652
rect 415 -653 416 -585
rect 765 -666 766 -652
rect 23 -666 24 -654
rect 450 -655 451 -585
rect 415 -666 416 -656
rect 744 -666 745 -656
rect 450 -666 451 -658
rect 471 -659 472 -585
rect 471 -666 472 -660
rect 520 -661 521 -585
rect 520 -666 521 -662
rect 569 -663 570 -585
rect 569 -666 570 -664
rect 821 -665 822 -585
rect 2 -676 3 -674
rect 89 -733 90 -675
rect 100 -676 101 -674
rect 100 -733 101 -675
rect 100 -676 101 -674
rect 100 -733 101 -675
rect 142 -676 143 -674
rect 418 -676 419 -674
rect 425 -733 426 -675
rect 506 -676 507 -674
rect 520 -676 521 -674
rect 523 -733 524 -675
rect 551 -733 552 -675
rect 660 -676 661 -674
rect 751 -676 752 -674
rect 751 -733 752 -675
rect 751 -676 752 -674
rect 751 -733 752 -675
rect 765 -676 766 -674
rect 765 -733 766 -675
rect 765 -676 766 -674
rect 765 -733 766 -675
rect 779 -676 780 -674
rect 786 -733 787 -675
rect 16 -678 17 -674
rect 68 -678 69 -674
rect 142 -733 143 -677
rect 163 -678 164 -674
rect 177 -678 178 -674
rect 177 -733 178 -677
rect 177 -678 178 -674
rect 177 -733 178 -677
rect 184 -678 185 -674
rect 348 -678 349 -674
rect 415 -678 416 -674
rect 436 -678 437 -674
rect 446 -733 447 -677
rect 527 -678 528 -674
rect 625 -678 626 -674
rect 625 -733 626 -677
rect 625 -678 626 -674
rect 625 -733 626 -677
rect 639 -678 640 -674
rect 639 -733 640 -677
rect 639 -678 640 -674
rect 639 -733 640 -677
rect 660 -733 661 -677
rect 674 -678 675 -674
rect 779 -733 780 -677
rect 807 -733 808 -677
rect 16 -733 17 -679
rect 93 -680 94 -674
rect 107 -680 108 -674
rect 436 -733 437 -679
rect 450 -733 451 -679
rect 485 -680 486 -674
rect 499 -680 500 -674
rect 502 -712 503 -679
rect 527 -733 528 -679
rect 709 -680 710 -674
rect 51 -682 52 -674
rect 86 -682 87 -674
rect 107 -733 108 -681
rect 268 -682 269 -674
rect 271 -682 272 -674
rect 667 -682 668 -674
rect 37 -684 38 -674
rect 51 -733 52 -683
rect 58 -733 59 -683
rect 121 -684 122 -674
rect 149 -684 150 -674
rect 184 -733 185 -683
rect 212 -684 213 -674
rect 317 -684 318 -674
rect 415 -733 416 -683
rect 429 -684 430 -674
rect 453 -684 454 -674
rect 653 -684 654 -674
rect 9 -686 10 -674
rect 317 -733 318 -685
rect 457 -733 458 -685
rect 464 -686 465 -674
rect 471 -686 472 -674
rect 800 -733 801 -685
rect 37 -733 38 -687
rect 79 -688 80 -674
rect 93 -733 94 -687
rect 271 -733 272 -687
rect 296 -688 297 -674
rect 772 -688 773 -674
rect 61 -690 62 -674
rect 170 -690 171 -674
rect 198 -690 199 -674
rect 296 -733 297 -689
rect 310 -690 311 -674
rect 429 -733 430 -689
rect 443 -690 444 -674
rect 471 -733 472 -689
rect 485 -733 486 -689
rect 492 -690 493 -674
rect 499 -733 500 -689
rect 513 -690 514 -674
rect 604 -690 605 -674
rect 667 -733 668 -689
rect 772 -733 773 -689
rect 793 -733 794 -689
rect 12 -733 13 -691
rect 310 -733 311 -691
rect 443 -733 444 -691
rect 737 -692 738 -674
rect 68 -733 69 -693
rect 79 -733 80 -693
rect 114 -694 115 -674
rect 121 -733 122 -693
rect 135 -694 136 -674
rect 149 -733 150 -693
rect 156 -694 157 -674
rect 156 -733 157 -693
rect 156 -694 157 -674
rect 156 -733 157 -693
rect 170 -733 171 -693
rect 261 -694 262 -674
rect 268 -733 269 -693
rect 366 -733 367 -693
rect 460 -694 461 -674
rect 737 -733 738 -693
rect 72 -696 73 -674
rect 163 -733 164 -695
rect 198 -733 199 -695
rect 240 -696 241 -674
rect 261 -733 262 -695
rect 303 -696 304 -674
rect 464 -733 465 -695
rect 534 -696 535 -674
rect 583 -696 584 -674
rect 604 -733 605 -695
rect 646 -696 647 -674
rect 674 -733 675 -695
rect 23 -698 24 -674
rect 72 -733 73 -697
rect 114 -733 115 -697
rect 128 -698 129 -674
rect 135 -733 136 -697
rect 229 -698 230 -674
rect 233 -698 234 -674
rect 289 -733 290 -697
rect 303 -733 304 -697
rect 369 -698 370 -674
rect 492 -733 493 -697
rect 569 -698 570 -674
rect 583 -733 584 -697
rect 611 -698 612 -674
rect 646 -733 647 -697
rect 702 -698 703 -674
rect 23 -733 24 -699
rect 191 -700 192 -674
rect 212 -733 213 -699
rect 254 -700 255 -674
rect 513 -733 514 -699
rect 555 -700 556 -674
rect 590 -700 591 -674
rect 611 -733 612 -699
rect 618 -700 619 -674
rect 702 -733 703 -699
rect 44 -702 45 -674
rect 128 -733 129 -701
rect 191 -733 192 -701
rect 205 -702 206 -674
rect 226 -733 227 -701
rect 709 -733 710 -701
rect 44 -733 45 -703
rect 65 -704 66 -674
rect 205 -733 206 -703
rect 219 -704 220 -674
rect 229 -733 230 -703
rect 380 -704 381 -674
rect 534 -733 535 -703
rect 782 -733 783 -703
rect 30 -706 31 -674
rect 65 -733 66 -705
rect 219 -733 220 -705
rect 408 -706 409 -674
rect 544 -706 545 -674
rect 590 -733 591 -705
rect 618 -733 619 -705
rect 688 -706 689 -674
rect 30 -733 31 -707
rect 324 -708 325 -674
rect 345 -733 346 -707
rect 408 -733 409 -707
rect 555 -733 556 -707
rect 562 -708 563 -674
rect 597 -708 598 -674
rect 688 -733 689 -707
rect 233 -733 234 -709
rect 247 -710 248 -674
rect 254 -733 255 -709
rect 338 -710 339 -674
rect 380 -733 381 -709
rect 695 -710 696 -674
rect 240 -733 241 -711
rect 275 -712 276 -674
rect 324 -733 325 -711
rect 359 -712 360 -674
rect 562 -733 563 -711
rect 597 -733 598 -711
rect 632 -712 633 -674
rect 653 -733 654 -711
rect 681 -712 682 -674
rect 695 -733 696 -711
rect 716 -712 717 -674
rect 166 -733 167 -713
rect 359 -733 360 -713
rect 478 -714 479 -674
rect 716 -733 717 -713
rect 247 -733 248 -715
rect 331 -716 332 -674
rect 338 -733 339 -715
rect 352 -716 353 -674
rect 478 -733 479 -715
rect 548 -716 549 -674
rect 576 -716 577 -674
rect 632 -733 633 -715
rect 681 -733 682 -715
rect 723 -716 724 -674
rect 275 -733 276 -717
rect 282 -718 283 -674
rect 331 -733 332 -717
rect 387 -718 388 -674
rect 530 -733 531 -717
rect 576 -733 577 -717
rect 723 -733 724 -717
rect 744 -718 745 -674
rect 282 -733 283 -719
rect 394 -720 395 -674
rect 744 -733 745 -719
rect 758 -720 759 -674
rect 320 -733 321 -721
rect 387 -733 388 -721
rect 394 -733 395 -721
rect 506 -733 507 -721
rect 730 -722 731 -674
rect 758 -733 759 -721
rect 131 -733 132 -723
rect 730 -733 731 -723
rect 352 -733 353 -725
rect 373 -726 374 -674
rect 373 -733 374 -727
rect 401 -728 402 -674
rect 401 -733 402 -729
rect 422 -730 423 -674
rect 422 -733 423 -731
rect 541 -733 542 -731
rect 2 -804 3 -742
rect 226 -804 227 -742
rect 268 -743 269 -741
rect 275 -743 276 -741
rect 289 -743 290 -741
rect 348 -743 349 -741
rect 397 -743 398 -741
rect 464 -743 465 -741
rect 481 -804 482 -742
rect 569 -743 570 -741
rect 572 -743 573 -741
rect 737 -743 738 -741
rect 765 -743 766 -741
rect 765 -804 766 -742
rect 765 -743 766 -741
rect 765 -804 766 -742
rect 782 -743 783 -741
rect 786 -743 787 -741
rect 793 -743 794 -741
rect 807 -743 808 -741
rect 9 -804 10 -744
rect 128 -804 129 -744
rect 166 -745 167 -741
rect 219 -745 220 -741
rect 268 -804 269 -744
rect 387 -745 388 -741
rect 422 -745 423 -741
rect 702 -745 703 -741
rect 737 -804 738 -744
rect 744 -745 745 -741
rect 16 -804 17 -746
rect 58 -747 59 -741
rect 65 -804 66 -746
rect 72 -747 73 -741
rect 79 -747 80 -741
rect 317 -747 318 -741
rect 345 -747 346 -741
rect 688 -747 689 -741
rect 702 -804 703 -746
rect 723 -747 724 -741
rect 744 -804 745 -746
rect 751 -747 752 -741
rect 30 -749 31 -741
rect 229 -749 230 -741
rect 275 -804 276 -748
rect 296 -749 297 -741
rect 310 -749 311 -741
rect 345 -804 346 -748
rect 366 -749 367 -741
rect 464 -804 465 -748
rect 506 -749 507 -741
rect 569 -804 570 -748
rect 576 -749 577 -741
rect 786 -804 787 -748
rect 19 -751 20 -741
rect 366 -804 367 -750
rect 376 -804 377 -750
rect 506 -804 507 -750
rect 513 -751 514 -741
rect 513 -804 514 -750
rect 513 -751 514 -741
rect 513 -804 514 -750
rect 520 -804 521 -750
rect 555 -751 556 -741
rect 562 -751 563 -741
rect 562 -804 563 -750
rect 562 -751 563 -741
rect 562 -804 563 -750
rect 600 -804 601 -750
rect 660 -751 661 -741
rect 751 -804 752 -750
rect 758 -751 759 -741
rect 30 -804 31 -752
rect 44 -753 45 -741
rect 58 -804 59 -752
rect 121 -753 122 -741
rect 184 -753 185 -741
rect 215 -804 216 -752
rect 233 -753 234 -741
rect 296 -804 297 -752
rect 310 -804 311 -752
rect 352 -753 353 -741
rect 380 -753 381 -741
rect 688 -804 689 -752
rect 758 -804 759 -752
rect 772 -753 773 -741
rect 40 -804 41 -754
rect 163 -804 164 -754
rect 184 -804 185 -754
rect 212 -755 213 -741
rect 282 -755 283 -741
rect 387 -804 388 -754
rect 408 -755 409 -741
rect 422 -804 423 -754
rect 446 -755 447 -741
rect 723 -804 724 -754
rect 772 -804 773 -754
rect 779 -804 780 -754
rect 44 -804 45 -756
rect 411 -804 412 -756
rect 450 -757 451 -741
rect 453 -757 454 -741
rect 530 -757 531 -741
rect 639 -757 640 -741
rect 653 -757 654 -741
rect 653 -804 654 -756
rect 653 -757 654 -741
rect 653 -804 654 -756
rect 72 -804 73 -758
rect 177 -759 178 -741
rect 198 -759 199 -741
rect 201 -777 202 -758
rect 205 -759 206 -741
rect 219 -804 220 -758
rect 247 -759 248 -741
rect 282 -804 283 -758
rect 289 -804 290 -758
rect 373 -759 374 -741
rect 450 -804 451 -758
rect 492 -759 493 -741
rect 541 -759 542 -741
rect 576 -804 577 -758
rect 618 -759 619 -741
rect 660 -804 661 -758
rect 75 -804 76 -760
rect 205 -804 206 -760
rect 233 -804 234 -760
rect 247 -804 248 -760
rect 320 -761 321 -741
rect 618 -804 619 -760
rect 625 -761 626 -741
rect 625 -804 626 -760
rect 625 -761 626 -741
rect 625 -804 626 -760
rect 632 -761 633 -741
rect 639 -804 640 -760
rect 79 -804 80 -762
rect 303 -763 304 -741
rect 331 -763 332 -741
rect 352 -804 353 -762
rect 359 -763 360 -741
rect 380 -804 381 -762
rect 485 -763 486 -741
rect 492 -804 493 -762
rect 534 -763 535 -741
rect 541 -804 542 -762
rect 548 -763 549 -741
rect 604 -763 605 -741
rect 86 -765 87 -741
rect 383 -765 384 -741
rect 471 -765 472 -741
rect 534 -804 535 -764
rect 551 -804 552 -764
rect 667 -765 668 -741
rect 86 -804 87 -766
rect 100 -767 101 -741
rect 107 -767 108 -741
rect 121 -804 122 -766
rect 177 -804 178 -766
rect 261 -767 262 -741
rect 303 -804 304 -766
rect 338 -767 339 -741
rect 359 -804 360 -766
rect 457 -767 458 -741
rect 471 -804 472 -766
rect 478 -767 479 -741
rect 555 -804 556 -766
rect 590 -767 591 -741
rect 597 -767 598 -741
rect 632 -804 633 -766
rect 667 -804 668 -766
rect 695 -767 696 -741
rect 89 -769 90 -741
rect 681 -769 682 -741
rect 695 -804 696 -768
rect 709 -769 710 -741
rect 93 -771 94 -741
rect 317 -804 318 -770
rect 324 -771 325 -741
rect 338 -804 339 -770
rect 362 -804 363 -770
rect 590 -804 591 -770
rect 646 -771 647 -741
rect 681 -804 682 -770
rect 23 -773 24 -741
rect 93 -804 94 -772
rect 100 -804 101 -772
rect 149 -773 150 -741
rect 170 -773 171 -741
rect 261 -804 262 -772
rect 373 -804 374 -772
rect 716 -773 717 -741
rect 23 -804 24 -774
rect 135 -775 136 -741
rect 149 -804 150 -774
rect 191 -775 192 -741
rect 198 -804 199 -774
rect 254 -775 255 -741
rect 324 -804 325 -774
rect 404 -804 405 -774
rect 597 -804 598 -774
rect 646 -804 647 -774
rect 674 -775 675 -741
rect 716 -804 717 -774
rect 730 -775 731 -741
rect 51 -777 52 -741
rect 170 -804 171 -776
rect 191 -804 192 -776
rect 443 -777 444 -741
rect 453 -804 454 -776
rect 485 -804 486 -776
rect 548 -804 549 -776
rect 730 -804 731 -776
rect 51 -804 52 -778
rect 425 -779 426 -741
rect 443 -804 444 -778
rect 527 -779 528 -741
rect 583 -779 584 -741
rect 604 -804 605 -778
rect 107 -804 108 -780
rect 114 -781 115 -741
rect 135 -804 136 -780
rect 142 -781 143 -741
rect 159 -804 160 -780
rect 527 -804 528 -780
rect 37 -783 38 -741
rect 114 -804 115 -782
rect 142 -804 143 -782
rect 156 -783 157 -741
rect 212 -804 213 -782
rect 331 -804 332 -782
rect 457 -804 458 -782
rect 800 -783 801 -741
rect 37 -804 38 -784
rect 611 -785 612 -741
rect 254 -804 255 -786
rect 674 -804 675 -786
rect 285 -804 286 -788
rect 611 -804 612 -788
rect 478 -804 479 -790
rect 709 -804 710 -790
rect 499 -793 500 -741
rect 583 -804 584 -792
rect 436 -795 437 -741
rect 499 -804 500 -794
rect 429 -797 430 -741
rect 436 -804 437 -796
rect 415 -799 416 -741
rect 429 -804 430 -798
rect 401 -801 402 -741
rect 415 -804 416 -800
rect 68 -803 69 -741
rect 401 -804 402 -802
rect 23 -814 24 -812
rect 156 -814 157 -812
rect 170 -814 171 -812
rect 250 -814 251 -812
rect 254 -859 255 -813
rect 275 -814 276 -812
rect 282 -814 283 -812
rect 296 -814 297 -812
rect 310 -859 311 -813
rect 380 -814 381 -812
rect 394 -859 395 -813
rect 429 -814 430 -812
rect 450 -814 451 -812
rect 450 -859 451 -813
rect 450 -814 451 -812
rect 450 -859 451 -813
rect 478 -859 479 -813
rect 527 -814 528 -812
rect 544 -859 545 -813
rect 681 -814 682 -812
rect 737 -814 738 -812
rect 737 -859 738 -813
rect 737 -814 738 -812
rect 737 -859 738 -813
rect 9 -816 10 -812
rect 23 -859 24 -815
rect 30 -816 31 -812
rect 40 -816 41 -812
rect 65 -816 66 -812
rect 131 -816 132 -812
rect 156 -859 157 -815
rect 233 -816 234 -812
rect 240 -816 241 -812
rect 257 -816 258 -812
rect 261 -816 262 -812
rect 261 -859 262 -815
rect 261 -816 262 -812
rect 261 -859 262 -815
rect 271 -859 272 -815
rect 443 -816 444 -812
rect 481 -816 482 -812
rect 562 -816 563 -812
rect 597 -816 598 -812
rect 744 -816 745 -812
rect 9 -859 10 -817
rect 128 -818 129 -812
rect 177 -818 178 -812
rect 212 -859 213 -817
rect 219 -818 220 -812
rect 222 -834 223 -817
rect 226 -818 227 -812
rect 376 -818 377 -812
rect 397 -818 398 -812
rect 485 -818 486 -812
rect 513 -818 514 -812
rect 527 -859 528 -817
rect 548 -818 549 -812
rect 646 -818 647 -812
rect 744 -859 745 -817
rect 786 -818 787 -812
rect 16 -820 17 -812
rect 65 -859 66 -819
rect 72 -820 73 -812
rect 86 -820 87 -812
rect 93 -820 94 -812
rect 226 -859 227 -819
rect 240 -859 241 -819
rect 422 -820 423 -812
rect 429 -859 430 -819
rect 457 -820 458 -812
rect 485 -859 486 -819
rect 569 -820 570 -812
rect 618 -820 619 -812
rect 765 -820 766 -812
rect 86 -859 87 -821
rect 114 -822 115 -812
rect 117 -859 118 -821
rect 159 -822 160 -812
rect 184 -822 185 -812
rect 233 -859 234 -821
rect 275 -859 276 -821
rect 331 -822 332 -812
rect 345 -822 346 -812
rect 401 -859 402 -821
rect 408 -859 409 -821
rect 502 -859 503 -821
rect 513 -859 514 -821
rect 520 -822 521 -812
rect 548 -859 549 -821
rect 604 -822 605 -812
rect 618 -859 619 -821
rect 702 -822 703 -812
rect 75 -824 76 -812
rect 114 -859 115 -823
rect 121 -824 122 -812
rect 128 -859 129 -823
rect 135 -824 136 -812
rect 177 -859 178 -823
rect 184 -859 185 -823
rect 205 -824 206 -812
rect 219 -859 220 -823
rect 303 -824 304 -812
rect 331 -859 332 -823
rect 338 -824 339 -812
rect 345 -859 346 -823
rect 590 -824 591 -812
rect 646 -859 647 -823
rect 716 -824 717 -812
rect 93 -859 94 -825
rect 107 -826 108 -812
rect 110 -859 111 -825
rect 191 -826 192 -812
rect 205 -859 206 -825
rect 268 -826 269 -812
rect 282 -859 283 -825
rect 436 -826 437 -812
rect 443 -859 444 -825
rect 506 -826 507 -812
rect 562 -859 563 -825
rect 611 -826 612 -812
rect 702 -859 703 -825
rect 751 -826 752 -812
rect 72 -859 73 -827
rect 107 -859 108 -827
rect 121 -859 122 -827
rect 149 -828 150 -812
rect 191 -859 192 -827
rect 324 -828 325 -812
rect 338 -859 339 -827
rect 387 -828 388 -812
rect 404 -828 405 -812
rect 506 -859 507 -827
rect 569 -859 570 -827
rect 632 -828 633 -812
rect 751 -859 752 -827
rect 758 -828 759 -812
rect 79 -830 80 -812
rect 268 -859 269 -829
rect 296 -859 297 -829
rect 317 -830 318 -812
rect 348 -859 349 -829
rect 688 -830 689 -812
rect 758 -859 759 -829
rect 779 -830 780 -812
rect 51 -832 52 -812
rect 79 -859 80 -831
rect 100 -832 101 -812
rect 149 -859 150 -831
rect 163 -832 164 -812
rect 317 -859 318 -831
rect 359 -859 360 -831
rect 390 -859 391 -831
rect 411 -832 412 -812
rect 583 -832 584 -812
rect 590 -859 591 -831
rect 639 -832 640 -812
rect 688 -859 689 -831
rect 726 -859 727 -831
rect 30 -859 31 -833
rect 51 -859 52 -833
rect 142 -834 143 -812
rect 163 -859 164 -833
rect 303 -859 304 -833
rect 366 -834 367 -812
rect 520 -859 521 -833
rect 583 -859 584 -833
rect 653 -834 654 -812
rect 44 -836 45 -812
rect 100 -859 101 -835
rect 247 -836 248 -812
rect 387 -859 388 -835
rect 422 -859 423 -835
rect 492 -836 493 -812
rect 611 -859 612 -835
rect 674 -836 675 -812
rect 44 -859 45 -837
rect 138 -859 139 -837
rect 198 -838 199 -812
rect 247 -859 248 -837
rect 324 -859 325 -837
rect 366 -859 367 -837
rect 373 -838 374 -812
rect 597 -859 598 -837
rect 632 -859 633 -837
rect 660 -838 661 -812
rect 58 -840 59 -812
rect 142 -859 143 -839
rect 198 -859 199 -839
rect 289 -840 290 -812
rect 373 -859 374 -839
rect 464 -840 465 -812
rect 492 -859 493 -839
rect 607 -859 608 -839
rect 639 -859 640 -839
rect 667 -840 668 -812
rect 58 -859 59 -841
rect 173 -859 174 -841
rect 264 -859 265 -841
rect 464 -859 465 -841
rect 653 -859 654 -841
rect 695 -842 696 -812
rect 289 -859 290 -843
rect 352 -844 353 -812
rect 380 -859 381 -843
rect 660 -859 661 -843
rect 667 -859 668 -843
rect 723 -844 724 -812
rect 352 -859 353 -845
rect 415 -846 416 -812
rect 436 -859 437 -845
rect 471 -846 472 -812
rect 695 -859 696 -845
rect 730 -846 731 -812
rect 415 -859 416 -847
rect 541 -848 542 -812
rect 457 -859 458 -849
rect 534 -850 535 -812
rect 471 -859 472 -851
rect 499 -852 500 -812
rect 534 -859 535 -851
rect 555 -852 556 -812
rect 555 -859 556 -853
rect 576 -854 577 -812
rect 576 -859 577 -855
rect 625 -856 626 -812
rect 625 -859 626 -857
rect 709 -858 710 -812
rect 9 -869 10 -867
rect 397 -912 398 -868
rect 471 -869 472 -867
rect 523 -912 524 -868
rect 544 -869 545 -867
rect 583 -869 584 -867
rect 604 -869 605 -867
rect 730 -869 731 -867
rect 733 -869 734 -867
rect 737 -869 738 -867
rect 747 -912 748 -868
rect 751 -869 752 -867
rect 19 -871 20 -867
rect 23 -871 24 -867
rect 51 -912 52 -870
rect 93 -871 94 -867
rect 114 -912 115 -870
rect 117 -871 118 -867
rect 124 -912 125 -870
rect 478 -871 479 -867
rect 499 -912 500 -870
rect 534 -871 535 -867
rect 583 -912 584 -870
rect 597 -871 598 -867
rect 604 -912 605 -870
rect 639 -871 640 -867
rect 663 -912 664 -870
rect 688 -871 689 -867
rect 726 -871 727 -867
rect 758 -871 759 -867
rect 54 -873 55 -867
rect 107 -873 108 -867
rect 135 -873 136 -867
rect 177 -873 178 -867
rect 180 -912 181 -872
rect 275 -873 276 -867
rect 282 -873 283 -867
rect 383 -873 384 -867
rect 387 -912 388 -872
rect 422 -873 423 -867
rect 502 -873 503 -867
rect 632 -873 633 -867
rect 674 -912 675 -872
rect 702 -873 703 -867
rect 30 -875 31 -867
rect 282 -912 283 -874
rect 317 -875 318 -867
rect 380 -912 381 -874
rect 390 -875 391 -867
rect 450 -875 451 -867
rect 520 -875 521 -867
rect 597 -912 598 -874
rect 632 -912 633 -874
rect 646 -875 647 -867
rect 681 -875 682 -867
rect 744 -875 745 -867
rect 58 -877 59 -867
rect 177 -912 178 -876
rect 212 -877 213 -867
rect 299 -912 300 -876
rect 317 -912 318 -876
rect 338 -877 339 -867
rect 345 -912 346 -876
rect 541 -877 542 -867
rect 642 -912 643 -876
rect 646 -912 647 -876
rect 681 -912 682 -876
rect 695 -877 696 -867
rect 58 -912 59 -878
rect 86 -879 87 -867
rect 93 -912 94 -878
rect 110 -879 111 -867
rect 121 -879 122 -867
rect 135 -912 136 -878
rect 142 -879 143 -867
rect 145 -893 146 -878
rect 149 -879 150 -867
rect 170 -879 171 -867
rect 257 -912 258 -878
rect 303 -879 304 -867
rect 352 -879 353 -867
rect 369 -879 370 -867
rect 401 -879 402 -867
rect 422 -912 423 -878
rect 450 -912 451 -878
rect 527 -879 528 -867
rect 534 -912 535 -878
rect 576 -879 577 -867
rect 684 -879 685 -867
rect 716 -912 717 -878
rect 65 -881 66 -867
rect 348 -881 349 -867
rect 352 -912 353 -880
rect 394 -881 395 -867
rect 401 -912 402 -880
rect 443 -881 444 -867
rect 527 -912 528 -880
rect 569 -881 570 -867
rect 576 -912 577 -880
rect 618 -881 619 -867
rect 65 -912 66 -882
rect 219 -883 220 -867
rect 261 -912 262 -882
rect 373 -883 374 -867
rect 394 -912 395 -882
rect 653 -883 654 -867
rect 79 -885 80 -867
rect 149 -912 150 -884
rect 163 -885 164 -867
rect 163 -912 164 -884
rect 163 -885 164 -867
rect 163 -912 164 -884
rect 170 -912 171 -884
rect 310 -885 311 -867
rect 366 -885 367 -867
rect 443 -912 444 -884
rect 492 -885 493 -867
rect 569 -912 570 -884
rect 618 -912 619 -884
rect 667 -885 668 -867
rect 79 -912 80 -886
rect 240 -887 241 -867
rect 271 -887 272 -867
rect 296 -887 297 -867
rect 303 -912 304 -886
rect 331 -887 332 -867
rect 373 -912 374 -886
rect 478 -912 479 -886
rect 541 -912 542 -886
rect 562 -887 563 -867
rect 86 -912 87 -888
rect 138 -889 139 -867
rect 142 -912 143 -888
rect 191 -889 192 -867
rect 198 -889 199 -867
rect 240 -912 241 -888
rect 271 -912 272 -888
rect 376 -912 377 -888
rect 464 -889 465 -867
rect 492 -912 493 -888
rect 555 -889 556 -867
rect 667 -912 668 -888
rect 100 -891 101 -867
rect 212 -912 213 -890
rect 219 -912 220 -890
rect 254 -891 255 -867
rect 275 -912 276 -890
rect 324 -891 325 -867
rect 331 -912 332 -890
rect 436 -891 437 -867
rect 562 -912 563 -890
rect 590 -891 591 -867
rect 72 -893 73 -867
rect 100 -912 101 -892
rect 107 -912 108 -892
rect 128 -893 129 -867
rect 191 -912 192 -892
rect 198 -912 199 -892
rect 233 -893 234 -867
rect 289 -893 290 -867
rect 338 -912 339 -892
rect 415 -893 416 -867
rect 436 -912 437 -892
rect 590 -912 591 -892
rect 611 -893 612 -867
rect 72 -912 73 -894
rect 226 -895 227 -867
rect 289 -912 290 -894
rect 408 -895 409 -867
rect 415 -912 416 -894
rect 467 -912 468 -894
rect 611 -912 612 -894
rect 625 -895 626 -867
rect 40 -897 41 -867
rect 226 -912 227 -896
rect 310 -912 311 -896
rect 359 -897 360 -867
rect 408 -912 409 -896
rect 429 -897 430 -867
rect 625 -912 626 -896
rect 660 -897 661 -867
rect 128 -912 129 -898
rect 156 -899 157 -867
rect 173 -899 174 -867
rect 555 -912 556 -898
rect 156 -912 157 -900
rect 359 -912 360 -900
rect 429 -912 430 -900
rect 457 -901 458 -867
rect 506 -901 507 -867
rect 660 -912 661 -900
rect 184 -903 185 -867
rect 233 -912 234 -902
rect 457 -912 458 -902
rect 485 -903 486 -867
rect 506 -912 507 -902
rect 548 -903 549 -867
rect 184 -912 185 -904
rect 247 -905 248 -867
rect 296 -912 297 -904
rect 548 -912 549 -904
rect 44 -907 45 -867
rect 247 -912 248 -906
rect 485 -912 486 -906
rect 513 -907 514 -867
rect 44 -912 45 -908
rect 205 -909 206 -867
rect 208 -912 209 -908
rect 513 -912 514 -908
rect 205 -912 206 -910
rect 471 -912 472 -910
rect 44 -922 45 -920
rect 453 -971 454 -921
rect 464 -922 465 -920
rect 492 -922 493 -920
rect 520 -922 521 -920
rect 576 -922 577 -920
rect 646 -922 647 -920
rect 653 -922 654 -920
rect 660 -971 661 -921
rect 674 -922 675 -920
rect 716 -922 717 -920
rect 744 -922 745 -920
rect 51 -924 52 -920
rect 121 -924 122 -920
rect 135 -924 136 -920
rect 135 -971 136 -923
rect 135 -924 136 -920
rect 135 -971 136 -923
rect 163 -924 164 -920
rect 163 -971 164 -923
rect 163 -924 164 -920
rect 163 -971 164 -923
rect 170 -924 171 -920
rect 177 -971 178 -923
rect 191 -924 192 -920
rect 205 -924 206 -920
rect 219 -924 220 -920
rect 268 -924 269 -920
rect 282 -924 283 -920
rect 313 -971 314 -923
rect 320 -971 321 -923
rect 422 -924 423 -920
rect 464 -971 465 -923
rect 555 -924 556 -920
rect 674 -971 675 -923
rect 681 -924 682 -920
rect 72 -971 73 -925
rect 93 -926 94 -920
rect 103 -971 104 -925
rect 121 -971 122 -925
rect 142 -926 143 -920
rect 219 -971 220 -925
rect 226 -926 227 -920
rect 425 -971 426 -925
rect 492 -971 493 -925
rect 569 -926 570 -920
rect 107 -928 108 -920
rect 156 -928 157 -920
rect 159 -928 160 -920
rect 170 -971 171 -927
rect 184 -928 185 -920
rect 205 -971 206 -927
rect 240 -928 241 -920
rect 324 -928 325 -920
rect 394 -971 395 -927
rect 429 -928 430 -920
rect 499 -928 500 -920
rect 576 -971 577 -927
rect 86 -930 87 -920
rect 107 -971 108 -929
rect 128 -930 129 -920
rect 142 -971 143 -929
rect 184 -971 185 -929
rect 233 -930 234 -920
rect 240 -971 241 -929
rect 352 -930 353 -920
rect 499 -971 500 -929
rect 618 -930 619 -920
rect 58 -932 59 -920
rect 86 -971 87 -931
rect 100 -932 101 -920
rect 128 -971 129 -931
rect 191 -971 192 -931
rect 366 -932 367 -920
rect 527 -932 528 -920
rect 569 -971 570 -931
rect 618 -971 619 -931
rect 639 -932 640 -920
rect 114 -934 115 -920
rect 233 -971 234 -933
rect 254 -934 255 -920
rect 429 -971 430 -933
rect 450 -934 451 -920
rect 527 -971 528 -933
rect 541 -934 542 -920
rect 642 -934 643 -920
rect 198 -936 199 -920
rect 541 -971 542 -935
rect 555 -971 556 -935
rect 611 -936 612 -920
rect 149 -938 150 -920
rect 198 -971 199 -937
rect 254 -971 255 -937
rect 436 -938 437 -920
rect 534 -938 535 -920
rect 611 -971 612 -937
rect 149 -971 150 -939
rect 226 -971 227 -939
rect 268 -971 269 -939
rect 317 -940 318 -920
rect 324 -971 325 -939
rect 471 -940 472 -920
rect 156 -971 157 -941
rect 317 -971 318 -941
rect 352 -971 353 -941
rect 415 -942 416 -920
rect 436 -971 437 -941
rect 457 -942 458 -920
rect 471 -971 472 -941
rect 485 -942 486 -920
rect 275 -944 276 -920
rect 282 -971 283 -943
rect 289 -944 290 -920
rect 299 -944 300 -920
rect 310 -944 311 -920
rect 544 -971 545 -943
rect 79 -946 80 -920
rect 289 -971 290 -945
rect 296 -971 297 -945
rect 338 -946 339 -920
rect 366 -971 367 -945
rect 632 -946 633 -920
rect 79 -971 80 -947
rect 303 -948 304 -920
rect 338 -971 339 -947
rect 359 -948 360 -920
rect 408 -948 409 -920
rect 534 -971 535 -947
rect 275 -971 276 -949
rect 345 -950 346 -920
rect 359 -971 360 -949
rect 380 -950 381 -920
rect 408 -971 409 -949
rect 443 -950 444 -920
rect 457 -971 458 -949
rect 583 -950 584 -920
rect 247 -952 248 -920
rect 345 -971 346 -951
rect 380 -971 381 -951
rect 387 -952 388 -920
rect 443 -971 444 -951
rect 513 -952 514 -920
rect 583 -971 584 -951
rect 597 -952 598 -920
rect 212 -954 213 -920
rect 247 -971 248 -953
rect 303 -971 304 -953
rect 369 -954 370 -920
rect 478 -954 479 -920
rect 485 -971 486 -953
rect 513 -971 514 -953
rect 562 -954 563 -920
rect 65 -956 66 -920
rect 212 -971 213 -955
rect 331 -956 332 -920
rect 597 -971 598 -955
rect 65 -971 66 -957
rect 257 -958 258 -920
rect 261 -958 262 -920
rect 331 -971 332 -957
rect 478 -971 479 -957
rect 548 -958 549 -920
rect 261 -971 262 -959
rect 401 -960 402 -920
rect 506 -960 507 -920
rect 562 -971 563 -959
rect 373 -971 374 -961
rect 401 -971 402 -961
rect 506 -971 507 -961
rect 628 -971 629 -961
rect 548 -971 549 -963
rect 590 -964 591 -920
rect 590 -971 591 -965
rect 625 -966 626 -920
rect 604 -968 605 -920
rect 625 -971 626 -967
rect 604 -971 605 -969
rect 667 -970 668 -920
rect 65 -981 66 -979
rect 229 -981 230 -979
rect 254 -981 255 -979
rect 418 -981 419 -979
rect 422 -981 423 -979
rect 492 -981 493 -979
rect 523 -981 524 -979
rect 527 -981 528 -979
rect 544 -1010 545 -980
rect 569 -981 570 -979
rect 576 -981 577 -979
rect 579 -985 580 -980
rect 607 -1010 608 -980
rect 611 -981 612 -979
rect 649 -1010 650 -980
rect 660 -981 661 -979
rect 670 -1010 671 -980
rect 674 -981 675 -979
rect 72 -983 73 -979
rect 96 -983 97 -979
rect 100 -983 101 -979
rect 250 -1010 251 -982
rect 254 -1010 255 -982
rect 362 -1010 363 -982
rect 373 -983 374 -979
rect 443 -983 444 -979
rect 453 -983 454 -979
rect 499 -983 500 -979
rect 527 -1010 528 -982
rect 534 -983 535 -979
rect 548 -983 549 -979
rect 548 -1010 549 -982
rect 548 -983 549 -979
rect 548 -1010 549 -982
rect 555 -983 556 -979
rect 569 -1010 570 -982
rect 576 -1010 577 -982
rect 590 -983 591 -979
rect 611 -1010 612 -982
rect 618 -983 619 -979
rect 79 -985 80 -979
rect 198 -1010 199 -984
rect 212 -985 213 -979
rect 369 -985 370 -979
rect 380 -985 381 -979
rect 446 -1010 447 -984
rect 464 -985 465 -979
rect 464 -1010 465 -984
rect 464 -985 465 -979
rect 464 -1010 465 -984
rect 471 -985 472 -979
rect 499 -1010 500 -984
rect 590 -1010 591 -984
rect 93 -987 94 -979
rect 100 -1010 101 -986
rect 107 -987 108 -979
rect 128 -987 129 -979
rect 149 -987 150 -979
rect 149 -1010 150 -986
rect 149 -987 150 -979
rect 149 -1010 150 -986
rect 170 -987 171 -979
rect 201 -987 202 -979
rect 264 -1010 265 -986
rect 324 -987 325 -979
rect 331 -987 332 -979
rect 331 -1010 332 -986
rect 331 -987 332 -979
rect 331 -1010 332 -986
rect 352 -987 353 -979
rect 390 -987 391 -979
rect 394 -987 395 -979
rect 422 -1010 423 -986
rect 425 -987 426 -979
rect 436 -987 437 -979
rect 439 -1010 440 -986
rect 506 -987 507 -979
rect 86 -989 87 -979
rect 170 -1010 171 -988
rect 191 -989 192 -979
rect 226 -989 227 -979
rect 240 -989 241 -979
rect 352 -1010 353 -988
rect 369 -1010 370 -988
rect 597 -989 598 -979
rect 117 -991 118 -979
rect 121 -991 122 -979
rect 177 -991 178 -979
rect 240 -1010 241 -990
rect 268 -991 269 -979
rect 373 -1010 374 -990
rect 380 -1010 381 -990
rect 450 -991 451 -979
rect 492 -1010 493 -990
rect 513 -991 514 -979
rect 163 -993 164 -979
rect 177 -1010 178 -992
rect 184 -993 185 -979
rect 268 -1010 269 -992
rect 296 -993 297 -979
rect 394 -1010 395 -992
rect 401 -993 402 -979
rect 401 -1010 402 -992
rect 401 -993 402 -979
rect 401 -1010 402 -992
rect 429 -993 430 -979
rect 646 -1010 647 -992
rect 156 -995 157 -979
rect 163 -1010 164 -994
rect 184 -1010 185 -994
rect 205 -995 206 -979
rect 226 -1010 227 -994
rect 289 -995 290 -979
rect 303 -995 304 -979
rect 436 -1010 437 -994
rect 450 -1010 451 -994
rect 478 -995 479 -979
rect 506 -1010 507 -994
rect 583 -995 584 -979
rect 142 -997 143 -979
rect 156 -1010 157 -996
rect 191 -1010 192 -996
rect 282 -997 283 -979
rect 310 -1010 311 -996
rect 345 -997 346 -979
rect 429 -1010 430 -996
rect 485 -997 486 -979
rect 562 -997 563 -979
rect 583 -1010 584 -996
rect 135 -999 136 -979
rect 142 -1010 143 -998
rect 205 -1010 206 -998
rect 275 -999 276 -979
rect 282 -1010 283 -998
rect 366 -999 367 -979
rect 233 -1001 234 -979
rect 275 -1010 276 -1000
rect 317 -1010 318 -1000
rect 457 -1001 458 -979
rect 219 -1003 220 -979
rect 233 -1010 234 -1002
rect 261 -1003 262 -979
rect 289 -1010 290 -1002
rect 324 -1010 325 -1002
rect 338 -1003 339 -979
rect 345 -1010 346 -1002
rect 408 -1003 409 -979
rect 457 -1010 458 -1002
rect 604 -1003 605 -979
rect 219 -1010 220 -1004
rect 247 -1005 248 -979
rect 338 -1010 339 -1004
rect 359 -1005 360 -979
rect 408 -1010 409 -1004
rect 415 -1005 416 -979
rect 247 -1010 248 -1006
rect 303 -1010 304 -1006
rect 313 -1007 314 -979
rect 415 -1010 416 -1006
rect 359 -1010 360 -1008
rect 387 -1010 388 -1008
rect 100 -1020 101 -1018
rect 100 -1039 101 -1019
rect 100 -1020 101 -1018
rect 100 -1039 101 -1019
rect 114 -1039 115 -1019
rect 173 -1039 174 -1019
rect 198 -1020 199 -1018
rect 348 -1020 349 -1018
rect 352 -1020 353 -1018
rect 460 -1020 461 -1018
rect 478 -1039 479 -1019
rect 506 -1020 507 -1018
rect 548 -1020 549 -1018
rect 548 -1039 549 -1019
rect 548 -1020 549 -1018
rect 548 -1039 549 -1019
rect 562 -1039 563 -1019
rect 576 -1020 577 -1018
rect 583 -1020 584 -1018
rect 583 -1039 584 -1019
rect 583 -1020 584 -1018
rect 583 -1039 584 -1019
rect 590 -1020 591 -1018
rect 590 -1039 591 -1019
rect 590 -1020 591 -1018
rect 590 -1039 591 -1019
rect 604 -1020 605 -1018
rect 611 -1020 612 -1018
rect 128 -1039 129 -1021
rect 163 -1022 164 -1018
rect 198 -1039 199 -1021
rect 219 -1022 220 -1018
rect 229 -1039 230 -1021
rect 247 -1022 248 -1018
rect 268 -1022 269 -1018
rect 366 -1022 367 -1018
rect 373 -1022 374 -1018
rect 429 -1039 430 -1021
rect 436 -1039 437 -1021
rect 450 -1022 451 -1018
rect 457 -1039 458 -1021
rect 464 -1022 465 -1018
rect 485 -1039 486 -1021
rect 492 -1022 493 -1018
rect 499 -1022 500 -1018
rect 527 -1022 528 -1018
rect 569 -1022 570 -1018
rect 569 -1039 570 -1021
rect 569 -1022 570 -1018
rect 569 -1039 570 -1021
rect 135 -1039 136 -1023
rect 149 -1024 150 -1018
rect 163 -1039 164 -1023
rect 177 -1024 178 -1018
rect 191 -1024 192 -1018
rect 247 -1039 248 -1023
rect 275 -1024 276 -1018
rect 317 -1024 318 -1018
rect 366 -1039 367 -1023
rect 380 -1024 381 -1018
rect 387 -1024 388 -1018
rect 387 -1039 388 -1023
rect 387 -1024 388 -1018
rect 387 -1039 388 -1023
rect 394 -1024 395 -1018
rect 474 -1039 475 -1023
rect 149 -1039 150 -1025
rect 156 -1026 157 -1018
rect 177 -1039 178 -1025
rect 219 -1039 220 -1025
rect 226 -1026 227 -1018
rect 268 -1039 269 -1025
rect 289 -1026 290 -1018
rect 359 -1026 360 -1018
rect 373 -1039 374 -1025
rect 415 -1026 416 -1018
rect 418 -1039 419 -1025
rect 422 -1026 423 -1018
rect 142 -1028 143 -1018
rect 156 -1039 157 -1027
rect 184 -1028 185 -1018
rect 191 -1039 192 -1027
rect 205 -1028 206 -1018
rect 306 -1039 307 -1027
rect 317 -1039 318 -1027
rect 338 -1028 339 -1018
rect 394 -1039 395 -1027
rect 401 -1028 402 -1018
rect 408 -1028 409 -1018
rect 408 -1039 409 -1027
rect 408 -1028 409 -1018
rect 408 -1039 409 -1027
rect 422 -1039 423 -1027
rect 443 -1028 444 -1018
rect 124 -1039 125 -1029
rect 142 -1039 143 -1029
rect 170 -1030 171 -1018
rect 205 -1039 206 -1029
rect 215 -1030 216 -1018
rect 233 -1030 234 -1018
rect 240 -1030 241 -1018
rect 243 -1039 244 -1029
rect 254 -1030 255 -1018
rect 289 -1039 290 -1029
rect 296 -1039 297 -1029
rect 310 -1030 311 -1018
rect 439 -1030 440 -1018
rect 443 -1039 444 -1029
rect 170 -1039 171 -1031
rect 282 -1032 283 -1018
rect 299 -1032 300 -1018
rect 303 -1032 304 -1018
rect 310 -1039 311 -1031
rect 324 -1032 325 -1018
rect 215 -1039 216 -1033
rect 254 -1039 255 -1033
rect 233 -1039 234 -1035
rect 264 -1036 265 -1018
rect 261 -1038 262 -1018
rect 264 -1039 265 -1037
rect 100 -1049 101 -1047
rect 107 -1060 108 -1048
rect 128 -1049 129 -1047
rect 194 -1060 195 -1048
rect 198 -1049 199 -1047
rect 212 -1049 213 -1047
rect 219 -1049 220 -1047
rect 226 -1060 227 -1048
rect 247 -1049 248 -1047
rect 303 -1049 304 -1047
rect 366 -1049 367 -1047
rect 380 -1060 381 -1048
rect 383 -1049 384 -1047
rect 387 -1049 388 -1047
rect 394 -1049 395 -1047
rect 404 -1049 405 -1047
rect 408 -1049 409 -1047
rect 411 -1060 412 -1048
rect 415 -1049 416 -1047
rect 429 -1049 430 -1047
rect 443 -1049 444 -1047
rect 453 -1060 454 -1048
rect 457 -1049 458 -1047
rect 457 -1060 458 -1048
rect 457 -1049 458 -1047
rect 457 -1060 458 -1048
rect 471 -1049 472 -1047
rect 485 -1049 486 -1047
rect 541 -1049 542 -1047
rect 548 -1049 549 -1047
rect 562 -1049 563 -1047
rect 562 -1060 563 -1048
rect 562 -1049 563 -1047
rect 562 -1060 563 -1048
rect 579 -1049 580 -1047
rect 583 -1049 584 -1047
rect 142 -1051 143 -1047
rect 173 -1051 174 -1047
rect 180 -1051 181 -1047
rect 233 -1051 234 -1047
rect 254 -1051 255 -1047
rect 275 -1051 276 -1047
rect 278 -1051 279 -1047
rect 296 -1051 297 -1047
rect 299 -1060 300 -1050
rect 310 -1051 311 -1047
rect 376 -1051 377 -1047
rect 422 -1051 423 -1047
rect 429 -1060 430 -1050
rect 436 -1051 437 -1047
rect 443 -1060 444 -1050
rect 478 -1051 479 -1047
rect 569 -1051 570 -1047
rect 583 -1060 584 -1050
rect 142 -1060 143 -1052
rect 156 -1053 157 -1047
rect 163 -1053 164 -1047
rect 184 -1053 185 -1047
rect 191 -1053 192 -1047
rect 198 -1060 199 -1052
rect 205 -1053 206 -1047
rect 233 -1060 234 -1052
rect 268 -1053 269 -1047
rect 282 -1060 283 -1052
rect 285 -1053 286 -1047
rect 317 -1053 318 -1047
rect 579 -1060 580 -1052
rect 590 -1053 591 -1047
rect 149 -1055 150 -1047
rect 163 -1060 164 -1054
rect 289 -1055 290 -1047
rect 296 -1060 297 -1054
rect 135 -1057 136 -1047
rect 149 -1060 150 -1056
rect 114 -1059 115 -1047
rect 135 -1060 136 -1058
rect 100 -1070 101 -1068
rect 107 -1070 108 -1068
rect 149 -1070 150 -1068
rect 159 -1070 160 -1068
rect 163 -1070 164 -1068
rect 170 -1070 171 -1068
rect 198 -1070 199 -1068
rect 205 -1070 206 -1068
rect 215 -1070 216 -1068
rect 233 -1070 234 -1068
rect 380 -1070 381 -1068
rect 394 -1070 395 -1068
rect 429 -1070 430 -1068
rect 439 -1070 440 -1068
rect 446 -1070 447 -1068
rect 457 -1070 458 -1068
rect 576 -1070 577 -1068
rect 583 -1070 584 -1068
rect 219 -1072 220 -1068
rect 226 -1072 227 -1068
<< labels >>
rlabel pdiffusion 3 -10 3 -10 0 cellNo=16
rlabel pdiffusion 10 -10 10 -10 0 cellNo=108
rlabel pdiffusion 17 -10 17 -10 0 cellNo=231
rlabel pdiffusion 24 -10 24 -10 0 cellNo=295
rlabel pdiffusion 115 -10 115 -10 0 cellNo=186
rlabel pdiffusion 122 -10 122 -10 0 feedthrough
rlabel pdiffusion 129 -10 129 -10 0 cellNo=18
rlabel pdiffusion 136 -10 136 -10 0 feedthrough
rlabel pdiffusion 143 -10 143 -10 0 cellNo=139
rlabel pdiffusion 150 -10 150 -10 0 cellNo=352
rlabel pdiffusion 157 -10 157 -10 0 feedthrough
rlabel pdiffusion 164 -10 164 -10 0 cellNo=190
rlabel pdiffusion 171 -10 171 -10 0 cellNo=57
rlabel pdiffusion 178 -10 178 -10 0 feedthrough
rlabel pdiffusion 185 -10 185 -10 0 cellNo=59
rlabel pdiffusion 192 -10 192 -10 0 feedthrough
rlabel pdiffusion 199 -10 199 -10 0 cellNo=319
rlabel pdiffusion 206 -10 206 -10 0 cellNo=5
rlabel pdiffusion 213 -10 213 -10 0 cellNo=172
rlabel pdiffusion 234 -10 234 -10 0 cellNo=9
rlabel pdiffusion 248 -10 248 -10 0 feedthrough
rlabel pdiffusion 297 -10 297 -10 0 feedthrough
rlabel pdiffusion 311 -10 311 -10 0 cellNo=294
rlabel pdiffusion 318 -10 318 -10 0 feedthrough
rlabel pdiffusion 332 -10 332 -10 0 feedthrough
rlabel pdiffusion 339 -10 339 -10 0 cellNo=275
rlabel pdiffusion 346 -10 346 -10 0 cellNo=8
rlabel pdiffusion 353 -10 353 -10 0 feedthrough
rlabel pdiffusion 374 -10 374 -10 0 cellNo=226
rlabel pdiffusion 423 -10 423 -10 0 cellNo=15
rlabel pdiffusion 3 -29 3 -29 0 cellNo=47
rlabel pdiffusion 10 -29 10 -29 0 cellNo=116
rlabel pdiffusion 66 -29 66 -29 0 cellNo=176
rlabel pdiffusion 73 -29 73 -29 0 feedthrough
rlabel pdiffusion 80 -29 80 -29 0 feedthrough
rlabel pdiffusion 87 -29 87 -29 0 cellNo=97
rlabel pdiffusion 94 -29 94 -29 0 cellNo=373
rlabel pdiffusion 101 -29 101 -29 0 feedthrough
rlabel pdiffusion 108 -29 108 -29 0 feedthrough
rlabel pdiffusion 115 -29 115 -29 0 cellNo=3
rlabel pdiffusion 122 -29 122 -29 0 cellNo=130
rlabel pdiffusion 129 -29 129 -29 0 cellNo=114
rlabel pdiffusion 136 -29 136 -29 0 feedthrough
rlabel pdiffusion 143 -29 143 -29 0 feedthrough
rlabel pdiffusion 150 -29 150 -29 0 feedthrough
rlabel pdiffusion 157 -29 157 -29 0 cellNo=161
rlabel pdiffusion 164 -29 164 -29 0 cellNo=258
rlabel pdiffusion 171 -29 171 -29 0 feedthrough
rlabel pdiffusion 178 -29 178 -29 0 feedthrough
rlabel pdiffusion 185 -29 185 -29 0 feedthrough
rlabel pdiffusion 192 -29 192 -29 0 feedthrough
rlabel pdiffusion 199 -29 199 -29 0 cellNo=195
rlabel pdiffusion 206 -29 206 -29 0 cellNo=93
rlabel pdiffusion 213 -29 213 -29 0 feedthrough
rlabel pdiffusion 220 -29 220 -29 0 cellNo=205
rlabel pdiffusion 227 -29 227 -29 0 cellNo=257
rlabel pdiffusion 234 -29 234 -29 0 feedthrough
rlabel pdiffusion 241 -29 241 -29 0 feedthrough
rlabel pdiffusion 248 -29 248 -29 0 cellNo=33
rlabel pdiffusion 255 -29 255 -29 0 feedthrough
rlabel pdiffusion 262 -29 262 -29 0 cellNo=302
rlabel pdiffusion 283 -29 283 -29 0 feedthrough
rlabel pdiffusion 297 -29 297 -29 0 feedthrough
rlabel pdiffusion 304 -29 304 -29 0 feedthrough
rlabel pdiffusion 311 -29 311 -29 0 cellNo=144
rlabel pdiffusion 325 -29 325 -29 0 cellNo=291
rlabel pdiffusion 332 -29 332 -29 0 feedthrough
rlabel pdiffusion 346 -29 346 -29 0 feedthrough
rlabel pdiffusion 353 -29 353 -29 0 feedthrough
rlabel pdiffusion 395 -29 395 -29 0 feedthrough
rlabel pdiffusion 402 -29 402 -29 0 cellNo=29
rlabel pdiffusion 430 -29 430 -29 0 feedthrough
rlabel pdiffusion 437 -29 437 -29 0 feedthrough
rlabel pdiffusion 486 -29 486 -29 0 cellNo=123
rlabel pdiffusion 556 -29 556 -29 0 feedthrough
rlabel pdiffusion 3 -58 3 -58 0 cellNo=42
rlabel pdiffusion 10 -58 10 -58 0 cellNo=92
rlabel pdiffusion 17 -58 17 -58 0 cellNo=253
rlabel pdiffusion 24 -58 24 -58 0 cellNo=312
rlabel pdiffusion 52 -58 52 -58 0 feedthrough
rlabel pdiffusion 59 -58 59 -58 0 cellNo=75
rlabel pdiffusion 66 -58 66 -58 0 feedthrough
rlabel pdiffusion 73 -58 73 -58 0 feedthrough
rlabel pdiffusion 80 -58 80 -58 0 cellNo=14
rlabel pdiffusion 87 -58 87 -58 0 feedthrough
rlabel pdiffusion 94 -58 94 -58 0 feedthrough
rlabel pdiffusion 101 -58 101 -58 0 cellNo=244
rlabel pdiffusion 108 -58 108 -58 0 feedthrough
rlabel pdiffusion 115 -58 115 -58 0 feedthrough
rlabel pdiffusion 122 -58 122 -58 0 feedthrough
rlabel pdiffusion 129 -58 129 -58 0 cellNo=113
rlabel pdiffusion 136 -58 136 -58 0 feedthrough
rlabel pdiffusion 143 -58 143 -58 0 feedthrough
rlabel pdiffusion 150 -58 150 -58 0 feedthrough
rlabel pdiffusion 157 -58 157 -58 0 cellNo=229
rlabel pdiffusion 164 -58 164 -58 0 feedthrough
rlabel pdiffusion 171 -58 171 -58 0 feedthrough
rlabel pdiffusion 178 -58 178 -58 0 feedthrough
rlabel pdiffusion 185 -58 185 -58 0 feedthrough
rlabel pdiffusion 192 -58 192 -58 0 cellNo=7
rlabel pdiffusion 199 -58 199 -58 0 feedthrough
rlabel pdiffusion 206 -58 206 -58 0 feedthrough
rlabel pdiffusion 213 -58 213 -58 0 cellNo=61
rlabel pdiffusion 220 -58 220 -58 0 feedthrough
rlabel pdiffusion 227 -58 227 -58 0 cellNo=67
rlabel pdiffusion 234 -58 234 -58 0 feedthrough
rlabel pdiffusion 241 -58 241 -58 0 cellNo=177
rlabel pdiffusion 248 -58 248 -58 0 feedthrough
rlabel pdiffusion 255 -58 255 -58 0 feedthrough
rlabel pdiffusion 262 -58 262 -58 0 feedthrough
rlabel pdiffusion 269 -58 269 -58 0 feedthrough
rlabel pdiffusion 276 -58 276 -58 0 feedthrough
rlabel pdiffusion 283 -58 283 -58 0 cellNo=189
rlabel pdiffusion 290 -58 290 -58 0 feedthrough
rlabel pdiffusion 297 -58 297 -58 0 feedthrough
rlabel pdiffusion 304 -58 304 -58 0 cellNo=88
rlabel pdiffusion 311 -58 311 -58 0 cellNo=41
rlabel pdiffusion 318 -58 318 -58 0 cellNo=109
rlabel pdiffusion 325 -58 325 -58 0 feedthrough
rlabel pdiffusion 332 -58 332 -58 0 feedthrough
rlabel pdiffusion 339 -58 339 -58 0 feedthrough
rlabel pdiffusion 346 -58 346 -58 0 feedthrough
rlabel pdiffusion 353 -58 353 -58 0 feedthrough
rlabel pdiffusion 360 -58 360 -58 0 feedthrough
rlabel pdiffusion 367 -58 367 -58 0 feedthrough
rlabel pdiffusion 374 -58 374 -58 0 feedthrough
rlabel pdiffusion 381 -58 381 -58 0 cellNo=191
rlabel pdiffusion 388 -58 388 -58 0 feedthrough
rlabel pdiffusion 395 -58 395 -58 0 feedthrough
rlabel pdiffusion 402 -58 402 -58 0 cellNo=132
rlabel pdiffusion 416 -58 416 -58 0 feedthrough
rlabel pdiffusion 444 -58 444 -58 0 feedthrough
rlabel pdiffusion 451 -58 451 -58 0 feedthrough
rlabel pdiffusion 458 -58 458 -58 0 cellNo=95
rlabel pdiffusion 577 -58 577 -58 0 feedthrough
rlabel pdiffusion 31 -97 31 -97 0 feedthrough
rlabel pdiffusion 38 -97 38 -97 0 feedthrough
rlabel pdiffusion 45 -97 45 -97 0 feedthrough
rlabel pdiffusion 52 -97 52 -97 0 feedthrough
rlabel pdiffusion 59 -97 59 -97 0 feedthrough
rlabel pdiffusion 66 -97 66 -97 0 cellNo=293
rlabel pdiffusion 73 -97 73 -97 0 feedthrough
rlabel pdiffusion 80 -97 80 -97 0 cellNo=266
rlabel pdiffusion 87 -97 87 -97 0 feedthrough
rlabel pdiffusion 94 -97 94 -97 0 cellNo=38
rlabel pdiffusion 101 -97 101 -97 0 feedthrough
rlabel pdiffusion 108 -97 108 -97 0 feedthrough
rlabel pdiffusion 115 -97 115 -97 0 feedthrough
rlabel pdiffusion 122 -97 122 -97 0 cellNo=198
rlabel pdiffusion 129 -97 129 -97 0 cellNo=187
rlabel pdiffusion 136 -97 136 -97 0 feedthrough
rlabel pdiffusion 143 -97 143 -97 0 feedthrough
rlabel pdiffusion 150 -97 150 -97 0 cellNo=284
rlabel pdiffusion 157 -97 157 -97 0 cellNo=337
rlabel pdiffusion 164 -97 164 -97 0 feedthrough
rlabel pdiffusion 171 -97 171 -97 0 feedthrough
rlabel pdiffusion 178 -97 178 -97 0 feedthrough
rlabel pdiffusion 185 -97 185 -97 0 feedthrough
rlabel pdiffusion 192 -97 192 -97 0 feedthrough
rlabel pdiffusion 199 -97 199 -97 0 feedthrough
rlabel pdiffusion 206 -97 206 -97 0 feedthrough
rlabel pdiffusion 213 -97 213 -97 0 feedthrough
rlabel pdiffusion 220 -97 220 -97 0 feedthrough
rlabel pdiffusion 227 -97 227 -97 0 feedthrough
rlabel pdiffusion 234 -97 234 -97 0 feedthrough
rlabel pdiffusion 241 -97 241 -97 0 cellNo=222
rlabel pdiffusion 248 -97 248 -97 0 feedthrough
rlabel pdiffusion 255 -97 255 -97 0 cellNo=73
rlabel pdiffusion 262 -97 262 -97 0 feedthrough
rlabel pdiffusion 269 -97 269 -97 0 feedthrough
rlabel pdiffusion 276 -97 276 -97 0 feedthrough
rlabel pdiffusion 283 -97 283 -97 0 cellNo=308
rlabel pdiffusion 290 -97 290 -97 0 feedthrough
rlabel pdiffusion 297 -97 297 -97 0 feedthrough
rlabel pdiffusion 304 -97 304 -97 0 feedthrough
rlabel pdiffusion 311 -97 311 -97 0 cellNo=245
rlabel pdiffusion 318 -97 318 -97 0 cellNo=78
rlabel pdiffusion 325 -97 325 -97 0 feedthrough
rlabel pdiffusion 332 -97 332 -97 0 feedthrough
rlabel pdiffusion 339 -97 339 -97 0 feedthrough
rlabel pdiffusion 346 -97 346 -97 0 feedthrough
rlabel pdiffusion 353 -97 353 -97 0 cellNo=72
rlabel pdiffusion 360 -97 360 -97 0 feedthrough
rlabel pdiffusion 367 -97 367 -97 0 cellNo=24
rlabel pdiffusion 374 -97 374 -97 0 cellNo=98
rlabel pdiffusion 381 -97 381 -97 0 feedthrough
rlabel pdiffusion 388 -97 388 -97 0 feedthrough
rlabel pdiffusion 395 -97 395 -97 0 feedthrough
rlabel pdiffusion 402 -97 402 -97 0 feedthrough
rlabel pdiffusion 409 -97 409 -97 0 feedthrough
rlabel pdiffusion 416 -97 416 -97 0 feedthrough
rlabel pdiffusion 423 -97 423 -97 0 cellNo=62
rlabel pdiffusion 430 -97 430 -97 0 feedthrough
rlabel pdiffusion 437 -97 437 -97 0 feedthrough
rlabel pdiffusion 444 -97 444 -97 0 cellNo=285
rlabel pdiffusion 451 -97 451 -97 0 feedthrough
rlabel pdiffusion 458 -97 458 -97 0 cellNo=35
rlabel pdiffusion 465 -97 465 -97 0 feedthrough
rlabel pdiffusion 472 -97 472 -97 0 feedthrough
rlabel pdiffusion 479 -97 479 -97 0 feedthrough
rlabel pdiffusion 493 -97 493 -97 0 feedthrough
rlabel pdiffusion 521 -97 521 -97 0 cellNo=80
rlabel pdiffusion 528 -97 528 -97 0 cellNo=60
rlabel pdiffusion 577 -97 577 -97 0 feedthrough
rlabel pdiffusion 591 -97 591 -97 0 feedthrough
rlabel pdiffusion 3 -148 3 -148 0 cellNo=169
rlabel pdiffusion 10 -148 10 -148 0 feedthrough
rlabel pdiffusion 17 -148 17 -148 0 feedthrough
rlabel pdiffusion 24 -148 24 -148 0 cellNo=334
rlabel pdiffusion 31 -148 31 -148 0 feedthrough
rlabel pdiffusion 38 -148 38 -148 0 feedthrough
rlabel pdiffusion 45 -148 45 -148 0 feedthrough
rlabel pdiffusion 52 -148 52 -148 0 feedthrough
rlabel pdiffusion 59 -148 59 -148 0 feedthrough
rlabel pdiffusion 66 -148 66 -148 0 feedthrough
rlabel pdiffusion 73 -148 73 -148 0 cellNo=36
rlabel pdiffusion 80 -148 80 -148 0 cellNo=43
rlabel pdiffusion 87 -148 87 -148 0 cellNo=70
rlabel pdiffusion 94 -148 94 -148 0 cellNo=194
rlabel pdiffusion 101 -148 101 -148 0 feedthrough
rlabel pdiffusion 108 -148 108 -148 0 feedthrough
rlabel pdiffusion 115 -148 115 -148 0 feedthrough
rlabel pdiffusion 122 -148 122 -148 0 feedthrough
rlabel pdiffusion 129 -148 129 -148 0 feedthrough
rlabel pdiffusion 136 -148 136 -148 0 feedthrough
rlabel pdiffusion 143 -148 143 -148 0 feedthrough
rlabel pdiffusion 150 -148 150 -148 0 feedthrough
rlabel pdiffusion 157 -148 157 -148 0 feedthrough
rlabel pdiffusion 164 -148 164 -148 0 cellNo=289
rlabel pdiffusion 171 -148 171 -148 0 cellNo=282
rlabel pdiffusion 178 -148 178 -148 0 feedthrough
rlabel pdiffusion 185 -148 185 -148 0 feedthrough
rlabel pdiffusion 192 -148 192 -148 0 feedthrough
rlabel pdiffusion 199 -148 199 -148 0 feedthrough
rlabel pdiffusion 206 -148 206 -148 0 feedthrough
rlabel pdiffusion 213 -148 213 -148 0 feedthrough
rlabel pdiffusion 220 -148 220 -148 0 cellNo=214
rlabel pdiffusion 227 -148 227 -148 0 feedthrough
rlabel pdiffusion 234 -148 234 -148 0 feedthrough
rlabel pdiffusion 241 -148 241 -148 0 feedthrough
rlabel pdiffusion 248 -148 248 -148 0 feedthrough
rlabel pdiffusion 255 -148 255 -148 0 cellNo=6
rlabel pdiffusion 262 -148 262 -148 0 cellNo=211
rlabel pdiffusion 269 -148 269 -148 0 feedthrough
rlabel pdiffusion 276 -148 276 -148 0 cellNo=350
rlabel pdiffusion 283 -148 283 -148 0 feedthrough
rlabel pdiffusion 290 -148 290 -148 0 cellNo=311
rlabel pdiffusion 297 -148 297 -148 0 feedthrough
rlabel pdiffusion 304 -148 304 -148 0 feedthrough
rlabel pdiffusion 311 -148 311 -148 0 cellNo=126
rlabel pdiffusion 318 -148 318 -148 0 cellNo=252
rlabel pdiffusion 325 -148 325 -148 0 feedthrough
rlabel pdiffusion 332 -148 332 -148 0 feedthrough
rlabel pdiffusion 339 -148 339 -148 0 feedthrough
rlabel pdiffusion 346 -148 346 -148 0 feedthrough
rlabel pdiffusion 353 -148 353 -148 0 feedthrough
rlabel pdiffusion 360 -148 360 -148 0 feedthrough
rlabel pdiffusion 367 -148 367 -148 0 feedthrough
rlabel pdiffusion 374 -148 374 -148 0 feedthrough
rlabel pdiffusion 381 -148 381 -148 0 feedthrough
rlabel pdiffusion 388 -148 388 -148 0 feedthrough
rlabel pdiffusion 395 -148 395 -148 0 feedthrough
rlabel pdiffusion 402 -148 402 -148 0 feedthrough
rlabel pdiffusion 409 -148 409 -148 0 feedthrough
rlabel pdiffusion 416 -148 416 -148 0 cellNo=117
rlabel pdiffusion 423 -148 423 -148 0 feedthrough
rlabel pdiffusion 430 -148 430 -148 0 feedthrough
rlabel pdiffusion 437 -148 437 -148 0 feedthrough
rlabel pdiffusion 444 -148 444 -148 0 feedthrough
rlabel pdiffusion 451 -148 451 -148 0 feedthrough
rlabel pdiffusion 458 -148 458 -148 0 feedthrough
rlabel pdiffusion 465 -148 465 -148 0 feedthrough
rlabel pdiffusion 472 -148 472 -148 0 cellNo=254
rlabel pdiffusion 479 -148 479 -148 0 feedthrough
rlabel pdiffusion 486 -148 486 -148 0 feedthrough
rlabel pdiffusion 493 -148 493 -148 0 feedthrough
rlabel pdiffusion 500 -148 500 -148 0 cellNo=255
rlabel pdiffusion 507 -148 507 -148 0 feedthrough
rlabel pdiffusion 514 -148 514 -148 0 feedthrough
rlabel pdiffusion 521 -148 521 -148 0 feedthrough
rlabel pdiffusion 528 -148 528 -148 0 feedthrough
rlabel pdiffusion 535 -148 535 -148 0 feedthrough
rlabel pdiffusion 542 -148 542 -148 0 feedthrough
rlabel pdiffusion 549 -148 549 -148 0 feedthrough
rlabel pdiffusion 556 -148 556 -148 0 feedthrough
rlabel pdiffusion 563 -148 563 -148 0 feedthrough
rlabel pdiffusion 570 -148 570 -148 0 feedthrough
rlabel pdiffusion 577 -148 577 -148 0 feedthrough
rlabel pdiffusion 584 -148 584 -148 0 cellNo=376
rlabel pdiffusion 591 -148 591 -148 0 feedthrough
rlabel pdiffusion 598 -148 598 -148 0 feedthrough
rlabel pdiffusion 605 -148 605 -148 0 feedthrough
rlabel pdiffusion 612 -148 612 -148 0 feedthrough
rlabel pdiffusion 619 -148 619 -148 0 feedthrough
rlabel pdiffusion 626 -148 626 -148 0 cellNo=23
rlabel pdiffusion 3 -209 3 -209 0 cellNo=102
rlabel pdiffusion 10 -209 10 -209 0 cellNo=118
rlabel pdiffusion 17 -209 17 -209 0 feedthrough
rlabel pdiffusion 24 -209 24 -209 0 feedthrough
rlabel pdiffusion 31 -209 31 -209 0 feedthrough
rlabel pdiffusion 38 -209 38 -209 0 feedthrough
rlabel pdiffusion 45 -209 45 -209 0 feedthrough
rlabel pdiffusion 52 -209 52 -209 0 feedthrough
rlabel pdiffusion 59 -209 59 -209 0 feedthrough
rlabel pdiffusion 66 -209 66 -209 0 feedthrough
rlabel pdiffusion 73 -209 73 -209 0 cellNo=101
rlabel pdiffusion 80 -209 80 -209 0 feedthrough
rlabel pdiffusion 87 -209 87 -209 0 feedthrough
rlabel pdiffusion 94 -209 94 -209 0 cellNo=84
rlabel pdiffusion 101 -209 101 -209 0 cellNo=119
rlabel pdiffusion 108 -209 108 -209 0 feedthrough
rlabel pdiffusion 115 -209 115 -209 0 feedthrough
rlabel pdiffusion 122 -209 122 -209 0 feedthrough
rlabel pdiffusion 129 -209 129 -209 0 feedthrough
rlabel pdiffusion 136 -209 136 -209 0 cellNo=166
rlabel pdiffusion 143 -209 143 -209 0 feedthrough
rlabel pdiffusion 150 -209 150 -209 0 feedthrough
rlabel pdiffusion 157 -209 157 -209 0 feedthrough
rlabel pdiffusion 164 -209 164 -209 0 feedthrough
rlabel pdiffusion 171 -209 171 -209 0 feedthrough
rlabel pdiffusion 178 -209 178 -209 0 cellNo=283
rlabel pdiffusion 185 -209 185 -209 0 feedthrough
rlabel pdiffusion 192 -209 192 -209 0 feedthrough
rlabel pdiffusion 199 -209 199 -209 0 feedthrough
rlabel pdiffusion 206 -209 206 -209 0 cellNo=77
rlabel pdiffusion 213 -209 213 -209 0 cellNo=242
rlabel pdiffusion 220 -209 220 -209 0 feedthrough
rlabel pdiffusion 227 -209 227 -209 0 feedthrough
rlabel pdiffusion 234 -209 234 -209 0 feedthrough
rlabel pdiffusion 241 -209 241 -209 0 feedthrough
rlabel pdiffusion 248 -209 248 -209 0 feedthrough
rlabel pdiffusion 255 -209 255 -209 0 feedthrough
rlabel pdiffusion 262 -209 262 -209 0 feedthrough
rlabel pdiffusion 269 -209 269 -209 0 feedthrough
rlabel pdiffusion 276 -209 276 -209 0 cellNo=55
rlabel pdiffusion 283 -209 283 -209 0 feedthrough
rlabel pdiffusion 290 -209 290 -209 0 feedthrough
rlabel pdiffusion 297 -209 297 -209 0 cellNo=356
rlabel pdiffusion 304 -209 304 -209 0 cellNo=197
rlabel pdiffusion 311 -209 311 -209 0 feedthrough
rlabel pdiffusion 318 -209 318 -209 0 cellNo=278
rlabel pdiffusion 325 -209 325 -209 0 cellNo=120
rlabel pdiffusion 332 -209 332 -209 0 cellNo=184
rlabel pdiffusion 339 -209 339 -209 0 cellNo=288
rlabel pdiffusion 346 -209 346 -209 0 feedthrough
rlabel pdiffusion 353 -209 353 -209 0 feedthrough
rlabel pdiffusion 360 -209 360 -209 0 feedthrough
rlabel pdiffusion 367 -209 367 -209 0 cellNo=149
rlabel pdiffusion 374 -209 374 -209 0 feedthrough
rlabel pdiffusion 381 -209 381 -209 0 feedthrough
rlabel pdiffusion 388 -209 388 -209 0 cellNo=135
rlabel pdiffusion 395 -209 395 -209 0 feedthrough
rlabel pdiffusion 402 -209 402 -209 0 feedthrough
rlabel pdiffusion 409 -209 409 -209 0 feedthrough
rlabel pdiffusion 416 -209 416 -209 0 feedthrough
rlabel pdiffusion 423 -209 423 -209 0 feedthrough
rlabel pdiffusion 430 -209 430 -209 0 feedthrough
rlabel pdiffusion 437 -209 437 -209 0 feedthrough
rlabel pdiffusion 444 -209 444 -209 0 cellNo=175
rlabel pdiffusion 451 -209 451 -209 0 feedthrough
rlabel pdiffusion 458 -209 458 -209 0 feedthrough
rlabel pdiffusion 465 -209 465 -209 0 feedthrough
rlabel pdiffusion 472 -209 472 -209 0 feedthrough
rlabel pdiffusion 479 -209 479 -209 0 feedthrough
rlabel pdiffusion 486 -209 486 -209 0 cellNo=310
rlabel pdiffusion 493 -209 493 -209 0 feedthrough
rlabel pdiffusion 500 -209 500 -209 0 feedthrough
rlabel pdiffusion 507 -209 507 -209 0 feedthrough
rlabel pdiffusion 514 -209 514 -209 0 feedthrough
rlabel pdiffusion 521 -209 521 -209 0 feedthrough
rlabel pdiffusion 528 -209 528 -209 0 feedthrough
rlabel pdiffusion 535 -209 535 -209 0 feedthrough
rlabel pdiffusion 542 -209 542 -209 0 feedthrough
rlabel pdiffusion 549 -209 549 -209 0 feedthrough
rlabel pdiffusion 556 -209 556 -209 0 feedthrough
rlabel pdiffusion 563 -209 563 -209 0 feedthrough
rlabel pdiffusion 570 -209 570 -209 0 feedthrough
rlabel pdiffusion 577 -209 577 -209 0 feedthrough
rlabel pdiffusion 584 -209 584 -209 0 feedthrough
rlabel pdiffusion 591 -209 591 -209 0 feedthrough
rlabel pdiffusion 598 -209 598 -209 0 feedthrough
rlabel pdiffusion 605 -209 605 -209 0 feedthrough
rlabel pdiffusion 612 -209 612 -209 0 feedthrough
rlabel pdiffusion 619 -209 619 -209 0 feedthrough
rlabel pdiffusion 626 -209 626 -209 0 feedthrough
rlabel pdiffusion 633 -209 633 -209 0 feedthrough
rlabel pdiffusion 640 -209 640 -209 0 feedthrough
rlabel pdiffusion 647 -209 647 -209 0 feedthrough
rlabel pdiffusion 654 -209 654 -209 0 feedthrough
rlabel pdiffusion 661 -209 661 -209 0 feedthrough
rlabel pdiffusion 668 -209 668 -209 0 feedthrough
rlabel pdiffusion 675 -209 675 -209 0 feedthrough
rlabel pdiffusion 3 -274 3 -274 0 feedthrough
rlabel pdiffusion 10 -274 10 -274 0 cellNo=203
rlabel pdiffusion 17 -274 17 -274 0 feedthrough
rlabel pdiffusion 24 -274 24 -274 0 feedthrough
rlabel pdiffusion 31 -274 31 -274 0 cellNo=147
rlabel pdiffusion 38 -274 38 -274 0 feedthrough
rlabel pdiffusion 45 -274 45 -274 0 feedthrough
rlabel pdiffusion 52 -274 52 -274 0 cellNo=152
rlabel pdiffusion 59 -274 59 -274 0 feedthrough
rlabel pdiffusion 66 -274 66 -274 0 feedthrough
rlabel pdiffusion 73 -274 73 -274 0 feedthrough
rlabel pdiffusion 80 -274 80 -274 0 cellNo=112
rlabel pdiffusion 87 -274 87 -274 0 feedthrough
rlabel pdiffusion 94 -274 94 -274 0 feedthrough
rlabel pdiffusion 101 -274 101 -274 0 cellNo=264
rlabel pdiffusion 108 -274 108 -274 0 cellNo=287
rlabel pdiffusion 115 -274 115 -274 0 cellNo=301
rlabel pdiffusion 122 -274 122 -274 0 feedthrough
rlabel pdiffusion 129 -274 129 -274 0 feedthrough
rlabel pdiffusion 136 -274 136 -274 0 feedthrough
rlabel pdiffusion 143 -274 143 -274 0 feedthrough
rlabel pdiffusion 150 -274 150 -274 0 cellNo=140
rlabel pdiffusion 157 -274 157 -274 0 feedthrough
rlabel pdiffusion 164 -274 164 -274 0 feedthrough
rlabel pdiffusion 171 -274 171 -274 0 feedthrough
rlabel pdiffusion 178 -274 178 -274 0 feedthrough
rlabel pdiffusion 185 -274 185 -274 0 feedthrough
rlabel pdiffusion 192 -274 192 -274 0 feedthrough
rlabel pdiffusion 199 -274 199 -274 0 feedthrough
rlabel pdiffusion 206 -274 206 -274 0 feedthrough
rlabel pdiffusion 213 -274 213 -274 0 feedthrough
rlabel pdiffusion 220 -274 220 -274 0 feedthrough
rlabel pdiffusion 227 -274 227 -274 0 feedthrough
rlabel pdiffusion 234 -274 234 -274 0 feedthrough
rlabel pdiffusion 241 -274 241 -274 0 cellNo=32
rlabel pdiffusion 248 -274 248 -274 0 cellNo=370
rlabel pdiffusion 255 -274 255 -274 0 feedthrough
rlabel pdiffusion 262 -274 262 -274 0 cellNo=268
rlabel pdiffusion 269 -274 269 -274 0 feedthrough
rlabel pdiffusion 276 -274 276 -274 0 cellNo=200
rlabel pdiffusion 283 -274 283 -274 0 feedthrough
rlabel pdiffusion 290 -274 290 -274 0 cellNo=199
rlabel pdiffusion 297 -274 297 -274 0 cellNo=246
rlabel pdiffusion 304 -274 304 -274 0 feedthrough
rlabel pdiffusion 311 -274 311 -274 0 cellNo=188
rlabel pdiffusion 318 -274 318 -274 0 feedthrough
rlabel pdiffusion 325 -274 325 -274 0 feedthrough
rlabel pdiffusion 332 -274 332 -274 0 feedthrough
rlabel pdiffusion 339 -274 339 -274 0 feedthrough
rlabel pdiffusion 346 -274 346 -274 0 feedthrough
rlabel pdiffusion 353 -274 353 -274 0 feedthrough
rlabel pdiffusion 360 -274 360 -274 0 feedthrough
rlabel pdiffusion 367 -274 367 -274 0 cellNo=383
rlabel pdiffusion 374 -274 374 -274 0 feedthrough
rlabel pdiffusion 381 -274 381 -274 0 cellNo=82
rlabel pdiffusion 388 -274 388 -274 0 feedthrough
rlabel pdiffusion 395 -274 395 -274 0 feedthrough
rlabel pdiffusion 402 -274 402 -274 0 feedthrough
rlabel pdiffusion 409 -274 409 -274 0 feedthrough
rlabel pdiffusion 416 -274 416 -274 0 feedthrough
rlabel pdiffusion 423 -274 423 -274 0 feedthrough
rlabel pdiffusion 430 -274 430 -274 0 feedthrough
rlabel pdiffusion 437 -274 437 -274 0 feedthrough
rlabel pdiffusion 444 -274 444 -274 0 feedthrough
rlabel pdiffusion 451 -274 451 -274 0 feedthrough
rlabel pdiffusion 458 -274 458 -274 0 feedthrough
rlabel pdiffusion 465 -274 465 -274 0 cellNo=83
rlabel pdiffusion 472 -274 472 -274 0 feedthrough
rlabel pdiffusion 479 -274 479 -274 0 feedthrough
rlabel pdiffusion 486 -274 486 -274 0 feedthrough
rlabel pdiffusion 493 -274 493 -274 0 feedthrough
rlabel pdiffusion 500 -274 500 -274 0 feedthrough
rlabel pdiffusion 507 -274 507 -274 0 feedthrough
rlabel pdiffusion 514 -274 514 -274 0 feedthrough
rlabel pdiffusion 521 -274 521 -274 0 feedthrough
rlabel pdiffusion 528 -274 528 -274 0 feedthrough
rlabel pdiffusion 535 -274 535 -274 0 feedthrough
rlabel pdiffusion 542 -274 542 -274 0 feedthrough
rlabel pdiffusion 549 -274 549 -274 0 feedthrough
rlabel pdiffusion 556 -274 556 -274 0 feedthrough
rlabel pdiffusion 563 -274 563 -274 0 feedthrough
rlabel pdiffusion 570 -274 570 -274 0 feedthrough
rlabel pdiffusion 577 -274 577 -274 0 feedthrough
rlabel pdiffusion 584 -274 584 -274 0 feedthrough
rlabel pdiffusion 591 -274 591 -274 0 feedthrough
rlabel pdiffusion 598 -274 598 -274 0 feedthrough
rlabel pdiffusion 605 -274 605 -274 0 feedthrough
rlabel pdiffusion 612 -274 612 -274 0 feedthrough
rlabel pdiffusion 619 -274 619 -274 0 feedthrough
rlabel pdiffusion 626 -274 626 -274 0 feedthrough
rlabel pdiffusion 633 -274 633 -274 0 feedthrough
rlabel pdiffusion 640 -274 640 -274 0 feedthrough
rlabel pdiffusion 647 -274 647 -274 0 feedthrough
rlabel pdiffusion 654 -274 654 -274 0 feedthrough
rlabel pdiffusion 661 -274 661 -274 0 feedthrough
rlabel pdiffusion 668 -274 668 -274 0 feedthrough
rlabel pdiffusion 675 -274 675 -274 0 feedthrough
rlabel pdiffusion 682 -274 682 -274 0 feedthrough
rlabel pdiffusion 689 -274 689 -274 0 feedthrough
rlabel pdiffusion 696 -274 696 -274 0 feedthrough
rlabel pdiffusion 703 -274 703 -274 0 feedthrough
rlabel pdiffusion 710 -274 710 -274 0 cellNo=223
rlabel pdiffusion 717 -274 717 -274 0 feedthrough
rlabel pdiffusion 724 -274 724 -274 0 feedthrough
rlabel pdiffusion 731 -274 731 -274 0 cellNo=121
rlabel pdiffusion 3 -341 3 -341 0 cellNo=209
rlabel pdiffusion 10 -341 10 -341 0 cellNo=235
rlabel pdiffusion 17 -341 17 -341 0 feedthrough
rlabel pdiffusion 24 -341 24 -341 0 cellNo=31
rlabel pdiffusion 31 -341 31 -341 0 feedthrough
rlabel pdiffusion 38 -341 38 -341 0 feedthrough
rlabel pdiffusion 45 -341 45 -341 0 cellNo=11
rlabel pdiffusion 52 -341 52 -341 0 cellNo=106
rlabel pdiffusion 59 -341 59 -341 0 cellNo=94
rlabel pdiffusion 66 -341 66 -341 0 feedthrough
rlabel pdiffusion 73 -341 73 -341 0 feedthrough
rlabel pdiffusion 80 -341 80 -341 0 feedthrough
rlabel pdiffusion 87 -341 87 -341 0 feedthrough
rlabel pdiffusion 94 -341 94 -341 0 feedthrough
rlabel pdiffusion 101 -341 101 -341 0 feedthrough
rlabel pdiffusion 108 -341 108 -341 0 cellNo=323
rlabel pdiffusion 115 -341 115 -341 0 feedthrough
rlabel pdiffusion 122 -341 122 -341 0 feedthrough
rlabel pdiffusion 129 -341 129 -341 0 feedthrough
rlabel pdiffusion 136 -341 136 -341 0 feedthrough
rlabel pdiffusion 143 -341 143 -341 0 feedthrough
rlabel pdiffusion 150 -341 150 -341 0 feedthrough
rlabel pdiffusion 157 -341 157 -341 0 feedthrough
rlabel pdiffusion 164 -341 164 -341 0 cellNo=170
rlabel pdiffusion 171 -341 171 -341 0 feedthrough
rlabel pdiffusion 178 -341 178 -341 0 feedthrough
rlabel pdiffusion 185 -341 185 -341 0 cellNo=233
rlabel pdiffusion 192 -341 192 -341 0 feedthrough
rlabel pdiffusion 199 -341 199 -341 0 feedthrough
rlabel pdiffusion 206 -341 206 -341 0 feedthrough
rlabel pdiffusion 213 -341 213 -341 0 feedthrough
rlabel pdiffusion 220 -341 220 -341 0 feedthrough
rlabel pdiffusion 227 -341 227 -341 0 cellNo=90
rlabel pdiffusion 234 -341 234 -341 0 feedthrough
rlabel pdiffusion 241 -341 241 -341 0 feedthrough
rlabel pdiffusion 248 -341 248 -341 0 feedthrough
rlabel pdiffusion 255 -341 255 -341 0 cellNo=74
rlabel pdiffusion 262 -341 262 -341 0 feedthrough
rlabel pdiffusion 269 -341 269 -341 0 feedthrough
rlabel pdiffusion 276 -341 276 -341 0 cellNo=34
rlabel pdiffusion 283 -341 283 -341 0 cellNo=201
rlabel pdiffusion 290 -341 290 -341 0 feedthrough
rlabel pdiffusion 297 -341 297 -341 0 cellNo=384
rlabel pdiffusion 304 -341 304 -341 0 feedthrough
rlabel pdiffusion 311 -341 311 -341 0 feedthrough
rlabel pdiffusion 318 -341 318 -341 0 feedthrough
rlabel pdiffusion 325 -341 325 -341 0 cellNo=25
rlabel pdiffusion 332 -341 332 -341 0 feedthrough
rlabel pdiffusion 339 -341 339 -341 0 feedthrough
rlabel pdiffusion 346 -341 346 -341 0 cellNo=304
rlabel pdiffusion 353 -341 353 -341 0 feedthrough
rlabel pdiffusion 360 -341 360 -341 0 cellNo=158
rlabel pdiffusion 367 -341 367 -341 0 cellNo=146
rlabel pdiffusion 374 -341 374 -341 0 feedthrough
rlabel pdiffusion 381 -341 381 -341 0 feedthrough
rlabel pdiffusion 388 -341 388 -341 0 feedthrough
rlabel pdiffusion 395 -341 395 -341 0 feedthrough
rlabel pdiffusion 402 -341 402 -341 0 cellNo=110
rlabel pdiffusion 409 -341 409 -341 0 feedthrough
rlabel pdiffusion 416 -341 416 -341 0 feedthrough
rlabel pdiffusion 423 -341 423 -341 0 feedthrough
rlabel pdiffusion 430 -341 430 -341 0 cellNo=332
rlabel pdiffusion 437 -341 437 -341 0 feedthrough
rlabel pdiffusion 444 -341 444 -341 0 feedthrough
rlabel pdiffusion 451 -341 451 -341 0 feedthrough
rlabel pdiffusion 458 -341 458 -341 0 feedthrough
rlabel pdiffusion 465 -341 465 -341 0 feedthrough
rlabel pdiffusion 472 -341 472 -341 0 feedthrough
rlabel pdiffusion 479 -341 479 -341 0 feedthrough
rlabel pdiffusion 486 -341 486 -341 0 feedthrough
rlabel pdiffusion 493 -341 493 -341 0 feedthrough
rlabel pdiffusion 500 -341 500 -341 0 feedthrough
rlabel pdiffusion 507 -341 507 -341 0 feedthrough
rlabel pdiffusion 514 -341 514 -341 0 feedthrough
rlabel pdiffusion 521 -341 521 -341 0 feedthrough
rlabel pdiffusion 528 -341 528 -341 0 feedthrough
rlabel pdiffusion 535 -341 535 -341 0 feedthrough
rlabel pdiffusion 542 -341 542 -341 0 feedthrough
rlabel pdiffusion 549 -341 549 -341 0 feedthrough
rlabel pdiffusion 556 -341 556 -341 0 feedthrough
rlabel pdiffusion 563 -341 563 -341 0 feedthrough
rlabel pdiffusion 570 -341 570 -341 0 feedthrough
rlabel pdiffusion 577 -341 577 -341 0 feedthrough
rlabel pdiffusion 584 -341 584 -341 0 feedthrough
rlabel pdiffusion 591 -341 591 -341 0 feedthrough
rlabel pdiffusion 598 -341 598 -341 0 feedthrough
rlabel pdiffusion 605 -341 605 -341 0 feedthrough
rlabel pdiffusion 612 -341 612 -341 0 feedthrough
rlabel pdiffusion 619 -341 619 -341 0 feedthrough
rlabel pdiffusion 626 -341 626 -341 0 feedthrough
rlabel pdiffusion 633 -341 633 -341 0 feedthrough
rlabel pdiffusion 640 -341 640 -341 0 feedthrough
rlabel pdiffusion 647 -341 647 -341 0 feedthrough
rlabel pdiffusion 654 -341 654 -341 0 feedthrough
rlabel pdiffusion 661 -341 661 -341 0 feedthrough
rlabel pdiffusion 668 -341 668 -341 0 feedthrough
rlabel pdiffusion 675 -341 675 -341 0 feedthrough
rlabel pdiffusion 682 -341 682 -341 0 feedthrough
rlabel pdiffusion 689 -341 689 -341 0 feedthrough
rlabel pdiffusion 696 -341 696 -341 0 feedthrough
rlabel pdiffusion 703 -341 703 -341 0 feedthrough
rlabel pdiffusion 710 -341 710 -341 0 feedthrough
rlabel pdiffusion 717 -341 717 -341 0 feedthrough
rlabel pdiffusion 724 -341 724 -341 0 feedthrough
rlabel pdiffusion 731 -341 731 -341 0 feedthrough
rlabel pdiffusion 738 -341 738 -341 0 feedthrough
rlabel pdiffusion 3 -420 3 -420 0 cellNo=286
rlabel pdiffusion 10 -420 10 -420 0 cellNo=230
rlabel pdiffusion 17 -420 17 -420 0 feedthrough
rlabel pdiffusion 24 -420 24 -420 0 feedthrough
rlabel pdiffusion 31 -420 31 -420 0 feedthrough
rlabel pdiffusion 38 -420 38 -420 0 feedthrough
rlabel pdiffusion 45 -420 45 -420 0 feedthrough
rlabel pdiffusion 52 -420 52 -420 0 feedthrough
rlabel pdiffusion 59 -420 59 -420 0 cellNo=180
rlabel pdiffusion 66 -420 66 -420 0 feedthrough
rlabel pdiffusion 73 -420 73 -420 0 feedthrough
rlabel pdiffusion 80 -420 80 -420 0 feedthrough
rlabel pdiffusion 87 -420 87 -420 0 feedthrough
rlabel pdiffusion 94 -420 94 -420 0 feedthrough
rlabel pdiffusion 101 -420 101 -420 0 feedthrough
rlabel pdiffusion 108 -420 108 -420 0 cellNo=193
rlabel pdiffusion 115 -420 115 -420 0 feedthrough
rlabel pdiffusion 122 -420 122 -420 0 cellNo=27
rlabel pdiffusion 129 -420 129 -420 0 feedthrough
rlabel pdiffusion 136 -420 136 -420 0 feedthrough
rlabel pdiffusion 143 -420 143 -420 0 feedthrough
rlabel pdiffusion 150 -420 150 -420 0 feedthrough
rlabel pdiffusion 157 -420 157 -420 0 feedthrough
rlabel pdiffusion 164 -420 164 -420 0 feedthrough
rlabel pdiffusion 171 -420 171 -420 0 feedthrough
rlabel pdiffusion 178 -420 178 -420 0 feedthrough
rlabel pdiffusion 185 -420 185 -420 0 feedthrough
rlabel pdiffusion 192 -420 192 -420 0 feedthrough
rlabel pdiffusion 199 -420 199 -420 0 feedthrough
rlabel pdiffusion 206 -420 206 -420 0 feedthrough
rlabel pdiffusion 213 -420 213 -420 0 feedthrough
rlabel pdiffusion 220 -420 220 -420 0 cellNo=213
rlabel pdiffusion 227 -420 227 -420 0 feedthrough
rlabel pdiffusion 234 -420 234 -420 0 feedthrough
rlabel pdiffusion 241 -420 241 -420 0 feedthrough
rlabel pdiffusion 248 -420 248 -420 0 feedthrough
rlabel pdiffusion 255 -420 255 -420 0 feedthrough
rlabel pdiffusion 262 -420 262 -420 0 feedthrough
rlabel pdiffusion 269 -420 269 -420 0 feedthrough
rlabel pdiffusion 276 -420 276 -420 0 feedthrough
rlabel pdiffusion 283 -420 283 -420 0 feedthrough
rlabel pdiffusion 290 -420 290 -420 0 cellNo=56
rlabel pdiffusion 297 -420 297 -420 0 feedthrough
rlabel pdiffusion 304 -420 304 -420 0 feedthrough
rlabel pdiffusion 311 -420 311 -420 0 feedthrough
rlabel pdiffusion 318 -420 318 -420 0 feedthrough
rlabel pdiffusion 325 -420 325 -420 0 feedthrough
rlabel pdiffusion 332 -420 332 -420 0 cellNo=171
rlabel pdiffusion 339 -420 339 -420 0 cellNo=228
rlabel pdiffusion 346 -420 346 -420 0 cellNo=51
rlabel pdiffusion 353 -420 353 -420 0 feedthrough
rlabel pdiffusion 360 -420 360 -420 0 feedthrough
rlabel pdiffusion 367 -420 367 -420 0 feedthrough
rlabel pdiffusion 374 -420 374 -420 0 cellNo=164
rlabel pdiffusion 381 -420 381 -420 0 cellNo=10
rlabel pdiffusion 388 -420 388 -420 0 feedthrough
rlabel pdiffusion 395 -420 395 -420 0 cellNo=137
rlabel pdiffusion 402 -420 402 -420 0 cellNo=168
rlabel pdiffusion 409 -420 409 -420 0 feedthrough
rlabel pdiffusion 416 -420 416 -420 0 cellNo=162
rlabel pdiffusion 423 -420 423 -420 0 feedthrough
rlabel pdiffusion 430 -420 430 -420 0 cellNo=17
rlabel pdiffusion 437 -420 437 -420 0 feedthrough
rlabel pdiffusion 444 -420 444 -420 0 feedthrough
rlabel pdiffusion 451 -420 451 -420 0 feedthrough
rlabel pdiffusion 458 -420 458 -420 0 feedthrough
rlabel pdiffusion 465 -420 465 -420 0 feedthrough
rlabel pdiffusion 472 -420 472 -420 0 cellNo=19
rlabel pdiffusion 479 -420 479 -420 0 feedthrough
rlabel pdiffusion 486 -420 486 -420 0 feedthrough
rlabel pdiffusion 493 -420 493 -420 0 feedthrough
rlabel pdiffusion 500 -420 500 -420 0 feedthrough
rlabel pdiffusion 507 -420 507 -420 0 cellNo=178
rlabel pdiffusion 514 -420 514 -420 0 feedthrough
rlabel pdiffusion 521 -420 521 -420 0 cellNo=141
rlabel pdiffusion 528 -420 528 -420 0 feedthrough
rlabel pdiffusion 535 -420 535 -420 0 feedthrough
rlabel pdiffusion 542 -420 542 -420 0 feedthrough
rlabel pdiffusion 549 -420 549 -420 0 feedthrough
rlabel pdiffusion 556 -420 556 -420 0 cellNo=127
rlabel pdiffusion 563 -420 563 -420 0 feedthrough
rlabel pdiffusion 570 -420 570 -420 0 feedthrough
rlabel pdiffusion 577 -420 577 -420 0 feedthrough
rlabel pdiffusion 584 -420 584 -420 0 feedthrough
rlabel pdiffusion 591 -420 591 -420 0 feedthrough
rlabel pdiffusion 598 -420 598 -420 0 feedthrough
rlabel pdiffusion 605 -420 605 -420 0 feedthrough
rlabel pdiffusion 612 -420 612 -420 0 feedthrough
rlabel pdiffusion 619 -420 619 -420 0 feedthrough
rlabel pdiffusion 626 -420 626 -420 0 feedthrough
rlabel pdiffusion 633 -420 633 -420 0 feedthrough
rlabel pdiffusion 640 -420 640 -420 0 feedthrough
rlabel pdiffusion 647 -420 647 -420 0 feedthrough
rlabel pdiffusion 654 -420 654 -420 0 feedthrough
rlabel pdiffusion 661 -420 661 -420 0 feedthrough
rlabel pdiffusion 668 -420 668 -420 0 feedthrough
rlabel pdiffusion 675 -420 675 -420 0 feedthrough
rlabel pdiffusion 682 -420 682 -420 0 feedthrough
rlabel pdiffusion 689 -420 689 -420 0 feedthrough
rlabel pdiffusion 696 -420 696 -420 0 feedthrough
rlabel pdiffusion 703 -420 703 -420 0 feedthrough
rlabel pdiffusion 710 -420 710 -420 0 feedthrough
rlabel pdiffusion 717 -420 717 -420 0 feedthrough
rlabel pdiffusion 724 -420 724 -420 0 feedthrough
rlabel pdiffusion 731 -420 731 -420 0 feedthrough
rlabel pdiffusion 738 -420 738 -420 0 feedthrough
rlabel pdiffusion 745 -420 745 -420 0 feedthrough
rlabel pdiffusion 752 -420 752 -420 0 feedthrough
rlabel pdiffusion 759 -420 759 -420 0 feedthrough
rlabel pdiffusion 766 -420 766 -420 0 feedthrough
rlabel pdiffusion 773 -420 773 -420 0 feedthrough
rlabel pdiffusion 780 -420 780 -420 0 feedthrough
rlabel pdiffusion 787 -420 787 -420 0 feedthrough
rlabel pdiffusion 794 -420 794 -420 0 feedthrough
rlabel pdiffusion 801 -420 801 -420 0 feedthrough
rlabel pdiffusion 808 -420 808 -420 0 feedthrough
rlabel pdiffusion 815 -420 815 -420 0 feedthrough
rlabel pdiffusion 3 -513 3 -513 0 cellNo=369
rlabel pdiffusion 10 -513 10 -513 0 feedthrough
rlabel pdiffusion 17 -513 17 -513 0 feedthrough
rlabel pdiffusion 24 -513 24 -513 0 feedthrough
rlabel pdiffusion 31 -513 31 -513 0 feedthrough
rlabel pdiffusion 38 -513 38 -513 0 feedthrough
rlabel pdiffusion 45 -513 45 -513 0 cellNo=160
rlabel pdiffusion 52 -513 52 -513 0 feedthrough
rlabel pdiffusion 59 -513 59 -513 0 cellNo=142
rlabel pdiffusion 66 -513 66 -513 0 feedthrough
rlabel pdiffusion 73 -513 73 -513 0 feedthrough
rlabel pdiffusion 80 -513 80 -513 0 feedthrough
rlabel pdiffusion 87 -513 87 -513 0 feedthrough
rlabel pdiffusion 94 -513 94 -513 0 feedthrough
rlabel pdiffusion 101 -513 101 -513 0 cellNo=216
rlabel pdiffusion 108 -513 108 -513 0 feedthrough
rlabel pdiffusion 115 -513 115 -513 0 feedthrough
rlabel pdiffusion 122 -513 122 -513 0 feedthrough
rlabel pdiffusion 129 -513 129 -513 0 feedthrough
rlabel pdiffusion 136 -513 136 -513 0 cellNo=58
rlabel pdiffusion 143 -513 143 -513 0 feedthrough
rlabel pdiffusion 150 -513 150 -513 0 feedthrough
rlabel pdiffusion 157 -513 157 -513 0 feedthrough
rlabel pdiffusion 164 -513 164 -513 0 feedthrough
rlabel pdiffusion 171 -513 171 -513 0 feedthrough
rlabel pdiffusion 178 -513 178 -513 0 feedthrough
rlabel pdiffusion 185 -513 185 -513 0 feedthrough
rlabel pdiffusion 192 -513 192 -513 0 feedthrough
rlabel pdiffusion 199 -513 199 -513 0 feedthrough
rlabel pdiffusion 206 -513 206 -513 0 feedthrough
rlabel pdiffusion 213 -513 213 -513 0 feedthrough
rlabel pdiffusion 220 -513 220 -513 0 cellNo=30
rlabel pdiffusion 227 -513 227 -513 0 cellNo=307
rlabel pdiffusion 234 -513 234 -513 0 feedthrough
rlabel pdiffusion 241 -513 241 -513 0 feedthrough
rlabel pdiffusion 248 -513 248 -513 0 feedthrough
rlabel pdiffusion 255 -513 255 -513 0 feedthrough
rlabel pdiffusion 262 -513 262 -513 0 cellNo=239
rlabel pdiffusion 269 -513 269 -513 0 feedthrough
rlabel pdiffusion 276 -513 276 -513 0 feedthrough
rlabel pdiffusion 283 -513 283 -513 0 feedthrough
rlabel pdiffusion 290 -513 290 -513 0 feedthrough
rlabel pdiffusion 297 -513 297 -513 0 feedthrough
rlabel pdiffusion 304 -513 304 -513 0 cellNo=207
rlabel pdiffusion 311 -513 311 -513 0 cellNo=99
rlabel pdiffusion 318 -513 318 -513 0 feedthrough
rlabel pdiffusion 325 -513 325 -513 0 feedthrough
rlabel pdiffusion 332 -513 332 -513 0 feedthrough
rlabel pdiffusion 339 -513 339 -513 0 feedthrough
rlabel pdiffusion 346 -513 346 -513 0 feedthrough
rlabel pdiffusion 353 -513 353 -513 0 cellNo=272
rlabel pdiffusion 360 -513 360 -513 0 feedthrough
rlabel pdiffusion 367 -513 367 -513 0 cellNo=111
rlabel pdiffusion 374 -513 374 -513 0 feedthrough
rlabel pdiffusion 381 -513 381 -513 0 cellNo=13
rlabel pdiffusion 388 -513 388 -513 0 cellNo=96
rlabel pdiffusion 395 -513 395 -513 0 feedthrough
rlabel pdiffusion 402 -513 402 -513 0 cellNo=71
rlabel pdiffusion 409 -513 409 -513 0 cellNo=196
rlabel pdiffusion 416 -513 416 -513 0 feedthrough
rlabel pdiffusion 423 -513 423 -513 0 feedthrough
rlabel pdiffusion 430 -513 430 -513 0 cellNo=22
rlabel pdiffusion 437 -513 437 -513 0 feedthrough
rlabel pdiffusion 444 -513 444 -513 0 feedthrough
rlabel pdiffusion 451 -513 451 -513 0 feedthrough
rlabel pdiffusion 458 -513 458 -513 0 feedthrough
rlabel pdiffusion 465 -513 465 -513 0 feedthrough
rlabel pdiffusion 472 -513 472 -513 0 cellNo=12
rlabel pdiffusion 479 -513 479 -513 0 feedthrough
rlabel pdiffusion 486 -513 486 -513 0 feedthrough
rlabel pdiffusion 493 -513 493 -513 0 cellNo=133
rlabel pdiffusion 500 -513 500 -513 0 feedthrough
rlabel pdiffusion 507 -513 507 -513 0 feedthrough
rlabel pdiffusion 514 -513 514 -513 0 feedthrough
rlabel pdiffusion 521 -513 521 -513 0 feedthrough
rlabel pdiffusion 528 -513 528 -513 0 feedthrough
rlabel pdiffusion 535 -513 535 -513 0 feedthrough
rlabel pdiffusion 542 -513 542 -513 0 feedthrough
rlabel pdiffusion 549 -513 549 -513 0 feedthrough
rlabel pdiffusion 556 -513 556 -513 0 cellNo=182
rlabel pdiffusion 563 -513 563 -513 0 feedthrough
rlabel pdiffusion 570 -513 570 -513 0 feedthrough
rlabel pdiffusion 577 -513 577 -513 0 feedthrough
rlabel pdiffusion 584 -513 584 -513 0 feedthrough
rlabel pdiffusion 591 -513 591 -513 0 feedthrough
rlabel pdiffusion 598 -513 598 -513 0 feedthrough
rlabel pdiffusion 605 -513 605 -513 0 feedthrough
rlabel pdiffusion 612 -513 612 -513 0 feedthrough
rlabel pdiffusion 619 -513 619 -513 0 feedthrough
rlabel pdiffusion 626 -513 626 -513 0 feedthrough
rlabel pdiffusion 633 -513 633 -513 0 feedthrough
rlabel pdiffusion 640 -513 640 -513 0 feedthrough
rlabel pdiffusion 647 -513 647 -513 0 feedthrough
rlabel pdiffusion 654 -513 654 -513 0 feedthrough
rlabel pdiffusion 661 -513 661 -513 0 feedthrough
rlabel pdiffusion 668 -513 668 -513 0 feedthrough
rlabel pdiffusion 675 -513 675 -513 0 feedthrough
rlabel pdiffusion 682 -513 682 -513 0 feedthrough
rlabel pdiffusion 689 -513 689 -513 0 feedthrough
rlabel pdiffusion 696 -513 696 -513 0 feedthrough
rlabel pdiffusion 703 -513 703 -513 0 feedthrough
rlabel pdiffusion 710 -513 710 -513 0 feedthrough
rlabel pdiffusion 717 -513 717 -513 0 feedthrough
rlabel pdiffusion 724 -513 724 -513 0 feedthrough
rlabel pdiffusion 731 -513 731 -513 0 feedthrough
rlabel pdiffusion 738 -513 738 -513 0 feedthrough
rlabel pdiffusion 745 -513 745 -513 0 feedthrough
rlabel pdiffusion 752 -513 752 -513 0 feedthrough
rlabel pdiffusion 759 -513 759 -513 0 feedthrough
rlabel pdiffusion 766 -513 766 -513 0 feedthrough
rlabel pdiffusion 773 -513 773 -513 0 feedthrough
rlabel pdiffusion 780 -513 780 -513 0 feedthrough
rlabel pdiffusion 787 -513 787 -513 0 feedthrough
rlabel pdiffusion 794 -513 794 -513 0 feedthrough
rlabel pdiffusion 801 -513 801 -513 0 feedthrough
rlabel pdiffusion 3 -582 3 -582 0 cellNo=279
rlabel pdiffusion 10 -582 10 -582 0 feedthrough
rlabel pdiffusion 17 -582 17 -582 0 feedthrough
rlabel pdiffusion 24 -582 24 -582 0 cellNo=54
rlabel pdiffusion 31 -582 31 -582 0 feedthrough
rlabel pdiffusion 38 -582 38 -582 0 feedthrough
rlabel pdiffusion 45 -582 45 -582 0 feedthrough
rlabel pdiffusion 52 -582 52 -582 0 cellNo=276
rlabel pdiffusion 59 -582 59 -582 0 feedthrough
rlabel pdiffusion 66 -582 66 -582 0 feedthrough
rlabel pdiffusion 73 -582 73 -582 0 feedthrough
rlabel pdiffusion 80 -582 80 -582 0 feedthrough
rlabel pdiffusion 87 -582 87 -582 0 feedthrough
rlabel pdiffusion 94 -582 94 -582 0 feedthrough
rlabel pdiffusion 101 -582 101 -582 0 feedthrough
rlabel pdiffusion 108 -582 108 -582 0 cellNo=238
rlabel pdiffusion 115 -582 115 -582 0 feedthrough
rlabel pdiffusion 122 -582 122 -582 0 cellNo=157
rlabel pdiffusion 129 -582 129 -582 0 cellNo=271
rlabel pdiffusion 136 -582 136 -582 0 cellNo=218
rlabel pdiffusion 143 -582 143 -582 0 feedthrough
rlabel pdiffusion 150 -582 150 -582 0 feedthrough
rlabel pdiffusion 157 -582 157 -582 0 feedthrough
rlabel pdiffusion 164 -582 164 -582 0 feedthrough
rlabel pdiffusion 171 -582 171 -582 0 feedthrough
rlabel pdiffusion 178 -582 178 -582 0 feedthrough
rlabel pdiffusion 185 -582 185 -582 0 feedthrough
rlabel pdiffusion 192 -582 192 -582 0 feedthrough
rlabel pdiffusion 199 -582 199 -582 0 feedthrough
rlabel pdiffusion 206 -582 206 -582 0 feedthrough
rlabel pdiffusion 213 -582 213 -582 0 feedthrough
rlabel pdiffusion 220 -582 220 -582 0 feedthrough
rlabel pdiffusion 227 -582 227 -582 0 feedthrough
rlabel pdiffusion 234 -582 234 -582 0 feedthrough
rlabel pdiffusion 241 -582 241 -582 0 feedthrough
rlabel pdiffusion 248 -582 248 -582 0 feedthrough
rlabel pdiffusion 255 -582 255 -582 0 cellNo=91
rlabel pdiffusion 262 -582 262 -582 0 feedthrough
rlabel pdiffusion 269 -582 269 -582 0 feedthrough
rlabel pdiffusion 276 -582 276 -582 0 feedthrough
rlabel pdiffusion 283 -582 283 -582 0 feedthrough
rlabel pdiffusion 290 -582 290 -582 0 feedthrough
rlabel pdiffusion 297 -582 297 -582 0 cellNo=219
rlabel pdiffusion 304 -582 304 -582 0 feedthrough
rlabel pdiffusion 311 -582 311 -582 0 cellNo=53
rlabel pdiffusion 318 -582 318 -582 0 cellNo=314
rlabel pdiffusion 325 -582 325 -582 0 feedthrough
rlabel pdiffusion 332 -582 332 -582 0 cellNo=273
rlabel pdiffusion 339 -582 339 -582 0 feedthrough
rlabel pdiffusion 346 -582 346 -582 0 feedthrough
rlabel pdiffusion 353 -582 353 -582 0 feedthrough
rlabel pdiffusion 360 -582 360 -582 0 feedthrough
rlabel pdiffusion 367 -582 367 -582 0 feedthrough
rlabel pdiffusion 374 -582 374 -582 0 feedthrough
rlabel pdiffusion 381 -582 381 -582 0 cellNo=50
rlabel pdiffusion 388 -582 388 -582 0 feedthrough
rlabel pdiffusion 395 -582 395 -582 0 feedthrough
rlabel pdiffusion 402 -582 402 -582 0 feedthrough
rlabel pdiffusion 409 -582 409 -582 0 feedthrough
rlabel pdiffusion 416 -582 416 -582 0 cellNo=318
rlabel pdiffusion 423 -582 423 -582 0 feedthrough
rlabel pdiffusion 430 -582 430 -582 0 feedthrough
rlabel pdiffusion 437 -582 437 -582 0 feedthrough
rlabel pdiffusion 444 -582 444 -582 0 feedthrough
rlabel pdiffusion 451 -582 451 -582 0 feedthrough
rlabel pdiffusion 458 -582 458 -582 0 cellNo=167
rlabel pdiffusion 465 -582 465 -582 0 cellNo=115
rlabel pdiffusion 472 -582 472 -582 0 feedthrough
rlabel pdiffusion 479 -582 479 -582 0 feedthrough
rlabel pdiffusion 486 -582 486 -582 0 cellNo=64
rlabel pdiffusion 493 -582 493 -582 0 feedthrough
rlabel pdiffusion 500 -582 500 -582 0 feedthrough
rlabel pdiffusion 507 -582 507 -582 0 cellNo=150
rlabel pdiffusion 514 -582 514 -582 0 cellNo=202
rlabel pdiffusion 521 -582 521 -582 0 feedthrough
rlabel pdiffusion 528 -582 528 -582 0 feedthrough
rlabel pdiffusion 535 -582 535 -582 0 feedthrough
rlabel pdiffusion 542 -582 542 -582 0 feedthrough
rlabel pdiffusion 549 -582 549 -582 0 cellNo=28
rlabel pdiffusion 556 -582 556 -582 0 feedthrough
rlabel pdiffusion 563 -582 563 -582 0 feedthrough
rlabel pdiffusion 570 -582 570 -582 0 feedthrough
rlabel pdiffusion 577 -582 577 -582 0 feedthrough
rlabel pdiffusion 584 -582 584 -582 0 feedthrough
rlabel pdiffusion 591 -582 591 -582 0 feedthrough
rlabel pdiffusion 598 -582 598 -582 0 feedthrough
rlabel pdiffusion 605 -582 605 -582 0 feedthrough
rlabel pdiffusion 612 -582 612 -582 0 feedthrough
rlabel pdiffusion 619 -582 619 -582 0 feedthrough
rlabel pdiffusion 626 -582 626 -582 0 feedthrough
rlabel pdiffusion 633 -582 633 -582 0 feedthrough
rlabel pdiffusion 640 -582 640 -582 0 feedthrough
rlabel pdiffusion 647 -582 647 -582 0 feedthrough
rlabel pdiffusion 654 -582 654 -582 0 feedthrough
rlabel pdiffusion 661 -582 661 -582 0 feedthrough
rlabel pdiffusion 668 -582 668 -582 0 feedthrough
rlabel pdiffusion 675 -582 675 -582 0 feedthrough
rlabel pdiffusion 682 -582 682 -582 0 feedthrough
rlabel pdiffusion 689 -582 689 -582 0 feedthrough
rlabel pdiffusion 696 -582 696 -582 0 feedthrough
rlabel pdiffusion 703 -582 703 -582 0 feedthrough
rlabel pdiffusion 710 -582 710 -582 0 feedthrough
rlabel pdiffusion 717 -582 717 -582 0 feedthrough
rlabel pdiffusion 724 -582 724 -582 0 feedthrough
rlabel pdiffusion 731 -582 731 -582 0 feedthrough
rlabel pdiffusion 738 -582 738 -582 0 feedthrough
rlabel pdiffusion 745 -582 745 -582 0 feedthrough
rlabel pdiffusion 752 -582 752 -582 0 feedthrough
rlabel pdiffusion 759 -582 759 -582 0 feedthrough
rlabel pdiffusion 766 -582 766 -582 0 feedthrough
rlabel pdiffusion 773 -582 773 -582 0 feedthrough
rlabel pdiffusion 780 -582 780 -582 0 feedthrough
rlabel pdiffusion 787 -582 787 -582 0 feedthrough
rlabel pdiffusion 794 -582 794 -582 0 feedthrough
rlabel pdiffusion 801 -582 801 -582 0 feedthrough
rlabel pdiffusion 808 -582 808 -582 0 feedthrough
rlabel pdiffusion 815 -582 815 -582 0 feedthrough
rlabel pdiffusion 822 -582 822 -582 0 feedthrough
rlabel pdiffusion 3 -671 3 -671 0 feedthrough
rlabel pdiffusion 10 -671 10 -671 0 feedthrough
rlabel pdiffusion 17 -671 17 -671 0 feedthrough
rlabel pdiffusion 24 -671 24 -671 0 feedthrough
rlabel pdiffusion 31 -671 31 -671 0 feedthrough
rlabel pdiffusion 38 -671 38 -671 0 feedthrough
rlabel pdiffusion 45 -671 45 -671 0 feedthrough
rlabel pdiffusion 52 -671 52 -671 0 cellNo=66
rlabel pdiffusion 59 -671 59 -671 0 cellNo=154
rlabel pdiffusion 66 -671 66 -671 0 cellNo=315
rlabel pdiffusion 73 -671 73 -671 0 feedthrough
rlabel pdiffusion 80 -671 80 -671 0 feedthrough
rlabel pdiffusion 87 -671 87 -671 0 feedthrough
rlabel pdiffusion 94 -671 94 -671 0 feedthrough
rlabel pdiffusion 101 -671 101 -671 0 feedthrough
rlabel pdiffusion 108 -671 108 -671 0 cellNo=262
rlabel pdiffusion 115 -671 115 -671 0 cellNo=63
rlabel pdiffusion 122 -671 122 -671 0 feedthrough
rlabel pdiffusion 129 -671 129 -671 0 feedthrough
rlabel pdiffusion 136 -671 136 -671 0 feedthrough
rlabel pdiffusion 143 -671 143 -671 0 cellNo=40
rlabel pdiffusion 150 -671 150 -671 0 feedthrough
rlabel pdiffusion 157 -671 157 -671 0 feedthrough
rlabel pdiffusion 164 -671 164 -671 0 feedthrough
rlabel pdiffusion 171 -671 171 -671 0 feedthrough
rlabel pdiffusion 178 -671 178 -671 0 feedthrough
rlabel pdiffusion 185 -671 185 -671 0 feedthrough
rlabel pdiffusion 192 -671 192 -671 0 feedthrough
rlabel pdiffusion 199 -671 199 -671 0 feedthrough
rlabel pdiffusion 206 -671 206 -671 0 feedthrough
rlabel pdiffusion 213 -671 213 -671 0 cellNo=155
rlabel pdiffusion 220 -671 220 -671 0 feedthrough
rlabel pdiffusion 227 -671 227 -671 0 cellNo=265
rlabel pdiffusion 234 -671 234 -671 0 feedthrough
rlabel pdiffusion 241 -671 241 -671 0 feedthrough
rlabel pdiffusion 248 -671 248 -671 0 feedthrough
rlabel pdiffusion 255 -671 255 -671 0 feedthrough
rlabel pdiffusion 262 -671 262 -671 0 feedthrough
rlabel pdiffusion 269 -671 269 -671 0 cellNo=37
rlabel pdiffusion 276 -671 276 -671 0 feedthrough
rlabel pdiffusion 283 -671 283 -671 0 feedthrough
rlabel pdiffusion 290 -671 290 -671 0 cellNo=105
rlabel pdiffusion 297 -671 297 -671 0 cellNo=232
rlabel pdiffusion 304 -671 304 -671 0 feedthrough
rlabel pdiffusion 311 -671 311 -671 0 feedthrough
rlabel pdiffusion 318 -671 318 -671 0 feedthrough
rlabel pdiffusion 325 -671 325 -671 0 feedthrough
rlabel pdiffusion 332 -671 332 -671 0 feedthrough
rlabel pdiffusion 339 -671 339 -671 0 feedthrough
rlabel pdiffusion 346 -671 346 -671 0 cellNo=21
rlabel pdiffusion 353 -671 353 -671 0 feedthrough
rlabel pdiffusion 360 -671 360 -671 0 feedthrough
rlabel pdiffusion 367 -671 367 -671 0 cellNo=89
rlabel pdiffusion 374 -671 374 -671 0 feedthrough
rlabel pdiffusion 381 -671 381 -671 0 cellNo=122
rlabel pdiffusion 388 -671 388 -671 0 feedthrough
rlabel pdiffusion 395 -671 395 -671 0 feedthrough
rlabel pdiffusion 402 -671 402 -671 0 feedthrough
rlabel pdiffusion 409 -671 409 -671 0 feedthrough
rlabel pdiffusion 416 -671 416 -671 0 cellNo=151
rlabel pdiffusion 423 -671 423 -671 0 feedthrough
rlabel pdiffusion 430 -671 430 -671 0 feedthrough
rlabel pdiffusion 437 -671 437 -671 0 feedthrough
rlabel pdiffusion 444 -671 444 -671 0 feedthrough
rlabel pdiffusion 451 -671 451 -671 0 cellNo=85
rlabel pdiffusion 458 -671 458 -671 0 cellNo=249
rlabel pdiffusion 465 -671 465 -671 0 feedthrough
rlabel pdiffusion 472 -671 472 -671 0 feedthrough
rlabel pdiffusion 479 -671 479 -671 0 feedthrough
rlabel pdiffusion 486 -671 486 -671 0 feedthrough
rlabel pdiffusion 493 -671 493 -671 0 feedthrough
rlabel pdiffusion 500 -671 500 -671 0 feedthrough
rlabel pdiffusion 507 -671 507 -671 0 feedthrough
rlabel pdiffusion 514 -671 514 -671 0 feedthrough
rlabel pdiffusion 521 -671 521 -671 0 feedthrough
rlabel pdiffusion 528 -671 528 -671 0 feedthrough
rlabel pdiffusion 535 -671 535 -671 0 feedthrough
rlabel pdiffusion 542 -671 542 -671 0 cellNo=347
rlabel pdiffusion 549 -671 549 -671 0 feedthrough
rlabel pdiffusion 556 -671 556 -671 0 feedthrough
rlabel pdiffusion 563 -671 563 -671 0 feedthrough
rlabel pdiffusion 570 -671 570 -671 0 feedthrough
rlabel pdiffusion 577 -671 577 -671 0 feedthrough
rlabel pdiffusion 584 -671 584 -671 0 feedthrough
rlabel pdiffusion 591 -671 591 -671 0 feedthrough
rlabel pdiffusion 598 -671 598 -671 0 feedthrough
rlabel pdiffusion 605 -671 605 -671 0 feedthrough
rlabel pdiffusion 612 -671 612 -671 0 feedthrough
rlabel pdiffusion 619 -671 619 -671 0 feedthrough
rlabel pdiffusion 626 -671 626 -671 0 feedthrough
rlabel pdiffusion 633 -671 633 -671 0 feedthrough
rlabel pdiffusion 640 -671 640 -671 0 feedthrough
rlabel pdiffusion 647 -671 647 -671 0 feedthrough
rlabel pdiffusion 654 -671 654 -671 0 feedthrough
rlabel pdiffusion 661 -671 661 -671 0 feedthrough
rlabel pdiffusion 668 -671 668 -671 0 feedthrough
rlabel pdiffusion 675 -671 675 -671 0 feedthrough
rlabel pdiffusion 682 -671 682 -671 0 feedthrough
rlabel pdiffusion 689 -671 689 -671 0 feedthrough
rlabel pdiffusion 696 -671 696 -671 0 feedthrough
rlabel pdiffusion 703 -671 703 -671 0 feedthrough
rlabel pdiffusion 710 -671 710 -671 0 feedthrough
rlabel pdiffusion 717 -671 717 -671 0 feedthrough
rlabel pdiffusion 724 -671 724 -671 0 feedthrough
rlabel pdiffusion 731 -671 731 -671 0 feedthrough
rlabel pdiffusion 738 -671 738 -671 0 feedthrough
rlabel pdiffusion 745 -671 745 -671 0 feedthrough
rlabel pdiffusion 752 -671 752 -671 0 feedthrough
rlabel pdiffusion 759 -671 759 -671 0 feedthrough
rlabel pdiffusion 766 -671 766 -671 0 feedthrough
rlabel pdiffusion 773 -671 773 -671 0 feedthrough
rlabel pdiffusion 780 -671 780 -671 0 feedthrough
rlabel pdiffusion 787 -671 787 -671 0 cellNo=134
rlabel pdiffusion 794 -671 794 -671 0 cellNo=221
rlabel pdiffusion 10 -738 10 -738 0 cellNo=81
rlabel pdiffusion 17 -738 17 -738 0 cellNo=76
rlabel pdiffusion 24 -738 24 -738 0 feedthrough
rlabel pdiffusion 31 -738 31 -738 0 feedthrough
rlabel pdiffusion 38 -738 38 -738 0 feedthrough
rlabel pdiffusion 45 -738 45 -738 0 feedthrough
rlabel pdiffusion 52 -738 52 -738 0 feedthrough
rlabel pdiffusion 59 -738 59 -738 0 feedthrough
rlabel pdiffusion 66 -738 66 -738 0 cellNo=100
rlabel pdiffusion 73 -738 73 -738 0 feedthrough
rlabel pdiffusion 80 -738 80 -738 0 feedthrough
rlabel pdiffusion 87 -738 87 -738 0 cellNo=179
rlabel pdiffusion 94 -738 94 -738 0 feedthrough
rlabel pdiffusion 101 -738 101 -738 0 feedthrough
rlabel pdiffusion 108 -738 108 -738 0 feedthrough
rlabel pdiffusion 115 -738 115 -738 0 feedthrough
rlabel pdiffusion 122 -738 122 -738 0 feedthrough
rlabel pdiffusion 129 -738 129 -738 0 cellNo=247
rlabel pdiffusion 136 -738 136 -738 0 feedthrough
rlabel pdiffusion 143 -738 143 -738 0 feedthrough
rlabel pdiffusion 150 -738 150 -738 0 feedthrough
rlabel pdiffusion 157 -738 157 -738 0 feedthrough
rlabel pdiffusion 164 -738 164 -738 0 cellNo=361
rlabel pdiffusion 171 -738 171 -738 0 feedthrough
rlabel pdiffusion 178 -738 178 -738 0 feedthrough
rlabel pdiffusion 185 -738 185 -738 0 feedthrough
rlabel pdiffusion 192 -738 192 -738 0 feedthrough
rlabel pdiffusion 199 -738 199 -738 0 feedthrough
rlabel pdiffusion 206 -738 206 -738 0 feedthrough
rlabel pdiffusion 213 -738 213 -738 0 feedthrough
rlabel pdiffusion 220 -738 220 -738 0 feedthrough
rlabel pdiffusion 227 -738 227 -738 0 cellNo=309
rlabel pdiffusion 234 -738 234 -738 0 feedthrough
rlabel pdiffusion 241 -738 241 -738 0 feedthrough
rlabel pdiffusion 248 -738 248 -738 0 feedthrough
rlabel pdiffusion 255 -738 255 -738 0 feedthrough
rlabel pdiffusion 262 -738 262 -738 0 feedthrough
rlabel pdiffusion 269 -738 269 -738 0 cellNo=4
rlabel pdiffusion 276 -738 276 -738 0 feedthrough
rlabel pdiffusion 283 -738 283 -738 0 feedthrough
rlabel pdiffusion 290 -738 290 -738 0 feedthrough
rlabel pdiffusion 297 -738 297 -738 0 feedthrough
rlabel pdiffusion 304 -738 304 -738 0 feedthrough
rlabel pdiffusion 311 -738 311 -738 0 feedthrough
rlabel pdiffusion 318 -738 318 -738 0 cellNo=290
rlabel pdiffusion 325 -738 325 -738 0 feedthrough
rlabel pdiffusion 332 -738 332 -738 0 feedthrough
rlabel pdiffusion 339 -738 339 -738 0 feedthrough
rlabel pdiffusion 346 -738 346 -738 0 cellNo=173
rlabel pdiffusion 353 -738 353 -738 0 feedthrough
rlabel pdiffusion 360 -738 360 -738 0 feedthrough
rlabel pdiffusion 367 -738 367 -738 0 feedthrough
rlabel pdiffusion 374 -738 374 -738 0 feedthrough
rlabel pdiffusion 381 -738 381 -738 0 cellNo=243
rlabel pdiffusion 388 -738 388 -738 0 feedthrough
rlabel pdiffusion 395 -738 395 -738 0 cellNo=263
rlabel pdiffusion 402 -738 402 -738 0 feedthrough
rlabel pdiffusion 409 -738 409 -738 0 feedthrough
rlabel pdiffusion 416 -738 416 -738 0 feedthrough
rlabel pdiffusion 423 -738 423 -738 0 cellNo=345
rlabel pdiffusion 430 -738 430 -738 0 feedthrough
rlabel pdiffusion 437 -738 437 -738 0 feedthrough
rlabel pdiffusion 444 -738 444 -738 0 cellNo=236
rlabel pdiffusion 451 -738 451 -738 0 feedthrough
rlabel pdiffusion 458 -738 458 -738 0 feedthrough
rlabel pdiffusion 465 -738 465 -738 0 feedthrough
rlabel pdiffusion 472 -738 472 -738 0 feedthrough
rlabel pdiffusion 479 -738 479 -738 0 feedthrough
rlabel pdiffusion 486 -738 486 -738 0 feedthrough
rlabel pdiffusion 493 -738 493 -738 0 feedthrough
rlabel pdiffusion 500 -738 500 -738 0 feedthrough
rlabel pdiffusion 507 -738 507 -738 0 feedthrough
rlabel pdiffusion 514 -738 514 -738 0 feedthrough
rlabel pdiffusion 521 -738 521 -738 0 cellNo=336
rlabel pdiffusion 528 -738 528 -738 0 cellNo=86
rlabel pdiffusion 535 -738 535 -738 0 feedthrough
rlabel pdiffusion 542 -738 542 -738 0 feedthrough
rlabel pdiffusion 549 -738 549 -738 0 cellNo=260
rlabel pdiffusion 556 -738 556 -738 0 feedthrough
rlabel pdiffusion 563 -738 563 -738 0 feedthrough
rlabel pdiffusion 570 -738 570 -738 0 cellNo=2
rlabel pdiffusion 577 -738 577 -738 0 feedthrough
rlabel pdiffusion 584 -738 584 -738 0 feedthrough
rlabel pdiffusion 591 -738 591 -738 0 feedthrough
rlabel pdiffusion 598 -738 598 -738 0 feedthrough
rlabel pdiffusion 605 -738 605 -738 0 feedthrough
rlabel pdiffusion 612 -738 612 -738 0 feedthrough
rlabel pdiffusion 619 -738 619 -738 0 feedthrough
rlabel pdiffusion 626 -738 626 -738 0 feedthrough
rlabel pdiffusion 633 -738 633 -738 0 feedthrough
rlabel pdiffusion 640 -738 640 -738 0 feedthrough
rlabel pdiffusion 647 -738 647 -738 0 feedthrough
rlabel pdiffusion 654 -738 654 -738 0 feedthrough
rlabel pdiffusion 661 -738 661 -738 0 feedthrough
rlabel pdiffusion 668 -738 668 -738 0 feedthrough
rlabel pdiffusion 675 -738 675 -738 0 feedthrough
rlabel pdiffusion 682 -738 682 -738 0 feedthrough
rlabel pdiffusion 689 -738 689 -738 0 feedthrough
rlabel pdiffusion 696 -738 696 -738 0 feedthrough
rlabel pdiffusion 703 -738 703 -738 0 feedthrough
rlabel pdiffusion 710 -738 710 -738 0 feedthrough
rlabel pdiffusion 717 -738 717 -738 0 feedthrough
rlabel pdiffusion 724 -738 724 -738 0 feedthrough
rlabel pdiffusion 731 -738 731 -738 0 feedthrough
rlabel pdiffusion 738 -738 738 -738 0 feedthrough
rlabel pdiffusion 745 -738 745 -738 0 feedthrough
rlabel pdiffusion 752 -738 752 -738 0 feedthrough
rlabel pdiffusion 759 -738 759 -738 0 feedthrough
rlabel pdiffusion 766 -738 766 -738 0 feedthrough
rlabel pdiffusion 773 -738 773 -738 0 feedthrough
rlabel pdiffusion 780 -738 780 -738 0 cellNo=338
rlabel pdiffusion 787 -738 787 -738 0 feedthrough
rlabel pdiffusion 794 -738 794 -738 0 cellNo=313
rlabel pdiffusion 801 -738 801 -738 0 feedthrough
rlabel pdiffusion 808 -738 808 -738 0 feedthrough
rlabel pdiffusion 3 -809 3 -809 0 cellNo=52
rlabel pdiffusion 10 -809 10 -809 0 feedthrough
rlabel pdiffusion 17 -809 17 -809 0 feedthrough
rlabel pdiffusion 24 -809 24 -809 0 feedthrough
rlabel pdiffusion 31 -809 31 -809 0 feedthrough
rlabel pdiffusion 38 -809 38 -809 0 cellNo=215
rlabel pdiffusion 45 -809 45 -809 0 feedthrough
rlabel pdiffusion 52 -809 52 -809 0 feedthrough
rlabel pdiffusion 59 -809 59 -809 0 feedthrough
rlabel pdiffusion 66 -809 66 -809 0 feedthrough
rlabel pdiffusion 73 -809 73 -809 0 cellNo=277
rlabel pdiffusion 80 -809 80 -809 0 feedthrough
rlabel pdiffusion 87 -809 87 -809 0 feedthrough
rlabel pdiffusion 94 -809 94 -809 0 feedthrough
rlabel pdiffusion 101 -809 101 -809 0 feedthrough
rlabel pdiffusion 108 -809 108 -809 0 feedthrough
rlabel pdiffusion 115 -809 115 -809 0 feedthrough
rlabel pdiffusion 122 -809 122 -809 0 feedthrough
rlabel pdiffusion 129 -809 129 -809 0 cellNo=163
rlabel pdiffusion 136 -809 136 -809 0 feedthrough
rlabel pdiffusion 143 -809 143 -809 0 feedthrough
rlabel pdiffusion 150 -809 150 -809 0 feedthrough
rlabel pdiffusion 157 -809 157 -809 0 cellNo=181
rlabel pdiffusion 164 -809 164 -809 0 feedthrough
rlabel pdiffusion 171 -809 171 -809 0 feedthrough
rlabel pdiffusion 178 -809 178 -809 0 feedthrough
rlabel pdiffusion 185 -809 185 -809 0 feedthrough
rlabel pdiffusion 192 -809 192 -809 0 feedthrough
rlabel pdiffusion 199 -809 199 -809 0 feedthrough
rlabel pdiffusion 206 -809 206 -809 0 feedthrough
rlabel pdiffusion 213 -809 213 -809 0 cellNo=124
rlabel pdiffusion 220 -809 220 -809 0 feedthrough
rlabel pdiffusion 227 -809 227 -809 0 feedthrough
rlabel pdiffusion 234 -809 234 -809 0 feedthrough
rlabel pdiffusion 241 -809 241 -809 0 feedthrough
rlabel pdiffusion 248 -809 248 -809 0 cellNo=107
rlabel pdiffusion 255 -809 255 -809 0 cellNo=317
rlabel pdiffusion 262 -809 262 -809 0 feedthrough
rlabel pdiffusion 269 -809 269 -809 0 feedthrough
rlabel pdiffusion 276 -809 276 -809 0 feedthrough
rlabel pdiffusion 283 -809 283 -809 0 cellNo=256
rlabel pdiffusion 290 -809 290 -809 0 feedthrough
rlabel pdiffusion 297 -809 297 -809 0 feedthrough
rlabel pdiffusion 304 -809 304 -809 0 feedthrough
rlabel pdiffusion 311 -809 311 -809 0 cellNo=280
rlabel pdiffusion 318 -809 318 -809 0 feedthrough
rlabel pdiffusion 325 -809 325 -809 0 feedthrough
rlabel pdiffusion 332 -809 332 -809 0 feedthrough
rlabel pdiffusion 339 -809 339 -809 0 feedthrough
rlabel pdiffusion 346 -809 346 -809 0 feedthrough
rlabel pdiffusion 353 -809 353 -809 0 feedthrough
rlabel pdiffusion 360 -809 360 -809 0 cellNo=153
rlabel pdiffusion 367 -809 367 -809 0 feedthrough
rlabel pdiffusion 374 -809 374 -809 0 cellNo=1
rlabel pdiffusion 381 -809 381 -809 0 feedthrough
rlabel pdiffusion 388 -809 388 -809 0 feedthrough
rlabel pdiffusion 395 -809 395 -809 0 cellNo=259
rlabel pdiffusion 402 -809 402 -809 0 cellNo=377
rlabel pdiffusion 409 -809 409 -809 0 cellNo=125
rlabel pdiffusion 416 -809 416 -809 0 feedthrough
rlabel pdiffusion 423 -809 423 -809 0 feedthrough
rlabel pdiffusion 430 -809 430 -809 0 feedthrough
rlabel pdiffusion 437 -809 437 -809 0 feedthrough
rlabel pdiffusion 444 -809 444 -809 0 feedthrough
rlabel pdiffusion 451 -809 451 -809 0 feedthrough
rlabel pdiffusion 458 -809 458 -809 0 feedthrough
rlabel pdiffusion 465 -809 465 -809 0 feedthrough
rlabel pdiffusion 472 -809 472 -809 0 feedthrough
rlabel pdiffusion 479 -809 479 -809 0 cellNo=45
rlabel pdiffusion 486 -809 486 -809 0 feedthrough
rlabel pdiffusion 493 -809 493 -809 0 feedthrough
rlabel pdiffusion 500 -809 500 -809 0 feedthrough
rlabel pdiffusion 507 -809 507 -809 0 feedthrough
rlabel pdiffusion 514 -809 514 -809 0 feedthrough
rlabel pdiffusion 521 -809 521 -809 0 feedthrough
rlabel pdiffusion 528 -809 528 -809 0 feedthrough
rlabel pdiffusion 535 -809 535 -809 0 feedthrough
rlabel pdiffusion 542 -809 542 -809 0 feedthrough
rlabel pdiffusion 549 -809 549 -809 0 cellNo=306
rlabel pdiffusion 556 -809 556 -809 0 feedthrough
rlabel pdiffusion 563 -809 563 -809 0 feedthrough
rlabel pdiffusion 570 -809 570 -809 0 feedthrough
rlabel pdiffusion 577 -809 577 -809 0 feedthrough
rlabel pdiffusion 584 -809 584 -809 0 feedthrough
rlabel pdiffusion 591 -809 591 -809 0 feedthrough
rlabel pdiffusion 598 -809 598 -809 0 cellNo=224
rlabel pdiffusion 605 -809 605 -809 0 feedthrough
rlabel pdiffusion 612 -809 612 -809 0 feedthrough
rlabel pdiffusion 619 -809 619 -809 0 cellNo=339
rlabel pdiffusion 626 -809 626 -809 0 feedthrough
rlabel pdiffusion 633 -809 633 -809 0 feedthrough
rlabel pdiffusion 640 -809 640 -809 0 feedthrough
rlabel pdiffusion 647 -809 647 -809 0 feedthrough
rlabel pdiffusion 654 -809 654 -809 0 feedthrough
rlabel pdiffusion 661 -809 661 -809 0 feedthrough
rlabel pdiffusion 668 -809 668 -809 0 feedthrough
rlabel pdiffusion 675 -809 675 -809 0 feedthrough
rlabel pdiffusion 682 -809 682 -809 0 feedthrough
rlabel pdiffusion 689 -809 689 -809 0 feedthrough
rlabel pdiffusion 696 -809 696 -809 0 feedthrough
rlabel pdiffusion 703 -809 703 -809 0 feedthrough
rlabel pdiffusion 710 -809 710 -809 0 feedthrough
rlabel pdiffusion 717 -809 717 -809 0 feedthrough
rlabel pdiffusion 724 -809 724 -809 0 feedthrough
rlabel pdiffusion 731 -809 731 -809 0 feedthrough
rlabel pdiffusion 738 -809 738 -809 0 feedthrough
rlabel pdiffusion 745 -809 745 -809 0 feedthrough
rlabel pdiffusion 752 -809 752 -809 0 feedthrough
rlabel pdiffusion 759 -809 759 -809 0 feedthrough
rlabel pdiffusion 766 -809 766 -809 0 feedthrough
rlabel pdiffusion 773 -809 773 -809 0 cellNo=204
rlabel pdiffusion 780 -809 780 -809 0 feedthrough
rlabel pdiffusion 787 -809 787 -809 0 feedthrough
rlabel pdiffusion 3 -864 3 -864 0 cellNo=131
rlabel pdiffusion 10 -864 10 -864 0 feedthrough
rlabel pdiffusion 17 -864 17 -864 0 cellNo=303
rlabel pdiffusion 24 -864 24 -864 0 feedthrough
rlabel pdiffusion 31 -864 31 -864 0 feedthrough
rlabel pdiffusion 38 -864 38 -864 0 cellNo=281
rlabel pdiffusion 45 -864 45 -864 0 feedthrough
rlabel pdiffusion 52 -864 52 -864 0 cellNo=234
rlabel pdiffusion 59 -864 59 -864 0 feedthrough
rlabel pdiffusion 66 -864 66 -864 0 feedthrough
rlabel pdiffusion 73 -864 73 -864 0 feedthrough
rlabel pdiffusion 80 -864 80 -864 0 feedthrough
rlabel pdiffusion 87 -864 87 -864 0 feedthrough
rlabel pdiffusion 94 -864 94 -864 0 feedthrough
rlabel pdiffusion 101 -864 101 -864 0 feedthrough
rlabel pdiffusion 108 -864 108 -864 0 cellNo=367
rlabel pdiffusion 115 -864 115 -864 0 cellNo=46
rlabel pdiffusion 122 -864 122 -864 0 feedthrough
rlabel pdiffusion 129 -864 129 -864 0 feedthrough
rlabel pdiffusion 136 -864 136 -864 0 cellNo=387
rlabel pdiffusion 143 -864 143 -864 0 feedthrough
rlabel pdiffusion 150 -864 150 -864 0 feedthrough
rlabel pdiffusion 157 -864 157 -864 0 feedthrough
rlabel pdiffusion 164 -864 164 -864 0 feedthrough
rlabel pdiffusion 171 -864 171 -864 0 cellNo=79
rlabel pdiffusion 178 -864 178 -864 0 feedthrough
rlabel pdiffusion 185 -864 185 -864 0 feedthrough
rlabel pdiffusion 192 -864 192 -864 0 feedthrough
rlabel pdiffusion 199 -864 199 -864 0 feedthrough
rlabel pdiffusion 206 -864 206 -864 0 feedthrough
rlabel pdiffusion 213 -864 213 -864 0 feedthrough
rlabel pdiffusion 220 -864 220 -864 0 feedthrough
rlabel pdiffusion 227 -864 227 -864 0 feedthrough
rlabel pdiffusion 234 -864 234 -864 0 feedthrough
rlabel pdiffusion 241 -864 241 -864 0 feedthrough
rlabel pdiffusion 248 -864 248 -864 0 feedthrough
rlabel pdiffusion 255 -864 255 -864 0 feedthrough
rlabel pdiffusion 262 -864 262 -864 0 cellNo=380
rlabel pdiffusion 269 -864 269 -864 0 cellNo=210
rlabel pdiffusion 276 -864 276 -864 0 feedthrough
rlabel pdiffusion 283 -864 283 -864 0 feedthrough
rlabel pdiffusion 290 -864 290 -864 0 feedthrough
rlabel pdiffusion 297 -864 297 -864 0 feedthrough
rlabel pdiffusion 304 -864 304 -864 0 feedthrough
rlabel pdiffusion 311 -864 311 -864 0 feedthrough
rlabel pdiffusion 318 -864 318 -864 0 feedthrough
rlabel pdiffusion 325 -864 325 -864 0 feedthrough
rlabel pdiffusion 332 -864 332 -864 0 feedthrough
rlabel pdiffusion 339 -864 339 -864 0 feedthrough
rlabel pdiffusion 346 -864 346 -864 0 cellNo=353
rlabel pdiffusion 353 -864 353 -864 0 feedthrough
rlabel pdiffusion 360 -864 360 -864 0 feedthrough
rlabel pdiffusion 367 -864 367 -864 0 cellNo=145
rlabel pdiffusion 374 -864 374 -864 0 feedthrough
rlabel pdiffusion 381 -864 381 -864 0 cellNo=398
rlabel pdiffusion 388 -864 388 -864 0 cellNo=296
rlabel pdiffusion 395 -864 395 -864 0 feedthrough
rlabel pdiffusion 402 -864 402 -864 0 feedthrough
rlabel pdiffusion 409 -864 409 -864 0 feedthrough
rlabel pdiffusion 416 -864 416 -864 0 feedthrough
rlabel pdiffusion 423 -864 423 -864 0 feedthrough
rlabel pdiffusion 430 -864 430 -864 0 feedthrough
rlabel pdiffusion 437 -864 437 -864 0 feedthrough
rlabel pdiffusion 444 -864 444 -864 0 feedthrough
rlabel pdiffusion 451 -864 451 -864 0 feedthrough
rlabel pdiffusion 458 -864 458 -864 0 feedthrough
rlabel pdiffusion 465 -864 465 -864 0 feedthrough
rlabel pdiffusion 472 -864 472 -864 0 feedthrough
rlabel pdiffusion 479 -864 479 -864 0 feedthrough
rlabel pdiffusion 486 -864 486 -864 0 feedthrough
rlabel pdiffusion 493 -864 493 -864 0 feedthrough
rlabel pdiffusion 500 -864 500 -864 0 cellNo=385
rlabel pdiffusion 507 -864 507 -864 0 feedthrough
rlabel pdiffusion 514 -864 514 -864 0 feedthrough
rlabel pdiffusion 521 -864 521 -864 0 feedthrough
rlabel pdiffusion 528 -864 528 -864 0 feedthrough
rlabel pdiffusion 535 -864 535 -864 0 feedthrough
rlabel pdiffusion 542 -864 542 -864 0 cellNo=217
rlabel pdiffusion 549 -864 549 -864 0 feedthrough
rlabel pdiffusion 556 -864 556 -864 0 feedthrough
rlabel pdiffusion 563 -864 563 -864 0 feedthrough
rlabel pdiffusion 570 -864 570 -864 0 feedthrough
rlabel pdiffusion 577 -864 577 -864 0 feedthrough
rlabel pdiffusion 584 -864 584 -864 0 feedthrough
rlabel pdiffusion 591 -864 591 -864 0 feedthrough
rlabel pdiffusion 598 -864 598 -864 0 feedthrough
rlabel pdiffusion 605 -864 605 -864 0 cellNo=267
rlabel pdiffusion 612 -864 612 -864 0 feedthrough
rlabel pdiffusion 619 -864 619 -864 0 feedthrough
rlabel pdiffusion 626 -864 626 -864 0 feedthrough
rlabel pdiffusion 633 -864 633 -864 0 feedthrough
rlabel pdiffusion 640 -864 640 -864 0 feedthrough
rlabel pdiffusion 647 -864 647 -864 0 feedthrough
rlabel pdiffusion 654 -864 654 -864 0 feedthrough
rlabel pdiffusion 661 -864 661 -864 0 feedthrough
rlabel pdiffusion 668 -864 668 -864 0 feedthrough
rlabel pdiffusion 682 -864 682 -864 0 cellNo=208
rlabel pdiffusion 689 -864 689 -864 0 feedthrough
rlabel pdiffusion 696 -864 696 -864 0 feedthrough
rlabel pdiffusion 703 -864 703 -864 0 feedthrough
rlabel pdiffusion 724 -864 724 -864 0 cellNo=185
rlabel pdiffusion 731 -864 731 -864 0 cellNo=328
rlabel pdiffusion 738 -864 738 -864 0 feedthrough
rlabel pdiffusion 745 -864 745 -864 0 feedthrough
rlabel pdiffusion 752 -864 752 -864 0 feedthrough
rlabel pdiffusion 759 -864 759 -864 0 feedthrough
rlabel pdiffusion 3 -917 3 -917 0 cellNo=128
rlabel pdiffusion 45 -917 45 -917 0 feedthrough
rlabel pdiffusion 52 -917 52 -917 0 feedthrough
rlabel pdiffusion 59 -917 59 -917 0 feedthrough
rlabel pdiffusion 66 -917 66 -917 0 feedthrough
rlabel pdiffusion 73 -917 73 -917 0 cellNo=48
rlabel pdiffusion 80 -917 80 -917 0 feedthrough
rlabel pdiffusion 87 -917 87 -917 0 feedthrough
rlabel pdiffusion 94 -917 94 -917 0 feedthrough
rlabel pdiffusion 101 -917 101 -917 0 feedthrough
rlabel pdiffusion 108 -917 108 -917 0 feedthrough
rlabel pdiffusion 115 -917 115 -917 0 feedthrough
rlabel pdiffusion 122 -917 122 -917 0 cellNo=103
rlabel pdiffusion 129 -917 129 -917 0 feedthrough
rlabel pdiffusion 136 -917 136 -917 0 feedthrough
rlabel pdiffusion 143 -917 143 -917 0 feedthrough
rlabel pdiffusion 150 -917 150 -917 0 feedthrough
rlabel pdiffusion 157 -917 157 -917 0 cellNo=104
rlabel pdiffusion 164 -917 164 -917 0 feedthrough
rlabel pdiffusion 171 -917 171 -917 0 feedthrough
rlabel pdiffusion 178 -917 178 -917 0 cellNo=250
rlabel pdiffusion 185 -917 185 -917 0 feedthrough
rlabel pdiffusion 192 -917 192 -917 0 feedthrough
rlabel pdiffusion 199 -917 199 -917 0 cellNo=297
rlabel pdiffusion 206 -917 206 -917 0 cellNo=251
rlabel pdiffusion 213 -917 213 -917 0 feedthrough
rlabel pdiffusion 220 -917 220 -917 0 feedthrough
rlabel pdiffusion 227 -917 227 -917 0 feedthrough
rlabel pdiffusion 234 -917 234 -917 0 feedthrough
rlabel pdiffusion 241 -917 241 -917 0 feedthrough
rlabel pdiffusion 248 -917 248 -917 0 feedthrough
rlabel pdiffusion 255 -917 255 -917 0 cellNo=274
rlabel pdiffusion 262 -917 262 -917 0 feedthrough
rlabel pdiffusion 269 -917 269 -917 0 cellNo=26
rlabel pdiffusion 276 -917 276 -917 0 feedthrough
rlabel pdiffusion 283 -917 283 -917 0 feedthrough
rlabel pdiffusion 290 -917 290 -917 0 feedthrough
rlabel pdiffusion 297 -917 297 -917 0 cellNo=143
rlabel pdiffusion 304 -917 304 -917 0 feedthrough
rlabel pdiffusion 311 -917 311 -917 0 feedthrough
rlabel pdiffusion 318 -917 318 -917 0 feedthrough
rlabel pdiffusion 325 -917 325 -917 0 cellNo=320
rlabel pdiffusion 332 -917 332 -917 0 feedthrough
rlabel pdiffusion 339 -917 339 -917 0 feedthrough
rlabel pdiffusion 346 -917 346 -917 0 feedthrough
rlabel pdiffusion 353 -917 353 -917 0 feedthrough
rlabel pdiffusion 360 -917 360 -917 0 feedthrough
rlabel pdiffusion 367 -917 367 -917 0 cellNo=159
rlabel pdiffusion 374 -917 374 -917 0 cellNo=316
rlabel pdiffusion 381 -917 381 -917 0 feedthrough
rlabel pdiffusion 388 -917 388 -917 0 feedthrough
rlabel pdiffusion 395 -917 395 -917 0 cellNo=325
rlabel pdiffusion 402 -917 402 -917 0 feedthrough
rlabel pdiffusion 409 -917 409 -917 0 feedthrough
rlabel pdiffusion 416 -917 416 -917 0 feedthrough
rlabel pdiffusion 423 -917 423 -917 0 feedthrough
rlabel pdiffusion 430 -917 430 -917 0 feedthrough
rlabel pdiffusion 437 -917 437 -917 0 feedthrough
rlabel pdiffusion 444 -917 444 -917 0 feedthrough
rlabel pdiffusion 451 -917 451 -917 0 feedthrough
rlabel pdiffusion 458 -917 458 -917 0 feedthrough
rlabel pdiffusion 465 -917 465 -917 0 cellNo=87
rlabel pdiffusion 472 -917 472 -917 0 feedthrough
rlabel pdiffusion 479 -917 479 -917 0 feedthrough
rlabel pdiffusion 486 -917 486 -917 0 feedthrough
rlabel pdiffusion 493 -917 493 -917 0 feedthrough
rlabel pdiffusion 500 -917 500 -917 0 feedthrough
rlabel pdiffusion 507 -917 507 -917 0 feedthrough
rlabel pdiffusion 514 -917 514 -917 0 feedthrough
rlabel pdiffusion 521 -917 521 -917 0 cellNo=227
rlabel pdiffusion 528 -917 528 -917 0 feedthrough
rlabel pdiffusion 535 -917 535 -917 0 feedthrough
rlabel pdiffusion 542 -917 542 -917 0 feedthrough
rlabel pdiffusion 549 -917 549 -917 0 feedthrough
rlabel pdiffusion 556 -917 556 -917 0 feedthrough
rlabel pdiffusion 563 -917 563 -917 0 feedthrough
rlabel pdiffusion 570 -917 570 -917 0 feedthrough
rlabel pdiffusion 577 -917 577 -917 0 feedthrough
rlabel pdiffusion 584 -917 584 -917 0 feedthrough
rlabel pdiffusion 591 -917 591 -917 0 feedthrough
rlabel pdiffusion 598 -917 598 -917 0 feedthrough
rlabel pdiffusion 605 -917 605 -917 0 feedthrough
rlabel pdiffusion 612 -917 612 -917 0 feedthrough
rlabel pdiffusion 619 -917 619 -917 0 feedthrough
rlabel pdiffusion 626 -917 626 -917 0 feedthrough
rlabel pdiffusion 633 -917 633 -917 0 feedthrough
rlabel pdiffusion 640 -917 640 -917 0 cellNo=44
rlabel pdiffusion 647 -917 647 -917 0 feedthrough
rlabel pdiffusion 654 -917 654 -917 0 cellNo=355
rlabel pdiffusion 661 -917 661 -917 0 cellNo=292
rlabel pdiffusion 668 -917 668 -917 0 feedthrough
rlabel pdiffusion 675 -917 675 -917 0 feedthrough
rlabel pdiffusion 682 -917 682 -917 0 feedthrough
rlabel pdiffusion 717 -917 717 -917 0 feedthrough
rlabel pdiffusion 745 -917 745 -917 0 cellNo=300
rlabel pdiffusion 3 -976 3 -976 0 cellNo=241
rlabel pdiffusion 10 -976 10 -976 0 cellNo=324
rlabel pdiffusion 17 -976 17 -976 0 cellNo=351
rlabel pdiffusion 66 -976 66 -976 0 feedthrough
rlabel pdiffusion 73 -976 73 -976 0 feedthrough
rlabel pdiffusion 80 -976 80 -976 0 feedthrough
rlabel pdiffusion 87 -976 87 -976 0 feedthrough
rlabel pdiffusion 94 -976 94 -976 0 cellNo=349
rlabel pdiffusion 101 -976 101 -976 0 cellNo=299
rlabel pdiffusion 108 -976 108 -976 0 cellNo=346
rlabel pdiffusion 115 -976 115 -976 0 cellNo=69
rlabel pdiffusion 122 -976 122 -976 0 feedthrough
rlabel pdiffusion 129 -976 129 -976 0 feedthrough
rlabel pdiffusion 136 -976 136 -976 0 feedthrough
rlabel pdiffusion 143 -976 143 -976 0 feedthrough
rlabel pdiffusion 150 -976 150 -976 0 feedthrough
rlabel pdiffusion 157 -976 157 -976 0 feedthrough
rlabel pdiffusion 164 -976 164 -976 0 feedthrough
rlabel pdiffusion 171 -976 171 -976 0 feedthrough
rlabel pdiffusion 178 -976 178 -976 0 feedthrough
rlabel pdiffusion 185 -976 185 -976 0 feedthrough
rlabel pdiffusion 192 -976 192 -976 0 feedthrough
rlabel pdiffusion 199 -976 199 -976 0 cellNo=39
rlabel pdiffusion 206 -976 206 -976 0 feedthrough
rlabel pdiffusion 213 -976 213 -976 0 feedthrough
rlabel pdiffusion 220 -976 220 -976 0 feedthrough
rlabel pdiffusion 227 -976 227 -976 0 cellNo=396
rlabel pdiffusion 234 -976 234 -976 0 feedthrough
rlabel pdiffusion 241 -976 241 -976 0 feedthrough
rlabel pdiffusion 248 -976 248 -976 0 feedthrough
rlabel pdiffusion 255 -976 255 -976 0 feedthrough
rlabel pdiffusion 262 -976 262 -976 0 feedthrough
rlabel pdiffusion 269 -976 269 -976 0 feedthrough
rlabel pdiffusion 276 -976 276 -976 0 feedthrough
rlabel pdiffusion 283 -976 283 -976 0 feedthrough
rlabel pdiffusion 290 -976 290 -976 0 feedthrough
rlabel pdiffusion 297 -976 297 -976 0 feedthrough
rlabel pdiffusion 304 -976 304 -976 0 feedthrough
rlabel pdiffusion 311 -976 311 -976 0 cellNo=371
rlabel pdiffusion 318 -976 318 -976 0 cellNo=322
rlabel pdiffusion 325 -976 325 -976 0 feedthrough
rlabel pdiffusion 332 -976 332 -976 0 feedthrough
rlabel pdiffusion 339 -976 339 -976 0 feedthrough
rlabel pdiffusion 346 -976 346 -976 0 feedthrough
rlabel pdiffusion 353 -976 353 -976 0 feedthrough
rlabel pdiffusion 360 -976 360 -976 0 feedthrough
rlabel pdiffusion 367 -976 367 -976 0 cellNo=386
rlabel pdiffusion 374 -976 374 -976 0 cellNo=374
rlabel pdiffusion 381 -976 381 -976 0 feedthrough
rlabel pdiffusion 388 -976 388 -976 0 cellNo=192
rlabel pdiffusion 395 -976 395 -976 0 feedthrough
rlabel pdiffusion 402 -976 402 -976 0 feedthrough
rlabel pdiffusion 409 -976 409 -976 0 feedthrough
rlabel pdiffusion 416 -976 416 -976 0 cellNo=206
rlabel pdiffusion 423 -976 423 -976 0 cellNo=390
rlabel pdiffusion 430 -976 430 -976 0 feedthrough
rlabel pdiffusion 437 -976 437 -976 0 feedthrough
rlabel pdiffusion 444 -976 444 -976 0 feedthrough
rlabel pdiffusion 451 -976 451 -976 0 cellNo=329
rlabel pdiffusion 458 -976 458 -976 0 feedthrough
rlabel pdiffusion 465 -976 465 -976 0 feedthrough
rlabel pdiffusion 472 -976 472 -976 0 feedthrough
rlabel pdiffusion 479 -976 479 -976 0 feedthrough
rlabel pdiffusion 486 -976 486 -976 0 feedthrough
rlabel pdiffusion 493 -976 493 -976 0 feedthrough
rlabel pdiffusion 500 -976 500 -976 0 feedthrough
rlabel pdiffusion 507 -976 507 -976 0 feedthrough
rlabel pdiffusion 514 -976 514 -976 0 feedthrough
rlabel pdiffusion 521 -976 521 -976 0 cellNo=368
rlabel pdiffusion 528 -976 528 -976 0 feedthrough
rlabel pdiffusion 535 -976 535 -976 0 feedthrough
rlabel pdiffusion 542 -976 542 -976 0 cellNo=261
rlabel pdiffusion 549 -976 549 -976 0 feedthrough
rlabel pdiffusion 556 -976 556 -976 0 feedthrough
rlabel pdiffusion 563 -976 563 -976 0 feedthrough
rlabel pdiffusion 570 -976 570 -976 0 feedthrough
rlabel pdiffusion 577 -976 577 -976 0 feedthrough
rlabel pdiffusion 584 -976 584 -976 0 feedthrough
rlabel pdiffusion 591 -976 591 -976 0 feedthrough
rlabel pdiffusion 598 -976 598 -976 0 feedthrough
rlabel pdiffusion 605 -976 605 -976 0 feedthrough
rlabel pdiffusion 612 -976 612 -976 0 feedthrough
rlabel pdiffusion 619 -976 619 -976 0 feedthrough
rlabel pdiffusion 626 -976 626 -976 0 cellNo=248
rlabel pdiffusion 661 -976 661 -976 0 feedthrough
rlabel pdiffusion 675 -976 675 -976 0 feedthrough
rlabel pdiffusion 3 -1015 3 -1015 0 cellNo=148
rlabel pdiffusion 10 -1015 10 -1015 0 cellNo=360
rlabel pdiffusion 101 -1015 101 -1015 0 feedthrough
rlabel pdiffusion 143 -1015 143 -1015 0 feedthrough
rlabel pdiffusion 150 -1015 150 -1015 0 feedthrough
rlabel pdiffusion 157 -1015 157 -1015 0 feedthrough
rlabel pdiffusion 164 -1015 164 -1015 0 feedthrough
rlabel pdiffusion 171 -1015 171 -1015 0 feedthrough
rlabel pdiffusion 178 -1015 178 -1015 0 feedthrough
rlabel pdiffusion 185 -1015 185 -1015 0 feedthrough
rlabel pdiffusion 192 -1015 192 -1015 0 feedthrough
rlabel pdiffusion 199 -1015 199 -1015 0 feedthrough
rlabel pdiffusion 206 -1015 206 -1015 0 feedthrough
rlabel pdiffusion 213 -1015 213 -1015 0 cellNo=343
rlabel pdiffusion 220 -1015 220 -1015 0 feedthrough
rlabel pdiffusion 227 -1015 227 -1015 0 feedthrough
rlabel pdiffusion 234 -1015 234 -1015 0 feedthrough
rlabel pdiffusion 241 -1015 241 -1015 0 feedthrough
rlabel pdiffusion 248 -1015 248 -1015 0 cellNo=305
rlabel pdiffusion 255 -1015 255 -1015 0 feedthrough
rlabel pdiffusion 262 -1015 262 -1015 0 cellNo=220
rlabel pdiffusion 269 -1015 269 -1015 0 feedthrough
rlabel pdiffusion 276 -1015 276 -1015 0 feedthrough
rlabel pdiffusion 283 -1015 283 -1015 0 feedthrough
rlabel pdiffusion 290 -1015 290 -1015 0 feedthrough
rlabel pdiffusion 297 -1015 297 -1015 0 cellNo=341
rlabel pdiffusion 304 -1015 304 -1015 0 feedthrough
rlabel pdiffusion 311 -1015 311 -1015 0 feedthrough
rlabel pdiffusion 318 -1015 318 -1015 0 cellNo=357
rlabel pdiffusion 325 -1015 325 -1015 0 feedthrough
rlabel pdiffusion 332 -1015 332 -1015 0 cellNo=330
rlabel pdiffusion 339 -1015 339 -1015 0 feedthrough
rlabel pdiffusion 346 -1015 346 -1015 0 cellNo=354
rlabel pdiffusion 353 -1015 353 -1015 0 feedthrough
rlabel pdiffusion 360 -1015 360 -1015 0 cellNo=49
rlabel pdiffusion 367 -1015 367 -1015 0 cellNo=20
rlabel pdiffusion 374 -1015 374 -1015 0 feedthrough
rlabel pdiffusion 381 -1015 381 -1015 0 feedthrough
rlabel pdiffusion 388 -1015 388 -1015 0 feedthrough
rlabel pdiffusion 395 -1015 395 -1015 0 feedthrough
rlabel pdiffusion 402 -1015 402 -1015 0 feedthrough
rlabel pdiffusion 409 -1015 409 -1015 0 feedthrough
rlabel pdiffusion 416 -1015 416 -1015 0 feedthrough
rlabel pdiffusion 423 -1015 423 -1015 0 feedthrough
rlabel pdiffusion 430 -1015 430 -1015 0 cellNo=344
rlabel pdiffusion 437 -1015 437 -1015 0 cellNo=65
rlabel pdiffusion 444 -1015 444 -1015 0 cellNo=270
rlabel pdiffusion 451 -1015 451 -1015 0 feedthrough
rlabel pdiffusion 458 -1015 458 -1015 0 cellNo=327
rlabel pdiffusion 465 -1015 465 -1015 0 feedthrough
rlabel pdiffusion 493 -1015 493 -1015 0 feedthrough
rlabel pdiffusion 500 -1015 500 -1015 0 feedthrough
rlabel pdiffusion 507 -1015 507 -1015 0 feedthrough
rlabel pdiffusion 528 -1015 528 -1015 0 cellNo=183
rlabel pdiffusion 542 -1015 542 -1015 0 cellNo=359
rlabel pdiffusion 549 -1015 549 -1015 0 feedthrough
rlabel pdiffusion 570 -1015 570 -1015 0 feedthrough
rlabel pdiffusion 577 -1015 577 -1015 0 feedthrough
rlabel pdiffusion 584 -1015 584 -1015 0 feedthrough
rlabel pdiffusion 591 -1015 591 -1015 0 feedthrough
rlabel pdiffusion 605 -1015 605 -1015 0 cellNo=342
rlabel pdiffusion 612 -1015 612 -1015 0 feedthrough
rlabel pdiffusion 647 -1015 647 -1015 0 cellNo=331
rlabel pdiffusion 668 -1015 668 -1015 0 cellNo=358
rlabel pdiffusion 3 -1044 3 -1044 0 cellNo=362
rlabel pdiffusion 10 -1044 10 -1044 0 cellNo=375
rlabel pdiffusion 101 -1044 101 -1044 0 feedthrough
rlabel pdiffusion 115 -1044 115 -1044 0 feedthrough
rlabel pdiffusion 122 -1044 122 -1044 0 cellNo=364
rlabel pdiffusion 129 -1044 129 -1044 0 feedthrough
rlabel pdiffusion 136 -1044 136 -1044 0 feedthrough
rlabel pdiffusion 143 -1044 143 -1044 0 feedthrough
rlabel pdiffusion 150 -1044 150 -1044 0 feedthrough
rlabel pdiffusion 157 -1044 157 -1044 0 feedthrough
rlabel pdiffusion 164 -1044 164 -1044 0 feedthrough
rlabel pdiffusion 171 -1044 171 -1044 0 cellNo=340
rlabel pdiffusion 178 -1044 178 -1044 0 cellNo=397
rlabel pdiffusion 185 -1044 185 -1044 0 cellNo=129
rlabel pdiffusion 192 -1044 192 -1044 0 feedthrough
rlabel pdiffusion 199 -1044 199 -1044 0 feedthrough
rlabel pdiffusion 206 -1044 206 -1044 0 feedthrough
rlabel pdiffusion 213 -1044 213 -1044 0 cellNo=372
rlabel pdiffusion 220 -1044 220 -1044 0 feedthrough
rlabel pdiffusion 227 -1044 227 -1044 0 cellNo=298
rlabel pdiffusion 234 -1044 234 -1044 0 feedthrough
rlabel pdiffusion 241 -1044 241 -1044 0 cellNo=136
rlabel pdiffusion 248 -1044 248 -1044 0 feedthrough
rlabel pdiffusion 255 -1044 255 -1044 0 feedthrough
rlabel pdiffusion 262 -1044 262 -1044 0 cellNo=138
rlabel pdiffusion 269 -1044 269 -1044 0 feedthrough
rlabel pdiffusion 276 -1044 276 -1044 0 cellNo=321
rlabel pdiffusion 283 -1044 283 -1044 0 cellNo=363
rlabel pdiffusion 290 -1044 290 -1044 0 feedthrough
rlabel pdiffusion 297 -1044 297 -1044 0 feedthrough
rlabel pdiffusion 304 -1044 304 -1044 0 cellNo=366
rlabel pdiffusion 311 -1044 311 -1044 0 feedthrough
rlabel pdiffusion 318 -1044 318 -1044 0 feedthrough
rlabel pdiffusion 367 -1044 367 -1044 0 feedthrough
rlabel pdiffusion 374 -1044 374 -1044 0 cellNo=378
rlabel pdiffusion 381 -1044 381 -1044 0 cellNo=348
rlabel pdiffusion 388 -1044 388 -1044 0 feedthrough
rlabel pdiffusion 395 -1044 395 -1044 0 feedthrough
rlabel pdiffusion 402 -1044 402 -1044 0 cellNo=335
rlabel pdiffusion 409 -1044 409 -1044 0 feedthrough
rlabel pdiffusion 416 -1044 416 -1044 0 cellNo=326
rlabel pdiffusion 423 -1044 423 -1044 0 feedthrough
rlabel pdiffusion 430 -1044 430 -1044 0 feedthrough
rlabel pdiffusion 437 -1044 437 -1044 0 feedthrough
rlabel pdiffusion 444 -1044 444 -1044 0 feedthrough
rlabel pdiffusion 458 -1044 458 -1044 0 feedthrough
rlabel pdiffusion 472 -1044 472 -1044 0 cellNo=156
rlabel pdiffusion 479 -1044 479 -1044 0 feedthrough
rlabel pdiffusion 486 -1044 486 -1044 0 feedthrough
rlabel pdiffusion 542 -1044 542 -1044 0 cellNo=379
rlabel pdiffusion 549 -1044 549 -1044 0 feedthrough
rlabel pdiffusion 563 -1044 563 -1044 0 feedthrough
rlabel pdiffusion 570 -1044 570 -1044 0 feedthrough
rlabel pdiffusion 577 -1044 577 -1044 0 cellNo=365
rlabel pdiffusion 584 -1044 584 -1044 0 feedthrough
rlabel pdiffusion 591 -1044 591 -1044 0 feedthrough
rlabel pdiffusion 3 -1065 3 -1065 0 cellNo=165
rlabel pdiffusion 10 -1065 10 -1065 0 cellNo=392
rlabel pdiffusion 101 -1065 101 -1065 0 cellNo=174
rlabel pdiffusion 108 -1065 108 -1065 0 feedthrough
rlabel pdiffusion 136 -1065 136 -1065 0 cellNo=333
rlabel pdiffusion 143 -1065 143 -1065 0 cellNo=225
rlabel pdiffusion 150 -1065 150 -1065 0 feedthrough
rlabel pdiffusion 157 -1065 157 -1065 0 cellNo=269
rlabel pdiffusion 164 -1065 164 -1065 0 feedthrough
rlabel pdiffusion 171 -1065 171 -1065 0 cellNo=237
rlabel pdiffusion 192 -1065 192 -1065 0 cellNo=381
rlabel pdiffusion 199 -1065 199 -1065 0 feedthrough
rlabel pdiffusion 206 -1065 206 -1065 0 cellNo=395
rlabel pdiffusion 213 -1065 213 -1065 0 cellNo=388
rlabel pdiffusion 220 -1065 220 -1065 0 cellNo=212
rlabel pdiffusion 227 -1065 227 -1065 0 feedthrough
rlabel pdiffusion 234 -1065 234 -1065 0 feedthrough
rlabel pdiffusion 283 -1065 283 -1065 0 cellNo=400
rlabel pdiffusion 297 -1065 297 -1065 0 cellNo=391
rlabel pdiffusion 381 -1065 381 -1065 0 feedthrough
rlabel pdiffusion 395 -1065 395 -1065 0 cellNo=394
rlabel pdiffusion 409 -1065 409 -1065 0 cellNo=382
rlabel pdiffusion 430 -1065 430 -1065 0 feedthrough
rlabel pdiffusion 437 -1065 437 -1065 0 cellNo=399
rlabel pdiffusion 444 -1065 444 -1065 0 cellNo=389
rlabel pdiffusion 451 -1065 451 -1065 0 cellNo=393
rlabel pdiffusion 458 -1065 458 -1065 0 feedthrough
rlabel pdiffusion 563 -1065 563 -1065 0 cellNo=68
rlabel pdiffusion 577 -1065 577 -1065 0 cellNo=240
rlabel pdiffusion 584 -1065 584 -1065 0 feedthrough
rlabel polysilicon 114 -6 114 -6 0 1
rlabel polysilicon 121 -6 121 -6 0 1
rlabel polysilicon 121 -12 121 -12 0 3
rlabel polysilicon 128 -6 128 -6 0 1
rlabel polysilicon 131 -6 131 -6 0 2
rlabel polysilicon 135 -6 135 -6 0 1
rlabel polysilicon 135 -12 135 -12 0 3
rlabel polysilicon 142 -6 142 -6 0 1
rlabel polysilicon 149 -6 149 -6 0 1
rlabel polysilicon 156 -6 156 -6 0 1
rlabel polysilicon 156 -12 156 -12 0 3
rlabel polysilicon 163 -6 163 -6 0 1
rlabel polysilicon 166 -6 166 -6 0 2
rlabel polysilicon 173 -12 173 -12 0 4
rlabel polysilicon 177 -6 177 -6 0 1
rlabel polysilicon 177 -12 177 -12 0 3
rlabel polysilicon 184 -12 184 -12 0 3
rlabel polysilicon 187 -12 187 -12 0 4
rlabel polysilicon 191 -6 191 -6 0 1
rlabel polysilicon 191 -12 191 -12 0 3
rlabel polysilicon 198 -6 198 -6 0 1
rlabel polysilicon 201 -12 201 -12 0 4
rlabel polysilicon 208 -6 208 -6 0 2
rlabel polysilicon 215 -12 215 -12 0 4
rlabel polysilicon 236 -6 236 -6 0 2
rlabel polysilicon 236 -12 236 -12 0 4
rlabel polysilicon 247 -6 247 -6 0 1
rlabel polysilicon 247 -12 247 -12 0 3
rlabel polysilicon 296 -6 296 -6 0 1
rlabel polysilicon 296 -12 296 -12 0 3
rlabel polysilicon 313 -6 313 -6 0 2
rlabel polysilicon 313 -12 313 -12 0 4
rlabel polysilicon 317 -6 317 -6 0 1
rlabel polysilicon 317 -12 317 -12 0 3
rlabel polysilicon 331 -6 331 -6 0 1
rlabel polysilicon 331 -12 331 -12 0 3
rlabel polysilicon 338 -6 338 -6 0 1
rlabel polysilicon 348 -6 348 -6 0 2
rlabel polysilicon 352 -6 352 -6 0 1
rlabel polysilicon 352 -12 352 -12 0 3
rlabel polysilicon 373 -6 373 -6 0 1
rlabel polysilicon 373 -12 373 -12 0 3
rlabel polysilicon 422 -12 422 -12 0 3
rlabel polysilicon 65 -31 65 -31 0 3
rlabel polysilicon 72 -25 72 -25 0 1
rlabel polysilicon 72 -31 72 -31 0 3
rlabel polysilicon 79 -25 79 -25 0 1
rlabel polysilicon 79 -31 79 -31 0 3
rlabel polysilicon 89 -25 89 -25 0 2
rlabel polysilicon 96 -25 96 -25 0 2
rlabel polysilicon 96 -31 96 -31 0 4
rlabel polysilicon 100 -25 100 -25 0 1
rlabel polysilicon 100 -31 100 -31 0 3
rlabel polysilicon 107 -25 107 -25 0 1
rlabel polysilicon 107 -31 107 -31 0 3
rlabel polysilicon 117 -25 117 -25 0 2
rlabel polysilicon 117 -31 117 -31 0 4
rlabel polysilicon 121 -31 121 -31 0 3
rlabel polysilicon 128 -25 128 -25 0 1
rlabel polysilicon 131 -25 131 -25 0 2
rlabel polysilicon 135 -25 135 -25 0 1
rlabel polysilicon 135 -31 135 -31 0 3
rlabel polysilicon 142 -25 142 -25 0 1
rlabel polysilicon 142 -31 142 -31 0 3
rlabel polysilicon 149 -25 149 -25 0 1
rlabel polysilicon 149 -31 149 -31 0 3
rlabel polysilicon 156 -25 156 -25 0 1
rlabel polysilicon 159 -25 159 -25 0 2
rlabel polysilicon 159 -31 159 -31 0 4
rlabel polysilicon 166 -31 166 -31 0 4
rlabel polysilicon 170 -25 170 -25 0 1
rlabel polysilicon 170 -31 170 -31 0 3
rlabel polysilicon 177 -25 177 -25 0 1
rlabel polysilicon 177 -31 177 -31 0 3
rlabel polysilicon 184 -25 184 -25 0 1
rlabel polysilicon 184 -31 184 -31 0 3
rlabel polysilicon 191 -25 191 -25 0 1
rlabel polysilicon 191 -31 191 -31 0 3
rlabel polysilicon 198 -25 198 -25 0 1
rlabel polysilicon 205 -31 205 -31 0 3
rlabel polysilicon 212 -25 212 -25 0 1
rlabel polysilicon 212 -31 212 -31 0 3
rlabel polysilicon 219 -25 219 -25 0 1
rlabel polysilicon 222 -31 222 -31 0 4
rlabel polysilicon 229 -25 229 -25 0 2
rlabel polysilicon 226 -31 226 -31 0 3
rlabel polysilicon 233 -25 233 -25 0 1
rlabel polysilicon 233 -31 233 -31 0 3
rlabel polysilicon 240 -25 240 -25 0 1
rlabel polysilicon 240 -31 240 -31 0 3
rlabel polysilicon 250 -31 250 -31 0 4
rlabel polysilicon 254 -25 254 -25 0 1
rlabel polysilicon 254 -31 254 -31 0 3
rlabel polysilicon 261 -31 261 -31 0 3
rlabel polysilicon 264 -31 264 -31 0 4
rlabel polysilicon 282 -25 282 -25 0 1
rlabel polysilicon 282 -31 282 -31 0 3
rlabel polysilicon 296 -25 296 -25 0 1
rlabel polysilicon 296 -31 296 -31 0 3
rlabel polysilicon 303 -25 303 -25 0 1
rlabel polysilicon 303 -31 303 -31 0 3
rlabel polysilicon 313 -31 313 -31 0 4
rlabel polysilicon 327 -31 327 -31 0 4
rlabel polysilicon 331 -25 331 -25 0 1
rlabel polysilicon 331 -31 331 -31 0 3
rlabel polysilicon 345 -25 345 -25 0 1
rlabel polysilicon 345 -31 345 -31 0 3
rlabel polysilicon 352 -25 352 -25 0 1
rlabel polysilicon 352 -31 352 -31 0 3
rlabel polysilicon 394 -25 394 -25 0 1
rlabel polysilicon 394 -31 394 -31 0 3
rlabel polysilicon 404 -25 404 -25 0 2
rlabel polysilicon 429 -25 429 -25 0 1
rlabel polysilicon 429 -31 429 -31 0 3
rlabel polysilicon 436 -25 436 -25 0 1
rlabel polysilicon 436 -31 436 -31 0 3
rlabel polysilicon 485 -25 485 -25 0 1
rlabel polysilicon 488 -31 488 -31 0 4
rlabel polysilicon 555 -25 555 -25 0 1
rlabel polysilicon 555 -31 555 -31 0 3
rlabel polysilicon 51 -54 51 -54 0 1
rlabel polysilicon 51 -60 51 -60 0 3
rlabel polysilicon 58 -54 58 -54 0 1
rlabel polysilicon 65 -54 65 -54 0 1
rlabel polysilicon 65 -60 65 -60 0 3
rlabel polysilicon 72 -54 72 -54 0 1
rlabel polysilicon 72 -60 72 -60 0 3
rlabel polysilicon 82 -60 82 -60 0 4
rlabel polysilicon 86 -54 86 -54 0 1
rlabel polysilicon 86 -60 86 -60 0 3
rlabel polysilicon 93 -54 93 -54 0 1
rlabel polysilicon 93 -60 93 -60 0 3
rlabel polysilicon 100 -54 100 -54 0 1
rlabel polysilicon 100 -60 100 -60 0 3
rlabel polysilicon 107 -54 107 -54 0 1
rlabel polysilicon 107 -60 107 -60 0 3
rlabel polysilicon 114 -54 114 -54 0 1
rlabel polysilicon 114 -60 114 -60 0 3
rlabel polysilicon 121 -54 121 -54 0 1
rlabel polysilicon 121 -60 121 -60 0 3
rlabel polysilicon 128 -60 128 -60 0 3
rlabel polysilicon 131 -60 131 -60 0 4
rlabel polysilicon 135 -54 135 -54 0 1
rlabel polysilicon 135 -60 135 -60 0 3
rlabel polysilicon 142 -54 142 -54 0 1
rlabel polysilicon 142 -60 142 -60 0 3
rlabel polysilicon 149 -54 149 -54 0 1
rlabel polysilicon 149 -60 149 -60 0 3
rlabel polysilicon 156 -54 156 -54 0 1
rlabel polysilicon 159 -54 159 -54 0 2
rlabel polysilicon 163 -54 163 -54 0 1
rlabel polysilicon 163 -60 163 -60 0 3
rlabel polysilicon 170 -54 170 -54 0 1
rlabel polysilicon 170 -60 170 -60 0 3
rlabel polysilicon 177 -54 177 -54 0 1
rlabel polysilicon 177 -60 177 -60 0 3
rlabel polysilicon 184 -54 184 -54 0 1
rlabel polysilicon 184 -60 184 -60 0 3
rlabel polysilicon 194 -54 194 -54 0 2
rlabel polysilicon 191 -60 191 -60 0 3
rlabel polysilicon 198 -54 198 -54 0 1
rlabel polysilicon 198 -60 198 -60 0 3
rlabel polysilicon 205 -54 205 -54 0 1
rlabel polysilicon 205 -60 205 -60 0 3
rlabel polysilicon 215 -54 215 -54 0 2
rlabel polysilicon 215 -60 215 -60 0 4
rlabel polysilicon 219 -54 219 -54 0 1
rlabel polysilicon 219 -60 219 -60 0 3
rlabel polysilicon 226 -54 226 -54 0 1
rlabel polysilicon 229 -60 229 -60 0 4
rlabel polysilicon 233 -54 233 -54 0 1
rlabel polysilicon 233 -60 233 -60 0 3
rlabel polysilicon 240 -60 240 -60 0 3
rlabel polysilicon 243 -60 243 -60 0 4
rlabel polysilicon 247 -54 247 -54 0 1
rlabel polysilicon 247 -60 247 -60 0 3
rlabel polysilicon 254 -54 254 -54 0 1
rlabel polysilicon 254 -60 254 -60 0 3
rlabel polysilicon 261 -54 261 -54 0 1
rlabel polysilicon 261 -60 261 -60 0 3
rlabel polysilicon 268 -54 268 -54 0 1
rlabel polysilicon 268 -60 268 -60 0 3
rlabel polysilicon 275 -54 275 -54 0 1
rlabel polysilicon 275 -60 275 -60 0 3
rlabel polysilicon 285 -54 285 -54 0 2
rlabel polysilicon 285 -60 285 -60 0 4
rlabel polysilicon 289 -54 289 -54 0 1
rlabel polysilicon 289 -60 289 -60 0 3
rlabel polysilicon 296 -54 296 -54 0 1
rlabel polysilicon 296 -60 296 -60 0 3
rlabel polysilicon 303 -54 303 -54 0 1
rlabel polysilicon 313 -60 313 -60 0 4
rlabel polysilicon 317 -54 317 -54 0 1
rlabel polysilicon 324 -54 324 -54 0 1
rlabel polysilicon 324 -60 324 -60 0 3
rlabel polysilicon 331 -54 331 -54 0 1
rlabel polysilicon 331 -60 331 -60 0 3
rlabel polysilicon 338 -54 338 -54 0 1
rlabel polysilicon 338 -60 338 -60 0 3
rlabel polysilicon 345 -54 345 -54 0 1
rlabel polysilicon 345 -60 345 -60 0 3
rlabel polysilicon 352 -54 352 -54 0 1
rlabel polysilicon 352 -60 352 -60 0 3
rlabel polysilicon 359 -54 359 -54 0 1
rlabel polysilicon 359 -60 359 -60 0 3
rlabel polysilicon 366 -54 366 -54 0 1
rlabel polysilicon 366 -60 366 -60 0 3
rlabel polysilicon 373 -54 373 -54 0 1
rlabel polysilicon 373 -60 373 -60 0 3
rlabel polysilicon 380 -54 380 -54 0 1
rlabel polysilicon 387 -54 387 -54 0 1
rlabel polysilicon 387 -60 387 -60 0 3
rlabel polysilicon 394 -54 394 -54 0 1
rlabel polysilicon 394 -60 394 -60 0 3
rlabel polysilicon 404 -54 404 -54 0 2
rlabel polysilicon 401 -60 401 -60 0 3
rlabel polysilicon 415 -54 415 -54 0 1
rlabel polysilicon 415 -60 415 -60 0 3
rlabel polysilicon 443 -54 443 -54 0 1
rlabel polysilicon 443 -60 443 -60 0 3
rlabel polysilicon 450 -54 450 -54 0 1
rlabel polysilicon 450 -60 450 -60 0 3
rlabel polysilicon 457 -60 457 -60 0 3
rlabel polysilicon 576 -54 576 -54 0 1
rlabel polysilicon 576 -60 576 -60 0 3
rlabel polysilicon 30 -93 30 -93 0 1
rlabel polysilicon 30 -99 30 -99 0 3
rlabel polysilicon 37 -93 37 -93 0 1
rlabel polysilicon 37 -99 37 -99 0 3
rlabel polysilicon 44 -93 44 -93 0 1
rlabel polysilicon 44 -99 44 -99 0 3
rlabel polysilicon 51 -93 51 -93 0 1
rlabel polysilicon 51 -99 51 -99 0 3
rlabel polysilicon 58 -93 58 -93 0 1
rlabel polysilicon 58 -99 58 -99 0 3
rlabel polysilicon 65 -93 65 -93 0 1
rlabel polysilicon 68 -99 68 -99 0 4
rlabel polysilicon 72 -93 72 -93 0 1
rlabel polysilicon 72 -99 72 -99 0 3
rlabel polysilicon 79 -93 79 -93 0 1
rlabel polysilicon 79 -99 79 -99 0 3
rlabel polysilicon 86 -93 86 -93 0 1
rlabel polysilicon 86 -99 86 -99 0 3
rlabel polysilicon 96 -93 96 -93 0 2
rlabel polysilicon 96 -99 96 -99 0 4
rlabel polysilicon 100 -93 100 -93 0 1
rlabel polysilicon 100 -99 100 -99 0 3
rlabel polysilicon 107 -93 107 -93 0 1
rlabel polysilicon 107 -99 107 -99 0 3
rlabel polysilicon 114 -93 114 -93 0 1
rlabel polysilicon 114 -99 114 -99 0 3
rlabel polysilicon 121 -99 121 -99 0 3
rlabel polysilicon 124 -99 124 -99 0 4
rlabel polysilicon 128 -93 128 -93 0 1
rlabel polysilicon 131 -93 131 -93 0 2
rlabel polysilicon 135 -93 135 -93 0 1
rlabel polysilicon 135 -99 135 -99 0 3
rlabel polysilicon 142 -93 142 -93 0 1
rlabel polysilicon 142 -99 142 -99 0 3
rlabel polysilicon 152 -93 152 -93 0 2
rlabel polysilicon 149 -99 149 -99 0 3
rlabel polysilicon 156 -93 156 -93 0 1
rlabel polysilicon 156 -99 156 -99 0 3
rlabel polysilicon 159 -99 159 -99 0 4
rlabel polysilicon 163 -93 163 -93 0 1
rlabel polysilicon 163 -99 163 -99 0 3
rlabel polysilicon 170 -93 170 -93 0 1
rlabel polysilicon 170 -99 170 -99 0 3
rlabel polysilicon 177 -93 177 -93 0 1
rlabel polysilicon 177 -99 177 -99 0 3
rlabel polysilicon 184 -93 184 -93 0 1
rlabel polysilicon 184 -99 184 -99 0 3
rlabel polysilicon 191 -93 191 -93 0 1
rlabel polysilicon 191 -99 191 -99 0 3
rlabel polysilicon 198 -93 198 -93 0 1
rlabel polysilicon 198 -99 198 -99 0 3
rlabel polysilicon 205 -93 205 -93 0 1
rlabel polysilicon 205 -99 205 -99 0 3
rlabel polysilicon 212 -93 212 -93 0 1
rlabel polysilicon 212 -99 212 -99 0 3
rlabel polysilicon 219 -93 219 -93 0 1
rlabel polysilicon 219 -99 219 -99 0 3
rlabel polysilicon 226 -93 226 -93 0 1
rlabel polysilicon 226 -99 226 -99 0 3
rlabel polysilicon 233 -93 233 -93 0 1
rlabel polysilicon 233 -99 233 -99 0 3
rlabel polysilicon 240 -93 240 -93 0 1
rlabel polysilicon 240 -99 240 -99 0 3
rlabel polysilicon 243 -99 243 -99 0 4
rlabel polysilicon 247 -93 247 -93 0 1
rlabel polysilicon 247 -99 247 -99 0 3
rlabel polysilicon 257 -99 257 -99 0 4
rlabel polysilicon 261 -93 261 -93 0 1
rlabel polysilicon 261 -99 261 -99 0 3
rlabel polysilicon 268 -93 268 -93 0 1
rlabel polysilicon 268 -99 268 -99 0 3
rlabel polysilicon 275 -93 275 -93 0 1
rlabel polysilicon 275 -99 275 -99 0 3
rlabel polysilicon 282 -99 282 -99 0 3
rlabel polysilicon 289 -93 289 -93 0 1
rlabel polysilicon 289 -99 289 -99 0 3
rlabel polysilicon 296 -93 296 -93 0 1
rlabel polysilicon 296 -99 296 -99 0 3
rlabel polysilicon 303 -93 303 -93 0 1
rlabel polysilicon 303 -99 303 -99 0 3
rlabel polysilicon 313 -93 313 -93 0 2
rlabel polysilicon 313 -99 313 -99 0 4
rlabel polysilicon 320 -99 320 -99 0 4
rlabel polysilicon 324 -93 324 -93 0 1
rlabel polysilicon 324 -99 324 -99 0 3
rlabel polysilicon 331 -93 331 -93 0 1
rlabel polysilicon 331 -99 331 -99 0 3
rlabel polysilicon 338 -93 338 -93 0 1
rlabel polysilicon 338 -99 338 -99 0 3
rlabel polysilicon 345 -93 345 -93 0 1
rlabel polysilicon 345 -99 345 -99 0 3
rlabel polysilicon 355 -99 355 -99 0 4
rlabel polysilicon 359 -93 359 -93 0 1
rlabel polysilicon 359 -99 359 -99 0 3
rlabel polysilicon 369 -93 369 -93 0 2
rlabel polysilicon 366 -99 366 -99 0 3
rlabel polysilicon 373 -93 373 -93 0 1
rlabel polysilicon 373 -99 373 -99 0 3
rlabel polysilicon 380 -93 380 -93 0 1
rlabel polysilicon 380 -99 380 -99 0 3
rlabel polysilicon 387 -93 387 -93 0 1
rlabel polysilicon 387 -99 387 -99 0 3
rlabel polysilicon 394 -93 394 -93 0 1
rlabel polysilicon 394 -99 394 -99 0 3
rlabel polysilicon 401 -93 401 -93 0 1
rlabel polysilicon 401 -99 401 -99 0 3
rlabel polysilicon 408 -93 408 -93 0 1
rlabel polysilicon 408 -99 408 -99 0 3
rlabel polysilicon 415 -93 415 -93 0 1
rlabel polysilicon 415 -99 415 -99 0 3
rlabel polysilicon 425 -93 425 -93 0 2
rlabel polysilicon 429 -93 429 -93 0 1
rlabel polysilicon 429 -99 429 -99 0 3
rlabel polysilicon 436 -93 436 -93 0 1
rlabel polysilicon 436 -99 436 -99 0 3
rlabel polysilicon 443 -99 443 -99 0 3
rlabel polysilicon 446 -99 446 -99 0 4
rlabel polysilicon 450 -93 450 -93 0 1
rlabel polysilicon 450 -99 450 -99 0 3
rlabel polysilicon 457 -93 457 -93 0 1
rlabel polysilicon 460 -99 460 -99 0 4
rlabel polysilicon 464 -93 464 -93 0 1
rlabel polysilicon 464 -99 464 -99 0 3
rlabel polysilicon 471 -93 471 -93 0 1
rlabel polysilicon 471 -99 471 -99 0 3
rlabel polysilicon 478 -93 478 -93 0 1
rlabel polysilicon 478 -99 478 -99 0 3
rlabel polysilicon 492 -93 492 -93 0 1
rlabel polysilicon 492 -99 492 -99 0 3
rlabel polysilicon 523 -99 523 -99 0 4
rlabel polysilicon 527 -93 527 -93 0 1
rlabel polysilicon 530 -93 530 -93 0 2
rlabel polysilicon 576 -93 576 -93 0 1
rlabel polysilicon 576 -99 576 -99 0 3
rlabel polysilicon 590 -93 590 -93 0 1
rlabel polysilicon 590 -99 590 -99 0 3
rlabel polysilicon 9 -144 9 -144 0 1
rlabel polysilicon 9 -150 9 -150 0 3
rlabel polysilicon 16 -144 16 -144 0 1
rlabel polysilicon 16 -150 16 -150 0 3
rlabel polysilicon 26 -144 26 -144 0 2
rlabel polysilicon 30 -144 30 -144 0 1
rlabel polysilicon 30 -150 30 -150 0 3
rlabel polysilicon 37 -144 37 -144 0 1
rlabel polysilicon 37 -150 37 -150 0 3
rlabel polysilicon 44 -144 44 -144 0 1
rlabel polysilicon 44 -150 44 -150 0 3
rlabel polysilicon 51 -144 51 -144 0 1
rlabel polysilicon 51 -150 51 -150 0 3
rlabel polysilicon 58 -144 58 -144 0 1
rlabel polysilicon 58 -150 58 -150 0 3
rlabel polysilicon 65 -144 65 -144 0 1
rlabel polysilicon 65 -150 65 -150 0 3
rlabel polysilicon 72 -144 72 -144 0 1
rlabel polysilicon 75 -144 75 -144 0 2
rlabel polysilicon 72 -150 72 -150 0 3
rlabel polysilicon 79 -150 79 -150 0 3
rlabel polysilicon 82 -150 82 -150 0 4
rlabel polysilicon 86 -144 86 -144 0 1
rlabel polysilicon 86 -150 86 -150 0 3
rlabel polysilicon 93 -144 93 -144 0 1
rlabel polysilicon 96 -150 96 -150 0 4
rlabel polysilicon 100 -144 100 -144 0 1
rlabel polysilicon 100 -150 100 -150 0 3
rlabel polysilicon 107 -144 107 -144 0 1
rlabel polysilicon 107 -150 107 -150 0 3
rlabel polysilicon 114 -144 114 -144 0 1
rlabel polysilicon 114 -150 114 -150 0 3
rlabel polysilicon 121 -144 121 -144 0 1
rlabel polysilicon 121 -150 121 -150 0 3
rlabel polysilicon 128 -144 128 -144 0 1
rlabel polysilicon 128 -150 128 -150 0 3
rlabel polysilicon 135 -144 135 -144 0 1
rlabel polysilicon 135 -150 135 -150 0 3
rlabel polysilicon 142 -144 142 -144 0 1
rlabel polysilicon 142 -150 142 -150 0 3
rlabel polysilicon 149 -144 149 -144 0 1
rlabel polysilicon 149 -150 149 -150 0 3
rlabel polysilicon 156 -144 156 -144 0 1
rlabel polysilicon 156 -150 156 -150 0 3
rlabel polysilicon 166 -144 166 -144 0 2
rlabel polysilicon 170 -144 170 -144 0 1
rlabel polysilicon 173 -144 173 -144 0 2
rlabel polysilicon 170 -150 170 -150 0 3
rlabel polysilicon 173 -150 173 -150 0 4
rlabel polysilicon 177 -144 177 -144 0 1
rlabel polysilicon 177 -150 177 -150 0 3
rlabel polysilicon 184 -144 184 -144 0 1
rlabel polysilicon 184 -150 184 -150 0 3
rlabel polysilicon 191 -144 191 -144 0 1
rlabel polysilicon 191 -150 191 -150 0 3
rlabel polysilicon 198 -144 198 -144 0 1
rlabel polysilicon 198 -150 198 -150 0 3
rlabel polysilicon 205 -144 205 -144 0 1
rlabel polysilicon 205 -150 205 -150 0 3
rlabel polysilicon 212 -144 212 -144 0 1
rlabel polysilicon 212 -150 212 -150 0 3
rlabel polysilicon 219 -144 219 -144 0 1
rlabel polysilicon 222 -144 222 -144 0 2
rlabel polysilicon 219 -150 219 -150 0 3
rlabel polysilicon 222 -150 222 -150 0 4
rlabel polysilicon 226 -144 226 -144 0 1
rlabel polysilicon 226 -150 226 -150 0 3
rlabel polysilicon 233 -144 233 -144 0 1
rlabel polysilicon 233 -150 233 -150 0 3
rlabel polysilicon 240 -144 240 -144 0 1
rlabel polysilicon 240 -150 240 -150 0 3
rlabel polysilicon 247 -144 247 -144 0 1
rlabel polysilicon 247 -150 247 -150 0 3
rlabel polysilicon 257 -144 257 -144 0 2
rlabel polysilicon 257 -150 257 -150 0 4
rlabel polysilicon 261 -144 261 -144 0 1
rlabel polysilicon 261 -150 261 -150 0 3
rlabel polysilicon 268 -144 268 -144 0 1
rlabel polysilicon 268 -150 268 -150 0 3
rlabel polysilicon 275 -144 275 -144 0 1
rlabel polysilicon 278 -150 278 -150 0 4
rlabel polysilicon 282 -144 282 -144 0 1
rlabel polysilicon 282 -150 282 -150 0 3
rlabel polysilicon 289 -144 289 -144 0 1
rlabel polysilicon 292 -150 292 -150 0 4
rlabel polysilicon 296 -144 296 -144 0 1
rlabel polysilicon 296 -150 296 -150 0 3
rlabel polysilicon 303 -144 303 -144 0 1
rlabel polysilicon 303 -150 303 -150 0 3
rlabel polysilicon 310 -144 310 -144 0 1
rlabel polysilicon 313 -144 313 -144 0 2
rlabel polysilicon 313 -150 313 -150 0 4
rlabel polysilicon 320 -144 320 -144 0 2
rlabel polysilicon 317 -150 317 -150 0 3
rlabel polysilicon 320 -150 320 -150 0 4
rlabel polysilicon 324 -144 324 -144 0 1
rlabel polysilicon 324 -150 324 -150 0 3
rlabel polysilicon 331 -144 331 -144 0 1
rlabel polysilicon 331 -150 331 -150 0 3
rlabel polysilicon 338 -144 338 -144 0 1
rlabel polysilicon 338 -150 338 -150 0 3
rlabel polysilicon 345 -144 345 -144 0 1
rlabel polysilicon 345 -150 345 -150 0 3
rlabel polysilicon 352 -144 352 -144 0 1
rlabel polysilicon 352 -150 352 -150 0 3
rlabel polysilicon 359 -144 359 -144 0 1
rlabel polysilicon 359 -150 359 -150 0 3
rlabel polysilicon 366 -144 366 -144 0 1
rlabel polysilicon 366 -150 366 -150 0 3
rlabel polysilicon 373 -144 373 -144 0 1
rlabel polysilicon 373 -150 373 -150 0 3
rlabel polysilicon 380 -144 380 -144 0 1
rlabel polysilicon 380 -150 380 -150 0 3
rlabel polysilicon 387 -144 387 -144 0 1
rlabel polysilicon 387 -150 387 -150 0 3
rlabel polysilicon 394 -144 394 -144 0 1
rlabel polysilicon 394 -150 394 -150 0 3
rlabel polysilicon 401 -144 401 -144 0 1
rlabel polysilicon 401 -150 401 -150 0 3
rlabel polysilicon 408 -144 408 -144 0 1
rlabel polysilicon 408 -150 408 -150 0 3
rlabel polysilicon 415 -144 415 -144 0 1
rlabel polysilicon 415 -150 415 -150 0 3
rlabel polysilicon 418 -150 418 -150 0 4
rlabel polysilicon 422 -144 422 -144 0 1
rlabel polysilicon 422 -150 422 -150 0 3
rlabel polysilicon 429 -144 429 -144 0 1
rlabel polysilicon 429 -150 429 -150 0 3
rlabel polysilicon 436 -144 436 -144 0 1
rlabel polysilicon 436 -150 436 -150 0 3
rlabel polysilicon 443 -144 443 -144 0 1
rlabel polysilicon 443 -150 443 -150 0 3
rlabel polysilicon 450 -144 450 -144 0 1
rlabel polysilicon 450 -150 450 -150 0 3
rlabel polysilicon 457 -144 457 -144 0 1
rlabel polysilicon 457 -150 457 -150 0 3
rlabel polysilicon 464 -144 464 -144 0 1
rlabel polysilicon 464 -150 464 -150 0 3
rlabel polysilicon 474 -144 474 -144 0 2
rlabel polysilicon 471 -150 471 -150 0 3
rlabel polysilicon 478 -144 478 -144 0 1
rlabel polysilicon 478 -150 478 -150 0 3
rlabel polysilicon 485 -144 485 -144 0 1
rlabel polysilicon 485 -150 485 -150 0 3
rlabel polysilicon 492 -144 492 -144 0 1
rlabel polysilicon 492 -150 492 -150 0 3
rlabel polysilicon 499 -144 499 -144 0 1
rlabel polysilicon 506 -144 506 -144 0 1
rlabel polysilicon 506 -150 506 -150 0 3
rlabel polysilicon 513 -144 513 -144 0 1
rlabel polysilicon 513 -150 513 -150 0 3
rlabel polysilicon 520 -144 520 -144 0 1
rlabel polysilicon 520 -150 520 -150 0 3
rlabel polysilicon 527 -144 527 -144 0 1
rlabel polysilicon 527 -150 527 -150 0 3
rlabel polysilicon 534 -144 534 -144 0 1
rlabel polysilicon 534 -150 534 -150 0 3
rlabel polysilicon 541 -144 541 -144 0 1
rlabel polysilicon 541 -150 541 -150 0 3
rlabel polysilicon 548 -144 548 -144 0 1
rlabel polysilicon 548 -150 548 -150 0 3
rlabel polysilicon 555 -144 555 -144 0 1
rlabel polysilicon 555 -150 555 -150 0 3
rlabel polysilicon 562 -144 562 -144 0 1
rlabel polysilicon 562 -150 562 -150 0 3
rlabel polysilicon 569 -144 569 -144 0 1
rlabel polysilicon 569 -150 569 -150 0 3
rlabel polysilicon 576 -144 576 -144 0 1
rlabel polysilicon 576 -150 576 -150 0 3
rlabel polysilicon 586 -144 586 -144 0 2
rlabel polysilicon 583 -150 583 -150 0 3
rlabel polysilicon 586 -150 586 -150 0 4
rlabel polysilicon 590 -144 590 -144 0 1
rlabel polysilicon 590 -150 590 -150 0 3
rlabel polysilicon 597 -144 597 -144 0 1
rlabel polysilicon 597 -150 597 -150 0 3
rlabel polysilicon 604 -144 604 -144 0 1
rlabel polysilicon 604 -150 604 -150 0 3
rlabel polysilicon 611 -144 611 -144 0 1
rlabel polysilicon 611 -150 611 -150 0 3
rlabel polysilicon 618 -144 618 -144 0 1
rlabel polysilicon 618 -150 618 -150 0 3
rlabel polysilicon 625 -150 625 -150 0 3
rlabel polysilicon 628 -150 628 -150 0 4
rlabel polysilicon 16 -205 16 -205 0 1
rlabel polysilicon 16 -211 16 -211 0 3
rlabel polysilicon 23 -205 23 -205 0 1
rlabel polysilicon 23 -211 23 -211 0 3
rlabel polysilicon 30 -205 30 -205 0 1
rlabel polysilicon 30 -211 30 -211 0 3
rlabel polysilicon 37 -205 37 -205 0 1
rlabel polysilicon 37 -211 37 -211 0 3
rlabel polysilicon 44 -205 44 -205 0 1
rlabel polysilicon 44 -211 44 -211 0 3
rlabel polysilicon 51 -205 51 -205 0 1
rlabel polysilicon 51 -211 51 -211 0 3
rlabel polysilicon 58 -205 58 -205 0 1
rlabel polysilicon 58 -211 58 -211 0 3
rlabel polysilicon 65 -205 65 -205 0 1
rlabel polysilicon 65 -211 65 -211 0 3
rlabel polysilicon 75 -211 75 -211 0 4
rlabel polysilicon 79 -205 79 -205 0 1
rlabel polysilicon 79 -211 79 -211 0 3
rlabel polysilicon 86 -205 86 -205 0 1
rlabel polysilicon 86 -211 86 -211 0 3
rlabel polysilicon 93 -205 93 -205 0 1
rlabel polysilicon 96 -205 96 -205 0 2
rlabel polysilicon 96 -211 96 -211 0 4
rlabel polysilicon 100 -205 100 -205 0 1
rlabel polysilicon 107 -205 107 -205 0 1
rlabel polysilicon 107 -211 107 -211 0 3
rlabel polysilicon 114 -205 114 -205 0 1
rlabel polysilicon 114 -211 114 -211 0 3
rlabel polysilicon 121 -205 121 -205 0 1
rlabel polysilicon 121 -211 121 -211 0 3
rlabel polysilicon 128 -205 128 -205 0 1
rlabel polysilicon 128 -211 128 -211 0 3
rlabel polysilicon 135 -205 135 -205 0 1
rlabel polysilicon 138 -205 138 -205 0 2
rlabel polysilicon 135 -211 135 -211 0 3
rlabel polysilicon 142 -205 142 -205 0 1
rlabel polysilicon 142 -211 142 -211 0 3
rlabel polysilicon 149 -205 149 -205 0 1
rlabel polysilicon 149 -211 149 -211 0 3
rlabel polysilicon 156 -205 156 -205 0 1
rlabel polysilicon 156 -211 156 -211 0 3
rlabel polysilicon 163 -205 163 -205 0 1
rlabel polysilicon 163 -211 163 -211 0 3
rlabel polysilicon 170 -205 170 -205 0 1
rlabel polysilicon 170 -211 170 -211 0 3
rlabel polysilicon 177 -205 177 -205 0 1
rlabel polysilicon 180 -205 180 -205 0 2
rlabel polysilicon 177 -211 177 -211 0 3
rlabel polysilicon 180 -211 180 -211 0 4
rlabel polysilicon 184 -205 184 -205 0 1
rlabel polysilicon 184 -211 184 -211 0 3
rlabel polysilicon 191 -205 191 -205 0 1
rlabel polysilicon 191 -211 191 -211 0 3
rlabel polysilicon 198 -205 198 -205 0 1
rlabel polysilicon 198 -211 198 -211 0 3
rlabel polysilicon 208 -205 208 -205 0 2
rlabel polysilicon 212 -205 212 -205 0 1
rlabel polysilicon 215 -205 215 -205 0 2
rlabel polysilicon 219 -205 219 -205 0 1
rlabel polysilicon 219 -211 219 -211 0 3
rlabel polysilicon 226 -205 226 -205 0 1
rlabel polysilicon 226 -211 226 -211 0 3
rlabel polysilicon 233 -205 233 -205 0 1
rlabel polysilicon 233 -211 233 -211 0 3
rlabel polysilicon 240 -205 240 -205 0 1
rlabel polysilicon 240 -211 240 -211 0 3
rlabel polysilicon 247 -205 247 -205 0 1
rlabel polysilicon 247 -211 247 -211 0 3
rlabel polysilicon 254 -205 254 -205 0 1
rlabel polysilicon 254 -211 254 -211 0 3
rlabel polysilicon 261 -205 261 -205 0 1
rlabel polysilicon 261 -211 261 -211 0 3
rlabel polysilicon 268 -205 268 -205 0 1
rlabel polysilicon 268 -211 268 -211 0 3
rlabel polysilicon 278 -205 278 -205 0 2
rlabel polysilicon 275 -211 275 -211 0 3
rlabel polysilicon 278 -211 278 -211 0 4
rlabel polysilicon 282 -205 282 -205 0 1
rlabel polysilicon 282 -211 282 -211 0 3
rlabel polysilicon 289 -205 289 -205 0 1
rlabel polysilicon 289 -211 289 -211 0 3
rlabel polysilicon 296 -205 296 -205 0 1
rlabel polysilicon 299 -205 299 -205 0 2
rlabel polysilicon 299 -211 299 -211 0 4
rlabel polysilicon 306 -205 306 -205 0 2
rlabel polysilicon 310 -205 310 -205 0 1
rlabel polysilicon 310 -211 310 -211 0 3
rlabel polysilicon 317 -205 317 -205 0 1
rlabel polysilicon 317 -211 317 -211 0 3
rlabel polysilicon 327 -211 327 -211 0 4
rlabel polysilicon 331 -205 331 -205 0 1
rlabel polysilicon 334 -205 334 -205 0 2
rlabel polysilicon 331 -211 331 -211 0 3
rlabel polysilicon 341 -205 341 -205 0 2
rlabel polysilicon 341 -211 341 -211 0 4
rlabel polysilicon 345 -205 345 -205 0 1
rlabel polysilicon 345 -211 345 -211 0 3
rlabel polysilicon 352 -205 352 -205 0 1
rlabel polysilicon 352 -211 352 -211 0 3
rlabel polysilicon 359 -205 359 -205 0 1
rlabel polysilicon 359 -211 359 -211 0 3
rlabel polysilicon 369 -205 369 -205 0 2
rlabel polysilicon 366 -211 366 -211 0 3
rlabel polysilicon 369 -211 369 -211 0 4
rlabel polysilicon 373 -205 373 -205 0 1
rlabel polysilicon 373 -211 373 -211 0 3
rlabel polysilicon 380 -205 380 -205 0 1
rlabel polysilicon 380 -211 380 -211 0 3
rlabel polysilicon 387 -205 387 -205 0 1
rlabel polysilicon 390 -205 390 -205 0 2
rlabel polysilicon 387 -211 387 -211 0 3
rlabel polysilicon 394 -205 394 -205 0 1
rlabel polysilicon 394 -211 394 -211 0 3
rlabel polysilicon 401 -205 401 -205 0 1
rlabel polysilicon 401 -211 401 -211 0 3
rlabel polysilicon 408 -205 408 -205 0 1
rlabel polysilicon 408 -211 408 -211 0 3
rlabel polysilicon 415 -205 415 -205 0 1
rlabel polysilicon 415 -211 415 -211 0 3
rlabel polysilicon 422 -205 422 -205 0 1
rlabel polysilicon 422 -211 422 -211 0 3
rlabel polysilicon 429 -205 429 -205 0 1
rlabel polysilicon 429 -211 429 -211 0 3
rlabel polysilicon 436 -205 436 -205 0 1
rlabel polysilicon 436 -211 436 -211 0 3
rlabel polysilicon 443 -211 443 -211 0 3
rlabel polysilicon 446 -211 446 -211 0 4
rlabel polysilicon 450 -205 450 -205 0 1
rlabel polysilicon 450 -211 450 -211 0 3
rlabel polysilicon 457 -205 457 -205 0 1
rlabel polysilicon 457 -211 457 -211 0 3
rlabel polysilicon 464 -205 464 -205 0 1
rlabel polysilicon 464 -211 464 -211 0 3
rlabel polysilicon 471 -205 471 -205 0 1
rlabel polysilicon 471 -211 471 -211 0 3
rlabel polysilicon 478 -205 478 -205 0 1
rlabel polysilicon 478 -211 478 -211 0 3
rlabel polysilicon 488 -205 488 -205 0 2
rlabel polysilicon 488 -211 488 -211 0 4
rlabel polysilicon 492 -205 492 -205 0 1
rlabel polysilicon 492 -211 492 -211 0 3
rlabel polysilicon 499 -205 499 -205 0 1
rlabel polysilicon 499 -211 499 -211 0 3
rlabel polysilicon 506 -205 506 -205 0 1
rlabel polysilicon 506 -211 506 -211 0 3
rlabel polysilicon 513 -205 513 -205 0 1
rlabel polysilicon 513 -211 513 -211 0 3
rlabel polysilicon 520 -205 520 -205 0 1
rlabel polysilicon 520 -211 520 -211 0 3
rlabel polysilicon 527 -205 527 -205 0 1
rlabel polysilicon 527 -211 527 -211 0 3
rlabel polysilicon 534 -205 534 -205 0 1
rlabel polysilicon 534 -211 534 -211 0 3
rlabel polysilicon 541 -205 541 -205 0 1
rlabel polysilicon 541 -211 541 -211 0 3
rlabel polysilicon 548 -205 548 -205 0 1
rlabel polysilicon 548 -211 548 -211 0 3
rlabel polysilicon 555 -205 555 -205 0 1
rlabel polysilicon 555 -211 555 -211 0 3
rlabel polysilicon 562 -205 562 -205 0 1
rlabel polysilicon 562 -211 562 -211 0 3
rlabel polysilicon 569 -205 569 -205 0 1
rlabel polysilicon 569 -211 569 -211 0 3
rlabel polysilicon 576 -205 576 -205 0 1
rlabel polysilicon 576 -211 576 -211 0 3
rlabel polysilicon 583 -205 583 -205 0 1
rlabel polysilicon 583 -211 583 -211 0 3
rlabel polysilicon 590 -205 590 -205 0 1
rlabel polysilicon 590 -211 590 -211 0 3
rlabel polysilicon 597 -205 597 -205 0 1
rlabel polysilicon 597 -211 597 -211 0 3
rlabel polysilicon 604 -205 604 -205 0 1
rlabel polysilicon 604 -211 604 -211 0 3
rlabel polysilicon 611 -205 611 -205 0 1
rlabel polysilicon 611 -211 611 -211 0 3
rlabel polysilicon 618 -205 618 -205 0 1
rlabel polysilicon 618 -211 618 -211 0 3
rlabel polysilicon 625 -205 625 -205 0 1
rlabel polysilicon 625 -211 625 -211 0 3
rlabel polysilicon 632 -205 632 -205 0 1
rlabel polysilicon 632 -211 632 -211 0 3
rlabel polysilicon 639 -205 639 -205 0 1
rlabel polysilicon 639 -211 639 -211 0 3
rlabel polysilicon 646 -205 646 -205 0 1
rlabel polysilicon 646 -211 646 -211 0 3
rlabel polysilicon 653 -205 653 -205 0 1
rlabel polysilicon 653 -211 653 -211 0 3
rlabel polysilicon 660 -205 660 -205 0 1
rlabel polysilicon 660 -211 660 -211 0 3
rlabel polysilicon 667 -205 667 -205 0 1
rlabel polysilicon 667 -211 667 -211 0 3
rlabel polysilicon 674 -205 674 -205 0 1
rlabel polysilicon 674 -211 674 -211 0 3
rlabel polysilicon 2 -270 2 -270 0 1
rlabel polysilicon 2 -276 2 -276 0 3
rlabel polysilicon 9 -270 9 -270 0 1
rlabel polysilicon 16 -270 16 -270 0 1
rlabel polysilicon 16 -276 16 -276 0 3
rlabel polysilicon 23 -270 23 -270 0 1
rlabel polysilicon 23 -276 23 -276 0 3
rlabel polysilicon 30 -270 30 -270 0 1
rlabel polysilicon 33 -270 33 -270 0 2
rlabel polysilicon 33 -276 33 -276 0 4
rlabel polysilicon 37 -270 37 -270 0 1
rlabel polysilicon 37 -276 37 -276 0 3
rlabel polysilicon 44 -270 44 -270 0 1
rlabel polysilicon 44 -276 44 -276 0 3
rlabel polysilicon 51 -270 51 -270 0 1
rlabel polysilicon 54 -270 54 -270 0 2
rlabel polysilicon 51 -276 51 -276 0 3
rlabel polysilicon 54 -276 54 -276 0 4
rlabel polysilicon 58 -270 58 -270 0 1
rlabel polysilicon 58 -276 58 -276 0 3
rlabel polysilicon 65 -270 65 -270 0 1
rlabel polysilicon 65 -276 65 -276 0 3
rlabel polysilicon 72 -270 72 -270 0 1
rlabel polysilicon 72 -276 72 -276 0 3
rlabel polysilicon 79 -270 79 -270 0 1
rlabel polysilicon 82 -270 82 -270 0 2
rlabel polysilicon 82 -276 82 -276 0 4
rlabel polysilicon 86 -270 86 -270 0 1
rlabel polysilicon 86 -276 86 -276 0 3
rlabel polysilicon 93 -270 93 -270 0 1
rlabel polysilicon 93 -276 93 -276 0 3
rlabel polysilicon 100 -270 100 -270 0 1
rlabel polysilicon 103 -270 103 -270 0 2
rlabel polysilicon 107 -270 107 -270 0 1
rlabel polysilicon 107 -276 107 -276 0 3
rlabel polysilicon 110 -276 110 -276 0 4
rlabel polysilicon 117 -270 117 -270 0 2
rlabel polysilicon 114 -276 114 -276 0 3
rlabel polysilicon 121 -270 121 -270 0 1
rlabel polysilicon 121 -276 121 -276 0 3
rlabel polysilicon 128 -270 128 -270 0 1
rlabel polysilicon 128 -276 128 -276 0 3
rlabel polysilicon 135 -270 135 -270 0 1
rlabel polysilicon 135 -276 135 -276 0 3
rlabel polysilicon 142 -270 142 -270 0 1
rlabel polysilicon 142 -276 142 -276 0 3
rlabel polysilicon 152 -270 152 -270 0 2
rlabel polysilicon 156 -270 156 -270 0 1
rlabel polysilicon 156 -276 156 -276 0 3
rlabel polysilicon 163 -270 163 -270 0 1
rlabel polysilicon 163 -276 163 -276 0 3
rlabel polysilicon 170 -270 170 -270 0 1
rlabel polysilicon 170 -276 170 -276 0 3
rlabel polysilicon 177 -270 177 -270 0 1
rlabel polysilicon 177 -276 177 -276 0 3
rlabel polysilicon 184 -270 184 -270 0 1
rlabel polysilicon 184 -276 184 -276 0 3
rlabel polysilicon 191 -270 191 -270 0 1
rlabel polysilicon 191 -276 191 -276 0 3
rlabel polysilicon 198 -270 198 -270 0 1
rlabel polysilicon 198 -276 198 -276 0 3
rlabel polysilicon 205 -270 205 -270 0 1
rlabel polysilicon 205 -276 205 -276 0 3
rlabel polysilicon 212 -270 212 -270 0 1
rlabel polysilicon 212 -276 212 -276 0 3
rlabel polysilicon 219 -270 219 -270 0 1
rlabel polysilicon 219 -276 219 -276 0 3
rlabel polysilicon 226 -270 226 -270 0 1
rlabel polysilicon 226 -276 226 -276 0 3
rlabel polysilicon 233 -270 233 -270 0 1
rlabel polysilicon 233 -276 233 -276 0 3
rlabel polysilicon 243 -270 243 -270 0 2
rlabel polysilicon 240 -276 240 -276 0 3
rlabel polysilicon 247 -270 247 -270 0 1
rlabel polysilicon 250 -270 250 -270 0 2
rlabel polysilicon 247 -276 247 -276 0 3
rlabel polysilicon 250 -276 250 -276 0 4
rlabel polysilicon 254 -270 254 -270 0 1
rlabel polysilicon 254 -276 254 -276 0 3
rlabel polysilicon 264 -270 264 -270 0 2
rlabel polysilicon 261 -276 261 -276 0 3
rlabel polysilicon 264 -276 264 -276 0 4
rlabel polysilicon 268 -270 268 -270 0 1
rlabel polysilicon 268 -276 268 -276 0 3
rlabel polysilicon 278 -270 278 -270 0 2
rlabel polysilicon 275 -276 275 -276 0 3
rlabel polysilicon 278 -276 278 -276 0 4
rlabel polysilicon 282 -270 282 -270 0 1
rlabel polysilicon 282 -276 282 -276 0 3
rlabel polysilicon 289 -270 289 -270 0 1
rlabel polysilicon 292 -270 292 -270 0 2
rlabel polysilicon 292 -276 292 -276 0 4
rlabel polysilicon 296 -270 296 -270 0 1
rlabel polysilicon 299 -270 299 -270 0 2
rlabel polysilicon 296 -276 296 -276 0 3
rlabel polysilicon 299 -276 299 -276 0 4
rlabel polysilicon 303 -270 303 -270 0 1
rlabel polysilicon 303 -276 303 -276 0 3
rlabel polysilicon 310 -270 310 -270 0 1
rlabel polysilicon 313 -270 313 -270 0 2
rlabel polysilicon 310 -276 310 -276 0 3
rlabel polysilicon 313 -276 313 -276 0 4
rlabel polysilicon 317 -270 317 -270 0 1
rlabel polysilicon 317 -276 317 -276 0 3
rlabel polysilicon 324 -270 324 -270 0 1
rlabel polysilicon 324 -276 324 -276 0 3
rlabel polysilicon 331 -270 331 -270 0 1
rlabel polysilicon 331 -276 331 -276 0 3
rlabel polysilicon 338 -270 338 -270 0 1
rlabel polysilicon 338 -276 338 -276 0 3
rlabel polysilicon 345 -270 345 -270 0 1
rlabel polysilicon 345 -276 345 -276 0 3
rlabel polysilicon 352 -270 352 -270 0 1
rlabel polysilicon 352 -276 352 -276 0 3
rlabel polysilicon 359 -270 359 -270 0 1
rlabel polysilicon 359 -276 359 -276 0 3
rlabel polysilicon 369 -270 369 -270 0 2
rlabel polysilicon 369 -276 369 -276 0 4
rlabel polysilicon 373 -270 373 -270 0 1
rlabel polysilicon 373 -276 373 -276 0 3
rlabel polysilicon 380 -270 380 -270 0 1
rlabel polysilicon 383 -270 383 -270 0 2
rlabel polysilicon 380 -276 380 -276 0 3
rlabel polysilicon 383 -276 383 -276 0 4
rlabel polysilicon 387 -270 387 -270 0 1
rlabel polysilicon 387 -276 387 -276 0 3
rlabel polysilicon 394 -270 394 -270 0 1
rlabel polysilicon 394 -276 394 -276 0 3
rlabel polysilicon 401 -270 401 -270 0 1
rlabel polysilicon 401 -276 401 -276 0 3
rlabel polysilicon 408 -270 408 -270 0 1
rlabel polysilicon 408 -276 408 -276 0 3
rlabel polysilicon 415 -270 415 -270 0 1
rlabel polysilicon 415 -276 415 -276 0 3
rlabel polysilicon 422 -270 422 -270 0 1
rlabel polysilicon 422 -276 422 -276 0 3
rlabel polysilicon 429 -270 429 -270 0 1
rlabel polysilicon 429 -276 429 -276 0 3
rlabel polysilicon 436 -270 436 -270 0 1
rlabel polysilicon 436 -276 436 -276 0 3
rlabel polysilicon 443 -270 443 -270 0 1
rlabel polysilicon 443 -276 443 -276 0 3
rlabel polysilicon 450 -270 450 -270 0 1
rlabel polysilicon 450 -276 450 -276 0 3
rlabel polysilicon 457 -270 457 -270 0 1
rlabel polysilicon 457 -276 457 -276 0 3
rlabel polysilicon 467 -276 467 -276 0 4
rlabel polysilicon 471 -270 471 -270 0 1
rlabel polysilicon 471 -276 471 -276 0 3
rlabel polysilicon 478 -270 478 -270 0 1
rlabel polysilicon 478 -276 478 -276 0 3
rlabel polysilicon 485 -270 485 -270 0 1
rlabel polysilicon 485 -276 485 -276 0 3
rlabel polysilicon 492 -270 492 -270 0 1
rlabel polysilicon 492 -276 492 -276 0 3
rlabel polysilicon 499 -270 499 -270 0 1
rlabel polysilicon 499 -276 499 -276 0 3
rlabel polysilicon 506 -270 506 -270 0 1
rlabel polysilicon 506 -276 506 -276 0 3
rlabel polysilicon 513 -270 513 -270 0 1
rlabel polysilicon 513 -276 513 -276 0 3
rlabel polysilicon 520 -270 520 -270 0 1
rlabel polysilicon 520 -276 520 -276 0 3
rlabel polysilicon 527 -270 527 -270 0 1
rlabel polysilicon 527 -276 527 -276 0 3
rlabel polysilicon 534 -270 534 -270 0 1
rlabel polysilicon 534 -276 534 -276 0 3
rlabel polysilicon 541 -270 541 -270 0 1
rlabel polysilicon 541 -276 541 -276 0 3
rlabel polysilicon 548 -270 548 -270 0 1
rlabel polysilicon 548 -276 548 -276 0 3
rlabel polysilicon 555 -270 555 -270 0 1
rlabel polysilicon 555 -276 555 -276 0 3
rlabel polysilicon 562 -270 562 -270 0 1
rlabel polysilicon 562 -276 562 -276 0 3
rlabel polysilicon 569 -270 569 -270 0 1
rlabel polysilicon 569 -276 569 -276 0 3
rlabel polysilicon 576 -270 576 -270 0 1
rlabel polysilicon 576 -276 576 -276 0 3
rlabel polysilicon 583 -270 583 -270 0 1
rlabel polysilicon 583 -276 583 -276 0 3
rlabel polysilicon 590 -270 590 -270 0 1
rlabel polysilicon 590 -276 590 -276 0 3
rlabel polysilicon 597 -270 597 -270 0 1
rlabel polysilicon 597 -276 597 -276 0 3
rlabel polysilicon 604 -270 604 -270 0 1
rlabel polysilicon 604 -276 604 -276 0 3
rlabel polysilicon 611 -270 611 -270 0 1
rlabel polysilicon 611 -276 611 -276 0 3
rlabel polysilicon 618 -270 618 -270 0 1
rlabel polysilicon 618 -276 618 -276 0 3
rlabel polysilicon 625 -270 625 -270 0 1
rlabel polysilicon 625 -276 625 -276 0 3
rlabel polysilicon 632 -270 632 -270 0 1
rlabel polysilicon 632 -276 632 -276 0 3
rlabel polysilicon 639 -270 639 -270 0 1
rlabel polysilicon 639 -276 639 -276 0 3
rlabel polysilicon 646 -270 646 -270 0 1
rlabel polysilicon 646 -276 646 -276 0 3
rlabel polysilicon 653 -270 653 -270 0 1
rlabel polysilicon 653 -276 653 -276 0 3
rlabel polysilicon 660 -270 660 -270 0 1
rlabel polysilicon 660 -276 660 -276 0 3
rlabel polysilicon 667 -270 667 -270 0 1
rlabel polysilicon 667 -276 667 -276 0 3
rlabel polysilicon 674 -270 674 -270 0 1
rlabel polysilicon 674 -276 674 -276 0 3
rlabel polysilicon 681 -270 681 -270 0 1
rlabel polysilicon 681 -276 681 -276 0 3
rlabel polysilicon 688 -270 688 -270 0 1
rlabel polysilicon 688 -276 688 -276 0 3
rlabel polysilicon 695 -270 695 -270 0 1
rlabel polysilicon 695 -276 695 -276 0 3
rlabel polysilicon 702 -270 702 -270 0 1
rlabel polysilicon 702 -276 702 -276 0 3
rlabel polysilicon 712 -270 712 -270 0 2
rlabel polysilicon 709 -276 709 -276 0 3
rlabel polysilicon 716 -270 716 -270 0 1
rlabel polysilicon 716 -276 716 -276 0 3
rlabel polysilicon 723 -270 723 -270 0 1
rlabel polysilicon 723 -276 723 -276 0 3
rlabel polysilicon 730 -270 730 -270 0 1
rlabel polysilicon 16 -337 16 -337 0 1
rlabel polysilicon 16 -343 16 -343 0 3
rlabel polysilicon 26 -337 26 -337 0 2
rlabel polysilicon 26 -343 26 -343 0 4
rlabel polysilicon 30 -337 30 -337 0 1
rlabel polysilicon 30 -343 30 -343 0 3
rlabel polysilicon 37 -337 37 -337 0 1
rlabel polysilicon 37 -343 37 -343 0 3
rlabel polysilicon 44 -337 44 -337 0 1
rlabel polysilicon 47 -337 47 -337 0 2
rlabel polysilicon 47 -343 47 -343 0 4
rlabel polysilicon 51 -337 51 -337 0 1
rlabel polysilicon 54 -337 54 -337 0 2
rlabel polysilicon 54 -343 54 -343 0 4
rlabel polysilicon 58 -337 58 -337 0 1
rlabel polysilicon 58 -343 58 -343 0 3
rlabel polysilicon 61 -343 61 -343 0 4
rlabel polysilicon 65 -337 65 -337 0 1
rlabel polysilicon 65 -343 65 -343 0 3
rlabel polysilicon 72 -337 72 -337 0 1
rlabel polysilicon 72 -343 72 -343 0 3
rlabel polysilicon 79 -337 79 -337 0 1
rlabel polysilicon 79 -343 79 -343 0 3
rlabel polysilicon 86 -337 86 -337 0 1
rlabel polysilicon 86 -343 86 -343 0 3
rlabel polysilicon 93 -337 93 -337 0 1
rlabel polysilicon 93 -343 93 -343 0 3
rlabel polysilicon 100 -337 100 -337 0 1
rlabel polysilicon 100 -343 100 -343 0 3
rlabel polysilicon 110 -337 110 -337 0 2
rlabel polysilicon 110 -343 110 -343 0 4
rlabel polysilicon 114 -337 114 -337 0 1
rlabel polysilicon 114 -343 114 -343 0 3
rlabel polysilicon 121 -337 121 -337 0 1
rlabel polysilicon 121 -343 121 -343 0 3
rlabel polysilicon 128 -337 128 -337 0 1
rlabel polysilicon 128 -343 128 -343 0 3
rlabel polysilicon 135 -337 135 -337 0 1
rlabel polysilicon 135 -343 135 -343 0 3
rlabel polysilicon 142 -337 142 -337 0 1
rlabel polysilicon 142 -343 142 -343 0 3
rlabel polysilicon 149 -337 149 -337 0 1
rlabel polysilicon 149 -343 149 -343 0 3
rlabel polysilicon 156 -337 156 -337 0 1
rlabel polysilicon 156 -343 156 -343 0 3
rlabel polysilicon 163 -343 163 -343 0 3
rlabel polysilicon 170 -337 170 -337 0 1
rlabel polysilicon 170 -343 170 -343 0 3
rlabel polysilicon 177 -337 177 -337 0 1
rlabel polysilicon 177 -343 177 -343 0 3
rlabel polysilicon 184 -337 184 -337 0 1
rlabel polysilicon 187 -337 187 -337 0 2
rlabel polysilicon 187 -343 187 -343 0 4
rlabel polysilicon 191 -337 191 -337 0 1
rlabel polysilicon 191 -343 191 -343 0 3
rlabel polysilicon 198 -337 198 -337 0 1
rlabel polysilicon 198 -343 198 -343 0 3
rlabel polysilicon 205 -337 205 -337 0 1
rlabel polysilicon 205 -343 205 -343 0 3
rlabel polysilicon 212 -337 212 -337 0 1
rlabel polysilicon 212 -343 212 -343 0 3
rlabel polysilicon 219 -337 219 -337 0 1
rlabel polysilicon 219 -343 219 -343 0 3
rlabel polysilicon 226 -337 226 -337 0 1
rlabel polysilicon 226 -343 226 -343 0 3
rlabel polysilicon 229 -343 229 -343 0 4
rlabel polysilicon 233 -337 233 -337 0 1
rlabel polysilicon 233 -343 233 -343 0 3
rlabel polysilicon 240 -337 240 -337 0 1
rlabel polysilicon 240 -343 240 -343 0 3
rlabel polysilicon 247 -337 247 -337 0 1
rlabel polysilicon 247 -343 247 -343 0 3
rlabel polysilicon 257 -337 257 -337 0 2
rlabel polysilicon 254 -343 254 -343 0 3
rlabel polysilicon 261 -337 261 -337 0 1
rlabel polysilicon 261 -343 261 -343 0 3
rlabel polysilicon 268 -337 268 -337 0 1
rlabel polysilicon 268 -343 268 -343 0 3
rlabel polysilicon 275 -337 275 -337 0 1
rlabel polysilicon 278 -337 278 -337 0 2
rlabel polysilicon 278 -343 278 -343 0 4
rlabel polysilicon 282 -337 282 -337 0 1
rlabel polysilicon 282 -343 282 -343 0 3
rlabel polysilicon 285 -343 285 -343 0 4
rlabel polysilicon 289 -337 289 -337 0 1
rlabel polysilicon 289 -343 289 -343 0 3
rlabel polysilicon 299 -337 299 -337 0 2
rlabel polysilicon 296 -343 296 -343 0 3
rlabel polysilicon 299 -343 299 -343 0 4
rlabel polysilicon 303 -337 303 -337 0 1
rlabel polysilicon 303 -343 303 -343 0 3
rlabel polysilicon 310 -337 310 -337 0 1
rlabel polysilicon 310 -343 310 -343 0 3
rlabel polysilicon 317 -337 317 -337 0 1
rlabel polysilicon 317 -343 317 -343 0 3
rlabel polysilicon 324 -337 324 -337 0 1
rlabel polysilicon 327 -337 327 -337 0 2
rlabel polysilicon 331 -337 331 -337 0 1
rlabel polysilicon 331 -343 331 -343 0 3
rlabel polysilicon 338 -337 338 -337 0 1
rlabel polysilicon 338 -343 338 -343 0 3
rlabel polysilicon 345 -337 345 -337 0 1
rlabel polysilicon 348 -337 348 -337 0 2
rlabel polysilicon 345 -343 345 -343 0 3
rlabel polysilicon 348 -343 348 -343 0 4
rlabel polysilicon 352 -337 352 -337 0 1
rlabel polysilicon 352 -343 352 -343 0 3
rlabel polysilicon 362 -337 362 -337 0 2
rlabel polysilicon 366 -343 366 -343 0 3
rlabel polysilicon 369 -343 369 -343 0 4
rlabel polysilicon 373 -337 373 -337 0 1
rlabel polysilicon 373 -343 373 -343 0 3
rlabel polysilicon 380 -337 380 -337 0 1
rlabel polysilicon 380 -343 380 -343 0 3
rlabel polysilicon 387 -337 387 -337 0 1
rlabel polysilicon 387 -343 387 -343 0 3
rlabel polysilicon 394 -337 394 -337 0 1
rlabel polysilicon 394 -343 394 -343 0 3
rlabel polysilicon 401 -337 401 -337 0 1
rlabel polysilicon 401 -343 401 -343 0 3
rlabel polysilicon 408 -337 408 -337 0 1
rlabel polysilicon 408 -343 408 -343 0 3
rlabel polysilicon 415 -337 415 -337 0 1
rlabel polysilicon 415 -343 415 -343 0 3
rlabel polysilicon 422 -337 422 -337 0 1
rlabel polysilicon 422 -343 422 -343 0 3
rlabel polysilicon 429 -337 429 -337 0 1
rlabel polysilicon 432 -337 432 -337 0 2
rlabel polysilicon 429 -343 429 -343 0 3
rlabel polysilicon 436 -337 436 -337 0 1
rlabel polysilicon 436 -343 436 -343 0 3
rlabel polysilicon 443 -337 443 -337 0 1
rlabel polysilicon 443 -343 443 -343 0 3
rlabel polysilicon 450 -337 450 -337 0 1
rlabel polysilicon 450 -343 450 -343 0 3
rlabel polysilicon 457 -337 457 -337 0 1
rlabel polysilicon 457 -343 457 -343 0 3
rlabel polysilicon 464 -337 464 -337 0 1
rlabel polysilicon 464 -343 464 -343 0 3
rlabel polysilicon 471 -337 471 -337 0 1
rlabel polysilicon 471 -343 471 -343 0 3
rlabel polysilicon 478 -337 478 -337 0 1
rlabel polysilicon 478 -343 478 -343 0 3
rlabel polysilicon 485 -337 485 -337 0 1
rlabel polysilicon 485 -343 485 -343 0 3
rlabel polysilicon 492 -337 492 -337 0 1
rlabel polysilicon 492 -343 492 -343 0 3
rlabel polysilicon 499 -337 499 -337 0 1
rlabel polysilicon 499 -343 499 -343 0 3
rlabel polysilicon 506 -337 506 -337 0 1
rlabel polysilicon 506 -343 506 -343 0 3
rlabel polysilicon 513 -337 513 -337 0 1
rlabel polysilicon 513 -343 513 -343 0 3
rlabel polysilicon 520 -337 520 -337 0 1
rlabel polysilicon 520 -343 520 -343 0 3
rlabel polysilicon 527 -337 527 -337 0 1
rlabel polysilicon 527 -343 527 -343 0 3
rlabel polysilicon 534 -337 534 -337 0 1
rlabel polysilicon 534 -343 534 -343 0 3
rlabel polysilicon 541 -337 541 -337 0 1
rlabel polysilicon 541 -343 541 -343 0 3
rlabel polysilicon 548 -337 548 -337 0 1
rlabel polysilicon 548 -343 548 -343 0 3
rlabel polysilicon 555 -337 555 -337 0 1
rlabel polysilicon 555 -343 555 -343 0 3
rlabel polysilicon 562 -337 562 -337 0 1
rlabel polysilicon 562 -343 562 -343 0 3
rlabel polysilicon 569 -337 569 -337 0 1
rlabel polysilicon 569 -343 569 -343 0 3
rlabel polysilicon 576 -337 576 -337 0 1
rlabel polysilicon 576 -343 576 -343 0 3
rlabel polysilicon 583 -337 583 -337 0 1
rlabel polysilicon 583 -343 583 -343 0 3
rlabel polysilicon 590 -337 590 -337 0 1
rlabel polysilicon 590 -343 590 -343 0 3
rlabel polysilicon 597 -337 597 -337 0 1
rlabel polysilicon 597 -343 597 -343 0 3
rlabel polysilicon 604 -337 604 -337 0 1
rlabel polysilicon 604 -343 604 -343 0 3
rlabel polysilicon 611 -337 611 -337 0 1
rlabel polysilicon 611 -343 611 -343 0 3
rlabel polysilicon 618 -337 618 -337 0 1
rlabel polysilicon 618 -343 618 -343 0 3
rlabel polysilicon 625 -337 625 -337 0 1
rlabel polysilicon 625 -343 625 -343 0 3
rlabel polysilicon 632 -337 632 -337 0 1
rlabel polysilicon 632 -343 632 -343 0 3
rlabel polysilicon 639 -337 639 -337 0 1
rlabel polysilicon 639 -343 639 -343 0 3
rlabel polysilicon 646 -337 646 -337 0 1
rlabel polysilicon 646 -343 646 -343 0 3
rlabel polysilicon 653 -337 653 -337 0 1
rlabel polysilicon 653 -343 653 -343 0 3
rlabel polysilicon 660 -337 660 -337 0 1
rlabel polysilicon 660 -343 660 -343 0 3
rlabel polysilicon 667 -337 667 -337 0 1
rlabel polysilicon 667 -343 667 -343 0 3
rlabel polysilicon 674 -337 674 -337 0 1
rlabel polysilicon 674 -343 674 -343 0 3
rlabel polysilicon 681 -337 681 -337 0 1
rlabel polysilicon 681 -343 681 -343 0 3
rlabel polysilicon 688 -337 688 -337 0 1
rlabel polysilicon 688 -343 688 -343 0 3
rlabel polysilicon 695 -337 695 -337 0 1
rlabel polysilicon 695 -343 695 -343 0 3
rlabel polysilicon 702 -337 702 -337 0 1
rlabel polysilicon 702 -343 702 -343 0 3
rlabel polysilicon 709 -337 709 -337 0 1
rlabel polysilicon 709 -343 709 -343 0 3
rlabel polysilicon 716 -337 716 -337 0 1
rlabel polysilicon 716 -343 716 -343 0 3
rlabel polysilicon 723 -337 723 -337 0 1
rlabel polysilicon 723 -343 723 -343 0 3
rlabel polysilicon 730 -337 730 -337 0 1
rlabel polysilicon 730 -343 730 -343 0 3
rlabel polysilicon 737 -337 737 -337 0 1
rlabel polysilicon 737 -343 737 -343 0 3
rlabel polysilicon 2 -416 2 -416 0 1
rlabel polysilicon 5 -416 5 -416 0 2
rlabel polysilicon 9 -422 9 -422 0 3
rlabel polysilicon 16 -416 16 -416 0 1
rlabel polysilicon 16 -422 16 -422 0 3
rlabel polysilicon 23 -416 23 -416 0 1
rlabel polysilicon 23 -422 23 -422 0 3
rlabel polysilicon 30 -416 30 -416 0 1
rlabel polysilicon 30 -422 30 -422 0 3
rlabel polysilicon 37 -416 37 -416 0 1
rlabel polysilicon 37 -422 37 -422 0 3
rlabel polysilicon 44 -416 44 -416 0 1
rlabel polysilicon 44 -422 44 -422 0 3
rlabel polysilicon 51 -416 51 -416 0 1
rlabel polysilicon 51 -422 51 -422 0 3
rlabel polysilicon 58 -422 58 -422 0 3
rlabel polysilicon 65 -416 65 -416 0 1
rlabel polysilicon 65 -422 65 -422 0 3
rlabel polysilicon 72 -416 72 -416 0 1
rlabel polysilicon 72 -422 72 -422 0 3
rlabel polysilicon 79 -416 79 -416 0 1
rlabel polysilicon 79 -422 79 -422 0 3
rlabel polysilicon 86 -416 86 -416 0 1
rlabel polysilicon 86 -422 86 -422 0 3
rlabel polysilicon 93 -416 93 -416 0 1
rlabel polysilicon 93 -422 93 -422 0 3
rlabel polysilicon 100 -416 100 -416 0 1
rlabel polysilicon 100 -422 100 -422 0 3
rlabel polysilicon 107 -416 107 -416 0 1
rlabel polysilicon 110 -416 110 -416 0 2
rlabel polysilicon 107 -422 107 -422 0 3
rlabel polysilicon 110 -422 110 -422 0 4
rlabel polysilicon 114 -416 114 -416 0 1
rlabel polysilicon 114 -422 114 -422 0 3
rlabel polysilicon 124 -416 124 -416 0 2
rlabel polysilicon 124 -422 124 -422 0 4
rlabel polysilicon 128 -416 128 -416 0 1
rlabel polysilicon 128 -422 128 -422 0 3
rlabel polysilicon 135 -416 135 -416 0 1
rlabel polysilicon 135 -422 135 -422 0 3
rlabel polysilicon 142 -416 142 -416 0 1
rlabel polysilicon 142 -422 142 -422 0 3
rlabel polysilicon 149 -416 149 -416 0 1
rlabel polysilicon 149 -422 149 -422 0 3
rlabel polysilicon 156 -416 156 -416 0 1
rlabel polysilicon 156 -422 156 -422 0 3
rlabel polysilicon 163 -416 163 -416 0 1
rlabel polysilicon 163 -422 163 -422 0 3
rlabel polysilicon 170 -416 170 -416 0 1
rlabel polysilicon 170 -422 170 -422 0 3
rlabel polysilicon 177 -416 177 -416 0 1
rlabel polysilicon 177 -422 177 -422 0 3
rlabel polysilicon 184 -416 184 -416 0 1
rlabel polysilicon 184 -422 184 -422 0 3
rlabel polysilicon 191 -416 191 -416 0 1
rlabel polysilicon 191 -422 191 -422 0 3
rlabel polysilicon 198 -416 198 -416 0 1
rlabel polysilicon 198 -422 198 -422 0 3
rlabel polysilicon 205 -416 205 -416 0 1
rlabel polysilicon 205 -422 205 -422 0 3
rlabel polysilicon 212 -416 212 -416 0 1
rlabel polysilicon 212 -422 212 -422 0 3
rlabel polysilicon 219 -416 219 -416 0 1
rlabel polysilicon 222 -416 222 -416 0 2
rlabel polysilicon 219 -422 219 -422 0 3
rlabel polysilicon 222 -422 222 -422 0 4
rlabel polysilicon 226 -416 226 -416 0 1
rlabel polysilicon 226 -422 226 -422 0 3
rlabel polysilicon 233 -416 233 -416 0 1
rlabel polysilicon 233 -422 233 -422 0 3
rlabel polysilicon 240 -416 240 -416 0 1
rlabel polysilicon 240 -422 240 -422 0 3
rlabel polysilicon 247 -416 247 -416 0 1
rlabel polysilicon 247 -422 247 -422 0 3
rlabel polysilicon 254 -416 254 -416 0 1
rlabel polysilicon 254 -422 254 -422 0 3
rlabel polysilicon 261 -416 261 -416 0 1
rlabel polysilicon 261 -422 261 -422 0 3
rlabel polysilicon 268 -416 268 -416 0 1
rlabel polysilicon 268 -422 268 -422 0 3
rlabel polysilicon 275 -416 275 -416 0 1
rlabel polysilicon 275 -422 275 -422 0 3
rlabel polysilicon 282 -416 282 -416 0 1
rlabel polysilicon 282 -422 282 -422 0 3
rlabel polysilicon 289 -416 289 -416 0 1
rlabel polysilicon 292 -416 292 -416 0 2
rlabel polysilicon 296 -416 296 -416 0 1
rlabel polysilicon 296 -422 296 -422 0 3
rlabel polysilicon 303 -416 303 -416 0 1
rlabel polysilicon 303 -422 303 -422 0 3
rlabel polysilicon 310 -416 310 -416 0 1
rlabel polysilicon 310 -422 310 -422 0 3
rlabel polysilicon 317 -416 317 -416 0 1
rlabel polysilicon 317 -422 317 -422 0 3
rlabel polysilicon 324 -416 324 -416 0 1
rlabel polysilicon 324 -422 324 -422 0 3
rlabel polysilicon 331 -416 331 -416 0 1
rlabel polysilicon 334 -416 334 -416 0 2
rlabel polysilicon 331 -422 331 -422 0 3
rlabel polysilicon 334 -422 334 -422 0 4
rlabel polysilicon 338 -416 338 -416 0 1
rlabel polysilicon 341 -416 341 -416 0 2
rlabel polysilicon 338 -422 338 -422 0 3
rlabel polysilicon 345 -416 345 -416 0 1
rlabel polysilicon 348 -416 348 -416 0 2
rlabel polysilicon 345 -422 345 -422 0 3
rlabel polysilicon 348 -422 348 -422 0 4
rlabel polysilicon 352 -416 352 -416 0 1
rlabel polysilicon 352 -422 352 -422 0 3
rlabel polysilicon 359 -416 359 -416 0 1
rlabel polysilicon 359 -422 359 -422 0 3
rlabel polysilicon 366 -416 366 -416 0 1
rlabel polysilicon 366 -422 366 -422 0 3
rlabel polysilicon 373 -416 373 -416 0 1
rlabel polysilicon 376 -416 376 -416 0 2
rlabel polysilicon 380 -416 380 -416 0 1
rlabel polysilicon 383 -416 383 -416 0 2
rlabel polysilicon 380 -422 380 -422 0 3
rlabel polysilicon 383 -422 383 -422 0 4
rlabel polysilicon 387 -416 387 -416 0 1
rlabel polysilicon 387 -422 387 -422 0 3
rlabel polysilicon 394 -416 394 -416 0 1
rlabel polysilicon 397 -416 397 -416 0 2
rlabel polysilicon 394 -422 394 -422 0 3
rlabel polysilicon 401 -416 401 -416 0 1
rlabel polysilicon 404 -416 404 -416 0 2
rlabel polysilicon 404 -422 404 -422 0 4
rlabel polysilicon 408 -416 408 -416 0 1
rlabel polysilicon 408 -422 408 -422 0 3
rlabel polysilicon 415 -416 415 -416 0 1
rlabel polysilicon 418 -416 418 -416 0 2
rlabel polysilicon 415 -422 415 -422 0 3
rlabel polysilicon 418 -422 418 -422 0 4
rlabel polysilicon 422 -416 422 -416 0 1
rlabel polysilicon 422 -422 422 -422 0 3
rlabel polysilicon 432 -416 432 -416 0 2
rlabel polysilicon 432 -422 432 -422 0 4
rlabel polysilicon 436 -416 436 -416 0 1
rlabel polysilicon 436 -422 436 -422 0 3
rlabel polysilicon 443 -416 443 -416 0 1
rlabel polysilicon 443 -422 443 -422 0 3
rlabel polysilicon 450 -416 450 -416 0 1
rlabel polysilicon 450 -422 450 -422 0 3
rlabel polysilicon 457 -416 457 -416 0 1
rlabel polysilicon 457 -422 457 -422 0 3
rlabel polysilicon 464 -416 464 -416 0 1
rlabel polysilicon 464 -422 464 -422 0 3
rlabel polysilicon 474 -416 474 -416 0 2
rlabel polysilicon 471 -422 471 -422 0 3
rlabel polysilicon 474 -422 474 -422 0 4
rlabel polysilicon 478 -416 478 -416 0 1
rlabel polysilicon 478 -422 478 -422 0 3
rlabel polysilicon 485 -416 485 -416 0 1
rlabel polysilicon 485 -422 485 -422 0 3
rlabel polysilicon 492 -416 492 -416 0 1
rlabel polysilicon 492 -422 492 -422 0 3
rlabel polysilicon 499 -416 499 -416 0 1
rlabel polysilicon 499 -422 499 -422 0 3
rlabel polysilicon 506 -422 506 -422 0 3
rlabel polysilicon 513 -416 513 -416 0 1
rlabel polysilicon 513 -422 513 -422 0 3
rlabel polysilicon 523 -416 523 -416 0 2
rlabel polysilicon 520 -422 520 -422 0 3
rlabel polysilicon 523 -422 523 -422 0 4
rlabel polysilicon 527 -416 527 -416 0 1
rlabel polysilicon 527 -422 527 -422 0 3
rlabel polysilicon 534 -416 534 -416 0 1
rlabel polysilicon 534 -422 534 -422 0 3
rlabel polysilicon 541 -416 541 -416 0 1
rlabel polysilicon 541 -422 541 -422 0 3
rlabel polysilicon 548 -416 548 -416 0 1
rlabel polysilicon 548 -422 548 -422 0 3
rlabel polysilicon 558 -416 558 -416 0 2
rlabel polysilicon 555 -422 555 -422 0 3
rlabel polysilicon 562 -416 562 -416 0 1
rlabel polysilicon 562 -422 562 -422 0 3
rlabel polysilicon 569 -416 569 -416 0 1
rlabel polysilicon 569 -422 569 -422 0 3
rlabel polysilicon 576 -416 576 -416 0 1
rlabel polysilicon 576 -422 576 -422 0 3
rlabel polysilicon 583 -416 583 -416 0 1
rlabel polysilicon 590 -416 590 -416 0 1
rlabel polysilicon 590 -422 590 -422 0 3
rlabel polysilicon 597 -416 597 -416 0 1
rlabel polysilicon 597 -422 597 -422 0 3
rlabel polysilicon 604 -416 604 -416 0 1
rlabel polysilicon 604 -422 604 -422 0 3
rlabel polysilicon 611 -416 611 -416 0 1
rlabel polysilicon 611 -422 611 -422 0 3
rlabel polysilicon 618 -416 618 -416 0 1
rlabel polysilicon 618 -422 618 -422 0 3
rlabel polysilicon 625 -416 625 -416 0 1
rlabel polysilicon 625 -422 625 -422 0 3
rlabel polysilicon 632 -416 632 -416 0 1
rlabel polysilicon 632 -422 632 -422 0 3
rlabel polysilicon 639 -416 639 -416 0 1
rlabel polysilicon 639 -422 639 -422 0 3
rlabel polysilicon 646 -416 646 -416 0 1
rlabel polysilicon 646 -422 646 -422 0 3
rlabel polysilicon 653 -416 653 -416 0 1
rlabel polysilicon 653 -422 653 -422 0 3
rlabel polysilicon 660 -416 660 -416 0 1
rlabel polysilicon 660 -422 660 -422 0 3
rlabel polysilicon 667 -416 667 -416 0 1
rlabel polysilicon 667 -422 667 -422 0 3
rlabel polysilicon 674 -416 674 -416 0 1
rlabel polysilicon 674 -422 674 -422 0 3
rlabel polysilicon 681 -416 681 -416 0 1
rlabel polysilicon 681 -422 681 -422 0 3
rlabel polysilicon 688 -416 688 -416 0 1
rlabel polysilicon 688 -422 688 -422 0 3
rlabel polysilicon 695 -416 695 -416 0 1
rlabel polysilicon 695 -422 695 -422 0 3
rlabel polysilicon 702 -416 702 -416 0 1
rlabel polysilicon 702 -422 702 -422 0 3
rlabel polysilicon 705 -422 705 -422 0 4
rlabel polysilicon 709 -416 709 -416 0 1
rlabel polysilicon 709 -422 709 -422 0 3
rlabel polysilicon 716 -416 716 -416 0 1
rlabel polysilicon 716 -422 716 -422 0 3
rlabel polysilicon 723 -416 723 -416 0 1
rlabel polysilicon 723 -422 723 -422 0 3
rlabel polysilicon 730 -416 730 -416 0 1
rlabel polysilicon 730 -422 730 -422 0 3
rlabel polysilicon 737 -416 737 -416 0 1
rlabel polysilicon 737 -422 737 -422 0 3
rlabel polysilicon 744 -416 744 -416 0 1
rlabel polysilicon 744 -422 744 -422 0 3
rlabel polysilicon 751 -416 751 -416 0 1
rlabel polysilicon 751 -422 751 -422 0 3
rlabel polysilicon 758 -416 758 -416 0 1
rlabel polysilicon 758 -422 758 -422 0 3
rlabel polysilicon 765 -416 765 -416 0 1
rlabel polysilicon 765 -422 765 -422 0 3
rlabel polysilicon 772 -416 772 -416 0 1
rlabel polysilicon 772 -422 772 -422 0 3
rlabel polysilicon 779 -416 779 -416 0 1
rlabel polysilicon 779 -422 779 -422 0 3
rlabel polysilicon 786 -416 786 -416 0 1
rlabel polysilicon 786 -422 786 -422 0 3
rlabel polysilicon 793 -416 793 -416 0 1
rlabel polysilicon 793 -422 793 -422 0 3
rlabel polysilicon 800 -416 800 -416 0 1
rlabel polysilicon 800 -422 800 -422 0 3
rlabel polysilicon 807 -416 807 -416 0 1
rlabel polysilicon 807 -422 807 -422 0 3
rlabel polysilicon 814 -416 814 -416 0 1
rlabel polysilicon 814 -422 814 -422 0 3
rlabel polysilicon 9 -509 9 -509 0 1
rlabel polysilicon 9 -515 9 -515 0 3
rlabel polysilicon 16 -509 16 -509 0 1
rlabel polysilicon 16 -515 16 -515 0 3
rlabel polysilicon 23 -509 23 -509 0 1
rlabel polysilicon 23 -515 23 -515 0 3
rlabel polysilicon 30 -509 30 -509 0 1
rlabel polysilicon 30 -515 30 -515 0 3
rlabel polysilicon 37 -509 37 -509 0 1
rlabel polysilicon 37 -515 37 -515 0 3
rlabel polysilicon 44 -509 44 -509 0 1
rlabel polysilicon 47 -509 47 -509 0 2
rlabel polysilicon 47 -515 47 -515 0 4
rlabel polysilicon 51 -509 51 -509 0 1
rlabel polysilicon 51 -515 51 -515 0 3
rlabel polysilicon 58 -509 58 -509 0 1
rlabel polysilicon 61 -509 61 -509 0 2
rlabel polysilicon 61 -515 61 -515 0 4
rlabel polysilicon 65 -509 65 -509 0 1
rlabel polysilicon 65 -515 65 -515 0 3
rlabel polysilicon 72 -509 72 -509 0 1
rlabel polysilicon 72 -515 72 -515 0 3
rlabel polysilicon 79 -509 79 -509 0 1
rlabel polysilicon 79 -515 79 -515 0 3
rlabel polysilicon 86 -509 86 -509 0 1
rlabel polysilicon 86 -515 86 -515 0 3
rlabel polysilicon 93 -509 93 -509 0 1
rlabel polysilicon 93 -515 93 -515 0 3
rlabel polysilicon 100 -509 100 -509 0 1
rlabel polysilicon 100 -515 100 -515 0 3
rlabel polysilicon 103 -515 103 -515 0 4
rlabel polysilicon 107 -509 107 -509 0 1
rlabel polysilicon 107 -515 107 -515 0 3
rlabel polysilicon 114 -509 114 -509 0 1
rlabel polysilicon 114 -515 114 -515 0 3
rlabel polysilicon 121 -509 121 -509 0 1
rlabel polysilicon 121 -515 121 -515 0 3
rlabel polysilicon 128 -509 128 -509 0 1
rlabel polysilicon 128 -515 128 -515 0 3
rlabel polysilicon 138 -509 138 -509 0 2
rlabel polysilicon 135 -515 135 -515 0 3
rlabel polysilicon 142 -509 142 -509 0 1
rlabel polysilicon 142 -515 142 -515 0 3
rlabel polysilicon 149 -509 149 -509 0 1
rlabel polysilicon 149 -515 149 -515 0 3
rlabel polysilicon 156 -509 156 -509 0 1
rlabel polysilicon 156 -515 156 -515 0 3
rlabel polysilicon 163 -509 163 -509 0 1
rlabel polysilicon 163 -515 163 -515 0 3
rlabel polysilicon 170 -509 170 -509 0 1
rlabel polysilicon 170 -515 170 -515 0 3
rlabel polysilicon 177 -509 177 -509 0 1
rlabel polysilicon 177 -515 177 -515 0 3
rlabel polysilicon 184 -509 184 -509 0 1
rlabel polysilicon 184 -515 184 -515 0 3
rlabel polysilicon 191 -509 191 -509 0 1
rlabel polysilicon 191 -515 191 -515 0 3
rlabel polysilicon 198 -509 198 -509 0 1
rlabel polysilicon 198 -515 198 -515 0 3
rlabel polysilicon 205 -509 205 -509 0 1
rlabel polysilicon 205 -515 205 -515 0 3
rlabel polysilicon 212 -509 212 -509 0 1
rlabel polysilicon 212 -515 212 -515 0 3
rlabel polysilicon 222 -509 222 -509 0 2
rlabel polysilicon 219 -515 219 -515 0 3
rlabel polysilicon 222 -515 222 -515 0 4
rlabel polysilicon 226 -515 226 -515 0 3
rlabel polysilicon 233 -509 233 -509 0 1
rlabel polysilicon 233 -515 233 -515 0 3
rlabel polysilicon 240 -509 240 -509 0 1
rlabel polysilicon 240 -515 240 -515 0 3
rlabel polysilicon 247 -509 247 -509 0 1
rlabel polysilicon 247 -515 247 -515 0 3
rlabel polysilicon 254 -509 254 -509 0 1
rlabel polysilicon 254 -515 254 -515 0 3
rlabel polysilicon 264 -509 264 -509 0 2
rlabel polysilicon 261 -515 261 -515 0 3
rlabel polysilicon 264 -515 264 -515 0 4
rlabel polysilicon 268 -509 268 -509 0 1
rlabel polysilicon 268 -515 268 -515 0 3
rlabel polysilicon 275 -509 275 -509 0 1
rlabel polysilicon 275 -515 275 -515 0 3
rlabel polysilicon 282 -509 282 -509 0 1
rlabel polysilicon 282 -515 282 -515 0 3
rlabel polysilicon 289 -509 289 -509 0 1
rlabel polysilicon 289 -515 289 -515 0 3
rlabel polysilicon 296 -509 296 -509 0 1
rlabel polysilicon 296 -515 296 -515 0 3
rlabel polysilicon 303 -509 303 -509 0 1
rlabel polysilicon 306 -515 306 -515 0 4
rlabel polysilicon 310 -509 310 -509 0 1
rlabel polysilicon 310 -515 310 -515 0 3
rlabel polysilicon 313 -515 313 -515 0 4
rlabel polysilicon 317 -509 317 -509 0 1
rlabel polysilicon 317 -515 317 -515 0 3
rlabel polysilicon 324 -509 324 -509 0 1
rlabel polysilicon 324 -515 324 -515 0 3
rlabel polysilicon 331 -509 331 -509 0 1
rlabel polysilicon 331 -515 331 -515 0 3
rlabel polysilicon 338 -509 338 -509 0 1
rlabel polysilicon 338 -515 338 -515 0 3
rlabel polysilicon 345 -509 345 -509 0 1
rlabel polysilicon 345 -515 345 -515 0 3
rlabel polysilicon 355 -509 355 -509 0 2
rlabel polysilicon 359 -509 359 -509 0 1
rlabel polysilicon 359 -515 359 -515 0 3
rlabel polysilicon 366 -509 366 -509 0 1
rlabel polysilicon 366 -515 366 -515 0 3
rlabel polysilicon 369 -515 369 -515 0 4
rlabel polysilicon 373 -509 373 -509 0 1
rlabel polysilicon 373 -515 373 -515 0 3
rlabel polysilicon 380 -509 380 -509 0 1
rlabel polysilicon 383 -509 383 -509 0 2
rlabel polysilicon 383 -515 383 -515 0 4
rlabel polysilicon 387 -515 387 -515 0 3
rlabel polysilicon 390 -515 390 -515 0 4
rlabel polysilicon 394 -509 394 -509 0 1
rlabel polysilicon 394 -515 394 -515 0 3
rlabel polysilicon 401 -509 401 -509 0 1
rlabel polysilicon 404 -509 404 -509 0 2
rlabel polysilicon 401 -515 401 -515 0 3
rlabel polysilicon 411 -515 411 -515 0 4
rlabel polysilicon 415 -509 415 -509 0 1
rlabel polysilicon 415 -515 415 -515 0 3
rlabel polysilicon 422 -509 422 -509 0 1
rlabel polysilicon 422 -515 422 -515 0 3
rlabel polysilicon 429 -515 429 -515 0 3
rlabel polysilicon 432 -515 432 -515 0 4
rlabel polysilicon 436 -509 436 -509 0 1
rlabel polysilicon 436 -515 436 -515 0 3
rlabel polysilicon 443 -509 443 -509 0 1
rlabel polysilicon 443 -515 443 -515 0 3
rlabel polysilicon 450 -509 450 -509 0 1
rlabel polysilicon 450 -515 450 -515 0 3
rlabel polysilicon 457 -509 457 -509 0 1
rlabel polysilicon 457 -515 457 -515 0 3
rlabel polysilicon 464 -509 464 -509 0 1
rlabel polysilicon 464 -515 464 -515 0 3
rlabel polysilicon 474 -509 474 -509 0 2
rlabel polysilicon 474 -515 474 -515 0 4
rlabel polysilicon 478 -509 478 -509 0 1
rlabel polysilicon 478 -515 478 -515 0 3
rlabel polysilicon 485 -509 485 -509 0 1
rlabel polysilicon 485 -515 485 -515 0 3
rlabel polysilicon 492 -509 492 -509 0 1
rlabel polysilicon 492 -515 492 -515 0 3
rlabel polysilicon 495 -515 495 -515 0 4
rlabel polysilicon 499 -509 499 -509 0 1
rlabel polysilicon 499 -515 499 -515 0 3
rlabel polysilicon 506 -509 506 -509 0 1
rlabel polysilicon 506 -515 506 -515 0 3
rlabel polysilicon 513 -509 513 -509 0 1
rlabel polysilicon 513 -515 513 -515 0 3
rlabel polysilicon 520 -509 520 -509 0 1
rlabel polysilicon 520 -515 520 -515 0 3
rlabel polysilicon 527 -509 527 -509 0 1
rlabel polysilicon 527 -515 527 -515 0 3
rlabel polysilicon 534 -509 534 -509 0 1
rlabel polysilicon 534 -515 534 -515 0 3
rlabel polysilicon 541 -509 541 -509 0 1
rlabel polysilicon 541 -515 541 -515 0 3
rlabel polysilicon 548 -509 548 -509 0 1
rlabel polysilicon 548 -515 548 -515 0 3
rlabel polysilicon 558 -509 558 -509 0 2
rlabel polysilicon 558 -515 558 -515 0 4
rlabel polysilicon 562 -509 562 -509 0 1
rlabel polysilicon 562 -515 562 -515 0 3
rlabel polysilicon 569 -509 569 -509 0 1
rlabel polysilicon 569 -515 569 -515 0 3
rlabel polysilicon 576 -509 576 -509 0 1
rlabel polysilicon 576 -515 576 -515 0 3
rlabel polysilicon 583 -515 583 -515 0 3
rlabel polysilicon 590 -509 590 -509 0 1
rlabel polysilicon 590 -515 590 -515 0 3
rlabel polysilicon 597 -509 597 -509 0 1
rlabel polysilicon 597 -515 597 -515 0 3
rlabel polysilicon 604 -509 604 -509 0 1
rlabel polysilicon 604 -515 604 -515 0 3
rlabel polysilicon 611 -509 611 -509 0 1
rlabel polysilicon 611 -515 611 -515 0 3
rlabel polysilicon 618 -509 618 -509 0 1
rlabel polysilicon 618 -515 618 -515 0 3
rlabel polysilicon 625 -509 625 -509 0 1
rlabel polysilicon 625 -515 625 -515 0 3
rlabel polysilicon 632 -509 632 -509 0 1
rlabel polysilicon 632 -515 632 -515 0 3
rlabel polysilicon 639 -509 639 -509 0 1
rlabel polysilicon 639 -515 639 -515 0 3
rlabel polysilicon 646 -509 646 -509 0 1
rlabel polysilicon 646 -515 646 -515 0 3
rlabel polysilicon 653 -509 653 -509 0 1
rlabel polysilicon 653 -515 653 -515 0 3
rlabel polysilicon 660 -509 660 -509 0 1
rlabel polysilicon 660 -515 660 -515 0 3
rlabel polysilicon 667 -509 667 -509 0 1
rlabel polysilicon 667 -515 667 -515 0 3
rlabel polysilicon 674 -509 674 -509 0 1
rlabel polysilicon 674 -515 674 -515 0 3
rlabel polysilicon 681 -509 681 -509 0 1
rlabel polysilicon 681 -515 681 -515 0 3
rlabel polysilicon 688 -509 688 -509 0 1
rlabel polysilicon 688 -515 688 -515 0 3
rlabel polysilicon 695 -509 695 -509 0 1
rlabel polysilicon 695 -515 695 -515 0 3
rlabel polysilicon 702 -509 702 -509 0 1
rlabel polysilicon 705 -509 705 -509 0 2
rlabel polysilicon 702 -515 702 -515 0 3
rlabel polysilicon 709 -509 709 -509 0 1
rlabel polysilicon 709 -515 709 -515 0 3
rlabel polysilicon 716 -509 716 -509 0 1
rlabel polysilicon 716 -515 716 -515 0 3
rlabel polysilicon 723 -509 723 -509 0 1
rlabel polysilicon 723 -515 723 -515 0 3
rlabel polysilicon 730 -509 730 -509 0 1
rlabel polysilicon 730 -515 730 -515 0 3
rlabel polysilicon 737 -509 737 -509 0 1
rlabel polysilicon 737 -515 737 -515 0 3
rlabel polysilicon 744 -509 744 -509 0 1
rlabel polysilicon 744 -515 744 -515 0 3
rlabel polysilicon 751 -509 751 -509 0 1
rlabel polysilicon 751 -515 751 -515 0 3
rlabel polysilicon 758 -509 758 -509 0 1
rlabel polysilicon 758 -515 758 -515 0 3
rlabel polysilicon 765 -509 765 -509 0 1
rlabel polysilicon 765 -515 765 -515 0 3
rlabel polysilicon 772 -509 772 -509 0 1
rlabel polysilicon 772 -515 772 -515 0 3
rlabel polysilicon 779 -509 779 -509 0 1
rlabel polysilicon 779 -515 779 -515 0 3
rlabel polysilicon 786 -509 786 -509 0 1
rlabel polysilicon 786 -515 786 -515 0 3
rlabel polysilicon 793 -509 793 -509 0 1
rlabel polysilicon 793 -515 793 -515 0 3
rlabel polysilicon 800 -509 800 -509 0 1
rlabel polysilicon 800 -515 800 -515 0 3
rlabel polysilicon 9 -578 9 -578 0 1
rlabel polysilicon 9 -584 9 -584 0 3
rlabel polysilicon 16 -578 16 -578 0 1
rlabel polysilicon 16 -584 16 -584 0 3
rlabel polysilicon 23 -578 23 -578 0 1
rlabel polysilicon 23 -584 23 -584 0 3
rlabel polysilicon 26 -584 26 -584 0 4
rlabel polysilicon 30 -578 30 -578 0 1
rlabel polysilicon 30 -584 30 -584 0 3
rlabel polysilicon 37 -578 37 -578 0 1
rlabel polysilicon 37 -584 37 -584 0 3
rlabel polysilicon 44 -578 44 -578 0 1
rlabel polysilicon 44 -584 44 -584 0 3
rlabel polysilicon 54 -578 54 -578 0 2
rlabel polysilicon 58 -578 58 -578 0 1
rlabel polysilicon 58 -584 58 -584 0 3
rlabel polysilicon 65 -578 65 -578 0 1
rlabel polysilicon 65 -584 65 -584 0 3
rlabel polysilicon 72 -578 72 -578 0 1
rlabel polysilicon 72 -584 72 -584 0 3
rlabel polysilicon 79 -578 79 -578 0 1
rlabel polysilicon 79 -584 79 -584 0 3
rlabel polysilicon 86 -578 86 -578 0 1
rlabel polysilicon 86 -584 86 -584 0 3
rlabel polysilicon 93 -578 93 -578 0 1
rlabel polysilicon 93 -584 93 -584 0 3
rlabel polysilicon 100 -578 100 -578 0 1
rlabel polysilicon 100 -584 100 -584 0 3
rlabel polysilicon 110 -578 110 -578 0 2
rlabel polysilicon 107 -584 107 -584 0 3
rlabel polysilicon 110 -584 110 -584 0 4
rlabel polysilicon 114 -578 114 -578 0 1
rlabel polysilicon 114 -584 114 -584 0 3
rlabel polysilicon 121 -584 121 -584 0 3
rlabel polysilicon 124 -584 124 -584 0 4
rlabel polysilicon 128 -578 128 -578 0 1
rlabel polysilicon 131 -578 131 -578 0 2
rlabel polysilicon 135 -578 135 -578 0 1
rlabel polysilicon 135 -584 135 -584 0 3
rlabel polysilicon 138 -584 138 -584 0 4
rlabel polysilicon 142 -578 142 -578 0 1
rlabel polysilicon 142 -584 142 -584 0 3
rlabel polysilicon 149 -578 149 -578 0 1
rlabel polysilicon 149 -584 149 -584 0 3
rlabel polysilicon 156 -578 156 -578 0 1
rlabel polysilicon 156 -584 156 -584 0 3
rlabel polysilicon 163 -578 163 -578 0 1
rlabel polysilicon 163 -584 163 -584 0 3
rlabel polysilicon 170 -578 170 -578 0 1
rlabel polysilicon 170 -584 170 -584 0 3
rlabel polysilicon 177 -578 177 -578 0 1
rlabel polysilicon 177 -584 177 -584 0 3
rlabel polysilicon 184 -578 184 -578 0 1
rlabel polysilicon 184 -584 184 -584 0 3
rlabel polysilicon 191 -578 191 -578 0 1
rlabel polysilicon 191 -584 191 -584 0 3
rlabel polysilicon 198 -578 198 -578 0 1
rlabel polysilicon 198 -584 198 -584 0 3
rlabel polysilicon 205 -578 205 -578 0 1
rlabel polysilicon 205 -584 205 -584 0 3
rlabel polysilicon 212 -578 212 -578 0 1
rlabel polysilicon 212 -584 212 -584 0 3
rlabel polysilicon 219 -578 219 -578 0 1
rlabel polysilicon 219 -584 219 -584 0 3
rlabel polysilicon 226 -578 226 -578 0 1
rlabel polysilicon 226 -584 226 -584 0 3
rlabel polysilicon 233 -578 233 -578 0 1
rlabel polysilicon 233 -584 233 -584 0 3
rlabel polysilicon 240 -578 240 -578 0 1
rlabel polysilicon 240 -584 240 -584 0 3
rlabel polysilicon 247 -578 247 -578 0 1
rlabel polysilicon 247 -584 247 -584 0 3
rlabel polysilicon 254 -578 254 -578 0 1
rlabel polysilicon 257 -578 257 -578 0 2
rlabel polysilicon 254 -584 254 -584 0 3
rlabel polysilicon 257 -584 257 -584 0 4
rlabel polysilicon 261 -578 261 -578 0 1
rlabel polysilicon 261 -584 261 -584 0 3
rlabel polysilicon 268 -578 268 -578 0 1
rlabel polysilicon 268 -584 268 -584 0 3
rlabel polysilicon 275 -578 275 -578 0 1
rlabel polysilicon 275 -584 275 -584 0 3
rlabel polysilicon 282 -578 282 -578 0 1
rlabel polysilicon 282 -584 282 -584 0 3
rlabel polysilicon 289 -578 289 -578 0 1
rlabel polysilicon 289 -584 289 -584 0 3
rlabel polysilicon 296 -584 296 -584 0 3
rlabel polysilicon 303 -578 303 -578 0 1
rlabel polysilicon 303 -584 303 -584 0 3
rlabel polysilicon 313 -578 313 -578 0 2
rlabel polysilicon 310 -584 310 -584 0 3
rlabel polysilicon 313 -584 313 -584 0 4
rlabel polysilicon 317 -578 317 -578 0 1
rlabel polysilicon 317 -584 317 -584 0 3
rlabel polysilicon 320 -584 320 -584 0 4
rlabel polysilicon 324 -578 324 -578 0 1
rlabel polysilicon 324 -584 324 -584 0 3
rlabel polysilicon 331 -578 331 -578 0 1
rlabel polysilicon 334 -578 334 -578 0 2
rlabel polysilicon 331 -584 331 -584 0 3
rlabel polysilicon 334 -584 334 -584 0 4
rlabel polysilicon 338 -578 338 -578 0 1
rlabel polysilicon 338 -584 338 -584 0 3
rlabel polysilicon 345 -578 345 -578 0 1
rlabel polysilicon 345 -584 345 -584 0 3
rlabel polysilicon 352 -578 352 -578 0 1
rlabel polysilicon 352 -584 352 -584 0 3
rlabel polysilicon 359 -578 359 -578 0 1
rlabel polysilicon 359 -584 359 -584 0 3
rlabel polysilicon 366 -578 366 -578 0 1
rlabel polysilicon 366 -584 366 -584 0 3
rlabel polysilicon 373 -578 373 -578 0 1
rlabel polysilicon 373 -584 373 -584 0 3
rlabel polysilicon 380 -578 380 -578 0 1
rlabel polysilicon 383 -578 383 -578 0 2
rlabel polysilicon 380 -584 380 -584 0 3
rlabel polysilicon 383 -584 383 -584 0 4
rlabel polysilicon 387 -578 387 -578 0 1
rlabel polysilicon 387 -584 387 -584 0 3
rlabel polysilicon 394 -578 394 -578 0 1
rlabel polysilicon 394 -584 394 -584 0 3
rlabel polysilicon 401 -578 401 -578 0 1
rlabel polysilicon 401 -584 401 -584 0 3
rlabel polysilicon 408 -578 408 -578 0 1
rlabel polysilicon 408 -584 408 -584 0 3
rlabel polysilicon 415 -578 415 -578 0 1
rlabel polysilicon 418 -578 418 -578 0 2
rlabel polysilicon 415 -584 415 -584 0 3
rlabel polysilicon 422 -578 422 -578 0 1
rlabel polysilicon 422 -584 422 -584 0 3
rlabel polysilicon 429 -578 429 -578 0 1
rlabel polysilicon 429 -584 429 -584 0 3
rlabel polysilicon 436 -578 436 -578 0 1
rlabel polysilicon 436 -584 436 -584 0 3
rlabel polysilicon 443 -578 443 -578 0 1
rlabel polysilicon 443 -584 443 -584 0 3
rlabel polysilicon 450 -578 450 -578 0 1
rlabel polysilicon 450 -584 450 -584 0 3
rlabel polysilicon 457 -578 457 -578 0 1
rlabel polysilicon 460 -584 460 -584 0 4
rlabel polysilicon 464 -578 464 -578 0 1
rlabel polysilicon 467 -578 467 -578 0 2
rlabel polysilicon 464 -584 464 -584 0 3
rlabel polysilicon 467 -584 467 -584 0 4
rlabel polysilicon 471 -578 471 -578 0 1
rlabel polysilicon 471 -584 471 -584 0 3
rlabel polysilicon 478 -578 478 -578 0 1
rlabel polysilicon 478 -584 478 -584 0 3
rlabel polysilicon 485 -578 485 -578 0 1
rlabel polysilicon 488 -578 488 -578 0 2
rlabel polysilicon 485 -584 485 -584 0 3
rlabel polysilicon 492 -578 492 -578 0 1
rlabel polysilicon 492 -584 492 -584 0 3
rlabel polysilicon 499 -578 499 -578 0 1
rlabel polysilicon 499 -584 499 -584 0 3
rlabel polysilicon 506 -578 506 -578 0 1
rlabel polysilicon 506 -584 506 -584 0 3
rlabel polysilicon 509 -584 509 -584 0 4
rlabel polysilicon 513 -584 513 -584 0 3
rlabel polysilicon 516 -584 516 -584 0 4
rlabel polysilicon 520 -578 520 -578 0 1
rlabel polysilicon 520 -584 520 -584 0 3
rlabel polysilicon 527 -578 527 -578 0 1
rlabel polysilicon 527 -584 527 -584 0 3
rlabel polysilicon 534 -578 534 -578 0 1
rlabel polysilicon 534 -584 534 -584 0 3
rlabel polysilicon 541 -578 541 -578 0 1
rlabel polysilicon 541 -584 541 -584 0 3
rlabel polysilicon 551 -578 551 -578 0 2
rlabel polysilicon 548 -584 548 -584 0 3
rlabel polysilicon 555 -578 555 -578 0 1
rlabel polysilicon 555 -584 555 -584 0 3
rlabel polysilicon 562 -578 562 -578 0 1
rlabel polysilicon 562 -584 562 -584 0 3
rlabel polysilicon 569 -578 569 -578 0 1
rlabel polysilicon 569 -584 569 -584 0 3
rlabel polysilicon 576 -578 576 -578 0 1
rlabel polysilicon 576 -584 576 -584 0 3
rlabel polysilicon 583 -578 583 -578 0 1
rlabel polysilicon 583 -584 583 -584 0 3
rlabel polysilicon 590 -578 590 -578 0 1
rlabel polysilicon 590 -584 590 -584 0 3
rlabel polysilicon 597 -578 597 -578 0 1
rlabel polysilicon 597 -584 597 -584 0 3
rlabel polysilicon 604 -578 604 -578 0 1
rlabel polysilicon 604 -584 604 -584 0 3
rlabel polysilicon 611 -578 611 -578 0 1
rlabel polysilicon 611 -584 611 -584 0 3
rlabel polysilicon 618 -578 618 -578 0 1
rlabel polysilicon 618 -584 618 -584 0 3
rlabel polysilicon 625 -578 625 -578 0 1
rlabel polysilicon 625 -584 625 -584 0 3
rlabel polysilicon 632 -578 632 -578 0 1
rlabel polysilicon 632 -584 632 -584 0 3
rlabel polysilicon 639 -578 639 -578 0 1
rlabel polysilicon 639 -584 639 -584 0 3
rlabel polysilicon 646 -578 646 -578 0 1
rlabel polysilicon 646 -584 646 -584 0 3
rlabel polysilicon 653 -578 653 -578 0 1
rlabel polysilicon 653 -584 653 -584 0 3
rlabel polysilicon 660 -578 660 -578 0 1
rlabel polysilicon 660 -584 660 -584 0 3
rlabel polysilicon 667 -578 667 -578 0 1
rlabel polysilicon 667 -584 667 -584 0 3
rlabel polysilicon 674 -578 674 -578 0 1
rlabel polysilicon 674 -584 674 -584 0 3
rlabel polysilicon 681 -578 681 -578 0 1
rlabel polysilicon 681 -584 681 -584 0 3
rlabel polysilicon 688 -578 688 -578 0 1
rlabel polysilicon 688 -584 688 -584 0 3
rlabel polysilicon 695 -578 695 -578 0 1
rlabel polysilicon 695 -584 695 -584 0 3
rlabel polysilicon 702 -578 702 -578 0 1
rlabel polysilicon 702 -584 702 -584 0 3
rlabel polysilicon 709 -578 709 -578 0 1
rlabel polysilicon 709 -584 709 -584 0 3
rlabel polysilicon 716 -578 716 -578 0 1
rlabel polysilicon 716 -584 716 -584 0 3
rlabel polysilicon 723 -578 723 -578 0 1
rlabel polysilicon 723 -584 723 -584 0 3
rlabel polysilicon 730 -578 730 -578 0 1
rlabel polysilicon 730 -584 730 -584 0 3
rlabel polysilicon 737 -578 737 -578 0 1
rlabel polysilicon 737 -584 737 -584 0 3
rlabel polysilicon 744 -578 744 -578 0 1
rlabel polysilicon 744 -584 744 -584 0 3
rlabel polysilicon 751 -578 751 -578 0 1
rlabel polysilicon 751 -584 751 -584 0 3
rlabel polysilicon 758 -578 758 -578 0 1
rlabel polysilicon 758 -584 758 -584 0 3
rlabel polysilicon 765 -578 765 -578 0 1
rlabel polysilicon 765 -584 765 -584 0 3
rlabel polysilicon 772 -578 772 -578 0 1
rlabel polysilicon 772 -584 772 -584 0 3
rlabel polysilicon 779 -578 779 -578 0 1
rlabel polysilicon 779 -584 779 -584 0 3
rlabel polysilicon 786 -578 786 -578 0 1
rlabel polysilicon 786 -584 786 -584 0 3
rlabel polysilicon 793 -578 793 -578 0 1
rlabel polysilicon 793 -584 793 -584 0 3
rlabel polysilicon 800 -578 800 -578 0 1
rlabel polysilicon 800 -584 800 -584 0 3
rlabel polysilicon 807 -578 807 -578 0 1
rlabel polysilicon 807 -584 807 -584 0 3
rlabel polysilicon 814 -578 814 -578 0 1
rlabel polysilicon 814 -584 814 -584 0 3
rlabel polysilicon 821 -578 821 -578 0 1
rlabel polysilicon 821 -584 821 -584 0 3
rlabel polysilicon 2 -667 2 -667 0 1
rlabel polysilicon 2 -673 2 -673 0 3
rlabel polysilicon 9 -667 9 -667 0 1
rlabel polysilicon 9 -673 9 -673 0 3
rlabel polysilicon 16 -667 16 -667 0 1
rlabel polysilicon 16 -673 16 -673 0 3
rlabel polysilicon 23 -667 23 -667 0 1
rlabel polysilicon 23 -673 23 -673 0 3
rlabel polysilicon 30 -667 30 -667 0 1
rlabel polysilicon 30 -673 30 -673 0 3
rlabel polysilicon 37 -667 37 -667 0 1
rlabel polysilicon 37 -673 37 -673 0 3
rlabel polysilicon 44 -667 44 -667 0 1
rlabel polysilicon 44 -673 44 -673 0 3
rlabel polysilicon 51 -667 51 -667 0 1
rlabel polysilicon 54 -667 54 -667 0 2
rlabel polysilicon 51 -673 51 -673 0 3
rlabel polysilicon 58 -667 58 -667 0 1
rlabel polysilicon 61 -667 61 -667 0 2
rlabel polysilicon 61 -673 61 -673 0 4
rlabel polysilicon 68 -667 68 -667 0 2
rlabel polysilicon 65 -673 65 -673 0 3
rlabel polysilicon 68 -673 68 -673 0 4
rlabel polysilicon 72 -667 72 -667 0 1
rlabel polysilicon 72 -673 72 -673 0 3
rlabel polysilicon 79 -667 79 -667 0 1
rlabel polysilicon 79 -673 79 -673 0 3
rlabel polysilicon 86 -667 86 -667 0 1
rlabel polysilicon 86 -673 86 -673 0 3
rlabel polysilicon 93 -667 93 -667 0 1
rlabel polysilicon 93 -673 93 -673 0 3
rlabel polysilicon 100 -667 100 -667 0 1
rlabel polysilicon 100 -673 100 -673 0 3
rlabel polysilicon 107 -667 107 -667 0 1
rlabel polysilicon 110 -667 110 -667 0 2
rlabel polysilicon 107 -673 107 -673 0 3
rlabel polysilicon 114 -667 114 -667 0 1
rlabel polysilicon 114 -673 114 -673 0 3
rlabel polysilicon 121 -667 121 -667 0 1
rlabel polysilicon 121 -673 121 -673 0 3
rlabel polysilicon 128 -667 128 -667 0 1
rlabel polysilicon 128 -673 128 -673 0 3
rlabel polysilicon 135 -667 135 -667 0 1
rlabel polysilicon 135 -673 135 -673 0 3
rlabel polysilicon 142 -667 142 -667 0 1
rlabel polysilicon 142 -673 142 -673 0 3
rlabel polysilicon 149 -667 149 -667 0 1
rlabel polysilicon 149 -673 149 -673 0 3
rlabel polysilicon 156 -667 156 -667 0 1
rlabel polysilicon 156 -673 156 -673 0 3
rlabel polysilicon 163 -667 163 -667 0 1
rlabel polysilicon 163 -673 163 -673 0 3
rlabel polysilicon 170 -667 170 -667 0 1
rlabel polysilicon 170 -673 170 -673 0 3
rlabel polysilicon 177 -667 177 -667 0 1
rlabel polysilicon 177 -673 177 -673 0 3
rlabel polysilicon 184 -667 184 -667 0 1
rlabel polysilicon 184 -673 184 -673 0 3
rlabel polysilicon 191 -667 191 -667 0 1
rlabel polysilicon 191 -673 191 -673 0 3
rlabel polysilicon 198 -667 198 -667 0 1
rlabel polysilicon 198 -673 198 -673 0 3
rlabel polysilicon 205 -667 205 -667 0 1
rlabel polysilicon 205 -673 205 -673 0 3
rlabel polysilicon 212 -667 212 -667 0 1
rlabel polysilicon 215 -667 215 -667 0 2
rlabel polysilicon 212 -673 212 -673 0 3
rlabel polysilicon 219 -667 219 -667 0 1
rlabel polysilicon 219 -673 219 -673 0 3
rlabel polysilicon 226 -667 226 -667 0 1
rlabel polysilicon 229 -667 229 -667 0 2
rlabel polysilicon 229 -673 229 -673 0 4
rlabel polysilicon 233 -667 233 -667 0 1
rlabel polysilicon 233 -673 233 -673 0 3
rlabel polysilicon 240 -667 240 -667 0 1
rlabel polysilicon 240 -673 240 -673 0 3
rlabel polysilicon 247 -667 247 -667 0 1
rlabel polysilicon 247 -673 247 -673 0 3
rlabel polysilicon 254 -667 254 -667 0 1
rlabel polysilicon 254 -673 254 -673 0 3
rlabel polysilicon 261 -667 261 -667 0 1
rlabel polysilicon 261 -673 261 -673 0 3
rlabel polysilicon 268 -667 268 -667 0 1
rlabel polysilicon 271 -667 271 -667 0 2
rlabel polysilicon 268 -673 268 -673 0 3
rlabel polysilicon 271 -673 271 -673 0 4
rlabel polysilicon 275 -667 275 -667 0 1
rlabel polysilicon 275 -673 275 -673 0 3
rlabel polysilicon 282 -667 282 -667 0 1
rlabel polysilicon 282 -673 282 -673 0 3
rlabel polysilicon 289 -667 289 -667 0 1
rlabel polysilicon 292 -667 292 -667 0 2
rlabel polysilicon 296 -667 296 -667 0 1
rlabel polysilicon 299 -667 299 -667 0 2
rlabel polysilicon 296 -673 296 -673 0 3
rlabel polysilicon 303 -667 303 -667 0 1
rlabel polysilicon 303 -673 303 -673 0 3
rlabel polysilicon 310 -667 310 -667 0 1
rlabel polysilicon 310 -673 310 -673 0 3
rlabel polysilicon 317 -667 317 -667 0 1
rlabel polysilicon 317 -673 317 -673 0 3
rlabel polysilicon 324 -667 324 -667 0 1
rlabel polysilicon 324 -673 324 -673 0 3
rlabel polysilicon 331 -667 331 -667 0 1
rlabel polysilicon 331 -673 331 -673 0 3
rlabel polysilicon 338 -667 338 -667 0 1
rlabel polysilicon 338 -673 338 -673 0 3
rlabel polysilicon 345 -667 345 -667 0 1
rlabel polysilicon 348 -667 348 -667 0 2
rlabel polysilicon 348 -673 348 -673 0 4
rlabel polysilicon 352 -667 352 -667 0 1
rlabel polysilicon 352 -673 352 -673 0 3
rlabel polysilicon 359 -667 359 -667 0 1
rlabel polysilicon 359 -673 359 -673 0 3
rlabel polysilicon 366 -667 366 -667 0 1
rlabel polysilicon 369 -667 369 -667 0 2
rlabel polysilicon 369 -673 369 -673 0 4
rlabel polysilicon 373 -667 373 -667 0 1
rlabel polysilicon 373 -673 373 -673 0 3
rlabel polysilicon 383 -667 383 -667 0 2
rlabel polysilicon 380 -673 380 -673 0 3
rlabel polysilicon 387 -667 387 -667 0 1
rlabel polysilicon 387 -673 387 -673 0 3
rlabel polysilicon 394 -667 394 -667 0 1
rlabel polysilicon 394 -673 394 -673 0 3
rlabel polysilicon 401 -667 401 -667 0 1
rlabel polysilicon 401 -673 401 -673 0 3
rlabel polysilicon 408 -667 408 -667 0 1
rlabel polysilicon 408 -673 408 -673 0 3
rlabel polysilicon 415 -667 415 -667 0 1
rlabel polysilicon 415 -673 415 -673 0 3
rlabel polysilicon 418 -673 418 -673 0 4
rlabel polysilicon 422 -667 422 -667 0 1
rlabel polysilicon 422 -673 422 -673 0 3
rlabel polysilicon 429 -667 429 -667 0 1
rlabel polysilicon 429 -673 429 -673 0 3
rlabel polysilicon 436 -667 436 -667 0 1
rlabel polysilicon 436 -673 436 -673 0 3
rlabel polysilicon 443 -667 443 -667 0 1
rlabel polysilicon 443 -673 443 -673 0 3
rlabel polysilicon 450 -667 450 -667 0 1
rlabel polysilicon 453 -667 453 -667 0 2
rlabel polysilicon 453 -673 453 -673 0 4
rlabel polysilicon 457 -667 457 -667 0 1
rlabel polysilicon 460 -667 460 -667 0 2
rlabel polysilicon 460 -673 460 -673 0 4
rlabel polysilicon 464 -667 464 -667 0 1
rlabel polysilicon 464 -673 464 -673 0 3
rlabel polysilicon 471 -667 471 -667 0 1
rlabel polysilicon 471 -673 471 -673 0 3
rlabel polysilicon 478 -667 478 -667 0 1
rlabel polysilicon 478 -673 478 -673 0 3
rlabel polysilicon 485 -667 485 -667 0 1
rlabel polysilicon 485 -673 485 -673 0 3
rlabel polysilicon 492 -667 492 -667 0 1
rlabel polysilicon 492 -673 492 -673 0 3
rlabel polysilicon 499 -667 499 -667 0 1
rlabel polysilicon 499 -673 499 -673 0 3
rlabel polysilicon 506 -667 506 -667 0 1
rlabel polysilicon 506 -673 506 -673 0 3
rlabel polysilicon 513 -667 513 -667 0 1
rlabel polysilicon 513 -673 513 -673 0 3
rlabel polysilicon 520 -667 520 -667 0 1
rlabel polysilicon 520 -673 520 -673 0 3
rlabel polysilicon 527 -667 527 -667 0 1
rlabel polysilicon 527 -673 527 -673 0 3
rlabel polysilicon 534 -667 534 -667 0 1
rlabel polysilicon 534 -673 534 -673 0 3
rlabel polysilicon 544 -673 544 -673 0 4
rlabel polysilicon 548 -667 548 -667 0 1
rlabel polysilicon 548 -673 548 -673 0 3
rlabel polysilicon 555 -667 555 -667 0 1
rlabel polysilicon 555 -673 555 -673 0 3
rlabel polysilicon 562 -667 562 -667 0 1
rlabel polysilicon 562 -673 562 -673 0 3
rlabel polysilicon 569 -667 569 -667 0 1
rlabel polysilicon 569 -673 569 -673 0 3
rlabel polysilicon 576 -667 576 -667 0 1
rlabel polysilicon 576 -673 576 -673 0 3
rlabel polysilicon 583 -667 583 -667 0 1
rlabel polysilicon 583 -673 583 -673 0 3
rlabel polysilicon 590 -667 590 -667 0 1
rlabel polysilicon 590 -673 590 -673 0 3
rlabel polysilicon 597 -667 597 -667 0 1
rlabel polysilicon 597 -673 597 -673 0 3
rlabel polysilicon 604 -667 604 -667 0 1
rlabel polysilicon 604 -673 604 -673 0 3
rlabel polysilicon 611 -667 611 -667 0 1
rlabel polysilicon 611 -673 611 -673 0 3
rlabel polysilicon 618 -667 618 -667 0 1
rlabel polysilicon 618 -673 618 -673 0 3
rlabel polysilicon 625 -667 625 -667 0 1
rlabel polysilicon 625 -673 625 -673 0 3
rlabel polysilicon 632 -667 632 -667 0 1
rlabel polysilicon 632 -673 632 -673 0 3
rlabel polysilicon 639 -667 639 -667 0 1
rlabel polysilicon 639 -673 639 -673 0 3
rlabel polysilicon 646 -667 646 -667 0 1
rlabel polysilicon 646 -673 646 -673 0 3
rlabel polysilicon 653 -667 653 -667 0 1
rlabel polysilicon 653 -673 653 -673 0 3
rlabel polysilicon 660 -667 660 -667 0 1
rlabel polysilicon 660 -673 660 -673 0 3
rlabel polysilicon 667 -667 667 -667 0 1
rlabel polysilicon 667 -673 667 -673 0 3
rlabel polysilicon 674 -667 674 -667 0 1
rlabel polysilicon 674 -673 674 -673 0 3
rlabel polysilicon 681 -667 681 -667 0 1
rlabel polysilicon 681 -673 681 -673 0 3
rlabel polysilicon 688 -667 688 -667 0 1
rlabel polysilicon 688 -673 688 -673 0 3
rlabel polysilicon 695 -667 695 -667 0 1
rlabel polysilicon 695 -673 695 -673 0 3
rlabel polysilicon 702 -667 702 -667 0 1
rlabel polysilicon 702 -673 702 -673 0 3
rlabel polysilicon 709 -667 709 -667 0 1
rlabel polysilicon 709 -673 709 -673 0 3
rlabel polysilicon 716 -667 716 -667 0 1
rlabel polysilicon 716 -673 716 -673 0 3
rlabel polysilicon 723 -667 723 -667 0 1
rlabel polysilicon 723 -673 723 -673 0 3
rlabel polysilicon 730 -667 730 -667 0 1
rlabel polysilicon 730 -673 730 -673 0 3
rlabel polysilicon 737 -667 737 -667 0 1
rlabel polysilicon 737 -673 737 -673 0 3
rlabel polysilicon 744 -667 744 -667 0 1
rlabel polysilicon 744 -673 744 -673 0 3
rlabel polysilicon 751 -667 751 -667 0 1
rlabel polysilicon 751 -673 751 -673 0 3
rlabel polysilicon 758 -667 758 -667 0 1
rlabel polysilicon 758 -673 758 -673 0 3
rlabel polysilicon 765 -667 765 -667 0 1
rlabel polysilicon 765 -673 765 -673 0 3
rlabel polysilicon 772 -667 772 -667 0 1
rlabel polysilicon 772 -673 772 -673 0 3
rlabel polysilicon 779 -667 779 -667 0 1
rlabel polysilicon 779 -673 779 -673 0 3
rlabel polysilicon 786 -667 786 -667 0 1
rlabel polysilicon 793 -667 793 -667 0 1
rlabel polysilicon 12 -734 12 -734 0 2
rlabel polysilicon 16 -734 16 -734 0 1
rlabel polysilicon 19 -740 19 -740 0 4
rlabel polysilicon 23 -734 23 -734 0 1
rlabel polysilicon 23 -740 23 -740 0 3
rlabel polysilicon 30 -734 30 -734 0 1
rlabel polysilicon 30 -740 30 -740 0 3
rlabel polysilicon 37 -734 37 -734 0 1
rlabel polysilicon 37 -740 37 -740 0 3
rlabel polysilicon 44 -734 44 -734 0 1
rlabel polysilicon 44 -740 44 -740 0 3
rlabel polysilicon 51 -734 51 -734 0 1
rlabel polysilicon 51 -740 51 -740 0 3
rlabel polysilicon 58 -734 58 -734 0 1
rlabel polysilicon 58 -740 58 -740 0 3
rlabel polysilicon 65 -734 65 -734 0 1
rlabel polysilicon 68 -734 68 -734 0 2
rlabel polysilicon 68 -740 68 -740 0 4
rlabel polysilicon 72 -734 72 -734 0 1
rlabel polysilicon 72 -740 72 -740 0 3
rlabel polysilicon 79 -734 79 -734 0 1
rlabel polysilicon 79 -740 79 -740 0 3
rlabel polysilicon 89 -734 89 -734 0 2
rlabel polysilicon 86 -740 86 -740 0 3
rlabel polysilicon 89 -740 89 -740 0 4
rlabel polysilicon 93 -734 93 -734 0 1
rlabel polysilicon 93 -740 93 -740 0 3
rlabel polysilicon 100 -734 100 -734 0 1
rlabel polysilicon 100 -740 100 -740 0 3
rlabel polysilicon 107 -734 107 -734 0 1
rlabel polysilicon 107 -740 107 -740 0 3
rlabel polysilicon 114 -734 114 -734 0 1
rlabel polysilicon 114 -740 114 -740 0 3
rlabel polysilicon 121 -734 121 -734 0 1
rlabel polysilicon 121 -740 121 -740 0 3
rlabel polysilicon 128 -734 128 -734 0 1
rlabel polysilicon 131 -734 131 -734 0 2
rlabel polysilicon 135 -734 135 -734 0 1
rlabel polysilicon 135 -740 135 -740 0 3
rlabel polysilicon 142 -734 142 -734 0 1
rlabel polysilicon 142 -740 142 -740 0 3
rlabel polysilicon 149 -734 149 -734 0 1
rlabel polysilicon 149 -740 149 -740 0 3
rlabel polysilicon 156 -734 156 -734 0 1
rlabel polysilicon 156 -740 156 -740 0 3
rlabel polysilicon 163 -734 163 -734 0 1
rlabel polysilicon 166 -734 166 -734 0 2
rlabel polysilicon 166 -740 166 -740 0 4
rlabel polysilicon 170 -734 170 -734 0 1
rlabel polysilicon 170 -740 170 -740 0 3
rlabel polysilicon 177 -734 177 -734 0 1
rlabel polysilicon 177 -740 177 -740 0 3
rlabel polysilicon 184 -734 184 -734 0 1
rlabel polysilicon 184 -740 184 -740 0 3
rlabel polysilicon 191 -734 191 -734 0 1
rlabel polysilicon 191 -740 191 -740 0 3
rlabel polysilicon 198 -734 198 -734 0 1
rlabel polysilicon 198 -740 198 -740 0 3
rlabel polysilicon 205 -734 205 -734 0 1
rlabel polysilicon 205 -740 205 -740 0 3
rlabel polysilicon 212 -734 212 -734 0 1
rlabel polysilicon 212 -740 212 -740 0 3
rlabel polysilicon 219 -734 219 -734 0 1
rlabel polysilicon 219 -740 219 -740 0 3
rlabel polysilicon 226 -734 226 -734 0 1
rlabel polysilicon 229 -734 229 -734 0 2
rlabel polysilicon 229 -740 229 -740 0 4
rlabel polysilicon 233 -734 233 -734 0 1
rlabel polysilicon 233 -740 233 -740 0 3
rlabel polysilicon 240 -734 240 -734 0 1
rlabel polysilicon 247 -734 247 -734 0 1
rlabel polysilicon 247 -740 247 -740 0 3
rlabel polysilicon 254 -734 254 -734 0 1
rlabel polysilicon 254 -740 254 -740 0 3
rlabel polysilicon 261 -734 261 -734 0 1
rlabel polysilicon 261 -740 261 -740 0 3
rlabel polysilicon 268 -734 268 -734 0 1
rlabel polysilicon 271 -734 271 -734 0 2
rlabel polysilicon 268 -740 268 -740 0 3
rlabel polysilicon 275 -734 275 -734 0 1
rlabel polysilicon 275 -740 275 -740 0 3
rlabel polysilicon 282 -734 282 -734 0 1
rlabel polysilicon 282 -740 282 -740 0 3
rlabel polysilicon 289 -734 289 -734 0 1
rlabel polysilicon 289 -740 289 -740 0 3
rlabel polysilicon 296 -734 296 -734 0 1
rlabel polysilicon 296 -740 296 -740 0 3
rlabel polysilicon 303 -734 303 -734 0 1
rlabel polysilicon 303 -740 303 -740 0 3
rlabel polysilicon 310 -734 310 -734 0 1
rlabel polysilicon 310 -740 310 -740 0 3
rlabel polysilicon 317 -734 317 -734 0 1
rlabel polysilicon 320 -734 320 -734 0 2
rlabel polysilicon 317 -740 317 -740 0 3
rlabel polysilicon 320 -740 320 -740 0 4
rlabel polysilicon 324 -734 324 -734 0 1
rlabel polysilicon 324 -740 324 -740 0 3
rlabel polysilicon 331 -734 331 -734 0 1
rlabel polysilicon 331 -740 331 -740 0 3
rlabel polysilicon 338 -734 338 -734 0 1
rlabel polysilicon 338 -740 338 -740 0 3
rlabel polysilicon 345 -734 345 -734 0 1
rlabel polysilicon 345 -740 345 -740 0 3
rlabel polysilicon 348 -740 348 -740 0 4
rlabel polysilicon 352 -734 352 -734 0 1
rlabel polysilicon 352 -740 352 -740 0 3
rlabel polysilicon 359 -734 359 -734 0 1
rlabel polysilicon 359 -740 359 -740 0 3
rlabel polysilicon 366 -734 366 -734 0 1
rlabel polysilicon 366 -740 366 -740 0 3
rlabel polysilicon 373 -734 373 -734 0 1
rlabel polysilicon 373 -740 373 -740 0 3
rlabel polysilicon 380 -734 380 -734 0 1
rlabel polysilicon 380 -740 380 -740 0 3
rlabel polysilicon 383 -740 383 -740 0 4
rlabel polysilicon 387 -734 387 -734 0 1
rlabel polysilicon 387 -740 387 -740 0 3
rlabel polysilicon 394 -734 394 -734 0 1
rlabel polysilicon 397 -740 397 -740 0 4
rlabel polysilicon 401 -734 401 -734 0 1
rlabel polysilicon 401 -740 401 -740 0 3
rlabel polysilicon 408 -734 408 -734 0 1
rlabel polysilicon 408 -740 408 -740 0 3
rlabel polysilicon 415 -734 415 -734 0 1
rlabel polysilicon 415 -740 415 -740 0 3
rlabel polysilicon 422 -734 422 -734 0 1
rlabel polysilicon 425 -734 425 -734 0 2
rlabel polysilicon 422 -740 422 -740 0 3
rlabel polysilicon 425 -740 425 -740 0 4
rlabel polysilicon 429 -734 429 -734 0 1
rlabel polysilicon 429 -740 429 -740 0 3
rlabel polysilicon 436 -734 436 -734 0 1
rlabel polysilicon 436 -740 436 -740 0 3
rlabel polysilicon 443 -734 443 -734 0 1
rlabel polysilicon 446 -734 446 -734 0 2
rlabel polysilicon 443 -740 443 -740 0 3
rlabel polysilicon 446 -740 446 -740 0 4
rlabel polysilicon 450 -734 450 -734 0 1
rlabel polysilicon 450 -740 450 -740 0 3
rlabel polysilicon 453 -740 453 -740 0 4
rlabel polysilicon 457 -734 457 -734 0 1
rlabel polysilicon 457 -740 457 -740 0 3
rlabel polysilicon 464 -734 464 -734 0 1
rlabel polysilicon 464 -740 464 -740 0 3
rlabel polysilicon 471 -734 471 -734 0 1
rlabel polysilicon 471 -740 471 -740 0 3
rlabel polysilicon 478 -734 478 -734 0 1
rlabel polysilicon 478 -740 478 -740 0 3
rlabel polysilicon 485 -734 485 -734 0 1
rlabel polysilicon 485 -740 485 -740 0 3
rlabel polysilicon 492 -734 492 -734 0 1
rlabel polysilicon 492 -740 492 -740 0 3
rlabel polysilicon 499 -734 499 -734 0 1
rlabel polysilicon 499 -740 499 -740 0 3
rlabel polysilicon 506 -734 506 -734 0 1
rlabel polysilicon 506 -740 506 -740 0 3
rlabel polysilicon 513 -734 513 -734 0 1
rlabel polysilicon 513 -740 513 -740 0 3
rlabel polysilicon 523 -734 523 -734 0 2
rlabel polysilicon 527 -734 527 -734 0 1
rlabel polysilicon 530 -734 530 -734 0 2
rlabel polysilicon 527 -740 527 -740 0 3
rlabel polysilicon 530 -740 530 -740 0 4
rlabel polysilicon 534 -734 534 -734 0 1
rlabel polysilicon 534 -740 534 -740 0 3
rlabel polysilicon 541 -734 541 -734 0 1
rlabel polysilicon 541 -740 541 -740 0 3
rlabel polysilicon 551 -734 551 -734 0 2
rlabel polysilicon 548 -740 548 -740 0 3
rlabel polysilicon 555 -734 555 -734 0 1
rlabel polysilicon 555 -740 555 -740 0 3
rlabel polysilicon 562 -734 562 -734 0 1
rlabel polysilicon 562 -740 562 -740 0 3
rlabel polysilicon 569 -740 569 -740 0 3
rlabel polysilicon 572 -740 572 -740 0 4
rlabel polysilicon 576 -734 576 -734 0 1
rlabel polysilicon 576 -740 576 -740 0 3
rlabel polysilicon 583 -734 583 -734 0 1
rlabel polysilicon 583 -740 583 -740 0 3
rlabel polysilicon 590 -734 590 -734 0 1
rlabel polysilicon 590 -740 590 -740 0 3
rlabel polysilicon 597 -734 597 -734 0 1
rlabel polysilicon 597 -740 597 -740 0 3
rlabel polysilicon 604 -734 604 -734 0 1
rlabel polysilicon 604 -740 604 -740 0 3
rlabel polysilicon 611 -734 611 -734 0 1
rlabel polysilicon 611 -740 611 -740 0 3
rlabel polysilicon 618 -734 618 -734 0 1
rlabel polysilicon 618 -740 618 -740 0 3
rlabel polysilicon 625 -734 625 -734 0 1
rlabel polysilicon 625 -740 625 -740 0 3
rlabel polysilicon 632 -734 632 -734 0 1
rlabel polysilicon 632 -740 632 -740 0 3
rlabel polysilicon 639 -734 639 -734 0 1
rlabel polysilicon 639 -740 639 -740 0 3
rlabel polysilicon 646 -734 646 -734 0 1
rlabel polysilicon 646 -740 646 -740 0 3
rlabel polysilicon 653 -734 653 -734 0 1
rlabel polysilicon 653 -740 653 -740 0 3
rlabel polysilicon 660 -734 660 -734 0 1
rlabel polysilicon 660 -740 660 -740 0 3
rlabel polysilicon 667 -734 667 -734 0 1
rlabel polysilicon 667 -740 667 -740 0 3
rlabel polysilicon 674 -734 674 -734 0 1
rlabel polysilicon 674 -740 674 -740 0 3
rlabel polysilicon 681 -734 681 -734 0 1
rlabel polysilicon 681 -740 681 -740 0 3
rlabel polysilicon 688 -734 688 -734 0 1
rlabel polysilicon 688 -740 688 -740 0 3
rlabel polysilicon 695 -734 695 -734 0 1
rlabel polysilicon 695 -740 695 -740 0 3
rlabel polysilicon 702 -734 702 -734 0 1
rlabel polysilicon 702 -740 702 -740 0 3
rlabel polysilicon 709 -734 709 -734 0 1
rlabel polysilicon 709 -740 709 -740 0 3
rlabel polysilicon 716 -734 716 -734 0 1
rlabel polysilicon 716 -740 716 -740 0 3
rlabel polysilicon 723 -734 723 -734 0 1
rlabel polysilicon 723 -740 723 -740 0 3
rlabel polysilicon 730 -734 730 -734 0 1
rlabel polysilicon 730 -740 730 -740 0 3
rlabel polysilicon 737 -734 737 -734 0 1
rlabel polysilicon 737 -740 737 -740 0 3
rlabel polysilicon 744 -734 744 -734 0 1
rlabel polysilicon 744 -740 744 -740 0 3
rlabel polysilicon 751 -734 751 -734 0 1
rlabel polysilicon 751 -740 751 -740 0 3
rlabel polysilicon 758 -734 758 -734 0 1
rlabel polysilicon 758 -740 758 -740 0 3
rlabel polysilicon 765 -734 765 -734 0 1
rlabel polysilicon 765 -740 765 -740 0 3
rlabel polysilicon 772 -734 772 -734 0 1
rlabel polysilicon 772 -740 772 -740 0 3
rlabel polysilicon 779 -734 779 -734 0 1
rlabel polysilicon 782 -734 782 -734 0 2
rlabel polysilicon 782 -740 782 -740 0 4
rlabel polysilicon 786 -734 786 -734 0 1
rlabel polysilicon 786 -740 786 -740 0 3
rlabel polysilicon 793 -734 793 -734 0 1
rlabel polysilicon 793 -740 793 -740 0 3
rlabel polysilicon 800 -734 800 -734 0 1
rlabel polysilicon 800 -740 800 -740 0 3
rlabel polysilicon 807 -734 807 -734 0 1
rlabel polysilicon 807 -740 807 -740 0 3
rlabel polysilicon 2 -805 2 -805 0 1
rlabel polysilicon 9 -805 9 -805 0 1
rlabel polysilicon 9 -811 9 -811 0 3
rlabel polysilicon 16 -805 16 -805 0 1
rlabel polysilicon 16 -811 16 -811 0 3
rlabel polysilicon 23 -805 23 -805 0 1
rlabel polysilicon 23 -811 23 -811 0 3
rlabel polysilicon 30 -805 30 -805 0 1
rlabel polysilicon 30 -811 30 -811 0 3
rlabel polysilicon 37 -805 37 -805 0 1
rlabel polysilicon 40 -805 40 -805 0 2
rlabel polysilicon 40 -811 40 -811 0 4
rlabel polysilicon 44 -805 44 -805 0 1
rlabel polysilicon 44 -811 44 -811 0 3
rlabel polysilicon 51 -805 51 -805 0 1
rlabel polysilicon 51 -811 51 -811 0 3
rlabel polysilicon 58 -805 58 -805 0 1
rlabel polysilicon 58 -811 58 -811 0 3
rlabel polysilicon 65 -805 65 -805 0 1
rlabel polysilicon 65 -811 65 -811 0 3
rlabel polysilicon 72 -805 72 -805 0 1
rlabel polysilicon 75 -805 75 -805 0 2
rlabel polysilicon 72 -811 72 -811 0 3
rlabel polysilicon 75 -811 75 -811 0 4
rlabel polysilicon 79 -805 79 -805 0 1
rlabel polysilicon 79 -811 79 -811 0 3
rlabel polysilicon 86 -805 86 -805 0 1
rlabel polysilicon 86 -811 86 -811 0 3
rlabel polysilicon 93 -805 93 -805 0 1
rlabel polysilicon 93 -811 93 -811 0 3
rlabel polysilicon 100 -805 100 -805 0 1
rlabel polysilicon 100 -811 100 -811 0 3
rlabel polysilicon 107 -805 107 -805 0 1
rlabel polysilicon 107 -811 107 -811 0 3
rlabel polysilicon 114 -805 114 -805 0 1
rlabel polysilicon 114 -811 114 -811 0 3
rlabel polysilicon 121 -805 121 -805 0 1
rlabel polysilicon 121 -811 121 -811 0 3
rlabel polysilicon 128 -805 128 -805 0 1
rlabel polysilicon 128 -811 128 -811 0 3
rlabel polysilicon 131 -811 131 -811 0 4
rlabel polysilicon 135 -805 135 -805 0 1
rlabel polysilicon 135 -811 135 -811 0 3
rlabel polysilicon 142 -805 142 -805 0 1
rlabel polysilicon 142 -811 142 -811 0 3
rlabel polysilicon 149 -805 149 -805 0 1
rlabel polysilicon 149 -811 149 -811 0 3
rlabel polysilicon 159 -805 159 -805 0 2
rlabel polysilicon 156 -811 156 -811 0 3
rlabel polysilicon 159 -811 159 -811 0 4
rlabel polysilicon 163 -805 163 -805 0 1
rlabel polysilicon 163 -811 163 -811 0 3
rlabel polysilicon 170 -805 170 -805 0 1
rlabel polysilicon 170 -811 170 -811 0 3
rlabel polysilicon 177 -805 177 -805 0 1
rlabel polysilicon 177 -811 177 -811 0 3
rlabel polysilicon 184 -805 184 -805 0 1
rlabel polysilicon 184 -811 184 -811 0 3
rlabel polysilicon 191 -805 191 -805 0 1
rlabel polysilicon 191 -811 191 -811 0 3
rlabel polysilicon 198 -805 198 -805 0 1
rlabel polysilicon 198 -811 198 -811 0 3
rlabel polysilicon 205 -805 205 -805 0 1
rlabel polysilicon 205 -811 205 -811 0 3
rlabel polysilicon 212 -805 212 -805 0 1
rlabel polysilicon 215 -805 215 -805 0 2
rlabel polysilicon 219 -805 219 -805 0 1
rlabel polysilicon 219 -811 219 -811 0 3
rlabel polysilicon 226 -805 226 -805 0 1
rlabel polysilicon 226 -811 226 -811 0 3
rlabel polysilicon 233 -805 233 -805 0 1
rlabel polysilicon 233 -811 233 -811 0 3
rlabel polysilicon 240 -811 240 -811 0 3
rlabel polysilicon 247 -805 247 -805 0 1
rlabel polysilicon 247 -811 247 -811 0 3
rlabel polysilicon 250 -811 250 -811 0 4
rlabel polysilicon 254 -805 254 -805 0 1
rlabel polysilicon 257 -811 257 -811 0 4
rlabel polysilicon 261 -805 261 -805 0 1
rlabel polysilicon 261 -811 261 -811 0 3
rlabel polysilicon 268 -805 268 -805 0 1
rlabel polysilicon 268 -811 268 -811 0 3
rlabel polysilicon 275 -805 275 -805 0 1
rlabel polysilicon 275 -811 275 -811 0 3
rlabel polysilicon 282 -805 282 -805 0 1
rlabel polysilicon 285 -805 285 -805 0 2
rlabel polysilicon 282 -811 282 -811 0 3
rlabel polysilicon 289 -805 289 -805 0 1
rlabel polysilicon 289 -811 289 -811 0 3
rlabel polysilicon 296 -805 296 -805 0 1
rlabel polysilicon 296 -811 296 -811 0 3
rlabel polysilicon 303 -805 303 -805 0 1
rlabel polysilicon 303 -811 303 -811 0 3
rlabel polysilicon 310 -805 310 -805 0 1
rlabel polysilicon 317 -805 317 -805 0 1
rlabel polysilicon 317 -811 317 -811 0 3
rlabel polysilicon 324 -805 324 -805 0 1
rlabel polysilicon 324 -811 324 -811 0 3
rlabel polysilicon 331 -805 331 -805 0 1
rlabel polysilicon 331 -811 331 -811 0 3
rlabel polysilicon 338 -805 338 -805 0 1
rlabel polysilicon 338 -811 338 -811 0 3
rlabel polysilicon 345 -805 345 -805 0 1
rlabel polysilicon 345 -811 345 -811 0 3
rlabel polysilicon 352 -805 352 -805 0 1
rlabel polysilicon 352 -811 352 -811 0 3
rlabel polysilicon 359 -805 359 -805 0 1
rlabel polysilicon 362 -805 362 -805 0 2
rlabel polysilicon 366 -805 366 -805 0 1
rlabel polysilicon 366 -811 366 -811 0 3
rlabel polysilicon 373 -805 373 -805 0 1
rlabel polysilicon 376 -805 376 -805 0 2
rlabel polysilicon 373 -811 373 -811 0 3
rlabel polysilicon 376 -811 376 -811 0 4
rlabel polysilicon 380 -805 380 -805 0 1
rlabel polysilicon 380 -811 380 -811 0 3
rlabel polysilicon 387 -805 387 -805 0 1
rlabel polysilicon 387 -811 387 -811 0 3
rlabel polysilicon 397 -811 397 -811 0 4
rlabel polysilicon 401 -805 401 -805 0 1
rlabel polysilicon 404 -805 404 -805 0 2
rlabel polysilicon 404 -811 404 -811 0 4
rlabel polysilicon 411 -805 411 -805 0 2
rlabel polysilicon 411 -811 411 -811 0 4
rlabel polysilicon 415 -805 415 -805 0 1
rlabel polysilicon 415 -811 415 -811 0 3
rlabel polysilicon 422 -805 422 -805 0 1
rlabel polysilicon 422 -811 422 -811 0 3
rlabel polysilicon 429 -805 429 -805 0 1
rlabel polysilicon 429 -811 429 -811 0 3
rlabel polysilicon 436 -805 436 -805 0 1
rlabel polysilicon 436 -811 436 -811 0 3
rlabel polysilicon 443 -805 443 -805 0 1
rlabel polysilicon 443 -811 443 -811 0 3
rlabel polysilicon 450 -805 450 -805 0 1
rlabel polysilicon 453 -805 453 -805 0 2
rlabel polysilicon 450 -811 450 -811 0 3
rlabel polysilicon 457 -805 457 -805 0 1
rlabel polysilicon 457 -811 457 -811 0 3
rlabel polysilicon 464 -805 464 -805 0 1
rlabel polysilicon 464 -811 464 -811 0 3
rlabel polysilicon 471 -805 471 -805 0 1
rlabel polysilicon 471 -811 471 -811 0 3
rlabel polysilicon 478 -805 478 -805 0 1
rlabel polysilicon 481 -805 481 -805 0 2
rlabel polysilicon 481 -811 481 -811 0 4
rlabel polysilicon 485 -805 485 -805 0 1
rlabel polysilicon 485 -811 485 -811 0 3
rlabel polysilicon 492 -805 492 -805 0 1
rlabel polysilicon 492 -811 492 -811 0 3
rlabel polysilicon 499 -805 499 -805 0 1
rlabel polysilicon 499 -811 499 -811 0 3
rlabel polysilicon 506 -805 506 -805 0 1
rlabel polysilicon 506 -811 506 -811 0 3
rlabel polysilicon 513 -805 513 -805 0 1
rlabel polysilicon 513 -811 513 -811 0 3
rlabel polysilicon 520 -805 520 -805 0 1
rlabel polysilicon 520 -811 520 -811 0 3
rlabel polysilicon 527 -805 527 -805 0 1
rlabel polysilicon 527 -811 527 -811 0 3
rlabel polysilicon 534 -805 534 -805 0 1
rlabel polysilicon 534 -811 534 -811 0 3
rlabel polysilicon 541 -805 541 -805 0 1
rlabel polysilicon 541 -811 541 -811 0 3
rlabel polysilicon 548 -805 548 -805 0 1
rlabel polysilicon 551 -805 551 -805 0 2
rlabel polysilicon 548 -811 548 -811 0 3
rlabel polysilicon 555 -805 555 -805 0 1
rlabel polysilicon 555 -811 555 -811 0 3
rlabel polysilicon 562 -805 562 -805 0 1
rlabel polysilicon 562 -811 562 -811 0 3
rlabel polysilicon 569 -805 569 -805 0 1
rlabel polysilicon 569 -811 569 -811 0 3
rlabel polysilicon 576 -805 576 -805 0 1
rlabel polysilicon 576 -811 576 -811 0 3
rlabel polysilicon 583 -805 583 -805 0 1
rlabel polysilicon 583 -811 583 -811 0 3
rlabel polysilicon 590 -805 590 -805 0 1
rlabel polysilicon 590 -811 590 -811 0 3
rlabel polysilicon 597 -805 597 -805 0 1
rlabel polysilicon 600 -805 600 -805 0 2
rlabel polysilicon 597 -811 597 -811 0 3
rlabel polysilicon 604 -805 604 -805 0 1
rlabel polysilicon 604 -811 604 -811 0 3
rlabel polysilicon 611 -805 611 -805 0 1
rlabel polysilicon 611 -811 611 -811 0 3
rlabel polysilicon 618 -805 618 -805 0 1
rlabel polysilicon 618 -811 618 -811 0 3
rlabel polysilicon 625 -805 625 -805 0 1
rlabel polysilicon 625 -811 625 -811 0 3
rlabel polysilicon 632 -805 632 -805 0 1
rlabel polysilicon 632 -811 632 -811 0 3
rlabel polysilicon 639 -805 639 -805 0 1
rlabel polysilicon 639 -811 639 -811 0 3
rlabel polysilicon 646 -805 646 -805 0 1
rlabel polysilicon 646 -811 646 -811 0 3
rlabel polysilicon 653 -805 653 -805 0 1
rlabel polysilicon 653 -811 653 -811 0 3
rlabel polysilicon 660 -805 660 -805 0 1
rlabel polysilicon 660 -811 660 -811 0 3
rlabel polysilicon 667 -805 667 -805 0 1
rlabel polysilicon 667 -811 667 -811 0 3
rlabel polysilicon 674 -805 674 -805 0 1
rlabel polysilicon 674 -811 674 -811 0 3
rlabel polysilicon 681 -805 681 -805 0 1
rlabel polysilicon 681 -811 681 -811 0 3
rlabel polysilicon 688 -805 688 -805 0 1
rlabel polysilicon 688 -811 688 -811 0 3
rlabel polysilicon 695 -805 695 -805 0 1
rlabel polysilicon 695 -811 695 -811 0 3
rlabel polysilicon 702 -805 702 -805 0 1
rlabel polysilicon 702 -811 702 -811 0 3
rlabel polysilicon 709 -805 709 -805 0 1
rlabel polysilicon 709 -811 709 -811 0 3
rlabel polysilicon 716 -805 716 -805 0 1
rlabel polysilicon 716 -811 716 -811 0 3
rlabel polysilicon 723 -805 723 -805 0 1
rlabel polysilicon 723 -811 723 -811 0 3
rlabel polysilicon 730 -805 730 -805 0 1
rlabel polysilicon 730 -811 730 -811 0 3
rlabel polysilicon 737 -805 737 -805 0 1
rlabel polysilicon 737 -811 737 -811 0 3
rlabel polysilicon 744 -805 744 -805 0 1
rlabel polysilicon 744 -811 744 -811 0 3
rlabel polysilicon 751 -805 751 -805 0 1
rlabel polysilicon 751 -811 751 -811 0 3
rlabel polysilicon 758 -805 758 -805 0 1
rlabel polysilicon 758 -811 758 -811 0 3
rlabel polysilicon 765 -805 765 -805 0 1
rlabel polysilicon 765 -811 765 -811 0 3
rlabel polysilicon 772 -805 772 -805 0 1
rlabel polysilicon 779 -805 779 -805 0 1
rlabel polysilicon 779 -811 779 -811 0 3
rlabel polysilicon 786 -805 786 -805 0 1
rlabel polysilicon 786 -811 786 -811 0 3
rlabel polysilicon 9 -860 9 -860 0 1
rlabel polysilicon 9 -866 9 -866 0 3
rlabel polysilicon 19 -866 19 -866 0 4
rlabel polysilicon 23 -860 23 -860 0 1
rlabel polysilicon 23 -866 23 -866 0 3
rlabel polysilicon 30 -860 30 -860 0 1
rlabel polysilicon 30 -866 30 -866 0 3
rlabel polysilicon 40 -866 40 -866 0 4
rlabel polysilicon 44 -860 44 -860 0 1
rlabel polysilicon 44 -866 44 -866 0 3
rlabel polysilicon 51 -860 51 -860 0 1
rlabel polysilicon 54 -866 54 -866 0 4
rlabel polysilicon 58 -860 58 -860 0 1
rlabel polysilicon 58 -866 58 -866 0 3
rlabel polysilicon 65 -860 65 -860 0 1
rlabel polysilicon 65 -866 65 -866 0 3
rlabel polysilicon 72 -860 72 -860 0 1
rlabel polysilicon 72 -866 72 -866 0 3
rlabel polysilicon 79 -860 79 -860 0 1
rlabel polysilicon 79 -866 79 -866 0 3
rlabel polysilicon 86 -860 86 -860 0 1
rlabel polysilicon 86 -866 86 -866 0 3
rlabel polysilicon 93 -860 93 -860 0 1
rlabel polysilicon 93 -866 93 -866 0 3
rlabel polysilicon 100 -860 100 -860 0 1
rlabel polysilicon 100 -866 100 -866 0 3
rlabel polysilicon 107 -860 107 -860 0 1
rlabel polysilicon 110 -860 110 -860 0 2
rlabel polysilicon 107 -866 107 -866 0 3
rlabel polysilicon 110 -866 110 -866 0 4
rlabel polysilicon 114 -860 114 -860 0 1
rlabel polysilicon 117 -860 117 -860 0 2
rlabel polysilicon 117 -866 117 -866 0 4
rlabel polysilicon 121 -860 121 -860 0 1
rlabel polysilicon 121 -866 121 -866 0 3
rlabel polysilicon 128 -860 128 -860 0 1
rlabel polysilicon 128 -866 128 -866 0 3
rlabel polysilicon 138 -860 138 -860 0 2
rlabel polysilicon 135 -866 135 -866 0 3
rlabel polysilicon 138 -866 138 -866 0 4
rlabel polysilicon 142 -860 142 -860 0 1
rlabel polysilicon 142 -866 142 -866 0 3
rlabel polysilicon 149 -860 149 -860 0 1
rlabel polysilicon 149 -866 149 -866 0 3
rlabel polysilicon 156 -860 156 -860 0 1
rlabel polysilicon 156 -866 156 -866 0 3
rlabel polysilicon 163 -860 163 -860 0 1
rlabel polysilicon 163 -866 163 -866 0 3
rlabel polysilicon 173 -860 173 -860 0 2
rlabel polysilicon 170 -866 170 -866 0 3
rlabel polysilicon 173 -866 173 -866 0 4
rlabel polysilicon 177 -860 177 -860 0 1
rlabel polysilicon 177 -866 177 -866 0 3
rlabel polysilicon 184 -860 184 -860 0 1
rlabel polysilicon 184 -866 184 -866 0 3
rlabel polysilicon 191 -860 191 -860 0 1
rlabel polysilicon 191 -866 191 -866 0 3
rlabel polysilicon 198 -860 198 -860 0 1
rlabel polysilicon 198 -866 198 -866 0 3
rlabel polysilicon 205 -860 205 -860 0 1
rlabel polysilicon 205 -866 205 -866 0 3
rlabel polysilicon 212 -860 212 -860 0 1
rlabel polysilicon 212 -866 212 -866 0 3
rlabel polysilicon 219 -860 219 -860 0 1
rlabel polysilicon 219 -866 219 -866 0 3
rlabel polysilicon 226 -860 226 -860 0 1
rlabel polysilicon 226 -866 226 -866 0 3
rlabel polysilicon 233 -860 233 -860 0 1
rlabel polysilicon 233 -866 233 -866 0 3
rlabel polysilicon 240 -860 240 -860 0 1
rlabel polysilicon 240 -866 240 -866 0 3
rlabel polysilicon 247 -860 247 -860 0 1
rlabel polysilicon 247 -866 247 -866 0 3
rlabel polysilicon 254 -860 254 -860 0 1
rlabel polysilicon 254 -866 254 -866 0 3
rlabel polysilicon 261 -860 261 -860 0 1
rlabel polysilicon 264 -860 264 -860 0 2
rlabel polysilicon 268 -860 268 -860 0 1
rlabel polysilicon 271 -860 271 -860 0 2
rlabel polysilicon 271 -866 271 -866 0 4
rlabel polysilicon 275 -860 275 -860 0 1
rlabel polysilicon 275 -866 275 -866 0 3
rlabel polysilicon 282 -860 282 -860 0 1
rlabel polysilicon 282 -866 282 -866 0 3
rlabel polysilicon 289 -860 289 -860 0 1
rlabel polysilicon 289 -866 289 -866 0 3
rlabel polysilicon 296 -860 296 -860 0 1
rlabel polysilicon 296 -866 296 -866 0 3
rlabel polysilicon 303 -860 303 -860 0 1
rlabel polysilicon 303 -866 303 -866 0 3
rlabel polysilicon 310 -860 310 -860 0 1
rlabel polysilicon 310 -866 310 -866 0 3
rlabel polysilicon 317 -860 317 -860 0 1
rlabel polysilicon 317 -866 317 -866 0 3
rlabel polysilicon 324 -860 324 -860 0 1
rlabel polysilicon 324 -866 324 -866 0 3
rlabel polysilicon 331 -860 331 -860 0 1
rlabel polysilicon 331 -866 331 -866 0 3
rlabel polysilicon 338 -860 338 -860 0 1
rlabel polysilicon 338 -866 338 -866 0 3
rlabel polysilicon 345 -860 345 -860 0 1
rlabel polysilicon 348 -860 348 -860 0 2
rlabel polysilicon 348 -866 348 -866 0 4
rlabel polysilicon 352 -860 352 -860 0 1
rlabel polysilicon 352 -866 352 -866 0 3
rlabel polysilicon 359 -860 359 -860 0 1
rlabel polysilicon 359 -866 359 -866 0 3
rlabel polysilicon 366 -860 366 -860 0 1
rlabel polysilicon 366 -866 366 -866 0 3
rlabel polysilicon 369 -866 369 -866 0 4
rlabel polysilicon 373 -860 373 -860 0 1
rlabel polysilicon 373 -866 373 -866 0 3
rlabel polysilicon 380 -860 380 -860 0 1
rlabel polysilicon 383 -866 383 -866 0 4
rlabel polysilicon 387 -860 387 -860 0 1
rlabel polysilicon 390 -860 390 -860 0 2
rlabel polysilicon 390 -866 390 -866 0 4
rlabel polysilicon 394 -860 394 -860 0 1
rlabel polysilicon 394 -866 394 -866 0 3
rlabel polysilicon 401 -860 401 -860 0 1
rlabel polysilicon 401 -866 401 -866 0 3
rlabel polysilicon 408 -860 408 -860 0 1
rlabel polysilicon 408 -866 408 -866 0 3
rlabel polysilicon 415 -860 415 -860 0 1
rlabel polysilicon 415 -866 415 -866 0 3
rlabel polysilicon 422 -860 422 -860 0 1
rlabel polysilicon 422 -866 422 -866 0 3
rlabel polysilicon 429 -860 429 -860 0 1
rlabel polysilicon 429 -866 429 -866 0 3
rlabel polysilicon 436 -860 436 -860 0 1
rlabel polysilicon 436 -866 436 -866 0 3
rlabel polysilicon 443 -860 443 -860 0 1
rlabel polysilicon 443 -866 443 -866 0 3
rlabel polysilicon 450 -860 450 -860 0 1
rlabel polysilicon 450 -866 450 -866 0 3
rlabel polysilicon 457 -860 457 -860 0 1
rlabel polysilicon 457 -866 457 -866 0 3
rlabel polysilicon 464 -860 464 -860 0 1
rlabel polysilicon 464 -866 464 -866 0 3
rlabel polysilicon 471 -860 471 -860 0 1
rlabel polysilicon 471 -866 471 -866 0 3
rlabel polysilicon 478 -860 478 -860 0 1
rlabel polysilicon 478 -866 478 -866 0 3
rlabel polysilicon 485 -860 485 -860 0 1
rlabel polysilicon 485 -866 485 -866 0 3
rlabel polysilicon 492 -860 492 -860 0 1
rlabel polysilicon 492 -866 492 -866 0 3
rlabel polysilicon 502 -860 502 -860 0 2
rlabel polysilicon 502 -866 502 -866 0 4
rlabel polysilicon 506 -860 506 -860 0 1
rlabel polysilicon 506 -866 506 -866 0 3
rlabel polysilicon 513 -860 513 -860 0 1
rlabel polysilicon 513 -866 513 -866 0 3
rlabel polysilicon 520 -860 520 -860 0 1
rlabel polysilicon 520 -866 520 -866 0 3
rlabel polysilicon 527 -860 527 -860 0 1
rlabel polysilicon 527 -866 527 -866 0 3
rlabel polysilicon 534 -860 534 -860 0 1
rlabel polysilicon 534 -866 534 -866 0 3
rlabel polysilicon 544 -860 544 -860 0 2
rlabel polysilicon 541 -866 541 -866 0 3
rlabel polysilicon 544 -866 544 -866 0 4
rlabel polysilicon 548 -860 548 -860 0 1
rlabel polysilicon 548 -866 548 -866 0 3
rlabel polysilicon 555 -860 555 -860 0 1
rlabel polysilicon 555 -866 555 -866 0 3
rlabel polysilicon 562 -860 562 -860 0 1
rlabel polysilicon 562 -866 562 -866 0 3
rlabel polysilicon 569 -860 569 -860 0 1
rlabel polysilicon 569 -866 569 -866 0 3
rlabel polysilicon 576 -860 576 -860 0 1
rlabel polysilicon 576 -866 576 -866 0 3
rlabel polysilicon 583 -860 583 -860 0 1
rlabel polysilicon 583 -866 583 -866 0 3
rlabel polysilicon 590 -860 590 -860 0 1
rlabel polysilicon 590 -866 590 -866 0 3
rlabel polysilicon 597 -860 597 -860 0 1
rlabel polysilicon 597 -866 597 -866 0 3
rlabel polysilicon 607 -860 607 -860 0 2
rlabel polysilicon 604 -866 604 -866 0 3
rlabel polysilicon 611 -860 611 -860 0 1
rlabel polysilicon 611 -866 611 -866 0 3
rlabel polysilicon 618 -860 618 -860 0 1
rlabel polysilicon 618 -866 618 -866 0 3
rlabel polysilicon 625 -860 625 -860 0 1
rlabel polysilicon 625 -866 625 -866 0 3
rlabel polysilicon 632 -860 632 -860 0 1
rlabel polysilicon 632 -866 632 -866 0 3
rlabel polysilicon 639 -860 639 -860 0 1
rlabel polysilicon 639 -866 639 -866 0 3
rlabel polysilicon 646 -860 646 -860 0 1
rlabel polysilicon 646 -866 646 -866 0 3
rlabel polysilicon 653 -860 653 -860 0 1
rlabel polysilicon 653 -866 653 -866 0 3
rlabel polysilicon 660 -860 660 -860 0 1
rlabel polysilicon 660 -866 660 -866 0 3
rlabel polysilicon 667 -860 667 -860 0 1
rlabel polysilicon 667 -866 667 -866 0 3
rlabel polysilicon 681 -866 681 -866 0 3
rlabel polysilicon 684 -866 684 -866 0 4
rlabel polysilicon 688 -860 688 -860 0 1
rlabel polysilicon 688 -866 688 -866 0 3
rlabel polysilicon 695 -860 695 -860 0 1
rlabel polysilicon 695 -866 695 -866 0 3
rlabel polysilicon 702 -860 702 -860 0 1
rlabel polysilicon 702 -866 702 -866 0 3
rlabel polysilicon 726 -860 726 -860 0 2
rlabel polysilicon 726 -866 726 -866 0 4
rlabel polysilicon 730 -866 730 -866 0 3
rlabel polysilicon 733 -866 733 -866 0 4
rlabel polysilicon 737 -860 737 -860 0 1
rlabel polysilicon 737 -866 737 -866 0 3
rlabel polysilicon 744 -860 744 -860 0 1
rlabel polysilicon 744 -866 744 -866 0 3
rlabel polysilicon 751 -860 751 -860 0 1
rlabel polysilicon 751 -866 751 -866 0 3
rlabel polysilicon 758 -860 758 -860 0 1
rlabel polysilicon 758 -866 758 -866 0 3
rlabel polysilicon 44 -913 44 -913 0 1
rlabel polysilicon 44 -919 44 -919 0 3
rlabel polysilicon 51 -913 51 -913 0 1
rlabel polysilicon 51 -919 51 -919 0 3
rlabel polysilicon 58 -913 58 -913 0 1
rlabel polysilicon 58 -919 58 -919 0 3
rlabel polysilicon 65 -913 65 -913 0 1
rlabel polysilicon 65 -919 65 -919 0 3
rlabel polysilicon 72 -913 72 -913 0 1
rlabel polysilicon 79 -913 79 -913 0 1
rlabel polysilicon 79 -919 79 -919 0 3
rlabel polysilicon 86 -913 86 -913 0 1
rlabel polysilicon 86 -919 86 -919 0 3
rlabel polysilicon 93 -913 93 -913 0 1
rlabel polysilicon 93 -919 93 -919 0 3
rlabel polysilicon 100 -913 100 -913 0 1
rlabel polysilicon 100 -919 100 -919 0 3
rlabel polysilicon 107 -913 107 -913 0 1
rlabel polysilicon 107 -919 107 -919 0 3
rlabel polysilicon 114 -913 114 -913 0 1
rlabel polysilicon 114 -919 114 -919 0 3
rlabel polysilicon 124 -913 124 -913 0 2
rlabel polysilicon 121 -919 121 -919 0 3
rlabel polysilicon 128 -913 128 -913 0 1
rlabel polysilicon 128 -919 128 -919 0 3
rlabel polysilicon 135 -913 135 -913 0 1
rlabel polysilicon 135 -919 135 -919 0 3
rlabel polysilicon 142 -913 142 -913 0 1
rlabel polysilicon 142 -919 142 -919 0 3
rlabel polysilicon 149 -913 149 -913 0 1
rlabel polysilicon 149 -919 149 -919 0 3
rlabel polysilicon 156 -913 156 -913 0 1
rlabel polysilicon 156 -919 156 -919 0 3
rlabel polysilicon 159 -919 159 -919 0 4
rlabel polysilicon 163 -913 163 -913 0 1
rlabel polysilicon 163 -919 163 -919 0 3
rlabel polysilicon 170 -913 170 -913 0 1
rlabel polysilicon 170 -919 170 -919 0 3
rlabel polysilicon 177 -913 177 -913 0 1
rlabel polysilicon 180 -913 180 -913 0 2
rlabel polysilicon 184 -913 184 -913 0 1
rlabel polysilicon 184 -919 184 -919 0 3
rlabel polysilicon 191 -913 191 -913 0 1
rlabel polysilicon 191 -919 191 -919 0 3
rlabel polysilicon 198 -913 198 -913 0 1
rlabel polysilicon 198 -919 198 -919 0 3
rlabel polysilicon 205 -913 205 -913 0 1
rlabel polysilicon 208 -913 208 -913 0 2
rlabel polysilicon 205 -919 205 -919 0 3
rlabel polysilicon 212 -913 212 -913 0 1
rlabel polysilicon 212 -919 212 -919 0 3
rlabel polysilicon 219 -913 219 -913 0 1
rlabel polysilicon 219 -919 219 -919 0 3
rlabel polysilicon 226 -913 226 -913 0 1
rlabel polysilicon 226 -919 226 -919 0 3
rlabel polysilicon 233 -913 233 -913 0 1
rlabel polysilicon 233 -919 233 -919 0 3
rlabel polysilicon 240 -913 240 -913 0 1
rlabel polysilicon 240 -919 240 -919 0 3
rlabel polysilicon 247 -913 247 -913 0 1
rlabel polysilicon 247 -919 247 -919 0 3
rlabel polysilicon 257 -913 257 -913 0 2
rlabel polysilicon 254 -919 254 -919 0 3
rlabel polysilicon 257 -919 257 -919 0 4
rlabel polysilicon 261 -913 261 -913 0 1
rlabel polysilicon 261 -919 261 -919 0 3
rlabel polysilicon 271 -913 271 -913 0 2
rlabel polysilicon 268 -919 268 -919 0 3
rlabel polysilicon 275 -913 275 -913 0 1
rlabel polysilicon 275 -919 275 -919 0 3
rlabel polysilicon 282 -913 282 -913 0 1
rlabel polysilicon 282 -919 282 -919 0 3
rlabel polysilicon 289 -913 289 -913 0 1
rlabel polysilicon 289 -919 289 -919 0 3
rlabel polysilicon 296 -913 296 -913 0 1
rlabel polysilicon 299 -913 299 -913 0 2
rlabel polysilicon 299 -919 299 -919 0 4
rlabel polysilicon 303 -913 303 -913 0 1
rlabel polysilicon 303 -919 303 -919 0 3
rlabel polysilicon 310 -913 310 -913 0 1
rlabel polysilicon 310 -919 310 -919 0 3
rlabel polysilicon 317 -913 317 -913 0 1
rlabel polysilicon 317 -919 317 -919 0 3
rlabel polysilicon 324 -919 324 -919 0 3
rlabel polysilicon 331 -913 331 -913 0 1
rlabel polysilicon 331 -919 331 -919 0 3
rlabel polysilicon 338 -913 338 -913 0 1
rlabel polysilicon 338 -919 338 -919 0 3
rlabel polysilicon 345 -913 345 -913 0 1
rlabel polysilicon 345 -919 345 -919 0 3
rlabel polysilicon 352 -913 352 -913 0 1
rlabel polysilicon 352 -919 352 -919 0 3
rlabel polysilicon 359 -913 359 -913 0 1
rlabel polysilicon 359 -919 359 -919 0 3
rlabel polysilicon 366 -919 366 -919 0 3
rlabel polysilicon 369 -919 369 -919 0 4
rlabel polysilicon 373 -913 373 -913 0 1
rlabel polysilicon 376 -913 376 -913 0 2
rlabel polysilicon 380 -913 380 -913 0 1
rlabel polysilicon 380 -919 380 -919 0 3
rlabel polysilicon 387 -913 387 -913 0 1
rlabel polysilicon 387 -919 387 -919 0 3
rlabel polysilicon 394 -913 394 -913 0 1
rlabel polysilicon 397 -913 397 -913 0 2
rlabel polysilicon 401 -913 401 -913 0 1
rlabel polysilicon 401 -919 401 -919 0 3
rlabel polysilicon 408 -913 408 -913 0 1
rlabel polysilicon 408 -919 408 -919 0 3
rlabel polysilicon 415 -913 415 -913 0 1
rlabel polysilicon 415 -919 415 -919 0 3
rlabel polysilicon 422 -913 422 -913 0 1
rlabel polysilicon 422 -919 422 -919 0 3
rlabel polysilicon 429 -913 429 -913 0 1
rlabel polysilicon 429 -919 429 -919 0 3
rlabel polysilicon 436 -913 436 -913 0 1
rlabel polysilicon 436 -919 436 -919 0 3
rlabel polysilicon 443 -913 443 -913 0 1
rlabel polysilicon 443 -919 443 -919 0 3
rlabel polysilicon 450 -913 450 -913 0 1
rlabel polysilicon 450 -919 450 -919 0 3
rlabel polysilicon 457 -913 457 -913 0 1
rlabel polysilicon 457 -919 457 -919 0 3
rlabel polysilicon 467 -913 467 -913 0 2
rlabel polysilicon 464 -919 464 -919 0 3
rlabel polysilicon 471 -913 471 -913 0 1
rlabel polysilicon 471 -919 471 -919 0 3
rlabel polysilicon 478 -913 478 -913 0 1
rlabel polysilicon 478 -919 478 -919 0 3
rlabel polysilicon 485 -913 485 -913 0 1
rlabel polysilicon 485 -919 485 -919 0 3
rlabel polysilicon 492 -913 492 -913 0 1
rlabel polysilicon 492 -919 492 -919 0 3
rlabel polysilicon 499 -913 499 -913 0 1
rlabel polysilicon 499 -919 499 -919 0 3
rlabel polysilicon 506 -913 506 -913 0 1
rlabel polysilicon 506 -919 506 -919 0 3
rlabel polysilicon 513 -913 513 -913 0 1
rlabel polysilicon 513 -919 513 -919 0 3
rlabel polysilicon 523 -913 523 -913 0 2
rlabel polysilicon 520 -919 520 -919 0 3
rlabel polysilicon 527 -913 527 -913 0 1
rlabel polysilicon 527 -919 527 -919 0 3
rlabel polysilicon 534 -913 534 -913 0 1
rlabel polysilicon 534 -919 534 -919 0 3
rlabel polysilicon 541 -913 541 -913 0 1
rlabel polysilicon 541 -919 541 -919 0 3
rlabel polysilicon 548 -913 548 -913 0 1
rlabel polysilicon 548 -919 548 -919 0 3
rlabel polysilicon 555 -913 555 -913 0 1
rlabel polysilicon 555 -919 555 -919 0 3
rlabel polysilicon 562 -913 562 -913 0 1
rlabel polysilicon 562 -919 562 -919 0 3
rlabel polysilicon 569 -913 569 -913 0 1
rlabel polysilicon 569 -919 569 -919 0 3
rlabel polysilicon 576 -913 576 -913 0 1
rlabel polysilicon 576 -919 576 -919 0 3
rlabel polysilicon 583 -913 583 -913 0 1
rlabel polysilicon 583 -919 583 -919 0 3
rlabel polysilicon 590 -913 590 -913 0 1
rlabel polysilicon 590 -919 590 -919 0 3
rlabel polysilicon 597 -913 597 -913 0 1
rlabel polysilicon 597 -919 597 -919 0 3
rlabel polysilicon 604 -913 604 -913 0 1
rlabel polysilicon 604 -919 604 -919 0 3
rlabel polysilicon 611 -913 611 -913 0 1
rlabel polysilicon 611 -919 611 -919 0 3
rlabel polysilicon 618 -913 618 -913 0 1
rlabel polysilicon 618 -919 618 -919 0 3
rlabel polysilicon 625 -913 625 -913 0 1
rlabel polysilicon 625 -919 625 -919 0 3
rlabel polysilicon 632 -913 632 -913 0 1
rlabel polysilicon 632 -919 632 -919 0 3
rlabel polysilicon 642 -913 642 -913 0 2
rlabel polysilicon 639 -919 639 -919 0 3
rlabel polysilicon 642 -919 642 -919 0 4
rlabel polysilicon 646 -913 646 -913 0 1
rlabel polysilicon 646 -919 646 -919 0 3
rlabel polysilicon 653 -919 653 -919 0 3
rlabel polysilicon 660 -913 660 -913 0 1
rlabel polysilicon 663 -913 663 -913 0 2
rlabel polysilicon 667 -913 667 -913 0 1
rlabel polysilicon 667 -919 667 -919 0 3
rlabel polysilicon 674 -913 674 -913 0 1
rlabel polysilicon 674 -919 674 -919 0 3
rlabel polysilicon 681 -913 681 -913 0 1
rlabel polysilicon 681 -919 681 -919 0 3
rlabel polysilicon 716 -913 716 -913 0 1
rlabel polysilicon 716 -919 716 -919 0 3
rlabel polysilicon 747 -913 747 -913 0 2
rlabel polysilicon 744 -919 744 -919 0 3
rlabel polysilicon 65 -972 65 -972 0 1
rlabel polysilicon 65 -978 65 -978 0 3
rlabel polysilicon 72 -972 72 -972 0 1
rlabel polysilicon 72 -978 72 -978 0 3
rlabel polysilicon 79 -972 79 -972 0 1
rlabel polysilicon 79 -978 79 -978 0 3
rlabel polysilicon 86 -972 86 -972 0 1
rlabel polysilicon 86 -978 86 -978 0 3
rlabel polysilicon 93 -978 93 -978 0 3
rlabel polysilicon 96 -978 96 -978 0 4
rlabel polysilicon 103 -972 103 -972 0 2
rlabel polysilicon 100 -978 100 -978 0 3
rlabel polysilicon 107 -972 107 -972 0 1
rlabel polysilicon 107 -978 107 -978 0 3
rlabel polysilicon 117 -978 117 -978 0 4
rlabel polysilicon 121 -972 121 -972 0 1
rlabel polysilicon 121 -978 121 -978 0 3
rlabel polysilicon 128 -972 128 -972 0 1
rlabel polysilicon 128 -978 128 -978 0 3
rlabel polysilicon 135 -972 135 -972 0 1
rlabel polysilicon 135 -978 135 -978 0 3
rlabel polysilicon 142 -972 142 -972 0 1
rlabel polysilicon 142 -978 142 -978 0 3
rlabel polysilicon 149 -972 149 -972 0 1
rlabel polysilicon 149 -978 149 -978 0 3
rlabel polysilicon 156 -972 156 -972 0 1
rlabel polysilicon 156 -978 156 -978 0 3
rlabel polysilicon 163 -972 163 -972 0 1
rlabel polysilicon 163 -978 163 -978 0 3
rlabel polysilicon 170 -972 170 -972 0 1
rlabel polysilicon 170 -978 170 -978 0 3
rlabel polysilicon 177 -972 177 -972 0 1
rlabel polysilicon 177 -978 177 -978 0 3
rlabel polysilicon 184 -972 184 -972 0 1
rlabel polysilicon 184 -978 184 -978 0 3
rlabel polysilicon 191 -972 191 -972 0 1
rlabel polysilicon 191 -978 191 -978 0 3
rlabel polysilicon 198 -972 198 -972 0 1
rlabel polysilicon 201 -978 201 -978 0 4
rlabel polysilicon 205 -972 205 -972 0 1
rlabel polysilicon 205 -978 205 -978 0 3
rlabel polysilicon 212 -972 212 -972 0 1
rlabel polysilicon 212 -978 212 -978 0 3
rlabel polysilicon 219 -972 219 -972 0 1
rlabel polysilicon 219 -978 219 -978 0 3
rlabel polysilicon 226 -972 226 -972 0 1
rlabel polysilicon 226 -978 226 -978 0 3
rlabel polysilicon 229 -978 229 -978 0 4
rlabel polysilicon 233 -972 233 -972 0 1
rlabel polysilicon 233 -978 233 -978 0 3
rlabel polysilicon 240 -972 240 -972 0 1
rlabel polysilicon 240 -978 240 -978 0 3
rlabel polysilicon 247 -972 247 -972 0 1
rlabel polysilicon 247 -978 247 -978 0 3
rlabel polysilicon 254 -972 254 -972 0 1
rlabel polysilicon 254 -978 254 -978 0 3
rlabel polysilicon 261 -972 261 -972 0 1
rlabel polysilicon 261 -978 261 -978 0 3
rlabel polysilicon 268 -972 268 -972 0 1
rlabel polysilicon 268 -978 268 -978 0 3
rlabel polysilicon 275 -972 275 -972 0 1
rlabel polysilicon 275 -978 275 -978 0 3
rlabel polysilicon 282 -972 282 -972 0 1
rlabel polysilicon 282 -978 282 -978 0 3
rlabel polysilicon 289 -972 289 -972 0 1
rlabel polysilicon 289 -978 289 -978 0 3
rlabel polysilicon 296 -972 296 -972 0 1
rlabel polysilicon 296 -978 296 -978 0 3
rlabel polysilicon 303 -972 303 -972 0 1
rlabel polysilicon 303 -978 303 -978 0 3
rlabel polysilicon 313 -972 313 -972 0 2
rlabel polysilicon 313 -978 313 -978 0 4
rlabel polysilicon 317 -972 317 -972 0 1
rlabel polysilicon 320 -972 320 -972 0 2
rlabel polysilicon 324 -972 324 -972 0 1
rlabel polysilicon 324 -978 324 -978 0 3
rlabel polysilicon 331 -972 331 -972 0 1
rlabel polysilicon 331 -978 331 -978 0 3
rlabel polysilicon 338 -972 338 -972 0 1
rlabel polysilicon 338 -978 338 -978 0 3
rlabel polysilicon 345 -972 345 -972 0 1
rlabel polysilicon 345 -978 345 -978 0 3
rlabel polysilicon 352 -972 352 -972 0 1
rlabel polysilicon 352 -978 352 -978 0 3
rlabel polysilicon 359 -972 359 -972 0 1
rlabel polysilicon 359 -978 359 -978 0 3
rlabel polysilicon 366 -972 366 -972 0 1
rlabel polysilicon 366 -978 366 -978 0 3
rlabel polysilicon 369 -978 369 -978 0 4
rlabel polysilicon 373 -972 373 -972 0 1
rlabel polysilicon 373 -978 373 -978 0 3
rlabel polysilicon 380 -972 380 -972 0 1
rlabel polysilicon 380 -978 380 -978 0 3
rlabel polysilicon 390 -978 390 -978 0 4
rlabel polysilicon 394 -972 394 -972 0 1
rlabel polysilicon 394 -978 394 -978 0 3
rlabel polysilicon 401 -972 401 -972 0 1
rlabel polysilicon 401 -978 401 -978 0 3
rlabel polysilicon 408 -972 408 -972 0 1
rlabel polysilicon 408 -978 408 -978 0 3
rlabel polysilicon 415 -978 415 -978 0 3
rlabel polysilicon 418 -978 418 -978 0 4
rlabel polysilicon 425 -972 425 -972 0 2
rlabel polysilicon 422 -978 422 -978 0 3
rlabel polysilicon 425 -978 425 -978 0 4
rlabel polysilicon 429 -972 429 -972 0 1
rlabel polysilicon 429 -978 429 -978 0 3
rlabel polysilicon 436 -972 436 -972 0 1
rlabel polysilicon 436 -978 436 -978 0 3
rlabel polysilicon 443 -972 443 -972 0 1
rlabel polysilicon 443 -978 443 -978 0 3
rlabel polysilicon 453 -972 453 -972 0 2
rlabel polysilicon 450 -978 450 -978 0 3
rlabel polysilicon 453 -978 453 -978 0 4
rlabel polysilicon 457 -972 457 -972 0 1
rlabel polysilicon 457 -978 457 -978 0 3
rlabel polysilicon 464 -972 464 -972 0 1
rlabel polysilicon 464 -978 464 -978 0 3
rlabel polysilicon 471 -972 471 -972 0 1
rlabel polysilicon 471 -978 471 -978 0 3
rlabel polysilicon 478 -972 478 -972 0 1
rlabel polysilicon 478 -978 478 -978 0 3
rlabel polysilicon 485 -972 485 -972 0 1
rlabel polysilicon 485 -978 485 -978 0 3
rlabel polysilicon 492 -972 492 -972 0 1
rlabel polysilicon 492 -978 492 -978 0 3
rlabel polysilicon 499 -972 499 -972 0 1
rlabel polysilicon 499 -978 499 -978 0 3
rlabel polysilicon 506 -972 506 -972 0 1
rlabel polysilicon 506 -978 506 -978 0 3
rlabel polysilicon 513 -972 513 -972 0 1
rlabel polysilicon 513 -978 513 -978 0 3
rlabel polysilicon 523 -978 523 -978 0 4
rlabel polysilicon 527 -972 527 -972 0 1
rlabel polysilicon 527 -978 527 -978 0 3
rlabel polysilicon 534 -972 534 -972 0 1
rlabel polysilicon 534 -978 534 -978 0 3
rlabel polysilicon 541 -972 541 -972 0 1
rlabel polysilicon 544 -972 544 -972 0 2
rlabel polysilicon 548 -972 548 -972 0 1
rlabel polysilicon 548 -978 548 -978 0 3
rlabel polysilicon 555 -972 555 -972 0 1
rlabel polysilicon 555 -978 555 -978 0 3
rlabel polysilicon 562 -972 562 -972 0 1
rlabel polysilicon 562 -978 562 -978 0 3
rlabel polysilicon 569 -972 569 -972 0 1
rlabel polysilicon 569 -978 569 -978 0 3
rlabel polysilicon 576 -972 576 -972 0 1
rlabel polysilicon 576 -978 576 -978 0 3
rlabel polysilicon 583 -972 583 -972 0 1
rlabel polysilicon 583 -978 583 -978 0 3
rlabel polysilicon 590 -972 590 -972 0 1
rlabel polysilicon 590 -978 590 -978 0 3
rlabel polysilicon 597 -972 597 -972 0 1
rlabel polysilicon 597 -978 597 -978 0 3
rlabel polysilicon 604 -972 604 -972 0 1
rlabel polysilicon 604 -978 604 -978 0 3
rlabel polysilicon 611 -972 611 -972 0 1
rlabel polysilicon 611 -978 611 -978 0 3
rlabel polysilicon 618 -972 618 -972 0 1
rlabel polysilicon 618 -978 618 -978 0 3
rlabel polysilicon 625 -972 625 -972 0 1
rlabel polysilicon 628 -972 628 -972 0 2
rlabel polysilicon 660 -972 660 -972 0 1
rlabel polysilicon 660 -978 660 -978 0 3
rlabel polysilicon 674 -972 674 -972 0 1
rlabel polysilicon 674 -978 674 -978 0 3
rlabel polysilicon 100 -1011 100 -1011 0 1
rlabel polysilicon 100 -1017 100 -1017 0 3
rlabel polysilicon 142 -1011 142 -1011 0 1
rlabel polysilicon 142 -1017 142 -1017 0 3
rlabel polysilicon 149 -1011 149 -1011 0 1
rlabel polysilicon 149 -1017 149 -1017 0 3
rlabel polysilicon 156 -1011 156 -1011 0 1
rlabel polysilicon 156 -1017 156 -1017 0 3
rlabel polysilicon 163 -1011 163 -1011 0 1
rlabel polysilicon 163 -1017 163 -1017 0 3
rlabel polysilicon 170 -1011 170 -1011 0 1
rlabel polysilicon 170 -1017 170 -1017 0 3
rlabel polysilicon 177 -1011 177 -1011 0 1
rlabel polysilicon 177 -1017 177 -1017 0 3
rlabel polysilicon 184 -1011 184 -1011 0 1
rlabel polysilicon 184 -1017 184 -1017 0 3
rlabel polysilicon 191 -1011 191 -1011 0 1
rlabel polysilicon 191 -1017 191 -1017 0 3
rlabel polysilicon 198 -1011 198 -1011 0 1
rlabel polysilicon 198 -1017 198 -1017 0 3
rlabel polysilicon 205 -1011 205 -1011 0 1
rlabel polysilicon 205 -1017 205 -1017 0 3
rlabel polysilicon 215 -1017 215 -1017 0 4
rlabel polysilicon 219 -1011 219 -1011 0 1
rlabel polysilicon 219 -1017 219 -1017 0 3
rlabel polysilicon 226 -1011 226 -1011 0 1
rlabel polysilicon 226 -1017 226 -1017 0 3
rlabel polysilicon 233 -1011 233 -1011 0 1
rlabel polysilicon 233 -1017 233 -1017 0 3
rlabel polysilicon 240 -1011 240 -1011 0 1
rlabel polysilicon 240 -1017 240 -1017 0 3
rlabel polysilicon 247 -1011 247 -1011 0 1
rlabel polysilicon 250 -1011 250 -1011 0 2
rlabel polysilicon 247 -1017 247 -1017 0 3
rlabel polysilicon 254 -1011 254 -1011 0 1
rlabel polysilicon 254 -1017 254 -1017 0 3
rlabel polysilicon 264 -1011 264 -1011 0 2
rlabel polysilicon 261 -1017 261 -1017 0 3
rlabel polysilicon 264 -1017 264 -1017 0 4
rlabel polysilicon 268 -1011 268 -1011 0 1
rlabel polysilicon 268 -1017 268 -1017 0 3
rlabel polysilicon 275 -1011 275 -1011 0 1
rlabel polysilicon 275 -1017 275 -1017 0 3
rlabel polysilicon 282 -1011 282 -1011 0 1
rlabel polysilicon 282 -1017 282 -1017 0 3
rlabel polysilicon 289 -1011 289 -1011 0 1
rlabel polysilicon 289 -1017 289 -1017 0 3
rlabel polysilicon 299 -1017 299 -1017 0 4
rlabel polysilicon 303 -1011 303 -1011 0 1
rlabel polysilicon 303 -1017 303 -1017 0 3
rlabel polysilicon 310 -1011 310 -1011 0 1
rlabel polysilicon 310 -1017 310 -1017 0 3
rlabel polysilicon 317 -1011 317 -1011 0 1
rlabel polysilicon 317 -1017 317 -1017 0 3
rlabel polysilicon 324 -1011 324 -1011 0 1
rlabel polysilicon 324 -1017 324 -1017 0 3
rlabel polysilicon 331 -1011 331 -1011 0 1
rlabel polysilicon 338 -1011 338 -1011 0 1
rlabel polysilicon 338 -1017 338 -1017 0 3
rlabel polysilicon 345 -1011 345 -1011 0 1
rlabel polysilicon 348 -1017 348 -1017 0 4
rlabel polysilicon 352 -1011 352 -1011 0 1
rlabel polysilicon 352 -1017 352 -1017 0 3
rlabel polysilicon 359 -1011 359 -1011 0 1
rlabel polysilicon 362 -1011 362 -1011 0 2
rlabel polysilicon 359 -1017 359 -1017 0 3
rlabel polysilicon 369 -1011 369 -1011 0 2
rlabel polysilicon 366 -1017 366 -1017 0 3
rlabel polysilicon 373 -1011 373 -1011 0 1
rlabel polysilicon 373 -1017 373 -1017 0 3
rlabel polysilicon 380 -1011 380 -1011 0 1
rlabel polysilicon 380 -1017 380 -1017 0 3
rlabel polysilicon 387 -1011 387 -1011 0 1
rlabel polysilicon 387 -1017 387 -1017 0 3
rlabel polysilicon 394 -1011 394 -1011 0 1
rlabel polysilicon 394 -1017 394 -1017 0 3
rlabel polysilicon 401 -1011 401 -1011 0 1
rlabel polysilicon 401 -1017 401 -1017 0 3
rlabel polysilicon 408 -1011 408 -1011 0 1
rlabel polysilicon 408 -1017 408 -1017 0 3
rlabel polysilicon 415 -1011 415 -1011 0 1
rlabel polysilicon 415 -1017 415 -1017 0 3
rlabel polysilicon 422 -1011 422 -1011 0 1
rlabel polysilicon 422 -1017 422 -1017 0 3
rlabel polysilicon 429 -1011 429 -1011 0 1
rlabel polysilicon 436 -1011 436 -1011 0 1
rlabel polysilicon 439 -1011 439 -1011 0 2
rlabel polysilicon 439 -1017 439 -1017 0 4
rlabel polysilicon 446 -1011 446 -1011 0 2
rlabel polysilicon 443 -1017 443 -1017 0 3
rlabel polysilicon 450 -1011 450 -1011 0 1
rlabel polysilicon 450 -1017 450 -1017 0 3
rlabel polysilicon 457 -1011 457 -1011 0 1
rlabel polysilicon 460 -1017 460 -1017 0 4
rlabel polysilicon 464 -1011 464 -1011 0 1
rlabel polysilicon 464 -1017 464 -1017 0 3
rlabel polysilicon 492 -1011 492 -1011 0 1
rlabel polysilicon 492 -1017 492 -1017 0 3
rlabel polysilicon 499 -1011 499 -1011 0 1
rlabel polysilicon 499 -1017 499 -1017 0 3
rlabel polysilicon 506 -1011 506 -1011 0 1
rlabel polysilicon 506 -1017 506 -1017 0 3
rlabel polysilicon 527 -1011 527 -1011 0 1
rlabel polysilicon 527 -1017 527 -1017 0 3
rlabel polysilicon 544 -1011 544 -1011 0 2
rlabel polysilicon 548 -1011 548 -1011 0 1
rlabel polysilicon 548 -1017 548 -1017 0 3
rlabel polysilicon 569 -1011 569 -1011 0 1
rlabel polysilicon 569 -1017 569 -1017 0 3
rlabel polysilicon 576 -1011 576 -1011 0 1
rlabel polysilicon 576 -1017 576 -1017 0 3
rlabel polysilicon 583 -1011 583 -1011 0 1
rlabel polysilicon 583 -1017 583 -1017 0 3
rlabel polysilicon 590 -1011 590 -1011 0 1
rlabel polysilicon 590 -1017 590 -1017 0 3
rlabel polysilicon 607 -1011 607 -1011 0 2
rlabel polysilicon 604 -1017 604 -1017 0 3
rlabel polysilicon 611 -1011 611 -1011 0 1
rlabel polysilicon 611 -1017 611 -1017 0 3
rlabel polysilicon 646 -1011 646 -1011 0 1
rlabel polysilicon 649 -1011 649 -1011 0 2
rlabel polysilicon 670 -1011 670 -1011 0 2
rlabel polysilicon 100 -1040 100 -1040 0 1
rlabel polysilicon 100 -1046 100 -1046 0 3
rlabel polysilicon 114 -1040 114 -1040 0 1
rlabel polysilicon 114 -1046 114 -1046 0 3
rlabel polysilicon 124 -1040 124 -1040 0 2
rlabel polysilicon 128 -1040 128 -1040 0 1
rlabel polysilicon 128 -1046 128 -1046 0 3
rlabel polysilicon 135 -1040 135 -1040 0 1
rlabel polysilicon 135 -1046 135 -1046 0 3
rlabel polysilicon 142 -1040 142 -1040 0 1
rlabel polysilicon 142 -1046 142 -1046 0 3
rlabel polysilicon 149 -1040 149 -1040 0 1
rlabel polysilicon 149 -1046 149 -1046 0 3
rlabel polysilicon 156 -1040 156 -1040 0 1
rlabel polysilicon 156 -1046 156 -1046 0 3
rlabel polysilicon 163 -1040 163 -1040 0 1
rlabel polysilicon 163 -1046 163 -1046 0 3
rlabel polysilicon 170 -1040 170 -1040 0 1
rlabel polysilicon 173 -1040 173 -1040 0 2
rlabel polysilicon 173 -1046 173 -1046 0 4
rlabel polysilicon 177 -1040 177 -1040 0 1
rlabel polysilicon 180 -1046 180 -1046 0 4
rlabel polysilicon 184 -1046 184 -1046 0 3
rlabel polysilicon 191 -1040 191 -1040 0 1
rlabel polysilicon 191 -1046 191 -1046 0 3
rlabel polysilicon 198 -1040 198 -1040 0 1
rlabel polysilicon 198 -1046 198 -1046 0 3
rlabel polysilicon 205 -1040 205 -1040 0 1
rlabel polysilicon 205 -1046 205 -1046 0 3
rlabel polysilicon 215 -1040 215 -1040 0 2
rlabel polysilicon 212 -1046 212 -1046 0 3
rlabel polysilicon 219 -1040 219 -1040 0 1
rlabel polysilicon 219 -1046 219 -1046 0 3
rlabel polysilicon 229 -1040 229 -1040 0 2
rlabel polysilicon 233 -1040 233 -1040 0 1
rlabel polysilicon 233 -1046 233 -1046 0 3
rlabel polysilicon 243 -1040 243 -1040 0 2
rlabel polysilicon 247 -1040 247 -1040 0 1
rlabel polysilicon 247 -1046 247 -1046 0 3
rlabel polysilicon 254 -1040 254 -1040 0 1
rlabel polysilicon 254 -1046 254 -1046 0 3
rlabel polysilicon 264 -1040 264 -1040 0 2
rlabel polysilicon 268 -1040 268 -1040 0 1
rlabel polysilicon 268 -1046 268 -1046 0 3
rlabel polysilicon 275 -1046 275 -1046 0 3
rlabel polysilicon 278 -1046 278 -1046 0 4
rlabel polysilicon 285 -1046 285 -1046 0 4
rlabel polysilicon 289 -1040 289 -1040 0 1
rlabel polysilicon 289 -1046 289 -1046 0 3
rlabel polysilicon 296 -1040 296 -1040 0 1
rlabel polysilicon 296 -1046 296 -1046 0 3
rlabel polysilicon 306 -1040 306 -1040 0 2
rlabel polysilicon 303 -1046 303 -1046 0 3
rlabel polysilicon 310 -1040 310 -1040 0 1
rlabel polysilicon 310 -1046 310 -1046 0 3
rlabel polysilicon 317 -1040 317 -1040 0 1
rlabel polysilicon 317 -1046 317 -1046 0 3
rlabel polysilicon 366 -1040 366 -1040 0 1
rlabel polysilicon 366 -1046 366 -1046 0 3
rlabel polysilicon 373 -1040 373 -1040 0 1
rlabel polysilicon 376 -1046 376 -1046 0 4
rlabel polysilicon 383 -1046 383 -1046 0 4
rlabel polysilicon 387 -1040 387 -1040 0 1
rlabel polysilicon 387 -1046 387 -1046 0 3
rlabel polysilicon 394 -1040 394 -1040 0 1
rlabel polysilicon 394 -1046 394 -1046 0 3
rlabel polysilicon 404 -1046 404 -1046 0 4
rlabel polysilicon 408 -1040 408 -1040 0 1
rlabel polysilicon 408 -1046 408 -1046 0 3
rlabel polysilicon 418 -1040 418 -1040 0 2
rlabel polysilicon 415 -1046 415 -1046 0 3
rlabel polysilicon 422 -1040 422 -1040 0 1
rlabel polysilicon 422 -1046 422 -1046 0 3
rlabel polysilicon 429 -1040 429 -1040 0 1
rlabel polysilicon 429 -1046 429 -1046 0 3
rlabel polysilicon 436 -1040 436 -1040 0 1
rlabel polysilicon 436 -1046 436 -1046 0 3
rlabel polysilicon 443 -1040 443 -1040 0 1
rlabel polysilicon 443 -1046 443 -1046 0 3
rlabel polysilicon 457 -1040 457 -1040 0 1
rlabel polysilicon 457 -1046 457 -1046 0 3
rlabel polysilicon 474 -1040 474 -1040 0 2
rlabel polysilicon 471 -1046 471 -1046 0 3
rlabel polysilicon 478 -1040 478 -1040 0 1
rlabel polysilicon 478 -1046 478 -1046 0 3
rlabel polysilicon 485 -1040 485 -1040 0 1
rlabel polysilicon 485 -1046 485 -1046 0 3
rlabel polysilicon 541 -1046 541 -1046 0 3
rlabel polysilicon 548 -1040 548 -1040 0 1
rlabel polysilicon 548 -1046 548 -1046 0 3
rlabel polysilicon 562 -1040 562 -1040 0 1
rlabel polysilicon 562 -1046 562 -1046 0 3
rlabel polysilicon 569 -1040 569 -1040 0 1
rlabel polysilicon 569 -1046 569 -1046 0 3
rlabel polysilicon 579 -1046 579 -1046 0 4
rlabel polysilicon 583 -1040 583 -1040 0 1
rlabel polysilicon 583 -1046 583 -1046 0 3
rlabel polysilicon 590 -1040 590 -1040 0 1
rlabel polysilicon 590 -1046 590 -1046 0 3
rlabel polysilicon 100 -1067 100 -1067 0 3
rlabel polysilicon 107 -1061 107 -1061 0 1
rlabel polysilicon 107 -1067 107 -1067 0 3
rlabel polysilicon 135 -1061 135 -1061 0 1
rlabel polysilicon 142 -1061 142 -1061 0 1
rlabel polysilicon 149 -1061 149 -1061 0 1
rlabel polysilicon 149 -1067 149 -1067 0 3
rlabel polysilicon 159 -1067 159 -1067 0 4
rlabel polysilicon 163 -1061 163 -1061 0 1
rlabel polysilicon 163 -1067 163 -1067 0 3
rlabel polysilicon 170 -1067 170 -1067 0 3
rlabel polysilicon 194 -1061 194 -1061 0 2
rlabel polysilicon 198 -1061 198 -1061 0 1
rlabel polysilicon 198 -1067 198 -1067 0 3
rlabel polysilicon 205 -1067 205 -1067 0 3
rlabel polysilicon 215 -1067 215 -1067 0 4
rlabel polysilicon 219 -1067 219 -1067 0 3
rlabel polysilicon 226 -1061 226 -1061 0 1
rlabel polysilicon 226 -1067 226 -1067 0 3
rlabel polysilicon 233 -1061 233 -1061 0 1
rlabel polysilicon 233 -1067 233 -1067 0 3
rlabel polysilicon 282 -1061 282 -1061 0 1
rlabel polysilicon 296 -1061 296 -1061 0 1
rlabel polysilicon 299 -1061 299 -1061 0 2
rlabel polysilicon 380 -1061 380 -1061 0 1
rlabel polysilicon 380 -1067 380 -1067 0 3
rlabel polysilicon 394 -1067 394 -1067 0 3
rlabel polysilicon 411 -1061 411 -1061 0 2
rlabel polysilicon 429 -1061 429 -1061 0 1
rlabel polysilicon 429 -1067 429 -1067 0 3
rlabel polysilicon 439 -1067 439 -1067 0 4
rlabel polysilicon 443 -1061 443 -1061 0 1
rlabel polysilicon 446 -1067 446 -1067 0 4
rlabel polysilicon 453 -1061 453 -1061 0 2
rlabel polysilicon 457 -1061 457 -1061 0 1
rlabel polysilicon 457 -1067 457 -1067 0 3
rlabel polysilicon 562 -1061 562 -1061 0 1
rlabel polysilicon 579 -1061 579 -1061 0 2
rlabel polysilicon 576 -1067 576 -1067 0 3
rlabel polysilicon 583 -1061 583 -1061 0 1
rlabel polysilicon 583 -1067 583 -1067 0 3
rlabel metal2 114 1 114 1 0 net=1727
rlabel metal2 128 1 128 1 0 net=291
rlabel metal2 156 1 156 1 0 net=963
rlabel metal2 177 1 177 1 0 net=1189
rlabel metal2 236 1 236 1 0 net=521
rlabel metal2 296 1 296 1 0 net=2479
rlabel metal2 317 1 317 1 0 net=2007
rlabel metal2 131 -1 131 -1 0 net=259
rlabel metal2 191 -1 191 -1 0 net=425
rlabel metal2 331 -1 331 -1 0 net=2185
rlabel metal2 348 -1 348 -1 0 net=2207
rlabel metal2 135 -3 135 -3 0 net=1559
rlabel metal2 72 -14 72 -14 0 net=2793
rlabel metal2 100 -14 100 -14 0 net=615
rlabel metal2 131 -14 131 -14 0 net=859
rlabel metal2 156 -14 156 -14 0 net=964
rlabel metal2 187 -14 187 -14 0 net=67
rlabel metal2 247 -14 247 -14 0 net=523
rlabel metal2 296 -14 296 -14 0 net=2481
rlabel metal2 331 -14 331 -14 0 net=2187
rlabel metal2 352 -14 352 -14 0 net=2209
rlabel metal2 352 -14 352 -14 0 net=2209
rlabel metal2 373 -14 373 -14 0 net=1309
rlabel metal2 485 -14 485 -14 0 net=2535
rlabel metal2 79 -16 79 -16 0 net=1695
rlabel metal2 107 -16 107 -16 0 net=1561
rlabel metal2 142 -16 142 -16 0 net=427
rlabel metal2 201 -16 201 -16 0 net=1617
rlabel metal2 215 -16 215 -16 0 net=2769
rlabel metal2 296 -16 296 -16 0 net=2009
rlabel metal2 394 -16 394 -16 0 net=1909
rlabel metal2 422 -16 422 -16 0 net=3031
rlabel metal2 117 -18 117 -18 0 net=1728
rlabel metal2 135 -18 135 -18 0 net=515
rlabel metal2 170 -18 170 -18 0 net=1191
rlabel metal2 184 -18 184 -18 0 net=1283
rlabel metal2 219 -18 219 -18 0 net=2033
rlabel metal2 313 -18 313 -18 0 net=1675
rlabel metal2 156 -20 156 -20 0 net=2353
rlabel metal2 229 -20 229 -20 0 net=2343
rlabel metal2 173 -22 173 -22 0 net=1615
rlabel metal2 51 -33 51 -33 0 net=1825
rlabel metal2 65 -33 65 -33 0 net=1257
rlabel metal2 79 -33 79 -33 0 net=1697
rlabel metal2 96 -33 96 -33 0 net=671
rlabel metal2 149 -33 149 -33 0 net=861
rlabel metal2 166 -33 166 -33 0 net=1192
rlabel metal2 184 -33 184 -33 0 net=1285
rlabel metal2 184 -33 184 -33 0 net=1285
rlabel metal2 191 -33 191 -33 0 net=2354
rlabel metal2 233 -33 233 -33 0 net=2771
rlabel metal2 275 -33 275 -33 0 net=1241
rlabel metal2 345 -33 345 -33 0 net=2189
rlabel metal2 387 -33 387 -33 0 net=1911
rlabel metal2 415 -33 415 -33 0 net=2105
rlabel metal2 555 -33 555 -33 0 net=2537
rlabel metal2 65 -35 65 -35 0 net=2795
rlabel metal2 86 -35 86 -35 0 net=617
rlabel metal2 107 -35 107 -35 0 net=1563
rlabel metal2 212 -35 212 -35 0 net=1619
rlabel metal2 233 -35 233 -35 0 net=1343
rlabel metal2 254 -35 254 -35 0 net=524
rlabel metal2 285 -35 285 -35 0 net=2891
rlabel metal2 352 -35 352 -35 0 net=2211
rlabel metal2 380 -35 380 -35 0 net=1961
rlabel metal2 429 -35 429 -35 0 net=3033
rlabel metal2 100 -37 100 -37 0 net=106
rlabel metal2 149 -37 149 -37 0 net=745
rlabel metal2 240 -37 240 -37 0 net=2345
rlabel metal2 261 -37 261 -37 0 net=2347
rlabel metal2 261 -37 261 -37 0 net=2347
rlabel metal2 289 -37 289 -37 0 net=1197
rlabel metal2 327 -37 327 -37 0 net=2901
rlabel metal2 359 -37 359 -37 0 net=915
rlabel metal2 436 -37 436 -37 0 net=1311
rlabel metal2 107 -39 107 -39 0 net=749
rlabel metal2 296 -39 296 -39 0 net=2011
rlabel metal2 296 -39 296 -39 0 net=2011
rlabel metal2 303 -39 303 -39 0 net=2483
rlabel metal2 331 -39 331 -39 0 net=1677
rlabel metal2 156 -41 156 -41 0 net=571
rlabel metal2 254 -41 254 -41 0 net=1215
rlabel metal2 159 -43 159 -43 0 net=1616
rlabel metal2 194 -43 194 -43 0 net=1817
rlabel metal2 282 -43 282 -43 0 net=2035
rlabel metal2 121 -45 121 -45 0 net=367
rlabel metal2 177 -45 177 -45 0 net=2197
rlabel metal2 121 -47 121 -47 0 net=517
rlabel metal2 135 -49 135 -49 0 net=429
rlabel metal2 142 -51 142 -51 0 net=909
rlabel metal2 30 -62 30 -62 0 net=409
rlabel metal2 156 -62 156 -62 0 net=1564
rlabel metal2 191 -62 191 -62 0 net=2772
rlabel metal2 366 -62 366 -62 0 net=2191
rlabel metal2 425 -62 425 -62 0 net=1877
rlabel metal2 471 -62 471 -62 0 net=1989
rlabel metal2 530 -62 530 -62 0 net=2323
rlabel metal2 37 -64 37 -64 0 net=1827
rlabel metal2 58 -64 58 -64 0 net=1079
rlabel metal2 93 -64 93 -64 0 net=1699
rlabel metal2 233 -64 233 -64 0 net=1345
rlabel metal2 373 -64 373 -64 0 net=2213
rlabel metal2 443 -64 443 -64 0 net=3035
rlabel metal2 576 -64 576 -64 0 net=2539
rlabel metal2 576 -64 576 -64 0 net=2539
rlabel metal2 44 -66 44 -66 0 net=431
rlabel metal2 142 -66 142 -66 0 net=911
rlabel metal2 240 -66 240 -66 0 net=2346
rlabel metal2 261 -66 261 -66 0 net=2348
rlabel metal2 303 -66 303 -66 0 net=1151
rlabel metal2 380 -66 380 -66 0 net=1913
rlabel metal2 401 -66 401 -66 0 net=2617
rlabel metal2 51 -68 51 -68 0 net=519
rlabel metal2 131 -68 131 -68 0 net=1725
rlabel metal2 198 -68 198 -68 0 net=573
rlabel metal2 198 -68 198 -68 0 net=573
rlabel metal2 205 -68 205 -68 0 net=1819
rlabel metal2 240 -68 240 -68 0 net=1216
rlabel metal2 261 -68 261 -68 0 net=1199
rlabel metal2 387 -68 387 -68 0 net=1963
rlabel metal2 401 -68 401 -68 0 net=2107
rlabel metal2 450 -68 450 -68 0 net=1313
rlabel metal2 450 -68 450 -68 0 net=1313
rlabel metal2 457 -68 457 -68 0 net=185
rlabel metal2 457 -68 457 -68 0 net=185
rlabel metal2 65 -70 65 -70 0 net=2796
rlabel metal2 100 -70 100 -70 0 net=2198
rlabel metal2 289 -70 289 -70 0 net=917
rlabel metal2 72 -72 72 -72 0 net=1258
rlabel metal2 86 -72 86 -72 0 net=619
rlabel metal2 107 -72 107 -72 0 net=751
rlabel metal2 107 -72 107 -72 0 net=751
rlabel metal2 114 -72 114 -72 0 net=673
rlabel metal2 114 -72 114 -72 0 net=673
rlabel metal2 128 -72 128 -72 0 net=1217
rlabel metal2 324 -72 324 -72 0 net=2485
rlabel metal2 65 -74 65 -74 0 net=1033
rlabel metal2 128 -74 128 -74 0 net=2417
rlabel metal2 313 -74 313 -74 0 net=1843
rlabel metal2 331 -74 331 -74 0 net=2037
rlabel metal2 72 -76 72 -76 0 net=875
rlabel metal2 296 -76 296 -76 0 net=2013
rlabel metal2 345 -76 345 -76 0 net=2903
rlabel metal2 131 -78 131 -78 0 net=799
rlabel metal2 142 -78 142 -78 0 net=1287
rlabel metal2 219 -78 219 -78 0 net=1621
rlabel metal2 313 -78 313 -78 0 net=2751
rlabel metal2 149 -80 149 -80 0 net=747
rlabel metal2 219 -80 219 -80 0 net=871
rlabel metal2 345 -80 345 -80 0 net=1369
rlabel metal2 163 -82 163 -82 0 net=863
rlabel metal2 163 -84 163 -84 0 net=663
rlabel metal2 184 -86 184 -86 0 net=1243
rlabel metal2 275 -88 275 -88 0 net=2893
rlabel metal2 338 -90 338 -90 0 net=1679
rlabel metal2 9 -101 9 -101 0 net=1829
rlabel metal2 51 -101 51 -101 0 net=520
rlabel metal2 128 -101 128 -101 0 net=581
rlabel metal2 282 -101 282 -101 0 net=2349
rlabel metal2 555 -101 555 -101 0 net=2541
rlabel metal2 590 -101 590 -101 0 net=2325
rlabel metal2 16 -103 16 -103 0 net=1081
rlabel metal2 65 -103 65 -103 0 net=621
rlabel metal2 121 -103 121 -103 0 net=701
rlabel metal2 170 -103 170 -103 0 net=1726
rlabel metal2 331 -103 331 -103 0 net=2015
rlabel metal2 460 -103 460 -103 0 net=2071
rlabel metal2 26 -105 26 -105 0 net=202
rlabel metal2 75 -105 75 -105 0 net=545
rlabel metal2 173 -105 173 -105 0 net=748
rlabel metal2 240 -105 240 -105 0 net=2603
rlabel metal2 30 -107 30 -107 0 net=410
rlabel metal2 100 -107 100 -107 0 net=753
rlabel metal2 149 -107 149 -107 0 net=1403
rlabel metal2 243 -107 243 -107 0 net=1346
rlabel metal2 282 -107 282 -107 0 net=919
rlabel metal2 313 -107 313 -107 0 net=2904
rlabel metal2 366 -107 366 -107 0 net=2589
rlabel metal2 37 -109 37 -109 0 net=711
rlabel metal2 86 -109 86 -109 0 net=1035
rlabel metal2 191 -109 191 -109 0 net=575
rlabel metal2 226 -109 226 -109 0 net=1701
rlabel metal2 275 -109 275 -109 0 net=2894
rlabel metal2 338 -109 338 -109 0 net=1681
rlabel metal2 366 -109 366 -109 0 net=1315
rlabel metal2 478 -109 478 -109 0 net=2619
rlabel metal2 30 -111 30 -111 0 net=807
rlabel metal2 345 -111 345 -111 0 net=1371
rlabel metal2 355 -111 355 -111 0 net=2895
rlabel metal2 51 -113 51 -113 0 net=1715
rlabel metal2 107 -113 107 -113 0 net=675
rlabel metal2 142 -113 142 -113 0 net=1289
rlabel metal2 345 -113 345 -113 0 net=2109
rlabel metal2 415 -113 415 -113 0 net=2487
rlabel metal2 58 -115 58 -115 0 net=541
rlabel metal2 114 -115 114 -115 0 net=697
rlabel metal2 142 -115 142 -115 0 net=665
rlabel metal2 198 -115 198 -115 0 net=913
rlabel metal2 226 -115 226 -115 0 net=1121
rlabel metal2 492 -115 492 -115 0 net=3037
rlabel metal2 205 -117 205 -117 0 net=865
rlabel metal2 233 -117 233 -117 0 net=1821
rlabel metal2 415 -117 415 -117 0 net=2649
rlabel metal2 499 -117 499 -117 0 net=2277
rlabel metal2 520 -117 520 -117 0 net=2263
rlabel metal2 135 -119 135 -119 0 net=801
rlabel metal2 247 -119 247 -119 0 net=2419
rlabel metal2 44 -121 44 -121 0 net=433
rlabel metal2 205 -121 205 -121 0 net=873
rlabel metal2 247 -121 247 -121 0 net=1153
rlabel metal2 373 -121 373 -121 0 net=2333
rlabel metal2 44 -123 44 -123 0 net=877
rlabel metal2 184 -123 184 -123 0 net=1245
rlabel metal2 320 -123 320 -123 0 net=1419
rlabel metal2 387 -123 387 -123 0 net=1965
rlabel metal2 72 -125 72 -125 0 net=1363
rlabel metal2 394 -125 394 -125 0 net=2039
rlabel metal2 159 -127 159 -127 0 net=815
rlabel metal2 219 -127 219 -127 0 net=141
rlabel metal2 261 -127 261 -127 0 net=1200
rlabel metal2 324 -127 324 -127 0 net=1845
rlabel metal2 422 -127 422 -127 0 net=1879
rlabel metal2 170 -129 170 -129 0 net=140
rlabel metal2 296 -129 296 -129 0 net=1623
rlabel metal2 408 -129 408 -129 0 net=2193
rlabel metal2 177 -131 177 -131 0 net=1219
rlabel metal2 310 -131 310 -131 0 net=1111
rlabel metal2 408 -131 408 -131 0 net=1991
rlabel metal2 166 -133 166 -133 0 net=595
rlabel metal2 429 -133 429 -133 0 net=2215
rlabel metal2 429 -135 429 -135 0 net=1787
rlabel metal2 436 -137 436 -137 0 net=2753
rlabel metal2 380 -139 380 -139 0 net=1915
rlabel metal2 443 -139 443 -139 0 net=2373
rlabel metal2 257 -141 257 -141 0 net=1475
rlabel metal2 443 -141 443 -141 0 net=1573
rlabel metal2 23 -152 23 -152 0 net=577
rlabel metal2 205 -152 205 -152 0 net=874
rlabel metal2 261 -152 261 -152 0 net=2590
rlabel metal2 611 -152 611 -152 0 net=3039
rlabel metal2 51 -154 51 -154 0 net=1716
rlabel metal2 184 -154 184 -154 0 net=816
rlabel metal2 450 -154 450 -154 0 net=1967
rlabel metal2 450 -154 450 -154 0 net=1967
rlabel metal2 464 -154 464 -154 0 net=2195
rlabel metal2 51 -156 51 -156 0 net=583
rlabel metal2 142 -156 142 -156 0 net=667
rlabel metal2 191 -156 191 -156 0 net=833
rlabel metal2 306 -156 306 -156 0 net=2040
rlabel metal2 618 -156 618 -156 0 net=2326
rlabel metal2 628 -156 628 -156 0 net=2849
rlabel metal2 65 -158 65 -158 0 net=622
rlabel metal2 100 -158 100 -158 0 net=755
rlabel metal2 135 -158 135 -158 0 net=435
rlabel metal2 156 -158 156 -158 0 net=547
rlabel metal2 173 -158 173 -158 0 net=914
rlabel metal2 212 -158 212 -158 0 net=867
rlabel metal2 313 -158 313 -158 0 net=2072
rlabel metal2 604 -158 604 -158 0 net=2897
rlabel metal2 58 -160 58 -160 0 net=543
rlabel metal2 72 -160 72 -160 0 net=95
rlabel metal2 198 -160 198 -160 0 net=1155
rlabel metal2 254 -160 254 -160 0 net=1221
rlabel metal2 334 -160 334 -160 0 net=1549
rlabel metal2 16 -162 16 -162 0 net=1083
rlabel metal2 79 -162 79 -162 0 net=1101
rlabel metal2 212 -162 212 -162 0 net=983
rlabel metal2 278 -162 278 -162 0 net=2488
rlabel metal2 541 -162 541 -162 0 net=2375
rlabel metal2 576 -162 576 -162 0 net=2621
rlabel metal2 16 -164 16 -164 0 net=879
rlabel metal2 79 -164 79 -164 0 net=677
rlabel metal2 135 -164 135 -164 0 net=218
rlabel metal2 387 -164 387 -164 0 net=1847
rlabel metal2 44 -166 44 -166 0 net=921
rlabel metal2 289 -166 289 -166 0 net=1113
rlabel metal2 387 -166 387 -166 0 net=2321
rlabel metal2 82 -168 82 -168 0 net=10
rlabel metal2 100 -168 100 -168 0 net=1822
rlabel metal2 436 -168 436 -168 0 net=1917
rlabel metal2 471 -168 471 -168 0 net=2631
rlabel metal2 86 -170 86 -170 0 net=1036
rlabel metal2 215 -170 215 -170 0 net=1624
rlabel metal2 457 -170 457 -170 0 net=2017
rlabel metal2 562 -170 562 -170 0 net=2605
rlabel metal2 86 -172 86 -172 0 net=699
rlabel metal2 149 -172 149 -172 0 net=2351
rlabel metal2 555 -172 555 -172 0 net=2543
rlabel metal2 107 -174 107 -174 0 net=703
rlabel metal2 219 -174 219 -174 0 net=1290
rlabel metal2 341 -174 341 -174 0 net=1937
rlabel metal2 485 -174 485 -174 0 net=2755
rlabel metal2 30 -176 30 -176 0 net=809
rlabel metal2 233 -176 233 -176 0 net=803
rlabel metal2 233 -176 233 -176 0 net=803
rlabel metal2 247 -176 247 -176 0 net=1201
rlabel metal2 30 -178 30 -178 0 net=1405
rlabel metal2 268 -178 268 -178 0 net=1703
rlabel metal2 422 -178 422 -178 0 net=1881
rlabel metal2 492 -178 492 -178 0 net=2651
rlabel metal2 37 -180 37 -180 0 net=713
rlabel metal2 222 -180 222 -180 0 net=2203
rlabel metal2 499 -180 499 -180 0 net=2335
rlabel metal2 520 -180 520 -180 0 net=2265
rlabel metal2 37 -182 37 -182 0 net=1145
rlabel metal2 114 -182 114 -182 0 net=1123
rlabel metal2 240 -182 240 -182 0 net=489
rlabel metal2 282 -182 282 -182 0 net=945
rlabel metal2 390 -182 390 -182 0 net=2987
rlabel metal2 177 -184 177 -184 0 net=597
rlabel metal2 296 -184 296 -184 0 net=1476
rlabel metal2 488 -184 488 -184 0 net=2905
rlabel metal2 520 -184 520 -184 0 net=1763
rlabel metal2 177 -186 177 -186 0 net=228
rlabel metal2 317 -186 317 -186 0 net=2383
rlabel metal2 268 -188 268 -188 0 net=899
rlabel metal2 320 -188 320 -188 0 net=1851
rlabel metal2 506 -188 506 -188 0 net=2279
rlabel metal2 548 -188 548 -188 0 net=2421
rlabel metal2 359 -190 359 -190 0 net=1683
rlabel metal2 331 -192 331 -192 0 net=1365
rlabel metal2 366 -192 366 -192 0 net=1317
rlabel metal2 415 -192 415 -192 0 net=2823
rlabel metal2 331 -194 331 -194 0 net=2399
rlabel metal2 345 -196 345 -196 0 net=2111
rlabel metal2 478 -196 478 -196 0 net=2217
rlabel metal2 170 -198 170 -198 0 net=1233
rlabel metal2 373 -198 373 -198 0 net=1421
rlabel metal2 408 -198 408 -198 0 net=1993
rlabel metal2 9 -200 9 -200 0 net=1831
rlabel metal2 352 -200 352 -200 0 net=1373
rlabel metal2 408 -200 408 -200 0 net=1789
rlabel metal2 303 -202 303 -202 0 net=1247
rlabel metal2 429 -202 429 -202 0 net=1575
rlabel metal2 23 -213 23 -213 0 net=579
rlabel metal2 219 -213 219 -213 0 net=811
rlabel metal2 219 -213 219 -213 0 net=811
rlabel metal2 275 -213 275 -213 0 net=2018
rlabel metal2 548 -213 548 -213 0 net=2825
rlabel metal2 23 -215 23 -215 0 net=1041
rlabel metal2 100 -215 100 -215 0 net=704
rlabel metal2 142 -215 142 -215 0 net=437
rlabel metal2 142 -215 142 -215 0 net=437
rlabel metal2 152 -215 152 -215 0 net=270
rlabel metal2 292 -215 292 -215 0 net=2199
rlabel metal2 548 -215 548 -215 0 net=2633
rlabel metal2 653 -215 653 -215 0 net=2989
rlabel metal2 44 -217 44 -217 0 net=923
rlabel metal2 103 -217 103 -217 0 net=804
rlabel metal2 296 -217 296 -217 0 net=1576
rlabel metal2 446 -217 446 -217 0 net=2377
rlabel metal2 660 -217 660 -217 0 net=3041
rlabel metal2 44 -219 44 -219 0 net=2089
rlabel metal2 58 -219 58 -219 0 net=1085
rlabel metal2 58 -219 58 -219 0 net=1085
rlabel metal2 65 -219 65 -219 0 net=544
rlabel metal2 86 -219 86 -219 0 net=700
rlabel metal2 156 -219 156 -219 0 net=1102
rlabel metal2 303 -219 303 -219 0 net=1249
rlabel metal2 369 -219 369 -219 0 net=2322
rlabel metal2 51 -221 51 -221 0 net=585
rlabel metal2 86 -221 86 -221 0 net=1017
rlabel metal2 313 -221 313 -221 0 net=2376
rlabel metal2 583 -221 583 -221 0 net=2423
rlabel metal2 51 -223 51 -223 0 net=2352
rlabel metal2 163 -223 163 -223 0 net=549
rlabel metal2 163 -223 163 -223 0 net=549
rlabel metal2 170 -223 170 -223 0 net=1833
rlabel metal2 331 -223 331 -223 0 net=2196
rlabel metal2 37 -225 37 -225 0 net=1147
rlabel metal2 338 -225 338 -225 0 net=1367
rlabel metal2 369 -225 369 -225 0 net=3003
rlabel metal2 590 -225 590 -225 0 net=2623
rlabel metal2 9 -227 9 -227 0 net=1063
rlabel metal2 65 -227 65 -227 0 net=953
rlabel metal2 128 -227 128 -227 0 net=757
rlabel metal2 177 -227 177 -227 0 net=868
rlabel metal2 341 -227 341 -227 0 net=1684
rlabel metal2 499 -227 499 -227 0 net=2337
rlabel metal2 611 -227 611 -227 0 net=2653
rlabel metal2 16 -229 16 -229 0 net=881
rlabel metal2 191 -229 191 -229 0 net=835
rlabel metal2 233 -229 233 -229 0 net=491
rlabel metal2 254 -229 254 -229 0 net=1223
rlabel metal2 387 -229 387 -229 0 net=2756
rlabel metal2 16 -231 16 -231 0 net=1087
rlabel metal2 128 -231 128 -231 0 net=669
rlabel metal2 191 -231 191 -231 0 net=599
rlabel metal2 254 -231 254 -231 0 net=901
rlabel metal2 299 -231 299 -231 0 net=2143
rlabel metal2 30 -233 30 -233 0 net=1406
rlabel metal2 345 -233 345 -233 0 net=1235
rlabel metal2 422 -233 422 -233 0 net=2205
rlabel metal2 33 -235 33 -235 0 net=539
rlabel metal2 247 -235 247 -235 0 net=1203
rlabel metal2 408 -235 408 -235 0 net=1791
rlabel metal2 457 -235 457 -235 0 net=1883
rlabel metal2 488 -235 488 -235 0 net=2606
rlabel metal2 79 -237 79 -237 0 net=679
rlabel metal2 198 -237 198 -237 0 net=1156
rlabel metal2 247 -237 247 -237 0 net=2773
rlabel metal2 2 -239 2 -239 0 net=2103
rlabel metal2 107 -239 107 -239 0 net=1361
rlabel metal2 464 -239 464 -239 0 net=1919
rlabel metal2 513 -239 513 -239 0 net=2907
rlabel metal2 121 -241 121 -241 0 net=715
rlabel metal2 198 -241 198 -241 0 net=1115
rlabel metal2 299 -241 299 -241 0 net=1643
rlabel metal2 471 -241 471 -241 0 net=1939
rlabel metal2 513 -241 513 -241 0 net=1849
rlabel metal2 121 -243 121 -243 0 net=555
rlabel metal2 268 -243 268 -243 0 net=947
rlabel metal2 327 -243 327 -243 0 net=2057
rlabel metal2 471 -243 471 -243 0 net=1995
rlabel metal2 527 -243 527 -243 0 net=2281
rlabel metal2 135 -245 135 -245 0 net=623
rlabel metal2 366 -245 366 -245 0 net=2087
rlabel metal2 555 -245 555 -245 0 net=2385
rlabel metal2 250 -247 250 -247 0 net=2515
rlabel metal2 562 -247 562 -247 0 net=2545
rlabel metal2 261 -249 261 -249 0 net=985
rlabel metal2 380 -249 380 -249 0 net=1423
rlabel metal2 436 -249 436 -249 0 net=1853
rlabel metal2 506 -249 506 -249 0 net=2219
rlabel metal2 576 -249 576 -249 0 net=2401
rlabel metal2 380 -251 380 -251 0 net=2850
rlabel metal2 383 -253 383 -253 0 net=2697
rlabel metal2 394 -255 394 -255 0 net=1705
rlabel metal2 506 -255 506 -255 0 net=1551
rlabel metal2 394 -257 394 -257 0 net=1319
rlabel metal2 541 -257 541 -257 0 net=2267
rlabel metal2 625 -257 625 -257 0 net=2899
rlabel metal2 373 -259 373 -259 0 net=1375
rlabel metal2 415 -259 415 -259 0 net=2113
rlabel metal2 646 -259 646 -259 0 net=2613
rlabel metal2 30 -261 30 -261 0 net=1253
rlabel metal2 443 -261 443 -261 0 net=2431
rlabel metal2 317 -263 317 -263 0 net=1625
rlabel metal2 443 -263 443 -263 0 net=1969
rlabel metal2 114 -265 114 -265 0 net=1125
rlabel metal2 450 -265 450 -265 0 net=1765
rlabel metal2 520 -267 520 -267 0 net=1823
rlabel metal2 23 -278 23 -278 0 net=1042
rlabel metal2 58 -278 58 -278 0 net=1086
rlabel metal2 128 -278 128 -278 0 net=670
rlabel metal2 289 -278 289 -278 0 net=1225
rlabel metal2 362 -278 362 -278 0 net=2114
rlabel metal2 569 -278 569 -278 0 net=3005
rlabel metal2 26 -280 26 -280 0 net=540
rlabel metal2 240 -280 240 -280 0 net=2088
rlabel metal2 534 -280 534 -280 0 net=2201
rlabel metal2 576 -280 576 -280 0 net=2269
rlabel metal2 576 -280 576 -280 0 net=2269
rlabel metal2 604 -280 604 -280 0 net=2387
rlabel metal2 604 -280 604 -280 0 net=2387
rlabel metal2 716 -280 716 -280 0 net=3043
rlabel metal2 2 -282 2 -282 0 net=2104
rlabel metal2 247 -282 247 -282 0 net=1250
rlabel metal2 310 -282 310 -282 0 net=1368
rlabel metal2 345 -282 345 -282 0 net=1205
rlabel metal2 373 -282 373 -282 0 net=1255
rlabel metal2 373 -282 373 -282 0 net=1255
rlabel metal2 380 -282 380 -282 0 net=2144
rlabel metal2 30 -284 30 -284 0 net=587
rlabel metal2 82 -284 82 -284 0 net=2900
rlabel metal2 16 -286 16 -286 0 net=1089
rlabel metal2 86 -286 86 -286 0 net=1019
rlabel metal2 310 -286 310 -286 0 net=1047
rlabel metal2 338 -286 338 -286 0 net=1627
rlabel metal2 422 -286 422 -286 0 net=1793
rlabel metal2 467 -286 467 -286 0 net=2634
rlabel metal2 639 -286 639 -286 0 net=2625
rlabel metal2 667 -286 667 -286 0 net=2775
rlabel metal2 16 -288 16 -288 0 net=837
rlabel metal2 212 -288 212 -288 0 net=580
rlabel metal2 292 -288 292 -288 0 net=2977
rlabel metal2 33 -290 33 -290 0 net=2145
rlabel metal2 541 -290 541 -290 0 net=2339
rlabel metal2 653 -290 653 -290 0 net=2699
rlabel metal2 37 -292 37 -292 0 net=1065
rlabel metal2 100 -292 100 -292 0 net=681
rlabel metal2 198 -292 198 -292 0 net=1116
rlabel metal2 380 -292 380 -292 0 net=1377
rlabel metal2 422 -292 422 -292 0 net=1553
rlabel metal2 548 -292 548 -292 0 net=2221
rlabel metal2 590 -292 590 -292 0 net=2403
rlabel metal2 44 -294 44 -294 0 net=2091
rlabel metal2 555 -294 555 -294 0 net=2517
rlabel metal2 47 -296 47 -296 0 net=1706
rlabel metal2 478 -296 478 -296 0 net=1855
rlabel metal2 478 -296 478 -296 0 net=1855
rlabel metal2 485 -296 485 -296 0 net=1885
rlabel metal2 485 -296 485 -296 0 net=1885
rlabel metal2 492 -296 492 -296 0 net=1921
rlabel metal2 492 -296 492 -296 0 net=1921
rlabel metal2 499 -296 499 -296 0 net=1941
rlabel metal2 555 -296 555 -296 0 net=2379
rlabel metal2 51 -298 51 -298 0 net=445
rlabel metal2 107 -298 107 -298 0 net=605
rlabel metal2 212 -298 212 -298 0 net=1513
rlabel metal2 394 -298 394 -298 0 net=1321
rlabel metal2 432 -298 432 -298 0 net=1824
rlabel metal2 562 -298 562 -298 0 net=2283
rlabel metal2 597 -298 597 -298 0 net=2433
rlabel metal2 54 -300 54 -300 0 net=116
rlabel metal2 121 -300 121 -300 0 net=557
rlabel metal2 135 -300 135 -300 0 net=625
rlabel metal2 156 -300 156 -300 0 net=759
rlabel metal2 257 -300 257 -300 0 net=2449
rlabel metal2 625 -300 625 -300 0 net=2547
rlabel metal2 58 -302 58 -302 0 net=189
rlabel metal2 345 -302 345 -302 0 net=2908
rlabel metal2 65 -304 65 -304 0 net=954
rlabel metal2 191 -304 191 -304 0 net=601
rlabel metal2 219 -304 219 -304 0 net=813
rlabel metal2 261 -304 261 -304 0 net=2783
rlabel metal2 65 -306 65 -306 0 net=949
rlabel metal2 299 -306 299 -306 0 net=2969
rlabel metal2 93 -308 93 -308 0 net=925
rlabel metal2 299 -308 299 -308 0 net=1850
rlabel metal2 583 -308 583 -308 0 net=2425
rlabel metal2 632 -308 632 -308 0 net=2615
rlabel metal2 110 -310 110 -310 0 net=641
rlabel metal2 121 -310 121 -310 0 net=965
rlabel metal2 394 -310 394 -310 0 net=1425
rlabel metal2 436 -310 436 -310 0 net=1585
rlabel metal2 135 -312 135 -312 0 net=717
rlabel metal2 191 -312 191 -312 0 net=987
rlabel metal2 401 -312 401 -312 0 net=2206
rlabel metal2 37 -314 37 -314 0 net=453
rlabel metal2 275 -314 275 -314 0 net=2729
rlabel metal2 646 -314 646 -314 0 net=2655
rlabel metal2 695 -314 695 -314 0 net=2991
rlabel metal2 44 -316 44 -316 0 net=2955
rlabel metal2 93 -318 93 -318 0 net=1171
rlabel metal2 443 -318 443 -318 0 net=1971
rlabel metal2 660 -318 660 -318 0 net=2827
rlabel metal2 142 -320 142 -320 0 net=439
rlabel metal2 177 -320 177 -320 0 net=883
rlabel metal2 275 -320 275 -320 0 net=1515
rlabel metal2 457 -320 457 -320 0 net=2059
rlabel metal2 142 -322 142 -322 0 net=501
rlabel metal2 324 -322 324 -322 0 net=1835
rlabel metal2 471 -322 471 -322 0 net=1997
rlabel metal2 156 -324 156 -324 0 net=493
rlabel metal2 324 -324 324 -324 0 net=1362
rlabel metal2 450 -324 450 -324 0 net=1767
rlabel metal2 51 -326 51 -326 0 net=1535
rlabel metal2 278 -326 278 -326 0 net=1525
rlabel metal2 429 -326 429 -326 0 net=1645
rlabel metal2 163 -328 163 -328 0 net=551
rlabel metal2 327 -328 327 -328 0 net=2951
rlabel metal2 177 -330 177 -330 0 net=903
rlabel metal2 331 -330 331 -330 0 net=1149
rlabel metal2 317 -332 317 -332 0 net=1127
rlabel metal2 429 -332 429 -332 0 net=2971
rlabel metal2 317 -334 317 -334 0 net=1237
rlabel metal2 5 -345 5 -345 0 net=1161
rlabel metal2 369 -345 369 -345 0 net=1856
rlabel metal2 555 -345 555 -345 0 net=2381
rlabel metal2 23 -347 23 -347 0 net=705
rlabel metal2 373 -347 373 -347 0 net=1256
rlabel metal2 373 -347 373 -347 0 net=1256
rlabel metal2 376 -347 376 -347 0 net=2995
rlabel metal2 26 -349 26 -349 0 net=1646
rlabel metal2 474 -349 474 -349 0 net=2887
rlabel metal2 30 -351 30 -351 0 net=589
rlabel metal2 187 -351 187 -351 0 net=814
rlabel metal2 261 -351 261 -351 0 net=885
rlabel metal2 261 -351 261 -351 0 net=885
rlabel metal2 268 -351 268 -351 0 net=926
rlabel metal2 282 -351 282 -351 0 net=2202
rlabel metal2 667 -351 667 -351 0 net=2777
rlabel metal2 30 -353 30 -353 0 net=495
rlabel metal2 219 -353 219 -353 0 net=552
rlabel metal2 268 -353 268 -353 0 net=1837
rlabel metal2 513 -353 513 -353 0 net=1999
rlabel metal2 583 -353 583 -353 0 net=2427
rlabel metal2 674 -353 674 -353 0 net=2785
rlabel metal2 2 -355 2 -355 0 net=2077
rlabel metal2 688 -355 688 -355 0 net=2953
rlabel metal2 44 -357 44 -357 0 net=741
rlabel metal2 408 -357 408 -357 0 net=1517
rlabel metal2 464 -357 464 -357 0 net=1795
rlabel metal2 527 -357 527 -357 0 net=2093
rlabel metal2 695 -357 695 -357 0 net=2957
rlabel metal2 47 -359 47 -359 0 net=158
rlabel metal2 324 -359 324 -359 0 net=1179
rlabel metal2 352 -359 352 -359 0 net=1207
rlabel metal2 408 -359 408 -359 0 net=1323
rlabel metal2 432 -359 432 -359 0 net=2992
rlabel metal2 730 -359 730 -359 0 net=3007
rlabel metal2 51 -361 51 -361 0 net=989
rlabel metal2 219 -361 219 -361 0 net=1150
rlabel metal2 485 -361 485 -361 0 net=1887
rlabel metal2 558 -361 558 -361 0 net=3051
rlabel metal2 54 -363 54 -363 0 net=92
rlabel metal2 415 -363 415 -363 0 net=3044
rlabel metal2 61 -365 61 -365 0 net=103
rlabel metal2 233 -365 233 -365 0 net=1536
rlabel metal2 422 -365 422 -365 0 net=1555
rlabel metal2 471 -365 471 -365 0 net=1769
rlabel metal2 562 -365 562 -365 0 net=2285
rlabel metal2 562 -365 562 -365 0 net=2285
rlabel metal2 618 -365 618 -365 0 net=2731
rlabel metal2 709 -365 709 -365 0 net=2973
rlabel metal2 72 -367 72 -367 0 net=1091
rlabel metal2 247 -367 247 -367 0 net=1629
rlabel metal2 345 -367 345 -367 0 net=2970
rlabel metal2 716 -367 716 -367 0 net=2979
rlabel metal2 72 -369 72 -369 0 net=447
rlabel metal2 93 -369 93 -369 0 net=1173
rlabel metal2 282 -369 282 -369 0 net=1129
rlabel metal2 338 -369 338 -369 0 net=1497
rlabel metal2 625 -369 625 -369 0 net=2549
rlabel metal2 37 -371 37 -371 0 net=454
rlabel metal2 348 -371 348 -371 0 net=2719
rlabel metal2 79 -373 79 -373 0 net=1067
rlabel metal2 226 -373 226 -373 0 net=1157
rlabel metal2 387 -373 387 -373 0 net=1527
rlabel metal2 429 -373 429 -373 0 net=2229
rlabel metal2 639 -373 639 -373 0 net=2627
rlabel metal2 79 -375 79 -375 0 net=905
rlabel metal2 226 -375 226 -375 0 net=1239
rlabel metal2 348 -375 348 -375 0 net=2743
rlabel metal2 86 -377 86 -377 0 net=719
rlabel metal2 149 -377 149 -377 0 net=627
rlabel metal2 149 -377 149 -377 0 net=627
rlabel metal2 285 -377 285 -377 0 net=38
rlabel metal2 541 -377 541 -377 0 net=2341
rlabel metal2 646 -377 646 -377 0 net=2657
rlabel metal2 93 -379 93 -379 0 net=525
rlabel metal2 436 -379 436 -379 0 net=1587
rlabel metal2 492 -379 492 -379 0 net=1923
rlabel metal2 576 -379 576 -379 0 net=2271
rlabel metal2 646 -379 646 -379 0 net=2829
rlabel metal2 681 -379 681 -379 0 net=2519
rlabel metal2 100 -381 100 -381 0 net=683
rlabel metal2 289 -381 289 -381 0 net=1227
rlabel metal2 394 -381 394 -381 0 net=1427
rlabel metal2 492 -381 492 -381 0 net=1973
rlabel metal2 520 -381 520 -381 0 net=2061
rlabel metal2 590 -381 590 -381 0 net=2405
rlabel metal2 100 -383 100 -383 0 net=607
rlabel metal2 292 -383 292 -383 0 net=1359
rlabel metal2 590 -383 590 -383 0 net=2435
rlabel metal2 611 -383 611 -383 0 net=2451
rlabel metal2 107 -385 107 -385 0 net=2616
rlabel metal2 653 -385 653 -385 0 net=2701
rlabel metal2 110 -387 110 -387 0 net=1291
rlabel metal2 296 -387 296 -387 0 net=1021
rlabel metal2 310 -387 310 -387 0 net=1049
rlabel metal2 534 -387 534 -387 0 net=2147
rlabel metal2 604 -387 604 -387 0 net=2389
rlabel metal2 110 -389 110 -389 0 net=1759
rlabel metal2 548 -389 548 -389 0 net=2223
rlabel metal2 121 -391 121 -391 0 net=967
rlabel metal2 222 -391 222 -391 0 net=1043
rlabel metal2 383 -391 383 -391 0 net=2167
rlabel metal2 124 -393 124 -393 0 net=1073
rlabel metal2 163 -393 163 -393 0 net=216
rlabel metal2 299 -393 299 -393 0 net=1977
rlabel metal2 114 -395 114 -395 0 net=643
rlabel metal2 303 -395 303 -395 0 net=1037
rlabel metal2 401 -395 401 -395 0 net=1891
rlabel metal2 37 -397 37 -397 0 net=1707
rlabel metal2 506 -397 506 -397 0 net=1943
rlabel metal2 114 -399 114 -399 0 net=761
rlabel metal2 128 -401 128 -401 0 net=559
rlabel metal2 240 -401 240 -401 0 net=1379
rlabel metal2 128 -403 128 -403 0 net=503
rlabel metal2 212 -403 212 -403 0 net=1514
rlabel metal2 16 -405 16 -405 0 net=839
rlabel metal2 16 -407 16 -407 0 net=603
rlabel metal2 142 -409 142 -409 0 net=441
rlabel metal2 198 -409 198 -409 0 net=1449
rlabel metal2 65 -411 65 -411 0 net=951
rlabel metal2 58 -413 58 -413 0 net=1259
rlabel metal2 9 -424 9 -424 0 net=990
rlabel metal2 58 -424 58 -424 0 net=2149
rlabel metal2 72 -424 72 -424 0 net=448
rlabel metal2 170 -424 170 -424 0 net=952
rlabel metal2 264 -424 264 -424 0 net=2786
rlabel metal2 9 -426 9 -426 0 net=743
rlabel metal2 47 -426 47 -426 0 net=2428
rlabel metal2 702 -426 702 -426 0 net=2629
rlabel metal2 51 -428 51 -428 0 net=609
rlabel metal2 107 -428 107 -428 0 net=2094
rlabel metal2 702 -428 702 -428 0 net=2779
rlabel metal2 58 -430 58 -430 0 net=2382
rlabel metal2 61 -432 61 -432 0 net=1838
rlabel metal2 275 -432 275 -432 0 net=1175
rlabel metal2 380 -432 380 -432 0 net=2406
rlabel metal2 730 -432 730 -432 0 net=2521
rlabel metal2 72 -434 72 -434 0 net=1451
rlabel metal2 205 -434 205 -434 0 net=969
rlabel metal2 334 -434 334 -434 0 net=2148
rlabel metal2 611 -434 611 -434 0 net=2391
rlabel metal2 716 -434 716 -434 0 net=2703
rlabel metal2 79 -436 79 -436 0 net=907
rlabel metal2 338 -436 338 -436 0 net=2224
rlabel metal2 79 -438 79 -438 0 net=1023
rlabel metal2 348 -438 348 -438 0 net=2720
rlabel metal2 86 -440 86 -440 0 net=721
rlabel metal2 163 -440 163 -440 0 net=645
rlabel metal2 233 -440 233 -440 0 net=1093
rlabel metal2 366 -440 366 -440 0 net=1208
rlabel metal2 394 -440 394 -440 0 net=2342
rlabel metal2 646 -440 646 -440 0 net=2831
rlabel metal2 44 -442 44 -442 0 net=1347
rlabel metal2 254 -442 254 -442 0 net=1293
rlabel metal2 387 -442 387 -442 0 net=1229
rlabel metal2 401 -442 401 -442 0 net=1978
rlabel metal2 709 -442 709 -442 0 net=2659
rlabel metal2 86 -444 86 -444 0 net=1163
rlabel metal2 404 -444 404 -444 0 net=2980
rlabel metal2 93 -446 93 -446 0 net=527
rlabel metal2 170 -446 170 -446 0 net=851
rlabel metal2 226 -446 226 -446 0 net=1240
rlabel metal2 436 -446 436 -446 0 net=1429
rlabel metal2 436 -446 436 -446 0 net=1429
rlabel metal2 443 -446 443 -446 0 net=1557
rlabel metal2 618 -446 618 -446 0 net=2231
rlabel metal2 695 -446 695 -446 0 net=2551
rlabel metal2 793 -446 793 -446 0 net=3009
rlabel metal2 93 -448 93 -448 0 net=957
rlabel metal2 352 -448 352 -448 0 net=1159
rlabel metal2 450 -448 450 -448 0 net=1499
rlabel metal2 450 -448 450 -448 0 net=1499
rlabel metal2 474 -448 474 -448 0 net=2954
rlabel metal2 100 -450 100 -450 0 net=268
rlabel metal2 474 -450 474 -450 0 net=2305
rlabel metal2 681 -450 681 -450 0 net=2453
rlabel metal2 772 -450 772 -450 0 net=2975
rlabel metal2 107 -452 107 -452 0 net=505
rlabel metal2 198 -452 198 -452 0 net=1051
rlabel metal2 324 -452 324 -452 0 net=1181
rlabel metal2 355 -452 355 -452 0 net=2123
rlabel metal2 625 -452 625 -452 0 net=2273
rlabel metal2 786 -452 786 -452 0 net=2997
rlabel metal2 30 -454 30 -454 0 net=497
rlabel metal2 191 -454 191 -454 0 net=1069
rlabel metal2 506 -454 506 -454 0 net=2041
rlabel metal2 604 -454 604 -454 0 net=2169
rlabel metal2 800 -454 800 -454 0 net=3053
rlabel metal2 30 -456 30 -456 0 net=1537
rlabel metal2 520 -456 520 -456 0 net=2744
rlabel metal2 37 -458 37 -458 0 net=1709
rlabel metal2 523 -458 523 -458 0 net=2888
rlabel metal2 37 -460 37 -460 0 net=629
rlabel metal2 212 -460 212 -460 0 net=841
rlabel metal2 261 -460 261 -460 0 net=887
rlabel metal2 303 -460 303 -460 0 net=1039
rlabel metal2 418 -460 418 -460 0 net=1743
rlabel metal2 541 -460 541 -460 0 net=1925
rlabel metal2 558 -460 558 -460 0 net=2803
rlabel metal2 765 -460 765 -460 0 net=2959
rlabel metal2 110 -462 110 -462 0 net=613
rlabel metal2 222 -462 222 -462 0 net=2981
rlabel metal2 135 -464 135 -464 0 net=685
rlabel metal2 247 -464 247 -464 0 net=1631
rlabel metal2 541 -464 541 -464 0 net=2079
rlabel metal2 590 -464 590 -464 0 net=2437
rlabel metal2 688 -464 688 -464 0 net=2733
rlabel metal2 149 -466 149 -466 0 net=779
rlabel metal2 562 -466 562 -466 0 net=2287
rlabel metal2 705 -466 705 -466 0 net=1
rlabel metal2 247 -468 247 -468 0 net=1131
rlabel metal2 303 -468 303 -468 0 net=1360
rlabel metal2 492 -468 492 -468 0 net=1975
rlabel metal2 569 -468 569 -468 0 net=2001
rlabel metal2 282 -470 282 -470 0 net=1045
rlabel metal2 380 -470 380 -470 0 net=2441
rlabel metal2 16 -472 16 -472 0 net=604
rlabel metal2 422 -472 422 -472 0 net=1529
rlabel metal2 492 -472 492 -472 0 net=2315
rlabel metal2 16 -474 16 -474 0 net=1109
rlabel metal2 422 -474 422 -474 0 net=1589
rlabel metal2 548 -474 548 -474 0 net=1945
rlabel metal2 576 -474 576 -474 0 net=2063
rlabel metal2 415 -476 415 -476 0 net=1875
rlabel metal2 527 -476 527 -476 0 net=1889
rlabel metal2 555 -476 555 -476 0 net=1947
rlabel metal2 408 -478 408 -478 0 net=1325
rlabel metal2 485 -478 485 -478 0 net=1771
rlabel metal2 485 -480 485 -480 0 net=1893
rlabel metal2 457 -482 457 -482 0 net=1519
rlabel metal2 457 -484 457 -484 0 net=1797
rlabel metal2 499 -486 499 -486 0 net=1761
rlabel metal2 331 -488 331 -488 0 net=1639
rlabel metal2 156 -490 156 -490 0 net=1075
rlabel metal2 156 -492 156 -492 0 net=591
rlabel metal2 142 -494 142 -494 0 net=443
rlabel metal2 142 -496 142 -496 0 net=561
rlabel metal2 23 -498 23 -498 0 net=707
rlabel metal2 23 -500 23 -500 0 net=1381
rlabel metal2 65 -502 65 -502 0 net=1261
rlabel metal2 65 -504 65 -504 0 net=763
rlabel metal2 114 -506 114 -506 0 net=1193
rlabel metal2 9 -517 9 -517 0 net=744
rlabel metal2 163 -517 163 -517 0 net=528
rlabel metal2 467 -517 467 -517 0 net=2976
rlabel metal2 793 -517 793 -517 0 net=3011
rlabel metal2 9 -519 9 -519 0 net=533
rlabel metal2 163 -519 163 -519 0 net=709
rlabel metal2 184 -519 184 -519 0 net=444
rlabel metal2 222 -519 222 -519 0 net=1520
rlabel metal2 555 -519 555 -519 0 net=1949
rlabel metal2 583 -519 583 -519 0 net=1927
rlabel metal2 16 -521 16 -521 0 net=1110
rlabel metal2 313 -521 313 -521 0 net=1160
rlabel metal2 380 -521 380 -521 0 net=314
rlabel metal2 618 -521 618 -521 0 net=2125
rlabel metal2 681 -521 681 -521 0 net=2439
rlabel metal2 681 -521 681 -521 0 net=2439
rlabel metal2 709 -521 709 -521 0 net=2553
rlabel metal2 709 -521 709 -521 0 net=2553
rlabel metal2 779 -521 779 -521 0 net=2983
rlabel metal2 800 -521 800 -521 0 net=3055
rlabel metal2 16 -523 16 -523 0 net=1501
rlabel metal2 471 -523 471 -523 0 net=1061
rlabel metal2 495 -523 495 -523 0 net=2780
rlabel metal2 758 -523 758 -523 0 net=2833
rlabel metal2 786 -523 786 -523 0 net=2999
rlabel metal2 44 -525 44 -525 0 net=927
rlabel metal2 135 -525 135 -525 0 net=1565
rlabel metal2 457 -525 457 -525 0 net=1799
rlabel metal2 520 -525 520 -525 0 net=1745
rlabel metal2 541 -525 541 -525 0 net=2081
rlabel metal2 618 -525 618 -525 0 net=2289
rlabel metal2 744 -525 744 -525 0 net=2523
rlabel metal2 765 -525 765 -525 0 net=2961
rlabel metal2 47 -527 47 -527 0 net=1076
rlabel metal2 383 -527 383 -527 0 net=1890
rlabel metal2 54 -529 54 -529 0 net=614
rlabel metal2 226 -529 226 -529 0 net=908
rlabel metal2 303 -529 303 -529 0 net=955
rlabel metal2 317 -529 317 -529 0 net=1040
rlabel metal2 383 -529 383 -529 0 net=1976
rlabel metal2 625 -529 625 -529 0 net=2151
rlabel metal2 58 -531 58 -531 0 net=959
rlabel metal2 131 -531 131 -531 0 net=935
rlabel metal2 212 -531 212 -531 0 net=687
rlabel metal2 233 -531 233 -531 0 net=1349
rlabel metal2 387 -531 387 -531 0 net=2429
rlabel metal2 61 -533 61 -533 0 net=449
rlabel metal2 121 -533 121 -533 0 net=723
rlabel metal2 240 -533 240 -533 0 net=1263
rlabel metal2 390 -533 390 -533 0 net=1762
rlabel metal2 520 -533 520 -533 0 net=1773
rlabel metal2 541 -533 541 -533 0 net=2003
rlabel metal2 625 -533 625 -533 0 net=2233
rlabel metal2 79 -535 79 -535 0 net=1025
rlabel metal2 240 -535 240 -535 0 net=1177
rlabel metal2 394 -535 394 -535 0 net=1231
rlabel metal2 429 -535 429 -535 0 net=2704
rlabel metal2 79 -537 79 -537 0 net=647
rlabel metal2 257 -537 257 -537 0 net=1046
rlabel metal2 310 -537 310 -537 0 net=2797
rlabel metal2 51 -539 51 -539 0 net=611
rlabel metal2 275 -539 275 -539 0 net=1685
rlabel metal2 345 -539 345 -539 0 net=1183
rlabel metal2 401 -539 401 -539 0 net=2051
rlabel metal2 639 -539 639 -539 0 net=2307
rlabel metal2 30 -541 30 -541 0 net=1539
rlabel metal2 401 -541 401 -541 0 net=1327
rlabel metal2 422 -541 422 -541 0 net=1591
rlabel metal2 457 -541 457 -541 0 net=2630
rlabel metal2 30 -543 30 -543 0 net=1053
rlabel metal2 282 -543 282 -543 0 net=1711
rlabel metal2 562 -543 562 -543 0 net=2043
rlabel metal2 86 -545 86 -545 0 net=1165
rlabel metal2 369 -545 369 -545 0 net=2593
rlabel metal2 86 -547 86 -547 0 net=659
rlabel metal2 317 -547 317 -547 0 net=2411
rlabel metal2 93 -549 93 -549 0 net=853
rlabel metal2 177 -549 177 -549 0 net=889
rlabel metal2 415 -549 415 -549 0 net=1558
rlabel metal2 114 -551 114 -551 0 net=1195
rlabel metal2 422 -551 422 -551 0 net=1431
rlabel metal2 474 -551 474 -551 0 net=1946
rlabel metal2 597 -551 597 -551 0 net=2171
rlabel metal2 23 -553 23 -553 0 net=1383
rlabel metal2 135 -553 135 -553 0 net=991
rlabel metal2 436 -553 436 -553 0 net=1531
rlabel metal2 478 -553 478 -553 0 net=1876
rlabel metal2 569 -553 569 -553 0 net=2065
rlabel metal2 611 -553 611 -553 0 net=2661
rlabel metal2 23 -555 23 -555 0 net=1070
rlabel metal2 411 -555 411 -555 0 net=2591
rlabel metal2 149 -557 149 -557 0 net=781
rlabel metal2 324 -557 324 -557 0 net=1095
rlabel metal2 443 -557 443 -557 0 net=1633
rlabel metal2 485 -557 485 -557 0 net=1895
rlabel metal2 604 -557 604 -557 0 net=2393
rlabel metal2 72 -559 72 -559 0 net=1453
rlabel metal2 488 -559 488 -559 0 net=2529
rlabel metal2 142 -561 142 -561 0 net=563
rlabel metal2 156 -561 156 -561 0 net=593
rlabel metal2 296 -561 296 -561 0 net=1295
rlabel metal2 499 -561 499 -561 0 net=1641
rlabel metal2 37 -563 37 -563 0 net=631
rlabel metal2 170 -563 170 -563 0 net=971
rlabel metal2 464 -563 464 -563 0 net=2599
rlabel metal2 506 -563 506 -563 0 net=2097
rlabel metal2 632 -563 632 -563 0 net=2275
rlabel metal2 674 -563 674 -563 0 net=2805
rlabel metal2 37 -565 37 -565 0 net=507
rlabel metal2 198 -565 198 -565 0 net=483
rlabel metal2 646 -565 646 -565 0 net=2317
rlabel metal2 737 -565 737 -565 0 net=2735
rlabel metal2 65 -567 65 -567 0 net=765
rlabel metal2 289 -567 289 -567 0 net=1103
rlabel metal2 667 -567 667 -567 0 net=2443
rlabel metal2 65 -569 65 -569 0 net=1133
rlabel metal2 418 -569 418 -569 0 net=2609
rlabel metal2 128 -571 128 -571 0 net=499
rlabel metal2 688 -571 688 -571 0 net=2455
rlabel metal2 72 -573 72 -573 0 net=529
rlabel metal2 247 -573 247 -573 0 net=843
rlabel metal2 334 -573 334 -573 0 net=2721
rlabel metal2 184 -575 184 -575 0 net=553
rlabel metal2 2 -586 2 -586 0 net=531
rlabel metal2 86 -586 86 -586 0 net=661
rlabel metal2 86 -586 86 -586 0 net=661
rlabel metal2 93 -586 93 -586 0 net=855
rlabel metal2 93 -586 93 -586 0 net=855
rlabel metal2 107 -586 107 -586 0 net=632
rlabel metal2 163 -586 163 -586 0 net=710
rlabel metal2 436 -586 436 -586 0 net=1533
rlabel metal2 436 -586 436 -586 0 net=1533
rlabel metal2 457 -586 457 -586 0 net=1950
rlabel metal2 9 -588 9 -588 0 net=534
rlabel metal2 296 -588 296 -588 0 net=1196
rlabel metal2 464 -588 464 -588 0 net=51
rlabel metal2 513 -588 513 -588 0 net=2276
rlabel metal2 9 -590 9 -590 0 net=2821
rlabel metal2 334 -590 334 -590 0 net=1642
rlabel metal2 54 -592 54 -592 0 net=1540
rlabel metal2 467 -592 467 -592 0 net=2052
rlabel metal2 730 -592 730 -592 0 net=3013
rlabel metal2 68 -594 68 -594 0 net=1712
rlabel metal2 299 -594 299 -594 0 net=500
rlabel metal2 485 -594 485 -594 0 net=2440
rlabel metal2 72 -596 72 -596 0 net=451
rlabel metal2 107 -596 107 -596 0 net=2152
rlabel metal2 100 -598 100 -598 0 net=1011
rlabel metal2 506 -598 506 -598 0 net=2126
rlabel metal2 110 -600 110 -600 0 net=554
rlabel metal2 205 -600 205 -600 0 net=612
rlabel metal2 271 -600 271 -600 0 net=1477
rlabel metal2 460 -600 460 -600 0 net=2685
rlabel metal2 110 -602 110 -602 0 net=1178
rlabel metal2 254 -602 254 -602 0 net=2567
rlabel metal2 653 -602 653 -602 0 net=2611
rlabel metal2 121 -604 121 -604 0 net=1232
rlabel metal2 506 -604 506 -604 0 net=2005
rlabel metal2 576 -604 576 -604 0 net=2663
rlabel metal2 737 -604 737 -604 0 net=2985
rlabel metal2 121 -606 121 -606 0 net=891
rlabel metal2 184 -606 184 -606 0 net=1635
rlabel metal2 513 -606 513 -606 0 net=2045
rlabel metal2 611 -606 611 -606 0 net=2457
rlabel metal2 26 -608 26 -608 0 net=2705
rlabel metal2 124 -610 124 -610 0 net=2430
rlabel metal2 128 -612 128 -612 0 net=973
rlabel metal2 177 -612 177 -612 0 net=1105
rlabel metal2 303 -612 303 -612 0 net=956
rlabel metal2 320 -612 320 -612 0 net=1521
rlabel metal2 478 -612 478 -612 0 net=1801
rlabel metal2 534 -612 534 -612 0 net=1747
rlabel metal2 562 -612 562 -612 0 net=2291
rlabel metal2 772 -612 772 -612 0 net=3001
rlabel metal2 138 -614 138 -614 0 net=766
rlabel metal2 149 -614 149 -614 0 net=565
rlabel metal2 331 -614 331 -614 0 net=1185
rlabel metal2 492 -614 492 -614 0 net=1897
rlabel metal2 534 -614 534 -614 0 net=2099
rlabel metal2 618 -614 618 -614 0 net=2531
rlabel metal2 37 -616 37 -616 0 net=508
rlabel metal2 156 -616 156 -616 0 net=467
rlabel metal2 303 -616 303 -616 0 net=1351
rlabel metal2 366 -616 366 -616 0 net=3056
rlabel metal2 30 -618 30 -618 0 net=1055
rlabel metal2 61 -618 61 -618 0 net=1117
rlabel metal2 163 -618 163 -618 0 net=689
rlabel metal2 240 -618 240 -618 0 net=845
rlabel metal2 282 -618 282 -618 0 net=1097
rlabel metal2 359 -618 359 -618 0 net=1433
rlabel metal2 527 -618 527 -618 0 net=2083
rlabel metal2 590 -618 590 -618 0 net=2413
rlabel metal2 702 -618 702 -618 0 net=2737
rlabel metal2 170 -620 170 -620 0 net=2647
rlabel metal2 289 -620 289 -620 0 net=1869
rlabel metal2 583 -620 583 -620 0 net=2395
rlabel metal2 751 -620 751 -620 0 net=2963
rlabel metal2 191 -622 191 -622 0 net=937
rlabel metal2 310 -622 310 -622 0 net=2234
rlabel metal2 191 -624 191 -624 0 net=1717
rlabel metal2 348 -624 348 -624 0 net=2757
rlabel metal2 205 -626 205 -626 0 net=725
rlabel metal2 275 -626 275 -626 0 net=1687
rlabel metal2 324 -626 324 -626 0 net=1167
rlabel metal2 373 -626 373 -626 0 net=1455
rlabel metal2 453 -626 453 -626 0 net=194
rlabel metal2 198 -628 198 -628 0 net=485
rlabel metal2 268 -628 268 -628 0 net=993
rlabel metal2 338 -628 338 -628 0 net=1297
rlabel metal2 422 -628 422 -628 0 net=1593
rlabel metal2 443 -628 443 -628 0 net=2129
rlabel metal2 548 -628 548 -628 0 net=2679
rlabel metal2 625 -628 625 -628 0 net=2555
rlabel metal2 65 -630 65 -630 0 net=1135
rlabel metal2 212 -630 212 -630 0 net=594
rlabel metal2 338 -630 338 -630 0 net=1265
rlabel metal2 548 -630 548 -630 0 net=2173
rlabel metal2 709 -630 709 -630 0 net=2835
rlabel metal2 30 -632 30 -632 0 net=461
rlabel metal2 215 -632 215 -632 0 net=2592
rlabel metal2 758 -632 758 -632 0 net=2525
rlabel metal2 219 -634 219 -634 0 net=1027
rlabel metal2 380 -634 380 -634 0 net=2857
rlabel metal2 758 -634 758 -634 0 net=2927
rlabel metal2 51 -636 51 -636 0 net=791
rlabel metal2 226 -636 226 -636 0 net=782
rlabel metal2 383 -636 383 -636 0 net=1661
rlabel metal2 597 -636 597 -636 0 net=2445
rlabel metal2 44 -638 44 -638 0 net=929
rlabel metal2 383 -638 383 -638 0 net=2259
rlabel metal2 646 -638 646 -638 0 net=2319
rlabel metal2 44 -640 44 -640 0 net=639
rlabel metal2 387 -640 387 -640 0 net=1329
rlabel metal2 646 -640 646 -640 0 net=2723
rlabel metal2 16 -642 16 -642 0 net=1503
rlabel metal2 499 -642 499 -642 0 net=2601
rlabel metal2 16 -644 16 -644 0 net=961
rlabel metal2 499 -644 499 -644 0 net=2309
rlabel metal2 58 -646 58 -646 0 net=330
rlabel metal2 639 -646 639 -646 0 net=2595
rlabel metal2 79 -648 79 -648 0 net=649
rlabel metal2 674 -648 674 -648 0 net=2807
rlabel metal2 79 -650 79 -650 0 net=1385
rlabel metal2 674 -650 674 -650 0 net=2799
rlabel metal2 23 -652 23 -652 0 net=190
rlabel metal2 415 -652 415 -652 0 net=3045
rlabel metal2 23 -654 23 -654 0 net=1567
rlabel metal2 415 -656 415 -656 0 net=2861
rlabel metal2 450 -658 450 -658 0 net=1062
rlabel metal2 471 -660 471 -660 0 net=1775
rlabel metal2 520 -662 520 -662 0 net=2067
rlabel metal2 569 -664 569 -664 0 net=1929
rlabel metal2 2 -675 2 -675 0 net=532
rlabel metal2 100 -675 100 -675 0 net=1013
rlabel metal2 100 -675 100 -675 0 net=1013
rlabel metal2 142 -675 142 -675 0 net=65
rlabel metal2 425 -675 425 -675 0 net=2006
rlabel metal2 520 -675 520 -675 0 net=2068
rlabel metal2 551 -675 551 -675 0 net=2758
rlabel metal2 751 -675 751 -675 0 net=2965
rlabel metal2 751 -675 751 -675 0 net=2965
rlabel metal2 765 -675 765 -675 0 net=3047
rlabel metal2 765 -675 765 -675 0 net=3047
rlabel metal2 779 -675 779 -675 0 net=2527
rlabel metal2 16 -677 16 -677 0 net=962
rlabel metal2 142 -677 142 -677 0 net=691
rlabel metal2 177 -677 177 -677 0 net=1107
rlabel metal2 177 -677 177 -677 0 net=1107
rlabel metal2 184 -677 184 -677 0 net=1636
rlabel metal2 415 -677 415 -677 0 net=1534
rlabel metal2 446 -677 446 -677 0 net=2084
rlabel metal2 625 -677 625 -677 0 net=2557
rlabel metal2 625 -677 625 -677 0 net=2557
rlabel metal2 639 -677 639 -677 0 net=2597
rlabel metal2 639 -677 639 -677 0 net=2597
rlabel metal2 660 -677 660 -677 0 net=2801
rlabel metal2 779 -677 779 -677 0 net=3057
rlabel metal2 16 -679 16 -679 0 net=856
rlabel metal2 107 -679 107 -679 0 net=2019
rlabel metal2 450 -679 450 -679 0 net=1871
rlabel metal2 499 -679 499 -679 0 net=2311
rlabel metal2 527 -679 527 -679 0 net=2836
rlabel metal2 51 -681 51 -681 0 net=662
rlabel metal2 107 -681 107 -681 0 net=417
rlabel metal2 271 -681 271 -681 0 net=2320
rlabel metal2 37 -683 37 -683 0 net=1057
rlabel metal2 58 -683 58 -683 0 net=893
rlabel metal2 149 -683 149 -683 0 net=1119
rlabel metal2 212 -683 212 -683 0 net=566
rlabel metal2 415 -683 415 -683 0 net=1663
rlabel metal2 453 -683 453 -683 0 net=2612
rlabel metal2 9 -685 9 -685 0 net=2822
rlabel metal2 457 -685 457 -685 0 net=2261
rlabel metal2 471 -685 471 -685 0 net=1777
rlabel metal2 37 -687 37 -687 0 net=1387
rlabel metal2 93 -687 93 -687 0 net=1209
rlabel metal2 296 -687 296 -687 0 net=3002
rlabel metal2 61 -689 61 -689 0 net=2648
rlabel metal2 198 -689 198 -689 0 net=1137
rlabel metal2 310 -689 310 -689 0 net=1689
rlabel metal2 443 -689 443 -689 0 net=2131
rlabel metal2 485 -689 485 -689 0 net=1899
rlabel metal2 499 -689 499 -689 0 net=2047
rlabel metal2 604 -689 604 -689 0 net=2681
rlabel metal2 772 -689 772 -689 0 net=3059
rlabel metal2 12 -691 12 -691 0 net=2363
rlabel metal2 443 -691 443 -691 0 net=2986
rlabel metal2 68 -693 68 -693 0 net=1637
rlabel metal2 114 -693 114 -693 0 net=783
rlabel metal2 135 -693 135 -693 0 net=651
rlabel metal2 156 -693 156 -693 0 net=469
rlabel metal2 156 -693 156 -693 0 net=469
rlabel metal2 170 -693 170 -693 0 net=931
rlabel metal2 268 -693 268 -693 0 net=1805
rlabel metal2 460 -693 460 -693 0 net=3025
rlabel metal2 72 -695 72 -695 0 net=452
rlabel metal2 198 -695 198 -695 0 net=847
rlabel metal2 261 -695 261 -695 0 net=1353
rlabel metal2 464 -695 464 -695 0 net=2101
rlabel metal2 583 -695 583 -695 0 net=2397
rlabel metal2 646 -695 646 -695 0 net=2725
rlabel metal2 23 -697 23 -697 0 net=1569
rlabel metal2 114 -697 114 -697 0 net=975
rlabel metal2 135 -697 135 -697 0 net=401
rlabel metal2 233 -697 233 -697 0 net=487
rlabel metal2 303 -697 303 -697 0 net=2225
rlabel metal2 492 -697 492 -697 0 net=1931
rlabel metal2 583 -697 583 -697 0 net=2459
rlabel metal2 646 -697 646 -697 0 net=2739
rlabel metal2 23 -699 23 -699 0 net=1719
rlabel metal2 212 -699 212 -699 0 net=939
rlabel metal2 513 -699 513 -699 0 net=1749
rlabel metal2 590 -699 590 -699 0 net=2415
rlabel metal2 618 -699 618 -699 0 net=2533
rlabel metal2 44 -701 44 -701 0 net=640
rlabel metal2 191 -701 191 -701 0 net=727
rlabel metal2 226 -701 226 -701 0 net=2851
rlabel metal2 44 -703 44 -703 0 net=535
rlabel metal2 205 -703 205 -703 0 net=793
rlabel metal2 229 -703 229 -703 0 net=207
rlabel metal2 534 -703 534 -703 0 net=2157
rlabel metal2 30 -705 30 -705 0 net=462
rlabel metal2 219 -705 219 -705 0 net=1523
rlabel metal2 544 -705 544 -705 0 net=2491
rlabel metal2 618 -705 618 -705 0 net=2707
rlabel metal2 30 -707 30 -707 0 net=1169
rlabel metal2 345 -707 345 -707 0 net=1647
rlabel metal2 555 -707 555 -707 0 net=2293
rlabel metal2 597 -707 597 -707 0 net=2447
rlabel metal2 233 -709 233 -709 0 net=1029
rlabel metal2 254 -709 254 -709 0 net=1267
rlabel metal2 380 -709 380 -709 0 net=2602
rlabel metal2 240 -711 240 -711 0 net=995
rlabel metal2 324 -711 324 -711 0 net=1435
rlabel metal2 597 -711 597 -711 0 net=2569
rlabel metal2 653 -711 653 -711 0 net=2687
rlabel metal2 695 -711 695 -711 0 net=2809
rlabel metal2 166 -713 166 -713 0 net=1463
rlabel metal2 478 -713 478 -713 0 net=1803
rlabel metal2 247 -715 247 -715 0 net=1187
rlabel metal2 338 -715 338 -715 0 net=1299
rlabel metal2 478 -715 478 -715 0 net=2175
rlabel metal2 576 -715 576 -715 0 net=2665
rlabel metal2 681 -715 681 -715 0 net=2859
rlabel metal2 275 -717 275 -717 0 net=1099
rlabel metal2 331 -717 331 -717 0 net=1331
rlabel metal2 530 -717 530 -717 0 net=2327
rlabel metal2 723 -717 723 -717 0 net=2863
rlabel metal2 282 -719 282 -719 0 net=1479
rlabel metal2 744 -719 744 -719 0 net=2929
rlabel metal2 320 -721 320 -721 0 net=1577
rlabel metal2 394 -721 394 -721 0 net=2235
rlabel metal2 730 -721 730 -721 0 net=3015
rlabel metal2 131 -723 131 -723 0 net=2909
rlabel metal2 352 -725 352 -725 0 net=1457
rlabel metal2 373 -727 373 -727 0 net=1505
rlabel metal2 401 -729 401 -729 0 net=1595
rlabel metal2 422 -731 422 -731 0 net=2245
rlabel metal2 2 -742 2 -742 0 net=569
rlabel metal2 268 -742 268 -742 0 net=1100
rlabel metal2 289 -742 289 -742 0 net=488
rlabel metal2 397 -742 397 -742 0 net=2102
rlabel metal2 481 -742 481 -742 0 net=400
rlabel metal2 572 -742 572 -742 0 net=3026
rlabel metal2 765 -742 765 -742 0 net=3049
rlabel metal2 765 -742 765 -742 0 net=3049
rlabel metal2 782 -742 782 -742 0 net=2528
rlabel metal2 793 -742 793 -742 0 net=3058
rlabel metal2 9 -744 9 -744 0 net=1839
rlabel metal2 166 -744 166 -744 0 net=1524
rlabel metal2 268 -744 268 -744 0 net=1579
rlabel metal2 422 -744 422 -744 0 net=2534
rlabel metal2 737 -744 737 -744 0 net=2931
rlabel metal2 16 -746 16 -746 0 net=895
rlabel metal2 65 -746 65 -746 0 net=1571
rlabel metal2 79 -746 79 -746 0 net=1638
rlabel metal2 345 -746 345 -746 0 net=2448
rlabel metal2 702 -746 702 -746 0 net=2865
rlabel metal2 744 -746 744 -746 0 net=2967
rlabel metal2 30 -748 30 -748 0 net=1170
rlabel metal2 275 -748 275 -748 0 net=1139
rlabel metal2 310 -748 310 -748 0 net=2365
rlabel metal2 366 -748 366 -748 0 net=1807
rlabel metal2 506 -748 506 -748 0 net=2237
rlabel metal2 576 -748 576 -748 0 net=2329
rlabel metal2 19 -750 19 -750 0 net=2635
rlabel metal2 376 -750 376 -750 0 net=1979
rlabel metal2 513 -750 513 -750 0 net=1751
rlabel metal2 513 -750 513 -750 0 net=1751
rlabel metal2 520 -750 520 -750 0 net=2295
rlabel metal2 562 -750 562 -750 0 net=2313
rlabel metal2 562 -750 562 -750 0 net=2313
rlabel metal2 600 -750 600 -750 0 net=2802
rlabel metal2 751 -750 751 -750 0 net=3017
rlabel metal2 30 -752 30 -752 0 net=537
rlabel metal2 58 -752 58 -752 0 net=785
rlabel metal2 184 -752 184 -752 0 net=1120
rlabel metal2 233 -752 233 -752 0 net=1031
rlabel metal2 310 -752 310 -752 0 net=1458
rlabel metal2 380 -752 380 -752 0 net=2889
rlabel metal2 758 -752 758 -752 0 net=3061
rlabel metal2 40 -754 40 -754 0 net=1857
rlabel metal2 184 -754 184 -754 0 net=941
rlabel metal2 282 -754 282 -754 0 net=1481
rlabel metal2 408 -754 408 -754 0 net=1649
rlabel metal2 446 -754 446 -754 0 net=2935
rlabel metal2 772 -754 772 -754 0 net=2053
rlabel metal2 44 -756 44 -756 0 net=1407
rlabel metal2 450 -756 450 -756 0 net=1873
rlabel metal2 530 -756 530 -756 0 net=2598
rlabel metal2 653 -756 653 -756 0 net=2689
rlabel metal2 653 -756 653 -756 0 net=2689
rlabel metal2 72 -758 72 -758 0 net=1108
rlabel metal2 198 -758 198 -758 0 net=849
rlabel metal2 205 -758 205 -758 0 net=795
rlabel metal2 247 -758 247 -758 0 net=1188
rlabel metal2 289 -758 289 -758 0 net=1507
rlabel metal2 450 -758 450 -758 0 net=1933
rlabel metal2 541 -758 541 -758 0 net=2247
rlabel metal2 618 -758 618 -758 0 net=2709
rlabel metal2 75 -760 75 -760 0 net=767
rlabel metal2 233 -760 233 -760 0 net=819
rlabel metal2 320 -760 320 -760 0 net=264
rlabel metal2 625 -760 625 -760 0 net=2559
rlabel metal2 625 -760 625 -760 0 net=2559
rlabel metal2 632 -760 632 -760 0 net=2667
rlabel metal2 79 -762 79 -762 0 net=2227
rlabel metal2 331 -762 331 -762 0 net=1333
rlabel metal2 359 -762 359 -762 0 net=1465
rlabel metal2 485 -762 485 -762 0 net=1901
rlabel metal2 534 -762 534 -762 0 net=2159
rlabel metal2 548 -762 548 -762 0 net=2398
rlabel metal2 86 -764 86 -764 0 net=256
rlabel metal2 471 -764 471 -764 0 net=2133
rlabel metal2 551 -764 551 -764 0 net=2682
rlabel metal2 86 -766 86 -766 0 net=1015
rlabel metal2 107 -766 107 -766 0 net=419
rlabel metal2 177 -766 177 -766 0 net=1355
rlabel metal2 303 -766 303 -766 0 net=1301
rlabel metal2 359 -766 359 -766 0 net=2262
rlabel metal2 471 -766 471 -766 0 net=2177
rlabel metal2 555 -766 555 -766 0 net=2493
rlabel metal2 597 -766 597 -766 0 net=2571
rlabel metal2 667 -766 667 -766 0 net=2811
rlabel metal2 89 -768 89 -768 0 net=2860
rlabel metal2 695 -768 695 -768 0 net=2853
rlabel metal2 93 -770 93 -770 0 net=1211
rlabel metal2 324 -770 324 -770 0 net=1437
rlabel metal2 362 -770 362 -770 0 net=2607
rlabel metal2 646 -770 646 -770 0 net=2741
rlabel metal2 23 -772 23 -772 0 net=1721
rlabel metal2 100 -772 100 -772 0 net=653
rlabel metal2 170 -772 170 -772 0 net=933
rlabel metal2 373 -772 373 -772 0 net=1804
rlabel metal2 23 -774 23 -774 0 net=403
rlabel metal2 149 -774 149 -774 0 net=729
rlabel metal2 198 -774 198 -774 0 net=997
rlabel metal2 254 -774 254 -774 0 net=1269
rlabel metal2 404 -774 404 -774 0 net=336
rlabel metal2 646 -774 646 -774 0 net=2727
rlabel metal2 716 -774 716 -774 0 net=2911
rlabel metal2 51 -776 51 -776 0 net=1059
rlabel metal2 191 -776 191 -776 0 net=869
rlabel metal2 453 -776 453 -776 0 net=1
rlabel metal2 548 -776 548 -776 0 net=2943
rlabel metal2 51 -778 51 -778 0 net=455
rlabel metal2 443 -778 443 -778 0 net=817
rlabel metal2 583 -778 583 -778 0 net=2461
rlabel metal2 107 -780 107 -780 0 net=977
rlabel metal2 135 -780 135 -780 0 net=693
rlabel metal2 159 -780 159 -780 0 net=2073
rlabel metal2 37 -782 37 -782 0 net=1389
rlabel metal2 142 -782 142 -782 0 net=471
rlabel metal2 212 -782 212 -782 0 net=1279
rlabel metal2 457 -782 457 -782 0 net=1779
rlabel metal2 37 -784 37 -784 0 net=2416
rlabel metal2 254 -786 254 -786 0 net=2837
rlabel metal2 285 -788 285 -788 0 net=2505
rlabel metal2 478 -790 478 -790 0 net=2873
rlabel metal2 499 -792 499 -792 0 net=2049
rlabel metal2 436 -794 436 -794 0 net=2021
rlabel metal2 429 -796 429 -796 0 net=1691
rlabel metal2 415 -798 415 -798 0 net=1665
rlabel metal2 401 -800 401 -800 0 net=1597
rlabel metal2 68 -802 68 -802 0 net=49
rlabel metal2 23 -813 23 -813 0 net=404
rlabel metal2 170 -813 170 -813 0 net=1060
rlabel metal2 254 -813 254 -813 0 net=1141
rlabel metal2 282 -813 282 -813 0 net=1032
rlabel metal2 310 -813 310 -813 0 net=1467
rlabel metal2 394 -813 394 -813 0 net=1667
rlabel metal2 450 -813 450 -813 0 net=1935
rlabel metal2 450 -813 450 -813 0 net=1935
rlabel metal2 478 -813 478 -813 0 net=2075
rlabel metal2 544 -813 544 -813 0 net=2742
rlabel metal2 737 -813 737 -813 0 net=2933
rlabel metal2 737 -813 737 -813 0 net=2933
rlabel metal2 9 -815 9 -815 0 net=1841
rlabel metal2 30 -815 30 -815 0 net=538
rlabel metal2 65 -815 65 -815 0 net=1572
rlabel metal2 156 -815 156 -815 0 net=821
rlabel metal2 240 -815 240 -815 0 net=850
rlabel metal2 261 -815 261 -815 0 net=934
rlabel metal2 261 -815 261 -815 0 net=934
rlabel metal2 271 -815 271 -815 0 net=818
rlabel metal2 481 -815 481 -815 0 net=2314
rlabel metal2 597 -815 597 -815 0 net=2968
rlabel metal2 9 -817 9 -817 0 net=805
rlabel metal2 177 -817 177 -817 0 net=1357
rlabel metal2 219 -817 219 -817 0 net=797
rlabel metal2 226 -817 226 -817 0 net=570
rlabel metal2 397 -817 397 -817 0 net=1874
rlabel metal2 513 -817 513 -817 0 net=1753
rlabel metal2 548 -817 548 -817 0 net=2728
rlabel metal2 744 -817 744 -817 0 net=2331
rlabel metal2 16 -819 16 -819 0 net=897
rlabel metal2 72 -819 72 -819 0 net=1016
rlabel metal2 93 -819 93 -819 0 net=1723
rlabel metal2 240 -819 240 -819 0 net=1651
rlabel metal2 429 -819 429 -819 0 net=1781
rlabel metal2 485 -819 485 -819 0 net=2239
rlabel metal2 618 -819 618 -819 0 net=3050
rlabel metal2 86 -821 86 -821 0 net=1391
rlabel metal2 117 -821 117 -821 0 net=363
rlabel metal2 184 -821 184 -821 0 net=943
rlabel metal2 275 -821 275 -821 0 net=1281
rlabel metal2 345 -821 345 -821 0 net=2367
rlabel metal2 408 -821 408 -821 0 net=2119
rlabel metal2 513 -821 513 -821 0 net=2297
rlabel metal2 548 -821 548 -821 0 net=2463
rlabel metal2 618 -821 618 -821 0 net=2867
rlabel metal2 75 -823 75 -823 0 net=91
rlabel metal2 121 -823 121 -823 0 net=421
rlabel metal2 135 -823 135 -823 0 net=695
rlabel metal2 184 -823 184 -823 0 net=769
rlabel metal2 219 -823 219 -823 0 net=1303
rlabel metal2 331 -823 331 -823 0 net=1439
rlabel metal2 345 -823 345 -823 0 net=2608
rlabel metal2 646 -823 646 -823 0 net=2913
rlabel metal2 93 -825 93 -825 0 net=979
rlabel metal2 110 -825 110 -825 0 net=870
rlabel metal2 205 -825 205 -825 0 net=1581
rlabel metal2 282 -825 282 -825 0 net=1693
rlabel metal2 443 -825 443 -825 0 net=1981
rlabel metal2 562 -825 562 -825 0 net=2507
rlabel metal2 702 -825 702 -825 0 net=3019
rlabel metal2 72 -827 72 -827 0 net=1729
rlabel metal2 121 -827 121 -827 0 net=731
rlabel metal2 191 -827 191 -827 0 net=1271
rlabel metal2 338 -827 338 -827 0 net=1483
rlabel metal2 404 -827 404 -827 0 net=2489
rlabel metal2 569 -827 569 -827 0 net=2573
rlabel metal2 751 -827 751 -827 0 net=3063
rlabel metal2 79 -829 79 -829 0 net=2228
rlabel metal2 296 -829 296 -829 0 net=1213
rlabel metal2 348 -829 348 -829 0 net=2890
rlabel metal2 758 -829 758 -829 0 net=2055
rlabel metal2 51 -831 51 -831 0 net=457
rlabel metal2 100 -831 100 -831 0 net=655
rlabel metal2 163 -831 163 -831 0 net=1859
rlabel metal2 359 -831 359 -831 0 net=1601
rlabel metal2 411 -831 411 -831 0 net=2050
rlabel metal2 590 -831 590 -831 0 net=2669
rlabel metal2 688 -831 688 -831 0 net=2993
rlabel metal2 30 -833 30 -833 0 net=2693
rlabel metal2 142 -833 142 -833 0 net=473
rlabel metal2 366 -833 366 -833 0 net=2637
rlabel metal2 583 -833 583 -833 0 net=2691
rlabel metal2 44 -835 44 -835 0 net=1409
rlabel metal2 247 -835 247 -835 0 net=210
rlabel metal2 422 -835 422 -835 0 net=1903
rlabel metal2 611 -835 611 -835 0 net=2839
rlabel metal2 44 -837 44 -837 0 net=1951
rlabel metal2 198 -837 198 -837 0 net=999
rlabel metal2 324 -837 324 -837 0 net=1605
rlabel metal2 373 -837 373 -837 0 net=2745
rlabel metal2 632 -837 632 -837 0 net=2711
rlabel metal2 58 -839 58 -839 0 net=787
rlabel metal2 198 -839 198 -839 0 net=1509
rlabel metal2 373 -839 373 -839 0 net=1809
rlabel metal2 492 -839 492 -839 0 net=2713
rlabel metal2 639 -839 639 -839 0 net=2813
rlabel metal2 58 -841 58 -841 0 net=465
rlabel metal2 264 -841 264 -841 0 net=2359
rlabel metal2 653 -841 653 -841 0 net=2855
rlabel metal2 289 -843 289 -843 0 net=1335
rlabel metal2 380 -843 380 -843 0 net=2917
rlabel metal2 667 -843 667 -843 0 net=2937
rlabel metal2 352 -845 352 -845 0 net=1599
rlabel metal2 436 -845 436 -845 0 net=2179
rlabel metal2 695 -845 695 -845 0 net=2945
rlabel metal2 415 -847 415 -847 0 net=2161
rlabel metal2 457 -849 457 -849 0 net=2135
rlabel metal2 471 -851 471 -851 0 net=2023
rlabel metal2 534 -851 534 -851 0 net=2495
rlabel metal2 555 -853 555 -853 0 net=2249
rlabel metal2 576 -855 576 -855 0 net=2561
rlabel metal2 625 -857 625 -857 0 net=2875
rlabel metal2 9 -868 9 -868 0 net=806
rlabel metal2 471 -868 471 -868 0 net=2024
rlabel metal2 544 -868 544 -868 0 net=2692
rlabel metal2 604 -868 604 -868 0 net=13
rlabel metal2 733 -868 733 -868 0 net=2934
rlabel metal2 747 -868 747 -868 0 net=3064
rlabel metal2 19 -870 19 -870 0 net=1842
rlabel metal2 51 -870 51 -870 0 net=981
rlabel metal2 114 -870 114 -870 0 net=509
rlabel metal2 124 -870 124 -870 0 net=2076
rlabel metal2 499 -870 499 -870 0 net=2497
rlabel metal2 583 -870 583 -870 0 net=2747
rlabel metal2 604 -870 604 -870 0 net=2815
rlabel metal2 663 -870 663 -870 0 net=2994
rlabel metal2 726 -870 726 -870 0 net=2056
rlabel metal2 54 -872 54 -872 0 net=104
rlabel metal2 135 -872 135 -872 0 net=696
rlabel metal2 180 -872 180 -872 0 net=1282
rlabel metal2 282 -872 282 -872 0 net=1694
rlabel metal2 387 -872 387 -872 0 net=1905
rlabel metal2 502 -872 502 -872 0 net=2712
rlabel metal2 674 -872 674 -872 0 net=3021
rlabel metal2 30 -874 30 -874 0 net=2695
rlabel metal2 317 -874 317 -874 0 net=1861
rlabel metal2 390 -874 390 -874 0 net=1936
rlabel metal2 520 -874 520 -874 0 net=2639
rlabel metal2 632 -874 632 -874 0 net=2915
rlabel metal2 681 -874 681 -874 0 net=2332
rlabel metal2 58 -876 58 -876 0 net=466
rlabel metal2 212 -876 212 -876 0 net=1358
rlabel metal2 317 -876 317 -876 0 net=1485
rlabel metal2 345 -876 345 -876 0 net=1735
rlabel metal2 642 -876 642 -876 0 net=463
rlabel metal2 681 -876 681 -876 0 net=2947
rlabel metal2 58 -878 58 -878 0 net=1393
rlabel metal2 93 -878 93 -878 0 net=2153
rlabel metal2 121 -878 121 -878 0 net=733
rlabel metal2 142 -878 142 -878 0 net=789
rlabel metal2 149 -878 149 -878 0 net=656
rlabel metal2 257 -878 257 -878 0 net=798
rlabel metal2 352 -878 352 -878 0 net=1600
rlabel metal2 401 -878 401 -878 0 net=2369
rlabel metal2 450 -878 450 -878 0 net=1755
rlabel metal2 534 -878 534 -878 0 net=2563
rlabel metal2 684 -878 684 -878 0 net=1447
rlabel metal2 65 -880 65 -880 0 net=898
rlabel metal2 352 -880 352 -880 0 net=1669
rlabel metal2 401 -880 401 -880 0 net=1983
rlabel metal2 527 -880 527 -880 0 net=2575
rlabel metal2 576 -880 576 -880 0 net=2869
rlabel metal2 65 -882 65 -882 0 net=1305
rlabel metal2 261 -882 261 -882 0 net=1811
rlabel metal2 394 -882 394 -882 0 net=2856
rlabel metal2 79 -884 79 -884 0 net=459
rlabel metal2 163 -884 163 -884 0 net=475
rlabel metal2 163 -884 163 -884 0 net=475
rlabel metal2 170 -884 170 -884 0 net=1469
rlabel metal2 366 -884 366 -884 0 net=2255
rlabel metal2 492 -884 492 -884 0 net=2715
rlabel metal2 618 -884 618 -884 0 net=2939
rlabel metal2 79 -886 79 -886 0 net=1653
rlabel metal2 271 -886 271 -886 0 net=1214
rlabel metal2 303 -886 303 -886 0 net=1441
rlabel metal2 373 -886 373 -886 0 net=2407
rlabel metal2 541 -886 541 -886 0 net=2509
rlabel metal2 86 -888 86 -888 0 net=1071
rlabel metal2 142 -888 142 -888 0 net=1273
rlabel metal2 198 -888 198 -888 0 net=1511
rlabel metal2 271 -888 271 -888 0 net=33
rlabel metal2 464 -888 464 -888 0 net=2361
rlabel metal2 555 -888 555 -888 0 net=2251
rlabel metal2 100 -890 100 -890 0 net=1411
rlabel metal2 219 -890 219 -890 0 net=1143
rlabel metal2 275 -890 275 -890 0 net=1607
rlabel metal2 331 -890 331 -890 0 net=2181
rlabel metal2 562 -890 562 -890 0 net=2671
rlabel metal2 72 -892 72 -892 0 net=1731
rlabel metal2 107 -892 107 -892 0 net=423
rlabel metal2 198 -892 198 -892 0 net=944
rlabel metal2 289 -892 289 -892 0 net=1337
rlabel metal2 415 -892 415 -892 0 net=2163
rlabel metal2 590 -892 590 -892 0 net=2841
rlabel metal2 72 -894 72 -894 0 net=1724
rlabel metal2 289 -894 289 -894 0 net=2121
rlabel metal2 415 -894 415 -894 0 net=2115
rlabel metal2 611 -894 611 -894 0 net=2877
rlabel metal2 40 -896 40 -896 0 net=1815
rlabel metal2 310 -896 310 -896 0 net=1603
rlabel metal2 408 -896 408 -896 0 net=1783
rlabel metal2 625 -896 625 -896 0 net=2919
rlabel metal2 128 -898 128 -898 0 net=823
rlabel metal2 173 -898 173 -898 0 net=2759
rlabel metal2 156 -900 156 -900 0 net=2025
rlabel metal2 429 -900 429 -900 0 net=2137
rlabel metal2 506 -900 506 -900 0 net=2490
rlabel metal2 184 -902 184 -902 0 net=771
rlabel metal2 457 -902 457 -902 0 net=2241
rlabel metal2 506 -902 506 -902 0 net=2465
rlabel metal2 184 -904 184 -904 0 net=1001
rlabel metal2 296 -904 296 -904 0 net=2579
rlabel metal2 44 -906 44 -906 0 net=1953
rlabel metal2 485 -906 485 -906 0 net=2299
rlabel metal2 44 -908 44 -908 0 net=1583
rlabel metal2 208 -908 208 -908 0 net=2511
rlabel metal2 205 -910 205 -910 0 net=2355
rlabel metal2 44 -921 44 -921 0 net=1584
rlabel metal2 464 -921 464 -921 0 net=2362
rlabel metal2 520 -921 520 -921 0 net=2870
rlabel metal2 646 -921 646 -921 0 net=464
rlabel metal2 660 -921 660 -921 0 net=3023
rlabel metal2 716 -921 716 -921 0 net=1448
rlabel metal2 51 -923 51 -923 0 net=982
rlabel metal2 135 -923 135 -923 0 net=735
rlabel metal2 135 -923 135 -923 0 net=735
rlabel metal2 163 -923 163 -923 0 net=477
rlabel metal2 163 -923 163 -923 0 net=477
rlabel metal2 170 -923 170 -923 0 net=1471
rlabel metal2 191 -923 191 -923 0 net=790
rlabel metal2 219 -923 219 -923 0 net=1144
rlabel metal2 282 -923 282 -923 0 net=2696
rlabel metal2 320 -923 320 -923 0 net=2370
rlabel metal2 464 -923 464 -923 0 net=2761
rlabel metal2 674 -923 674 -923 0 net=2949
rlabel metal2 72 -925 72 -925 0 net=2155
rlabel metal2 103 -925 103 -925 0 net=1741
rlabel metal2 142 -925 142 -925 0 net=1275
rlabel metal2 226 -925 226 -925 0 net=1816
rlabel metal2 492 -925 492 -925 0 net=2717
rlabel metal2 107 -927 107 -927 0 net=424
rlabel metal2 159 -927 159 -927 0 net=657
rlabel metal2 184 -927 184 -927 0 net=1003
rlabel metal2 240 -927 240 -927 0 net=1512
rlabel metal2 394 -927 394 -927 0 net=2139
rlabel metal2 499 -927 499 -927 0 net=2499
rlabel metal2 86 -929 86 -929 0 net=1072
rlabel metal2 128 -929 128 -929 0 net=825
rlabel metal2 184 -929 184 -929 0 net=773
rlabel metal2 240 -929 240 -929 0 net=1671
rlabel metal2 499 -929 499 -929 0 net=2941
rlabel metal2 58 -931 58 -931 0 net=1395
rlabel metal2 100 -931 100 -931 0 net=1733
rlabel metal2 191 -931 191 -931 0 net=777
rlabel metal2 527 -931 527 -931 0 net=2577
rlabel metal2 618 -931 618 -931 0 net=405
rlabel metal2 114 -933 114 -933 0 net=511
rlabel metal2 254 -933 254 -933 0 net=1077
rlabel metal2 450 -933 450 -933 0 net=1757
rlabel metal2 541 -933 541 -933 0 net=2510
rlabel metal2 198 -935 198 -935 0 net=170
rlabel metal2 555 -935 555 -935 0 net=2879
rlabel metal2 149 -937 149 -937 0 net=460
rlabel metal2 254 -937 254 -937 0 net=2165
rlabel metal2 534 -937 534 -937 0 net=2565
rlabel metal2 149 -939 149 -939 0 net=1541
rlabel metal2 268 -939 268 -939 0 net=1487
rlabel metal2 324 -939 324 -939 0 net=2357
rlabel metal2 156 -941 156 -941 0 net=633
rlabel metal2 352 -941 352 -941 0 net=2117
rlabel metal2 436 -941 436 -941 0 net=2243
rlabel metal2 471 -941 471 -941 0 net=2301
rlabel metal2 275 -943 275 -943 0 net=1609
rlabel metal2 289 -943 289 -943 0 net=2122
rlabel metal2 310 -943 310 -943 0 net=1604
rlabel metal2 79 -945 79 -945 0 net=1655
rlabel metal2 296 -945 296 -945 0 net=1339
rlabel metal2 366 -945 366 -945 0 net=2916
rlabel metal2 79 -947 79 -947 0 net=1443
rlabel metal2 338 -947 338 -947 0 net=2027
rlabel metal2 408 -947 408 -947 0 net=1785
rlabel metal2 275 -949 275 -949 0 net=1737
rlabel metal2 359 -949 359 -949 0 net=1863
rlabel metal2 408 -949 408 -949 0 net=2257
rlabel metal2 457 -949 457 -949 0 net=2749
rlabel metal2 247 -951 247 -951 0 net=1955
rlabel metal2 380 -951 380 -951 0 net=1907
rlabel metal2 443 -951 443 -951 0 net=2513
rlabel metal2 583 -951 583 -951 0 net=2641
rlabel metal2 212 -953 212 -953 0 net=1413
rlabel metal2 303 -953 303 -953 0 net=2683
rlabel metal2 478 -953 478 -953 0 net=2409
rlabel metal2 513 -953 513 -953 0 net=2673
rlabel metal2 65 -955 65 -955 0 net=1307
rlabel metal2 331 -955 331 -955 0 net=2183
rlabel metal2 65 -957 65 -957 0 net=2871
rlabel metal2 261 -957 261 -957 0 net=1813
rlabel metal2 478 -957 478 -957 0 net=2581
rlabel metal2 261 -959 261 -959 0 net=1985
rlabel metal2 506 -959 506 -959 0 net=2467
rlabel metal2 373 -961 373 -961 0 net=2787
rlabel metal2 506 -961 506 -961 0 net=2127
rlabel metal2 548 -963 548 -963 0 net=2843
rlabel metal2 590 -965 590 -965 0 net=2921
rlabel metal2 604 -967 604 -967 0 net=2816
rlabel metal2 604 -969 604 -969 0 net=2253
rlabel metal2 65 -980 65 -980 0 net=2872
rlabel metal2 254 -980 254 -980 0 net=2166
rlabel metal2 422 -980 422 -980 0 net=2718
rlabel metal2 523 -980 523 -980 0 net=1758
rlabel metal2 544 -980 544 -980 0 net=2578
rlabel metal2 576 -980 576 -980 0 net=2501
rlabel metal2 607 -980 607 -980 0 net=2566
rlabel metal2 649 -980 649 -980 0 net=3024
rlabel metal2 670 -980 670 -980 0 net=2950
rlabel metal2 72 -982 72 -982 0 net=2156
rlabel metal2 100 -982 100 -982 0 net=56
rlabel metal2 254 -982 254 -982 0 net=1493
rlabel metal2 373 -982 373 -982 0 net=2514
rlabel metal2 453 -982 453 -982 0 net=2942
rlabel metal2 527 -982 527 -982 0 net=1786
rlabel metal2 548 -982 548 -982 0 net=2845
rlabel metal2 548 -982 548 -982 0 net=2845
rlabel metal2 555 -982 555 -982 0 net=2881
rlabel metal2 576 -982 576 -982 0 net=2923
rlabel metal2 611 -982 611 -982 0 net=407
rlabel metal2 79 -984 79 -984 0 net=1445
rlabel metal2 212 -984 212 -984 0 net=1308
rlabel metal2 380 -984 380 -984 0 net=1908
rlabel metal2 464 -984 464 -984 0 net=2763
rlabel metal2 464 -984 464 -984 0 net=2763
rlabel metal2 471 -984 471 -984 0 net=2303
rlabel metal2 93 -986 93 -986 0 net=2473
rlabel metal2 107 -986 107 -986 0 net=1734
rlabel metal2 149 -986 149 -986 0 net=1543
rlabel metal2 149 -986 149 -986 0 net=1543
rlabel metal2 170 -986 170 -986 0 net=658
rlabel metal2 264 -986 264 -986 0 net=2358
rlabel metal2 331 -986 331 -986 0 net=1814
rlabel metal2 331 -986 331 -986 0 net=1814
rlabel metal2 352 -986 352 -986 0 net=2118
rlabel metal2 394 -986 394 -986 0 net=2141
rlabel metal2 425 -986 425 -986 0 net=2244
rlabel metal2 439 -986 439 -986 0 net=2128
rlabel metal2 86 -988 86 -988 0 net=1397
rlabel metal2 191 -988 191 -988 0 net=778
rlabel metal2 240 -988 240 -988 0 net=1673
rlabel metal2 369 -988 369 -988 0 net=2184
rlabel metal2 117 -990 117 -990 0 net=1742
rlabel metal2 177 -990 177 -990 0 net=1473
rlabel metal2 268 -990 268 -990 0 net=1489
rlabel metal2 380 -990 380 -990 0 net=411
rlabel metal2 492 -990 492 -990 0 net=2675
rlabel metal2 163 -992 163 -992 0 net=479
rlabel metal2 184 -992 184 -992 0 net=775
rlabel metal2 296 -992 296 -992 0 net=1341
rlabel metal2 401 -992 401 -992 0 net=2789
rlabel metal2 401 -992 401 -992 0 net=2789
rlabel metal2 429 -992 429 -992 0 net=1078
rlabel metal2 156 -994 156 -994 0 net=635
rlabel metal2 184 -994 184 -994 0 net=1005
rlabel metal2 226 -994 226 -994 0 net=1657
rlabel metal2 303 -994 303 -994 0 net=2684
rlabel metal2 450 -994 450 -994 0 net=2583
rlabel metal2 506 -994 506 -994 0 net=2643
rlabel metal2 142 -996 142 -996 0 net=827
rlabel metal2 191 -996 191 -996 0 net=1611
rlabel metal2 310 -996 310 -996 0 net=1957
rlabel metal2 429 -996 429 -996 0 net=2410
rlabel metal2 562 -996 562 -996 0 net=2469
rlabel metal2 135 -998 135 -998 0 net=737
rlabel metal2 205 -998 205 -998 0 net=1739
rlabel metal2 282 -998 282 -998 0 net=1713
rlabel metal2 233 -1000 233 -1000 0 net=513
rlabel metal2 317 -1000 317 -1000 0 net=2750
rlabel metal2 219 -1002 219 -1002 0 net=1277
rlabel metal2 261 -1002 261 -1002 0 net=1987
rlabel metal2 324 -1002 324 -1002 0 net=2029
rlabel metal2 345 -1002 345 -1002 0 net=2258
rlabel metal2 457 -1002 457 -1002 0 net=2254
rlabel metal2 219 -1004 219 -1004 0 net=1415
rlabel metal2 338 -1004 338 -1004 0 net=1865
rlabel metal2 408 -1004 408 -1004 0 net=2817
rlabel metal2 247 -1006 247 -1006 0 net=2781
rlabel metal2 313 -1006 313 -1006 0 net=2085
rlabel metal2 359 -1008 359 -1008 0 net=3027
rlabel metal2 100 -1019 100 -1019 0 net=2475
rlabel metal2 100 -1019 100 -1019 0 net=2475
rlabel metal2 114 -1019 114 -1019 0 net=857
rlabel metal2 198 -1019 198 -1019 0 net=1446
rlabel metal2 352 -1019 352 -1019 0 net=1674
rlabel metal2 478 -1019 478 -1019 0 net=2645
rlabel metal2 548 -1019 548 -1019 0 net=2847
rlabel metal2 548 -1019 548 -1019 0 net=2847
rlabel metal2 562 -1019 562 -1019 0 net=2925
rlabel metal2 583 -1019 583 -1019 0 net=2471
rlabel metal2 583 -1019 583 -1019 0 net=2471
rlabel metal2 590 -1019 590 -1019 0 net=2503
rlabel metal2 590 -1019 590 -1019 0 net=2503
rlabel metal2 604 -1019 604 -1019 0 net=408
rlabel metal2 128 -1021 128 -1021 0 net=637
rlabel metal2 198 -1021 198 -1021 0 net=1417
rlabel metal2 229 -1021 229 -1021 0 net=151
rlabel metal2 268 -1021 268 -1021 0 net=776
rlabel metal2 373 -1021 373 -1021 0 net=1491
rlabel metal2 436 -1021 436 -1021 0 net=2585
rlabel metal2 457 -1021 457 -1021 0 net=2765
rlabel metal2 485 -1021 485 -1021 0 net=2677
rlabel metal2 499 -1021 499 -1021 0 net=2304
rlabel metal2 569 -1021 569 -1021 0 net=2883
rlabel metal2 569 -1021 569 -1021 0 net=2883
rlabel metal2 135 -1023 135 -1023 0 net=1545
rlabel metal2 163 -1023 163 -1023 0 net=481
rlabel metal2 191 -1023 191 -1023 0 net=1613
rlabel metal2 275 -1023 275 -1023 0 net=514
rlabel metal2 366 -1023 366 -1023 0 net=413
rlabel metal2 387 -1023 387 -1023 0 net=3029
rlabel metal2 387 -1023 387 -1023 0 net=3029
rlabel metal2 394 -1023 394 -1023 0 net=1342
rlabel metal2 149 -1025 149 -1025 0 net=829
rlabel metal2 177 -1025 177 -1025 0 net=1459
rlabel metal2 226 -1025 226 -1025 0 net=1659
rlabel metal2 289 -1025 289 -1025 0 net=1988
rlabel metal2 373 -1025 373 -1025 0 net=2086
rlabel metal2 418 -1025 418 -1025 0 net=2142
rlabel metal2 142 -1027 142 -1027 0 net=739
rlabel metal2 184 -1027 184 -1027 0 net=1007
rlabel metal2 205 -1027 205 -1027 0 net=1740
rlabel metal2 317 -1027 317 -1027 0 net=1867
rlabel metal2 394 -1027 394 -1027 0 net=2791
rlabel metal2 408 -1027 408 -1027 0 net=2819
rlabel metal2 408 -1027 408 -1027 0 net=2819
rlabel metal2 422 -1027 422 -1027 0 net=567
rlabel metal2 124 -1029 124 -1029 0 net=2095
rlabel metal2 170 -1029 170 -1029 0 net=1399
rlabel metal2 215 -1029 215 -1029 0 net=1278
rlabel metal2 240 -1029 240 -1029 0 net=1474
rlabel metal2 254 -1029 254 -1029 0 net=1495
rlabel metal2 296 -1029 296 -1029 0 net=1959
rlabel metal2 439 -1029 439 -1029 0 net=2069
rlabel metal2 170 -1031 170 -1031 0 net=1714
rlabel metal2 299 -1031 299 -1031 0 net=2782
rlabel metal2 310 -1031 310 -1031 0 net=2031
rlabel metal2 215 -1033 215 -1033 0 net=1251
rlabel metal2 233 -1035 233 -1035 0 net=2371
rlabel metal2 261 -1037 261 -1037 0 net=306
rlabel metal2 100 -1048 100 -1048 0 net=2477
rlabel metal2 128 -1048 128 -1048 0 net=638
rlabel metal2 198 -1048 198 -1048 0 net=1418
rlabel metal2 219 -1048 219 -1048 0 net=1461
rlabel metal2 247 -1048 247 -1048 0 net=1614
rlabel metal2 366 -1048 366 -1048 0 net=415
rlabel metal2 383 -1048 383 -1048 0 net=3030
rlabel metal2 394 -1048 394 -1048 0 net=2792
rlabel metal2 408 -1048 408 -1048 0 net=2820
rlabel metal2 415 -1048 415 -1048 0 net=1492
rlabel metal2 443 -1048 443 -1048 0 net=2070
rlabel metal2 457 -1048 457 -1048 0 net=2767
rlabel metal2 457 -1048 457 -1048 0 net=2767
rlabel metal2 471 -1048 471 -1048 0 net=2678
rlabel metal2 541 -1048 541 -1048 0 net=2848
rlabel metal2 562 -1048 562 -1048 0 net=2926
rlabel metal2 562 -1048 562 -1048 0 net=2926
rlabel metal2 579 -1048 579 -1048 0 net=2472
rlabel metal2 142 -1050 142 -1050 0 net=2096
rlabel metal2 180 -1050 180 -1050 0 net=2372
rlabel metal2 254 -1050 254 -1050 0 net=1252
rlabel metal2 278 -1050 278 -1050 0 net=1960
rlabel metal2 299 -1050 299 -1050 0 net=2032
rlabel metal2 376 -1050 376 -1050 0 net=568
rlabel metal2 429 -1050 429 -1050 0 net=2587
rlabel metal2 443 -1050 443 -1050 0 net=2646
rlabel metal2 569 -1050 569 -1050 0 net=2885
rlabel metal2 142 -1052 142 -1052 0 net=740
rlabel metal2 163 -1052 163 -1052 0 net=482
rlabel metal2 191 -1052 191 -1052 0 net=1009
rlabel metal2 205 -1052 205 -1052 0 net=1401
rlabel metal2 268 -1052 268 -1052 0 net=1660
rlabel metal2 285 -1052 285 -1052 0 net=1868
rlabel metal2 579 -1052 579 -1052 0 net=2504
rlabel metal2 149 -1054 149 -1054 0 net=831
rlabel metal2 289 -1054 289 -1054 0 net=1496
rlabel metal2 135 -1056 135 -1056 0 net=1547
rlabel metal2 114 -1058 114 -1058 0 net=858
rlabel metal2 100 -1069 100 -1069 0 net=2478
rlabel metal2 149 -1069 149 -1069 0 net=1548
rlabel metal2 163 -1069 163 -1069 0 net=832
rlabel metal2 198 -1069 198 -1069 0 net=1010
rlabel metal2 215 -1069 215 -1069 0 net=1402
rlabel metal2 380 -1069 380 -1069 0 net=416
rlabel metal2 429 -1069 429 -1069 0 net=2588
rlabel metal2 446 -1069 446 -1069 0 net=2768
rlabel metal2 576 -1069 576 -1069 0 net=2886
rlabel metal2 219 -1071 219 -1071 0 net=1462
<< end >>
