magic
tech scmos
timestamp 1555071777 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 36 -10 42 -4
rect 43 -10 49 -4
rect 99 -10 105 -4
rect 106 -10 112 -4
rect 127 -10 133 -4
rect 134 -10 137 -4
rect 141 -10 147 -4
rect 148 -10 154 -4
rect 155 -10 158 -4
rect 162 -10 168 -4
rect 169 -10 175 -4
rect 176 -10 179 -4
rect 183 -10 189 -4
rect 190 -10 196 -4
rect 197 -10 200 -4
rect 204 -10 210 -4
rect 211 -10 214 -4
rect 1 -29 7 -23
rect 8 -29 14 -23
rect 15 -29 21 -23
rect 22 -29 28 -23
rect 29 -29 35 -23
rect 36 -29 42 -23
rect 78 -29 81 -23
rect 85 -29 91 -23
rect 92 -29 98 -23
rect 99 -29 105 -23
rect 106 -29 112 -23
rect 120 -29 123 -23
rect 127 -29 133 -23
rect 134 -29 137 -23
rect 141 -29 144 -23
rect 148 -29 154 -23
rect 155 -29 161 -23
rect 162 -29 168 -23
rect 169 -29 172 -23
rect 176 -29 182 -23
rect 183 -29 189 -23
rect 190 -29 196 -23
rect 197 -29 200 -23
rect 204 -29 210 -23
rect 211 -29 217 -23
rect 218 -29 221 -23
rect 225 -29 231 -23
rect 232 -29 235 -23
rect 1 -52 7 -46
rect 8 -52 14 -46
rect 15 -52 21 -46
rect 22 -52 28 -46
rect 29 -52 35 -46
rect 57 -52 63 -46
rect 64 -52 67 -46
rect 71 -52 74 -46
rect 78 -52 84 -46
rect 85 -52 91 -46
rect 92 -52 98 -46
rect 99 -52 102 -46
rect 106 -52 112 -46
rect 113 -52 116 -46
rect 120 -52 126 -46
rect 127 -52 133 -46
rect 134 -52 137 -46
rect 141 -52 147 -46
rect 148 -52 154 -46
rect 155 -52 158 -46
rect 162 -52 165 -46
rect 169 -52 175 -46
rect 176 -52 182 -46
rect 183 -52 186 -46
rect 190 -52 193 -46
rect 197 -52 203 -46
rect 204 -52 207 -46
rect 211 -52 217 -46
rect 218 -52 224 -46
rect 225 -52 228 -46
rect 232 -52 235 -46
rect 239 -52 242 -46
rect 246 -52 249 -46
rect 253 -52 256 -46
rect 260 -52 263 -46
rect 267 -52 273 -46
rect 274 -52 277 -46
rect 281 -52 284 -46
rect 1 -83 7 -77
rect 8 -83 14 -77
rect 15 -83 21 -77
rect 22 -83 28 -77
rect 29 -83 32 -77
rect 36 -83 42 -77
rect 43 -83 46 -77
rect 50 -83 53 -77
rect 57 -83 60 -77
rect 64 -83 67 -77
rect 71 -83 77 -77
rect 78 -83 81 -77
rect 85 -83 88 -77
rect 92 -83 95 -77
rect 99 -83 105 -77
rect 106 -83 112 -77
rect 113 -83 119 -77
rect 120 -83 123 -77
rect 127 -83 133 -77
rect 134 -83 140 -77
rect 141 -83 144 -77
rect 148 -83 151 -77
rect 155 -83 161 -77
rect 162 -83 165 -77
rect 169 -83 172 -77
rect 176 -83 182 -77
rect 183 -83 189 -77
rect 190 -83 193 -77
rect 197 -83 203 -77
rect 204 -83 210 -77
rect 211 -83 217 -77
rect 218 -83 221 -77
rect 225 -83 228 -77
rect 232 -83 235 -77
rect 239 -83 245 -77
rect 246 -83 252 -77
rect 253 -83 256 -77
rect 260 -83 263 -77
rect 267 -83 270 -77
rect 274 -83 277 -77
rect 281 -83 284 -77
rect 288 -83 291 -77
rect 295 -83 301 -77
rect 302 -83 305 -77
rect 1 -128 7 -122
rect 8 -128 14 -122
rect 15 -128 18 -122
rect 22 -128 28 -122
rect 29 -128 32 -122
rect 36 -128 39 -122
rect 43 -128 49 -122
rect 50 -128 53 -122
rect 57 -128 63 -122
rect 64 -128 70 -122
rect 71 -128 74 -122
rect 78 -128 84 -122
rect 85 -128 88 -122
rect 92 -128 95 -122
rect 99 -128 105 -122
rect 106 -128 109 -122
rect 113 -128 119 -122
rect 120 -128 126 -122
rect 127 -128 133 -122
rect 134 -128 140 -122
rect 141 -128 147 -122
rect 148 -128 154 -122
rect 155 -128 161 -122
rect 162 -128 168 -122
rect 169 -128 172 -122
rect 176 -128 182 -122
rect 183 -128 189 -122
rect 190 -128 196 -122
rect 197 -128 203 -122
rect 204 -128 210 -122
rect 211 -128 214 -122
rect 218 -128 221 -122
rect 225 -128 228 -122
rect 232 -128 238 -122
rect 239 -128 242 -122
rect 246 -128 249 -122
rect 253 -128 256 -122
rect 260 -128 263 -122
rect 267 -128 270 -122
rect 274 -128 277 -122
rect 281 -128 284 -122
rect 288 -128 291 -122
rect 295 -128 298 -122
rect 302 -128 305 -122
rect 309 -128 312 -122
rect 316 -128 319 -122
rect 323 -128 326 -122
rect 330 -128 333 -122
rect 1 -175 7 -169
rect 8 -175 14 -169
rect 15 -175 21 -169
rect 22 -175 28 -169
rect 29 -175 32 -169
rect 36 -175 42 -169
rect 43 -175 46 -169
rect 50 -175 56 -169
rect 57 -175 63 -169
rect 64 -175 67 -169
rect 71 -175 74 -169
rect 78 -175 81 -169
rect 85 -175 91 -169
rect 92 -175 95 -169
rect 99 -175 102 -169
rect 106 -175 112 -169
rect 113 -175 119 -169
rect 120 -175 126 -169
rect 127 -175 130 -169
rect 134 -175 140 -169
rect 141 -175 144 -169
rect 148 -175 154 -169
rect 155 -175 161 -169
rect 162 -175 168 -169
rect 169 -175 172 -169
rect 176 -175 179 -169
rect 183 -175 186 -169
rect 190 -175 196 -169
rect 197 -175 203 -169
rect 204 -175 210 -169
rect 211 -175 217 -169
rect 218 -175 221 -169
rect 225 -175 228 -169
rect 232 -175 238 -169
rect 239 -175 245 -169
rect 246 -175 249 -169
rect 253 -175 256 -169
rect 260 -175 263 -169
rect 267 -175 273 -169
rect 274 -175 277 -169
rect 281 -175 284 -169
rect 288 -175 291 -169
rect 295 -175 298 -169
rect 302 -175 305 -169
rect 309 -175 312 -169
rect 1 -212 7 -206
rect 8 -212 11 -206
rect 15 -212 18 -206
rect 22 -212 28 -206
rect 29 -212 35 -206
rect 36 -212 39 -206
rect 43 -212 46 -206
rect 50 -212 56 -206
rect 57 -212 60 -206
rect 64 -212 70 -206
rect 71 -212 77 -206
rect 78 -212 81 -206
rect 85 -212 91 -206
rect 92 -212 95 -206
rect 99 -212 102 -206
rect 106 -212 112 -206
rect 113 -212 119 -206
rect 120 -212 123 -206
rect 127 -212 130 -206
rect 134 -212 137 -206
rect 141 -212 147 -206
rect 148 -212 154 -206
rect 155 -212 161 -206
rect 162 -212 165 -206
rect 169 -212 172 -206
rect 176 -212 179 -206
rect 183 -212 189 -206
rect 190 -212 193 -206
rect 197 -212 200 -206
rect 204 -212 210 -206
rect 211 -212 217 -206
rect 218 -212 224 -206
rect 225 -212 228 -206
rect 232 -212 238 -206
rect 239 -212 242 -206
rect 246 -212 249 -206
rect 253 -212 256 -206
rect 260 -212 263 -206
rect 267 -212 273 -206
rect 274 -212 277 -206
rect 281 -212 287 -206
rect 288 -212 294 -206
rect 295 -212 298 -206
rect 302 -212 305 -206
rect 309 -212 312 -206
rect 316 -212 319 -206
rect 323 -212 326 -206
rect 330 -212 333 -206
rect 337 -212 340 -206
rect 344 -212 347 -206
rect 351 -212 354 -206
rect 358 -212 361 -206
rect 365 -212 368 -206
rect 372 -212 375 -206
rect 379 -212 382 -206
rect 386 -212 392 -206
rect 393 -212 396 -206
rect 8 -257 11 -251
rect 15 -257 18 -251
rect 22 -257 28 -251
rect 29 -257 32 -251
rect 36 -257 39 -251
rect 43 -257 46 -251
rect 50 -257 53 -251
rect 57 -257 60 -251
rect 64 -257 70 -251
rect 71 -257 77 -251
rect 78 -257 84 -251
rect 85 -257 88 -251
rect 92 -257 95 -251
rect 99 -257 105 -251
rect 106 -257 112 -251
rect 113 -257 116 -251
rect 120 -257 126 -251
rect 127 -257 130 -251
rect 134 -257 140 -251
rect 141 -257 144 -251
rect 148 -257 154 -251
rect 155 -257 161 -251
rect 162 -257 165 -251
rect 169 -257 172 -251
rect 176 -257 179 -251
rect 183 -257 186 -251
rect 190 -257 193 -251
rect 197 -257 203 -251
rect 204 -257 210 -251
rect 211 -257 217 -251
rect 218 -257 221 -251
rect 225 -257 231 -251
rect 232 -257 235 -251
rect 239 -257 242 -251
rect 246 -257 249 -251
rect 253 -257 256 -251
rect 260 -257 266 -251
rect 267 -257 270 -251
rect 274 -257 280 -251
rect 281 -257 284 -251
rect 288 -257 294 -251
rect 295 -257 298 -251
rect 302 -257 305 -251
rect 309 -257 312 -251
rect 316 -257 319 -251
rect 323 -257 326 -251
rect 330 -257 333 -251
rect 337 -257 340 -251
rect 344 -257 347 -251
rect 351 -257 354 -251
rect 358 -257 361 -251
rect 365 -257 371 -251
rect 372 -257 378 -251
rect 379 -257 382 -251
rect 1 -304 4 -298
rect 8 -304 11 -298
rect 15 -304 18 -298
rect 22 -304 25 -298
rect 29 -304 32 -298
rect 36 -304 39 -298
rect 43 -304 46 -298
rect 50 -304 56 -298
rect 57 -304 63 -298
rect 64 -304 67 -298
rect 71 -304 74 -298
rect 78 -304 84 -298
rect 85 -304 88 -298
rect 92 -304 95 -298
rect 99 -304 102 -298
rect 106 -304 109 -298
rect 113 -304 116 -298
rect 120 -304 126 -298
rect 127 -304 130 -298
rect 134 -304 140 -298
rect 141 -304 144 -298
rect 148 -304 151 -298
rect 155 -304 161 -298
rect 162 -304 168 -298
rect 169 -304 172 -298
rect 176 -304 179 -298
rect 183 -304 189 -298
rect 190 -304 193 -298
rect 197 -304 203 -298
rect 204 -304 210 -298
rect 211 -304 217 -298
rect 218 -304 221 -298
rect 225 -304 228 -298
rect 232 -304 238 -298
rect 239 -304 245 -298
rect 246 -304 252 -298
rect 253 -304 259 -298
rect 260 -304 263 -298
rect 267 -304 270 -298
rect 274 -304 277 -298
rect 281 -304 284 -298
rect 288 -304 291 -298
rect 295 -304 301 -298
rect 302 -304 305 -298
rect 309 -304 312 -298
rect 316 -304 319 -298
rect 323 -304 326 -298
rect 330 -304 333 -298
rect 337 -304 340 -298
rect 344 -304 347 -298
rect 351 -304 354 -298
rect 358 -304 361 -298
rect 365 -304 371 -298
rect 372 -304 378 -298
rect 379 -304 382 -298
rect 1 -345 4 -339
rect 8 -345 11 -339
rect 15 -345 18 -339
rect 22 -345 25 -339
rect 29 -345 32 -339
rect 36 -345 39 -339
rect 43 -345 49 -339
rect 50 -345 53 -339
rect 57 -345 63 -339
rect 64 -345 70 -339
rect 71 -345 74 -339
rect 78 -345 81 -339
rect 85 -345 91 -339
rect 92 -345 95 -339
rect 99 -345 105 -339
rect 106 -345 112 -339
rect 113 -345 119 -339
rect 120 -345 126 -339
rect 127 -345 130 -339
rect 134 -345 137 -339
rect 141 -345 147 -339
rect 148 -345 154 -339
rect 155 -345 161 -339
rect 162 -345 165 -339
rect 169 -345 175 -339
rect 176 -345 179 -339
rect 183 -345 186 -339
rect 190 -345 196 -339
rect 197 -345 200 -339
rect 204 -345 210 -339
rect 211 -345 217 -339
rect 218 -345 221 -339
rect 225 -345 228 -339
rect 232 -345 238 -339
rect 239 -345 245 -339
rect 246 -345 249 -339
rect 253 -345 256 -339
rect 260 -345 263 -339
rect 267 -345 270 -339
rect 274 -345 277 -339
rect 281 -345 284 -339
rect 288 -345 291 -339
rect 295 -345 298 -339
rect 302 -345 305 -339
rect 309 -345 312 -339
rect 316 -345 319 -339
rect 323 -345 326 -339
rect 330 -345 333 -339
rect 337 -345 343 -339
rect 344 -345 347 -339
rect 351 -345 354 -339
rect 358 -345 361 -339
rect 372 -345 378 -339
rect 386 -345 389 -339
rect 8 -390 11 -384
rect 15 -390 18 -384
rect 22 -390 25 -384
rect 29 -390 32 -384
rect 36 -390 39 -384
rect 43 -390 46 -384
rect 50 -390 53 -384
rect 57 -390 60 -384
rect 64 -390 70 -384
rect 71 -390 74 -384
rect 78 -390 84 -384
rect 85 -390 91 -384
rect 92 -390 98 -384
rect 99 -390 102 -384
rect 106 -390 109 -384
rect 113 -390 119 -384
rect 120 -390 123 -384
rect 127 -390 133 -384
rect 134 -390 137 -384
rect 141 -390 147 -384
rect 148 -390 154 -384
rect 155 -390 161 -384
rect 162 -390 165 -384
rect 169 -390 175 -384
rect 176 -390 179 -384
rect 183 -390 189 -384
rect 190 -390 196 -384
rect 197 -390 200 -384
rect 204 -390 207 -384
rect 211 -390 217 -384
rect 218 -390 224 -384
rect 225 -390 228 -384
rect 232 -390 235 -384
rect 239 -390 245 -384
rect 246 -390 249 -384
rect 253 -390 259 -384
rect 260 -390 263 -384
rect 267 -390 273 -384
rect 274 -390 277 -384
rect 281 -390 287 -384
rect 288 -390 291 -384
rect 295 -390 298 -384
rect 302 -390 305 -384
rect 309 -390 312 -384
rect 316 -390 319 -384
rect 323 -390 326 -384
rect 330 -390 333 -384
rect 337 -390 340 -384
rect 344 -390 347 -384
rect 351 -390 354 -384
rect 358 -390 361 -384
rect 365 -390 368 -384
rect 372 -390 375 -384
rect 379 -390 382 -384
rect 386 -390 389 -384
rect 393 -390 399 -384
rect 400 -390 403 -384
rect 407 -390 413 -384
rect 22 -429 25 -423
rect 29 -429 32 -423
rect 36 -429 42 -423
rect 43 -429 49 -423
rect 50 -429 56 -423
rect 57 -429 60 -423
rect 64 -429 70 -423
rect 71 -429 74 -423
rect 78 -429 81 -423
rect 85 -429 88 -423
rect 92 -429 98 -423
rect 99 -429 105 -423
rect 106 -429 112 -423
rect 113 -429 119 -423
rect 120 -429 123 -423
rect 127 -429 130 -423
rect 134 -429 140 -423
rect 141 -429 144 -423
rect 148 -429 151 -423
rect 155 -429 161 -423
rect 162 -429 168 -423
rect 169 -429 172 -423
rect 176 -429 179 -423
rect 183 -429 186 -423
rect 190 -429 196 -423
rect 197 -429 203 -423
rect 204 -429 210 -423
rect 211 -429 217 -423
rect 218 -429 221 -423
rect 225 -429 228 -423
rect 232 -429 235 -423
rect 239 -429 245 -423
rect 246 -429 252 -423
rect 253 -429 259 -423
rect 260 -429 263 -423
rect 267 -429 270 -423
rect 274 -429 277 -423
rect 281 -429 287 -423
rect 288 -429 291 -423
rect 295 -429 298 -423
rect 302 -429 305 -423
rect 309 -429 312 -423
rect 316 -429 319 -423
rect 323 -429 326 -423
rect 330 -429 333 -423
rect 337 -429 340 -423
rect 344 -429 347 -423
rect 351 -429 357 -423
rect 358 -429 364 -423
rect 365 -429 368 -423
rect 372 -429 375 -423
rect 379 -429 382 -423
rect 22 -462 28 -456
rect 29 -462 35 -456
rect 36 -462 39 -456
rect 43 -462 46 -456
rect 50 -462 53 -456
rect 57 -462 60 -456
rect 64 -462 70 -456
rect 71 -462 77 -456
rect 78 -462 81 -456
rect 85 -462 88 -456
rect 92 -462 95 -456
rect 99 -462 102 -456
rect 106 -462 109 -456
rect 113 -462 119 -456
rect 120 -462 126 -456
rect 127 -462 133 -456
rect 134 -462 140 -456
rect 141 -462 147 -456
rect 148 -462 151 -456
rect 155 -462 161 -456
rect 162 -462 165 -456
rect 169 -462 172 -456
rect 176 -462 179 -456
rect 183 -462 189 -456
rect 190 -462 196 -456
rect 197 -462 200 -456
rect 204 -462 207 -456
rect 211 -462 217 -456
rect 218 -462 221 -456
rect 225 -462 231 -456
rect 232 -462 235 -456
rect 239 -462 242 -456
rect 246 -462 252 -456
rect 253 -462 256 -456
rect 260 -462 263 -456
rect 267 -462 270 -456
rect 274 -462 277 -456
rect 281 -462 284 -456
rect 288 -462 291 -456
rect 295 -462 298 -456
rect 302 -462 308 -456
rect 309 -462 315 -456
rect 316 -462 322 -456
rect 330 -462 333 -456
rect 351 -462 354 -456
rect 358 -462 361 -456
rect 365 -462 368 -456
rect 372 -462 378 -456
rect 36 -499 39 -493
rect 43 -499 46 -493
rect 50 -499 53 -493
rect 57 -499 60 -493
rect 64 -499 70 -493
rect 71 -499 74 -493
rect 78 -499 81 -493
rect 85 -499 88 -493
rect 92 -499 98 -493
rect 99 -499 102 -493
rect 106 -499 112 -493
rect 113 -499 119 -493
rect 120 -499 123 -493
rect 127 -499 133 -493
rect 134 -499 137 -493
rect 141 -499 144 -493
rect 148 -499 151 -493
rect 155 -499 158 -493
rect 162 -499 165 -493
rect 169 -499 175 -493
rect 176 -499 179 -493
rect 183 -499 186 -493
rect 190 -499 196 -493
rect 197 -499 203 -493
rect 204 -499 210 -493
rect 211 -499 217 -493
rect 218 -499 224 -493
rect 225 -499 228 -493
rect 232 -499 235 -493
rect 239 -499 245 -493
rect 246 -499 249 -493
rect 253 -499 256 -493
rect 260 -499 263 -493
rect 267 -499 270 -493
rect 274 -499 277 -493
rect 281 -499 287 -493
rect 288 -499 291 -493
rect 295 -499 301 -493
rect 302 -499 305 -493
rect 309 -499 315 -493
rect 316 -499 322 -493
rect 323 -499 326 -493
rect 330 -499 333 -493
rect 337 -499 343 -493
rect 344 -499 350 -493
rect 351 -499 354 -493
rect 358 -499 364 -493
rect 15 -538 18 -532
rect 22 -538 28 -532
rect 29 -538 32 -532
rect 36 -538 39 -532
rect 43 -538 46 -532
rect 50 -538 53 -532
rect 57 -538 60 -532
rect 64 -538 67 -532
rect 71 -538 77 -532
rect 78 -538 81 -532
rect 85 -538 88 -532
rect 92 -538 98 -532
rect 99 -538 105 -532
rect 106 -538 112 -532
rect 113 -538 116 -532
rect 120 -538 126 -532
rect 127 -538 133 -532
rect 134 -538 137 -532
rect 141 -538 147 -532
rect 148 -538 154 -532
rect 155 -538 161 -532
rect 162 -538 168 -532
rect 169 -538 172 -532
rect 176 -538 179 -532
rect 183 -538 189 -532
rect 190 -538 196 -532
rect 197 -538 203 -532
rect 204 -538 210 -532
rect 211 -538 214 -532
rect 218 -538 224 -532
rect 225 -538 231 -532
rect 232 -538 235 -532
rect 239 -538 242 -532
rect 246 -538 249 -532
rect 253 -538 256 -532
rect 260 -538 263 -532
rect 267 -538 270 -532
rect 274 -538 280 -532
rect 281 -538 284 -532
rect 288 -538 291 -532
rect 295 -538 298 -532
rect 302 -538 305 -532
rect 309 -538 312 -532
rect 316 -538 319 -532
rect 323 -538 326 -532
rect 330 -538 333 -532
rect 337 -538 343 -532
rect 344 -538 350 -532
rect 351 -538 354 -532
rect 358 -538 361 -532
rect 365 -538 368 -532
rect 372 -538 375 -532
rect 8 -577 11 -571
rect 15 -577 18 -571
rect 22 -577 28 -571
rect 29 -577 35 -571
rect 36 -577 42 -571
rect 43 -577 49 -571
rect 50 -577 56 -571
rect 57 -577 60 -571
rect 64 -577 67 -571
rect 71 -577 74 -571
rect 78 -577 84 -571
rect 85 -577 88 -571
rect 92 -577 95 -571
rect 99 -577 102 -571
rect 106 -577 112 -571
rect 113 -577 116 -571
rect 120 -577 126 -571
rect 127 -577 133 -571
rect 134 -577 137 -571
rect 141 -577 147 -571
rect 148 -577 154 -571
rect 155 -577 161 -571
rect 162 -577 165 -571
rect 169 -577 175 -571
rect 176 -577 179 -571
rect 183 -577 189 -571
rect 190 -577 193 -571
rect 197 -577 200 -571
rect 204 -577 207 -571
rect 211 -577 214 -571
rect 218 -577 221 -571
rect 225 -577 228 -571
rect 232 -577 238 -571
rect 239 -577 242 -571
rect 246 -577 249 -571
rect 253 -577 259 -571
rect 260 -577 263 -571
rect 267 -577 270 -571
rect 274 -577 280 -571
rect 281 -577 284 -571
rect 288 -577 294 -571
rect 295 -577 298 -571
rect 302 -577 305 -571
rect 309 -577 315 -571
rect 323 -577 326 -571
rect 351 -577 357 -571
rect 358 -577 361 -571
rect 22 -608 28 -602
rect 29 -608 32 -602
rect 36 -608 42 -602
rect 43 -608 46 -602
rect 50 -608 53 -602
rect 57 -608 60 -602
rect 64 -608 67 -602
rect 71 -608 77 -602
rect 78 -608 84 -602
rect 85 -608 88 -602
rect 92 -608 98 -602
rect 99 -608 105 -602
rect 106 -608 109 -602
rect 113 -608 119 -602
rect 120 -608 123 -602
rect 127 -608 133 -602
rect 134 -608 140 -602
rect 141 -608 144 -602
rect 148 -608 154 -602
rect 155 -608 161 -602
rect 162 -608 165 -602
rect 169 -608 172 -602
rect 176 -608 182 -602
rect 183 -608 189 -602
rect 190 -608 193 -602
rect 197 -608 200 -602
rect 204 -608 207 -602
rect 211 -608 214 -602
rect 218 -608 221 -602
rect 225 -608 231 -602
rect 232 -608 235 -602
rect 239 -608 245 -602
rect 246 -608 249 -602
rect 253 -608 256 -602
rect 260 -608 263 -602
rect 267 -608 270 -602
rect 274 -608 280 -602
rect 281 -608 284 -602
rect 288 -608 291 -602
rect 302 -608 308 -602
rect 323 -608 326 -602
rect 22 -633 28 -627
rect 50 -633 53 -627
rect 64 -633 67 -627
rect 71 -633 77 -627
rect 78 -633 84 -627
rect 85 -633 91 -627
rect 92 -633 95 -627
rect 99 -633 105 -627
rect 106 -633 112 -627
rect 113 -633 119 -627
rect 120 -633 123 -627
rect 127 -633 130 -627
rect 134 -633 137 -627
rect 141 -633 147 -627
rect 148 -633 154 -627
rect 155 -633 158 -627
rect 162 -633 165 -627
rect 169 -633 175 -627
rect 176 -633 182 -627
rect 183 -633 189 -627
rect 190 -633 193 -627
rect 197 -633 200 -627
rect 204 -633 207 -627
rect 211 -633 214 -627
rect 218 -633 221 -627
rect 225 -633 228 -627
rect 232 -633 238 -627
rect 239 -633 242 -627
rect 246 -633 252 -627
rect 253 -633 259 -627
rect 260 -633 266 -627
rect 323 -633 329 -627
rect 29 -666 32 -660
rect 36 -666 39 -660
rect 43 -666 46 -660
rect 50 -666 53 -660
rect 57 -666 63 -660
rect 64 -666 70 -660
rect 71 -666 77 -660
rect 78 -666 81 -660
rect 85 -666 88 -660
rect 92 -666 98 -660
rect 99 -666 102 -660
rect 106 -666 109 -660
rect 113 -666 119 -660
rect 120 -666 126 -660
rect 127 -666 130 -660
rect 134 -666 140 -660
rect 141 -666 147 -660
rect 148 -666 151 -660
rect 155 -666 161 -660
rect 162 -666 165 -660
rect 169 -666 175 -660
rect 176 -666 182 -660
rect 183 -666 189 -660
rect 190 -666 196 -660
rect 197 -666 203 -660
rect 204 -666 210 -660
rect 211 -666 214 -660
rect 218 -666 221 -660
rect 225 -666 228 -660
rect 232 -666 235 -660
rect 239 -666 242 -660
rect 246 -666 249 -660
rect 253 -666 256 -660
rect 260 -666 263 -660
rect 267 -666 270 -660
rect 274 -666 277 -660
rect 281 -666 284 -660
rect 288 -666 291 -660
rect 295 -666 301 -660
rect 57 -699 63 -693
rect 71 -699 77 -693
rect 78 -699 81 -693
rect 85 -699 91 -693
rect 92 -699 95 -693
rect 99 -699 102 -693
rect 106 -699 112 -693
rect 113 -699 119 -693
rect 120 -699 123 -693
rect 127 -699 130 -693
rect 134 -699 140 -693
rect 141 -699 144 -693
rect 148 -699 154 -693
rect 155 -699 161 -693
rect 162 -699 165 -693
rect 169 -699 172 -693
rect 176 -699 182 -693
rect 183 -699 189 -693
rect 190 -699 196 -693
rect 197 -699 200 -693
rect 204 -699 207 -693
rect 211 -699 217 -693
rect 218 -699 221 -693
rect 225 -699 228 -693
rect 232 -699 235 -693
rect 239 -699 242 -693
rect 246 -699 252 -693
rect 253 -699 256 -693
rect 260 -699 266 -693
rect 267 -699 270 -693
rect 274 -699 280 -693
rect 113 -722 119 -716
rect 120 -722 123 -716
rect 127 -722 133 -716
rect 134 -722 140 -716
rect 141 -722 144 -716
rect 148 -722 154 -716
rect 162 -722 165 -716
rect 169 -722 175 -716
rect 176 -722 182 -716
rect 183 -722 186 -716
rect 190 -722 196 -716
rect 197 -722 200 -716
rect 204 -722 207 -716
rect 211 -722 217 -716
rect 225 -722 231 -716
rect 239 -722 242 -716
rect 113 -737 119 -731
rect 120 -737 123 -731
rect 127 -737 133 -731
rect 134 -737 137 -731
rect 155 -737 161 -731
rect 162 -737 168 -731
rect 169 -737 172 -731
rect 176 -737 179 -731
rect 183 -737 189 -731
rect 190 -737 193 -731
rect 120 -750 126 -744
rect 127 -750 130 -744
rect 148 -750 154 -744
rect 155 -750 161 -744
rect 162 -750 165 -744
rect 169 -750 172 -744
rect 183 -750 186 -744
rect 190 -750 196 -744
<< polysilicon >>
rect 103 -5 104 -3
rect 103 -11 104 -9
rect 107 -5 108 -3
rect 128 -5 129 -3
rect 135 -5 136 -3
rect 135 -11 136 -9
rect 142 -5 143 -3
rect 142 -11 143 -9
rect 149 -11 150 -9
rect 156 -5 157 -3
rect 156 -11 157 -9
rect 163 -11 164 -9
rect 173 -11 174 -9
rect 177 -5 178 -3
rect 177 -11 178 -9
rect 184 -11 185 -9
rect 191 -5 192 -3
rect 194 -5 195 -3
rect 198 -5 199 -3
rect 198 -11 199 -9
rect 205 -5 206 -3
rect 212 -5 213 -3
rect 212 -11 213 -9
rect 79 -24 80 -22
rect 79 -30 80 -28
rect 86 -30 87 -28
rect 89 -30 90 -28
rect 96 -24 97 -22
rect 93 -30 94 -28
rect 100 -24 101 -22
rect 100 -30 101 -28
rect 110 -24 111 -22
rect 107 -30 108 -28
rect 121 -24 122 -22
rect 121 -30 122 -28
rect 128 -30 129 -28
rect 135 -24 136 -22
rect 135 -30 136 -28
rect 142 -24 143 -22
rect 142 -30 143 -28
rect 149 -24 150 -22
rect 152 -24 153 -22
rect 149 -30 150 -28
rect 156 -24 157 -22
rect 156 -30 157 -28
rect 159 -30 160 -28
rect 166 -30 167 -28
rect 170 -24 171 -22
rect 170 -30 171 -28
rect 177 -30 178 -28
rect 184 -24 185 -22
rect 184 -30 185 -28
rect 187 -30 188 -28
rect 194 -24 195 -22
rect 191 -30 192 -28
rect 198 -24 199 -22
rect 198 -30 199 -28
rect 208 -24 209 -22
rect 215 -24 216 -22
rect 219 -24 220 -22
rect 219 -30 220 -28
rect 226 -24 227 -22
rect 229 -30 230 -28
rect 233 -24 234 -22
rect 233 -30 234 -28
rect 61 -53 62 -51
rect 65 -47 66 -45
rect 65 -53 66 -51
rect 72 -47 73 -45
rect 72 -53 73 -51
rect 79 -47 80 -45
rect 82 -53 83 -51
rect 86 -47 87 -45
rect 89 -47 90 -45
rect 89 -53 90 -51
rect 93 -47 94 -45
rect 96 -53 97 -51
rect 100 -47 101 -45
rect 100 -53 101 -51
rect 110 -47 111 -45
rect 110 -53 111 -51
rect 114 -47 115 -45
rect 114 -53 115 -51
rect 121 -53 122 -51
rect 124 -53 125 -51
rect 128 -47 129 -45
rect 131 -53 132 -51
rect 135 -47 136 -45
rect 135 -53 136 -51
rect 142 -53 143 -51
rect 145 -53 146 -51
rect 149 -47 150 -45
rect 152 -47 153 -45
rect 156 -47 157 -45
rect 156 -53 157 -51
rect 163 -47 164 -45
rect 163 -53 164 -51
rect 170 -47 171 -45
rect 173 -47 174 -45
rect 170 -53 171 -51
rect 180 -47 181 -45
rect 184 -47 185 -45
rect 184 -53 185 -51
rect 191 -47 192 -45
rect 191 -53 192 -51
rect 201 -47 202 -45
rect 198 -53 199 -51
rect 201 -53 202 -51
rect 205 -47 206 -45
rect 205 -53 206 -51
rect 215 -47 216 -45
rect 212 -53 213 -51
rect 219 -47 220 -45
rect 222 -53 223 -51
rect 226 -47 227 -45
rect 226 -53 227 -51
rect 233 -47 234 -45
rect 233 -53 234 -51
rect 240 -47 241 -45
rect 240 -53 241 -51
rect 247 -47 248 -45
rect 247 -53 248 -51
rect 254 -47 255 -45
rect 254 -53 255 -51
rect 261 -47 262 -45
rect 261 -53 262 -51
rect 271 -47 272 -45
rect 275 -47 276 -45
rect 275 -53 276 -51
rect 282 -47 283 -45
rect 282 -53 283 -51
rect 30 -78 31 -76
rect 30 -84 31 -82
rect 37 -84 38 -82
rect 44 -78 45 -76
rect 44 -84 45 -82
rect 51 -78 52 -76
rect 51 -84 52 -82
rect 58 -78 59 -76
rect 58 -84 59 -82
rect 65 -78 66 -76
rect 65 -84 66 -82
rect 72 -78 73 -76
rect 75 -78 76 -76
rect 79 -78 80 -76
rect 79 -84 80 -82
rect 86 -78 87 -76
rect 86 -84 87 -82
rect 93 -78 94 -76
rect 93 -84 94 -82
rect 100 -78 101 -76
rect 103 -78 104 -76
rect 100 -84 101 -82
rect 107 -84 108 -82
rect 110 -84 111 -82
rect 114 -78 115 -76
rect 117 -78 118 -76
rect 114 -84 115 -82
rect 117 -84 118 -82
rect 121 -78 122 -76
rect 121 -84 122 -82
rect 128 -84 129 -82
rect 135 -78 136 -76
rect 138 -78 139 -76
rect 138 -84 139 -82
rect 142 -78 143 -76
rect 142 -84 143 -82
rect 149 -78 150 -76
rect 149 -84 150 -82
rect 156 -78 157 -76
rect 159 -78 160 -76
rect 163 -78 164 -76
rect 163 -84 164 -82
rect 170 -78 171 -76
rect 170 -84 171 -82
rect 177 -78 178 -76
rect 180 -78 181 -76
rect 177 -84 178 -82
rect 180 -84 181 -82
rect 184 -78 185 -76
rect 187 -78 188 -76
rect 187 -84 188 -82
rect 191 -78 192 -76
rect 191 -84 192 -82
rect 198 -78 199 -76
rect 198 -84 199 -82
rect 201 -84 202 -82
rect 205 -84 206 -82
rect 208 -84 209 -82
rect 212 -78 213 -76
rect 219 -78 220 -76
rect 219 -84 220 -82
rect 226 -78 227 -76
rect 226 -84 227 -82
rect 233 -78 234 -76
rect 233 -84 234 -82
rect 243 -78 244 -76
rect 243 -84 244 -82
rect 250 -84 251 -82
rect 254 -78 255 -76
rect 254 -84 255 -82
rect 261 -78 262 -76
rect 261 -84 262 -82
rect 268 -78 269 -76
rect 268 -84 269 -82
rect 275 -78 276 -76
rect 275 -84 276 -82
rect 282 -78 283 -76
rect 282 -84 283 -82
rect 289 -78 290 -76
rect 289 -84 290 -82
rect 299 -84 300 -82
rect 303 -78 304 -76
rect 303 -84 304 -82
rect 16 -123 17 -121
rect 16 -129 17 -127
rect 26 -123 27 -121
rect 23 -129 24 -127
rect 30 -123 31 -121
rect 30 -129 31 -127
rect 37 -123 38 -121
rect 37 -129 38 -127
rect 47 -129 48 -127
rect 51 -123 52 -121
rect 51 -129 52 -127
rect 61 -129 62 -127
rect 65 -123 66 -121
rect 68 -123 69 -121
rect 65 -129 66 -127
rect 72 -123 73 -121
rect 72 -129 73 -127
rect 79 -123 80 -121
rect 79 -129 80 -127
rect 82 -129 83 -127
rect 86 -123 87 -121
rect 86 -129 87 -127
rect 93 -123 94 -121
rect 93 -129 94 -127
rect 100 -123 101 -121
rect 103 -123 104 -121
rect 100 -129 101 -127
rect 103 -129 104 -127
rect 107 -123 108 -121
rect 107 -129 108 -127
rect 117 -123 118 -121
rect 114 -129 115 -127
rect 117 -129 118 -127
rect 124 -123 125 -121
rect 128 -123 129 -121
rect 131 -123 132 -121
rect 128 -129 129 -127
rect 131 -129 132 -127
rect 135 -123 136 -121
rect 138 -123 139 -121
rect 135 -129 136 -127
rect 142 -129 143 -127
rect 145 -129 146 -127
rect 149 -123 150 -121
rect 152 -123 153 -121
rect 152 -129 153 -127
rect 159 -123 160 -121
rect 156 -129 157 -127
rect 159 -129 160 -127
rect 170 -123 171 -121
rect 170 -129 171 -127
rect 180 -123 181 -121
rect 177 -129 178 -127
rect 180 -129 181 -127
rect 184 -123 185 -121
rect 187 -123 188 -121
rect 184 -129 185 -127
rect 187 -129 188 -127
rect 194 -123 195 -121
rect 198 -123 199 -121
rect 201 -123 202 -121
rect 198 -129 199 -127
rect 201 -129 202 -127
rect 205 -123 206 -121
rect 208 -123 209 -121
rect 205 -129 206 -127
rect 212 -123 213 -121
rect 212 -129 213 -127
rect 219 -123 220 -121
rect 219 -129 220 -127
rect 226 -123 227 -121
rect 226 -129 227 -127
rect 236 -123 237 -121
rect 233 -129 234 -127
rect 236 -129 237 -127
rect 240 -123 241 -121
rect 240 -129 241 -127
rect 247 -123 248 -121
rect 247 -129 248 -127
rect 254 -123 255 -121
rect 254 -129 255 -127
rect 261 -123 262 -121
rect 261 -129 262 -127
rect 268 -123 269 -121
rect 268 -129 269 -127
rect 275 -123 276 -121
rect 275 -129 276 -127
rect 282 -123 283 -121
rect 282 -129 283 -127
rect 289 -123 290 -121
rect 289 -129 290 -127
rect 296 -123 297 -121
rect 296 -129 297 -127
rect 303 -123 304 -121
rect 303 -129 304 -127
rect 310 -123 311 -121
rect 310 -129 311 -127
rect 317 -123 318 -121
rect 317 -129 318 -127
rect 324 -123 325 -121
rect 324 -129 325 -127
rect 331 -123 332 -121
rect 331 -129 332 -127
rect 19 -176 20 -174
rect 23 -170 24 -168
rect 26 -170 27 -168
rect 30 -170 31 -168
rect 30 -176 31 -174
rect 37 -170 38 -168
rect 44 -170 45 -168
rect 44 -176 45 -174
rect 51 -176 52 -174
rect 61 -170 62 -168
rect 58 -176 59 -174
rect 65 -170 66 -168
rect 65 -176 66 -174
rect 72 -170 73 -168
rect 72 -176 73 -174
rect 79 -170 80 -168
rect 79 -176 80 -174
rect 89 -170 90 -168
rect 86 -176 87 -174
rect 93 -170 94 -168
rect 93 -176 94 -174
rect 100 -170 101 -168
rect 100 -176 101 -174
rect 110 -170 111 -168
rect 107 -176 108 -174
rect 110 -176 111 -174
rect 114 -170 115 -168
rect 117 -170 118 -168
rect 117 -176 118 -174
rect 124 -170 125 -168
rect 124 -176 125 -174
rect 128 -170 129 -168
rect 128 -176 129 -174
rect 135 -176 136 -174
rect 142 -170 143 -168
rect 142 -176 143 -174
rect 152 -170 153 -168
rect 149 -176 150 -174
rect 159 -170 160 -168
rect 156 -176 157 -174
rect 159 -176 160 -174
rect 166 -170 167 -168
rect 170 -170 171 -168
rect 170 -176 171 -174
rect 177 -170 178 -168
rect 177 -176 178 -174
rect 184 -170 185 -168
rect 184 -176 185 -174
rect 194 -170 195 -168
rect 194 -176 195 -174
rect 201 -170 202 -168
rect 201 -176 202 -174
rect 205 -170 206 -168
rect 205 -176 206 -174
rect 208 -176 209 -174
rect 212 -170 213 -168
rect 215 -170 216 -168
rect 219 -170 220 -168
rect 219 -176 220 -174
rect 226 -170 227 -168
rect 226 -176 227 -174
rect 233 -170 234 -168
rect 236 -170 237 -168
rect 243 -170 244 -168
rect 240 -176 241 -174
rect 243 -176 244 -174
rect 247 -170 248 -168
rect 247 -176 248 -174
rect 254 -170 255 -168
rect 254 -176 255 -174
rect 261 -170 262 -168
rect 261 -176 262 -174
rect 268 -176 269 -174
rect 275 -170 276 -168
rect 275 -176 276 -174
rect 282 -170 283 -168
rect 282 -176 283 -174
rect 289 -170 290 -168
rect 289 -176 290 -174
rect 296 -170 297 -168
rect 296 -176 297 -174
rect 303 -170 304 -168
rect 303 -176 304 -174
rect 310 -170 311 -168
rect 310 -176 311 -174
rect 9 -207 10 -205
rect 9 -213 10 -211
rect 16 -207 17 -205
rect 16 -213 17 -211
rect 23 -207 24 -205
rect 33 -207 34 -205
rect 37 -207 38 -205
rect 37 -213 38 -211
rect 44 -207 45 -205
rect 44 -213 45 -211
rect 51 -207 52 -205
rect 54 -207 55 -205
rect 54 -213 55 -211
rect 58 -207 59 -205
rect 58 -213 59 -211
rect 68 -207 69 -205
rect 72 -207 73 -205
rect 72 -213 73 -211
rect 75 -213 76 -211
rect 79 -207 80 -205
rect 79 -213 80 -211
rect 86 -207 87 -205
rect 89 -207 90 -205
rect 89 -213 90 -211
rect 93 -207 94 -205
rect 93 -213 94 -211
rect 100 -207 101 -205
rect 100 -213 101 -211
rect 107 -207 108 -205
rect 110 -213 111 -211
rect 114 -207 115 -205
rect 117 -207 118 -205
rect 114 -213 115 -211
rect 117 -213 118 -211
rect 121 -207 122 -205
rect 121 -213 122 -211
rect 128 -207 129 -205
rect 128 -213 129 -211
rect 135 -207 136 -205
rect 135 -213 136 -211
rect 145 -207 146 -205
rect 142 -213 143 -211
rect 149 -207 150 -205
rect 149 -213 150 -211
rect 156 -207 157 -205
rect 156 -213 157 -211
rect 163 -207 164 -205
rect 163 -213 164 -211
rect 170 -207 171 -205
rect 170 -213 171 -211
rect 177 -207 178 -205
rect 177 -213 178 -211
rect 184 -207 185 -205
rect 187 -213 188 -211
rect 191 -207 192 -205
rect 191 -213 192 -211
rect 198 -207 199 -205
rect 198 -213 199 -211
rect 205 -207 206 -205
rect 208 -213 209 -211
rect 212 -207 213 -205
rect 215 -207 216 -205
rect 215 -213 216 -211
rect 219 -207 220 -205
rect 222 -207 223 -205
rect 219 -213 220 -211
rect 222 -213 223 -211
rect 226 -207 227 -205
rect 226 -213 227 -211
rect 236 -207 237 -205
rect 233 -213 234 -211
rect 240 -207 241 -205
rect 240 -213 241 -211
rect 247 -207 248 -205
rect 247 -213 248 -211
rect 254 -207 255 -205
rect 254 -213 255 -211
rect 261 -207 262 -205
rect 261 -213 262 -211
rect 271 -207 272 -205
rect 268 -213 269 -211
rect 275 -207 276 -205
rect 275 -213 276 -211
rect 285 -207 286 -205
rect 285 -213 286 -211
rect 289 -207 290 -205
rect 292 -207 293 -205
rect 296 -207 297 -205
rect 296 -213 297 -211
rect 303 -207 304 -205
rect 303 -213 304 -211
rect 310 -207 311 -205
rect 310 -213 311 -211
rect 317 -207 318 -205
rect 317 -213 318 -211
rect 324 -207 325 -205
rect 324 -213 325 -211
rect 331 -207 332 -205
rect 331 -213 332 -211
rect 338 -207 339 -205
rect 338 -213 339 -211
rect 345 -207 346 -205
rect 345 -213 346 -211
rect 352 -207 353 -205
rect 352 -213 353 -211
rect 359 -207 360 -205
rect 359 -213 360 -211
rect 366 -207 367 -205
rect 366 -213 367 -211
rect 373 -207 374 -205
rect 373 -213 374 -211
rect 380 -207 381 -205
rect 380 -213 381 -211
rect 387 -207 388 -205
rect 394 -207 395 -205
rect 394 -213 395 -211
rect 9 -252 10 -250
rect 9 -258 10 -256
rect 16 -252 17 -250
rect 16 -258 17 -256
rect 26 -252 27 -250
rect 30 -252 31 -250
rect 30 -258 31 -256
rect 37 -252 38 -250
rect 37 -258 38 -256
rect 44 -252 45 -250
rect 44 -258 45 -256
rect 51 -252 52 -250
rect 51 -258 52 -256
rect 58 -252 59 -250
rect 58 -258 59 -256
rect 68 -258 69 -256
rect 72 -252 73 -250
rect 72 -258 73 -256
rect 75 -258 76 -256
rect 79 -252 80 -250
rect 82 -252 83 -250
rect 82 -258 83 -256
rect 86 -252 87 -250
rect 86 -258 87 -256
rect 93 -252 94 -250
rect 93 -258 94 -256
rect 100 -258 101 -256
rect 103 -258 104 -256
rect 110 -252 111 -250
rect 107 -258 108 -256
rect 114 -252 115 -250
rect 114 -258 115 -256
rect 121 -252 122 -250
rect 124 -252 125 -250
rect 124 -258 125 -256
rect 128 -252 129 -250
rect 128 -258 129 -256
rect 135 -258 136 -256
rect 138 -258 139 -256
rect 142 -252 143 -250
rect 142 -258 143 -256
rect 152 -252 153 -250
rect 152 -258 153 -256
rect 156 -252 157 -250
rect 159 -252 160 -250
rect 159 -258 160 -256
rect 163 -252 164 -250
rect 163 -258 164 -256
rect 170 -252 171 -250
rect 170 -258 171 -256
rect 177 -252 178 -250
rect 177 -258 178 -256
rect 184 -252 185 -250
rect 184 -258 185 -256
rect 191 -252 192 -250
rect 191 -258 192 -256
rect 198 -252 199 -250
rect 201 -252 202 -250
rect 198 -258 199 -256
rect 201 -258 202 -256
rect 208 -252 209 -250
rect 205 -258 206 -256
rect 208 -258 209 -256
rect 212 -252 213 -250
rect 215 -252 216 -250
rect 215 -258 216 -256
rect 219 -252 220 -250
rect 219 -258 220 -256
rect 226 -252 227 -250
rect 229 -252 230 -250
rect 226 -258 227 -256
rect 233 -252 234 -250
rect 233 -258 234 -256
rect 240 -252 241 -250
rect 240 -258 241 -256
rect 247 -252 248 -250
rect 247 -258 248 -256
rect 254 -252 255 -250
rect 254 -258 255 -256
rect 264 -258 265 -256
rect 268 -252 269 -250
rect 268 -258 269 -256
rect 275 -252 276 -250
rect 275 -258 276 -256
rect 282 -252 283 -250
rect 282 -258 283 -256
rect 289 -252 290 -250
rect 292 -252 293 -250
rect 289 -258 290 -256
rect 296 -252 297 -250
rect 296 -258 297 -256
rect 303 -252 304 -250
rect 303 -258 304 -256
rect 310 -252 311 -250
rect 310 -258 311 -256
rect 317 -252 318 -250
rect 317 -258 318 -256
rect 324 -252 325 -250
rect 324 -258 325 -256
rect 331 -252 332 -250
rect 331 -258 332 -256
rect 338 -252 339 -250
rect 338 -258 339 -256
rect 345 -252 346 -250
rect 345 -258 346 -256
rect 352 -252 353 -250
rect 352 -258 353 -256
rect 359 -252 360 -250
rect 359 -258 360 -256
rect 366 -258 367 -256
rect 369 -258 370 -256
rect 373 -252 374 -250
rect 380 -252 381 -250
rect 380 -258 381 -256
rect 2 -299 3 -297
rect 2 -305 3 -303
rect 9 -299 10 -297
rect 9 -305 10 -303
rect 16 -299 17 -297
rect 16 -305 17 -303
rect 23 -299 24 -297
rect 23 -305 24 -303
rect 30 -299 31 -297
rect 30 -305 31 -303
rect 37 -299 38 -297
rect 37 -305 38 -303
rect 44 -299 45 -297
rect 44 -305 45 -303
rect 51 -299 52 -297
rect 54 -299 55 -297
rect 61 -299 62 -297
rect 61 -305 62 -303
rect 65 -299 66 -297
rect 65 -305 66 -303
rect 72 -299 73 -297
rect 72 -305 73 -303
rect 79 -299 80 -297
rect 82 -305 83 -303
rect 86 -299 87 -297
rect 86 -305 87 -303
rect 93 -299 94 -297
rect 93 -305 94 -303
rect 100 -299 101 -297
rect 100 -305 101 -303
rect 107 -299 108 -297
rect 107 -305 108 -303
rect 114 -299 115 -297
rect 114 -305 115 -303
rect 121 -299 122 -297
rect 124 -299 125 -297
rect 124 -305 125 -303
rect 128 -299 129 -297
rect 128 -305 129 -303
rect 135 -305 136 -303
rect 138 -305 139 -303
rect 142 -299 143 -297
rect 142 -305 143 -303
rect 149 -299 150 -297
rect 149 -305 150 -303
rect 156 -299 157 -297
rect 159 -299 160 -297
rect 156 -305 157 -303
rect 159 -305 160 -303
rect 166 -299 167 -297
rect 163 -305 164 -303
rect 166 -305 167 -303
rect 170 -299 171 -297
rect 170 -305 171 -303
rect 177 -299 178 -297
rect 177 -305 178 -303
rect 184 -299 185 -297
rect 187 -299 188 -297
rect 187 -305 188 -303
rect 191 -299 192 -297
rect 191 -305 192 -303
rect 198 -299 199 -297
rect 201 -299 202 -297
rect 201 -305 202 -303
rect 205 -299 206 -297
rect 208 -299 209 -297
rect 208 -305 209 -303
rect 212 -299 213 -297
rect 215 -299 216 -297
rect 212 -305 213 -303
rect 215 -305 216 -303
rect 219 -299 220 -297
rect 219 -305 220 -303
rect 226 -299 227 -297
rect 226 -305 227 -303
rect 233 -305 234 -303
rect 236 -305 237 -303
rect 240 -299 241 -297
rect 240 -305 241 -303
rect 243 -305 244 -303
rect 247 -299 248 -297
rect 250 -299 251 -297
rect 250 -305 251 -303
rect 257 -299 258 -297
rect 254 -305 255 -303
rect 261 -299 262 -297
rect 261 -305 262 -303
rect 268 -299 269 -297
rect 268 -305 269 -303
rect 275 -299 276 -297
rect 275 -305 276 -303
rect 282 -299 283 -297
rect 282 -305 283 -303
rect 289 -299 290 -297
rect 289 -305 290 -303
rect 296 -299 297 -297
rect 299 -305 300 -303
rect 303 -299 304 -297
rect 303 -305 304 -303
rect 310 -299 311 -297
rect 310 -305 311 -303
rect 317 -299 318 -297
rect 317 -305 318 -303
rect 324 -299 325 -297
rect 324 -305 325 -303
rect 331 -299 332 -297
rect 331 -305 332 -303
rect 338 -299 339 -297
rect 338 -305 339 -303
rect 345 -299 346 -297
rect 345 -305 346 -303
rect 352 -299 353 -297
rect 352 -305 353 -303
rect 359 -299 360 -297
rect 359 -305 360 -303
rect 366 -299 367 -297
rect 369 -299 370 -297
rect 369 -305 370 -303
rect 376 -299 377 -297
rect 376 -305 377 -303
rect 380 -299 381 -297
rect 380 -305 381 -303
rect 2 -340 3 -338
rect 2 -346 3 -344
rect 9 -340 10 -338
rect 9 -346 10 -344
rect 16 -340 17 -338
rect 16 -346 17 -344
rect 23 -340 24 -338
rect 23 -346 24 -344
rect 30 -340 31 -338
rect 30 -346 31 -344
rect 37 -340 38 -338
rect 37 -346 38 -344
rect 44 -340 45 -338
rect 44 -346 45 -344
rect 51 -340 52 -338
rect 51 -346 52 -344
rect 61 -346 62 -344
rect 65 -340 66 -338
rect 68 -340 69 -338
rect 72 -340 73 -338
rect 72 -346 73 -344
rect 79 -340 80 -338
rect 79 -346 80 -344
rect 86 -340 87 -338
rect 89 -340 90 -338
rect 89 -346 90 -344
rect 93 -340 94 -338
rect 93 -346 94 -344
rect 100 -340 101 -338
rect 100 -346 101 -344
rect 110 -340 111 -338
rect 107 -346 108 -344
rect 110 -346 111 -344
rect 114 -340 115 -338
rect 117 -340 118 -338
rect 114 -346 115 -344
rect 117 -346 118 -344
rect 124 -340 125 -338
rect 121 -346 122 -344
rect 128 -340 129 -338
rect 128 -346 129 -344
rect 135 -340 136 -338
rect 135 -346 136 -344
rect 142 -340 143 -338
rect 145 -340 146 -338
rect 142 -346 143 -344
rect 145 -346 146 -344
rect 152 -340 153 -338
rect 149 -346 150 -344
rect 156 -340 157 -338
rect 159 -340 160 -338
rect 159 -346 160 -344
rect 163 -340 164 -338
rect 163 -346 164 -344
rect 173 -340 174 -338
rect 170 -346 171 -344
rect 173 -346 174 -344
rect 177 -340 178 -338
rect 177 -346 178 -344
rect 184 -340 185 -338
rect 184 -346 185 -344
rect 194 -340 195 -338
rect 191 -346 192 -344
rect 194 -346 195 -344
rect 198 -340 199 -338
rect 198 -346 199 -344
rect 205 -340 206 -338
rect 205 -346 206 -344
rect 208 -346 209 -344
rect 212 -346 213 -344
rect 219 -340 220 -338
rect 219 -346 220 -344
rect 226 -340 227 -338
rect 226 -346 227 -344
rect 236 -346 237 -344
rect 240 -340 241 -338
rect 240 -346 241 -344
rect 243 -346 244 -344
rect 247 -340 248 -338
rect 247 -346 248 -344
rect 254 -340 255 -338
rect 254 -346 255 -344
rect 261 -340 262 -338
rect 261 -346 262 -344
rect 268 -340 269 -338
rect 268 -346 269 -344
rect 275 -340 276 -338
rect 275 -346 276 -344
rect 282 -340 283 -338
rect 282 -346 283 -344
rect 289 -340 290 -338
rect 289 -346 290 -344
rect 296 -340 297 -338
rect 296 -346 297 -344
rect 303 -340 304 -338
rect 303 -346 304 -344
rect 310 -340 311 -338
rect 310 -346 311 -344
rect 317 -340 318 -338
rect 317 -346 318 -344
rect 324 -340 325 -338
rect 324 -346 325 -344
rect 331 -340 332 -338
rect 331 -346 332 -344
rect 338 -340 339 -338
rect 345 -340 346 -338
rect 345 -346 346 -344
rect 352 -340 353 -338
rect 352 -346 353 -344
rect 359 -340 360 -338
rect 359 -346 360 -344
rect 373 -340 374 -338
rect 387 -340 388 -338
rect 387 -346 388 -344
rect 9 -385 10 -383
rect 9 -391 10 -389
rect 16 -385 17 -383
rect 16 -391 17 -389
rect 23 -385 24 -383
rect 23 -391 24 -389
rect 30 -385 31 -383
rect 30 -391 31 -389
rect 37 -385 38 -383
rect 37 -391 38 -389
rect 44 -385 45 -383
rect 44 -391 45 -389
rect 51 -385 52 -383
rect 51 -391 52 -389
rect 58 -385 59 -383
rect 58 -391 59 -389
rect 65 -385 66 -383
rect 68 -385 69 -383
rect 65 -391 66 -389
rect 72 -385 73 -383
rect 72 -391 73 -389
rect 79 -385 80 -383
rect 79 -391 80 -389
rect 86 -385 87 -383
rect 89 -385 90 -383
rect 89 -391 90 -389
rect 93 -385 94 -383
rect 96 -385 97 -383
rect 100 -385 101 -383
rect 100 -391 101 -389
rect 107 -385 108 -383
rect 107 -391 108 -389
rect 114 -385 115 -383
rect 114 -391 115 -389
rect 117 -391 118 -389
rect 121 -385 122 -383
rect 121 -391 122 -389
rect 128 -385 129 -383
rect 128 -391 129 -389
rect 131 -391 132 -389
rect 135 -385 136 -383
rect 135 -391 136 -389
rect 142 -385 143 -383
rect 145 -385 146 -383
rect 142 -391 143 -389
rect 145 -391 146 -389
rect 149 -385 150 -383
rect 152 -385 153 -383
rect 149 -391 150 -389
rect 159 -385 160 -383
rect 156 -391 157 -389
rect 159 -391 160 -389
rect 163 -385 164 -383
rect 163 -391 164 -389
rect 170 -385 171 -383
rect 173 -385 174 -383
rect 170 -391 171 -389
rect 173 -391 174 -389
rect 177 -385 178 -383
rect 177 -391 178 -389
rect 187 -385 188 -383
rect 184 -391 185 -389
rect 191 -385 192 -383
rect 194 -391 195 -389
rect 198 -385 199 -383
rect 198 -391 199 -389
rect 205 -385 206 -383
rect 205 -391 206 -389
rect 212 -385 213 -383
rect 215 -385 216 -383
rect 212 -391 213 -389
rect 219 -385 220 -383
rect 222 -385 223 -383
rect 219 -391 220 -389
rect 222 -391 223 -389
rect 226 -385 227 -383
rect 226 -391 227 -389
rect 233 -385 234 -383
rect 233 -391 234 -389
rect 240 -385 241 -383
rect 243 -385 244 -383
rect 240 -391 241 -389
rect 243 -391 244 -389
rect 247 -385 248 -383
rect 247 -391 248 -389
rect 257 -385 258 -383
rect 261 -385 262 -383
rect 261 -391 262 -389
rect 271 -385 272 -383
rect 268 -391 269 -389
rect 275 -385 276 -383
rect 275 -391 276 -389
rect 285 -385 286 -383
rect 285 -391 286 -389
rect 289 -385 290 -383
rect 289 -391 290 -389
rect 296 -385 297 -383
rect 296 -391 297 -389
rect 303 -385 304 -383
rect 303 -391 304 -389
rect 310 -385 311 -383
rect 310 -391 311 -389
rect 317 -385 318 -383
rect 317 -391 318 -389
rect 324 -385 325 -383
rect 324 -391 325 -389
rect 331 -385 332 -383
rect 331 -391 332 -389
rect 338 -385 339 -383
rect 338 -391 339 -389
rect 345 -385 346 -383
rect 345 -391 346 -389
rect 352 -385 353 -383
rect 352 -391 353 -389
rect 359 -385 360 -383
rect 359 -391 360 -389
rect 366 -385 367 -383
rect 366 -391 367 -389
rect 373 -385 374 -383
rect 373 -391 374 -389
rect 380 -385 381 -383
rect 380 -391 381 -389
rect 387 -385 388 -383
rect 387 -391 388 -389
rect 397 -385 398 -383
rect 394 -391 395 -389
rect 401 -385 402 -383
rect 401 -391 402 -389
rect 411 -391 412 -389
rect 23 -424 24 -422
rect 23 -430 24 -428
rect 30 -424 31 -422
rect 30 -430 31 -428
rect 37 -424 38 -422
rect 47 -430 48 -428
rect 51 -430 52 -428
rect 58 -424 59 -422
rect 58 -430 59 -428
rect 65 -424 66 -422
rect 68 -424 69 -422
rect 65 -430 66 -428
rect 72 -424 73 -422
rect 72 -430 73 -428
rect 79 -424 80 -422
rect 79 -430 80 -428
rect 86 -424 87 -422
rect 86 -430 87 -428
rect 93 -424 94 -422
rect 93 -430 94 -428
rect 96 -430 97 -428
rect 100 -424 101 -422
rect 100 -430 101 -428
rect 110 -424 111 -422
rect 117 -424 118 -422
rect 114 -430 115 -428
rect 121 -424 122 -422
rect 121 -430 122 -428
rect 128 -424 129 -422
rect 128 -430 129 -428
rect 135 -424 136 -422
rect 142 -424 143 -422
rect 142 -430 143 -428
rect 149 -424 150 -422
rect 149 -430 150 -428
rect 156 -424 157 -422
rect 159 -424 160 -422
rect 159 -430 160 -428
rect 163 -424 164 -422
rect 170 -424 171 -422
rect 170 -430 171 -428
rect 177 -424 178 -422
rect 177 -430 178 -428
rect 184 -424 185 -422
rect 184 -430 185 -428
rect 191 -430 192 -428
rect 194 -430 195 -428
rect 198 -424 199 -422
rect 201 -424 202 -422
rect 198 -430 199 -428
rect 205 -424 206 -422
rect 208 -424 209 -422
rect 205 -430 206 -428
rect 215 -424 216 -422
rect 212 -430 213 -428
rect 215 -430 216 -428
rect 219 -424 220 -422
rect 219 -430 220 -428
rect 226 -424 227 -422
rect 226 -430 227 -428
rect 233 -424 234 -422
rect 233 -430 234 -428
rect 243 -424 244 -422
rect 247 -424 248 -422
rect 250 -424 251 -422
rect 247 -430 248 -428
rect 257 -424 258 -422
rect 254 -430 255 -428
rect 261 -424 262 -422
rect 261 -430 262 -428
rect 268 -424 269 -422
rect 268 -430 269 -428
rect 275 -424 276 -422
rect 275 -430 276 -428
rect 282 -424 283 -422
rect 285 -424 286 -422
rect 282 -430 283 -428
rect 289 -424 290 -422
rect 289 -430 290 -428
rect 296 -424 297 -422
rect 296 -430 297 -428
rect 303 -424 304 -422
rect 303 -430 304 -428
rect 310 -424 311 -422
rect 310 -430 311 -428
rect 317 -424 318 -422
rect 317 -430 318 -428
rect 324 -424 325 -422
rect 324 -430 325 -428
rect 331 -424 332 -422
rect 331 -430 332 -428
rect 338 -424 339 -422
rect 338 -430 339 -428
rect 345 -424 346 -422
rect 345 -430 346 -428
rect 352 -424 353 -422
rect 352 -430 353 -428
rect 355 -430 356 -428
rect 359 -424 360 -422
rect 362 -430 363 -428
rect 366 -424 367 -422
rect 366 -430 367 -428
rect 373 -424 374 -422
rect 373 -430 374 -428
rect 380 -424 381 -422
rect 380 -430 381 -428
rect 26 -463 27 -461
rect 33 -463 34 -461
rect 37 -457 38 -455
rect 37 -463 38 -461
rect 44 -457 45 -455
rect 44 -463 45 -461
rect 51 -457 52 -455
rect 51 -463 52 -461
rect 58 -457 59 -455
rect 58 -463 59 -461
rect 65 -457 66 -455
rect 68 -457 69 -455
rect 75 -457 76 -455
rect 72 -463 73 -461
rect 79 -457 80 -455
rect 79 -463 80 -461
rect 86 -457 87 -455
rect 86 -463 87 -461
rect 93 -457 94 -455
rect 93 -463 94 -461
rect 100 -457 101 -455
rect 100 -463 101 -461
rect 107 -457 108 -455
rect 107 -463 108 -461
rect 114 -457 115 -455
rect 117 -457 118 -455
rect 114 -463 115 -461
rect 117 -463 118 -461
rect 124 -457 125 -455
rect 121 -463 122 -461
rect 131 -457 132 -455
rect 128 -463 129 -461
rect 131 -463 132 -461
rect 135 -457 136 -455
rect 135 -463 136 -461
rect 138 -463 139 -461
rect 142 -457 143 -455
rect 145 -463 146 -461
rect 149 -457 150 -455
rect 149 -463 150 -461
rect 156 -457 157 -455
rect 159 -457 160 -455
rect 163 -457 164 -455
rect 163 -463 164 -461
rect 170 -457 171 -455
rect 170 -463 171 -461
rect 177 -457 178 -455
rect 177 -463 178 -461
rect 184 -457 185 -455
rect 187 -457 188 -455
rect 187 -463 188 -461
rect 191 -457 192 -455
rect 194 -457 195 -455
rect 191 -463 192 -461
rect 194 -463 195 -461
rect 198 -457 199 -455
rect 198 -463 199 -461
rect 205 -457 206 -455
rect 205 -463 206 -461
rect 212 -457 213 -455
rect 215 -457 216 -455
rect 212 -463 213 -461
rect 219 -457 220 -455
rect 219 -463 220 -461
rect 229 -457 230 -455
rect 226 -463 227 -461
rect 229 -463 230 -461
rect 233 -457 234 -455
rect 233 -463 234 -461
rect 240 -457 241 -455
rect 240 -463 241 -461
rect 250 -463 251 -461
rect 254 -457 255 -455
rect 254 -463 255 -461
rect 261 -457 262 -455
rect 261 -463 262 -461
rect 268 -457 269 -455
rect 268 -463 269 -461
rect 275 -457 276 -455
rect 275 -463 276 -461
rect 282 -457 283 -455
rect 282 -463 283 -461
rect 289 -457 290 -455
rect 289 -463 290 -461
rect 296 -457 297 -455
rect 296 -463 297 -461
rect 303 -457 304 -455
rect 306 -457 307 -455
rect 306 -463 307 -461
rect 313 -457 314 -455
rect 320 -457 321 -455
rect 317 -463 318 -461
rect 331 -457 332 -455
rect 331 -463 332 -461
rect 352 -457 353 -455
rect 352 -463 353 -461
rect 359 -457 360 -455
rect 359 -463 360 -461
rect 366 -457 367 -455
rect 366 -463 367 -461
rect 376 -463 377 -461
rect 37 -494 38 -492
rect 37 -500 38 -498
rect 44 -494 45 -492
rect 44 -500 45 -498
rect 51 -494 52 -492
rect 51 -500 52 -498
rect 58 -494 59 -492
rect 58 -500 59 -498
rect 65 -494 66 -492
rect 68 -494 69 -492
rect 65 -500 66 -498
rect 68 -500 69 -498
rect 72 -494 73 -492
rect 72 -500 73 -498
rect 79 -494 80 -492
rect 79 -500 80 -498
rect 86 -494 87 -492
rect 86 -500 87 -498
rect 93 -500 94 -498
rect 100 -494 101 -492
rect 100 -500 101 -498
rect 110 -494 111 -492
rect 107 -500 108 -498
rect 110 -500 111 -498
rect 114 -494 115 -492
rect 114 -500 115 -498
rect 121 -494 122 -492
rect 121 -500 122 -498
rect 128 -494 129 -492
rect 131 -494 132 -492
rect 135 -494 136 -492
rect 135 -500 136 -498
rect 142 -494 143 -492
rect 142 -500 143 -498
rect 149 -494 150 -492
rect 149 -500 150 -498
rect 156 -494 157 -492
rect 156 -500 157 -498
rect 163 -494 164 -492
rect 163 -500 164 -498
rect 170 -494 171 -492
rect 173 -494 174 -492
rect 173 -500 174 -498
rect 177 -494 178 -492
rect 177 -500 178 -498
rect 184 -494 185 -492
rect 184 -500 185 -498
rect 194 -500 195 -498
rect 198 -494 199 -492
rect 198 -500 199 -498
rect 201 -500 202 -498
rect 205 -494 206 -492
rect 208 -494 209 -492
rect 215 -494 216 -492
rect 212 -500 213 -498
rect 219 -500 220 -498
rect 226 -494 227 -492
rect 226 -500 227 -498
rect 233 -494 234 -492
rect 233 -500 234 -498
rect 240 -494 241 -492
rect 243 -494 244 -492
rect 240 -500 241 -498
rect 243 -500 244 -498
rect 247 -494 248 -492
rect 247 -500 248 -498
rect 254 -494 255 -492
rect 254 -500 255 -498
rect 261 -494 262 -492
rect 261 -500 262 -498
rect 268 -494 269 -492
rect 268 -500 269 -498
rect 275 -494 276 -492
rect 275 -500 276 -498
rect 282 -500 283 -498
rect 289 -494 290 -492
rect 289 -500 290 -498
rect 296 -500 297 -498
rect 299 -500 300 -498
rect 303 -494 304 -492
rect 303 -500 304 -498
rect 313 -500 314 -498
rect 320 -494 321 -492
rect 324 -494 325 -492
rect 324 -500 325 -498
rect 331 -494 332 -492
rect 331 -500 332 -498
rect 338 -494 339 -492
rect 341 -500 342 -498
rect 348 -494 349 -492
rect 348 -500 349 -498
rect 352 -494 353 -492
rect 352 -500 353 -498
rect 359 -494 360 -492
rect 16 -533 17 -531
rect 16 -539 17 -537
rect 26 -539 27 -537
rect 30 -533 31 -531
rect 30 -539 31 -537
rect 37 -533 38 -531
rect 37 -539 38 -537
rect 44 -533 45 -531
rect 44 -539 45 -537
rect 51 -533 52 -531
rect 51 -539 52 -537
rect 58 -533 59 -531
rect 58 -539 59 -537
rect 65 -533 66 -531
rect 65 -539 66 -537
rect 72 -533 73 -531
rect 79 -533 80 -531
rect 79 -539 80 -537
rect 86 -533 87 -531
rect 86 -539 87 -537
rect 93 -533 94 -531
rect 93 -539 94 -537
rect 100 -533 101 -531
rect 100 -539 101 -537
rect 103 -539 104 -537
rect 110 -533 111 -531
rect 110 -539 111 -537
rect 114 -533 115 -531
rect 114 -539 115 -537
rect 124 -539 125 -537
rect 131 -533 132 -531
rect 128 -539 129 -537
rect 131 -539 132 -537
rect 135 -533 136 -531
rect 135 -539 136 -537
rect 142 -533 143 -531
rect 145 -539 146 -537
rect 149 -533 150 -531
rect 149 -539 150 -537
rect 152 -539 153 -537
rect 156 -533 157 -531
rect 159 -533 160 -531
rect 156 -539 157 -537
rect 163 -533 164 -531
rect 166 -533 167 -531
rect 166 -539 167 -537
rect 170 -533 171 -531
rect 170 -539 171 -537
rect 177 -533 178 -531
rect 177 -539 178 -537
rect 184 -533 185 -531
rect 191 -533 192 -531
rect 194 -533 195 -531
rect 198 -533 199 -531
rect 201 -533 202 -531
rect 198 -539 199 -537
rect 201 -539 202 -537
rect 205 -533 206 -531
rect 208 -533 209 -531
rect 205 -539 206 -537
rect 208 -539 209 -537
rect 212 -533 213 -531
rect 212 -539 213 -537
rect 219 -533 220 -531
rect 222 -533 223 -531
rect 222 -539 223 -537
rect 226 -533 227 -531
rect 229 -533 230 -531
rect 229 -539 230 -537
rect 233 -533 234 -531
rect 233 -539 234 -537
rect 240 -533 241 -531
rect 240 -539 241 -537
rect 247 -533 248 -531
rect 247 -539 248 -537
rect 254 -533 255 -531
rect 254 -539 255 -537
rect 261 -533 262 -531
rect 261 -539 262 -537
rect 268 -533 269 -531
rect 268 -539 269 -537
rect 275 -539 276 -537
rect 278 -539 279 -537
rect 282 -533 283 -531
rect 282 -539 283 -537
rect 289 -533 290 -531
rect 289 -539 290 -537
rect 296 -533 297 -531
rect 296 -539 297 -537
rect 303 -533 304 -531
rect 303 -539 304 -537
rect 310 -533 311 -531
rect 310 -539 311 -537
rect 317 -533 318 -531
rect 317 -539 318 -537
rect 324 -533 325 -531
rect 324 -539 325 -537
rect 331 -533 332 -531
rect 331 -539 332 -537
rect 338 -533 339 -531
rect 341 -533 342 -531
rect 338 -539 339 -537
rect 345 -533 346 -531
rect 348 -533 349 -531
rect 345 -539 346 -537
rect 348 -539 349 -537
rect 352 -533 353 -531
rect 352 -539 353 -537
rect 359 -533 360 -531
rect 359 -539 360 -537
rect 366 -533 367 -531
rect 366 -539 367 -537
rect 373 -533 374 -531
rect 373 -539 374 -537
rect 9 -572 10 -570
rect 9 -578 10 -576
rect 16 -572 17 -570
rect 16 -578 17 -576
rect 23 -572 24 -570
rect 23 -578 24 -576
rect 33 -578 34 -576
rect 40 -578 41 -576
rect 44 -572 45 -570
rect 44 -578 45 -576
rect 51 -578 52 -576
rect 58 -572 59 -570
rect 58 -578 59 -576
rect 65 -572 66 -570
rect 65 -578 66 -576
rect 72 -572 73 -570
rect 72 -578 73 -576
rect 82 -572 83 -570
rect 79 -578 80 -576
rect 82 -578 83 -576
rect 86 -572 87 -570
rect 86 -578 87 -576
rect 93 -572 94 -570
rect 93 -578 94 -576
rect 100 -572 101 -570
rect 100 -578 101 -576
rect 107 -572 108 -570
rect 107 -578 108 -576
rect 110 -578 111 -576
rect 114 -572 115 -570
rect 114 -578 115 -576
rect 121 -572 122 -570
rect 124 -572 125 -570
rect 131 -572 132 -570
rect 131 -578 132 -576
rect 135 -572 136 -570
rect 135 -578 136 -576
rect 142 -572 143 -570
rect 145 -572 146 -570
rect 145 -578 146 -576
rect 152 -572 153 -570
rect 152 -578 153 -576
rect 159 -572 160 -570
rect 159 -578 160 -576
rect 163 -572 164 -570
rect 163 -578 164 -576
rect 170 -572 171 -570
rect 177 -572 178 -570
rect 177 -578 178 -576
rect 187 -578 188 -576
rect 191 -572 192 -570
rect 191 -578 192 -576
rect 198 -572 199 -570
rect 198 -578 199 -576
rect 205 -572 206 -570
rect 205 -578 206 -576
rect 212 -572 213 -570
rect 212 -578 213 -576
rect 219 -572 220 -570
rect 219 -578 220 -576
rect 226 -572 227 -570
rect 226 -578 227 -576
rect 236 -572 237 -570
rect 240 -572 241 -570
rect 240 -578 241 -576
rect 247 -572 248 -570
rect 247 -578 248 -576
rect 257 -578 258 -576
rect 261 -572 262 -570
rect 261 -578 262 -576
rect 268 -572 269 -570
rect 268 -578 269 -576
rect 275 -572 276 -570
rect 278 -572 279 -570
rect 282 -572 283 -570
rect 282 -578 283 -576
rect 289 -572 290 -570
rect 292 -572 293 -570
rect 296 -572 297 -570
rect 296 -578 297 -576
rect 303 -572 304 -570
rect 303 -578 304 -576
rect 310 -578 311 -576
rect 324 -572 325 -570
rect 324 -578 325 -576
rect 355 -578 356 -576
rect 359 -572 360 -570
rect 359 -578 360 -576
rect 23 -603 24 -601
rect 26 -609 27 -607
rect 30 -603 31 -601
rect 30 -609 31 -607
rect 40 -603 41 -601
rect 37 -609 38 -607
rect 44 -603 45 -601
rect 44 -609 45 -607
rect 51 -603 52 -601
rect 51 -609 52 -607
rect 58 -603 59 -601
rect 58 -609 59 -607
rect 65 -603 66 -601
rect 65 -609 66 -607
rect 75 -603 76 -601
rect 75 -609 76 -607
rect 79 -603 80 -601
rect 79 -609 80 -607
rect 82 -609 83 -607
rect 86 -603 87 -601
rect 86 -609 87 -607
rect 93 -603 94 -601
rect 96 -603 97 -601
rect 100 -603 101 -601
rect 100 -609 101 -607
rect 107 -603 108 -601
rect 107 -609 108 -607
rect 114 -603 115 -601
rect 114 -609 115 -607
rect 117 -609 118 -607
rect 121 -603 122 -601
rect 121 -609 122 -607
rect 128 -603 129 -601
rect 131 -609 132 -607
rect 135 -603 136 -601
rect 138 -603 139 -601
rect 135 -609 136 -607
rect 138 -609 139 -607
rect 142 -603 143 -601
rect 142 -609 143 -607
rect 149 -603 150 -601
rect 152 -603 153 -601
rect 149 -609 150 -607
rect 152 -609 153 -607
rect 156 -603 157 -601
rect 159 -603 160 -601
rect 156 -609 157 -607
rect 159 -609 160 -607
rect 163 -603 164 -601
rect 163 -609 164 -607
rect 170 -603 171 -601
rect 170 -609 171 -607
rect 177 -603 178 -601
rect 177 -609 178 -607
rect 180 -609 181 -607
rect 184 -603 185 -601
rect 187 -603 188 -601
rect 191 -603 192 -601
rect 191 -609 192 -607
rect 198 -603 199 -601
rect 198 -609 199 -607
rect 205 -603 206 -601
rect 205 -609 206 -607
rect 212 -603 213 -601
rect 212 -609 213 -607
rect 219 -603 220 -601
rect 219 -609 220 -607
rect 229 -603 230 -601
rect 226 -609 227 -607
rect 233 -603 234 -601
rect 233 -609 234 -607
rect 243 -609 244 -607
rect 247 -603 248 -601
rect 247 -609 248 -607
rect 254 -603 255 -601
rect 254 -609 255 -607
rect 261 -603 262 -601
rect 261 -609 262 -607
rect 268 -603 269 -601
rect 268 -609 269 -607
rect 278 -603 279 -601
rect 275 -609 276 -607
rect 282 -603 283 -601
rect 282 -609 283 -607
rect 289 -603 290 -601
rect 289 -609 290 -607
rect 303 -603 304 -601
rect 306 -603 307 -601
rect 324 -603 325 -601
rect 324 -609 325 -607
rect 26 -628 27 -626
rect 51 -628 52 -626
rect 51 -634 52 -632
rect 65 -628 66 -626
rect 65 -634 66 -632
rect 72 -628 73 -626
rect 75 -634 76 -632
rect 79 -628 80 -626
rect 82 -634 83 -632
rect 86 -628 87 -626
rect 93 -628 94 -626
rect 93 -634 94 -632
rect 103 -628 104 -626
rect 100 -634 101 -632
rect 107 -628 108 -626
rect 107 -634 108 -632
rect 114 -628 115 -626
rect 117 -628 118 -626
rect 121 -628 122 -626
rect 121 -634 122 -632
rect 128 -628 129 -626
rect 128 -634 129 -632
rect 135 -628 136 -626
rect 135 -634 136 -632
rect 142 -628 143 -626
rect 145 -628 146 -626
rect 145 -634 146 -632
rect 149 -634 150 -632
rect 152 -634 153 -632
rect 156 -628 157 -626
rect 156 -634 157 -632
rect 163 -628 164 -626
rect 163 -634 164 -632
rect 173 -628 174 -626
rect 180 -628 181 -626
rect 184 -628 185 -626
rect 187 -628 188 -626
rect 187 -634 188 -632
rect 191 -628 192 -626
rect 191 -634 192 -632
rect 198 -628 199 -626
rect 198 -634 199 -632
rect 205 -628 206 -626
rect 205 -634 206 -632
rect 212 -628 213 -626
rect 212 -634 213 -632
rect 219 -628 220 -626
rect 219 -634 220 -632
rect 226 -628 227 -626
rect 226 -634 227 -632
rect 233 -628 234 -626
rect 233 -634 234 -632
rect 236 -634 237 -632
rect 240 -628 241 -626
rect 240 -634 241 -632
rect 247 -628 248 -626
rect 247 -634 248 -632
rect 254 -628 255 -626
rect 257 -628 258 -626
rect 257 -634 258 -632
rect 261 -628 262 -626
rect 264 -628 265 -626
rect 324 -628 325 -626
rect 30 -661 31 -659
rect 30 -667 31 -665
rect 37 -661 38 -659
rect 37 -667 38 -665
rect 44 -661 45 -659
rect 44 -667 45 -665
rect 51 -661 52 -659
rect 51 -667 52 -665
rect 58 -667 59 -665
rect 61 -667 62 -665
rect 68 -661 69 -659
rect 68 -667 69 -665
rect 72 -661 73 -659
rect 75 -661 76 -659
rect 79 -661 80 -659
rect 79 -667 80 -665
rect 86 -661 87 -659
rect 86 -667 87 -665
rect 96 -661 97 -659
rect 93 -667 94 -665
rect 96 -667 97 -665
rect 100 -661 101 -659
rect 100 -667 101 -665
rect 107 -661 108 -659
rect 107 -667 108 -665
rect 117 -661 118 -659
rect 114 -667 115 -665
rect 117 -667 118 -665
rect 121 -661 122 -659
rect 124 -661 125 -659
rect 128 -661 129 -659
rect 128 -667 129 -665
rect 135 -661 136 -659
rect 138 -661 139 -659
rect 138 -667 139 -665
rect 142 -661 143 -659
rect 145 -667 146 -665
rect 149 -661 150 -659
rect 149 -667 150 -665
rect 156 -661 157 -659
rect 156 -667 157 -665
rect 159 -667 160 -665
rect 163 -661 164 -659
rect 163 -667 164 -665
rect 170 -661 171 -659
rect 173 -661 174 -659
rect 173 -667 174 -665
rect 177 -667 178 -665
rect 180 -667 181 -665
rect 184 -661 185 -659
rect 187 -661 188 -659
rect 184 -667 185 -665
rect 191 -661 192 -659
rect 191 -667 192 -665
rect 201 -661 202 -659
rect 201 -667 202 -665
rect 205 -667 206 -665
rect 208 -667 209 -665
rect 212 -661 213 -659
rect 212 -667 213 -665
rect 219 -661 220 -659
rect 219 -667 220 -665
rect 226 -661 227 -659
rect 226 -667 227 -665
rect 233 -661 234 -659
rect 233 -667 234 -665
rect 240 -661 241 -659
rect 240 -667 241 -665
rect 247 -661 248 -659
rect 247 -667 248 -665
rect 254 -661 255 -659
rect 254 -667 255 -665
rect 261 -661 262 -659
rect 261 -667 262 -665
rect 268 -661 269 -659
rect 268 -667 269 -665
rect 275 -661 276 -659
rect 275 -667 276 -665
rect 282 -661 283 -659
rect 282 -667 283 -665
rect 289 -661 290 -659
rect 289 -667 290 -665
rect 296 -661 297 -659
rect 61 -694 62 -692
rect 61 -700 62 -698
rect 72 -700 73 -698
rect 75 -700 76 -698
rect 79 -694 80 -692
rect 79 -700 80 -698
rect 89 -694 90 -692
rect 93 -694 94 -692
rect 93 -700 94 -698
rect 100 -694 101 -692
rect 100 -700 101 -698
rect 107 -694 108 -692
rect 110 -694 111 -692
rect 114 -700 115 -698
rect 117 -700 118 -698
rect 121 -694 122 -692
rect 121 -700 122 -698
rect 128 -694 129 -692
rect 128 -700 129 -698
rect 138 -694 139 -692
rect 142 -694 143 -692
rect 142 -700 143 -698
rect 152 -700 153 -698
rect 156 -694 157 -692
rect 163 -694 164 -692
rect 163 -700 164 -698
rect 170 -694 171 -692
rect 170 -700 171 -698
rect 177 -694 178 -692
rect 180 -694 181 -692
rect 177 -700 178 -698
rect 187 -694 188 -692
rect 187 -700 188 -698
rect 191 -694 192 -692
rect 194 -700 195 -698
rect 198 -694 199 -692
rect 198 -700 199 -698
rect 205 -694 206 -692
rect 205 -700 206 -698
rect 212 -694 213 -692
rect 219 -694 220 -692
rect 219 -700 220 -698
rect 226 -694 227 -692
rect 226 -700 227 -698
rect 233 -694 234 -692
rect 233 -700 234 -698
rect 240 -694 241 -692
rect 240 -700 241 -698
rect 247 -700 248 -698
rect 254 -694 255 -692
rect 254 -700 255 -698
rect 261 -700 262 -698
rect 268 -694 269 -692
rect 268 -700 269 -698
rect 278 -694 279 -692
rect 114 -723 115 -721
rect 121 -717 122 -715
rect 121 -723 122 -721
rect 131 -717 132 -715
rect 131 -723 132 -721
rect 135 -717 136 -715
rect 142 -717 143 -715
rect 142 -723 143 -721
rect 149 -717 150 -715
rect 163 -717 164 -715
rect 163 -723 164 -721
rect 170 -717 171 -715
rect 173 -717 174 -715
rect 173 -723 174 -721
rect 180 -717 181 -715
rect 177 -723 178 -721
rect 180 -723 181 -721
rect 184 -717 185 -715
rect 184 -723 185 -721
rect 194 -717 195 -715
rect 191 -723 192 -721
rect 194 -723 195 -721
rect 198 -717 199 -715
rect 198 -723 199 -721
rect 205 -717 206 -715
rect 205 -723 206 -721
rect 215 -717 216 -715
rect 229 -723 230 -721
rect 240 -717 241 -715
rect 240 -723 241 -721
rect 117 -732 118 -730
rect 121 -732 122 -730
rect 121 -738 122 -736
rect 131 -732 132 -730
rect 128 -738 129 -736
rect 135 -732 136 -730
rect 135 -738 136 -736
rect 159 -732 160 -730
rect 156 -738 157 -736
rect 166 -738 167 -736
rect 170 -732 171 -730
rect 170 -738 171 -736
rect 177 -732 178 -730
rect 177 -738 178 -736
rect 184 -732 185 -730
rect 187 -738 188 -736
rect 191 -732 192 -730
rect 191 -738 192 -736
rect 124 -751 125 -749
rect 128 -745 129 -743
rect 128 -751 129 -749
rect 149 -745 150 -743
rect 156 -751 157 -749
rect 159 -751 160 -749
rect 163 -745 164 -743
rect 163 -751 164 -749
rect 170 -745 171 -743
rect 170 -751 171 -749
rect 184 -745 185 -743
rect 184 -751 185 -749
rect 191 -751 192 -749
<< metal1 >>
rect 103 0 108 1
rect 128 0 136 1
rect 142 0 157 1
rect 177 0 192 1
rect 194 0 213 1
rect 198 -2 206 -1
rect 79 -13 97 -12
rect 100 -13 104 -12
rect 110 -13 122 -12
rect 135 -13 143 -12
rect 149 -13 157 -12
rect 170 -13 195 -12
rect 208 -13 234 -12
rect 135 -15 157 -14
rect 177 -15 185 -14
rect 212 -15 227 -14
rect 142 -17 174 -16
rect 184 -17 199 -16
rect 215 -17 220 -16
rect 149 -19 164 -18
rect 152 -21 199 -20
rect 65 -32 90 -31
rect 93 -32 97 -31
rect 114 -32 174 -31
rect 184 -32 248 -31
rect 271 -32 276 -31
rect 72 -34 111 -33
rect 142 -34 188 -33
rect 198 -34 227 -33
rect 229 -34 283 -33
rect 86 -36 90 -35
rect 93 -36 101 -35
rect 149 -36 171 -35
rect 180 -36 185 -35
rect 201 -36 255 -35
rect 86 -38 108 -37
rect 135 -38 150 -37
rect 152 -38 241 -37
rect 96 -40 101 -39
rect 121 -40 136 -39
rect 156 -40 164 -39
rect 215 -40 220 -39
rect 233 -40 262 -39
rect 156 -42 171 -41
rect 191 -42 234 -41
rect 159 -44 167 -43
rect 177 -44 192 -43
rect 205 -44 220 -43
rect 30 -55 76 -54
rect 82 -55 146 -54
rect 170 -55 262 -54
rect 44 -57 115 -56
rect 117 -57 150 -56
rect 163 -57 171 -56
rect 184 -57 262 -56
rect 51 -59 132 -58
rect 159 -59 164 -58
rect 187 -59 290 -58
rect 58 -61 157 -60
rect 191 -61 199 -60
rect 201 -61 241 -60
rect 243 -61 304 -60
rect 61 -63 90 -62
rect 93 -63 178 -62
rect 198 -63 227 -62
rect 233 -63 269 -62
rect 65 -65 87 -64
rect 100 -65 115 -64
rect 121 -65 136 -64
rect 142 -65 192 -64
rect 219 -65 276 -64
rect 65 -67 97 -66
rect 100 -67 139 -66
rect 180 -67 227 -66
rect 254 -67 276 -66
rect 72 -69 136 -68
rect 184 -69 234 -68
rect 72 -71 80 -70
rect 103 -71 143 -70
rect 212 -71 255 -70
rect 110 -73 125 -72
rect 205 -73 213 -72
rect 222 -73 283 -72
rect 121 -75 157 -74
rect 247 -75 283 -74
rect 16 -86 80 -85
rect 86 -86 101 -85
rect 103 -86 108 -85
rect 114 -86 136 -85
rect 170 -86 181 -85
rect 184 -86 195 -85
rect 201 -86 237 -85
rect 243 -86 283 -85
rect 299 -86 332 -85
rect 30 -88 325 -87
rect 26 -90 31 -89
rect 37 -90 80 -89
rect 100 -90 209 -89
rect 250 -90 290 -89
rect 37 -92 94 -91
rect 107 -92 125 -91
rect 131 -92 227 -91
rect 268 -92 311 -91
rect 44 -94 111 -93
rect 138 -94 283 -93
rect 51 -96 188 -95
rect 191 -96 241 -95
rect 275 -96 318 -95
rect 58 -98 129 -97
rect 142 -98 290 -97
rect 65 -100 87 -99
rect 93 -100 139 -99
rect 163 -100 171 -99
rect 177 -100 262 -99
rect 51 -102 66 -101
rect 68 -102 160 -101
rect 180 -102 213 -101
rect 219 -102 227 -101
rect 72 -104 118 -103
rect 128 -104 153 -103
rect 187 -104 262 -103
rect 117 -106 269 -105
rect 198 -108 276 -107
rect 198 -110 304 -109
rect 149 -112 304 -111
rect 121 -114 150 -113
rect 201 -114 234 -113
rect 205 -116 297 -115
rect 205 -118 248 -117
rect 208 -120 220 -119
rect 23 -131 146 -130
rect 159 -131 241 -130
rect 26 -133 31 -132
rect 37 -133 181 -132
rect 198 -133 248 -132
rect 23 -135 31 -134
rect 44 -135 52 -134
rect 61 -135 90 -134
rect 100 -135 283 -134
rect 37 -137 62 -136
rect 65 -137 325 -136
rect 47 -139 66 -138
rect 72 -139 83 -138
rect 86 -139 118 -138
rect 128 -139 244 -138
rect 72 -141 94 -140
rect 100 -141 108 -140
rect 110 -141 115 -140
rect 117 -141 125 -140
rect 128 -141 153 -140
rect 166 -141 195 -140
rect 205 -141 269 -140
rect 16 -143 115 -142
rect 135 -143 290 -142
rect 79 -145 94 -144
rect 142 -145 304 -144
rect 79 -147 153 -146
rect 170 -147 185 -146
rect 205 -147 311 -146
rect 131 -149 171 -148
rect 177 -149 188 -148
rect 201 -149 311 -148
rect 103 -151 178 -150
rect 201 -151 290 -150
rect 303 -151 332 -150
rect 142 -153 160 -152
rect 215 -153 297 -152
rect 156 -155 185 -154
rect 226 -155 230 -154
rect 233 -155 297 -154
rect 212 -157 234 -156
rect 236 -157 318 -156
rect 212 -159 248 -158
rect 226 -161 262 -160
rect 236 -163 283 -162
rect 254 -165 262 -164
rect 229 -167 255 -166
rect 16 -178 34 -177
rect 37 -178 69 -177
rect 72 -178 87 -177
rect 89 -178 111 -177
rect 121 -178 129 -177
rect 135 -178 143 -177
rect 145 -178 395 -177
rect 9 -180 87 -179
rect 149 -180 199 -179
rect 222 -180 297 -179
rect 303 -180 360 -179
rect 19 -182 59 -181
rect 72 -182 136 -181
rect 149 -182 185 -181
rect 191 -182 216 -181
rect 240 -182 262 -181
rect 268 -182 332 -181
rect 23 -184 31 -183
rect 44 -184 52 -183
rect 54 -184 59 -183
rect 79 -184 108 -183
rect 117 -184 241 -183
rect 243 -184 325 -183
rect 44 -186 185 -185
rect 194 -186 227 -185
rect 247 -186 262 -185
rect 271 -186 304 -185
rect 310 -186 374 -185
rect 51 -188 94 -187
rect 107 -188 237 -187
rect 247 -188 388 -187
rect 65 -190 80 -189
rect 93 -190 206 -189
rect 212 -190 311 -189
rect 117 -192 125 -191
rect 156 -192 164 -191
rect 170 -192 206 -191
rect 275 -192 297 -191
rect 114 -194 276 -193
rect 282 -194 339 -193
rect 128 -196 157 -195
rect 159 -196 220 -195
rect 285 -196 353 -195
rect 170 -198 209 -197
rect 219 -198 381 -197
rect 177 -200 227 -199
rect 289 -200 346 -199
rect 177 -202 255 -201
rect 289 -202 318 -201
rect 201 -204 255 -203
rect 292 -204 367 -203
rect 9 -215 143 -214
rect 149 -215 185 -214
rect 187 -215 346 -214
rect 9 -217 76 -216
rect 86 -217 101 -216
rect 114 -217 136 -216
rect 156 -217 171 -216
rect 177 -217 216 -216
rect 222 -217 374 -216
rect 16 -219 55 -218
rect 72 -219 80 -218
rect 93 -219 160 -218
rect 163 -219 234 -218
rect 261 -219 283 -218
rect 289 -219 325 -218
rect 16 -221 125 -220
rect 128 -221 143 -220
rect 170 -221 220 -220
rect 229 -221 360 -220
rect 26 -223 111 -222
rect 117 -223 381 -222
rect 30 -225 192 -224
rect 215 -225 297 -224
rect 366 -225 381 -224
rect 37 -227 164 -226
rect 191 -227 255 -226
rect 268 -227 339 -226
rect 37 -229 122 -228
rect 128 -229 213 -228
rect 219 -229 227 -228
rect 233 -229 248 -228
rect 254 -229 286 -228
rect 292 -229 346 -228
rect 44 -231 178 -230
rect 198 -231 269 -230
rect 296 -231 304 -230
rect 44 -233 83 -232
rect 89 -233 360 -232
rect 51 -235 59 -234
rect 72 -235 80 -234
rect 93 -235 111 -234
rect 114 -235 227 -234
rect 240 -235 325 -234
rect 58 -237 153 -236
rect 156 -237 248 -236
rect 303 -237 311 -236
rect 121 -239 395 -238
rect 198 -241 332 -240
rect 208 -243 339 -242
rect 208 -245 276 -244
rect 310 -245 318 -244
rect 331 -245 374 -244
rect 201 -247 318 -246
rect 240 -249 276 -248
rect 2 -260 125 -259
rect 138 -260 255 -259
rect 264 -260 297 -259
rect 359 -260 370 -259
rect 376 -260 381 -259
rect 9 -262 76 -261
rect 79 -262 108 -261
rect 121 -262 157 -261
rect 166 -262 262 -261
rect 275 -262 332 -261
rect 366 -262 370 -261
rect 9 -264 59 -263
rect 65 -264 129 -263
rect 149 -264 178 -263
rect 184 -264 258 -263
rect 275 -264 283 -263
rect 289 -264 353 -263
rect 366 -264 381 -263
rect 16 -266 101 -265
rect 107 -266 209 -265
rect 212 -266 220 -265
rect 247 -266 283 -265
rect 289 -266 318 -265
rect 16 -268 104 -267
rect 152 -268 192 -267
rect 205 -268 241 -267
rect 250 -268 332 -267
rect 37 -270 202 -269
rect 215 -270 360 -269
rect 23 -272 216 -271
rect 233 -272 241 -271
rect 296 -272 339 -271
rect 44 -274 125 -273
rect 163 -274 178 -273
rect 191 -274 227 -273
rect 303 -274 318 -273
rect 51 -276 55 -275
rect 68 -276 83 -275
rect 86 -276 129 -275
rect 170 -276 220 -275
rect 303 -276 325 -275
rect 37 -278 52 -277
rect 72 -278 87 -277
rect 93 -278 160 -277
rect 170 -278 185 -277
rect 198 -278 227 -277
rect 268 -278 325 -277
rect 30 -280 199 -279
rect 201 -280 353 -279
rect 30 -282 136 -281
rect 205 -282 269 -281
rect 310 -282 339 -281
rect 44 -284 160 -283
rect 61 -286 311 -285
rect 72 -288 209 -287
rect 93 -290 115 -289
rect 100 -292 188 -291
rect 114 -294 143 -293
rect 142 -296 248 -295
rect 9 -307 62 -306
rect 68 -307 73 -306
rect 79 -307 90 -306
rect 107 -307 216 -306
rect 240 -307 318 -306
rect 373 -307 377 -306
rect 380 -307 388 -306
rect 9 -309 38 -308
rect 72 -309 87 -308
rect 110 -309 171 -308
rect 173 -309 192 -308
rect 198 -309 241 -308
rect 250 -309 339 -308
rect 2 -311 87 -310
rect 124 -311 150 -310
rect 152 -311 227 -310
rect 296 -311 300 -310
rect 310 -311 370 -310
rect 2 -313 157 -312
rect 159 -313 304 -312
rect 16 -315 167 -314
rect 187 -315 360 -314
rect 23 -317 125 -316
rect 128 -317 185 -316
rect 205 -317 325 -316
rect 345 -317 360 -316
rect 23 -319 83 -318
rect 93 -319 157 -318
rect 208 -319 353 -318
rect 30 -321 136 -320
rect 138 -321 234 -320
rect 236 -321 311 -320
rect 324 -321 332 -320
rect 338 -321 353 -320
rect 30 -323 143 -322
rect 145 -323 248 -322
rect 254 -323 332 -322
rect 37 -325 115 -324
rect 135 -325 244 -324
rect 268 -325 346 -324
rect 44 -327 143 -326
rect 159 -327 255 -326
rect 261 -327 269 -326
rect 275 -327 304 -326
rect 44 -329 52 -328
rect 93 -329 118 -328
rect 163 -329 262 -328
rect 275 -329 290 -328
rect 100 -331 129 -330
rect 163 -331 202 -330
rect 212 -331 318 -330
rect 65 -333 101 -332
rect 219 -333 227 -332
rect 282 -333 290 -332
rect 16 -335 66 -334
rect 114 -335 220 -334
rect 194 -337 283 -336
rect 2 -348 146 -347
rect 170 -348 367 -347
rect 397 -348 402 -347
rect 9 -350 45 -349
rect 61 -350 188 -349
rect 194 -350 290 -349
rect 331 -350 339 -349
rect 16 -352 97 -351
rect 110 -352 227 -351
rect 236 -352 269 -351
rect 282 -352 381 -351
rect 16 -354 73 -353
rect 86 -354 118 -353
rect 170 -354 374 -353
rect 23 -356 115 -355
rect 177 -356 192 -355
rect 198 -356 213 -355
rect 215 -356 234 -355
rect 240 -356 346 -355
rect 23 -358 101 -357
rect 114 -358 185 -357
rect 191 -358 258 -357
rect 285 -358 360 -357
rect 30 -360 160 -359
rect 163 -360 178 -359
rect 198 -360 244 -359
rect 247 -360 346 -359
rect 30 -362 66 -361
rect 68 -362 90 -361
rect 93 -362 122 -361
rect 128 -362 164 -361
rect 205 -362 290 -361
rect 296 -362 360 -361
rect 9 -364 90 -363
rect 100 -364 150 -363
rect 208 -364 332 -363
rect 37 -366 174 -365
rect 212 -366 318 -365
rect 37 -368 136 -367
rect 149 -368 353 -367
rect 58 -370 129 -369
rect 135 -370 153 -369
rect 219 -370 227 -369
rect 240 -370 318 -369
rect 72 -372 94 -371
rect 121 -372 146 -371
rect 219 -372 297 -371
rect 79 -374 206 -373
rect 222 -374 304 -373
rect 44 -376 80 -375
rect 173 -376 304 -375
rect 243 -378 311 -377
rect 247 -380 255 -379
rect 261 -380 311 -379
rect 159 -382 262 -381
rect 271 -382 353 -381
rect 9 -393 160 -392
rect 170 -393 206 -392
rect 240 -393 276 -392
rect 282 -393 325 -392
rect 387 -393 395 -392
rect 401 -393 412 -392
rect 16 -395 118 -394
rect 131 -395 174 -394
rect 184 -395 209 -394
rect 268 -395 311 -394
rect 324 -395 367 -394
rect 23 -397 150 -396
rect 156 -397 178 -396
rect 194 -397 199 -396
rect 201 -397 220 -396
rect 261 -397 269 -396
rect 296 -397 367 -396
rect 23 -399 94 -398
rect 110 -399 178 -398
rect 198 -399 227 -398
rect 250 -399 262 -398
rect 296 -399 381 -398
rect 37 -401 129 -400
rect 142 -401 248 -400
rect 310 -401 353 -400
rect 30 -403 38 -402
rect 65 -403 118 -402
rect 128 -403 136 -402
rect 149 -403 223 -402
rect 226 -403 258 -402
rect 331 -403 381 -402
rect 30 -405 52 -404
rect 65 -405 234 -404
rect 285 -405 332 -404
rect 338 -405 353 -404
rect 68 -407 276 -406
rect 72 -409 216 -408
rect 233 -409 304 -408
rect 72 -411 122 -410
rect 135 -411 171 -410
rect 247 -411 339 -410
rect 79 -413 90 -412
rect 107 -413 143 -412
rect 156 -413 220 -412
rect 303 -413 346 -412
rect 44 -415 80 -414
rect 86 -415 101 -414
rect 114 -415 286 -414
rect 317 -415 346 -414
rect 100 -417 146 -416
rect 163 -417 185 -416
rect 317 -417 360 -416
rect 121 -419 160 -418
rect 163 -419 213 -418
rect 289 -419 360 -418
rect 205 -421 290 -420
rect 23 -432 48 -431
rect 65 -432 101 -431
rect 107 -432 129 -431
rect 142 -432 146 -431
rect 159 -432 185 -431
rect 191 -432 234 -431
rect 240 -432 269 -431
rect 306 -432 311 -431
rect 313 -432 339 -431
rect 352 -432 374 -431
rect 30 -434 69 -433
rect 72 -434 132 -433
rect 142 -434 150 -433
rect 163 -434 213 -433
rect 215 -434 318 -433
rect 320 -434 346 -433
rect 352 -434 367 -433
rect 37 -436 125 -435
rect 145 -436 150 -435
rect 170 -436 188 -435
rect 215 -436 332 -435
rect 359 -436 381 -435
rect 44 -438 52 -437
rect 86 -438 97 -437
rect 114 -438 122 -437
rect 170 -438 185 -437
rect 226 -438 234 -437
rect 247 -438 304 -437
rect 362 -438 367 -437
rect 51 -440 213 -439
rect 229 -440 325 -439
rect 65 -442 87 -441
rect 93 -442 101 -441
rect 177 -442 206 -441
rect 254 -442 262 -441
rect 268 -442 276 -441
rect 303 -442 332 -441
rect 75 -444 115 -443
rect 117 -444 255 -443
rect 275 -444 290 -443
rect 93 -446 160 -445
rect 198 -446 262 -445
rect 289 -446 297 -445
rect 135 -448 178 -447
rect 191 -448 297 -447
rect 194 -450 199 -449
rect 205 -450 356 -449
rect 194 -452 220 -451
rect 156 -454 220 -453
rect 26 -465 111 -464
rect 121 -465 199 -464
rect 212 -465 227 -464
rect 250 -465 276 -464
rect 296 -465 325 -464
rect 338 -465 353 -464
rect 366 -465 377 -464
rect 33 -467 73 -466
rect 79 -467 115 -466
rect 121 -467 209 -466
rect 215 -467 241 -466
rect 254 -467 353 -466
rect 37 -469 115 -468
rect 142 -469 206 -468
rect 240 -469 290 -468
rect 317 -469 360 -468
rect 37 -471 118 -470
rect 149 -471 157 -470
rect 177 -471 227 -470
rect 261 -471 304 -470
rect 331 -471 360 -470
rect 44 -473 69 -472
rect 72 -473 87 -472
rect 93 -473 136 -472
rect 177 -473 220 -472
rect 275 -473 321 -472
rect 331 -473 349 -472
rect 44 -475 66 -474
rect 86 -475 129 -474
rect 135 -475 164 -474
rect 184 -475 230 -474
rect 282 -475 290 -474
rect 58 -477 80 -476
rect 107 -477 139 -476
rect 163 -477 171 -476
rect 187 -477 269 -476
rect 51 -479 59 -478
rect 128 -479 150 -478
rect 170 -479 262 -478
rect 51 -481 132 -480
rect 173 -481 269 -480
rect 100 -483 132 -482
rect 191 -483 234 -482
rect 100 -485 146 -484
rect 194 -485 255 -484
rect 198 -487 248 -486
rect 205 -489 244 -488
rect 233 -491 307 -490
rect 16 -502 108 -501
rect 156 -502 174 -501
rect 177 -502 195 -501
rect 201 -502 206 -501
rect 222 -502 300 -501
rect 338 -502 360 -501
rect 30 -504 45 -503
rect 51 -504 244 -503
rect 268 -504 314 -503
rect 345 -504 349 -503
rect 352 -504 374 -503
rect 65 -506 80 -505
rect 86 -506 94 -505
rect 110 -506 157 -505
rect 159 -506 227 -505
rect 275 -506 297 -505
rect 317 -506 349 -505
rect 51 -508 94 -507
rect 163 -508 199 -507
rect 226 -508 290 -507
rect 296 -508 332 -507
rect 341 -508 353 -507
rect 44 -510 199 -509
rect 208 -510 332 -509
rect 341 -510 367 -509
rect 65 -512 143 -511
rect 149 -512 164 -511
rect 166 -512 311 -511
rect 68 -514 111 -513
rect 170 -514 241 -513
rect 282 -514 325 -513
rect 72 -516 132 -515
rect 191 -516 220 -515
rect 233 -516 241 -515
rect 247 -516 283 -515
rect 289 -516 304 -515
rect 37 -518 73 -517
rect 79 -518 150 -517
rect 194 -518 248 -517
rect 261 -518 325 -517
rect 37 -520 59 -519
rect 86 -520 101 -519
rect 114 -520 220 -519
rect 229 -520 304 -519
rect 58 -522 122 -521
rect 142 -522 234 -521
rect 100 -524 269 -523
rect 114 -526 136 -525
rect 201 -526 262 -525
rect 135 -528 185 -527
rect 177 -530 185 -529
rect 9 -541 108 -540
rect 121 -541 150 -540
rect 156 -541 220 -540
rect 222 -541 332 -540
rect 338 -541 374 -540
rect 16 -543 230 -542
rect 275 -543 290 -542
rect 348 -543 353 -542
rect 16 -545 52 -544
rect 58 -545 167 -544
rect 177 -545 206 -544
rect 208 -545 290 -544
rect 23 -547 27 -546
rect 37 -547 83 -546
rect 86 -547 104 -546
rect 131 -547 346 -546
rect 44 -549 125 -548
rect 142 -549 206 -548
rect 226 -549 262 -548
rect 275 -549 367 -548
rect 30 -551 45 -550
rect 58 -551 80 -550
rect 86 -551 111 -550
rect 114 -551 132 -550
rect 145 -551 248 -550
rect 254 -551 262 -550
rect 65 -553 153 -552
rect 177 -553 237 -552
rect 247 -553 279 -552
rect 65 -555 160 -554
rect 191 -555 234 -554
rect 268 -555 279 -554
rect 72 -557 136 -556
rect 201 -557 283 -556
rect 93 -559 241 -558
rect 268 -559 325 -558
rect 93 -561 146 -560
rect 240 -561 304 -560
rect 317 -561 325 -560
rect 100 -563 199 -562
rect 282 -563 293 -562
rect 303 -563 311 -562
rect 100 -565 129 -564
rect 135 -565 153 -564
rect 198 -565 213 -564
rect 114 -567 125 -566
rect 170 -567 213 -566
rect 163 -569 171 -568
rect 9 -580 157 -579
rect 159 -580 199 -579
rect 205 -580 234 -579
rect 257 -580 262 -579
rect 282 -580 311 -579
rect 355 -580 360 -579
rect 16 -582 52 -581
rect 65 -582 97 -581
rect 100 -582 111 -581
rect 135 -582 143 -581
rect 187 -582 192 -581
rect 198 -582 220 -581
rect 226 -582 255 -581
rect 261 -582 269 -581
rect 282 -582 307 -581
rect 30 -584 83 -583
rect 86 -584 146 -583
rect 163 -584 192 -583
rect 205 -584 230 -583
rect 268 -584 279 -583
rect 289 -584 304 -583
rect 51 -586 132 -585
rect 135 -586 139 -585
rect 163 -586 185 -585
rect 219 -586 241 -585
rect 296 -586 304 -585
rect 58 -588 66 -587
rect 72 -588 153 -587
rect 177 -588 188 -587
rect 58 -590 101 -589
rect 152 -590 213 -589
rect 75 -592 129 -591
rect 170 -592 178 -591
rect 212 -592 248 -591
rect 86 -594 115 -593
rect 159 -594 248 -593
rect 93 -596 108 -595
rect 114 -596 122 -595
rect 79 -598 94 -597
rect 107 -598 150 -597
rect 33 -600 80 -599
rect 30 -611 83 -610
rect 100 -611 104 -610
rect 114 -611 129 -610
rect 131 -611 150 -610
rect 156 -611 181 -610
rect 184 -611 213 -610
rect 226 -611 255 -610
rect 257 -611 283 -610
rect 37 -613 45 -612
rect 51 -613 118 -612
rect 135 -613 192 -612
rect 205 -613 227 -612
rect 233 -613 265 -612
rect 275 -613 290 -612
rect 51 -615 73 -614
rect 86 -615 118 -614
rect 135 -615 143 -614
rect 159 -615 199 -614
rect 205 -615 220 -614
rect 233 -615 262 -614
rect 58 -617 139 -616
rect 142 -617 157 -616
rect 163 -617 174 -616
rect 177 -617 181 -616
rect 187 -617 213 -616
rect 240 -617 248 -616
rect 261 -617 269 -616
rect 65 -619 87 -618
rect 114 -619 146 -618
rect 152 -619 220 -618
rect 243 -619 248 -618
rect 65 -621 108 -620
rect 121 -621 164 -620
rect 170 -621 199 -620
rect 79 -623 122 -622
rect 191 -623 255 -622
rect 75 -625 80 -624
rect 93 -625 108 -624
rect 30 -636 52 -635
rect 65 -636 108 -635
rect 121 -636 150 -635
rect 152 -636 192 -635
rect 201 -636 269 -635
rect 37 -638 73 -637
rect 82 -638 101 -637
rect 107 -638 118 -637
rect 124 -638 164 -637
rect 184 -638 241 -637
rect 247 -638 290 -637
rect 44 -640 76 -639
rect 96 -640 234 -639
rect 254 -640 258 -639
rect 51 -642 94 -641
rect 100 -642 122 -641
rect 135 -642 146 -641
rect 149 -642 188 -641
rect 205 -642 234 -641
rect 68 -644 80 -643
rect 128 -644 136 -643
rect 142 -644 262 -643
rect 75 -646 87 -645
rect 128 -646 139 -645
rect 156 -646 174 -645
rect 187 -646 297 -645
rect 156 -648 164 -647
rect 170 -648 248 -647
rect 212 -650 241 -649
rect 198 -652 213 -651
rect 219 -652 283 -651
rect 219 -654 237 -653
rect 226 -656 276 -655
rect 191 -658 227 -657
rect 37 -669 111 -668
rect 114 -669 143 -668
rect 156 -669 227 -668
rect 254 -669 279 -668
rect 44 -671 146 -670
rect 156 -671 164 -670
rect 173 -671 269 -670
rect 51 -673 118 -672
rect 121 -673 192 -672
rect 198 -673 213 -672
rect 247 -673 255 -672
rect 261 -673 269 -672
rect 58 -675 87 -674
rect 89 -675 139 -674
rect 159 -675 202 -674
rect 208 -675 276 -674
rect 61 -677 69 -676
rect 93 -677 185 -676
rect 187 -677 234 -676
rect 30 -679 62 -678
rect 93 -679 150 -678
rect 180 -679 283 -678
rect 96 -681 101 -680
rect 138 -681 164 -680
rect 180 -681 290 -680
rect 100 -683 108 -682
rect 191 -683 227 -682
rect 107 -685 171 -684
rect 212 -685 241 -684
rect 177 -687 241 -686
rect 219 -689 234 -688
rect 177 -691 220 -690
rect 61 -702 73 -701
rect 75 -702 80 -701
rect 100 -702 118 -701
rect 121 -702 178 -701
rect 184 -702 227 -701
rect 240 -702 262 -701
rect 114 -704 122 -703
rect 128 -704 136 -703
rect 142 -704 188 -703
rect 194 -704 199 -703
rect 240 -704 255 -703
rect 131 -706 143 -705
rect 149 -706 171 -705
rect 194 -706 220 -705
rect 247 -706 269 -705
rect 93 -708 171 -707
rect 198 -708 234 -707
rect 152 -710 206 -709
rect 163 -712 174 -711
rect 205 -712 216 -711
rect 163 -714 181 -713
rect 114 -725 132 -724
rect 135 -725 143 -724
rect 159 -725 178 -724
rect 180 -725 185 -724
rect 191 -725 206 -724
rect 229 -725 241 -724
rect 121 -727 132 -726
rect 163 -727 171 -726
rect 173 -727 199 -726
rect 117 -729 122 -728
rect 177 -729 185 -728
rect 191 -729 195 -728
rect 128 -740 136 -739
rect 149 -740 164 -739
rect 166 -740 171 -739
rect 177 -740 185 -739
rect 187 -740 192 -739
rect 121 -742 129 -741
rect 156 -742 171 -741
rect 124 -753 129 -752
rect 156 -753 171 -752
rect 184 -753 192 -752
rect 159 -755 164 -754
<< m2contact >>
rect 103 0 104 1
rect 107 0 108 1
rect 128 0 129 1
rect 135 0 136 1
rect 142 0 143 1
rect 156 0 157 1
rect 177 0 178 1
rect 191 0 192 1
rect 194 0 195 1
rect 212 0 213 1
rect 198 -2 199 -1
rect 205 -2 206 -1
rect 79 -13 80 -12
rect 96 -13 97 -12
rect 100 -13 101 -12
rect 103 -13 104 -12
rect 110 -13 111 -12
rect 121 -13 122 -12
rect 135 -13 136 -12
rect 142 -13 143 -12
rect 149 -13 150 -12
rect 156 -13 157 -12
rect 170 -13 171 -12
rect 194 -13 195 -12
rect 208 -13 209 -12
rect 233 -13 234 -12
rect 135 -15 136 -14
rect 156 -15 157 -14
rect 177 -15 178 -14
rect 184 -15 185 -14
rect 212 -15 213 -14
rect 226 -15 227 -14
rect 142 -17 143 -16
rect 173 -17 174 -16
rect 184 -17 185 -16
rect 198 -17 199 -16
rect 215 -17 216 -16
rect 219 -17 220 -16
rect 149 -19 150 -18
rect 163 -19 164 -18
rect 152 -21 153 -20
rect 198 -21 199 -20
rect 65 -32 66 -31
rect 89 -32 90 -31
rect 93 -32 94 -31
rect 96 -32 97 -31
rect 114 -32 115 -31
rect 173 -32 174 -31
rect 184 -32 185 -31
rect 247 -32 248 -31
rect 271 -32 272 -31
rect 275 -32 276 -31
rect 72 -34 73 -33
rect 110 -34 111 -33
rect 142 -34 143 -33
rect 187 -34 188 -33
rect 198 -34 199 -33
rect 226 -34 227 -33
rect 229 -34 230 -33
rect 282 -34 283 -33
rect 86 -36 87 -35
rect 89 -36 90 -35
rect 93 -36 94 -35
rect 100 -36 101 -35
rect 149 -36 150 -35
rect 170 -36 171 -35
rect 180 -36 181 -35
rect 184 -36 185 -35
rect 201 -36 202 -35
rect 254 -36 255 -35
rect 86 -38 87 -37
rect 107 -38 108 -37
rect 135 -38 136 -37
rect 149 -38 150 -37
rect 152 -38 153 -37
rect 240 -38 241 -37
rect 96 -40 97 -39
rect 100 -40 101 -39
rect 121 -40 122 -39
rect 135 -40 136 -39
rect 156 -40 157 -39
rect 163 -40 164 -39
rect 215 -40 216 -39
rect 219 -40 220 -39
rect 233 -40 234 -39
rect 261 -40 262 -39
rect 156 -42 157 -41
rect 170 -42 171 -41
rect 191 -42 192 -41
rect 233 -42 234 -41
rect 159 -44 160 -43
rect 166 -44 167 -43
rect 177 -44 178 -43
rect 191 -44 192 -43
rect 205 -44 206 -43
rect 219 -44 220 -43
rect 30 -55 31 -54
rect 75 -55 76 -54
rect 82 -55 83 -54
rect 145 -55 146 -54
rect 170 -55 171 -54
rect 261 -55 262 -54
rect 44 -57 45 -56
rect 114 -57 115 -56
rect 117 -57 118 -56
rect 149 -57 150 -56
rect 163 -57 164 -56
rect 170 -57 171 -56
rect 184 -57 185 -56
rect 261 -57 262 -56
rect 51 -59 52 -58
rect 131 -59 132 -58
rect 159 -59 160 -58
rect 163 -59 164 -58
rect 187 -59 188 -58
rect 289 -59 290 -58
rect 58 -61 59 -60
rect 156 -61 157 -60
rect 191 -61 192 -60
rect 198 -61 199 -60
rect 201 -61 202 -60
rect 240 -61 241 -60
rect 243 -61 244 -60
rect 303 -61 304 -60
rect 61 -63 62 -62
rect 89 -63 90 -62
rect 93 -63 94 -62
rect 177 -63 178 -62
rect 198 -63 199 -62
rect 226 -63 227 -62
rect 233 -63 234 -62
rect 268 -63 269 -62
rect 65 -65 66 -64
rect 86 -65 87 -64
rect 100 -65 101 -64
rect 114 -65 115 -64
rect 121 -65 122 -64
rect 135 -65 136 -64
rect 142 -65 143 -64
rect 191 -65 192 -64
rect 219 -65 220 -64
rect 275 -65 276 -64
rect 65 -67 66 -66
rect 96 -67 97 -66
rect 100 -67 101 -66
rect 138 -67 139 -66
rect 180 -67 181 -66
rect 226 -67 227 -66
rect 254 -67 255 -66
rect 275 -67 276 -66
rect 72 -69 73 -68
rect 135 -69 136 -68
rect 184 -69 185 -68
rect 233 -69 234 -68
rect 72 -71 73 -70
rect 79 -71 80 -70
rect 103 -71 104 -70
rect 142 -71 143 -70
rect 212 -71 213 -70
rect 254 -71 255 -70
rect 110 -73 111 -72
rect 124 -73 125 -72
rect 205 -73 206 -72
rect 212 -73 213 -72
rect 222 -73 223 -72
rect 282 -73 283 -72
rect 121 -75 122 -74
rect 156 -75 157 -74
rect 247 -75 248 -74
rect 282 -75 283 -74
rect 16 -86 17 -85
rect 79 -86 80 -85
rect 86 -86 87 -85
rect 100 -86 101 -85
rect 103 -86 104 -85
rect 107 -86 108 -85
rect 114 -86 115 -85
rect 135 -86 136 -85
rect 170 -86 171 -85
rect 180 -86 181 -85
rect 184 -86 185 -85
rect 194 -86 195 -85
rect 201 -86 202 -85
rect 236 -86 237 -85
rect 243 -86 244 -85
rect 282 -86 283 -85
rect 299 -86 300 -85
rect 331 -86 332 -85
rect 30 -88 31 -87
rect 324 -88 325 -87
rect 26 -90 27 -89
rect 30 -90 31 -89
rect 37 -90 38 -89
rect 79 -90 80 -89
rect 100 -90 101 -89
rect 208 -90 209 -89
rect 250 -90 251 -89
rect 289 -90 290 -89
rect 37 -92 38 -91
rect 93 -92 94 -91
rect 107 -92 108 -91
rect 124 -92 125 -91
rect 131 -92 132 -91
rect 226 -92 227 -91
rect 268 -92 269 -91
rect 310 -92 311 -91
rect 44 -94 45 -93
rect 110 -94 111 -93
rect 138 -94 139 -93
rect 282 -94 283 -93
rect 51 -96 52 -95
rect 187 -96 188 -95
rect 191 -96 192 -95
rect 240 -96 241 -95
rect 275 -96 276 -95
rect 317 -96 318 -95
rect 58 -98 59 -97
rect 128 -98 129 -97
rect 142 -98 143 -97
rect 289 -98 290 -97
rect 65 -100 66 -99
rect 86 -100 87 -99
rect 93 -100 94 -99
rect 138 -100 139 -99
rect 163 -100 164 -99
rect 170 -100 171 -99
rect 177 -100 178 -99
rect 261 -100 262 -99
rect 51 -102 52 -101
rect 65 -102 66 -101
rect 68 -102 69 -101
rect 159 -102 160 -101
rect 180 -102 181 -101
rect 212 -102 213 -101
rect 219 -102 220 -101
rect 226 -102 227 -101
rect 72 -104 73 -103
rect 117 -104 118 -103
rect 128 -104 129 -103
rect 152 -104 153 -103
rect 187 -104 188 -103
rect 261 -104 262 -103
rect 117 -106 118 -105
rect 268 -106 269 -105
rect 198 -108 199 -107
rect 275 -108 276 -107
rect 198 -110 199 -109
rect 303 -110 304 -109
rect 149 -112 150 -111
rect 303 -112 304 -111
rect 121 -114 122 -113
rect 149 -114 150 -113
rect 201 -114 202 -113
rect 233 -114 234 -113
rect 205 -116 206 -115
rect 296 -116 297 -115
rect 205 -118 206 -117
rect 247 -118 248 -117
rect 208 -120 209 -119
rect 219 -120 220 -119
rect 23 -131 24 -130
rect 145 -131 146 -130
rect 159 -131 160 -130
rect 240 -131 241 -130
rect 26 -133 27 -132
rect 30 -133 31 -132
rect 37 -133 38 -132
rect 180 -133 181 -132
rect 198 -133 199 -132
rect 247 -133 248 -132
rect 23 -135 24 -134
rect 30 -135 31 -134
rect 44 -135 45 -134
rect 51 -135 52 -134
rect 61 -135 62 -134
rect 89 -135 90 -134
rect 100 -135 101 -134
rect 282 -135 283 -134
rect 37 -137 38 -136
rect 61 -137 62 -136
rect 65 -137 66 -136
rect 324 -137 325 -136
rect 47 -139 48 -138
rect 65 -139 66 -138
rect 72 -139 73 -138
rect 82 -139 83 -138
rect 86 -139 87 -138
rect 117 -139 118 -138
rect 128 -139 129 -138
rect 243 -139 244 -138
rect 72 -141 73 -140
rect 93 -141 94 -140
rect 100 -141 101 -140
rect 107 -141 108 -140
rect 110 -141 111 -140
rect 114 -141 115 -140
rect 117 -141 118 -140
rect 124 -141 125 -140
rect 128 -141 129 -140
rect 152 -141 153 -140
rect 166 -141 167 -140
rect 194 -141 195 -140
rect 205 -141 206 -140
rect 268 -141 269 -140
rect 16 -143 17 -142
rect 114 -143 115 -142
rect 135 -143 136 -142
rect 289 -143 290 -142
rect 79 -145 80 -144
rect 93 -145 94 -144
rect 142 -145 143 -144
rect 303 -145 304 -144
rect 79 -147 80 -146
rect 152 -147 153 -146
rect 170 -147 171 -146
rect 184 -147 185 -146
rect 205 -147 206 -146
rect 310 -147 311 -146
rect 131 -149 132 -148
rect 170 -149 171 -148
rect 177 -149 178 -148
rect 187 -149 188 -148
rect 201 -149 202 -148
rect 310 -149 311 -148
rect 103 -151 104 -150
rect 177 -151 178 -150
rect 201 -151 202 -150
rect 289 -151 290 -150
rect 303 -151 304 -150
rect 331 -151 332 -150
rect 142 -153 143 -152
rect 159 -153 160 -152
rect 215 -153 216 -152
rect 296 -153 297 -152
rect 156 -155 157 -154
rect 184 -155 185 -154
rect 226 -155 227 -154
rect 229 -155 230 -154
rect 233 -155 234 -154
rect 296 -155 297 -154
rect 212 -157 213 -156
rect 233 -157 234 -156
rect 236 -157 237 -156
rect 317 -157 318 -156
rect 212 -159 213 -158
rect 247 -159 248 -158
rect 226 -161 227 -160
rect 261 -161 262 -160
rect 236 -163 237 -162
rect 282 -163 283 -162
rect 254 -165 255 -164
rect 261 -165 262 -164
rect 229 -167 230 -166
rect 254 -167 255 -166
rect 16 -178 17 -177
rect 33 -178 34 -177
rect 37 -178 38 -177
rect 68 -178 69 -177
rect 72 -178 73 -177
rect 86 -178 87 -177
rect 89 -178 90 -177
rect 110 -178 111 -177
rect 121 -178 122 -177
rect 128 -178 129 -177
rect 135 -178 136 -177
rect 142 -178 143 -177
rect 145 -178 146 -177
rect 394 -178 395 -177
rect 9 -180 10 -179
rect 86 -180 87 -179
rect 149 -180 150 -179
rect 198 -180 199 -179
rect 222 -180 223 -179
rect 296 -180 297 -179
rect 303 -180 304 -179
rect 359 -180 360 -179
rect 19 -182 20 -181
rect 58 -182 59 -181
rect 72 -182 73 -181
rect 135 -182 136 -181
rect 149 -182 150 -181
rect 184 -182 185 -181
rect 191 -182 192 -181
rect 215 -182 216 -181
rect 240 -182 241 -181
rect 261 -182 262 -181
rect 268 -182 269 -181
rect 331 -182 332 -181
rect 23 -184 24 -183
rect 30 -184 31 -183
rect 44 -184 45 -183
rect 51 -184 52 -183
rect 54 -184 55 -183
rect 58 -184 59 -183
rect 79 -184 80 -183
rect 107 -184 108 -183
rect 117 -184 118 -183
rect 240 -184 241 -183
rect 243 -184 244 -183
rect 324 -184 325 -183
rect 44 -186 45 -185
rect 184 -186 185 -185
rect 194 -186 195 -185
rect 226 -186 227 -185
rect 247 -186 248 -185
rect 261 -186 262 -185
rect 271 -186 272 -185
rect 303 -186 304 -185
rect 310 -186 311 -185
rect 373 -186 374 -185
rect 51 -188 52 -187
rect 93 -188 94 -187
rect 107 -188 108 -187
rect 236 -188 237 -187
rect 247 -188 248 -187
rect 387 -188 388 -187
rect 65 -190 66 -189
rect 79 -190 80 -189
rect 93 -190 94 -189
rect 205 -190 206 -189
rect 212 -190 213 -189
rect 310 -190 311 -189
rect 117 -192 118 -191
rect 124 -192 125 -191
rect 156 -192 157 -191
rect 163 -192 164 -191
rect 170 -192 171 -191
rect 205 -192 206 -191
rect 275 -192 276 -191
rect 296 -192 297 -191
rect 114 -194 115 -193
rect 275 -194 276 -193
rect 282 -194 283 -193
rect 338 -194 339 -193
rect 128 -196 129 -195
rect 156 -196 157 -195
rect 159 -196 160 -195
rect 219 -196 220 -195
rect 285 -196 286 -195
rect 352 -196 353 -195
rect 170 -198 171 -197
rect 208 -198 209 -197
rect 219 -198 220 -197
rect 380 -198 381 -197
rect 177 -200 178 -199
rect 226 -200 227 -199
rect 289 -200 290 -199
rect 345 -200 346 -199
rect 177 -202 178 -201
rect 254 -202 255 -201
rect 289 -202 290 -201
rect 317 -202 318 -201
rect 201 -204 202 -203
rect 254 -204 255 -203
rect 292 -204 293 -203
rect 366 -204 367 -203
rect 9 -215 10 -214
rect 142 -215 143 -214
rect 149 -215 150 -214
rect 184 -215 185 -214
rect 187 -215 188 -214
rect 345 -215 346 -214
rect 9 -217 10 -216
rect 75 -217 76 -216
rect 86 -217 87 -216
rect 100 -217 101 -216
rect 114 -217 115 -216
rect 135 -217 136 -216
rect 156 -217 157 -216
rect 170 -217 171 -216
rect 177 -217 178 -216
rect 215 -217 216 -216
rect 222 -217 223 -216
rect 373 -217 374 -216
rect 16 -219 17 -218
rect 54 -219 55 -218
rect 72 -219 73 -218
rect 79 -219 80 -218
rect 93 -219 94 -218
rect 159 -219 160 -218
rect 163 -219 164 -218
rect 233 -219 234 -218
rect 261 -219 262 -218
rect 282 -219 283 -218
rect 289 -219 290 -218
rect 324 -219 325 -218
rect 16 -221 17 -220
rect 124 -221 125 -220
rect 128 -221 129 -220
rect 142 -221 143 -220
rect 170 -221 171 -220
rect 219 -221 220 -220
rect 229 -221 230 -220
rect 359 -221 360 -220
rect 26 -223 27 -222
rect 110 -223 111 -222
rect 117 -223 118 -222
rect 380 -223 381 -222
rect 30 -225 31 -224
rect 191 -225 192 -224
rect 215 -225 216 -224
rect 296 -225 297 -224
rect 366 -225 367 -224
rect 380 -225 381 -224
rect 37 -227 38 -226
rect 163 -227 164 -226
rect 191 -227 192 -226
rect 254 -227 255 -226
rect 268 -227 269 -226
rect 338 -227 339 -226
rect 37 -229 38 -228
rect 121 -229 122 -228
rect 128 -229 129 -228
rect 212 -229 213 -228
rect 219 -229 220 -228
rect 226 -229 227 -228
rect 233 -229 234 -228
rect 247 -229 248 -228
rect 254 -229 255 -228
rect 285 -229 286 -228
rect 292 -229 293 -228
rect 345 -229 346 -228
rect 44 -231 45 -230
rect 177 -231 178 -230
rect 198 -231 199 -230
rect 268 -231 269 -230
rect 296 -231 297 -230
rect 303 -231 304 -230
rect 44 -233 45 -232
rect 82 -233 83 -232
rect 89 -233 90 -232
rect 359 -233 360 -232
rect 51 -235 52 -234
rect 58 -235 59 -234
rect 72 -235 73 -234
rect 79 -235 80 -234
rect 93 -235 94 -234
rect 110 -235 111 -234
rect 114 -235 115 -234
rect 226 -235 227 -234
rect 240 -235 241 -234
rect 324 -235 325 -234
rect 58 -237 59 -236
rect 152 -237 153 -236
rect 156 -237 157 -236
rect 247 -237 248 -236
rect 303 -237 304 -236
rect 310 -237 311 -236
rect 121 -239 122 -238
rect 394 -239 395 -238
rect 198 -241 199 -240
rect 331 -241 332 -240
rect 208 -243 209 -242
rect 338 -243 339 -242
rect 208 -245 209 -244
rect 275 -245 276 -244
rect 310 -245 311 -244
rect 317 -245 318 -244
rect 331 -245 332 -244
rect 373 -245 374 -244
rect 201 -247 202 -246
rect 317 -247 318 -246
rect 240 -249 241 -248
rect 275 -249 276 -248
rect 2 -260 3 -259
rect 124 -260 125 -259
rect 138 -260 139 -259
rect 254 -260 255 -259
rect 264 -260 265 -259
rect 296 -260 297 -259
rect 359 -260 360 -259
rect 369 -260 370 -259
rect 376 -260 377 -259
rect 380 -260 381 -259
rect 9 -262 10 -261
rect 75 -262 76 -261
rect 79 -262 80 -261
rect 107 -262 108 -261
rect 121 -262 122 -261
rect 156 -262 157 -261
rect 166 -262 167 -261
rect 261 -262 262 -261
rect 275 -262 276 -261
rect 331 -262 332 -261
rect 366 -262 367 -261
rect 369 -262 370 -261
rect 9 -264 10 -263
rect 58 -264 59 -263
rect 65 -264 66 -263
rect 128 -264 129 -263
rect 149 -264 150 -263
rect 177 -264 178 -263
rect 184 -264 185 -263
rect 257 -264 258 -263
rect 275 -264 276 -263
rect 282 -264 283 -263
rect 289 -264 290 -263
rect 352 -264 353 -263
rect 366 -264 367 -263
rect 380 -264 381 -263
rect 16 -266 17 -265
rect 100 -266 101 -265
rect 107 -266 108 -265
rect 208 -266 209 -265
rect 212 -266 213 -265
rect 219 -266 220 -265
rect 247 -266 248 -265
rect 282 -266 283 -265
rect 289 -266 290 -265
rect 317 -266 318 -265
rect 16 -268 17 -267
rect 103 -268 104 -267
rect 152 -268 153 -267
rect 191 -268 192 -267
rect 205 -268 206 -267
rect 240 -268 241 -267
rect 250 -268 251 -267
rect 331 -268 332 -267
rect 37 -270 38 -269
rect 201 -270 202 -269
rect 215 -270 216 -269
rect 359 -270 360 -269
rect 23 -272 24 -271
rect 215 -272 216 -271
rect 233 -272 234 -271
rect 240 -272 241 -271
rect 296 -272 297 -271
rect 338 -272 339 -271
rect 44 -274 45 -273
rect 124 -274 125 -273
rect 163 -274 164 -273
rect 177 -274 178 -273
rect 191 -274 192 -273
rect 226 -274 227 -273
rect 303 -274 304 -273
rect 317 -274 318 -273
rect 51 -276 52 -275
rect 54 -276 55 -275
rect 68 -276 69 -275
rect 82 -276 83 -275
rect 86 -276 87 -275
rect 128 -276 129 -275
rect 170 -276 171 -275
rect 219 -276 220 -275
rect 303 -276 304 -275
rect 324 -276 325 -275
rect 37 -278 38 -277
rect 51 -278 52 -277
rect 72 -278 73 -277
rect 86 -278 87 -277
rect 93 -278 94 -277
rect 159 -278 160 -277
rect 170 -278 171 -277
rect 184 -278 185 -277
rect 198 -278 199 -277
rect 226 -278 227 -277
rect 268 -278 269 -277
rect 324 -278 325 -277
rect 30 -280 31 -279
rect 198 -280 199 -279
rect 201 -280 202 -279
rect 352 -280 353 -279
rect 30 -282 31 -281
rect 135 -282 136 -281
rect 205 -282 206 -281
rect 268 -282 269 -281
rect 310 -282 311 -281
rect 338 -282 339 -281
rect 44 -284 45 -283
rect 159 -284 160 -283
rect 61 -286 62 -285
rect 310 -286 311 -285
rect 72 -288 73 -287
rect 208 -288 209 -287
rect 93 -290 94 -289
rect 114 -290 115 -289
rect 100 -292 101 -291
rect 187 -292 188 -291
rect 114 -294 115 -293
rect 142 -294 143 -293
rect 142 -296 143 -295
rect 247 -296 248 -295
rect 9 -307 10 -306
rect 61 -307 62 -306
rect 68 -307 69 -306
rect 72 -307 73 -306
rect 79 -307 80 -306
rect 89 -307 90 -306
rect 107 -307 108 -306
rect 215 -307 216 -306
rect 240 -307 241 -306
rect 317 -307 318 -306
rect 373 -307 374 -306
rect 376 -307 377 -306
rect 380 -307 381 -306
rect 387 -307 388 -306
rect 9 -309 10 -308
rect 37 -309 38 -308
rect 72 -309 73 -308
rect 86 -309 87 -308
rect 110 -309 111 -308
rect 170 -309 171 -308
rect 173 -309 174 -308
rect 191 -309 192 -308
rect 198 -309 199 -308
rect 240 -309 241 -308
rect 250 -309 251 -308
rect 338 -309 339 -308
rect 2 -311 3 -310
rect 86 -311 87 -310
rect 124 -311 125 -310
rect 149 -311 150 -310
rect 152 -311 153 -310
rect 226 -311 227 -310
rect 296 -311 297 -310
rect 299 -311 300 -310
rect 310 -311 311 -310
rect 369 -311 370 -310
rect 2 -313 3 -312
rect 156 -313 157 -312
rect 159 -313 160 -312
rect 303 -313 304 -312
rect 16 -315 17 -314
rect 166 -315 167 -314
rect 187 -315 188 -314
rect 359 -315 360 -314
rect 23 -317 24 -316
rect 124 -317 125 -316
rect 128 -317 129 -316
rect 184 -317 185 -316
rect 205 -317 206 -316
rect 324 -317 325 -316
rect 345 -317 346 -316
rect 359 -317 360 -316
rect 23 -319 24 -318
rect 82 -319 83 -318
rect 93 -319 94 -318
rect 156 -319 157 -318
rect 208 -319 209 -318
rect 352 -319 353 -318
rect 30 -321 31 -320
rect 135 -321 136 -320
rect 138 -321 139 -320
rect 233 -321 234 -320
rect 236 -321 237 -320
rect 310 -321 311 -320
rect 324 -321 325 -320
rect 331 -321 332 -320
rect 338 -321 339 -320
rect 352 -321 353 -320
rect 30 -323 31 -322
rect 142 -323 143 -322
rect 145 -323 146 -322
rect 247 -323 248 -322
rect 254 -323 255 -322
rect 331 -323 332 -322
rect 37 -325 38 -324
rect 114 -325 115 -324
rect 135 -325 136 -324
rect 243 -325 244 -324
rect 268 -325 269 -324
rect 345 -325 346 -324
rect 44 -327 45 -326
rect 142 -327 143 -326
rect 159 -327 160 -326
rect 254 -327 255 -326
rect 261 -327 262 -326
rect 268 -327 269 -326
rect 275 -327 276 -326
rect 303 -327 304 -326
rect 44 -329 45 -328
rect 51 -329 52 -328
rect 93 -329 94 -328
rect 117 -329 118 -328
rect 163 -329 164 -328
rect 261 -329 262 -328
rect 275 -329 276 -328
rect 289 -329 290 -328
rect 100 -331 101 -330
rect 128 -331 129 -330
rect 163 -331 164 -330
rect 201 -331 202 -330
rect 212 -331 213 -330
rect 317 -331 318 -330
rect 65 -333 66 -332
rect 100 -333 101 -332
rect 219 -333 220 -332
rect 226 -333 227 -332
rect 282 -333 283 -332
rect 289 -333 290 -332
rect 16 -335 17 -334
rect 65 -335 66 -334
rect 114 -335 115 -334
rect 219 -335 220 -334
rect 194 -337 195 -336
rect 282 -337 283 -336
rect 2 -348 3 -347
rect 145 -348 146 -347
rect 170 -348 171 -347
rect 366 -348 367 -347
rect 397 -348 398 -347
rect 401 -348 402 -347
rect 9 -350 10 -349
rect 44 -350 45 -349
rect 61 -350 62 -349
rect 187 -350 188 -349
rect 194 -350 195 -349
rect 289 -350 290 -349
rect 331 -350 332 -349
rect 338 -350 339 -349
rect 16 -352 17 -351
rect 96 -352 97 -351
rect 110 -352 111 -351
rect 226 -352 227 -351
rect 236 -352 237 -351
rect 268 -352 269 -351
rect 282 -352 283 -351
rect 380 -352 381 -351
rect 16 -354 17 -353
rect 72 -354 73 -353
rect 86 -354 87 -353
rect 117 -354 118 -353
rect 170 -354 171 -353
rect 373 -354 374 -353
rect 23 -356 24 -355
rect 114 -356 115 -355
rect 177 -356 178 -355
rect 191 -356 192 -355
rect 198 -356 199 -355
rect 212 -356 213 -355
rect 215 -356 216 -355
rect 233 -356 234 -355
rect 240 -356 241 -355
rect 345 -356 346 -355
rect 23 -358 24 -357
rect 100 -358 101 -357
rect 114 -358 115 -357
rect 184 -358 185 -357
rect 191 -358 192 -357
rect 257 -358 258 -357
rect 285 -358 286 -357
rect 359 -358 360 -357
rect 30 -360 31 -359
rect 159 -360 160 -359
rect 163 -360 164 -359
rect 177 -360 178 -359
rect 198 -360 199 -359
rect 243 -360 244 -359
rect 247 -360 248 -359
rect 345 -360 346 -359
rect 30 -362 31 -361
rect 65 -362 66 -361
rect 68 -362 69 -361
rect 89 -362 90 -361
rect 93 -362 94 -361
rect 121 -362 122 -361
rect 128 -362 129 -361
rect 163 -362 164 -361
rect 205 -362 206 -361
rect 289 -362 290 -361
rect 296 -362 297 -361
rect 359 -362 360 -361
rect 9 -364 10 -363
rect 89 -364 90 -363
rect 100 -364 101 -363
rect 149 -364 150 -363
rect 208 -364 209 -363
rect 331 -364 332 -363
rect 37 -366 38 -365
rect 173 -366 174 -365
rect 212 -366 213 -365
rect 317 -366 318 -365
rect 37 -368 38 -367
rect 135 -368 136 -367
rect 149 -368 150 -367
rect 352 -368 353 -367
rect 58 -370 59 -369
rect 128 -370 129 -369
rect 135 -370 136 -369
rect 152 -370 153 -369
rect 219 -370 220 -369
rect 226 -370 227 -369
rect 240 -370 241 -369
rect 317 -370 318 -369
rect 72 -372 73 -371
rect 93 -372 94 -371
rect 121 -372 122 -371
rect 145 -372 146 -371
rect 219 -372 220 -371
rect 296 -372 297 -371
rect 79 -374 80 -373
rect 205 -374 206 -373
rect 222 -374 223 -373
rect 303 -374 304 -373
rect 44 -376 45 -375
rect 79 -376 80 -375
rect 173 -376 174 -375
rect 303 -376 304 -375
rect 243 -378 244 -377
rect 310 -378 311 -377
rect 247 -380 248 -379
rect 254 -380 255 -379
rect 261 -380 262 -379
rect 310 -380 311 -379
rect 159 -382 160 -381
rect 261 -382 262 -381
rect 271 -382 272 -381
rect 352 -382 353 -381
rect 9 -393 10 -392
rect 159 -393 160 -392
rect 170 -393 171 -392
rect 205 -393 206 -392
rect 240 -393 241 -392
rect 275 -393 276 -392
rect 282 -393 283 -392
rect 324 -393 325 -392
rect 387 -393 388 -392
rect 394 -393 395 -392
rect 401 -393 402 -392
rect 411 -393 412 -392
rect 16 -395 17 -394
rect 117 -395 118 -394
rect 131 -395 132 -394
rect 173 -395 174 -394
rect 184 -395 185 -394
rect 208 -395 209 -394
rect 268 -395 269 -394
rect 310 -395 311 -394
rect 324 -395 325 -394
rect 366 -395 367 -394
rect 23 -397 24 -396
rect 149 -397 150 -396
rect 156 -397 157 -396
rect 177 -397 178 -396
rect 194 -397 195 -396
rect 198 -397 199 -396
rect 201 -397 202 -396
rect 219 -397 220 -396
rect 261 -397 262 -396
rect 268 -397 269 -396
rect 296 -397 297 -396
rect 366 -397 367 -396
rect 23 -399 24 -398
rect 93 -399 94 -398
rect 110 -399 111 -398
rect 177 -399 178 -398
rect 198 -399 199 -398
rect 226 -399 227 -398
rect 250 -399 251 -398
rect 261 -399 262 -398
rect 296 -399 297 -398
rect 380 -399 381 -398
rect 37 -401 38 -400
rect 128 -401 129 -400
rect 142 -401 143 -400
rect 247 -401 248 -400
rect 310 -401 311 -400
rect 352 -401 353 -400
rect 30 -403 31 -402
rect 37 -403 38 -402
rect 65 -403 66 -402
rect 117 -403 118 -402
rect 128 -403 129 -402
rect 135 -403 136 -402
rect 149 -403 150 -402
rect 222 -403 223 -402
rect 226 -403 227 -402
rect 257 -403 258 -402
rect 331 -403 332 -402
rect 380 -403 381 -402
rect 30 -405 31 -404
rect 51 -405 52 -404
rect 65 -405 66 -404
rect 233 -405 234 -404
rect 285 -405 286 -404
rect 331 -405 332 -404
rect 338 -405 339 -404
rect 352 -405 353 -404
rect 68 -407 69 -406
rect 275 -407 276 -406
rect 72 -409 73 -408
rect 215 -409 216 -408
rect 233 -409 234 -408
rect 303 -409 304 -408
rect 72 -411 73 -410
rect 121 -411 122 -410
rect 135 -411 136 -410
rect 170 -411 171 -410
rect 247 -411 248 -410
rect 338 -411 339 -410
rect 79 -413 80 -412
rect 89 -413 90 -412
rect 107 -413 108 -412
rect 142 -413 143 -412
rect 156 -413 157 -412
rect 219 -413 220 -412
rect 303 -413 304 -412
rect 345 -413 346 -412
rect 44 -415 45 -414
rect 79 -415 80 -414
rect 86 -415 87 -414
rect 100 -415 101 -414
rect 114 -415 115 -414
rect 285 -415 286 -414
rect 317 -415 318 -414
rect 345 -415 346 -414
rect 100 -417 101 -416
rect 145 -417 146 -416
rect 163 -417 164 -416
rect 184 -417 185 -416
rect 317 -417 318 -416
rect 359 -417 360 -416
rect 121 -419 122 -418
rect 159 -419 160 -418
rect 163 -419 164 -418
rect 212 -419 213 -418
rect 289 -419 290 -418
rect 359 -419 360 -418
rect 205 -421 206 -420
rect 289 -421 290 -420
rect 23 -432 24 -431
rect 47 -432 48 -431
rect 65 -432 66 -431
rect 100 -432 101 -431
rect 107 -432 108 -431
rect 128 -432 129 -431
rect 142 -432 143 -431
rect 145 -432 146 -431
rect 159 -432 160 -431
rect 184 -432 185 -431
rect 191 -432 192 -431
rect 233 -432 234 -431
rect 240 -432 241 -431
rect 268 -432 269 -431
rect 306 -432 307 -431
rect 310 -432 311 -431
rect 313 -432 314 -431
rect 338 -432 339 -431
rect 352 -432 353 -431
rect 373 -432 374 -431
rect 30 -434 31 -433
rect 68 -434 69 -433
rect 72 -434 73 -433
rect 131 -434 132 -433
rect 142 -434 143 -433
rect 149 -434 150 -433
rect 163 -434 164 -433
rect 212 -434 213 -433
rect 215 -434 216 -433
rect 317 -434 318 -433
rect 320 -434 321 -433
rect 345 -434 346 -433
rect 352 -434 353 -433
rect 366 -434 367 -433
rect 37 -436 38 -435
rect 124 -436 125 -435
rect 145 -436 146 -435
rect 149 -436 150 -435
rect 170 -436 171 -435
rect 187 -436 188 -435
rect 215 -436 216 -435
rect 331 -436 332 -435
rect 359 -436 360 -435
rect 380 -436 381 -435
rect 44 -438 45 -437
rect 51 -438 52 -437
rect 86 -438 87 -437
rect 96 -438 97 -437
rect 114 -438 115 -437
rect 121 -438 122 -437
rect 170 -438 171 -437
rect 184 -438 185 -437
rect 226 -438 227 -437
rect 233 -438 234 -437
rect 247 -438 248 -437
rect 303 -438 304 -437
rect 362 -438 363 -437
rect 366 -438 367 -437
rect 51 -440 52 -439
rect 212 -440 213 -439
rect 229 -440 230 -439
rect 324 -440 325 -439
rect 65 -442 66 -441
rect 86 -442 87 -441
rect 93 -442 94 -441
rect 100 -442 101 -441
rect 177 -442 178 -441
rect 205 -442 206 -441
rect 254 -442 255 -441
rect 261 -442 262 -441
rect 268 -442 269 -441
rect 275 -442 276 -441
rect 303 -442 304 -441
rect 331 -442 332 -441
rect 75 -444 76 -443
rect 114 -444 115 -443
rect 117 -444 118 -443
rect 254 -444 255 -443
rect 275 -444 276 -443
rect 289 -444 290 -443
rect 93 -446 94 -445
rect 159 -446 160 -445
rect 198 -446 199 -445
rect 261 -446 262 -445
rect 289 -446 290 -445
rect 296 -446 297 -445
rect 135 -448 136 -447
rect 177 -448 178 -447
rect 191 -448 192 -447
rect 296 -448 297 -447
rect 194 -450 195 -449
rect 198 -450 199 -449
rect 205 -450 206 -449
rect 355 -450 356 -449
rect 194 -452 195 -451
rect 219 -452 220 -451
rect 156 -454 157 -453
rect 219 -454 220 -453
rect 26 -465 27 -464
rect 110 -465 111 -464
rect 121 -465 122 -464
rect 198 -465 199 -464
rect 212 -465 213 -464
rect 226 -465 227 -464
rect 250 -465 251 -464
rect 275 -465 276 -464
rect 296 -465 297 -464
rect 324 -465 325 -464
rect 338 -465 339 -464
rect 352 -465 353 -464
rect 366 -465 367 -464
rect 376 -465 377 -464
rect 33 -467 34 -466
rect 72 -467 73 -466
rect 79 -467 80 -466
rect 114 -467 115 -466
rect 121 -467 122 -466
rect 208 -467 209 -466
rect 215 -467 216 -466
rect 240 -467 241 -466
rect 254 -467 255 -466
rect 352 -467 353 -466
rect 37 -469 38 -468
rect 114 -469 115 -468
rect 142 -469 143 -468
rect 205 -469 206 -468
rect 240 -469 241 -468
rect 289 -469 290 -468
rect 317 -469 318 -468
rect 359 -469 360 -468
rect 37 -471 38 -470
rect 117 -471 118 -470
rect 149 -471 150 -470
rect 156 -471 157 -470
rect 177 -471 178 -470
rect 226 -471 227 -470
rect 261 -471 262 -470
rect 303 -471 304 -470
rect 331 -471 332 -470
rect 359 -471 360 -470
rect 44 -473 45 -472
rect 68 -473 69 -472
rect 72 -473 73 -472
rect 86 -473 87 -472
rect 93 -473 94 -472
rect 135 -473 136 -472
rect 177 -473 178 -472
rect 219 -473 220 -472
rect 275 -473 276 -472
rect 320 -473 321 -472
rect 331 -473 332 -472
rect 348 -473 349 -472
rect 44 -475 45 -474
rect 65 -475 66 -474
rect 86 -475 87 -474
rect 128 -475 129 -474
rect 135 -475 136 -474
rect 163 -475 164 -474
rect 184 -475 185 -474
rect 229 -475 230 -474
rect 282 -475 283 -474
rect 289 -475 290 -474
rect 58 -477 59 -476
rect 79 -477 80 -476
rect 107 -477 108 -476
rect 138 -477 139 -476
rect 163 -477 164 -476
rect 170 -477 171 -476
rect 187 -477 188 -476
rect 268 -477 269 -476
rect 51 -479 52 -478
rect 58 -479 59 -478
rect 128 -479 129 -478
rect 149 -479 150 -478
rect 170 -479 171 -478
rect 261 -479 262 -478
rect 51 -481 52 -480
rect 131 -481 132 -480
rect 173 -481 174 -480
rect 268 -481 269 -480
rect 100 -483 101 -482
rect 131 -483 132 -482
rect 191 -483 192 -482
rect 233 -483 234 -482
rect 100 -485 101 -484
rect 145 -485 146 -484
rect 194 -485 195 -484
rect 254 -485 255 -484
rect 198 -487 199 -486
rect 247 -487 248 -486
rect 205 -489 206 -488
rect 243 -489 244 -488
rect 233 -491 234 -490
rect 306 -491 307 -490
rect 16 -502 17 -501
rect 107 -502 108 -501
rect 156 -502 157 -501
rect 173 -502 174 -501
rect 177 -502 178 -501
rect 194 -502 195 -501
rect 201 -502 202 -501
rect 205 -502 206 -501
rect 222 -502 223 -501
rect 299 -502 300 -501
rect 338 -502 339 -501
rect 359 -502 360 -501
rect 30 -504 31 -503
rect 44 -504 45 -503
rect 51 -504 52 -503
rect 243 -504 244 -503
rect 268 -504 269 -503
rect 313 -504 314 -503
rect 345 -504 346 -503
rect 348 -504 349 -503
rect 352 -504 353 -503
rect 373 -504 374 -503
rect 65 -506 66 -505
rect 79 -506 80 -505
rect 86 -506 87 -505
rect 93 -506 94 -505
rect 110 -506 111 -505
rect 156 -506 157 -505
rect 159 -506 160 -505
rect 226 -506 227 -505
rect 275 -506 276 -505
rect 296 -506 297 -505
rect 317 -506 318 -505
rect 348 -506 349 -505
rect 51 -508 52 -507
rect 93 -508 94 -507
rect 163 -508 164 -507
rect 198 -508 199 -507
rect 226 -508 227 -507
rect 289 -508 290 -507
rect 296 -508 297 -507
rect 331 -508 332 -507
rect 341 -508 342 -507
rect 352 -508 353 -507
rect 44 -510 45 -509
rect 198 -510 199 -509
rect 208 -510 209 -509
rect 331 -510 332 -509
rect 341 -510 342 -509
rect 366 -510 367 -509
rect 65 -512 66 -511
rect 142 -512 143 -511
rect 149 -512 150 -511
rect 163 -512 164 -511
rect 166 -512 167 -511
rect 310 -512 311 -511
rect 68 -514 69 -513
rect 110 -514 111 -513
rect 170 -514 171 -513
rect 240 -514 241 -513
rect 282 -514 283 -513
rect 324 -514 325 -513
rect 72 -516 73 -515
rect 131 -516 132 -515
rect 191 -516 192 -515
rect 219 -516 220 -515
rect 233 -516 234 -515
rect 240 -516 241 -515
rect 247 -516 248 -515
rect 282 -516 283 -515
rect 289 -516 290 -515
rect 303 -516 304 -515
rect 37 -518 38 -517
rect 72 -518 73 -517
rect 79 -518 80 -517
rect 149 -518 150 -517
rect 194 -518 195 -517
rect 247 -518 248 -517
rect 261 -518 262 -517
rect 324 -518 325 -517
rect 37 -520 38 -519
rect 58 -520 59 -519
rect 86 -520 87 -519
rect 100 -520 101 -519
rect 114 -520 115 -519
rect 219 -520 220 -519
rect 229 -520 230 -519
rect 303 -520 304 -519
rect 58 -522 59 -521
rect 121 -522 122 -521
rect 142 -522 143 -521
rect 233 -522 234 -521
rect 100 -524 101 -523
rect 268 -524 269 -523
rect 114 -526 115 -525
rect 135 -526 136 -525
rect 201 -526 202 -525
rect 261 -526 262 -525
rect 135 -528 136 -527
rect 184 -528 185 -527
rect 177 -530 178 -529
rect 184 -530 185 -529
rect 9 -541 10 -540
rect 107 -541 108 -540
rect 121 -541 122 -540
rect 149 -541 150 -540
rect 156 -541 157 -540
rect 219 -541 220 -540
rect 222 -541 223 -540
rect 331 -541 332 -540
rect 338 -541 339 -540
rect 373 -541 374 -540
rect 16 -543 17 -542
rect 229 -543 230 -542
rect 275 -543 276 -542
rect 289 -543 290 -542
rect 348 -543 349 -542
rect 352 -543 353 -542
rect 16 -545 17 -544
rect 51 -545 52 -544
rect 58 -545 59 -544
rect 166 -545 167 -544
rect 177 -545 178 -544
rect 205 -545 206 -544
rect 208 -545 209 -544
rect 289 -545 290 -544
rect 23 -547 24 -546
rect 26 -547 27 -546
rect 37 -547 38 -546
rect 82 -547 83 -546
rect 86 -547 87 -546
rect 103 -547 104 -546
rect 131 -547 132 -546
rect 345 -547 346 -546
rect 44 -549 45 -548
rect 124 -549 125 -548
rect 142 -549 143 -548
rect 205 -549 206 -548
rect 226 -549 227 -548
rect 261 -549 262 -548
rect 275 -549 276 -548
rect 366 -549 367 -548
rect 30 -551 31 -550
rect 44 -551 45 -550
rect 58 -551 59 -550
rect 79 -551 80 -550
rect 86 -551 87 -550
rect 110 -551 111 -550
rect 114 -551 115 -550
rect 131 -551 132 -550
rect 145 -551 146 -550
rect 247 -551 248 -550
rect 254 -551 255 -550
rect 261 -551 262 -550
rect 65 -553 66 -552
rect 152 -553 153 -552
rect 177 -553 178 -552
rect 236 -553 237 -552
rect 247 -553 248 -552
rect 278 -553 279 -552
rect 65 -555 66 -554
rect 159 -555 160 -554
rect 191 -555 192 -554
rect 233 -555 234 -554
rect 268 -555 269 -554
rect 278 -555 279 -554
rect 72 -557 73 -556
rect 135 -557 136 -556
rect 201 -557 202 -556
rect 282 -557 283 -556
rect 93 -559 94 -558
rect 240 -559 241 -558
rect 268 -559 269 -558
rect 324 -559 325 -558
rect 93 -561 94 -560
rect 145 -561 146 -560
rect 240 -561 241 -560
rect 303 -561 304 -560
rect 317 -561 318 -560
rect 324 -561 325 -560
rect 100 -563 101 -562
rect 198 -563 199 -562
rect 282 -563 283 -562
rect 292 -563 293 -562
rect 303 -563 304 -562
rect 310 -563 311 -562
rect 100 -565 101 -564
rect 128 -565 129 -564
rect 135 -565 136 -564
rect 152 -565 153 -564
rect 198 -565 199 -564
rect 212 -565 213 -564
rect 114 -567 115 -566
rect 124 -567 125 -566
rect 170 -567 171 -566
rect 212 -567 213 -566
rect 163 -569 164 -568
rect 170 -569 171 -568
rect 9 -580 10 -579
rect 156 -580 157 -579
rect 159 -580 160 -579
rect 198 -580 199 -579
rect 205 -580 206 -579
rect 233 -580 234 -579
rect 257 -580 258 -579
rect 261 -580 262 -579
rect 282 -580 283 -579
rect 310 -580 311 -579
rect 355 -580 356 -579
rect 359 -580 360 -579
rect 16 -582 17 -581
rect 51 -582 52 -581
rect 65 -582 66 -581
rect 96 -582 97 -581
rect 100 -582 101 -581
rect 110 -582 111 -581
rect 135 -582 136 -581
rect 142 -582 143 -581
rect 187 -582 188 -581
rect 191 -582 192 -581
rect 198 -582 199 -581
rect 219 -582 220 -581
rect 226 -582 227 -581
rect 254 -582 255 -581
rect 261 -582 262 -581
rect 268 -582 269 -581
rect 282 -582 283 -581
rect 306 -582 307 -581
rect 30 -584 31 -583
rect 82 -584 83 -583
rect 86 -584 87 -583
rect 145 -584 146 -583
rect 163 -584 164 -583
rect 191 -584 192 -583
rect 205 -584 206 -583
rect 229 -584 230 -583
rect 268 -584 269 -583
rect 278 -584 279 -583
rect 289 -584 290 -583
rect 303 -584 304 -583
rect 51 -586 52 -585
rect 131 -586 132 -585
rect 135 -586 136 -585
rect 138 -586 139 -585
rect 163 -586 164 -585
rect 184 -586 185 -585
rect 219 -586 220 -585
rect 240 -586 241 -585
rect 296 -586 297 -585
rect 303 -586 304 -585
rect 58 -588 59 -587
rect 65 -588 66 -587
rect 72 -588 73 -587
rect 152 -588 153 -587
rect 177 -588 178 -587
rect 187 -588 188 -587
rect 58 -590 59 -589
rect 100 -590 101 -589
rect 152 -590 153 -589
rect 212 -590 213 -589
rect 75 -592 76 -591
rect 128 -592 129 -591
rect 170 -592 171 -591
rect 177 -592 178 -591
rect 212 -592 213 -591
rect 247 -592 248 -591
rect 86 -594 87 -593
rect 114 -594 115 -593
rect 159 -594 160 -593
rect 247 -594 248 -593
rect 93 -596 94 -595
rect 107 -596 108 -595
rect 114 -596 115 -595
rect 121 -596 122 -595
rect 79 -598 80 -597
rect 93 -598 94 -597
rect 107 -598 108 -597
rect 149 -598 150 -597
rect 33 -600 34 -599
rect 79 -600 80 -599
rect 30 -611 31 -610
rect 82 -611 83 -610
rect 100 -611 101 -610
rect 103 -611 104 -610
rect 114 -611 115 -610
rect 128 -611 129 -610
rect 131 -611 132 -610
rect 149 -611 150 -610
rect 156 -611 157 -610
rect 180 -611 181 -610
rect 184 -611 185 -610
rect 212 -611 213 -610
rect 226 -611 227 -610
rect 254 -611 255 -610
rect 257 -611 258 -610
rect 282 -611 283 -610
rect 37 -613 38 -612
rect 44 -613 45 -612
rect 51 -613 52 -612
rect 117 -613 118 -612
rect 135 -613 136 -612
rect 191 -613 192 -612
rect 205 -613 206 -612
rect 226 -613 227 -612
rect 233 -613 234 -612
rect 264 -613 265 -612
rect 275 -613 276 -612
rect 289 -613 290 -612
rect 51 -615 52 -614
rect 72 -615 73 -614
rect 86 -615 87 -614
rect 117 -615 118 -614
rect 135 -615 136 -614
rect 142 -615 143 -614
rect 159 -615 160 -614
rect 198 -615 199 -614
rect 205 -615 206 -614
rect 219 -615 220 -614
rect 233 -615 234 -614
rect 261 -615 262 -614
rect 58 -617 59 -616
rect 138 -617 139 -616
rect 142 -617 143 -616
rect 156 -617 157 -616
rect 163 -617 164 -616
rect 173 -617 174 -616
rect 177 -617 178 -616
rect 180 -617 181 -616
rect 187 -617 188 -616
rect 212 -617 213 -616
rect 240 -617 241 -616
rect 247 -617 248 -616
rect 261 -617 262 -616
rect 268 -617 269 -616
rect 65 -619 66 -618
rect 86 -619 87 -618
rect 114 -619 115 -618
rect 145 -619 146 -618
rect 152 -619 153 -618
rect 219 -619 220 -618
rect 243 -619 244 -618
rect 247 -619 248 -618
rect 65 -621 66 -620
rect 107 -621 108 -620
rect 121 -621 122 -620
rect 163 -621 164 -620
rect 170 -621 171 -620
rect 198 -621 199 -620
rect 79 -623 80 -622
rect 121 -623 122 -622
rect 191 -623 192 -622
rect 254 -623 255 -622
rect 75 -625 76 -624
rect 79 -625 80 -624
rect 93 -625 94 -624
rect 107 -625 108 -624
rect 30 -636 31 -635
rect 51 -636 52 -635
rect 65 -636 66 -635
rect 107 -636 108 -635
rect 121 -636 122 -635
rect 149 -636 150 -635
rect 152 -636 153 -635
rect 191 -636 192 -635
rect 201 -636 202 -635
rect 268 -636 269 -635
rect 37 -638 38 -637
rect 72 -638 73 -637
rect 82 -638 83 -637
rect 100 -638 101 -637
rect 107 -638 108 -637
rect 117 -638 118 -637
rect 124 -638 125 -637
rect 163 -638 164 -637
rect 184 -638 185 -637
rect 240 -638 241 -637
rect 247 -638 248 -637
rect 289 -638 290 -637
rect 44 -640 45 -639
rect 75 -640 76 -639
rect 96 -640 97 -639
rect 233 -640 234 -639
rect 254 -640 255 -639
rect 257 -640 258 -639
rect 51 -642 52 -641
rect 93 -642 94 -641
rect 100 -642 101 -641
rect 121 -642 122 -641
rect 135 -642 136 -641
rect 145 -642 146 -641
rect 149 -642 150 -641
rect 187 -642 188 -641
rect 205 -642 206 -641
rect 233 -642 234 -641
rect 68 -644 69 -643
rect 79 -644 80 -643
rect 128 -644 129 -643
rect 135 -644 136 -643
rect 142 -644 143 -643
rect 261 -644 262 -643
rect 75 -646 76 -645
rect 86 -646 87 -645
rect 128 -646 129 -645
rect 138 -646 139 -645
rect 156 -646 157 -645
rect 173 -646 174 -645
rect 187 -646 188 -645
rect 296 -646 297 -645
rect 156 -648 157 -647
rect 163 -648 164 -647
rect 170 -648 171 -647
rect 247 -648 248 -647
rect 212 -650 213 -649
rect 240 -650 241 -649
rect 198 -652 199 -651
rect 212 -652 213 -651
rect 219 -652 220 -651
rect 282 -652 283 -651
rect 219 -654 220 -653
rect 236 -654 237 -653
rect 226 -656 227 -655
rect 275 -656 276 -655
rect 191 -658 192 -657
rect 226 -658 227 -657
rect 37 -669 38 -668
rect 110 -669 111 -668
rect 114 -669 115 -668
rect 142 -669 143 -668
rect 156 -669 157 -668
rect 226 -669 227 -668
rect 254 -669 255 -668
rect 278 -669 279 -668
rect 44 -671 45 -670
rect 145 -671 146 -670
rect 156 -671 157 -670
rect 163 -671 164 -670
rect 173 -671 174 -670
rect 268 -671 269 -670
rect 51 -673 52 -672
rect 117 -673 118 -672
rect 121 -673 122 -672
rect 191 -673 192 -672
rect 198 -673 199 -672
rect 212 -673 213 -672
rect 247 -673 248 -672
rect 254 -673 255 -672
rect 261 -673 262 -672
rect 268 -673 269 -672
rect 58 -675 59 -674
rect 86 -675 87 -674
rect 89 -675 90 -674
rect 138 -675 139 -674
rect 159 -675 160 -674
rect 201 -675 202 -674
rect 208 -675 209 -674
rect 275 -675 276 -674
rect 61 -677 62 -676
rect 68 -677 69 -676
rect 93 -677 94 -676
rect 184 -677 185 -676
rect 187 -677 188 -676
rect 233 -677 234 -676
rect 30 -679 31 -678
rect 61 -679 62 -678
rect 93 -679 94 -678
rect 149 -679 150 -678
rect 180 -679 181 -678
rect 282 -679 283 -678
rect 96 -681 97 -680
rect 100 -681 101 -680
rect 138 -681 139 -680
rect 163 -681 164 -680
rect 180 -681 181 -680
rect 289 -681 290 -680
rect 100 -683 101 -682
rect 107 -683 108 -682
rect 191 -683 192 -682
rect 226 -683 227 -682
rect 107 -685 108 -684
rect 170 -685 171 -684
rect 212 -685 213 -684
rect 240 -685 241 -684
rect 177 -687 178 -686
rect 240 -687 241 -686
rect 219 -689 220 -688
rect 233 -689 234 -688
rect 177 -691 178 -690
rect 219 -691 220 -690
rect 61 -702 62 -701
rect 72 -702 73 -701
rect 75 -702 76 -701
rect 79 -702 80 -701
rect 100 -702 101 -701
rect 117 -702 118 -701
rect 121 -702 122 -701
rect 177 -702 178 -701
rect 184 -702 185 -701
rect 226 -702 227 -701
rect 240 -702 241 -701
rect 261 -702 262 -701
rect 114 -704 115 -703
rect 121 -704 122 -703
rect 128 -704 129 -703
rect 135 -704 136 -703
rect 142 -704 143 -703
rect 187 -704 188 -703
rect 194 -704 195 -703
rect 198 -704 199 -703
rect 240 -704 241 -703
rect 254 -704 255 -703
rect 131 -706 132 -705
rect 142 -706 143 -705
rect 149 -706 150 -705
rect 170 -706 171 -705
rect 194 -706 195 -705
rect 219 -706 220 -705
rect 247 -706 248 -705
rect 268 -706 269 -705
rect 93 -708 94 -707
rect 170 -708 171 -707
rect 198 -708 199 -707
rect 233 -708 234 -707
rect 152 -710 153 -709
rect 205 -710 206 -709
rect 163 -712 164 -711
rect 173 -712 174 -711
rect 205 -712 206 -711
rect 215 -712 216 -711
rect 163 -714 164 -713
rect 180 -714 181 -713
rect 114 -725 115 -724
rect 131 -725 132 -724
rect 135 -725 136 -724
rect 142 -725 143 -724
rect 159 -725 160 -724
rect 177 -725 178 -724
rect 180 -725 181 -724
rect 184 -725 185 -724
rect 191 -725 192 -724
rect 205 -725 206 -724
rect 229 -725 230 -724
rect 240 -725 241 -724
rect 121 -727 122 -726
rect 131 -727 132 -726
rect 163 -727 164 -726
rect 170 -727 171 -726
rect 173 -727 174 -726
rect 198 -727 199 -726
rect 117 -729 118 -728
rect 121 -729 122 -728
rect 177 -729 178 -728
rect 184 -729 185 -728
rect 191 -729 192 -728
rect 194 -729 195 -728
rect 128 -740 129 -739
rect 135 -740 136 -739
rect 149 -740 150 -739
rect 163 -740 164 -739
rect 166 -740 167 -739
rect 170 -740 171 -739
rect 177 -740 178 -739
rect 184 -740 185 -739
rect 187 -740 188 -739
rect 191 -740 192 -739
rect 121 -742 122 -741
rect 128 -742 129 -741
rect 156 -742 157 -741
rect 170 -742 171 -741
rect 124 -753 125 -752
rect 128 -753 129 -752
rect 156 -753 157 -752
rect 170 -753 171 -752
rect 184 -753 185 -752
rect 191 -753 192 -752
rect 159 -755 160 -754
rect 163 -755 164 -754
<< metal2 >>
rect 103 -3 104 1
rect 107 -3 108 1
rect 128 -3 129 1
rect 135 -3 136 1
rect 142 -3 143 1
rect 156 -3 157 1
rect 177 -3 178 1
rect 191 -3 192 1
rect 194 -3 195 1
rect 212 -3 213 1
rect 198 -3 199 -1
rect 205 -3 206 -1
rect 79 -22 80 -12
rect 96 -22 97 -12
rect 100 -22 101 -12
rect 103 -13 104 -11
rect 110 -22 111 -12
rect 121 -22 122 -12
rect 135 -13 136 -11
rect 142 -13 143 -11
rect 149 -13 150 -11
rect 156 -13 157 -11
rect 170 -22 171 -12
rect 194 -22 195 -12
rect 208 -22 209 -12
rect 233 -22 234 -12
rect 135 -22 136 -14
rect 156 -22 157 -14
rect 177 -15 178 -11
rect 184 -15 185 -11
rect 212 -15 213 -11
rect 226 -22 227 -14
rect 142 -22 143 -16
rect 173 -17 174 -11
rect 184 -22 185 -16
rect 198 -17 199 -11
rect 215 -22 216 -16
rect 219 -22 220 -16
rect 149 -22 150 -18
rect 163 -19 164 -11
rect 152 -22 153 -20
rect 198 -22 199 -20
rect 65 -45 66 -31
rect 89 -32 90 -30
rect 93 -32 94 -30
rect 96 -40 97 -31
rect 114 -45 115 -31
rect 173 -45 174 -31
rect 184 -32 185 -30
rect 247 -45 248 -31
rect 271 -45 272 -31
rect 275 -45 276 -31
rect 72 -45 73 -33
rect 110 -45 111 -33
rect 128 -34 129 -30
rect 128 -45 129 -33
rect 128 -34 129 -30
rect 128 -45 129 -33
rect 142 -34 143 -30
rect 187 -34 188 -30
rect 198 -34 199 -30
rect 226 -45 227 -33
rect 229 -34 230 -30
rect 282 -45 283 -33
rect 79 -36 80 -30
rect 79 -45 80 -35
rect 79 -36 80 -30
rect 79 -45 80 -35
rect 86 -36 87 -30
rect 89 -45 90 -35
rect 93 -45 94 -35
rect 100 -36 101 -30
rect 149 -36 150 -30
rect 170 -36 171 -30
rect 180 -45 181 -35
rect 184 -45 185 -35
rect 201 -45 202 -35
rect 254 -45 255 -35
rect 86 -45 87 -37
rect 107 -38 108 -30
rect 135 -38 136 -30
rect 149 -45 150 -37
rect 152 -45 153 -37
rect 240 -45 241 -37
rect 100 -45 101 -39
rect 121 -40 122 -30
rect 135 -45 136 -39
rect 156 -40 157 -30
rect 163 -45 164 -39
rect 215 -45 216 -39
rect 219 -40 220 -30
rect 233 -40 234 -30
rect 261 -45 262 -39
rect 156 -45 157 -41
rect 170 -45 171 -41
rect 191 -42 192 -30
rect 233 -45 234 -41
rect 159 -44 160 -30
rect 166 -44 167 -30
rect 177 -44 178 -30
rect 191 -45 192 -43
rect 205 -45 206 -43
rect 219 -45 220 -43
rect 30 -76 31 -54
rect 75 -76 76 -54
rect 82 -55 83 -53
rect 145 -55 146 -53
rect 170 -55 171 -53
rect 261 -55 262 -53
rect 44 -76 45 -56
rect 114 -57 115 -53
rect 117 -76 118 -56
rect 149 -76 150 -56
rect 163 -57 164 -53
rect 170 -76 171 -56
rect 184 -57 185 -53
rect 261 -76 262 -56
rect 51 -76 52 -58
rect 131 -59 132 -53
rect 159 -76 160 -58
rect 163 -76 164 -58
rect 187 -76 188 -58
rect 289 -76 290 -58
rect 58 -76 59 -60
rect 156 -61 157 -53
rect 191 -61 192 -53
rect 198 -61 199 -53
rect 201 -61 202 -53
rect 240 -61 241 -53
rect 243 -76 244 -60
rect 303 -76 304 -60
rect 61 -63 62 -53
rect 89 -63 90 -53
rect 93 -76 94 -62
rect 177 -76 178 -62
rect 198 -76 199 -62
rect 226 -63 227 -53
rect 233 -63 234 -53
rect 268 -76 269 -62
rect 65 -65 66 -53
rect 86 -76 87 -64
rect 100 -65 101 -53
rect 114 -76 115 -64
rect 121 -65 122 -53
rect 135 -65 136 -53
rect 142 -65 143 -53
rect 191 -76 192 -64
rect 219 -76 220 -64
rect 275 -65 276 -53
rect 65 -76 66 -66
rect 96 -67 97 -53
rect 100 -76 101 -66
rect 138 -76 139 -66
rect 180 -76 181 -66
rect 226 -76 227 -66
rect 254 -67 255 -53
rect 275 -76 276 -66
rect 72 -69 73 -53
rect 135 -76 136 -68
rect 184 -76 185 -68
rect 233 -76 234 -68
rect 72 -76 73 -70
rect 79 -76 80 -70
rect 103 -76 104 -70
rect 142 -76 143 -70
rect 212 -71 213 -53
rect 254 -76 255 -70
rect 110 -73 111 -53
rect 124 -73 125 -53
rect 205 -73 206 -53
rect 212 -76 213 -72
rect 222 -73 223 -53
rect 282 -73 283 -53
rect 121 -76 122 -74
rect 156 -76 157 -74
rect 247 -75 248 -53
rect 282 -76 283 -74
rect 16 -121 17 -85
rect 79 -86 80 -84
rect 86 -86 87 -84
rect 100 -86 101 -84
rect 103 -121 104 -85
rect 107 -86 108 -84
rect 114 -86 115 -84
rect 135 -121 136 -85
rect 170 -86 171 -84
rect 180 -86 181 -84
rect 184 -121 185 -85
rect 194 -121 195 -85
rect 201 -86 202 -84
rect 236 -121 237 -85
rect 243 -86 244 -84
rect 282 -86 283 -84
rect 299 -86 300 -84
rect 331 -121 332 -85
rect 30 -88 31 -84
rect 324 -121 325 -87
rect 26 -121 27 -89
rect 30 -121 31 -89
rect 37 -90 38 -84
rect 79 -121 80 -89
rect 100 -121 101 -89
rect 208 -90 209 -84
rect 250 -90 251 -84
rect 289 -90 290 -84
rect 37 -121 38 -91
rect 93 -92 94 -84
rect 107 -121 108 -91
rect 124 -121 125 -91
rect 131 -121 132 -91
rect 226 -92 227 -84
rect 254 -92 255 -84
rect 254 -121 255 -91
rect 254 -92 255 -84
rect 254 -121 255 -91
rect 268 -92 269 -84
rect 310 -121 311 -91
rect 44 -94 45 -84
rect 110 -94 111 -84
rect 138 -94 139 -84
rect 282 -121 283 -93
rect 51 -96 52 -84
rect 187 -96 188 -84
rect 191 -96 192 -84
rect 240 -121 241 -95
rect 275 -96 276 -84
rect 317 -121 318 -95
rect 58 -98 59 -84
rect 128 -98 129 -84
rect 142 -98 143 -84
rect 289 -121 290 -97
rect 65 -100 66 -84
rect 86 -121 87 -99
rect 93 -121 94 -99
rect 138 -121 139 -99
rect 163 -100 164 -84
rect 170 -121 171 -99
rect 177 -100 178 -84
rect 261 -100 262 -84
rect 51 -121 52 -101
rect 65 -121 66 -101
rect 68 -121 69 -101
rect 159 -121 160 -101
rect 180 -121 181 -101
rect 212 -121 213 -101
rect 219 -102 220 -84
rect 226 -121 227 -101
rect 72 -121 73 -103
rect 117 -104 118 -84
rect 128 -121 129 -103
rect 152 -121 153 -103
rect 187 -121 188 -103
rect 261 -121 262 -103
rect 117 -121 118 -105
rect 268 -121 269 -105
rect 198 -108 199 -84
rect 275 -121 276 -107
rect 198 -121 199 -109
rect 303 -110 304 -84
rect 149 -112 150 -84
rect 303 -121 304 -111
rect 121 -114 122 -84
rect 149 -121 150 -113
rect 201 -121 202 -113
rect 233 -114 234 -84
rect 205 -116 206 -84
rect 296 -121 297 -115
rect 205 -121 206 -117
rect 247 -121 248 -117
rect 208 -121 209 -119
rect 219 -121 220 -119
rect 23 -131 24 -129
rect 145 -131 146 -129
rect 159 -131 160 -129
rect 240 -131 241 -129
rect 275 -131 276 -129
rect 275 -168 276 -130
rect 275 -131 276 -129
rect 275 -168 276 -130
rect 26 -168 27 -132
rect 30 -133 31 -129
rect 37 -133 38 -129
rect 180 -133 181 -129
rect 198 -133 199 -129
rect 247 -133 248 -129
rect 23 -168 24 -134
rect 30 -168 31 -134
rect 44 -168 45 -134
rect 51 -135 52 -129
rect 61 -135 62 -129
rect 89 -168 90 -134
rect 100 -135 101 -129
rect 282 -135 283 -129
rect 37 -168 38 -136
rect 61 -168 62 -136
rect 65 -137 66 -129
rect 324 -137 325 -129
rect 47 -139 48 -129
rect 65 -168 66 -138
rect 72 -139 73 -129
rect 82 -139 83 -129
rect 86 -139 87 -129
rect 117 -139 118 -129
rect 128 -139 129 -129
rect 243 -168 244 -138
rect 72 -168 73 -140
rect 93 -141 94 -129
rect 100 -168 101 -140
rect 107 -141 108 -129
rect 110 -168 111 -140
rect 114 -141 115 -129
rect 117 -168 118 -140
rect 124 -168 125 -140
rect 128 -168 129 -140
rect 152 -141 153 -129
rect 166 -168 167 -140
rect 194 -168 195 -140
rect 205 -141 206 -129
rect 268 -141 269 -129
rect 16 -143 17 -129
rect 114 -168 115 -142
rect 135 -143 136 -129
rect 289 -143 290 -129
rect 79 -145 80 -129
rect 93 -168 94 -144
rect 142 -145 143 -129
rect 303 -145 304 -129
rect 79 -168 80 -146
rect 152 -168 153 -146
rect 170 -147 171 -129
rect 184 -147 185 -129
rect 205 -168 206 -146
rect 310 -147 311 -129
rect 131 -149 132 -129
rect 170 -168 171 -148
rect 177 -149 178 -129
rect 187 -149 188 -129
rect 201 -149 202 -129
rect 310 -168 311 -148
rect 103 -151 104 -129
rect 177 -168 178 -150
rect 201 -168 202 -150
rect 289 -168 290 -150
rect 303 -168 304 -150
rect 331 -151 332 -129
rect 142 -168 143 -152
rect 159 -168 160 -152
rect 215 -168 216 -152
rect 296 -153 297 -129
rect 156 -155 157 -129
rect 184 -168 185 -154
rect 219 -155 220 -129
rect 219 -168 220 -154
rect 219 -155 220 -129
rect 219 -168 220 -154
rect 226 -155 227 -129
rect 229 -167 230 -154
rect 233 -155 234 -129
rect 296 -168 297 -154
rect 212 -157 213 -129
rect 233 -168 234 -156
rect 236 -157 237 -129
rect 317 -157 318 -129
rect 212 -168 213 -158
rect 247 -168 248 -158
rect 226 -168 227 -160
rect 261 -161 262 -129
rect 236 -168 237 -162
rect 282 -168 283 -162
rect 254 -165 255 -129
rect 261 -168 262 -164
rect 254 -168 255 -166
rect 16 -205 17 -177
rect 33 -205 34 -177
rect 37 -205 38 -177
rect 68 -205 69 -177
rect 72 -178 73 -176
rect 86 -178 87 -176
rect 89 -205 90 -177
rect 110 -178 111 -176
rect 121 -205 122 -177
rect 128 -178 129 -176
rect 135 -178 136 -176
rect 142 -178 143 -176
rect 145 -205 146 -177
rect 394 -205 395 -177
rect 9 -205 10 -179
rect 86 -205 87 -179
rect 100 -180 101 -176
rect 100 -205 101 -179
rect 100 -180 101 -176
rect 100 -205 101 -179
rect 149 -180 150 -176
rect 198 -205 199 -179
rect 222 -205 223 -179
rect 296 -180 297 -176
rect 303 -180 304 -176
rect 359 -205 360 -179
rect 19 -182 20 -176
rect 58 -182 59 -176
rect 72 -205 73 -181
rect 135 -205 136 -181
rect 149 -205 150 -181
rect 184 -182 185 -176
rect 191 -205 192 -181
rect 215 -205 216 -181
rect 240 -182 241 -176
rect 261 -182 262 -176
rect 268 -182 269 -176
rect 331 -205 332 -181
rect 23 -205 24 -183
rect 30 -184 31 -176
rect 44 -184 45 -176
rect 51 -184 52 -176
rect 54 -205 55 -183
rect 58 -205 59 -183
rect 79 -184 80 -176
rect 107 -184 108 -176
rect 117 -184 118 -176
rect 240 -205 241 -183
rect 243 -184 244 -176
rect 324 -205 325 -183
rect 44 -205 45 -185
rect 184 -205 185 -185
rect 194 -186 195 -176
rect 226 -186 227 -176
rect 247 -186 248 -176
rect 261 -205 262 -185
rect 271 -205 272 -185
rect 303 -205 304 -185
rect 310 -186 311 -176
rect 373 -205 374 -185
rect 51 -205 52 -187
rect 93 -188 94 -176
rect 107 -205 108 -187
rect 236 -205 237 -187
rect 247 -205 248 -187
rect 387 -205 388 -187
rect 65 -190 66 -176
rect 79 -205 80 -189
rect 93 -205 94 -189
rect 205 -190 206 -176
rect 212 -205 213 -189
rect 310 -205 311 -189
rect 117 -205 118 -191
rect 124 -192 125 -176
rect 156 -192 157 -176
rect 163 -205 164 -191
rect 170 -192 171 -176
rect 205 -205 206 -191
rect 275 -192 276 -176
rect 296 -205 297 -191
rect 114 -205 115 -193
rect 275 -205 276 -193
rect 282 -194 283 -176
rect 338 -205 339 -193
rect 128 -205 129 -195
rect 156 -205 157 -195
rect 159 -196 160 -176
rect 219 -196 220 -176
rect 285 -205 286 -195
rect 352 -205 353 -195
rect 170 -205 171 -197
rect 208 -198 209 -176
rect 219 -205 220 -197
rect 380 -205 381 -197
rect 177 -200 178 -176
rect 226 -205 227 -199
rect 289 -200 290 -176
rect 345 -205 346 -199
rect 177 -205 178 -201
rect 254 -202 255 -176
rect 289 -205 290 -201
rect 317 -205 318 -201
rect 201 -204 202 -176
rect 254 -205 255 -203
rect 292 -205 293 -203
rect 366 -205 367 -203
rect 9 -215 10 -213
rect 142 -215 143 -213
rect 149 -215 150 -213
rect 184 -250 185 -214
rect 187 -215 188 -213
rect 345 -215 346 -213
rect 352 -215 353 -213
rect 352 -250 353 -214
rect 352 -215 353 -213
rect 352 -250 353 -214
rect 9 -250 10 -216
rect 75 -217 76 -213
rect 86 -250 87 -216
rect 100 -217 101 -213
rect 114 -217 115 -213
rect 135 -217 136 -213
rect 156 -217 157 -213
rect 170 -217 171 -213
rect 177 -217 178 -213
rect 215 -217 216 -213
rect 222 -217 223 -213
rect 373 -217 374 -213
rect 16 -219 17 -213
rect 54 -219 55 -213
rect 72 -219 73 -213
rect 79 -219 80 -213
rect 93 -219 94 -213
rect 159 -250 160 -218
rect 163 -219 164 -213
rect 233 -219 234 -213
rect 261 -219 262 -213
rect 282 -250 283 -218
rect 289 -250 290 -218
rect 324 -219 325 -213
rect 16 -250 17 -220
rect 124 -250 125 -220
rect 128 -221 129 -213
rect 142 -250 143 -220
rect 170 -250 171 -220
rect 219 -221 220 -213
rect 229 -250 230 -220
rect 359 -221 360 -213
rect 26 -250 27 -222
rect 110 -223 111 -213
rect 117 -223 118 -213
rect 380 -223 381 -213
rect 30 -250 31 -224
rect 191 -225 192 -213
rect 215 -250 216 -224
rect 296 -225 297 -213
rect 366 -225 367 -213
rect 380 -250 381 -224
rect 37 -227 38 -213
rect 163 -250 164 -226
rect 191 -250 192 -226
rect 254 -227 255 -213
rect 268 -227 269 -213
rect 338 -227 339 -213
rect 37 -250 38 -228
rect 121 -229 122 -213
rect 128 -250 129 -228
rect 212 -250 213 -228
rect 219 -250 220 -228
rect 226 -229 227 -213
rect 233 -250 234 -228
rect 247 -229 248 -213
rect 254 -250 255 -228
rect 285 -229 286 -213
rect 292 -250 293 -228
rect 345 -250 346 -228
rect 44 -231 45 -213
rect 177 -250 178 -230
rect 198 -231 199 -213
rect 268 -250 269 -230
rect 296 -250 297 -230
rect 303 -231 304 -213
rect 44 -250 45 -232
rect 82 -250 83 -232
rect 89 -233 90 -213
rect 359 -250 360 -232
rect 51 -250 52 -234
rect 58 -235 59 -213
rect 72 -250 73 -234
rect 79 -250 80 -234
rect 93 -250 94 -234
rect 110 -250 111 -234
rect 114 -250 115 -234
rect 226 -250 227 -234
rect 240 -235 241 -213
rect 324 -250 325 -234
rect 58 -250 59 -236
rect 152 -250 153 -236
rect 156 -250 157 -236
rect 247 -250 248 -236
rect 303 -250 304 -236
rect 310 -237 311 -213
rect 121 -250 122 -238
rect 394 -239 395 -213
rect 198 -250 199 -240
rect 331 -241 332 -213
rect 208 -243 209 -213
rect 338 -250 339 -242
rect 208 -250 209 -244
rect 275 -245 276 -213
rect 310 -250 311 -244
rect 317 -245 318 -213
rect 331 -250 332 -244
rect 373 -250 374 -244
rect 201 -250 202 -246
rect 317 -250 318 -246
rect 240 -250 241 -248
rect 275 -250 276 -248
rect 2 -297 3 -259
rect 124 -260 125 -258
rect 138 -260 139 -258
rect 254 -260 255 -258
rect 264 -260 265 -258
rect 296 -260 297 -258
rect 345 -260 346 -258
rect 345 -297 346 -259
rect 345 -260 346 -258
rect 345 -297 346 -259
rect 359 -260 360 -258
rect 369 -260 370 -258
rect 376 -297 377 -259
rect 380 -260 381 -258
rect 9 -262 10 -258
rect 75 -262 76 -258
rect 79 -297 80 -261
rect 107 -262 108 -258
rect 121 -297 122 -261
rect 156 -297 157 -261
rect 166 -297 167 -261
rect 261 -297 262 -261
rect 275 -262 276 -258
rect 331 -262 332 -258
rect 366 -262 367 -258
rect 369 -297 370 -261
rect 9 -297 10 -263
rect 58 -264 59 -258
rect 65 -297 66 -263
rect 128 -264 129 -258
rect 149 -297 150 -263
rect 177 -264 178 -258
rect 184 -264 185 -258
rect 257 -297 258 -263
rect 275 -297 276 -263
rect 282 -264 283 -258
rect 289 -264 290 -258
rect 352 -264 353 -258
rect 366 -297 367 -263
rect 380 -297 381 -263
rect 16 -266 17 -258
rect 100 -266 101 -258
rect 107 -297 108 -265
rect 208 -266 209 -258
rect 212 -297 213 -265
rect 219 -266 220 -258
rect 247 -266 248 -258
rect 282 -297 283 -265
rect 289 -297 290 -265
rect 317 -266 318 -258
rect 16 -297 17 -267
rect 103 -268 104 -258
rect 152 -268 153 -258
rect 191 -268 192 -258
rect 205 -268 206 -258
rect 240 -268 241 -258
rect 250 -297 251 -267
rect 331 -297 332 -267
rect 37 -270 38 -258
rect 201 -270 202 -258
rect 215 -270 216 -258
rect 359 -297 360 -269
rect 23 -297 24 -271
rect 215 -297 216 -271
rect 233 -272 234 -258
rect 240 -297 241 -271
rect 296 -297 297 -271
rect 338 -272 339 -258
rect 44 -274 45 -258
rect 124 -297 125 -273
rect 163 -274 164 -258
rect 177 -297 178 -273
rect 191 -297 192 -273
rect 226 -274 227 -258
rect 303 -274 304 -258
rect 317 -297 318 -273
rect 51 -276 52 -258
rect 54 -297 55 -275
rect 68 -276 69 -258
rect 82 -276 83 -258
rect 86 -276 87 -258
rect 128 -297 129 -275
rect 170 -276 171 -258
rect 219 -297 220 -275
rect 303 -297 304 -275
rect 324 -276 325 -258
rect 37 -297 38 -277
rect 51 -297 52 -277
rect 72 -278 73 -258
rect 86 -297 87 -277
rect 93 -278 94 -258
rect 159 -278 160 -258
rect 170 -297 171 -277
rect 184 -297 185 -277
rect 198 -278 199 -258
rect 226 -297 227 -277
rect 268 -278 269 -258
rect 324 -297 325 -277
rect 30 -280 31 -258
rect 198 -297 199 -279
rect 201 -297 202 -279
rect 352 -297 353 -279
rect 30 -297 31 -281
rect 135 -282 136 -258
rect 205 -297 206 -281
rect 268 -297 269 -281
rect 310 -282 311 -258
rect 338 -297 339 -281
rect 44 -297 45 -283
rect 159 -297 160 -283
rect 61 -297 62 -285
rect 310 -297 311 -285
rect 72 -297 73 -287
rect 208 -297 209 -287
rect 93 -297 94 -289
rect 114 -290 115 -258
rect 100 -297 101 -291
rect 187 -297 188 -291
rect 114 -297 115 -293
rect 142 -294 143 -258
rect 142 -297 143 -295
rect 247 -297 248 -295
rect 9 -307 10 -305
rect 61 -307 62 -305
rect 68 -338 69 -306
rect 72 -307 73 -305
rect 79 -338 80 -306
rect 89 -338 90 -306
rect 107 -307 108 -305
rect 215 -307 216 -305
rect 240 -307 241 -305
rect 317 -307 318 -305
rect 373 -338 374 -306
rect 376 -307 377 -305
rect 380 -307 381 -305
rect 387 -338 388 -306
rect 9 -338 10 -308
rect 37 -309 38 -305
rect 72 -338 73 -308
rect 86 -309 87 -305
rect 110 -338 111 -308
rect 170 -309 171 -305
rect 173 -338 174 -308
rect 191 -309 192 -305
rect 198 -338 199 -308
rect 240 -338 241 -308
rect 250 -309 251 -305
rect 338 -309 339 -305
rect 2 -311 3 -305
rect 86 -338 87 -310
rect 124 -311 125 -305
rect 149 -311 150 -305
rect 152 -338 153 -310
rect 226 -311 227 -305
rect 296 -338 297 -310
rect 299 -311 300 -305
rect 310 -311 311 -305
rect 369 -311 370 -305
rect 2 -338 3 -312
rect 156 -313 157 -305
rect 159 -313 160 -305
rect 303 -313 304 -305
rect 16 -315 17 -305
rect 166 -315 167 -305
rect 177 -315 178 -305
rect 177 -338 178 -314
rect 177 -315 178 -305
rect 177 -338 178 -314
rect 187 -315 188 -305
rect 359 -315 360 -305
rect 23 -317 24 -305
rect 124 -338 125 -316
rect 128 -317 129 -305
rect 184 -338 185 -316
rect 205 -338 206 -316
rect 324 -317 325 -305
rect 345 -317 346 -305
rect 359 -338 360 -316
rect 23 -338 24 -318
rect 82 -319 83 -305
rect 93 -319 94 -305
rect 156 -338 157 -318
rect 208 -319 209 -305
rect 352 -319 353 -305
rect 30 -321 31 -305
rect 135 -321 136 -305
rect 138 -321 139 -305
rect 233 -321 234 -305
rect 236 -321 237 -305
rect 310 -338 311 -320
rect 324 -338 325 -320
rect 331 -321 332 -305
rect 338 -338 339 -320
rect 352 -338 353 -320
rect 30 -338 31 -322
rect 142 -323 143 -305
rect 145 -338 146 -322
rect 247 -338 248 -322
rect 254 -323 255 -305
rect 331 -338 332 -322
rect 37 -338 38 -324
rect 114 -325 115 -305
rect 135 -338 136 -324
rect 243 -325 244 -305
rect 268 -325 269 -305
rect 345 -338 346 -324
rect 44 -327 45 -305
rect 142 -338 143 -326
rect 159 -338 160 -326
rect 254 -338 255 -326
rect 261 -327 262 -305
rect 268 -338 269 -326
rect 275 -327 276 -305
rect 303 -338 304 -326
rect 44 -338 45 -328
rect 51 -338 52 -328
rect 93 -338 94 -328
rect 117 -338 118 -328
rect 163 -329 164 -305
rect 261 -338 262 -328
rect 275 -338 276 -328
rect 289 -329 290 -305
rect 100 -331 101 -305
rect 128 -338 129 -330
rect 163 -338 164 -330
rect 201 -331 202 -305
rect 212 -331 213 -305
rect 317 -338 318 -330
rect 65 -333 66 -305
rect 100 -338 101 -332
rect 219 -333 220 -305
rect 226 -338 227 -332
rect 282 -333 283 -305
rect 289 -338 290 -332
rect 16 -338 17 -334
rect 65 -338 66 -334
rect 114 -338 115 -334
rect 219 -338 220 -334
rect 194 -338 195 -336
rect 282 -338 283 -336
rect 2 -348 3 -346
rect 145 -348 146 -346
rect 170 -348 171 -346
rect 366 -383 367 -347
rect 387 -348 388 -346
rect 387 -383 388 -347
rect 387 -348 388 -346
rect 387 -383 388 -347
rect 397 -383 398 -347
rect 401 -383 402 -347
rect 9 -350 10 -346
rect 44 -350 45 -346
rect 51 -350 52 -346
rect 51 -383 52 -349
rect 51 -350 52 -346
rect 51 -383 52 -349
rect 61 -350 62 -346
rect 187 -383 188 -349
rect 194 -350 195 -346
rect 289 -350 290 -346
rect 324 -350 325 -346
rect 324 -383 325 -349
rect 324 -350 325 -346
rect 324 -383 325 -349
rect 331 -350 332 -346
rect 338 -383 339 -349
rect 16 -352 17 -346
rect 96 -383 97 -351
rect 107 -352 108 -346
rect 107 -383 108 -351
rect 107 -352 108 -346
rect 107 -383 108 -351
rect 110 -352 111 -346
rect 226 -352 227 -346
rect 236 -352 237 -346
rect 268 -352 269 -346
rect 275 -352 276 -346
rect 275 -383 276 -351
rect 275 -352 276 -346
rect 275 -383 276 -351
rect 282 -352 283 -346
rect 380 -383 381 -351
rect 16 -383 17 -353
rect 72 -354 73 -346
rect 86 -383 87 -353
rect 117 -354 118 -346
rect 142 -354 143 -346
rect 142 -383 143 -353
rect 142 -354 143 -346
rect 142 -383 143 -353
rect 170 -383 171 -353
rect 373 -383 374 -353
rect 23 -356 24 -346
rect 114 -356 115 -346
rect 177 -356 178 -346
rect 191 -356 192 -346
rect 198 -356 199 -346
rect 212 -356 213 -346
rect 215 -383 216 -355
rect 233 -383 234 -355
rect 240 -356 241 -346
rect 345 -356 346 -346
rect 23 -383 24 -357
rect 100 -358 101 -346
rect 114 -383 115 -357
rect 184 -358 185 -346
rect 191 -383 192 -357
rect 257 -383 258 -357
rect 285 -383 286 -357
rect 359 -358 360 -346
rect 30 -360 31 -346
rect 159 -360 160 -346
rect 163 -360 164 -346
rect 177 -383 178 -359
rect 198 -383 199 -359
rect 243 -360 244 -346
rect 247 -360 248 -346
rect 345 -383 346 -359
rect 30 -383 31 -361
rect 65 -383 66 -361
rect 68 -383 69 -361
rect 89 -362 90 -346
rect 93 -362 94 -346
rect 121 -362 122 -346
rect 128 -362 129 -346
rect 163 -383 164 -361
rect 205 -362 206 -346
rect 289 -383 290 -361
rect 296 -362 297 -346
rect 359 -383 360 -361
rect 9 -383 10 -363
rect 89 -383 90 -363
rect 100 -383 101 -363
rect 149 -364 150 -346
rect 208 -364 209 -346
rect 331 -383 332 -363
rect 37 -366 38 -346
rect 173 -366 174 -346
rect 212 -383 213 -365
rect 317 -366 318 -346
rect 37 -383 38 -367
rect 135 -368 136 -346
rect 149 -383 150 -367
rect 352 -368 353 -346
rect 58 -383 59 -369
rect 128 -383 129 -369
rect 135 -383 136 -369
rect 152 -383 153 -369
rect 219 -370 220 -346
rect 226 -383 227 -369
rect 240 -383 241 -369
rect 317 -383 318 -369
rect 72 -383 73 -371
rect 93 -383 94 -371
rect 121 -383 122 -371
rect 145 -383 146 -371
rect 219 -383 220 -371
rect 296 -383 297 -371
rect 79 -374 80 -346
rect 205 -383 206 -373
rect 222 -383 223 -373
rect 303 -374 304 -346
rect 44 -383 45 -375
rect 79 -383 80 -375
rect 173 -383 174 -375
rect 303 -383 304 -375
rect 243 -383 244 -377
rect 310 -378 311 -346
rect 247 -383 248 -379
rect 254 -380 255 -346
rect 261 -380 262 -346
rect 310 -383 311 -379
rect 159 -383 160 -381
rect 261 -383 262 -381
rect 271 -383 272 -381
rect 352 -383 353 -381
rect 9 -393 10 -391
rect 159 -393 160 -391
rect 170 -393 171 -391
rect 205 -393 206 -391
rect 240 -393 241 -391
rect 275 -393 276 -391
rect 282 -422 283 -392
rect 324 -393 325 -391
rect 373 -393 374 -391
rect 373 -422 374 -392
rect 373 -393 374 -391
rect 373 -422 374 -392
rect 387 -393 388 -391
rect 394 -393 395 -391
rect 401 -393 402 -391
rect 411 -393 412 -391
rect 16 -395 17 -391
rect 117 -395 118 -391
rect 131 -395 132 -391
rect 173 -395 174 -391
rect 184 -395 185 -391
rect 208 -422 209 -394
rect 243 -395 244 -391
rect 243 -422 244 -394
rect 243 -395 244 -391
rect 243 -422 244 -394
rect 268 -395 269 -391
rect 310 -395 311 -391
rect 324 -422 325 -394
rect 366 -395 367 -391
rect 23 -397 24 -391
rect 149 -397 150 -391
rect 156 -397 157 -391
rect 177 -397 178 -391
rect 194 -397 195 -391
rect 198 -397 199 -391
rect 201 -422 202 -396
rect 219 -397 220 -391
rect 261 -397 262 -391
rect 268 -422 269 -396
rect 296 -397 297 -391
rect 366 -422 367 -396
rect 23 -422 24 -398
rect 93 -422 94 -398
rect 110 -422 111 -398
rect 177 -422 178 -398
rect 198 -422 199 -398
rect 226 -399 227 -391
rect 250 -422 251 -398
rect 261 -422 262 -398
rect 296 -422 297 -398
rect 380 -399 381 -391
rect 37 -401 38 -391
rect 128 -401 129 -391
rect 142 -401 143 -391
rect 247 -401 248 -391
rect 310 -422 311 -400
rect 352 -401 353 -391
rect 30 -403 31 -391
rect 37 -422 38 -402
rect 58 -403 59 -391
rect 58 -422 59 -402
rect 58 -403 59 -391
rect 58 -422 59 -402
rect 65 -403 66 -391
rect 117 -422 118 -402
rect 128 -422 129 -402
rect 135 -403 136 -391
rect 149 -422 150 -402
rect 222 -403 223 -391
rect 226 -422 227 -402
rect 257 -422 258 -402
rect 331 -403 332 -391
rect 380 -422 381 -402
rect 30 -422 31 -404
rect 51 -405 52 -391
rect 65 -422 66 -404
rect 233 -405 234 -391
rect 285 -405 286 -391
rect 331 -422 332 -404
rect 338 -405 339 -391
rect 352 -422 353 -404
rect 68 -422 69 -406
rect 275 -422 276 -406
rect 72 -409 73 -391
rect 215 -422 216 -408
rect 233 -422 234 -408
rect 303 -409 304 -391
rect 72 -422 73 -410
rect 121 -411 122 -391
rect 135 -422 136 -410
rect 170 -422 171 -410
rect 247 -422 248 -410
rect 338 -422 339 -410
rect 79 -413 80 -391
rect 89 -413 90 -391
rect 107 -413 108 -391
rect 142 -422 143 -412
rect 156 -422 157 -412
rect 219 -422 220 -412
rect 303 -422 304 -412
rect 345 -413 346 -391
rect 44 -415 45 -391
rect 79 -422 80 -414
rect 86 -422 87 -414
rect 100 -415 101 -391
rect 114 -415 115 -391
rect 285 -422 286 -414
rect 317 -415 318 -391
rect 345 -422 346 -414
rect 100 -422 101 -416
rect 145 -417 146 -391
rect 163 -417 164 -391
rect 184 -422 185 -416
rect 317 -422 318 -416
rect 359 -417 360 -391
rect 121 -422 122 -418
rect 159 -422 160 -418
rect 163 -422 164 -418
rect 212 -419 213 -391
rect 289 -419 290 -391
rect 359 -422 360 -418
rect 205 -422 206 -420
rect 289 -422 290 -420
rect 23 -432 24 -430
rect 47 -432 48 -430
rect 58 -432 59 -430
rect 58 -455 59 -431
rect 58 -432 59 -430
rect 58 -455 59 -431
rect 65 -432 66 -430
rect 100 -432 101 -430
rect 107 -455 108 -431
rect 128 -432 129 -430
rect 142 -432 143 -430
rect 145 -436 146 -431
rect 159 -432 160 -430
rect 184 -432 185 -430
rect 191 -432 192 -430
rect 233 -432 234 -430
rect 240 -455 241 -431
rect 268 -432 269 -430
rect 282 -432 283 -430
rect 282 -455 283 -431
rect 282 -432 283 -430
rect 282 -455 283 -431
rect 306 -455 307 -431
rect 310 -432 311 -430
rect 313 -455 314 -431
rect 338 -432 339 -430
rect 352 -432 353 -430
rect 373 -432 374 -430
rect 30 -434 31 -430
rect 68 -455 69 -433
rect 72 -434 73 -430
rect 131 -455 132 -433
rect 142 -455 143 -433
rect 149 -434 150 -430
rect 163 -455 164 -433
rect 212 -434 213 -430
rect 215 -434 216 -430
rect 317 -434 318 -430
rect 320 -455 321 -433
rect 345 -434 346 -430
rect 352 -455 353 -433
rect 366 -434 367 -430
rect 37 -455 38 -435
rect 124 -455 125 -435
rect 149 -455 150 -435
rect 170 -436 171 -430
rect 187 -455 188 -435
rect 215 -455 216 -435
rect 331 -436 332 -430
rect 359 -455 360 -435
rect 380 -436 381 -430
rect 44 -455 45 -437
rect 51 -438 52 -430
rect 79 -438 80 -430
rect 79 -455 80 -437
rect 79 -438 80 -430
rect 79 -455 80 -437
rect 86 -438 87 -430
rect 96 -438 97 -430
rect 114 -438 115 -430
rect 121 -438 122 -430
rect 170 -455 171 -437
rect 184 -455 185 -437
rect 226 -438 227 -430
rect 233 -455 234 -437
rect 247 -438 248 -430
rect 303 -438 304 -430
rect 362 -438 363 -430
rect 366 -455 367 -437
rect 51 -455 52 -439
rect 212 -455 213 -439
rect 229 -455 230 -439
rect 324 -440 325 -430
rect 65 -455 66 -441
rect 86 -455 87 -441
rect 93 -442 94 -430
rect 100 -455 101 -441
rect 177 -442 178 -430
rect 205 -442 206 -430
rect 254 -442 255 -430
rect 261 -442 262 -430
rect 268 -455 269 -441
rect 275 -442 276 -430
rect 303 -455 304 -441
rect 331 -455 332 -441
rect 75 -455 76 -443
rect 114 -455 115 -443
rect 117 -455 118 -443
rect 254 -455 255 -443
rect 275 -455 276 -443
rect 289 -444 290 -430
rect 93 -455 94 -445
rect 159 -455 160 -445
rect 198 -446 199 -430
rect 261 -455 262 -445
rect 289 -455 290 -445
rect 296 -446 297 -430
rect 135 -455 136 -447
rect 177 -455 178 -447
rect 191 -455 192 -447
rect 296 -455 297 -447
rect 194 -450 195 -430
rect 198 -455 199 -449
rect 205 -455 206 -449
rect 355 -450 356 -430
rect 194 -455 195 -451
rect 219 -452 220 -430
rect 156 -455 157 -453
rect 219 -455 220 -453
rect 26 -465 27 -463
rect 110 -492 111 -464
rect 121 -465 122 -463
rect 198 -465 199 -463
rect 212 -465 213 -463
rect 226 -465 227 -463
rect 250 -465 251 -463
rect 275 -465 276 -463
rect 296 -465 297 -463
rect 324 -492 325 -464
rect 338 -492 339 -464
rect 352 -465 353 -463
rect 366 -465 367 -463
rect 376 -465 377 -463
rect 33 -467 34 -463
rect 72 -467 73 -463
rect 79 -467 80 -463
rect 114 -467 115 -463
rect 121 -492 122 -466
rect 208 -492 209 -466
rect 215 -492 216 -466
rect 240 -467 241 -463
rect 254 -467 255 -463
rect 352 -492 353 -466
rect 37 -469 38 -463
rect 114 -492 115 -468
rect 142 -492 143 -468
rect 205 -469 206 -463
rect 240 -492 241 -468
rect 289 -469 290 -463
rect 317 -469 318 -463
rect 359 -469 360 -463
rect 37 -492 38 -470
rect 117 -471 118 -463
rect 149 -471 150 -463
rect 156 -492 157 -470
rect 177 -471 178 -463
rect 226 -492 227 -470
rect 261 -471 262 -463
rect 303 -492 304 -470
rect 331 -471 332 -463
rect 359 -492 360 -470
rect 44 -473 45 -463
rect 68 -492 69 -472
rect 72 -492 73 -472
rect 86 -473 87 -463
rect 93 -473 94 -463
rect 135 -473 136 -463
rect 177 -492 178 -472
rect 219 -473 220 -463
rect 275 -492 276 -472
rect 320 -492 321 -472
rect 331 -492 332 -472
rect 348 -492 349 -472
rect 44 -492 45 -474
rect 65 -492 66 -474
rect 86 -492 87 -474
rect 128 -475 129 -463
rect 135 -492 136 -474
rect 163 -475 164 -463
rect 184 -492 185 -474
rect 229 -475 230 -463
rect 282 -475 283 -463
rect 289 -492 290 -474
rect 58 -477 59 -463
rect 79 -492 80 -476
rect 107 -477 108 -463
rect 138 -477 139 -463
rect 163 -492 164 -476
rect 170 -477 171 -463
rect 187 -477 188 -463
rect 268 -477 269 -463
rect 51 -479 52 -463
rect 58 -492 59 -478
rect 128 -492 129 -478
rect 149 -492 150 -478
rect 170 -492 171 -478
rect 261 -492 262 -478
rect 51 -492 52 -480
rect 131 -481 132 -463
rect 173 -492 174 -480
rect 268 -492 269 -480
rect 100 -483 101 -463
rect 131 -492 132 -482
rect 191 -483 192 -463
rect 233 -483 234 -463
rect 100 -492 101 -484
rect 145 -485 146 -463
rect 194 -485 195 -463
rect 254 -492 255 -484
rect 198 -492 199 -486
rect 247 -492 248 -486
rect 205 -492 206 -488
rect 243 -492 244 -488
rect 233 -492 234 -490
rect 306 -491 307 -463
rect 16 -531 17 -501
rect 107 -502 108 -500
rect 156 -502 157 -500
rect 173 -502 174 -500
rect 177 -502 178 -500
rect 194 -502 195 -500
rect 201 -502 202 -500
rect 205 -531 206 -501
rect 212 -502 213 -500
rect 212 -531 213 -501
rect 212 -502 213 -500
rect 212 -531 213 -501
rect 222 -531 223 -501
rect 299 -502 300 -500
rect 338 -531 339 -501
rect 359 -531 360 -501
rect 30 -531 31 -503
rect 44 -504 45 -500
rect 51 -504 52 -500
rect 243 -504 244 -500
rect 254 -504 255 -500
rect 254 -531 255 -503
rect 254 -504 255 -500
rect 254 -531 255 -503
rect 268 -504 269 -500
rect 313 -504 314 -500
rect 345 -531 346 -503
rect 348 -504 349 -500
rect 352 -504 353 -500
rect 373 -531 374 -503
rect 65 -506 66 -500
rect 79 -506 80 -500
rect 86 -506 87 -500
rect 93 -506 94 -500
rect 110 -506 111 -500
rect 156 -531 157 -505
rect 159 -531 160 -505
rect 226 -506 227 -500
rect 275 -506 276 -500
rect 296 -506 297 -500
rect 317 -531 318 -505
rect 348 -531 349 -505
rect 51 -531 52 -507
rect 93 -531 94 -507
rect 163 -508 164 -500
rect 198 -508 199 -500
rect 226 -531 227 -507
rect 289 -508 290 -500
rect 296 -531 297 -507
rect 331 -508 332 -500
rect 341 -508 342 -500
rect 352 -531 353 -507
rect 44 -531 45 -509
rect 198 -531 199 -509
rect 208 -531 209 -509
rect 331 -531 332 -509
rect 341 -531 342 -509
rect 366 -531 367 -509
rect 65 -531 66 -511
rect 142 -512 143 -500
rect 149 -512 150 -500
rect 163 -531 164 -511
rect 166 -531 167 -511
rect 310 -531 311 -511
rect 68 -514 69 -500
rect 110 -531 111 -513
rect 170 -531 171 -513
rect 240 -514 241 -500
rect 282 -514 283 -500
rect 324 -514 325 -500
rect 72 -516 73 -500
rect 131 -531 132 -515
rect 191 -531 192 -515
rect 219 -516 220 -500
rect 233 -516 234 -500
rect 240 -531 241 -515
rect 247 -516 248 -500
rect 282 -531 283 -515
rect 289 -531 290 -515
rect 303 -516 304 -500
rect 37 -518 38 -500
rect 72 -531 73 -517
rect 79 -531 80 -517
rect 149 -531 150 -517
rect 194 -531 195 -517
rect 247 -531 248 -517
rect 261 -518 262 -500
rect 324 -531 325 -517
rect 37 -531 38 -519
rect 58 -520 59 -500
rect 86 -531 87 -519
rect 100 -520 101 -500
rect 114 -520 115 -500
rect 219 -531 220 -519
rect 229 -531 230 -519
rect 303 -531 304 -519
rect 58 -531 59 -521
rect 121 -522 122 -500
rect 142 -531 143 -521
rect 233 -531 234 -521
rect 100 -531 101 -523
rect 268 -531 269 -523
rect 114 -531 115 -525
rect 135 -526 136 -500
rect 201 -531 202 -525
rect 261 -531 262 -525
rect 135 -531 136 -527
rect 184 -528 185 -500
rect 177 -531 178 -529
rect 184 -531 185 -529
rect 9 -570 10 -540
rect 107 -570 108 -540
rect 121 -570 122 -540
rect 149 -541 150 -539
rect 156 -541 157 -539
rect 219 -570 220 -540
rect 222 -541 223 -539
rect 331 -541 332 -539
rect 338 -541 339 -539
rect 373 -541 374 -539
rect 16 -543 17 -539
rect 229 -543 230 -539
rect 275 -543 276 -539
rect 289 -543 290 -539
rect 296 -543 297 -539
rect 296 -570 297 -542
rect 296 -543 297 -539
rect 296 -570 297 -542
rect 348 -543 349 -539
rect 352 -543 353 -539
rect 359 -543 360 -539
rect 359 -570 360 -542
rect 359 -543 360 -539
rect 359 -570 360 -542
rect 16 -570 17 -544
rect 51 -545 52 -539
rect 58 -545 59 -539
rect 166 -545 167 -539
rect 177 -545 178 -539
rect 205 -545 206 -539
rect 208 -545 209 -539
rect 289 -570 290 -544
rect 23 -570 24 -546
rect 26 -547 27 -539
rect 37 -547 38 -539
rect 82 -570 83 -546
rect 86 -547 87 -539
rect 103 -547 104 -539
rect 131 -547 132 -539
rect 345 -547 346 -539
rect 44 -549 45 -539
rect 124 -549 125 -539
rect 142 -570 143 -548
rect 205 -570 206 -548
rect 226 -570 227 -548
rect 261 -549 262 -539
rect 275 -570 276 -548
rect 366 -549 367 -539
rect 30 -551 31 -539
rect 44 -570 45 -550
rect 58 -570 59 -550
rect 79 -551 80 -539
rect 86 -570 87 -550
rect 110 -551 111 -539
rect 114 -551 115 -539
rect 131 -570 132 -550
rect 145 -551 146 -539
rect 247 -551 248 -539
rect 254 -551 255 -539
rect 261 -570 262 -550
rect 65 -553 66 -539
rect 152 -553 153 -539
rect 177 -570 178 -552
rect 236 -570 237 -552
rect 247 -570 248 -552
rect 278 -553 279 -539
rect 65 -570 66 -554
rect 159 -570 160 -554
rect 191 -570 192 -554
rect 233 -555 234 -539
rect 268 -555 269 -539
rect 278 -570 279 -554
rect 72 -570 73 -556
rect 135 -557 136 -539
rect 201 -557 202 -539
rect 282 -557 283 -539
rect 93 -559 94 -539
rect 240 -559 241 -539
rect 268 -570 269 -558
rect 324 -559 325 -539
rect 93 -570 94 -560
rect 145 -570 146 -560
rect 240 -570 241 -560
rect 303 -561 304 -539
rect 317 -561 318 -539
rect 324 -570 325 -560
rect 100 -563 101 -539
rect 198 -563 199 -539
rect 282 -570 283 -562
rect 292 -570 293 -562
rect 303 -570 304 -562
rect 310 -563 311 -539
rect 100 -570 101 -564
rect 128 -565 129 -539
rect 135 -570 136 -564
rect 152 -570 153 -564
rect 198 -570 199 -564
rect 212 -565 213 -539
rect 114 -570 115 -566
rect 124 -570 125 -566
rect 170 -567 171 -539
rect 212 -570 213 -566
rect 163 -570 164 -568
rect 170 -570 171 -568
rect 9 -580 10 -578
rect 156 -601 157 -579
rect 159 -580 160 -578
rect 198 -580 199 -578
rect 205 -580 206 -578
rect 233 -601 234 -579
rect 257 -580 258 -578
rect 261 -580 262 -578
rect 282 -580 283 -578
rect 310 -580 311 -578
rect 324 -580 325 -578
rect 324 -601 325 -579
rect 324 -580 325 -578
rect 324 -601 325 -579
rect 355 -580 356 -578
rect 359 -580 360 -578
rect 16 -582 17 -578
rect 51 -582 52 -578
rect 65 -582 66 -578
rect 96 -601 97 -581
rect 100 -582 101 -578
rect 110 -582 111 -578
rect 135 -582 136 -578
rect 142 -601 143 -581
rect 187 -582 188 -578
rect 191 -582 192 -578
rect 198 -601 199 -581
rect 219 -582 220 -578
rect 226 -582 227 -578
rect 254 -601 255 -581
rect 261 -601 262 -581
rect 268 -582 269 -578
rect 282 -601 283 -581
rect 306 -601 307 -581
rect 23 -584 24 -578
rect 23 -601 24 -583
rect 23 -584 24 -578
rect 23 -601 24 -583
rect 30 -601 31 -583
rect 82 -584 83 -578
rect 86 -584 87 -578
rect 145 -584 146 -578
rect 163 -584 164 -578
rect 191 -601 192 -583
rect 205 -601 206 -583
rect 229 -601 230 -583
rect 268 -601 269 -583
rect 278 -601 279 -583
rect 289 -601 290 -583
rect 303 -584 304 -578
rect 40 -586 41 -578
rect 40 -601 41 -585
rect 40 -586 41 -578
rect 40 -601 41 -585
rect 44 -586 45 -578
rect 44 -601 45 -585
rect 44 -586 45 -578
rect 44 -601 45 -585
rect 51 -601 52 -585
rect 131 -586 132 -578
rect 135 -601 136 -585
rect 138 -601 139 -585
rect 163 -601 164 -585
rect 184 -601 185 -585
rect 219 -601 220 -585
rect 240 -586 241 -578
rect 296 -586 297 -578
rect 303 -601 304 -585
rect 58 -588 59 -578
rect 65 -601 66 -587
rect 72 -588 73 -578
rect 152 -588 153 -578
rect 177 -588 178 -578
rect 187 -601 188 -587
rect 58 -601 59 -589
rect 100 -601 101 -589
rect 152 -601 153 -589
rect 212 -590 213 -578
rect 75 -601 76 -591
rect 128 -601 129 -591
rect 170 -601 171 -591
rect 177 -601 178 -591
rect 212 -601 213 -591
rect 247 -592 248 -578
rect 86 -601 87 -593
rect 114 -594 115 -578
rect 159 -601 160 -593
rect 247 -601 248 -593
rect 93 -596 94 -578
rect 107 -596 108 -578
rect 114 -601 115 -595
rect 121 -601 122 -595
rect 79 -598 80 -578
rect 93 -601 94 -597
rect 107 -601 108 -597
rect 149 -601 150 -597
rect 33 -600 34 -578
rect 79 -601 80 -599
rect 26 -611 27 -609
rect 26 -626 27 -610
rect 26 -611 27 -609
rect 26 -626 27 -610
rect 30 -611 31 -609
rect 82 -611 83 -609
rect 100 -611 101 -609
rect 103 -626 104 -610
rect 114 -611 115 -609
rect 128 -626 129 -610
rect 131 -611 132 -609
rect 149 -611 150 -609
rect 156 -611 157 -609
rect 180 -611 181 -609
rect 184 -626 185 -610
rect 212 -611 213 -609
rect 226 -611 227 -609
rect 254 -611 255 -609
rect 257 -626 258 -610
rect 282 -611 283 -609
rect 324 -611 325 -609
rect 324 -626 325 -610
rect 324 -611 325 -609
rect 324 -626 325 -610
rect 37 -613 38 -609
rect 44 -613 45 -609
rect 51 -613 52 -609
rect 117 -613 118 -609
rect 135 -613 136 -609
rect 191 -613 192 -609
rect 205 -613 206 -609
rect 226 -626 227 -612
rect 233 -613 234 -609
rect 264 -626 265 -612
rect 275 -613 276 -609
rect 289 -613 290 -609
rect 51 -626 52 -614
rect 72 -626 73 -614
rect 86 -615 87 -609
rect 117 -626 118 -614
rect 135 -626 136 -614
rect 142 -615 143 -609
rect 159 -615 160 -609
rect 198 -615 199 -609
rect 205 -626 206 -614
rect 219 -615 220 -609
rect 233 -626 234 -614
rect 261 -615 262 -609
rect 58 -617 59 -609
rect 138 -617 139 -609
rect 142 -626 143 -616
rect 156 -626 157 -616
rect 163 -617 164 -609
rect 173 -626 174 -616
rect 177 -617 178 -609
rect 180 -626 181 -616
rect 187 -626 188 -616
rect 212 -626 213 -616
rect 240 -626 241 -616
rect 247 -617 248 -609
rect 261 -626 262 -616
rect 268 -617 269 -609
rect 65 -619 66 -609
rect 86 -626 87 -618
rect 114 -626 115 -618
rect 145 -626 146 -618
rect 152 -619 153 -609
rect 219 -626 220 -618
rect 243 -619 244 -609
rect 247 -626 248 -618
rect 65 -626 66 -620
rect 107 -621 108 -609
rect 121 -621 122 -609
rect 163 -626 164 -620
rect 170 -621 171 -609
rect 198 -626 199 -620
rect 79 -623 80 -609
rect 121 -626 122 -622
rect 191 -626 192 -622
rect 254 -626 255 -622
rect 75 -625 76 -609
rect 79 -626 80 -624
rect 93 -626 94 -624
rect 107 -626 108 -624
rect 30 -659 31 -635
rect 51 -636 52 -634
rect 65 -636 66 -634
rect 107 -636 108 -634
rect 121 -636 122 -634
rect 149 -636 150 -634
rect 152 -636 153 -634
rect 191 -636 192 -634
rect 201 -659 202 -635
rect 268 -659 269 -635
rect 37 -659 38 -637
rect 72 -659 73 -637
rect 82 -638 83 -634
rect 100 -638 101 -634
rect 107 -659 108 -637
rect 117 -659 118 -637
rect 124 -659 125 -637
rect 163 -638 164 -634
rect 184 -659 185 -637
rect 240 -638 241 -634
rect 247 -638 248 -634
rect 289 -659 290 -637
rect 44 -659 45 -639
rect 75 -640 76 -634
rect 96 -659 97 -639
rect 233 -640 234 -634
rect 254 -659 255 -639
rect 257 -640 258 -634
rect 51 -659 52 -641
rect 93 -642 94 -634
rect 100 -659 101 -641
rect 121 -659 122 -641
rect 135 -642 136 -634
rect 145 -642 146 -634
rect 149 -659 150 -641
rect 187 -642 188 -634
rect 205 -642 206 -634
rect 233 -659 234 -641
rect 68 -659 69 -643
rect 79 -659 80 -643
rect 128 -644 129 -634
rect 135 -659 136 -643
rect 142 -659 143 -643
rect 261 -659 262 -643
rect 75 -659 76 -645
rect 86 -659 87 -645
rect 128 -659 129 -645
rect 138 -659 139 -645
rect 156 -646 157 -634
rect 173 -659 174 -645
rect 187 -659 188 -645
rect 296 -659 297 -645
rect 156 -659 157 -647
rect 163 -659 164 -647
rect 170 -659 171 -647
rect 247 -659 248 -647
rect 212 -650 213 -634
rect 240 -659 241 -649
rect 198 -652 199 -634
rect 212 -659 213 -651
rect 219 -652 220 -634
rect 282 -659 283 -651
rect 219 -659 220 -653
rect 236 -654 237 -634
rect 226 -656 227 -634
rect 275 -659 276 -655
rect 191 -659 192 -657
rect 226 -659 227 -657
rect 37 -669 38 -667
rect 110 -692 111 -668
rect 114 -669 115 -667
rect 142 -692 143 -668
rect 156 -669 157 -667
rect 226 -669 227 -667
rect 254 -669 255 -667
rect 278 -692 279 -668
rect 44 -671 45 -667
rect 145 -671 146 -667
rect 156 -692 157 -670
rect 163 -671 164 -667
rect 173 -671 174 -667
rect 268 -671 269 -667
rect 51 -673 52 -667
rect 117 -673 118 -667
rect 121 -692 122 -672
rect 191 -673 192 -667
rect 198 -692 199 -672
rect 212 -673 213 -667
rect 247 -673 248 -667
rect 254 -692 255 -672
rect 261 -673 262 -667
rect 268 -692 269 -672
rect 58 -675 59 -667
rect 86 -675 87 -667
rect 89 -692 90 -674
rect 138 -675 139 -667
rect 159 -675 160 -667
rect 201 -675 202 -667
rect 205 -675 206 -667
rect 205 -692 206 -674
rect 205 -675 206 -667
rect 205 -692 206 -674
rect 208 -675 209 -667
rect 275 -675 276 -667
rect 61 -677 62 -667
rect 68 -677 69 -667
rect 79 -677 80 -667
rect 79 -692 80 -676
rect 79 -677 80 -667
rect 79 -692 80 -676
rect 93 -677 94 -667
rect 184 -677 185 -667
rect 187 -692 188 -676
rect 233 -677 234 -667
rect 30 -679 31 -667
rect 61 -692 62 -678
rect 93 -692 94 -678
rect 149 -679 150 -667
rect 180 -679 181 -667
rect 282 -679 283 -667
rect 96 -681 97 -667
rect 100 -681 101 -667
rect 128 -681 129 -667
rect 128 -692 129 -680
rect 128 -681 129 -667
rect 128 -692 129 -680
rect 138 -692 139 -680
rect 163 -692 164 -680
rect 180 -692 181 -680
rect 289 -681 290 -667
rect 100 -692 101 -682
rect 107 -683 108 -667
rect 191 -692 192 -682
rect 226 -692 227 -682
rect 107 -692 108 -684
rect 170 -692 171 -684
rect 212 -692 213 -684
rect 240 -685 241 -667
rect 177 -687 178 -667
rect 240 -692 241 -686
rect 219 -689 220 -667
rect 233 -692 234 -688
rect 177 -692 178 -690
rect 219 -692 220 -690
rect 61 -702 62 -700
rect 72 -702 73 -700
rect 75 -702 76 -700
rect 79 -702 80 -700
rect 100 -702 101 -700
rect 117 -702 118 -700
rect 121 -702 122 -700
rect 177 -702 178 -700
rect 184 -715 185 -701
rect 226 -702 227 -700
rect 240 -702 241 -700
rect 261 -702 262 -700
rect 114 -704 115 -700
rect 121 -715 122 -703
rect 128 -704 129 -700
rect 135 -715 136 -703
rect 142 -704 143 -700
rect 187 -704 188 -700
rect 194 -704 195 -700
rect 198 -704 199 -700
rect 240 -715 241 -703
rect 254 -704 255 -700
rect 131 -715 132 -705
rect 142 -715 143 -705
rect 149 -715 150 -705
rect 170 -706 171 -700
rect 194 -715 195 -705
rect 219 -706 220 -700
rect 247 -706 248 -700
rect 268 -706 269 -700
rect 93 -708 94 -700
rect 170 -715 171 -707
rect 198 -715 199 -707
rect 233 -708 234 -700
rect 152 -710 153 -700
rect 205 -710 206 -700
rect 163 -712 164 -700
rect 173 -715 174 -711
rect 205 -715 206 -711
rect 215 -715 216 -711
rect 163 -715 164 -713
rect 180 -715 181 -713
rect 114 -725 115 -723
rect 131 -725 132 -723
rect 135 -730 136 -724
rect 142 -725 143 -723
rect 159 -730 160 -724
rect 177 -725 178 -723
rect 180 -725 181 -723
rect 184 -725 185 -723
rect 191 -725 192 -723
rect 205 -725 206 -723
rect 229 -725 230 -723
rect 240 -725 241 -723
rect 121 -727 122 -723
rect 131 -730 132 -726
rect 163 -727 164 -723
rect 170 -730 171 -726
rect 173 -727 174 -723
rect 198 -727 199 -723
rect 117 -730 118 -728
rect 121 -730 122 -728
rect 177 -730 178 -728
rect 184 -730 185 -728
rect 191 -730 192 -728
rect 194 -729 195 -723
rect 128 -740 129 -738
rect 135 -740 136 -738
rect 149 -743 150 -739
rect 163 -743 164 -739
rect 166 -740 167 -738
rect 170 -740 171 -738
rect 177 -740 178 -738
rect 184 -743 185 -739
rect 187 -740 188 -738
rect 191 -740 192 -738
rect 121 -742 122 -738
rect 128 -743 129 -741
rect 156 -742 157 -738
rect 170 -743 171 -741
rect 124 -753 125 -751
rect 128 -753 129 -751
rect 156 -753 157 -751
rect 170 -753 171 -751
rect 184 -753 185 -751
rect 191 -753 192 -751
rect 159 -755 160 -751
rect 163 -755 164 -751
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=16
rlabel pdiffusion 10 -8 10 -8 0 cellNo=108
rlabel pdiffusion 17 -8 17 -8 0 cellNo=42
rlabel pdiffusion 24 -8 24 -8 0 cellNo=312
rlabel pdiffusion 31 -8 31 -8 0 cellNo=128
rlabel pdiffusion 38 -8 38 -8 0 cellNo=253
rlabel pdiffusion 45 -8 45 -8 0 cellNo=369
rlabel pdiffusion 101 -8 101 -8 0 cellNo=3
rlabel pdiffusion 108 -8 108 -8 0 cellNo=186
rlabel pdiffusion 129 -8 129 -8 0 cellNo=225
rlabel pdiffusion 136 -8 136 -8 0 feedthrough
rlabel pdiffusion 143 -8 143 -8 0 cellNo=266
rlabel pdiffusion 150 -8 150 -8 0 cellNo=176
rlabel pdiffusion 157 -8 157 -8 0 feedthrough
rlabel pdiffusion 164 -8 164 -8 0 cellNo=180
rlabel pdiffusion 171 -8 171 -8 0 cellNo=33
rlabel pdiffusion 178 -8 178 -8 0 feedthrough
rlabel pdiffusion 185 -8 185 -8 0 cellNo=170
rlabel pdiffusion 192 -8 192 -8 0 cellNo=56
rlabel pdiffusion 199 -8 199 -8 0 feedthrough
rlabel pdiffusion 206 -8 206 -8 0 cellNo=88
rlabel pdiffusion 213 -8 213 -8 0 feedthrough
rlabel pdiffusion 3 -27 3 -27 0 cellNo=116
rlabel pdiffusion 10 -27 10 -27 0 cellNo=375
rlabel pdiffusion 17 -27 17 -27 0 cellNo=360
rlabel pdiffusion 24 -27 24 -27 0 cellNo=209
rlabel pdiffusion 31 -27 31 -27 0 cellNo=241
rlabel pdiffusion 38 -27 38 -27 0 cellNo=362
rlabel pdiffusion 80 -27 80 -27 0 feedthrough
rlabel pdiffusion 87 -27 87 -27 0 cellNo=198
rlabel pdiffusion 94 -27 94 -27 0 cellNo=284
rlabel pdiffusion 101 -27 101 -27 0 cellNo=244
rlabel pdiffusion 108 -27 108 -27 0 cellNo=257
rlabel pdiffusion 122 -27 122 -27 0 feedthrough
rlabel pdiffusion 129 -27 129 -27 0 cellNo=95
rlabel pdiffusion 136 -27 136 -27 0 feedthrough
rlabel pdiffusion 143 -27 143 -27 0 feedthrough
rlabel pdiffusion 150 -27 150 -27 0 cellNo=262
rlabel pdiffusion 157 -27 157 -27 0 cellNo=287
rlabel pdiffusion 164 -27 164 -27 0 cellNo=14
rlabel pdiffusion 171 -27 171 -27 0 feedthrough
rlabel pdiffusion 178 -27 178 -27 0 cellNo=219
rlabel pdiffusion 185 -27 185 -27 0 cellNo=222
rlabel pdiffusion 192 -27 192 -27 0 cellNo=227
rlabel pdiffusion 199 -27 199 -27 0 feedthrough
rlabel pdiffusion 206 -27 206 -27 0 cellNo=8
rlabel pdiffusion 213 -27 213 -27 0 cellNo=140
rlabel pdiffusion 220 -27 220 -27 0 feedthrough
rlabel pdiffusion 227 -27 227 -27 0 cellNo=207
rlabel pdiffusion 234 -27 234 -27 0 feedthrough
rlabel pdiffusion 3 -50 3 -50 0 cellNo=47
rlabel pdiffusion 10 -50 10 -50 0 cellNo=102
rlabel pdiffusion 17 -50 17 -50 0 cellNo=148
rlabel pdiffusion 24 -50 24 -50 0 cellNo=235
rlabel pdiffusion 31 -50 31 -50 0 cellNo=392
rlabel pdiffusion 59 -50 59 -50 0 cellNo=57
rlabel pdiffusion 66 -50 66 -50 0 feedthrough
rlabel pdiffusion 73 -50 73 -50 0 feedthrough
rlabel pdiffusion 80 -50 80 -50 0 cellNo=194
rlabel pdiffusion 87 -50 87 -50 0 cellNo=161
rlabel pdiffusion 94 -50 94 -50 0 cellNo=67
rlabel pdiffusion 101 -50 101 -50 0 feedthrough
rlabel pdiffusion 108 -50 108 -50 0 cellNo=6
rlabel pdiffusion 115 -50 115 -50 0 feedthrough
rlabel pdiffusion 122 -50 122 -50 0 cellNo=177
rlabel pdiffusion 129 -50 129 -50 0 cellNo=35
rlabel pdiffusion 136 -50 136 -50 0 feedthrough
rlabel pdiffusion 143 -50 143 -50 0 cellNo=43
rlabel pdiffusion 150 -50 150 -50 0 cellNo=25
rlabel pdiffusion 157 -50 157 -50 0 feedthrough
rlabel pdiffusion 164 -50 164 -50 0 feedthrough
rlabel pdiffusion 171 -50 171 -50 0 cellNo=228
rlabel pdiffusion 178 -50 178 -50 0 cellNo=359
rlabel pdiffusion 185 -50 185 -50 0 feedthrough
rlabel pdiffusion 192 -50 192 -50 0 feedthrough
rlabel pdiffusion 199 -50 199 -50 0 cellNo=19
rlabel pdiffusion 206 -50 206 -50 0 feedthrough
rlabel pdiffusion 213 -50 213 -50 0 cellNo=32
rlabel pdiffusion 220 -50 220 -50 0 cellNo=398
rlabel pdiffusion 227 -50 227 -50 0 feedthrough
rlabel pdiffusion 234 -50 234 -50 0 feedthrough
rlabel pdiffusion 241 -50 241 -50 0 feedthrough
rlabel pdiffusion 248 -50 248 -50 0 feedthrough
rlabel pdiffusion 255 -50 255 -50 0 feedthrough
rlabel pdiffusion 262 -50 262 -50 0 feedthrough
rlabel pdiffusion 269 -50 269 -50 0 cellNo=62
rlabel pdiffusion 276 -50 276 -50 0 feedthrough
rlabel pdiffusion 283 -50 283 -50 0 feedthrough
rlabel pdiffusion 3 -81 3 -81 0 cellNo=92
rlabel pdiffusion 10 -81 10 -81 0 cellNo=169
rlabel pdiffusion 17 -81 17 -81 0 cellNo=231
rlabel pdiffusion 24 -81 24 -81 0 cellNo=351
rlabel pdiffusion 31 -81 31 -81 0 feedthrough
rlabel pdiffusion 38 -81 38 -81 0 cellNo=237
rlabel pdiffusion 45 -81 45 -81 0 feedthrough
rlabel pdiffusion 52 -81 52 -81 0 feedthrough
rlabel pdiffusion 59 -81 59 -81 0 feedthrough
rlabel pdiffusion 66 -81 66 -81 0 feedthrough
rlabel pdiffusion 73 -81 73 -81 0 cellNo=164
rlabel pdiffusion 80 -81 80 -81 0 feedthrough
rlabel pdiffusion 87 -81 87 -81 0 feedthrough
rlabel pdiffusion 94 -81 94 -81 0 feedthrough
rlabel pdiffusion 101 -81 101 -81 0 cellNo=166
rlabel pdiffusion 108 -81 108 -81 0 cellNo=22
rlabel pdiffusion 115 -81 115 -81 0 cellNo=188
rlabel pdiffusion 122 -81 122 -81 0 feedthrough
rlabel pdiffusion 129 -81 129 -81 0 cellNo=320
rlabel pdiffusion 136 -81 136 -81 0 cellNo=356
rlabel pdiffusion 143 -81 143 -81 0 feedthrough
rlabel pdiffusion 150 -81 150 -81 0 feedthrough
rlabel pdiffusion 157 -81 157 -81 0 cellNo=114
rlabel pdiffusion 164 -81 164 -81 0 feedthrough
rlabel pdiffusion 171 -81 171 -81 0 feedthrough
rlabel pdiffusion 178 -81 178 -81 0 cellNo=91
rlabel pdiffusion 185 -81 185 -81 0 cellNo=126
rlabel pdiffusion 192 -81 192 -81 0 feedthrough
rlabel pdiffusion 199 -81 199 -81 0 cellNo=201
rlabel pdiffusion 206 -81 206 -81 0 cellNo=23
rlabel pdiffusion 213 -81 213 -81 0 cellNo=68
rlabel pdiffusion 220 -81 220 -81 0 feedthrough
rlabel pdiffusion 227 -81 227 -81 0 feedthrough
rlabel pdiffusion 234 -81 234 -81 0 feedthrough
rlabel pdiffusion 241 -81 241 -81 0 cellNo=310
rlabel pdiffusion 248 -81 248 -81 0 cellNo=291
rlabel pdiffusion 255 -81 255 -81 0 feedthrough
rlabel pdiffusion 262 -81 262 -81 0 feedthrough
rlabel pdiffusion 269 -81 269 -81 0 feedthrough
rlabel pdiffusion 276 -81 276 -81 0 feedthrough
rlabel pdiffusion 283 -81 283 -81 0 feedthrough
rlabel pdiffusion 290 -81 290 -81 0 feedthrough
rlabel pdiffusion 297 -81 297 -81 0 cellNo=196
rlabel pdiffusion 304 -81 304 -81 0 feedthrough
rlabel pdiffusion 3 -126 3 -126 0 cellNo=118
rlabel pdiffusion 10 -126 10 -126 0 cellNo=165
rlabel pdiffusion 17 -126 17 -126 0 feedthrough
rlabel pdiffusion 24 -126 24 -126 0 cellNo=26
rlabel pdiffusion 31 -126 31 -126 0 feedthrough
rlabel pdiffusion 38 -126 38 -126 0 feedthrough
rlabel pdiffusion 45 -126 45 -126 0 cellNo=343
rlabel pdiffusion 52 -126 52 -126 0 feedthrough
rlabel pdiffusion 59 -126 59 -126 0 cellNo=365
rlabel pdiffusion 66 -126 66 -126 0 cellNo=232
rlabel pdiffusion 73 -126 73 -126 0 feedthrough
rlabel pdiffusion 80 -126 80 -126 0 cellNo=107
rlabel pdiffusion 87 -126 87 -126 0 feedthrough
rlabel pdiffusion 94 -126 94 -126 0 feedthrough
rlabel pdiffusion 101 -126 101 -126 0 cellNo=82
rlabel pdiffusion 108 -126 108 -126 0 feedthrough
rlabel pdiffusion 115 -126 115 -126 0 cellNo=200
rlabel pdiffusion 122 -126 122 -126 0 cellNo=289
rlabel pdiffusion 129 -126 129 -126 0 cellNo=213
rlabel pdiffusion 136 -126 136 -126 0 cellNo=36
rlabel pdiffusion 143 -126 143 -126 0 cellNo=285
rlabel pdiffusion 150 -126 150 -126 0 cellNo=84
rlabel pdiffusion 157 -126 157 -126 0 cellNo=55
rlabel pdiffusion 164 -126 164 -126 0 cellNo=324
rlabel pdiffusion 171 -126 171 -126 0 feedthrough
rlabel pdiffusion 178 -126 178 -126 0 cellNo=238
rlabel pdiffusion 185 -126 185 -126 0 cellNo=283
rlabel pdiffusion 192 -126 192 -126 0 cellNo=77
rlabel pdiffusion 199 -126 199 -126 0 cellNo=304
rlabel pdiffusion 206 -126 206 -126 0 cellNo=256
rlabel pdiffusion 213 -126 213 -126 0 feedthrough
rlabel pdiffusion 220 -126 220 -126 0 feedthrough
rlabel pdiffusion 227 -126 227 -126 0 feedthrough
rlabel pdiffusion 234 -126 234 -126 0 cellNo=141
rlabel pdiffusion 241 -126 241 -126 0 feedthrough
rlabel pdiffusion 248 -126 248 -126 0 feedthrough
rlabel pdiffusion 255 -126 255 -126 0 feedthrough
rlabel pdiffusion 262 -126 262 -126 0 feedthrough
rlabel pdiffusion 269 -126 269 -126 0 feedthrough
rlabel pdiffusion 276 -126 276 -126 0 feedthrough
rlabel pdiffusion 283 -126 283 -126 0 feedthrough
rlabel pdiffusion 290 -126 290 -126 0 feedthrough
rlabel pdiffusion 297 -126 297 -126 0 feedthrough
rlabel pdiffusion 304 -126 304 -126 0 feedthrough
rlabel pdiffusion 311 -126 311 -126 0 feedthrough
rlabel pdiffusion 318 -126 318 -126 0 feedthrough
rlabel pdiffusion 325 -126 325 -126 0 feedthrough
rlabel pdiffusion 332 -126 332 -126 0 feedthrough
rlabel pdiffusion 3 -173 3 -173 0 cellNo=131
rlabel pdiffusion 10 -173 10 -173 0 cellNo=295
rlabel pdiffusion 17 -173 17 -173 0 cellNo=172
rlabel pdiffusion 24 -173 24 -173 0 cellNo=316
rlabel pdiffusion 31 -173 31 -173 0 feedthrough
rlabel pdiffusion 38 -173 38 -173 0 cellNo=119
rlabel pdiffusion 45 -173 45 -173 0 feedthrough
rlabel pdiffusion 52 -173 52 -173 0 cellNo=129
rlabel pdiffusion 59 -173 59 -173 0 cellNo=7
rlabel pdiffusion 66 -173 66 -173 0 feedthrough
rlabel pdiffusion 73 -173 73 -173 0 feedthrough
rlabel pdiffusion 80 -173 80 -173 0 feedthrough
rlabel pdiffusion 87 -173 87 -173 0 cellNo=74
rlabel pdiffusion 94 -173 94 -173 0 feedthrough
rlabel pdiffusion 101 -173 101 -173 0 feedthrough
rlabel pdiffusion 108 -173 108 -173 0 cellNo=217
rlabel pdiffusion 115 -173 115 -173 0 cellNo=147
rlabel pdiffusion 122 -173 122 -173 0 cellNo=31
rlabel pdiffusion 129 -173 129 -173 0 feedthrough
rlabel pdiffusion 136 -173 136 -173 0 cellNo=355
rlabel pdiffusion 143 -173 143 -173 0 feedthrough
rlabel pdiffusion 150 -173 150 -173 0 cellNo=366
rlabel pdiffusion 157 -173 157 -173 0 cellNo=44
rlabel pdiffusion 164 -173 164 -173 0 cellNo=97
rlabel pdiffusion 171 -173 171 -173 0 feedthrough
rlabel pdiffusion 178 -173 178 -173 0 feedthrough
rlabel pdiffusion 185 -173 185 -173 0 feedthrough
rlabel pdiffusion 192 -173 192 -173 0 cellNo=38
rlabel pdiffusion 199 -173 199 -173 0 cellNo=294
rlabel pdiffusion 206 -173 206 -173 0 cellNo=151
rlabel pdiffusion 213 -173 213 -173 0 cellNo=60
rlabel pdiffusion 220 -173 220 -173 0 feedthrough
rlabel pdiffusion 227 -173 227 -173 0 feedthrough
rlabel pdiffusion 234 -173 234 -173 0 cellNo=380
rlabel pdiffusion 241 -173 241 -173 0 cellNo=149
rlabel pdiffusion 248 -173 248 -173 0 feedthrough
rlabel pdiffusion 255 -173 255 -173 0 feedthrough
rlabel pdiffusion 262 -173 262 -173 0 feedthrough
rlabel pdiffusion 269 -173 269 -173 0 cellNo=308
rlabel pdiffusion 276 -173 276 -173 0 feedthrough
rlabel pdiffusion 283 -173 283 -173 0 feedthrough
rlabel pdiffusion 290 -173 290 -173 0 feedthrough
rlabel pdiffusion 297 -173 297 -173 0 feedthrough
rlabel pdiffusion 304 -173 304 -173 0 feedthrough
rlabel pdiffusion 311 -173 311 -173 0 feedthrough
rlabel pdiffusion 3 -210 3 -210 0 cellNo=279
rlabel pdiffusion 10 -210 10 -210 0 feedthrough
rlabel pdiffusion 17 -210 17 -210 0 feedthrough
rlabel pdiffusion 24 -210 24 -210 0 cellNo=344
rlabel pdiffusion 31 -210 31 -210 0 cellNo=29
rlabel pdiffusion 38 -210 38 -210 0 feedthrough
rlabel pdiffusion 45 -210 45 -210 0 feedthrough
rlabel pdiffusion 52 -210 52 -210 0 cellNo=296
rlabel pdiffusion 59 -210 59 -210 0 feedthrough
rlabel pdiffusion 66 -210 66 -210 0 cellNo=5
rlabel pdiffusion 73 -210 73 -210 0 cellNo=94
rlabel pdiffusion 80 -210 80 -210 0 feedthrough
rlabel pdiffusion 87 -210 87 -210 0 cellNo=249
rlabel pdiffusion 94 -210 94 -210 0 feedthrough
rlabel pdiffusion 101 -210 101 -210 0 feedthrough
rlabel pdiffusion 108 -210 108 -210 0 cellNo=123
rlabel pdiffusion 115 -210 115 -210 0 cellNo=246
rlabel pdiffusion 122 -210 122 -210 0 feedthrough
rlabel pdiffusion 129 -210 129 -210 0 feedthrough
rlabel pdiffusion 136 -210 136 -210 0 feedthrough
rlabel pdiffusion 143 -210 143 -210 0 cellNo=127
rlabel pdiffusion 150 -210 150 -210 0 cellNo=226
rlabel pdiffusion 157 -210 157 -210 0 cellNo=40
rlabel pdiffusion 164 -210 164 -210 0 feedthrough
rlabel pdiffusion 171 -210 171 -210 0 feedthrough
rlabel pdiffusion 178 -210 178 -210 0 feedthrough
rlabel pdiffusion 185 -210 185 -210 0 cellNo=350
rlabel pdiffusion 192 -210 192 -210 0 feedthrough
rlabel pdiffusion 199 -210 199 -210 0 feedthrough
rlabel pdiffusion 206 -210 206 -210 0 cellNo=76
rlabel pdiffusion 213 -210 213 -210 0 cellNo=13
rlabel pdiffusion 220 -210 220 -210 0 cellNo=51
rlabel pdiffusion 227 -210 227 -210 0 feedthrough
rlabel pdiffusion 234 -210 234 -210 0 cellNo=342
rlabel pdiffusion 241 -210 241 -210 0 feedthrough
rlabel pdiffusion 248 -210 248 -210 0 feedthrough
rlabel pdiffusion 255 -210 255 -210 0 feedthrough
rlabel pdiffusion 262 -210 262 -210 0 feedthrough
rlabel pdiffusion 269 -210 269 -210 0 cellNo=87
rlabel pdiffusion 276 -210 276 -210 0 feedthrough
rlabel pdiffusion 283 -210 283 -210 0 cellNo=245
rlabel pdiffusion 290 -210 290 -210 0 cellNo=292
rlabel pdiffusion 297 -210 297 -210 0 feedthrough
rlabel pdiffusion 304 -210 304 -210 0 feedthrough
rlabel pdiffusion 311 -210 311 -210 0 feedthrough
rlabel pdiffusion 318 -210 318 -210 0 feedthrough
rlabel pdiffusion 325 -210 325 -210 0 feedthrough
rlabel pdiffusion 332 -210 332 -210 0 feedthrough
rlabel pdiffusion 339 -210 339 -210 0 feedthrough
rlabel pdiffusion 346 -210 346 -210 0 feedthrough
rlabel pdiffusion 353 -210 353 -210 0 feedthrough
rlabel pdiffusion 360 -210 360 -210 0 feedthrough
rlabel pdiffusion 367 -210 367 -210 0 feedthrough
rlabel pdiffusion 374 -210 374 -210 0 feedthrough
rlabel pdiffusion 381 -210 381 -210 0 feedthrough
rlabel pdiffusion 388 -210 388 -210 0 cellNo=400
rlabel pdiffusion 395 -210 395 -210 0 feedthrough
rlabel pdiffusion 10 -255 10 -255 0 feedthrough
rlabel pdiffusion 17 -255 17 -255 0 feedthrough
rlabel pdiffusion 24 -255 24 -255 0 cellNo=158
rlabel pdiffusion 31 -255 31 -255 0 feedthrough
rlabel pdiffusion 38 -255 38 -255 0 feedthrough
rlabel pdiffusion 45 -255 45 -255 0 feedthrough
rlabel pdiffusion 52 -255 52 -255 0 feedthrough
rlabel pdiffusion 59 -255 59 -255 0 feedthrough
rlabel pdiffusion 66 -255 66 -255 0 cellNo=72
rlabel pdiffusion 73 -255 73 -255 0 cellNo=90
rlabel pdiffusion 80 -255 80 -255 0 cellNo=112
rlabel pdiffusion 87 -255 87 -255 0 feedthrough
rlabel pdiffusion 94 -255 94 -255 0 feedthrough
rlabel pdiffusion 101 -255 101 -255 0 cellNo=146
rlabel pdiffusion 108 -255 108 -255 0 cellNo=132
rlabel pdiffusion 115 -255 115 -255 0 feedthrough
rlabel pdiffusion 122 -255 122 -255 0 cellNo=89
rlabel pdiffusion 129 -255 129 -255 0 feedthrough
rlabel pdiffusion 136 -255 136 -255 0 cellNo=113
rlabel pdiffusion 143 -255 143 -255 0 feedthrough
rlabel pdiffusion 150 -255 150 -255 0 cellNo=288
rlabel pdiffusion 157 -255 157 -255 0 cellNo=34
rlabel pdiffusion 164 -255 164 -255 0 feedthrough
rlabel pdiffusion 171 -255 171 -255 0 feedthrough
rlabel pdiffusion 178 -255 178 -255 0 feedthrough
rlabel pdiffusion 185 -255 185 -255 0 feedthrough
rlabel pdiffusion 192 -255 192 -255 0 feedthrough
rlabel pdiffusion 199 -255 199 -255 0 cellNo=152
rlabel pdiffusion 206 -255 206 -255 0 cellNo=376
rlabel pdiffusion 213 -255 213 -255 0 cellNo=199
rlabel pdiffusion 220 -255 220 -255 0 feedthrough
rlabel pdiffusion 227 -255 227 -255 0 cellNo=155
rlabel pdiffusion 234 -255 234 -255 0 feedthrough
rlabel pdiffusion 241 -255 241 -255 0 feedthrough
rlabel pdiffusion 248 -255 248 -255 0 feedthrough
rlabel pdiffusion 255 -255 255 -255 0 feedthrough
rlabel pdiffusion 262 -255 262 -255 0 cellNo=192
rlabel pdiffusion 269 -255 269 -255 0 feedthrough
rlabel pdiffusion 276 -255 276 -255 0 cellNo=183
rlabel pdiffusion 283 -255 283 -255 0 feedthrough
rlabel pdiffusion 290 -255 290 -255 0 cellNo=135
rlabel pdiffusion 297 -255 297 -255 0 feedthrough
rlabel pdiffusion 304 -255 304 -255 0 feedthrough
rlabel pdiffusion 311 -255 311 -255 0 feedthrough
rlabel pdiffusion 318 -255 318 -255 0 feedthrough
rlabel pdiffusion 325 -255 325 -255 0 feedthrough
rlabel pdiffusion 332 -255 332 -255 0 feedthrough
rlabel pdiffusion 339 -255 339 -255 0 feedthrough
rlabel pdiffusion 346 -255 346 -255 0 feedthrough
rlabel pdiffusion 353 -255 353 -255 0 feedthrough
rlabel pdiffusion 360 -255 360 -255 0 feedthrough
rlabel pdiffusion 367 -255 367 -255 0 cellNo=2
rlabel pdiffusion 374 -255 374 -255 0 cellNo=255
rlabel pdiffusion 381 -255 381 -255 0 feedthrough
rlabel pdiffusion 3 -302 3 -302 0 feedthrough
rlabel pdiffusion 10 -302 10 -302 0 feedthrough
rlabel pdiffusion 17 -302 17 -302 0 feedthrough
rlabel pdiffusion 24 -302 24 -302 0 feedthrough
rlabel pdiffusion 31 -302 31 -302 0 feedthrough
rlabel pdiffusion 38 -302 38 -302 0 feedthrough
rlabel pdiffusion 45 -302 45 -302 0 feedthrough
rlabel pdiffusion 52 -302 52 -302 0 cellNo=261
rlabel pdiffusion 59 -302 59 -302 0 cellNo=12
rlabel pdiffusion 66 -302 66 -302 0 feedthrough
rlabel pdiffusion 73 -302 73 -302 0 feedthrough
rlabel pdiffusion 80 -302 80 -302 0 cellNo=167
rlabel pdiffusion 87 -302 87 -302 0 feedthrough
rlabel pdiffusion 94 -302 94 -302 0 feedthrough
rlabel pdiffusion 101 -302 101 -302 0 feedthrough
rlabel pdiffusion 108 -302 108 -302 0 feedthrough
rlabel pdiffusion 115 -302 115 -302 0 feedthrough
rlabel pdiffusion 122 -302 122 -302 0 cellNo=233
rlabel pdiffusion 129 -302 129 -302 0 feedthrough
rlabel pdiffusion 136 -302 136 -302 0 cellNo=157
rlabel pdiffusion 143 -302 143 -302 0 feedthrough
rlabel pdiffusion 150 -302 150 -302 0 feedthrough
rlabel pdiffusion 157 -302 157 -302 0 cellNo=171
rlabel pdiffusion 164 -302 164 -302 0 cellNo=252
rlabel pdiffusion 171 -302 171 -302 0 feedthrough
rlabel pdiffusion 178 -302 178 -302 0 feedthrough
rlabel pdiffusion 185 -302 185 -302 0 cellNo=168
rlabel pdiffusion 192 -302 192 -302 0 feedthrough
rlabel pdiffusion 199 -302 199 -302 0 cellNo=265
rlabel pdiffusion 206 -302 206 -302 0 cellNo=154
rlabel pdiffusion 213 -302 213 -302 0 cellNo=10
rlabel pdiffusion 220 -302 220 -302 0 feedthrough
rlabel pdiffusion 227 -302 227 -302 0 feedthrough
rlabel pdiffusion 234 -302 234 -302 0 cellNo=96
rlabel pdiffusion 241 -302 241 -302 0 cellNo=173
rlabel pdiffusion 248 -302 248 -302 0 cellNo=377
rlabel pdiffusion 255 -302 255 -302 0 cellNo=156
rlabel pdiffusion 262 -302 262 -302 0 feedthrough
rlabel pdiffusion 269 -302 269 -302 0 feedthrough
rlabel pdiffusion 276 -302 276 -302 0 feedthrough
rlabel pdiffusion 283 -302 283 -302 0 feedthrough
rlabel pdiffusion 290 -302 290 -302 0 feedthrough
rlabel pdiffusion 297 -302 297 -302 0 cellNo=389
rlabel pdiffusion 304 -302 304 -302 0 feedthrough
rlabel pdiffusion 311 -302 311 -302 0 feedthrough
rlabel pdiffusion 318 -302 318 -302 0 feedthrough
rlabel pdiffusion 325 -302 325 -302 0 feedthrough
rlabel pdiffusion 332 -302 332 -302 0 feedthrough
rlabel pdiffusion 339 -302 339 -302 0 feedthrough
rlabel pdiffusion 346 -302 346 -302 0 feedthrough
rlabel pdiffusion 353 -302 353 -302 0 feedthrough
rlabel pdiffusion 360 -302 360 -302 0 feedthrough
rlabel pdiffusion 367 -302 367 -302 0 cellNo=45
rlabel pdiffusion 374 -302 374 -302 0 cellNo=185
rlabel pdiffusion 381 -302 381 -302 0 feedthrough
rlabel pdiffusion 3 -343 3 -343 0 feedthrough
rlabel pdiffusion 10 -343 10 -343 0 feedthrough
rlabel pdiffusion 17 -343 17 -343 0 feedthrough
rlabel pdiffusion 24 -343 24 -343 0 feedthrough
rlabel pdiffusion 31 -343 31 -343 0 feedthrough
rlabel pdiffusion 38 -343 38 -343 0 feedthrough
rlabel pdiffusion 45 -343 45 -343 0 cellNo=297
rlabel pdiffusion 52 -343 52 -343 0 feedthrough
rlabel pdiffusion 59 -343 59 -343 0 cellNo=69
rlabel pdiffusion 66 -343 66 -343 0 cellNo=124
rlabel pdiffusion 73 -343 73 -343 0 feedthrough
rlabel pdiffusion 80 -343 80 -343 0 feedthrough
rlabel pdiffusion 87 -343 87 -343 0 cellNo=210
rlabel pdiffusion 94 -343 94 -343 0 feedthrough
rlabel pdiffusion 101 -343 101 -343 0 cellNo=98
rlabel pdiffusion 108 -343 108 -343 0 cellNo=315
rlabel pdiffusion 115 -343 115 -343 0 cellNo=277
rlabel pdiffusion 122 -343 122 -343 0 cellNo=20
rlabel pdiffusion 129 -343 129 -343 0 feedthrough
rlabel pdiffusion 136 -343 136 -343 0 feedthrough
rlabel pdiffusion 143 -343 143 -343 0 cellNo=273
rlabel pdiffusion 150 -343 150 -343 0 cellNo=58
rlabel pdiffusion 157 -343 157 -343 0 cellNo=100
rlabel pdiffusion 164 -343 164 -343 0 feedthrough
rlabel pdiffusion 171 -343 171 -343 0 cellNo=268
rlabel pdiffusion 178 -343 178 -343 0 feedthrough
rlabel pdiffusion 185 -343 185 -343 0 feedthrough
rlabel pdiffusion 192 -343 192 -343 0 cellNo=30
rlabel pdiffusion 199 -343 199 -343 0 feedthrough
rlabel pdiffusion 206 -343 206 -343 0 cellNo=145
rlabel pdiffusion 213 -343 213 -343 0 cellNo=395
rlabel pdiffusion 220 -343 220 -343 0 feedthrough
rlabel pdiffusion 227 -343 227 -343 0 feedthrough
rlabel pdiffusion 234 -343 234 -343 0 cellNo=144
rlabel pdiffusion 241 -343 241 -343 0 cellNo=218
rlabel pdiffusion 248 -343 248 -343 0 feedthrough
rlabel pdiffusion 255 -343 255 -343 0 feedthrough
rlabel pdiffusion 262 -343 262 -343 0 feedthrough
rlabel pdiffusion 269 -343 269 -343 0 feedthrough
rlabel pdiffusion 276 -343 276 -343 0 feedthrough
rlabel pdiffusion 283 -343 283 -343 0 feedthrough
rlabel pdiffusion 290 -343 290 -343 0 feedthrough
rlabel pdiffusion 297 -343 297 -343 0 feedthrough
rlabel pdiffusion 304 -343 304 -343 0 feedthrough
rlabel pdiffusion 311 -343 311 -343 0 feedthrough
rlabel pdiffusion 318 -343 318 -343 0 feedthrough
rlabel pdiffusion 325 -343 325 -343 0 feedthrough
rlabel pdiffusion 332 -343 332 -343 0 feedthrough
rlabel pdiffusion 339 -343 339 -343 0 cellNo=280
rlabel pdiffusion 346 -343 346 -343 0 feedthrough
rlabel pdiffusion 353 -343 353 -343 0 feedthrough
rlabel pdiffusion 360 -343 360 -343 0 feedthrough
rlabel pdiffusion 374 -343 374 -343 0 cellNo=204
rlabel pdiffusion 388 -343 388 -343 0 feedthrough
rlabel pdiffusion 10 -388 10 -388 0 feedthrough
rlabel pdiffusion 17 -388 17 -388 0 feedthrough
rlabel pdiffusion 24 -388 24 -388 0 feedthrough
rlabel pdiffusion 31 -388 31 -388 0 feedthrough
rlabel pdiffusion 38 -388 38 -388 0 feedthrough
rlabel pdiffusion 45 -388 45 -388 0 feedthrough
rlabel pdiffusion 52 -388 52 -388 0 feedthrough
rlabel pdiffusion 59 -388 59 -388 0 feedthrough
rlabel pdiffusion 66 -388 66 -388 0 cellNo=4
rlabel pdiffusion 73 -388 73 -388 0 feedthrough
rlabel pdiffusion 80 -388 80 -388 0 cellNo=357
rlabel pdiffusion 87 -388 87 -388 0 cellNo=46
rlabel pdiffusion 94 -388 94 -388 0 cellNo=250
rlabel pdiffusion 101 -388 101 -388 0 feedthrough
rlabel pdiffusion 108 -388 108 -388 0 feedthrough
rlabel pdiffusion 115 -388 115 -388 0 cellNo=99
rlabel pdiffusion 122 -388 122 -388 0 feedthrough
rlabel pdiffusion 129 -388 129 -388 0 cellNo=111
rlabel pdiffusion 136 -388 136 -388 0 feedthrough
rlabel pdiffusion 143 -388 143 -388 0 cellNo=290
rlabel pdiffusion 150 -388 150 -388 0 cellNo=137
rlabel pdiffusion 157 -388 157 -388 0 cellNo=181
rlabel pdiffusion 164 -388 164 -388 0 feedthrough
rlabel pdiffusion 171 -388 171 -388 0 cellNo=86
rlabel pdiffusion 178 -388 178 -388 0 feedthrough
rlabel pdiffusion 185 -388 185 -388 0 cellNo=299
rlabel pdiffusion 192 -388 192 -388 0 cellNo=205
rlabel pdiffusion 199 -388 199 -388 0 feedthrough
rlabel pdiffusion 206 -388 206 -388 0 feedthrough
rlabel pdiffusion 213 -388 213 -388 0 cellNo=184
rlabel pdiffusion 220 -388 220 -388 0 cellNo=345
rlabel pdiffusion 227 -388 227 -388 0 feedthrough
rlabel pdiffusion 234 -388 234 -388 0 feedthrough
rlabel pdiffusion 241 -388 241 -388 0 cellNo=193
rlabel pdiffusion 248 -388 248 -388 0 feedthrough
rlabel pdiffusion 255 -388 255 -388 0 cellNo=197
rlabel pdiffusion 262 -388 262 -388 0 feedthrough
rlabel pdiffusion 269 -388 269 -388 0 cellNo=260
rlabel pdiffusion 276 -388 276 -388 0 feedthrough
rlabel pdiffusion 283 -388 283 -388 0 cellNo=17
rlabel pdiffusion 290 -388 290 -388 0 feedthrough
rlabel pdiffusion 297 -388 297 -388 0 feedthrough
rlabel pdiffusion 304 -388 304 -388 0 feedthrough
rlabel pdiffusion 311 -388 311 -388 0 feedthrough
rlabel pdiffusion 318 -388 318 -388 0 feedthrough
rlabel pdiffusion 325 -388 325 -388 0 feedthrough
rlabel pdiffusion 332 -388 332 -388 0 feedthrough
rlabel pdiffusion 339 -388 339 -388 0 feedthrough
rlabel pdiffusion 346 -388 346 -388 0 feedthrough
rlabel pdiffusion 353 -388 353 -388 0 feedthrough
rlabel pdiffusion 360 -388 360 -388 0 feedthrough
rlabel pdiffusion 367 -388 367 -388 0 feedthrough
rlabel pdiffusion 374 -388 374 -388 0 feedthrough
rlabel pdiffusion 381 -388 381 -388 0 feedthrough
rlabel pdiffusion 388 -388 388 -388 0 feedthrough
rlabel pdiffusion 395 -388 395 -388 0 cellNo=240
rlabel pdiffusion 402 -388 402 -388 0 feedthrough
rlabel pdiffusion 409 -388 409 -388 0 cellNo=347
rlabel pdiffusion 24 -427 24 -427 0 feedthrough
rlabel pdiffusion 31 -427 31 -427 0 feedthrough
rlabel pdiffusion 38 -427 38 -427 0 cellNo=330
rlabel pdiffusion 45 -427 45 -427 0 cellNo=303
rlabel pdiffusion 52 -427 52 -427 0 cellNo=93
rlabel pdiffusion 59 -427 59 -427 0 feedthrough
rlabel pdiffusion 66 -427 66 -427 0 cellNo=318
rlabel pdiffusion 73 -427 73 -427 0 feedthrough
rlabel pdiffusion 80 -427 80 -427 0 feedthrough
rlabel pdiffusion 87 -427 87 -427 0 feedthrough
rlabel pdiffusion 94 -427 94 -427 0 cellNo=163
rlabel pdiffusion 101 -427 101 -427 0 cellNo=339
rlabel pdiffusion 108 -427 108 -427 0 cellNo=298
rlabel pdiffusion 115 -427 115 -427 0 cellNo=301
rlabel pdiffusion 122 -427 122 -427 0 feedthrough
rlabel pdiffusion 129 -427 129 -427 0 feedthrough
rlabel pdiffusion 136 -427 136 -427 0 cellNo=134
rlabel pdiffusion 143 -427 143 -427 0 feedthrough
rlabel pdiffusion 150 -427 150 -427 0 feedthrough
rlabel pdiffusion 157 -427 157 -427 0 cellNo=106
rlabel pdiffusion 164 -427 164 -427 0 cellNo=275
rlabel pdiffusion 171 -427 171 -427 0 feedthrough
rlabel pdiffusion 178 -427 178 -427 0 feedthrough
rlabel pdiffusion 185 -427 185 -427 0 feedthrough
rlabel pdiffusion 192 -427 192 -427 0 cellNo=208
rlabel pdiffusion 199 -427 199 -427 0 cellNo=64
rlabel pdiffusion 206 -427 206 -427 0 cellNo=305
rlabel pdiffusion 213 -427 213 -427 0 cellNo=79
rlabel pdiffusion 220 -427 220 -427 0 feedthrough
rlabel pdiffusion 227 -427 227 -427 0 feedthrough
rlabel pdiffusion 234 -427 234 -427 0 feedthrough
rlabel pdiffusion 241 -427 241 -427 0 cellNo=276
rlabel pdiffusion 248 -427 248 -427 0 cellNo=306
rlabel pdiffusion 255 -427 255 -427 0 cellNo=28
rlabel pdiffusion 262 -427 262 -427 0 feedthrough
rlabel pdiffusion 269 -427 269 -427 0 feedthrough
rlabel pdiffusion 276 -427 276 -427 0 feedthrough
rlabel pdiffusion 283 -427 283 -427 0 cellNo=224
rlabel pdiffusion 290 -427 290 -427 0 feedthrough
rlabel pdiffusion 297 -427 297 -427 0 feedthrough
rlabel pdiffusion 304 -427 304 -427 0 feedthrough
rlabel pdiffusion 311 -427 311 -427 0 feedthrough
rlabel pdiffusion 318 -427 318 -427 0 feedthrough
rlabel pdiffusion 325 -427 325 -427 0 feedthrough
rlabel pdiffusion 332 -427 332 -427 0 feedthrough
rlabel pdiffusion 339 -427 339 -427 0 feedthrough
rlabel pdiffusion 346 -427 346 -427 0 feedthrough
rlabel pdiffusion 353 -427 353 -427 0 cellNo=117
rlabel pdiffusion 360 -427 360 -427 0 cellNo=354
rlabel pdiffusion 367 -427 367 -427 0 feedthrough
rlabel pdiffusion 374 -427 374 -427 0 feedthrough
rlabel pdiffusion 381 -427 381 -427 0 feedthrough
rlabel pdiffusion 24 -460 24 -460 0 cellNo=41
rlabel pdiffusion 31 -460 31 -460 0 cellNo=83
rlabel pdiffusion 38 -460 38 -460 0 feedthrough
rlabel pdiffusion 45 -460 45 -460 0 feedthrough
rlabel pdiffusion 52 -460 52 -460 0 feedthrough
rlabel pdiffusion 59 -460 59 -460 0 feedthrough
rlabel pdiffusion 66 -460 66 -460 0 cellNo=271
rlabel pdiffusion 73 -460 73 -460 0 cellNo=254
rlabel pdiffusion 80 -460 80 -460 0 feedthrough
rlabel pdiffusion 87 -460 87 -460 0 feedthrough
rlabel pdiffusion 94 -460 94 -460 0 feedthrough
rlabel pdiffusion 101 -460 101 -460 0 feedthrough
rlabel pdiffusion 108 -460 108 -460 0 feedthrough
rlabel pdiffusion 115 -460 115 -460 0 cellNo=1
rlabel pdiffusion 122 -460 122 -460 0 cellNo=300
rlabel pdiffusion 129 -460 129 -460 0 cellNo=329
rlabel pdiffusion 136 -460 136 -460 0 cellNo=216
rlabel pdiffusion 143 -460 143 -460 0 cellNo=39
rlabel pdiffusion 150 -460 150 -460 0 feedthrough
rlabel pdiffusion 157 -460 157 -460 0 cellNo=105
rlabel pdiffusion 164 -460 164 -460 0 feedthrough
rlabel pdiffusion 171 -460 171 -460 0 feedthrough
rlabel pdiffusion 178 -460 178 -460 0 feedthrough
rlabel pdiffusion 185 -460 185 -460 0 cellNo=85
rlabel pdiffusion 192 -460 192 -460 0 cellNo=162
rlabel pdiffusion 199 -460 199 -460 0 feedthrough
rlabel pdiffusion 206 -460 206 -460 0 feedthrough
rlabel pdiffusion 213 -460 213 -460 0 cellNo=66
rlabel pdiffusion 220 -460 220 -460 0 feedthrough
rlabel pdiffusion 227 -460 227 -460 0 cellNo=239
rlabel pdiffusion 234 -460 234 -460 0 feedthrough
rlabel pdiffusion 241 -460 241 -460 0 feedthrough
rlabel pdiffusion 248 -460 248 -460 0 cellNo=341
rlabel pdiffusion 255 -460 255 -460 0 feedthrough
rlabel pdiffusion 262 -460 262 -460 0 feedthrough
rlabel pdiffusion 269 -460 269 -460 0 feedthrough
rlabel pdiffusion 276 -460 276 -460 0 feedthrough
rlabel pdiffusion 283 -460 283 -460 0 feedthrough
rlabel pdiffusion 290 -460 290 -460 0 feedthrough
rlabel pdiffusion 297 -460 297 -460 0 feedthrough
rlabel pdiffusion 304 -460 304 -460 0 cellNo=21
rlabel pdiffusion 311 -460 311 -460 0 cellNo=358
rlabel pdiffusion 318 -460 318 -460 0 cellNo=223
rlabel pdiffusion 332 -460 332 -460 0 feedthrough
rlabel pdiffusion 353 -460 353 -460 0 feedthrough
rlabel pdiffusion 360 -460 360 -460 0 feedthrough
rlabel pdiffusion 367 -460 367 -460 0 feedthrough
rlabel pdiffusion 374 -460 374 -460 0 cellNo=78
rlabel pdiffusion 38 -497 38 -497 0 feedthrough
rlabel pdiffusion 45 -497 45 -497 0 feedthrough
rlabel pdiffusion 52 -497 52 -497 0 feedthrough
rlabel pdiffusion 59 -497 59 -497 0 feedthrough
rlabel pdiffusion 66 -497 66 -497 0 cellNo=282
rlabel pdiffusion 73 -497 73 -497 0 feedthrough
rlabel pdiffusion 80 -497 80 -497 0 feedthrough
rlabel pdiffusion 87 -497 87 -497 0 feedthrough
rlabel pdiffusion 94 -497 94 -497 0 cellNo=394
rlabel pdiffusion 101 -497 101 -497 0 feedthrough
rlabel pdiffusion 108 -497 108 -497 0 cellNo=384
rlabel pdiffusion 115 -497 115 -497 0 cellNo=313
rlabel pdiffusion 122 -497 122 -497 0 feedthrough
rlabel pdiffusion 129 -497 129 -497 0 cellNo=325
rlabel pdiffusion 136 -497 136 -497 0 feedthrough
rlabel pdiffusion 143 -497 143 -497 0 feedthrough
rlabel pdiffusion 150 -497 150 -497 0 feedthrough
rlabel pdiffusion 157 -497 157 -497 0 feedthrough
rlabel pdiffusion 164 -497 164 -497 0 feedthrough
rlabel pdiffusion 171 -497 171 -497 0 cellNo=215
rlabel pdiffusion 178 -497 178 -497 0 feedthrough
rlabel pdiffusion 185 -497 185 -497 0 feedthrough
rlabel pdiffusion 192 -497 192 -497 0 cellNo=259
rlabel pdiffusion 199 -497 199 -497 0 cellNo=133
rlabel pdiffusion 206 -497 206 -497 0 cellNo=286
rlabel pdiffusion 213 -497 213 -497 0 cellNo=103
rlabel pdiffusion 220 -497 220 -497 0 cellNo=230
rlabel pdiffusion 227 -497 227 -497 0 feedthrough
rlabel pdiffusion 234 -497 234 -497 0 feedthrough
rlabel pdiffusion 241 -497 241 -497 0 cellNo=236
rlabel pdiffusion 248 -497 248 -497 0 feedthrough
rlabel pdiffusion 255 -497 255 -497 0 feedthrough
rlabel pdiffusion 262 -497 262 -497 0 feedthrough
rlabel pdiffusion 269 -497 269 -497 0 feedthrough
rlabel pdiffusion 276 -497 276 -497 0 feedthrough
rlabel pdiffusion 283 -497 283 -497 0 cellNo=15
rlabel pdiffusion 290 -497 290 -497 0 feedthrough
rlabel pdiffusion 297 -497 297 -497 0 cellNo=206
rlabel pdiffusion 304 -497 304 -497 0 feedthrough
rlabel pdiffusion 311 -497 311 -497 0 cellNo=363
rlabel pdiffusion 318 -497 318 -497 0 cellNo=382
rlabel pdiffusion 325 -497 325 -497 0 feedthrough
rlabel pdiffusion 332 -497 332 -497 0 feedthrough
rlabel pdiffusion 339 -497 339 -497 0 cellNo=327
rlabel pdiffusion 346 -497 346 -497 0 cellNo=182
rlabel pdiffusion 353 -497 353 -497 0 feedthrough
rlabel pdiffusion 360 -497 360 -497 0 cellNo=48
rlabel pdiffusion 17 -536 17 -536 0 feedthrough
rlabel pdiffusion 24 -536 24 -536 0 cellNo=101
rlabel pdiffusion 31 -536 31 -536 0 feedthrough
rlabel pdiffusion 38 -536 38 -536 0 feedthrough
rlabel pdiffusion 45 -536 45 -536 0 feedthrough
rlabel pdiffusion 52 -536 52 -536 0 feedthrough
rlabel pdiffusion 59 -536 59 -536 0 feedthrough
rlabel pdiffusion 66 -536 66 -536 0 feedthrough
rlabel pdiffusion 73 -536 73 -536 0 cellNo=52
rlabel pdiffusion 80 -536 80 -536 0 feedthrough
rlabel pdiffusion 87 -536 87 -536 0 feedthrough
rlabel pdiffusion 94 -536 94 -536 0 cellNo=278
rlabel pdiffusion 101 -536 101 -536 0 cellNo=104
rlabel pdiffusion 108 -536 108 -536 0 cellNo=61
rlabel pdiffusion 115 -536 115 -536 0 feedthrough
rlabel pdiffusion 122 -536 122 -536 0 cellNo=73
rlabel pdiffusion 129 -536 129 -536 0 cellNo=179
rlabel pdiffusion 136 -536 136 -536 0 feedthrough
rlabel pdiffusion 143 -536 143 -536 0 cellNo=319
rlabel pdiffusion 150 -536 150 -536 0 cellNo=337
rlabel pdiffusion 157 -536 157 -536 0 cellNo=71
rlabel pdiffusion 164 -536 164 -536 0 cellNo=309
rlabel pdiffusion 171 -536 171 -536 0 feedthrough
rlabel pdiffusion 178 -536 178 -536 0 feedthrough
rlabel pdiffusion 185 -536 185 -536 0 cellNo=109
rlabel pdiffusion 192 -536 192 -536 0 cellNo=242
rlabel pdiffusion 199 -536 199 -536 0 cellNo=37
rlabel pdiffusion 206 -536 206 -536 0 cellNo=370
rlabel pdiffusion 213 -536 213 -536 0 feedthrough
rlabel pdiffusion 220 -536 220 -536 0 cellNo=338
rlabel pdiffusion 227 -536 227 -536 0 cellNo=11
rlabel pdiffusion 234 -536 234 -536 0 feedthrough
rlabel pdiffusion 241 -536 241 -536 0 feedthrough
rlabel pdiffusion 248 -536 248 -536 0 feedthrough
rlabel pdiffusion 255 -536 255 -536 0 feedthrough
rlabel pdiffusion 262 -536 262 -536 0 feedthrough
rlabel pdiffusion 269 -536 269 -536 0 feedthrough
rlabel pdiffusion 276 -536 276 -536 0 cellNo=175
rlabel pdiffusion 283 -536 283 -536 0 feedthrough
rlabel pdiffusion 290 -536 290 -536 0 feedthrough
rlabel pdiffusion 297 -536 297 -536 0 feedthrough
rlabel pdiffusion 304 -536 304 -536 0 feedthrough
rlabel pdiffusion 311 -536 311 -536 0 feedthrough
rlabel pdiffusion 318 -536 318 -536 0 feedthrough
rlabel pdiffusion 325 -536 325 -536 0 feedthrough
rlabel pdiffusion 332 -536 332 -536 0 feedthrough
rlabel pdiffusion 339 -536 339 -536 0 cellNo=49
rlabel pdiffusion 346 -536 346 -536 0 cellNo=50
rlabel pdiffusion 353 -536 353 -536 0 feedthrough
rlabel pdiffusion 360 -536 360 -536 0 feedthrough
rlabel pdiffusion 367 -536 367 -536 0 feedthrough
rlabel pdiffusion 374 -536 374 -536 0 feedthrough
rlabel pdiffusion 10 -575 10 -575 0 feedthrough
rlabel pdiffusion 17 -575 17 -575 0 feedthrough
rlabel pdiffusion 24 -575 24 -575 0 cellNo=70
rlabel pdiffusion 31 -575 31 -575 0 cellNo=269
rlabel pdiffusion 38 -575 38 -575 0 cellNo=388
rlabel pdiffusion 45 -575 45 -575 0 cellNo=211
rlabel pdiffusion 52 -575 52 -575 0 cellNo=307
rlabel pdiffusion 59 -575 59 -575 0 feedthrough
rlabel pdiffusion 66 -575 66 -575 0 feedthrough
rlabel pdiffusion 73 -575 73 -575 0 feedthrough
rlabel pdiffusion 80 -575 80 -575 0 cellNo=274
rlabel pdiffusion 87 -575 87 -575 0 feedthrough
rlabel pdiffusion 94 -575 94 -575 0 feedthrough
rlabel pdiffusion 101 -575 101 -575 0 feedthrough
rlabel pdiffusion 108 -575 108 -575 0 cellNo=243
rlabel pdiffusion 115 -575 115 -575 0 feedthrough
rlabel pdiffusion 122 -575 122 -575 0 cellNo=264
rlabel pdiffusion 129 -575 129 -575 0 cellNo=323
rlabel pdiffusion 136 -575 136 -575 0 feedthrough
rlabel pdiffusion 143 -575 143 -575 0 cellNo=353
rlabel pdiffusion 150 -575 150 -575 0 cellNo=27
rlabel pdiffusion 157 -575 157 -575 0 cellNo=383
rlabel pdiffusion 164 -575 164 -575 0 feedthrough
rlabel pdiffusion 171 -575 171 -575 0 cellNo=195
rlabel pdiffusion 178 -575 178 -575 0 feedthrough
rlabel pdiffusion 185 -575 185 -575 0 cellNo=258
rlabel pdiffusion 192 -575 192 -575 0 feedthrough
rlabel pdiffusion 199 -575 199 -575 0 feedthrough
rlabel pdiffusion 206 -575 206 -575 0 feedthrough
rlabel pdiffusion 213 -575 213 -575 0 feedthrough
rlabel pdiffusion 220 -575 220 -575 0 feedthrough
rlabel pdiffusion 227 -575 227 -575 0 feedthrough
rlabel pdiffusion 234 -575 234 -575 0 cellNo=81
rlabel pdiffusion 241 -575 241 -575 0 feedthrough
rlabel pdiffusion 248 -575 248 -575 0 feedthrough
rlabel pdiffusion 255 -575 255 -575 0 cellNo=368
rlabel pdiffusion 262 -575 262 -575 0 feedthrough
rlabel pdiffusion 269 -575 269 -575 0 feedthrough
rlabel pdiffusion 276 -575 276 -575 0 cellNo=391
rlabel pdiffusion 283 -575 283 -575 0 feedthrough
rlabel pdiffusion 290 -575 290 -575 0 cellNo=229
rlabel pdiffusion 297 -575 297 -575 0 feedthrough
rlabel pdiffusion 304 -575 304 -575 0 feedthrough
rlabel pdiffusion 311 -575 311 -575 0 cellNo=130
rlabel pdiffusion 325 -575 325 -575 0 feedthrough
rlabel pdiffusion 353 -575 353 -575 0 cellNo=348
rlabel pdiffusion 360 -575 360 -575 0 feedthrough
rlabel pdiffusion 24 -606 24 -606 0 cellNo=293
rlabel pdiffusion 31 -606 31 -606 0 feedthrough
rlabel pdiffusion 38 -606 38 -606 0 cellNo=24
rlabel pdiffusion 45 -606 45 -606 0 feedthrough
rlabel pdiffusion 52 -606 52 -606 0 feedthrough
rlabel pdiffusion 59 -606 59 -606 0 feedthrough
rlabel pdiffusion 66 -606 66 -606 0 feedthrough
rlabel pdiffusion 73 -606 73 -606 0 cellNo=371
rlabel pdiffusion 80 -606 80 -606 0 cellNo=396
rlabel pdiffusion 87 -606 87 -606 0 feedthrough
rlabel pdiffusion 94 -606 94 -606 0 cellNo=331
rlabel pdiffusion 101 -606 101 -606 0 cellNo=110
rlabel pdiffusion 108 -606 108 -606 0 feedthrough
rlabel pdiffusion 115 -606 115 -606 0 cellNo=386
rlabel pdiffusion 122 -606 122 -606 0 feedthrough
rlabel pdiffusion 129 -606 129 -606 0 cellNo=234
rlabel pdiffusion 136 -606 136 -606 0 cellNo=214
rlabel pdiffusion 143 -606 143 -606 0 feedthrough
rlabel pdiffusion 150 -606 150 -606 0 cellNo=367
rlabel pdiffusion 157 -606 157 -606 0 cellNo=115
rlabel pdiffusion 164 -606 164 -606 0 feedthrough
rlabel pdiffusion 171 -606 171 -606 0 feedthrough
rlabel pdiffusion 178 -606 178 -606 0 cellNo=150
rlabel pdiffusion 185 -606 185 -606 0 cellNo=322
rlabel pdiffusion 192 -606 192 -606 0 feedthrough
rlabel pdiffusion 199 -606 199 -606 0 feedthrough
rlabel pdiffusion 206 -606 206 -606 0 feedthrough
rlabel pdiffusion 213 -606 213 -606 0 feedthrough
rlabel pdiffusion 220 -606 220 -606 0 feedthrough
rlabel pdiffusion 227 -606 227 -606 0 cellNo=326
rlabel pdiffusion 234 -606 234 -606 0 feedthrough
rlabel pdiffusion 241 -606 241 -606 0 cellNo=335
rlabel pdiffusion 248 -606 248 -606 0 feedthrough
rlabel pdiffusion 255 -606 255 -606 0 feedthrough
rlabel pdiffusion 262 -606 262 -606 0 feedthrough
rlabel pdiffusion 269 -606 269 -606 0 feedthrough
rlabel pdiffusion 276 -606 276 -606 0 cellNo=122
rlabel pdiffusion 283 -606 283 -606 0 feedthrough
rlabel pdiffusion 290 -606 290 -606 0 feedthrough
rlabel pdiffusion 304 -606 304 -606 0 cellNo=248
rlabel pdiffusion 325 -606 325 -606 0 feedthrough
rlabel pdiffusion 24 -631 24 -631 0 cellNo=334
rlabel pdiffusion 52 -631 52 -631 0 feedthrough
rlabel pdiffusion 66 -631 66 -631 0 feedthrough
rlabel pdiffusion 73 -631 73 -631 0 cellNo=311
rlabel pdiffusion 80 -631 80 -631 0 cellNo=378
rlabel pdiffusion 87 -631 87 -631 0 cellNo=139
rlabel pdiffusion 94 -631 94 -631 0 feedthrough
rlabel pdiffusion 101 -631 101 -631 0 cellNo=270
rlabel pdiffusion 108 -631 108 -631 0 cellNo=346
rlabel pdiffusion 115 -631 115 -631 0 cellNo=187
rlabel pdiffusion 122 -631 122 -631 0 feedthrough
rlabel pdiffusion 129 -631 129 -631 0 feedthrough
rlabel pdiffusion 136 -631 136 -631 0 feedthrough
rlabel pdiffusion 143 -631 143 -631 0 cellNo=160
rlabel pdiffusion 150 -631 150 -631 0 cellNo=159
rlabel pdiffusion 157 -631 157 -631 0 feedthrough
rlabel pdiffusion 164 -631 164 -631 0 feedthrough
rlabel pdiffusion 171 -631 171 -631 0 cellNo=381
rlabel pdiffusion 178 -631 178 -631 0 cellNo=272
rlabel pdiffusion 185 -631 185 -631 0 cellNo=142
rlabel pdiffusion 192 -631 192 -631 0 feedthrough
rlabel pdiffusion 199 -631 199 -631 0 feedthrough
rlabel pdiffusion 206 -631 206 -631 0 feedthrough
rlabel pdiffusion 213 -631 213 -631 0 feedthrough
rlabel pdiffusion 220 -631 220 -631 0 feedthrough
rlabel pdiffusion 227 -631 227 -631 0 feedthrough
rlabel pdiffusion 234 -631 234 -631 0 cellNo=314
rlabel pdiffusion 241 -631 241 -631 0 feedthrough
rlabel pdiffusion 248 -631 248 -631 0 cellNo=374
rlabel pdiffusion 255 -631 255 -631 0 cellNo=65
rlabel pdiffusion 262 -631 262 -631 0 cellNo=153
rlabel pdiffusion 325 -631 325 -631 0 cellNo=191
rlabel pdiffusion 31 -664 31 -664 0 feedthrough
rlabel pdiffusion 38 -664 38 -664 0 feedthrough
rlabel pdiffusion 45 -664 45 -664 0 feedthrough
rlabel pdiffusion 52 -664 52 -664 0 feedthrough
rlabel pdiffusion 59 -664 59 -664 0 cellNo=59
rlabel pdiffusion 66 -664 66 -664 0 cellNo=9
rlabel pdiffusion 73 -664 73 -664 0 cellNo=190
rlabel pdiffusion 80 -664 80 -664 0 feedthrough
rlabel pdiffusion 87 -664 87 -664 0 feedthrough
rlabel pdiffusion 94 -664 94 -664 0 cellNo=53
rlabel pdiffusion 101 -664 101 -664 0 feedthrough
rlabel pdiffusion 108 -664 108 -664 0 feedthrough
rlabel pdiffusion 115 -664 115 -664 0 cellNo=387
rlabel pdiffusion 122 -664 122 -664 0 cellNo=247
rlabel pdiffusion 129 -664 129 -664 0 feedthrough
rlabel pdiffusion 136 -664 136 -664 0 cellNo=340
rlabel pdiffusion 143 -664 143 -664 0 cellNo=317
rlabel pdiffusion 150 -664 150 -664 0 feedthrough
rlabel pdiffusion 157 -664 157 -664 0 cellNo=54
rlabel pdiffusion 164 -664 164 -664 0 feedthrough
rlabel pdiffusion 171 -664 171 -664 0 cellNo=143
rlabel pdiffusion 178 -664 178 -664 0 cellNo=349
rlabel pdiffusion 185 -664 185 -664 0 cellNo=332
rlabel pdiffusion 192 -664 192 -664 0 cellNo=63
rlabel pdiffusion 199 -664 199 -664 0 cellNo=385
rlabel pdiffusion 206 -664 206 -664 0 cellNo=202
rlabel pdiffusion 213 -664 213 -664 0 feedthrough
rlabel pdiffusion 220 -664 220 -664 0 feedthrough
rlabel pdiffusion 227 -664 227 -664 0 feedthrough
rlabel pdiffusion 234 -664 234 -664 0 feedthrough
rlabel pdiffusion 241 -664 241 -664 0 feedthrough
rlabel pdiffusion 248 -664 248 -664 0 feedthrough
rlabel pdiffusion 255 -664 255 -664 0 feedthrough
rlabel pdiffusion 262 -664 262 -664 0 feedthrough
rlabel pdiffusion 269 -664 269 -664 0 feedthrough
rlabel pdiffusion 276 -664 276 -664 0 feedthrough
rlabel pdiffusion 283 -664 283 -664 0 feedthrough
rlabel pdiffusion 290 -664 290 -664 0 feedthrough
rlabel pdiffusion 297 -664 297 -664 0 cellNo=121
rlabel pdiffusion 59 -697 59 -697 0 cellNo=189
rlabel pdiffusion 73 -697 73 -697 0 cellNo=302
rlabel pdiffusion 80 -697 80 -697 0 feedthrough
rlabel pdiffusion 87 -697 87 -697 0 cellNo=364
rlabel pdiffusion 94 -697 94 -697 0 feedthrough
rlabel pdiffusion 101 -697 101 -697 0 feedthrough
rlabel pdiffusion 108 -697 108 -697 0 cellNo=18
rlabel pdiffusion 115 -697 115 -697 0 cellNo=321
rlabel pdiffusion 122 -697 122 -697 0 feedthrough
rlabel pdiffusion 129 -697 129 -697 0 feedthrough
rlabel pdiffusion 136 -697 136 -697 0 cellNo=136
rlabel pdiffusion 143 -697 143 -697 0 feedthrough
rlabel pdiffusion 150 -697 150 -697 0 cellNo=80
rlabel pdiffusion 157 -697 157 -697 0 cellNo=203
rlabel pdiffusion 164 -697 164 -697 0 feedthrough
rlabel pdiffusion 171 -697 171 -697 0 feedthrough
rlabel pdiffusion 178 -697 178 -697 0 cellNo=251
rlabel pdiffusion 185 -697 185 -697 0 cellNo=373
rlabel pdiffusion 192 -697 192 -697 0 cellNo=263
rlabel pdiffusion 199 -697 199 -697 0 feedthrough
rlabel pdiffusion 206 -697 206 -697 0 feedthrough
rlabel pdiffusion 213 -697 213 -697 0 cellNo=75
rlabel pdiffusion 220 -697 220 -697 0 feedthrough
rlabel pdiffusion 227 -697 227 -697 0 feedthrough
rlabel pdiffusion 234 -697 234 -697 0 feedthrough
rlabel pdiffusion 241 -697 241 -697 0 feedthrough
rlabel pdiffusion 248 -697 248 -697 0 cellNo=379
rlabel pdiffusion 255 -697 255 -697 0 feedthrough
rlabel pdiffusion 262 -697 262 -697 0 cellNo=174
rlabel pdiffusion 269 -697 269 -697 0 feedthrough
rlabel pdiffusion 276 -697 276 -697 0 cellNo=393
rlabel pdiffusion 115 -720 115 -720 0 cellNo=178
rlabel pdiffusion 122 -720 122 -720 0 feedthrough
rlabel pdiffusion 129 -720 129 -720 0 cellNo=125
rlabel pdiffusion 136 -720 136 -720 0 cellNo=333
rlabel pdiffusion 143 -720 143 -720 0 feedthrough
rlabel pdiffusion 150 -720 150 -720 0 cellNo=352
rlabel pdiffusion 164 -720 164 -720 0 feedthrough
rlabel pdiffusion 171 -720 171 -720 0 cellNo=361
rlabel pdiffusion 178 -720 178 -720 0 cellNo=390
rlabel pdiffusion 185 -720 185 -720 0 feedthrough
rlabel pdiffusion 192 -720 192 -720 0 cellNo=220
rlabel pdiffusion 199 -720 199 -720 0 feedthrough
rlabel pdiffusion 206 -720 206 -720 0 feedthrough
rlabel pdiffusion 213 -720 213 -720 0 cellNo=138
rlabel pdiffusion 227 -720 227 -720 0 cellNo=399
rlabel pdiffusion 241 -720 241 -720 0 feedthrough
rlabel pdiffusion 115 -735 115 -735 0 cellNo=336
rlabel pdiffusion 122 -735 122 -735 0 feedthrough
rlabel pdiffusion 129 -735 129 -735 0 cellNo=372
rlabel pdiffusion 136 -735 136 -735 0 feedthrough
rlabel pdiffusion 157 -735 157 -735 0 cellNo=267
rlabel pdiffusion 164 -735 164 -735 0 cellNo=281
rlabel pdiffusion 171 -735 171 -735 0 feedthrough
rlabel pdiffusion 178 -735 178 -735 0 feedthrough
rlabel pdiffusion 185 -735 185 -735 0 cellNo=397
rlabel pdiffusion 192 -735 192 -735 0 feedthrough
rlabel pdiffusion 122 -748 122 -748 0 cellNo=120
rlabel pdiffusion 129 -748 129 -748 0 feedthrough
rlabel pdiffusion 150 -748 150 -748 0 cellNo=221
rlabel pdiffusion 157 -748 157 -748 0 cellNo=328
rlabel pdiffusion 164 -748 164 -748 0 feedthrough
rlabel pdiffusion 171 -748 171 -748 0 feedthrough
rlabel pdiffusion 185 -748 185 -748 0 feedthrough
rlabel pdiffusion 192 -748 192 -748 0 cellNo=212
rlabel polysilicon 103 -4 103 -4 0 2
rlabel polysilicon 103 -10 103 -10 0 4
rlabel polysilicon 107 -4 107 -4 0 1
rlabel polysilicon 128 -4 128 -4 0 1
rlabel polysilicon 135 -4 135 -4 0 1
rlabel polysilicon 135 -10 135 -10 0 3
rlabel polysilicon 142 -4 142 -4 0 1
rlabel polysilicon 142 -10 142 -10 0 3
rlabel polysilicon 149 -10 149 -10 0 3
rlabel polysilicon 156 -4 156 -4 0 1
rlabel polysilicon 156 -10 156 -10 0 3
rlabel polysilicon 163 -10 163 -10 0 3
rlabel polysilicon 173 -10 173 -10 0 4
rlabel polysilicon 177 -4 177 -4 0 1
rlabel polysilicon 177 -10 177 -10 0 3
rlabel polysilicon 184 -10 184 -10 0 3
rlabel polysilicon 191 -4 191 -4 0 1
rlabel polysilicon 194 -4 194 -4 0 2
rlabel polysilicon 198 -4 198 -4 0 1
rlabel polysilicon 198 -10 198 -10 0 3
rlabel polysilicon 205 -4 205 -4 0 1
rlabel polysilicon 212 -4 212 -4 0 1
rlabel polysilicon 212 -10 212 -10 0 3
rlabel polysilicon 79 -23 79 -23 0 1
rlabel polysilicon 79 -29 79 -29 0 3
rlabel polysilicon 86 -29 86 -29 0 3
rlabel polysilicon 89 -29 89 -29 0 4
rlabel polysilicon 96 -23 96 -23 0 2
rlabel polysilicon 93 -29 93 -29 0 3
rlabel polysilicon 100 -23 100 -23 0 1
rlabel polysilicon 100 -29 100 -29 0 3
rlabel polysilicon 110 -23 110 -23 0 2
rlabel polysilicon 107 -29 107 -29 0 3
rlabel polysilicon 121 -23 121 -23 0 1
rlabel polysilicon 121 -29 121 -29 0 3
rlabel polysilicon 128 -29 128 -29 0 3
rlabel polysilicon 135 -23 135 -23 0 1
rlabel polysilicon 135 -29 135 -29 0 3
rlabel polysilicon 142 -23 142 -23 0 1
rlabel polysilicon 142 -29 142 -29 0 3
rlabel polysilicon 149 -23 149 -23 0 1
rlabel polysilicon 152 -23 152 -23 0 2
rlabel polysilicon 149 -29 149 -29 0 3
rlabel polysilicon 156 -23 156 -23 0 1
rlabel polysilicon 156 -29 156 -29 0 3
rlabel polysilicon 159 -29 159 -29 0 4
rlabel polysilicon 166 -29 166 -29 0 4
rlabel polysilicon 170 -23 170 -23 0 1
rlabel polysilicon 170 -29 170 -29 0 3
rlabel polysilicon 177 -29 177 -29 0 3
rlabel polysilicon 184 -23 184 -23 0 1
rlabel polysilicon 184 -29 184 -29 0 3
rlabel polysilicon 187 -29 187 -29 0 4
rlabel polysilicon 194 -23 194 -23 0 2
rlabel polysilicon 191 -29 191 -29 0 3
rlabel polysilicon 198 -23 198 -23 0 1
rlabel polysilicon 198 -29 198 -29 0 3
rlabel polysilicon 208 -23 208 -23 0 2
rlabel polysilicon 215 -23 215 -23 0 2
rlabel polysilicon 219 -23 219 -23 0 1
rlabel polysilicon 219 -29 219 -29 0 3
rlabel polysilicon 226 -23 226 -23 0 1
rlabel polysilicon 229 -29 229 -29 0 4
rlabel polysilicon 233 -23 233 -23 0 1
rlabel polysilicon 233 -29 233 -29 0 3
rlabel polysilicon 61 -52 61 -52 0 4
rlabel polysilicon 65 -46 65 -46 0 1
rlabel polysilicon 65 -52 65 -52 0 3
rlabel polysilicon 72 -46 72 -46 0 1
rlabel polysilicon 72 -52 72 -52 0 3
rlabel polysilicon 79 -46 79 -46 0 1
rlabel polysilicon 82 -52 82 -52 0 4
rlabel polysilicon 86 -46 86 -46 0 1
rlabel polysilicon 89 -46 89 -46 0 2
rlabel polysilicon 89 -52 89 -52 0 4
rlabel polysilicon 93 -46 93 -46 0 1
rlabel polysilicon 96 -52 96 -52 0 4
rlabel polysilicon 100 -46 100 -46 0 1
rlabel polysilicon 100 -52 100 -52 0 3
rlabel polysilicon 110 -46 110 -46 0 2
rlabel polysilicon 110 -52 110 -52 0 4
rlabel polysilicon 114 -46 114 -46 0 1
rlabel polysilicon 114 -52 114 -52 0 3
rlabel polysilicon 121 -52 121 -52 0 3
rlabel polysilicon 124 -52 124 -52 0 4
rlabel polysilicon 128 -46 128 -46 0 1
rlabel polysilicon 131 -52 131 -52 0 4
rlabel polysilicon 135 -46 135 -46 0 1
rlabel polysilicon 135 -52 135 -52 0 3
rlabel polysilicon 142 -52 142 -52 0 3
rlabel polysilicon 145 -52 145 -52 0 4
rlabel polysilicon 149 -46 149 -46 0 1
rlabel polysilicon 152 -46 152 -46 0 2
rlabel polysilicon 156 -46 156 -46 0 1
rlabel polysilicon 156 -52 156 -52 0 3
rlabel polysilicon 163 -46 163 -46 0 1
rlabel polysilicon 163 -52 163 -52 0 3
rlabel polysilicon 170 -46 170 -46 0 1
rlabel polysilicon 173 -46 173 -46 0 2
rlabel polysilicon 170 -52 170 -52 0 3
rlabel polysilicon 180 -46 180 -46 0 2
rlabel polysilicon 184 -46 184 -46 0 1
rlabel polysilicon 184 -52 184 -52 0 3
rlabel polysilicon 191 -46 191 -46 0 1
rlabel polysilicon 191 -52 191 -52 0 3
rlabel polysilicon 201 -46 201 -46 0 2
rlabel polysilicon 198 -52 198 -52 0 3
rlabel polysilicon 201 -52 201 -52 0 4
rlabel polysilicon 205 -46 205 -46 0 1
rlabel polysilicon 205 -52 205 -52 0 3
rlabel polysilicon 215 -46 215 -46 0 2
rlabel polysilicon 212 -52 212 -52 0 3
rlabel polysilicon 219 -46 219 -46 0 1
rlabel polysilicon 222 -52 222 -52 0 4
rlabel polysilicon 226 -46 226 -46 0 1
rlabel polysilicon 226 -52 226 -52 0 3
rlabel polysilicon 233 -46 233 -46 0 1
rlabel polysilicon 233 -52 233 -52 0 3
rlabel polysilicon 240 -46 240 -46 0 1
rlabel polysilicon 240 -52 240 -52 0 3
rlabel polysilicon 247 -46 247 -46 0 1
rlabel polysilicon 247 -52 247 -52 0 3
rlabel polysilicon 254 -46 254 -46 0 1
rlabel polysilicon 254 -52 254 -52 0 3
rlabel polysilicon 261 -46 261 -46 0 1
rlabel polysilicon 261 -52 261 -52 0 3
rlabel polysilicon 271 -46 271 -46 0 2
rlabel polysilicon 275 -46 275 -46 0 1
rlabel polysilicon 275 -52 275 -52 0 3
rlabel polysilicon 282 -46 282 -46 0 1
rlabel polysilicon 282 -52 282 -52 0 3
rlabel polysilicon 30 -77 30 -77 0 1
rlabel polysilicon 30 -83 30 -83 0 3
rlabel polysilicon 37 -83 37 -83 0 3
rlabel polysilicon 44 -77 44 -77 0 1
rlabel polysilicon 44 -83 44 -83 0 3
rlabel polysilicon 51 -77 51 -77 0 1
rlabel polysilicon 51 -83 51 -83 0 3
rlabel polysilicon 58 -77 58 -77 0 1
rlabel polysilicon 58 -83 58 -83 0 3
rlabel polysilicon 65 -77 65 -77 0 1
rlabel polysilicon 65 -83 65 -83 0 3
rlabel polysilicon 72 -77 72 -77 0 1
rlabel polysilicon 75 -77 75 -77 0 2
rlabel polysilicon 79 -77 79 -77 0 1
rlabel polysilicon 79 -83 79 -83 0 3
rlabel polysilicon 86 -77 86 -77 0 1
rlabel polysilicon 86 -83 86 -83 0 3
rlabel polysilicon 93 -77 93 -77 0 1
rlabel polysilicon 93 -83 93 -83 0 3
rlabel polysilicon 100 -77 100 -77 0 1
rlabel polysilicon 103 -77 103 -77 0 2
rlabel polysilicon 100 -83 100 -83 0 3
rlabel polysilicon 107 -83 107 -83 0 3
rlabel polysilicon 110 -83 110 -83 0 4
rlabel polysilicon 114 -77 114 -77 0 1
rlabel polysilicon 117 -77 117 -77 0 2
rlabel polysilicon 114 -83 114 -83 0 3
rlabel polysilicon 117 -83 117 -83 0 4
rlabel polysilicon 121 -77 121 -77 0 1
rlabel polysilicon 121 -83 121 -83 0 3
rlabel polysilicon 128 -83 128 -83 0 3
rlabel polysilicon 135 -77 135 -77 0 1
rlabel polysilicon 138 -77 138 -77 0 2
rlabel polysilicon 138 -83 138 -83 0 4
rlabel polysilicon 142 -77 142 -77 0 1
rlabel polysilicon 142 -83 142 -83 0 3
rlabel polysilicon 149 -77 149 -77 0 1
rlabel polysilicon 149 -83 149 -83 0 3
rlabel polysilicon 156 -77 156 -77 0 1
rlabel polysilicon 159 -77 159 -77 0 2
rlabel polysilicon 163 -77 163 -77 0 1
rlabel polysilicon 163 -83 163 -83 0 3
rlabel polysilicon 170 -77 170 -77 0 1
rlabel polysilicon 170 -83 170 -83 0 3
rlabel polysilicon 177 -77 177 -77 0 1
rlabel polysilicon 180 -77 180 -77 0 2
rlabel polysilicon 177 -83 177 -83 0 3
rlabel polysilicon 180 -83 180 -83 0 4
rlabel polysilicon 184 -77 184 -77 0 1
rlabel polysilicon 187 -77 187 -77 0 2
rlabel polysilicon 187 -83 187 -83 0 4
rlabel polysilicon 191 -77 191 -77 0 1
rlabel polysilicon 191 -83 191 -83 0 3
rlabel polysilicon 198 -77 198 -77 0 1
rlabel polysilicon 198 -83 198 -83 0 3
rlabel polysilicon 201 -83 201 -83 0 4
rlabel polysilicon 205 -83 205 -83 0 3
rlabel polysilicon 208 -83 208 -83 0 4
rlabel polysilicon 212 -77 212 -77 0 1
rlabel polysilicon 219 -77 219 -77 0 1
rlabel polysilicon 219 -83 219 -83 0 3
rlabel polysilicon 226 -77 226 -77 0 1
rlabel polysilicon 226 -83 226 -83 0 3
rlabel polysilicon 233 -77 233 -77 0 1
rlabel polysilicon 233 -83 233 -83 0 3
rlabel polysilicon 243 -77 243 -77 0 2
rlabel polysilicon 243 -83 243 -83 0 4
rlabel polysilicon 250 -83 250 -83 0 4
rlabel polysilicon 254 -77 254 -77 0 1
rlabel polysilicon 254 -83 254 -83 0 3
rlabel polysilicon 261 -77 261 -77 0 1
rlabel polysilicon 261 -83 261 -83 0 3
rlabel polysilicon 268 -77 268 -77 0 1
rlabel polysilicon 268 -83 268 -83 0 3
rlabel polysilicon 275 -77 275 -77 0 1
rlabel polysilicon 275 -83 275 -83 0 3
rlabel polysilicon 282 -77 282 -77 0 1
rlabel polysilicon 282 -83 282 -83 0 3
rlabel polysilicon 289 -77 289 -77 0 1
rlabel polysilicon 289 -83 289 -83 0 3
rlabel polysilicon 299 -83 299 -83 0 4
rlabel polysilicon 303 -77 303 -77 0 1
rlabel polysilicon 303 -83 303 -83 0 3
rlabel polysilicon 16 -122 16 -122 0 1
rlabel polysilicon 16 -128 16 -128 0 3
rlabel polysilicon 26 -122 26 -122 0 2
rlabel polysilicon 23 -128 23 -128 0 3
rlabel polysilicon 30 -122 30 -122 0 1
rlabel polysilicon 30 -128 30 -128 0 3
rlabel polysilicon 37 -122 37 -122 0 1
rlabel polysilicon 37 -128 37 -128 0 3
rlabel polysilicon 47 -128 47 -128 0 4
rlabel polysilicon 51 -122 51 -122 0 1
rlabel polysilicon 51 -128 51 -128 0 3
rlabel polysilicon 61 -128 61 -128 0 4
rlabel polysilicon 65 -122 65 -122 0 1
rlabel polysilicon 68 -122 68 -122 0 2
rlabel polysilicon 65 -128 65 -128 0 3
rlabel polysilicon 72 -122 72 -122 0 1
rlabel polysilicon 72 -128 72 -128 0 3
rlabel polysilicon 79 -122 79 -122 0 1
rlabel polysilicon 79 -128 79 -128 0 3
rlabel polysilicon 82 -128 82 -128 0 4
rlabel polysilicon 86 -122 86 -122 0 1
rlabel polysilicon 86 -128 86 -128 0 3
rlabel polysilicon 93 -122 93 -122 0 1
rlabel polysilicon 93 -128 93 -128 0 3
rlabel polysilicon 100 -122 100 -122 0 1
rlabel polysilicon 103 -122 103 -122 0 2
rlabel polysilicon 100 -128 100 -128 0 3
rlabel polysilicon 103 -128 103 -128 0 4
rlabel polysilicon 107 -122 107 -122 0 1
rlabel polysilicon 107 -128 107 -128 0 3
rlabel polysilicon 117 -122 117 -122 0 2
rlabel polysilicon 114 -128 114 -128 0 3
rlabel polysilicon 117 -128 117 -128 0 4
rlabel polysilicon 124 -122 124 -122 0 2
rlabel polysilicon 128 -122 128 -122 0 1
rlabel polysilicon 131 -122 131 -122 0 2
rlabel polysilicon 128 -128 128 -128 0 3
rlabel polysilicon 131 -128 131 -128 0 4
rlabel polysilicon 135 -122 135 -122 0 1
rlabel polysilicon 138 -122 138 -122 0 2
rlabel polysilicon 135 -128 135 -128 0 3
rlabel polysilicon 142 -128 142 -128 0 3
rlabel polysilicon 145 -128 145 -128 0 4
rlabel polysilicon 149 -122 149 -122 0 1
rlabel polysilicon 152 -122 152 -122 0 2
rlabel polysilicon 152 -128 152 -128 0 4
rlabel polysilicon 159 -122 159 -122 0 2
rlabel polysilicon 156 -128 156 -128 0 3
rlabel polysilicon 159 -128 159 -128 0 4
rlabel polysilicon 170 -122 170 -122 0 1
rlabel polysilicon 170 -128 170 -128 0 3
rlabel polysilicon 180 -122 180 -122 0 2
rlabel polysilicon 177 -128 177 -128 0 3
rlabel polysilicon 180 -128 180 -128 0 4
rlabel polysilicon 184 -122 184 -122 0 1
rlabel polysilicon 187 -122 187 -122 0 2
rlabel polysilicon 184 -128 184 -128 0 3
rlabel polysilicon 187 -128 187 -128 0 4
rlabel polysilicon 194 -122 194 -122 0 2
rlabel polysilicon 198 -122 198 -122 0 1
rlabel polysilicon 201 -122 201 -122 0 2
rlabel polysilicon 198 -128 198 -128 0 3
rlabel polysilicon 201 -128 201 -128 0 4
rlabel polysilicon 205 -122 205 -122 0 1
rlabel polysilicon 208 -122 208 -122 0 2
rlabel polysilicon 205 -128 205 -128 0 3
rlabel polysilicon 212 -122 212 -122 0 1
rlabel polysilicon 212 -128 212 -128 0 3
rlabel polysilicon 219 -122 219 -122 0 1
rlabel polysilicon 219 -128 219 -128 0 3
rlabel polysilicon 226 -122 226 -122 0 1
rlabel polysilicon 226 -128 226 -128 0 3
rlabel polysilicon 236 -122 236 -122 0 2
rlabel polysilicon 233 -128 233 -128 0 3
rlabel polysilicon 236 -128 236 -128 0 4
rlabel polysilicon 240 -122 240 -122 0 1
rlabel polysilicon 240 -128 240 -128 0 3
rlabel polysilicon 247 -122 247 -122 0 1
rlabel polysilicon 247 -128 247 -128 0 3
rlabel polysilicon 254 -122 254 -122 0 1
rlabel polysilicon 254 -128 254 -128 0 3
rlabel polysilicon 261 -122 261 -122 0 1
rlabel polysilicon 261 -128 261 -128 0 3
rlabel polysilicon 268 -122 268 -122 0 1
rlabel polysilicon 268 -128 268 -128 0 3
rlabel polysilicon 275 -122 275 -122 0 1
rlabel polysilicon 275 -128 275 -128 0 3
rlabel polysilicon 282 -122 282 -122 0 1
rlabel polysilicon 282 -128 282 -128 0 3
rlabel polysilicon 289 -122 289 -122 0 1
rlabel polysilicon 289 -128 289 -128 0 3
rlabel polysilicon 296 -122 296 -122 0 1
rlabel polysilicon 296 -128 296 -128 0 3
rlabel polysilicon 303 -122 303 -122 0 1
rlabel polysilicon 303 -128 303 -128 0 3
rlabel polysilicon 310 -122 310 -122 0 1
rlabel polysilicon 310 -128 310 -128 0 3
rlabel polysilicon 317 -122 317 -122 0 1
rlabel polysilicon 317 -128 317 -128 0 3
rlabel polysilicon 324 -122 324 -122 0 1
rlabel polysilicon 324 -128 324 -128 0 3
rlabel polysilicon 331 -122 331 -122 0 1
rlabel polysilicon 331 -128 331 -128 0 3
rlabel polysilicon 19 -175 19 -175 0 4
rlabel polysilicon 23 -169 23 -169 0 1
rlabel polysilicon 26 -169 26 -169 0 2
rlabel polysilicon 30 -169 30 -169 0 1
rlabel polysilicon 30 -175 30 -175 0 3
rlabel polysilicon 37 -169 37 -169 0 1
rlabel polysilicon 44 -169 44 -169 0 1
rlabel polysilicon 44 -175 44 -175 0 3
rlabel polysilicon 51 -175 51 -175 0 3
rlabel polysilicon 61 -169 61 -169 0 2
rlabel polysilicon 58 -175 58 -175 0 3
rlabel polysilicon 65 -169 65 -169 0 1
rlabel polysilicon 65 -175 65 -175 0 3
rlabel polysilicon 72 -169 72 -169 0 1
rlabel polysilicon 72 -175 72 -175 0 3
rlabel polysilicon 79 -169 79 -169 0 1
rlabel polysilicon 79 -175 79 -175 0 3
rlabel polysilicon 89 -169 89 -169 0 2
rlabel polysilicon 86 -175 86 -175 0 3
rlabel polysilicon 93 -169 93 -169 0 1
rlabel polysilicon 93 -175 93 -175 0 3
rlabel polysilicon 100 -169 100 -169 0 1
rlabel polysilicon 100 -175 100 -175 0 3
rlabel polysilicon 110 -169 110 -169 0 2
rlabel polysilicon 107 -175 107 -175 0 3
rlabel polysilicon 110 -175 110 -175 0 4
rlabel polysilicon 114 -169 114 -169 0 1
rlabel polysilicon 117 -169 117 -169 0 2
rlabel polysilicon 117 -175 117 -175 0 4
rlabel polysilicon 124 -169 124 -169 0 2
rlabel polysilicon 124 -175 124 -175 0 4
rlabel polysilicon 128 -169 128 -169 0 1
rlabel polysilicon 128 -175 128 -175 0 3
rlabel polysilicon 135 -175 135 -175 0 3
rlabel polysilicon 142 -169 142 -169 0 1
rlabel polysilicon 142 -175 142 -175 0 3
rlabel polysilicon 152 -169 152 -169 0 2
rlabel polysilicon 149 -175 149 -175 0 3
rlabel polysilicon 159 -169 159 -169 0 2
rlabel polysilicon 156 -175 156 -175 0 3
rlabel polysilicon 159 -175 159 -175 0 4
rlabel polysilicon 166 -169 166 -169 0 2
rlabel polysilicon 170 -169 170 -169 0 1
rlabel polysilicon 170 -175 170 -175 0 3
rlabel polysilicon 177 -169 177 -169 0 1
rlabel polysilicon 177 -175 177 -175 0 3
rlabel polysilicon 184 -169 184 -169 0 1
rlabel polysilicon 184 -175 184 -175 0 3
rlabel polysilicon 194 -169 194 -169 0 2
rlabel polysilicon 194 -175 194 -175 0 4
rlabel polysilicon 201 -169 201 -169 0 2
rlabel polysilicon 201 -175 201 -175 0 4
rlabel polysilicon 205 -169 205 -169 0 1
rlabel polysilicon 205 -175 205 -175 0 3
rlabel polysilicon 208 -175 208 -175 0 4
rlabel polysilicon 212 -169 212 -169 0 1
rlabel polysilicon 215 -169 215 -169 0 2
rlabel polysilicon 219 -169 219 -169 0 1
rlabel polysilicon 219 -175 219 -175 0 3
rlabel polysilicon 226 -169 226 -169 0 1
rlabel polysilicon 226 -175 226 -175 0 3
rlabel polysilicon 233 -169 233 -169 0 1
rlabel polysilicon 236 -169 236 -169 0 2
rlabel polysilicon 243 -169 243 -169 0 2
rlabel polysilicon 240 -175 240 -175 0 3
rlabel polysilicon 243 -175 243 -175 0 4
rlabel polysilicon 247 -169 247 -169 0 1
rlabel polysilicon 247 -175 247 -175 0 3
rlabel polysilicon 254 -169 254 -169 0 1
rlabel polysilicon 254 -175 254 -175 0 3
rlabel polysilicon 261 -169 261 -169 0 1
rlabel polysilicon 261 -175 261 -175 0 3
rlabel polysilicon 268 -175 268 -175 0 3
rlabel polysilicon 275 -169 275 -169 0 1
rlabel polysilicon 275 -175 275 -175 0 3
rlabel polysilicon 282 -169 282 -169 0 1
rlabel polysilicon 282 -175 282 -175 0 3
rlabel polysilicon 289 -169 289 -169 0 1
rlabel polysilicon 289 -175 289 -175 0 3
rlabel polysilicon 296 -169 296 -169 0 1
rlabel polysilicon 296 -175 296 -175 0 3
rlabel polysilicon 303 -169 303 -169 0 1
rlabel polysilicon 303 -175 303 -175 0 3
rlabel polysilicon 310 -169 310 -169 0 1
rlabel polysilicon 310 -175 310 -175 0 3
rlabel polysilicon 9 -206 9 -206 0 1
rlabel polysilicon 9 -212 9 -212 0 3
rlabel polysilicon 16 -206 16 -206 0 1
rlabel polysilicon 16 -212 16 -212 0 3
rlabel polysilicon 23 -206 23 -206 0 1
rlabel polysilicon 33 -206 33 -206 0 2
rlabel polysilicon 37 -206 37 -206 0 1
rlabel polysilicon 37 -212 37 -212 0 3
rlabel polysilicon 44 -206 44 -206 0 1
rlabel polysilicon 44 -212 44 -212 0 3
rlabel polysilicon 51 -206 51 -206 0 1
rlabel polysilicon 54 -206 54 -206 0 2
rlabel polysilicon 54 -212 54 -212 0 4
rlabel polysilicon 58 -206 58 -206 0 1
rlabel polysilicon 58 -212 58 -212 0 3
rlabel polysilicon 68 -206 68 -206 0 2
rlabel polysilicon 72 -206 72 -206 0 1
rlabel polysilicon 72 -212 72 -212 0 3
rlabel polysilicon 75 -212 75 -212 0 4
rlabel polysilicon 79 -206 79 -206 0 1
rlabel polysilicon 79 -212 79 -212 0 3
rlabel polysilicon 86 -206 86 -206 0 1
rlabel polysilicon 89 -206 89 -206 0 2
rlabel polysilicon 89 -212 89 -212 0 4
rlabel polysilicon 93 -206 93 -206 0 1
rlabel polysilicon 93 -212 93 -212 0 3
rlabel polysilicon 100 -206 100 -206 0 1
rlabel polysilicon 100 -212 100 -212 0 3
rlabel polysilicon 107 -206 107 -206 0 1
rlabel polysilicon 110 -212 110 -212 0 4
rlabel polysilicon 114 -206 114 -206 0 1
rlabel polysilicon 117 -206 117 -206 0 2
rlabel polysilicon 114 -212 114 -212 0 3
rlabel polysilicon 117 -212 117 -212 0 4
rlabel polysilicon 121 -206 121 -206 0 1
rlabel polysilicon 121 -212 121 -212 0 3
rlabel polysilicon 128 -206 128 -206 0 1
rlabel polysilicon 128 -212 128 -212 0 3
rlabel polysilicon 135 -206 135 -206 0 1
rlabel polysilicon 135 -212 135 -212 0 3
rlabel polysilicon 145 -206 145 -206 0 2
rlabel polysilicon 142 -212 142 -212 0 3
rlabel polysilicon 149 -206 149 -206 0 1
rlabel polysilicon 149 -212 149 -212 0 3
rlabel polysilicon 156 -206 156 -206 0 1
rlabel polysilicon 156 -212 156 -212 0 3
rlabel polysilicon 163 -206 163 -206 0 1
rlabel polysilicon 163 -212 163 -212 0 3
rlabel polysilicon 170 -206 170 -206 0 1
rlabel polysilicon 170 -212 170 -212 0 3
rlabel polysilicon 177 -206 177 -206 0 1
rlabel polysilicon 177 -212 177 -212 0 3
rlabel polysilicon 184 -206 184 -206 0 1
rlabel polysilicon 187 -212 187 -212 0 4
rlabel polysilicon 191 -206 191 -206 0 1
rlabel polysilicon 191 -212 191 -212 0 3
rlabel polysilicon 198 -206 198 -206 0 1
rlabel polysilicon 198 -212 198 -212 0 3
rlabel polysilicon 205 -206 205 -206 0 1
rlabel polysilicon 208 -212 208 -212 0 4
rlabel polysilicon 212 -206 212 -206 0 1
rlabel polysilicon 215 -206 215 -206 0 2
rlabel polysilicon 215 -212 215 -212 0 4
rlabel polysilicon 219 -206 219 -206 0 1
rlabel polysilicon 222 -206 222 -206 0 2
rlabel polysilicon 219 -212 219 -212 0 3
rlabel polysilicon 222 -212 222 -212 0 4
rlabel polysilicon 226 -206 226 -206 0 1
rlabel polysilicon 226 -212 226 -212 0 3
rlabel polysilicon 236 -206 236 -206 0 2
rlabel polysilicon 233 -212 233 -212 0 3
rlabel polysilicon 240 -206 240 -206 0 1
rlabel polysilicon 240 -212 240 -212 0 3
rlabel polysilicon 247 -206 247 -206 0 1
rlabel polysilicon 247 -212 247 -212 0 3
rlabel polysilicon 254 -206 254 -206 0 1
rlabel polysilicon 254 -212 254 -212 0 3
rlabel polysilicon 261 -206 261 -206 0 1
rlabel polysilicon 261 -212 261 -212 0 3
rlabel polysilicon 271 -206 271 -206 0 2
rlabel polysilicon 268 -212 268 -212 0 3
rlabel polysilicon 275 -206 275 -206 0 1
rlabel polysilicon 275 -212 275 -212 0 3
rlabel polysilicon 285 -206 285 -206 0 2
rlabel polysilicon 285 -212 285 -212 0 4
rlabel polysilicon 289 -206 289 -206 0 1
rlabel polysilicon 292 -206 292 -206 0 2
rlabel polysilicon 296 -206 296 -206 0 1
rlabel polysilicon 296 -212 296 -212 0 3
rlabel polysilicon 303 -206 303 -206 0 1
rlabel polysilicon 303 -212 303 -212 0 3
rlabel polysilicon 310 -206 310 -206 0 1
rlabel polysilicon 310 -212 310 -212 0 3
rlabel polysilicon 317 -206 317 -206 0 1
rlabel polysilicon 317 -212 317 -212 0 3
rlabel polysilicon 324 -206 324 -206 0 1
rlabel polysilicon 324 -212 324 -212 0 3
rlabel polysilicon 331 -206 331 -206 0 1
rlabel polysilicon 331 -212 331 -212 0 3
rlabel polysilicon 338 -206 338 -206 0 1
rlabel polysilicon 338 -212 338 -212 0 3
rlabel polysilicon 345 -206 345 -206 0 1
rlabel polysilicon 345 -212 345 -212 0 3
rlabel polysilicon 352 -206 352 -206 0 1
rlabel polysilicon 352 -212 352 -212 0 3
rlabel polysilicon 359 -206 359 -206 0 1
rlabel polysilicon 359 -212 359 -212 0 3
rlabel polysilicon 366 -206 366 -206 0 1
rlabel polysilicon 366 -212 366 -212 0 3
rlabel polysilicon 373 -206 373 -206 0 1
rlabel polysilicon 373 -212 373 -212 0 3
rlabel polysilicon 380 -206 380 -206 0 1
rlabel polysilicon 380 -212 380 -212 0 3
rlabel polysilicon 387 -206 387 -206 0 1
rlabel polysilicon 394 -206 394 -206 0 1
rlabel polysilicon 394 -212 394 -212 0 3
rlabel polysilicon 9 -251 9 -251 0 1
rlabel polysilicon 9 -257 9 -257 0 3
rlabel polysilicon 16 -251 16 -251 0 1
rlabel polysilicon 16 -257 16 -257 0 3
rlabel polysilicon 26 -251 26 -251 0 2
rlabel polysilicon 30 -251 30 -251 0 1
rlabel polysilicon 30 -257 30 -257 0 3
rlabel polysilicon 37 -251 37 -251 0 1
rlabel polysilicon 37 -257 37 -257 0 3
rlabel polysilicon 44 -251 44 -251 0 1
rlabel polysilicon 44 -257 44 -257 0 3
rlabel polysilicon 51 -251 51 -251 0 1
rlabel polysilicon 51 -257 51 -257 0 3
rlabel polysilicon 58 -251 58 -251 0 1
rlabel polysilicon 58 -257 58 -257 0 3
rlabel polysilicon 68 -257 68 -257 0 4
rlabel polysilicon 72 -251 72 -251 0 1
rlabel polysilicon 72 -257 72 -257 0 3
rlabel polysilicon 75 -257 75 -257 0 4
rlabel polysilicon 79 -251 79 -251 0 1
rlabel polysilicon 82 -251 82 -251 0 2
rlabel polysilicon 82 -257 82 -257 0 4
rlabel polysilicon 86 -251 86 -251 0 1
rlabel polysilicon 86 -257 86 -257 0 3
rlabel polysilicon 93 -251 93 -251 0 1
rlabel polysilicon 93 -257 93 -257 0 3
rlabel polysilicon 100 -257 100 -257 0 3
rlabel polysilicon 103 -257 103 -257 0 4
rlabel polysilicon 110 -251 110 -251 0 2
rlabel polysilicon 107 -257 107 -257 0 3
rlabel polysilicon 114 -251 114 -251 0 1
rlabel polysilicon 114 -257 114 -257 0 3
rlabel polysilicon 121 -251 121 -251 0 1
rlabel polysilicon 124 -251 124 -251 0 2
rlabel polysilicon 124 -257 124 -257 0 4
rlabel polysilicon 128 -251 128 -251 0 1
rlabel polysilicon 128 -257 128 -257 0 3
rlabel polysilicon 135 -257 135 -257 0 3
rlabel polysilicon 138 -257 138 -257 0 4
rlabel polysilicon 142 -251 142 -251 0 1
rlabel polysilicon 142 -257 142 -257 0 3
rlabel polysilicon 152 -251 152 -251 0 2
rlabel polysilicon 152 -257 152 -257 0 4
rlabel polysilicon 156 -251 156 -251 0 1
rlabel polysilicon 159 -251 159 -251 0 2
rlabel polysilicon 159 -257 159 -257 0 4
rlabel polysilicon 163 -251 163 -251 0 1
rlabel polysilicon 163 -257 163 -257 0 3
rlabel polysilicon 170 -251 170 -251 0 1
rlabel polysilicon 170 -257 170 -257 0 3
rlabel polysilicon 177 -251 177 -251 0 1
rlabel polysilicon 177 -257 177 -257 0 3
rlabel polysilicon 184 -251 184 -251 0 1
rlabel polysilicon 184 -257 184 -257 0 3
rlabel polysilicon 191 -251 191 -251 0 1
rlabel polysilicon 191 -257 191 -257 0 3
rlabel polysilicon 198 -251 198 -251 0 1
rlabel polysilicon 201 -251 201 -251 0 2
rlabel polysilicon 198 -257 198 -257 0 3
rlabel polysilicon 201 -257 201 -257 0 4
rlabel polysilicon 208 -251 208 -251 0 2
rlabel polysilicon 205 -257 205 -257 0 3
rlabel polysilicon 208 -257 208 -257 0 4
rlabel polysilicon 212 -251 212 -251 0 1
rlabel polysilicon 215 -251 215 -251 0 2
rlabel polysilicon 215 -257 215 -257 0 4
rlabel polysilicon 219 -251 219 -251 0 1
rlabel polysilicon 219 -257 219 -257 0 3
rlabel polysilicon 226 -251 226 -251 0 1
rlabel polysilicon 229 -251 229 -251 0 2
rlabel polysilicon 226 -257 226 -257 0 3
rlabel polysilicon 233 -251 233 -251 0 1
rlabel polysilicon 233 -257 233 -257 0 3
rlabel polysilicon 240 -251 240 -251 0 1
rlabel polysilicon 240 -257 240 -257 0 3
rlabel polysilicon 247 -251 247 -251 0 1
rlabel polysilicon 247 -257 247 -257 0 3
rlabel polysilicon 254 -251 254 -251 0 1
rlabel polysilicon 254 -257 254 -257 0 3
rlabel polysilicon 264 -257 264 -257 0 4
rlabel polysilicon 268 -251 268 -251 0 1
rlabel polysilicon 268 -257 268 -257 0 3
rlabel polysilicon 275 -251 275 -251 0 1
rlabel polysilicon 275 -257 275 -257 0 3
rlabel polysilicon 282 -251 282 -251 0 1
rlabel polysilicon 282 -257 282 -257 0 3
rlabel polysilicon 289 -251 289 -251 0 1
rlabel polysilicon 292 -251 292 -251 0 2
rlabel polysilicon 289 -257 289 -257 0 3
rlabel polysilicon 296 -251 296 -251 0 1
rlabel polysilicon 296 -257 296 -257 0 3
rlabel polysilicon 303 -251 303 -251 0 1
rlabel polysilicon 303 -257 303 -257 0 3
rlabel polysilicon 310 -251 310 -251 0 1
rlabel polysilicon 310 -257 310 -257 0 3
rlabel polysilicon 317 -251 317 -251 0 1
rlabel polysilicon 317 -257 317 -257 0 3
rlabel polysilicon 324 -251 324 -251 0 1
rlabel polysilicon 324 -257 324 -257 0 3
rlabel polysilicon 331 -251 331 -251 0 1
rlabel polysilicon 331 -257 331 -257 0 3
rlabel polysilicon 338 -251 338 -251 0 1
rlabel polysilicon 338 -257 338 -257 0 3
rlabel polysilicon 345 -251 345 -251 0 1
rlabel polysilicon 345 -257 345 -257 0 3
rlabel polysilicon 352 -251 352 -251 0 1
rlabel polysilicon 352 -257 352 -257 0 3
rlabel polysilicon 359 -251 359 -251 0 1
rlabel polysilicon 359 -257 359 -257 0 3
rlabel polysilicon 366 -257 366 -257 0 3
rlabel polysilicon 369 -257 369 -257 0 4
rlabel polysilicon 373 -251 373 -251 0 1
rlabel polysilicon 380 -251 380 -251 0 1
rlabel polysilicon 380 -257 380 -257 0 3
rlabel polysilicon 2 -298 2 -298 0 1
rlabel polysilicon 2 -304 2 -304 0 3
rlabel polysilicon 9 -298 9 -298 0 1
rlabel polysilicon 9 -304 9 -304 0 3
rlabel polysilicon 16 -298 16 -298 0 1
rlabel polysilicon 16 -304 16 -304 0 3
rlabel polysilicon 23 -298 23 -298 0 1
rlabel polysilicon 23 -304 23 -304 0 3
rlabel polysilicon 30 -298 30 -298 0 1
rlabel polysilicon 30 -304 30 -304 0 3
rlabel polysilicon 37 -298 37 -298 0 1
rlabel polysilicon 37 -304 37 -304 0 3
rlabel polysilicon 44 -298 44 -298 0 1
rlabel polysilicon 44 -304 44 -304 0 3
rlabel polysilicon 51 -298 51 -298 0 1
rlabel polysilicon 54 -298 54 -298 0 2
rlabel polysilicon 61 -298 61 -298 0 2
rlabel polysilicon 61 -304 61 -304 0 4
rlabel polysilicon 65 -298 65 -298 0 1
rlabel polysilicon 65 -304 65 -304 0 3
rlabel polysilicon 72 -298 72 -298 0 1
rlabel polysilicon 72 -304 72 -304 0 3
rlabel polysilicon 79 -298 79 -298 0 1
rlabel polysilicon 82 -304 82 -304 0 4
rlabel polysilicon 86 -298 86 -298 0 1
rlabel polysilicon 86 -304 86 -304 0 3
rlabel polysilicon 93 -298 93 -298 0 1
rlabel polysilicon 93 -304 93 -304 0 3
rlabel polysilicon 100 -298 100 -298 0 1
rlabel polysilicon 100 -304 100 -304 0 3
rlabel polysilicon 107 -298 107 -298 0 1
rlabel polysilicon 107 -304 107 -304 0 3
rlabel polysilicon 114 -298 114 -298 0 1
rlabel polysilicon 114 -304 114 -304 0 3
rlabel polysilicon 121 -298 121 -298 0 1
rlabel polysilicon 124 -298 124 -298 0 2
rlabel polysilicon 124 -304 124 -304 0 4
rlabel polysilicon 128 -298 128 -298 0 1
rlabel polysilicon 128 -304 128 -304 0 3
rlabel polysilicon 135 -304 135 -304 0 3
rlabel polysilicon 138 -304 138 -304 0 4
rlabel polysilicon 142 -298 142 -298 0 1
rlabel polysilicon 142 -304 142 -304 0 3
rlabel polysilicon 149 -298 149 -298 0 1
rlabel polysilicon 149 -304 149 -304 0 3
rlabel polysilicon 156 -298 156 -298 0 1
rlabel polysilicon 159 -298 159 -298 0 2
rlabel polysilicon 156 -304 156 -304 0 3
rlabel polysilicon 159 -304 159 -304 0 4
rlabel polysilicon 166 -298 166 -298 0 2
rlabel polysilicon 163 -304 163 -304 0 3
rlabel polysilicon 166 -304 166 -304 0 4
rlabel polysilicon 170 -298 170 -298 0 1
rlabel polysilicon 170 -304 170 -304 0 3
rlabel polysilicon 177 -298 177 -298 0 1
rlabel polysilicon 177 -304 177 -304 0 3
rlabel polysilicon 184 -298 184 -298 0 1
rlabel polysilicon 187 -298 187 -298 0 2
rlabel polysilicon 187 -304 187 -304 0 4
rlabel polysilicon 191 -298 191 -298 0 1
rlabel polysilicon 191 -304 191 -304 0 3
rlabel polysilicon 198 -298 198 -298 0 1
rlabel polysilicon 201 -298 201 -298 0 2
rlabel polysilicon 201 -304 201 -304 0 4
rlabel polysilicon 205 -298 205 -298 0 1
rlabel polysilicon 208 -298 208 -298 0 2
rlabel polysilicon 208 -304 208 -304 0 4
rlabel polysilicon 212 -298 212 -298 0 1
rlabel polysilicon 215 -298 215 -298 0 2
rlabel polysilicon 212 -304 212 -304 0 3
rlabel polysilicon 215 -304 215 -304 0 4
rlabel polysilicon 219 -298 219 -298 0 1
rlabel polysilicon 219 -304 219 -304 0 3
rlabel polysilicon 226 -298 226 -298 0 1
rlabel polysilicon 226 -304 226 -304 0 3
rlabel polysilicon 233 -304 233 -304 0 3
rlabel polysilicon 236 -304 236 -304 0 4
rlabel polysilicon 240 -298 240 -298 0 1
rlabel polysilicon 240 -304 240 -304 0 3
rlabel polysilicon 243 -304 243 -304 0 4
rlabel polysilicon 247 -298 247 -298 0 1
rlabel polysilicon 250 -298 250 -298 0 2
rlabel polysilicon 250 -304 250 -304 0 4
rlabel polysilicon 257 -298 257 -298 0 2
rlabel polysilicon 254 -304 254 -304 0 3
rlabel polysilicon 261 -298 261 -298 0 1
rlabel polysilicon 261 -304 261 -304 0 3
rlabel polysilicon 268 -298 268 -298 0 1
rlabel polysilicon 268 -304 268 -304 0 3
rlabel polysilicon 275 -298 275 -298 0 1
rlabel polysilicon 275 -304 275 -304 0 3
rlabel polysilicon 282 -298 282 -298 0 1
rlabel polysilicon 282 -304 282 -304 0 3
rlabel polysilicon 289 -298 289 -298 0 1
rlabel polysilicon 289 -304 289 -304 0 3
rlabel polysilicon 296 -298 296 -298 0 1
rlabel polysilicon 299 -304 299 -304 0 4
rlabel polysilicon 303 -298 303 -298 0 1
rlabel polysilicon 303 -304 303 -304 0 3
rlabel polysilicon 310 -298 310 -298 0 1
rlabel polysilicon 310 -304 310 -304 0 3
rlabel polysilicon 317 -298 317 -298 0 1
rlabel polysilicon 317 -304 317 -304 0 3
rlabel polysilicon 324 -298 324 -298 0 1
rlabel polysilicon 324 -304 324 -304 0 3
rlabel polysilicon 331 -298 331 -298 0 1
rlabel polysilicon 331 -304 331 -304 0 3
rlabel polysilicon 338 -298 338 -298 0 1
rlabel polysilicon 338 -304 338 -304 0 3
rlabel polysilicon 345 -298 345 -298 0 1
rlabel polysilicon 345 -304 345 -304 0 3
rlabel polysilicon 352 -298 352 -298 0 1
rlabel polysilicon 352 -304 352 -304 0 3
rlabel polysilicon 359 -298 359 -298 0 1
rlabel polysilicon 359 -304 359 -304 0 3
rlabel polysilicon 366 -298 366 -298 0 1
rlabel polysilicon 369 -298 369 -298 0 2
rlabel polysilicon 369 -304 369 -304 0 4
rlabel polysilicon 376 -298 376 -298 0 2
rlabel polysilicon 376 -304 376 -304 0 4
rlabel polysilicon 380 -298 380 -298 0 1
rlabel polysilicon 380 -304 380 -304 0 3
rlabel polysilicon 2 -339 2 -339 0 1
rlabel polysilicon 2 -345 2 -345 0 3
rlabel polysilicon 9 -339 9 -339 0 1
rlabel polysilicon 9 -345 9 -345 0 3
rlabel polysilicon 16 -339 16 -339 0 1
rlabel polysilicon 16 -345 16 -345 0 3
rlabel polysilicon 23 -339 23 -339 0 1
rlabel polysilicon 23 -345 23 -345 0 3
rlabel polysilicon 30 -339 30 -339 0 1
rlabel polysilicon 30 -345 30 -345 0 3
rlabel polysilicon 37 -339 37 -339 0 1
rlabel polysilicon 37 -345 37 -345 0 3
rlabel polysilicon 44 -339 44 -339 0 1
rlabel polysilicon 44 -345 44 -345 0 3
rlabel polysilicon 51 -339 51 -339 0 1
rlabel polysilicon 51 -345 51 -345 0 3
rlabel polysilicon 61 -345 61 -345 0 4
rlabel polysilicon 65 -339 65 -339 0 1
rlabel polysilicon 68 -339 68 -339 0 2
rlabel polysilicon 72 -339 72 -339 0 1
rlabel polysilicon 72 -345 72 -345 0 3
rlabel polysilicon 79 -339 79 -339 0 1
rlabel polysilicon 79 -345 79 -345 0 3
rlabel polysilicon 86 -339 86 -339 0 1
rlabel polysilicon 89 -339 89 -339 0 2
rlabel polysilicon 89 -345 89 -345 0 4
rlabel polysilicon 93 -339 93 -339 0 1
rlabel polysilicon 93 -345 93 -345 0 3
rlabel polysilicon 100 -339 100 -339 0 1
rlabel polysilicon 100 -345 100 -345 0 3
rlabel polysilicon 110 -339 110 -339 0 2
rlabel polysilicon 107 -345 107 -345 0 3
rlabel polysilicon 110 -345 110 -345 0 4
rlabel polysilicon 114 -339 114 -339 0 1
rlabel polysilicon 117 -339 117 -339 0 2
rlabel polysilicon 114 -345 114 -345 0 3
rlabel polysilicon 117 -345 117 -345 0 4
rlabel polysilicon 124 -339 124 -339 0 2
rlabel polysilicon 121 -345 121 -345 0 3
rlabel polysilicon 128 -339 128 -339 0 1
rlabel polysilicon 128 -345 128 -345 0 3
rlabel polysilicon 135 -339 135 -339 0 1
rlabel polysilicon 135 -345 135 -345 0 3
rlabel polysilicon 142 -339 142 -339 0 1
rlabel polysilicon 145 -339 145 -339 0 2
rlabel polysilicon 142 -345 142 -345 0 3
rlabel polysilicon 145 -345 145 -345 0 4
rlabel polysilicon 152 -339 152 -339 0 2
rlabel polysilicon 149 -345 149 -345 0 3
rlabel polysilicon 156 -339 156 -339 0 1
rlabel polysilicon 159 -339 159 -339 0 2
rlabel polysilicon 159 -345 159 -345 0 4
rlabel polysilicon 163 -339 163 -339 0 1
rlabel polysilicon 163 -345 163 -345 0 3
rlabel polysilicon 173 -339 173 -339 0 2
rlabel polysilicon 170 -345 170 -345 0 3
rlabel polysilicon 173 -345 173 -345 0 4
rlabel polysilicon 177 -339 177 -339 0 1
rlabel polysilicon 177 -345 177 -345 0 3
rlabel polysilicon 184 -339 184 -339 0 1
rlabel polysilicon 184 -345 184 -345 0 3
rlabel polysilicon 194 -339 194 -339 0 2
rlabel polysilicon 191 -345 191 -345 0 3
rlabel polysilicon 194 -345 194 -345 0 4
rlabel polysilicon 198 -339 198 -339 0 1
rlabel polysilicon 198 -345 198 -345 0 3
rlabel polysilicon 205 -339 205 -339 0 1
rlabel polysilicon 205 -345 205 -345 0 3
rlabel polysilicon 208 -345 208 -345 0 4
rlabel polysilicon 212 -345 212 -345 0 3
rlabel polysilicon 219 -339 219 -339 0 1
rlabel polysilicon 219 -345 219 -345 0 3
rlabel polysilicon 226 -339 226 -339 0 1
rlabel polysilicon 226 -345 226 -345 0 3
rlabel polysilicon 236 -345 236 -345 0 4
rlabel polysilicon 240 -339 240 -339 0 1
rlabel polysilicon 240 -345 240 -345 0 3
rlabel polysilicon 243 -345 243 -345 0 4
rlabel polysilicon 247 -339 247 -339 0 1
rlabel polysilicon 247 -345 247 -345 0 3
rlabel polysilicon 254 -339 254 -339 0 1
rlabel polysilicon 254 -345 254 -345 0 3
rlabel polysilicon 261 -339 261 -339 0 1
rlabel polysilicon 261 -345 261 -345 0 3
rlabel polysilicon 268 -339 268 -339 0 1
rlabel polysilicon 268 -345 268 -345 0 3
rlabel polysilicon 275 -339 275 -339 0 1
rlabel polysilicon 275 -345 275 -345 0 3
rlabel polysilicon 282 -339 282 -339 0 1
rlabel polysilicon 282 -345 282 -345 0 3
rlabel polysilicon 289 -339 289 -339 0 1
rlabel polysilicon 289 -345 289 -345 0 3
rlabel polysilicon 296 -339 296 -339 0 1
rlabel polysilicon 296 -345 296 -345 0 3
rlabel polysilicon 303 -339 303 -339 0 1
rlabel polysilicon 303 -345 303 -345 0 3
rlabel polysilicon 310 -339 310 -339 0 1
rlabel polysilicon 310 -345 310 -345 0 3
rlabel polysilicon 317 -339 317 -339 0 1
rlabel polysilicon 317 -345 317 -345 0 3
rlabel polysilicon 324 -339 324 -339 0 1
rlabel polysilicon 324 -345 324 -345 0 3
rlabel polysilicon 331 -339 331 -339 0 1
rlabel polysilicon 331 -345 331 -345 0 3
rlabel polysilicon 338 -339 338 -339 0 1
rlabel polysilicon 345 -339 345 -339 0 1
rlabel polysilicon 345 -345 345 -345 0 3
rlabel polysilicon 352 -339 352 -339 0 1
rlabel polysilicon 352 -345 352 -345 0 3
rlabel polysilicon 359 -339 359 -339 0 1
rlabel polysilicon 359 -345 359 -345 0 3
rlabel polysilicon 373 -339 373 -339 0 1
rlabel polysilicon 387 -339 387 -339 0 1
rlabel polysilicon 387 -345 387 -345 0 3
rlabel polysilicon 9 -384 9 -384 0 1
rlabel polysilicon 9 -390 9 -390 0 3
rlabel polysilicon 16 -384 16 -384 0 1
rlabel polysilicon 16 -390 16 -390 0 3
rlabel polysilicon 23 -384 23 -384 0 1
rlabel polysilicon 23 -390 23 -390 0 3
rlabel polysilicon 30 -384 30 -384 0 1
rlabel polysilicon 30 -390 30 -390 0 3
rlabel polysilicon 37 -384 37 -384 0 1
rlabel polysilicon 37 -390 37 -390 0 3
rlabel polysilicon 44 -384 44 -384 0 1
rlabel polysilicon 44 -390 44 -390 0 3
rlabel polysilicon 51 -384 51 -384 0 1
rlabel polysilicon 51 -390 51 -390 0 3
rlabel polysilicon 58 -384 58 -384 0 1
rlabel polysilicon 58 -390 58 -390 0 3
rlabel polysilicon 65 -384 65 -384 0 1
rlabel polysilicon 68 -384 68 -384 0 2
rlabel polysilicon 65 -390 65 -390 0 3
rlabel polysilicon 72 -384 72 -384 0 1
rlabel polysilicon 72 -390 72 -390 0 3
rlabel polysilicon 79 -384 79 -384 0 1
rlabel polysilicon 79 -390 79 -390 0 3
rlabel polysilicon 86 -384 86 -384 0 1
rlabel polysilicon 89 -384 89 -384 0 2
rlabel polysilicon 89 -390 89 -390 0 4
rlabel polysilicon 93 -384 93 -384 0 1
rlabel polysilicon 96 -384 96 -384 0 2
rlabel polysilicon 100 -384 100 -384 0 1
rlabel polysilicon 100 -390 100 -390 0 3
rlabel polysilicon 107 -384 107 -384 0 1
rlabel polysilicon 107 -390 107 -390 0 3
rlabel polysilicon 114 -384 114 -384 0 1
rlabel polysilicon 114 -390 114 -390 0 3
rlabel polysilicon 117 -390 117 -390 0 4
rlabel polysilicon 121 -384 121 -384 0 1
rlabel polysilicon 121 -390 121 -390 0 3
rlabel polysilicon 128 -384 128 -384 0 1
rlabel polysilicon 128 -390 128 -390 0 3
rlabel polysilicon 131 -390 131 -390 0 4
rlabel polysilicon 135 -384 135 -384 0 1
rlabel polysilicon 135 -390 135 -390 0 3
rlabel polysilicon 142 -384 142 -384 0 1
rlabel polysilicon 145 -384 145 -384 0 2
rlabel polysilicon 142 -390 142 -390 0 3
rlabel polysilicon 145 -390 145 -390 0 4
rlabel polysilicon 149 -384 149 -384 0 1
rlabel polysilicon 152 -384 152 -384 0 2
rlabel polysilicon 149 -390 149 -390 0 3
rlabel polysilicon 159 -384 159 -384 0 2
rlabel polysilicon 156 -390 156 -390 0 3
rlabel polysilicon 159 -390 159 -390 0 4
rlabel polysilicon 163 -384 163 -384 0 1
rlabel polysilicon 163 -390 163 -390 0 3
rlabel polysilicon 170 -384 170 -384 0 1
rlabel polysilicon 173 -384 173 -384 0 2
rlabel polysilicon 170 -390 170 -390 0 3
rlabel polysilicon 173 -390 173 -390 0 4
rlabel polysilicon 177 -384 177 -384 0 1
rlabel polysilicon 177 -390 177 -390 0 3
rlabel polysilicon 187 -384 187 -384 0 2
rlabel polysilicon 184 -390 184 -390 0 3
rlabel polysilicon 191 -384 191 -384 0 1
rlabel polysilicon 194 -390 194 -390 0 4
rlabel polysilicon 198 -384 198 -384 0 1
rlabel polysilicon 198 -390 198 -390 0 3
rlabel polysilicon 205 -384 205 -384 0 1
rlabel polysilicon 205 -390 205 -390 0 3
rlabel polysilicon 212 -384 212 -384 0 1
rlabel polysilicon 215 -384 215 -384 0 2
rlabel polysilicon 212 -390 212 -390 0 3
rlabel polysilicon 219 -384 219 -384 0 1
rlabel polysilicon 222 -384 222 -384 0 2
rlabel polysilicon 219 -390 219 -390 0 3
rlabel polysilicon 222 -390 222 -390 0 4
rlabel polysilicon 226 -384 226 -384 0 1
rlabel polysilicon 226 -390 226 -390 0 3
rlabel polysilicon 233 -384 233 -384 0 1
rlabel polysilicon 233 -390 233 -390 0 3
rlabel polysilicon 240 -384 240 -384 0 1
rlabel polysilicon 243 -384 243 -384 0 2
rlabel polysilicon 240 -390 240 -390 0 3
rlabel polysilicon 243 -390 243 -390 0 4
rlabel polysilicon 247 -384 247 -384 0 1
rlabel polysilicon 247 -390 247 -390 0 3
rlabel polysilicon 257 -384 257 -384 0 2
rlabel polysilicon 261 -384 261 -384 0 1
rlabel polysilicon 261 -390 261 -390 0 3
rlabel polysilicon 271 -384 271 -384 0 2
rlabel polysilicon 268 -390 268 -390 0 3
rlabel polysilicon 275 -384 275 -384 0 1
rlabel polysilicon 275 -390 275 -390 0 3
rlabel polysilicon 285 -384 285 -384 0 2
rlabel polysilicon 285 -390 285 -390 0 4
rlabel polysilicon 289 -384 289 -384 0 1
rlabel polysilicon 289 -390 289 -390 0 3
rlabel polysilicon 296 -384 296 -384 0 1
rlabel polysilicon 296 -390 296 -390 0 3
rlabel polysilicon 303 -384 303 -384 0 1
rlabel polysilicon 303 -390 303 -390 0 3
rlabel polysilicon 310 -384 310 -384 0 1
rlabel polysilicon 310 -390 310 -390 0 3
rlabel polysilicon 317 -384 317 -384 0 1
rlabel polysilicon 317 -390 317 -390 0 3
rlabel polysilicon 324 -384 324 -384 0 1
rlabel polysilicon 324 -390 324 -390 0 3
rlabel polysilicon 331 -384 331 -384 0 1
rlabel polysilicon 331 -390 331 -390 0 3
rlabel polysilicon 338 -384 338 -384 0 1
rlabel polysilicon 338 -390 338 -390 0 3
rlabel polysilicon 345 -384 345 -384 0 1
rlabel polysilicon 345 -390 345 -390 0 3
rlabel polysilicon 352 -384 352 -384 0 1
rlabel polysilicon 352 -390 352 -390 0 3
rlabel polysilicon 359 -384 359 -384 0 1
rlabel polysilicon 359 -390 359 -390 0 3
rlabel polysilicon 366 -384 366 -384 0 1
rlabel polysilicon 366 -390 366 -390 0 3
rlabel polysilicon 373 -384 373 -384 0 1
rlabel polysilicon 373 -390 373 -390 0 3
rlabel polysilicon 380 -384 380 -384 0 1
rlabel polysilicon 380 -390 380 -390 0 3
rlabel polysilicon 387 -384 387 -384 0 1
rlabel polysilicon 387 -390 387 -390 0 3
rlabel polysilicon 397 -384 397 -384 0 2
rlabel polysilicon 394 -390 394 -390 0 3
rlabel polysilicon 401 -384 401 -384 0 1
rlabel polysilicon 401 -390 401 -390 0 3
rlabel polysilicon 411 -390 411 -390 0 4
rlabel polysilicon 23 -423 23 -423 0 1
rlabel polysilicon 23 -429 23 -429 0 3
rlabel polysilicon 30 -423 30 -423 0 1
rlabel polysilicon 30 -429 30 -429 0 3
rlabel polysilicon 37 -423 37 -423 0 1
rlabel polysilicon 47 -429 47 -429 0 4
rlabel polysilicon 51 -429 51 -429 0 3
rlabel polysilicon 58 -423 58 -423 0 1
rlabel polysilicon 58 -429 58 -429 0 3
rlabel polysilicon 65 -423 65 -423 0 1
rlabel polysilicon 68 -423 68 -423 0 2
rlabel polysilicon 65 -429 65 -429 0 3
rlabel polysilicon 72 -423 72 -423 0 1
rlabel polysilicon 72 -429 72 -429 0 3
rlabel polysilicon 79 -423 79 -423 0 1
rlabel polysilicon 79 -429 79 -429 0 3
rlabel polysilicon 86 -423 86 -423 0 1
rlabel polysilicon 86 -429 86 -429 0 3
rlabel polysilicon 93 -423 93 -423 0 1
rlabel polysilicon 93 -429 93 -429 0 3
rlabel polysilicon 96 -429 96 -429 0 4
rlabel polysilicon 100 -423 100 -423 0 1
rlabel polysilicon 100 -429 100 -429 0 3
rlabel polysilicon 110 -423 110 -423 0 2
rlabel polysilicon 117 -423 117 -423 0 2
rlabel polysilicon 114 -429 114 -429 0 3
rlabel polysilicon 121 -423 121 -423 0 1
rlabel polysilicon 121 -429 121 -429 0 3
rlabel polysilicon 128 -423 128 -423 0 1
rlabel polysilicon 128 -429 128 -429 0 3
rlabel polysilicon 135 -423 135 -423 0 1
rlabel polysilicon 142 -423 142 -423 0 1
rlabel polysilicon 142 -429 142 -429 0 3
rlabel polysilicon 149 -423 149 -423 0 1
rlabel polysilicon 149 -429 149 -429 0 3
rlabel polysilicon 156 -423 156 -423 0 1
rlabel polysilicon 159 -423 159 -423 0 2
rlabel polysilicon 159 -429 159 -429 0 4
rlabel polysilicon 163 -423 163 -423 0 1
rlabel polysilicon 170 -423 170 -423 0 1
rlabel polysilicon 170 -429 170 -429 0 3
rlabel polysilicon 177 -423 177 -423 0 1
rlabel polysilicon 177 -429 177 -429 0 3
rlabel polysilicon 184 -423 184 -423 0 1
rlabel polysilicon 184 -429 184 -429 0 3
rlabel polysilicon 191 -429 191 -429 0 3
rlabel polysilicon 194 -429 194 -429 0 4
rlabel polysilicon 198 -423 198 -423 0 1
rlabel polysilicon 201 -423 201 -423 0 2
rlabel polysilicon 198 -429 198 -429 0 3
rlabel polysilicon 205 -423 205 -423 0 1
rlabel polysilicon 208 -423 208 -423 0 2
rlabel polysilicon 205 -429 205 -429 0 3
rlabel polysilicon 215 -423 215 -423 0 2
rlabel polysilicon 212 -429 212 -429 0 3
rlabel polysilicon 215 -429 215 -429 0 4
rlabel polysilicon 219 -423 219 -423 0 1
rlabel polysilicon 219 -429 219 -429 0 3
rlabel polysilicon 226 -423 226 -423 0 1
rlabel polysilicon 226 -429 226 -429 0 3
rlabel polysilicon 233 -423 233 -423 0 1
rlabel polysilicon 233 -429 233 -429 0 3
rlabel polysilicon 243 -423 243 -423 0 2
rlabel polysilicon 247 -423 247 -423 0 1
rlabel polysilicon 250 -423 250 -423 0 2
rlabel polysilicon 247 -429 247 -429 0 3
rlabel polysilicon 257 -423 257 -423 0 2
rlabel polysilicon 254 -429 254 -429 0 3
rlabel polysilicon 261 -423 261 -423 0 1
rlabel polysilicon 261 -429 261 -429 0 3
rlabel polysilicon 268 -423 268 -423 0 1
rlabel polysilicon 268 -429 268 -429 0 3
rlabel polysilicon 275 -423 275 -423 0 1
rlabel polysilicon 275 -429 275 -429 0 3
rlabel polysilicon 282 -423 282 -423 0 1
rlabel polysilicon 285 -423 285 -423 0 2
rlabel polysilicon 282 -429 282 -429 0 3
rlabel polysilicon 289 -423 289 -423 0 1
rlabel polysilicon 289 -429 289 -429 0 3
rlabel polysilicon 296 -423 296 -423 0 1
rlabel polysilicon 296 -429 296 -429 0 3
rlabel polysilicon 303 -423 303 -423 0 1
rlabel polysilicon 303 -429 303 -429 0 3
rlabel polysilicon 310 -423 310 -423 0 1
rlabel polysilicon 310 -429 310 -429 0 3
rlabel polysilicon 317 -423 317 -423 0 1
rlabel polysilicon 317 -429 317 -429 0 3
rlabel polysilicon 324 -423 324 -423 0 1
rlabel polysilicon 324 -429 324 -429 0 3
rlabel polysilicon 331 -423 331 -423 0 1
rlabel polysilicon 331 -429 331 -429 0 3
rlabel polysilicon 338 -423 338 -423 0 1
rlabel polysilicon 338 -429 338 -429 0 3
rlabel polysilicon 345 -423 345 -423 0 1
rlabel polysilicon 345 -429 345 -429 0 3
rlabel polysilicon 352 -423 352 -423 0 1
rlabel polysilicon 352 -429 352 -429 0 3
rlabel polysilicon 355 -429 355 -429 0 4
rlabel polysilicon 359 -423 359 -423 0 1
rlabel polysilicon 362 -429 362 -429 0 4
rlabel polysilicon 366 -423 366 -423 0 1
rlabel polysilicon 366 -429 366 -429 0 3
rlabel polysilicon 373 -423 373 -423 0 1
rlabel polysilicon 373 -429 373 -429 0 3
rlabel polysilicon 380 -423 380 -423 0 1
rlabel polysilicon 380 -429 380 -429 0 3
rlabel polysilicon 26 -462 26 -462 0 4
rlabel polysilicon 33 -462 33 -462 0 4
rlabel polysilicon 37 -456 37 -456 0 1
rlabel polysilicon 37 -462 37 -462 0 3
rlabel polysilicon 44 -456 44 -456 0 1
rlabel polysilicon 44 -462 44 -462 0 3
rlabel polysilicon 51 -456 51 -456 0 1
rlabel polysilicon 51 -462 51 -462 0 3
rlabel polysilicon 58 -456 58 -456 0 1
rlabel polysilicon 58 -462 58 -462 0 3
rlabel polysilicon 65 -456 65 -456 0 1
rlabel polysilicon 68 -456 68 -456 0 2
rlabel polysilicon 75 -456 75 -456 0 2
rlabel polysilicon 72 -462 72 -462 0 3
rlabel polysilicon 79 -456 79 -456 0 1
rlabel polysilicon 79 -462 79 -462 0 3
rlabel polysilicon 86 -456 86 -456 0 1
rlabel polysilicon 86 -462 86 -462 0 3
rlabel polysilicon 93 -456 93 -456 0 1
rlabel polysilicon 93 -462 93 -462 0 3
rlabel polysilicon 100 -456 100 -456 0 1
rlabel polysilicon 100 -462 100 -462 0 3
rlabel polysilicon 107 -456 107 -456 0 1
rlabel polysilicon 107 -462 107 -462 0 3
rlabel polysilicon 114 -456 114 -456 0 1
rlabel polysilicon 117 -456 117 -456 0 2
rlabel polysilicon 114 -462 114 -462 0 3
rlabel polysilicon 117 -462 117 -462 0 4
rlabel polysilicon 124 -456 124 -456 0 2
rlabel polysilicon 121 -462 121 -462 0 3
rlabel polysilicon 131 -456 131 -456 0 2
rlabel polysilicon 128 -462 128 -462 0 3
rlabel polysilicon 131 -462 131 -462 0 4
rlabel polysilicon 135 -456 135 -456 0 1
rlabel polysilicon 135 -462 135 -462 0 3
rlabel polysilicon 138 -462 138 -462 0 4
rlabel polysilicon 142 -456 142 -456 0 1
rlabel polysilicon 145 -462 145 -462 0 4
rlabel polysilicon 149 -456 149 -456 0 1
rlabel polysilicon 149 -462 149 -462 0 3
rlabel polysilicon 156 -456 156 -456 0 1
rlabel polysilicon 159 -456 159 -456 0 2
rlabel polysilicon 163 -456 163 -456 0 1
rlabel polysilicon 163 -462 163 -462 0 3
rlabel polysilicon 170 -456 170 -456 0 1
rlabel polysilicon 170 -462 170 -462 0 3
rlabel polysilicon 177 -456 177 -456 0 1
rlabel polysilicon 177 -462 177 -462 0 3
rlabel polysilicon 184 -456 184 -456 0 1
rlabel polysilicon 187 -456 187 -456 0 2
rlabel polysilicon 187 -462 187 -462 0 4
rlabel polysilicon 191 -456 191 -456 0 1
rlabel polysilicon 194 -456 194 -456 0 2
rlabel polysilicon 191 -462 191 -462 0 3
rlabel polysilicon 194 -462 194 -462 0 4
rlabel polysilicon 198 -456 198 -456 0 1
rlabel polysilicon 198 -462 198 -462 0 3
rlabel polysilicon 205 -456 205 -456 0 1
rlabel polysilicon 205 -462 205 -462 0 3
rlabel polysilicon 212 -456 212 -456 0 1
rlabel polysilicon 215 -456 215 -456 0 2
rlabel polysilicon 212 -462 212 -462 0 3
rlabel polysilicon 219 -456 219 -456 0 1
rlabel polysilicon 219 -462 219 -462 0 3
rlabel polysilicon 229 -456 229 -456 0 2
rlabel polysilicon 226 -462 226 -462 0 3
rlabel polysilicon 229 -462 229 -462 0 4
rlabel polysilicon 233 -456 233 -456 0 1
rlabel polysilicon 233 -462 233 -462 0 3
rlabel polysilicon 240 -456 240 -456 0 1
rlabel polysilicon 240 -462 240 -462 0 3
rlabel polysilicon 250 -462 250 -462 0 4
rlabel polysilicon 254 -456 254 -456 0 1
rlabel polysilicon 254 -462 254 -462 0 3
rlabel polysilicon 261 -456 261 -456 0 1
rlabel polysilicon 261 -462 261 -462 0 3
rlabel polysilicon 268 -456 268 -456 0 1
rlabel polysilicon 268 -462 268 -462 0 3
rlabel polysilicon 275 -456 275 -456 0 1
rlabel polysilicon 275 -462 275 -462 0 3
rlabel polysilicon 282 -456 282 -456 0 1
rlabel polysilicon 282 -462 282 -462 0 3
rlabel polysilicon 289 -456 289 -456 0 1
rlabel polysilicon 289 -462 289 -462 0 3
rlabel polysilicon 296 -456 296 -456 0 1
rlabel polysilicon 296 -462 296 -462 0 3
rlabel polysilicon 303 -456 303 -456 0 1
rlabel polysilicon 306 -456 306 -456 0 2
rlabel polysilicon 306 -462 306 -462 0 4
rlabel polysilicon 313 -456 313 -456 0 2
rlabel polysilicon 320 -456 320 -456 0 2
rlabel polysilicon 317 -462 317 -462 0 3
rlabel polysilicon 331 -456 331 -456 0 1
rlabel polysilicon 331 -462 331 -462 0 3
rlabel polysilicon 352 -456 352 -456 0 1
rlabel polysilicon 352 -462 352 -462 0 3
rlabel polysilicon 359 -456 359 -456 0 1
rlabel polysilicon 359 -462 359 -462 0 3
rlabel polysilicon 366 -456 366 -456 0 1
rlabel polysilicon 366 -462 366 -462 0 3
rlabel polysilicon 376 -462 376 -462 0 4
rlabel polysilicon 37 -493 37 -493 0 1
rlabel polysilicon 37 -499 37 -499 0 3
rlabel polysilicon 44 -493 44 -493 0 1
rlabel polysilicon 44 -499 44 -499 0 3
rlabel polysilicon 51 -493 51 -493 0 1
rlabel polysilicon 51 -499 51 -499 0 3
rlabel polysilicon 58 -493 58 -493 0 1
rlabel polysilicon 58 -499 58 -499 0 3
rlabel polysilicon 65 -493 65 -493 0 1
rlabel polysilicon 68 -493 68 -493 0 2
rlabel polysilicon 65 -499 65 -499 0 3
rlabel polysilicon 68 -499 68 -499 0 4
rlabel polysilicon 72 -493 72 -493 0 1
rlabel polysilicon 72 -499 72 -499 0 3
rlabel polysilicon 79 -493 79 -493 0 1
rlabel polysilicon 79 -499 79 -499 0 3
rlabel polysilicon 86 -493 86 -493 0 1
rlabel polysilicon 86 -499 86 -499 0 3
rlabel polysilicon 93 -499 93 -499 0 3
rlabel polysilicon 100 -493 100 -493 0 1
rlabel polysilicon 100 -499 100 -499 0 3
rlabel polysilicon 110 -493 110 -493 0 2
rlabel polysilicon 107 -499 107 -499 0 3
rlabel polysilicon 110 -499 110 -499 0 4
rlabel polysilicon 114 -493 114 -493 0 1
rlabel polysilicon 114 -499 114 -499 0 3
rlabel polysilicon 121 -493 121 -493 0 1
rlabel polysilicon 121 -499 121 -499 0 3
rlabel polysilicon 128 -493 128 -493 0 1
rlabel polysilicon 131 -493 131 -493 0 2
rlabel polysilicon 135 -493 135 -493 0 1
rlabel polysilicon 135 -499 135 -499 0 3
rlabel polysilicon 142 -493 142 -493 0 1
rlabel polysilicon 142 -499 142 -499 0 3
rlabel polysilicon 149 -493 149 -493 0 1
rlabel polysilicon 149 -499 149 -499 0 3
rlabel polysilicon 156 -493 156 -493 0 1
rlabel polysilicon 156 -499 156 -499 0 3
rlabel polysilicon 163 -493 163 -493 0 1
rlabel polysilicon 163 -499 163 -499 0 3
rlabel polysilicon 170 -493 170 -493 0 1
rlabel polysilicon 173 -493 173 -493 0 2
rlabel polysilicon 173 -499 173 -499 0 4
rlabel polysilicon 177 -493 177 -493 0 1
rlabel polysilicon 177 -499 177 -499 0 3
rlabel polysilicon 184 -493 184 -493 0 1
rlabel polysilicon 184 -499 184 -499 0 3
rlabel polysilicon 194 -499 194 -499 0 4
rlabel polysilicon 198 -493 198 -493 0 1
rlabel polysilicon 198 -499 198 -499 0 3
rlabel polysilicon 201 -499 201 -499 0 4
rlabel polysilicon 205 -493 205 -493 0 1
rlabel polysilicon 208 -493 208 -493 0 2
rlabel polysilicon 215 -493 215 -493 0 2
rlabel polysilicon 212 -499 212 -499 0 3
rlabel polysilicon 219 -499 219 -499 0 3
rlabel polysilicon 226 -493 226 -493 0 1
rlabel polysilicon 226 -499 226 -499 0 3
rlabel polysilicon 233 -493 233 -493 0 1
rlabel polysilicon 233 -499 233 -499 0 3
rlabel polysilicon 240 -493 240 -493 0 1
rlabel polysilicon 243 -493 243 -493 0 2
rlabel polysilicon 240 -499 240 -499 0 3
rlabel polysilicon 243 -499 243 -499 0 4
rlabel polysilicon 247 -493 247 -493 0 1
rlabel polysilicon 247 -499 247 -499 0 3
rlabel polysilicon 254 -493 254 -493 0 1
rlabel polysilicon 254 -499 254 -499 0 3
rlabel polysilicon 261 -493 261 -493 0 1
rlabel polysilicon 261 -499 261 -499 0 3
rlabel polysilicon 268 -493 268 -493 0 1
rlabel polysilicon 268 -499 268 -499 0 3
rlabel polysilicon 275 -493 275 -493 0 1
rlabel polysilicon 275 -499 275 -499 0 3
rlabel polysilicon 282 -499 282 -499 0 3
rlabel polysilicon 289 -493 289 -493 0 1
rlabel polysilicon 289 -499 289 -499 0 3
rlabel polysilicon 296 -499 296 -499 0 3
rlabel polysilicon 299 -499 299 -499 0 4
rlabel polysilicon 303 -493 303 -493 0 1
rlabel polysilicon 303 -499 303 -499 0 3
rlabel polysilicon 313 -499 313 -499 0 4
rlabel polysilicon 320 -493 320 -493 0 2
rlabel polysilicon 324 -493 324 -493 0 1
rlabel polysilicon 324 -499 324 -499 0 3
rlabel polysilicon 331 -493 331 -493 0 1
rlabel polysilicon 331 -499 331 -499 0 3
rlabel polysilicon 338 -493 338 -493 0 1
rlabel polysilicon 341 -499 341 -499 0 4
rlabel polysilicon 348 -493 348 -493 0 2
rlabel polysilicon 348 -499 348 -499 0 4
rlabel polysilicon 352 -493 352 -493 0 1
rlabel polysilicon 352 -499 352 -499 0 3
rlabel polysilicon 359 -493 359 -493 0 1
rlabel polysilicon 16 -532 16 -532 0 1
rlabel polysilicon 16 -538 16 -538 0 3
rlabel polysilicon 26 -538 26 -538 0 4
rlabel polysilicon 30 -532 30 -532 0 1
rlabel polysilicon 30 -538 30 -538 0 3
rlabel polysilicon 37 -532 37 -532 0 1
rlabel polysilicon 37 -538 37 -538 0 3
rlabel polysilicon 44 -532 44 -532 0 1
rlabel polysilicon 44 -538 44 -538 0 3
rlabel polysilicon 51 -532 51 -532 0 1
rlabel polysilicon 51 -538 51 -538 0 3
rlabel polysilicon 58 -532 58 -532 0 1
rlabel polysilicon 58 -538 58 -538 0 3
rlabel polysilicon 65 -532 65 -532 0 1
rlabel polysilicon 65 -538 65 -538 0 3
rlabel polysilicon 72 -532 72 -532 0 1
rlabel polysilicon 79 -532 79 -532 0 1
rlabel polysilicon 79 -538 79 -538 0 3
rlabel polysilicon 86 -532 86 -532 0 1
rlabel polysilicon 86 -538 86 -538 0 3
rlabel polysilicon 93 -532 93 -532 0 1
rlabel polysilicon 93 -538 93 -538 0 3
rlabel polysilicon 100 -532 100 -532 0 1
rlabel polysilicon 100 -538 100 -538 0 3
rlabel polysilicon 103 -538 103 -538 0 4
rlabel polysilicon 110 -532 110 -532 0 2
rlabel polysilicon 110 -538 110 -538 0 4
rlabel polysilicon 114 -532 114 -532 0 1
rlabel polysilicon 114 -538 114 -538 0 3
rlabel polysilicon 124 -538 124 -538 0 4
rlabel polysilicon 131 -532 131 -532 0 2
rlabel polysilicon 128 -538 128 -538 0 3
rlabel polysilicon 131 -538 131 -538 0 4
rlabel polysilicon 135 -532 135 -532 0 1
rlabel polysilicon 135 -538 135 -538 0 3
rlabel polysilicon 142 -532 142 -532 0 1
rlabel polysilicon 145 -538 145 -538 0 4
rlabel polysilicon 149 -532 149 -532 0 1
rlabel polysilicon 149 -538 149 -538 0 3
rlabel polysilicon 152 -538 152 -538 0 4
rlabel polysilicon 156 -532 156 -532 0 1
rlabel polysilicon 159 -532 159 -532 0 2
rlabel polysilicon 156 -538 156 -538 0 3
rlabel polysilicon 163 -532 163 -532 0 1
rlabel polysilicon 166 -532 166 -532 0 2
rlabel polysilicon 166 -538 166 -538 0 4
rlabel polysilicon 170 -532 170 -532 0 1
rlabel polysilicon 170 -538 170 -538 0 3
rlabel polysilicon 177 -532 177 -532 0 1
rlabel polysilicon 177 -538 177 -538 0 3
rlabel polysilicon 184 -532 184 -532 0 1
rlabel polysilicon 191 -532 191 -532 0 1
rlabel polysilicon 194 -532 194 -532 0 2
rlabel polysilicon 198 -532 198 -532 0 1
rlabel polysilicon 201 -532 201 -532 0 2
rlabel polysilicon 198 -538 198 -538 0 3
rlabel polysilicon 201 -538 201 -538 0 4
rlabel polysilicon 205 -532 205 -532 0 1
rlabel polysilicon 208 -532 208 -532 0 2
rlabel polysilicon 205 -538 205 -538 0 3
rlabel polysilicon 208 -538 208 -538 0 4
rlabel polysilicon 212 -532 212 -532 0 1
rlabel polysilicon 212 -538 212 -538 0 3
rlabel polysilicon 219 -532 219 -532 0 1
rlabel polysilicon 222 -532 222 -532 0 2
rlabel polysilicon 222 -538 222 -538 0 4
rlabel polysilicon 226 -532 226 -532 0 1
rlabel polysilicon 229 -532 229 -532 0 2
rlabel polysilicon 229 -538 229 -538 0 4
rlabel polysilicon 233 -532 233 -532 0 1
rlabel polysilicon 233 -538 233 -538 0 3
rlabel polysilicon 240 -532 240 -532 0 1
rlabel polysilicon 240 -538 240 -538 0 3
rlabel polysilicon 247 -532 247 -532 0 1
rlabel polysilicon 247 -538 247 -538 0 3
rlabel polysilicon 254 -532 254 -532 0 1
rlabel polysilicon 254 -538 254 -538 0 3
rlabel polysilicon 261 -532 261 -532 0 1
rlabel polysilicon 261 -538 261 -538 0 3
rlabel polysilicon 268 -532 268 -532 0 1
rlabel polysilicon 268 -538 268 -538 0 3
rlabel polysilicon 275 -538 275 -538 0 3
rlabel polysilicon 278 -538 278 -538 0 4
rlabel polysilicon 282 -532 282 -532 0 1
rlabel polysilicon 282 -538 282 -538 0 3
rlabel polysilicon 289 -532 289 -532 0 1
rlabel polysilicon 289 -538 289 -538 0 3
rlabel polysilicon 296 -532 296 -532 0 1
rlabel polysilicon 296 -538 296 -538 0 3
rlabel polysilicon 303 -532 303 -532 0 1
rlabel polysilicon 303 -538 303 -538 0 3
rlabel polysilicon 310 -532 310 -532 0 1
rlabel polysilicon 310 -538 310 -538 0 3
rlabel polysilicon 317 -532 317 -532 0 1
rlabel polysilicon 317 -538 317 -538 0 3
rlabel polysilicon 324 -532 324 -532 0 1
rlabel polysilicon 324 -538 324 -538 0 3
rlabel polysilicon 331 -532 331 -532 0 1
rlabel polysilicon 331 -538 331 -538 0 3
rlabel polysilicon 338 -532 338 -532 0 1
rlabel polysilicon 341 -532 341 -532 0 2
rlabel polysilicon 338 -538 338 -538 0 3
rlabel polysilicon 345 -532 345 -532 0 1
rlabel polysilicon 348 -532 348 -532 0 2
rlabel polysilicon 345 -538 345 -538 0 3
rlabel polysilicon 348 -538 348 -538 0 4
rlabel polysilicon 352 -532 352 -532 0 1
rlabel polysilicon 352 -538 352 -538 0 3
rlabel polysilicon 359 -532 359 -532 0 1
rlabel polysilicon 359 -538 359 -538 0 3
rlabel polysilicon 366 -532 366 -532 0 1
rlabel polysilicon 366 -538 366 -538 0 3
rlabel polysilicon 373 -532 373 -532 0 1
rlabel polysilicon 373 -538 373 -538 0 3
rlabel polysilicon 9 -571 9 -571 0 1
rlabel polysilicon 9 -577 9 -577 0 3
rlabel polysilicon 16 -571 16 -571 0 1
rlabel polysilicon 16 -577 16 -577 0 3
rlabel polysilicon 23 -571 23 -571 0 1
rlabel polysilicon 23 -577 23 -577 0 3
rlabel polysilicon 33 -577 33 -577 0 4
rlabel polysilicon 40 -577 40 -577 0 4
rlabel polysilicon 44 -571 44 -571 0 1
rlabel polysilicon 44 -577 44 -577 0 3
rlabel polysilicon 51 -577 51 -577 0 3
rlabel polysilicon 58 -571 58 -571 0 1
rlabel polysilicon 58 -577 58 -577 0 3
rlabel polysilicon 65 -571 65 -571 0 1
rlabel polysilicon 65 -577 65 -577 0 3
rlabel polysilicon 72 -571 72 -571 0 1
rlabel polysilicon 72 -577 72 -577 0 3
rlabel polysilicon 82 -571 82 -571 0 2
rlabel polysilicon 79 -577 79 -577 0 3
rlabel polysilicon 82 -577 82 -577 0 4
rlabel polysilicon 86 -571 86 -571 0 1
rlabel polysilicon 86 -577 86 -577 0 3
rlabel polysilicon 93 -571 93 -571 0 1
rlabel polysilicon 93 -577 93 -577 0 3
rlabel polysilicon 100 -571 100 -571 0 1
rlabel polysilicon 100 -577 100 -577 0 3
rlabel polysilicon 107 -571 107 -571 0 1
rlabel polysilicon 107 -577 107 -577 0 3
rlabel polysilicon 110 -577 110 -577 0 4
rlabel polysilicon 114 -571 114 -571 0 1
rlabel polysilicon 114 -577 114 -577 0 3
rlabel polysilicon 121 -571 121 -571 0 1
rlabel polysilicon 124 -571 124 -571 0 2
rlabel polysilicon 131 -571 131 -571 0 2
rlabel polysilicon 131 -577 131 -577 0 4
rlabel polysilicon 135 -571 135 -571 0 1
rlabel polysilicon 135 -577 135 -577 0 3
rlabel polysilicon 142 -571 142 -571 0 1
rlabel polysilicon 145 -571 145 -571 0 2
rlabel polysilicon 145 -577 145 -577 0 4
rlabel polysilicon 152 -571 152 -571 0 2
rlabel polysilicon 152 -577 152 -577 0 4
rlabel polysilicon 159 -571 159 -571 0 2
rlabel polysilicon 159 -577 159 -577 0 4
rlabel polysilicon 163 -571 163 -571 0 1
rlabel polysilicon 163 -577 163 -577 0 3
rlabel polysilicon 170 -571 170 -571 0 1
rlabel polysilicon 177 -571 177 -571 0 1
rlabel polysilicon 177 -577 177 -577 0 3
rlabel polysilicon 187 -577 187 -577 0 4
rlabel polysilicon 191 -571 191 -571 0 1
rlabel polysilicon 191 -577 191 -577 0 3
rlabel polysilicon 198 -571 198 -571 0 1
rlabel polysilicon 198 -577 198 -577 0 3
rlabel polysilicon 205 -571 205 -571 0 1
rlabel polysilicon 205 -577 205 -577 0 3
rlabel polysilicon 212 -571 212 -571 0 1
rlabel polysilicon 212 -577 212 -577 0 3
rlabel polysilicon 219 -571 219 -571 0 1
rlabel polysilicon 219 -577 219 -577 0 3
rlabel polysilicon 226 -571 226 -571 0 1
rlabel polysilicon 226 -577 226 -577 0 3
rlabel polysilicon 236 -571 236 -571 0 2
rlabel polysilicon 240 -571 240 -571 0 1
rlabel polysilicon 240 -577 240 -577 0 3
rlabel polysilicon 247 -571 247 -571 0 1
rlabel polysilicon 247 -577 247 -577 0 3
rlabel polysilicon 257 -577 257 -577 0 4
rlabel polysilicon 261 -571 261 -571 0 1
rlabel polysilicon 261 -577 261 -577 0 3
rlabel polysilicon 268 -571 268 -571 0 1
rlabel polysilicon 268 -577 268 -577 0 3
rlabel polysilicon 275 -571 275 -571 0 1
rlabel polysilicon 278 -571 278 -571 0 2
rlabel polysilicon 282 -571 282 -571 0 1
rlabel polysilicon 282 -577 282 -577 0 3
rlabel polysilicon 289 -571 289 -571 0 1
rlabel polysilicon 292 -571 292 -571 0 2
rlabel polysilicon 296 -571 296 -571 0 1
rlabel polysilicon 296 -577 296 -577 0 3
rlabel polysilicon 303 -571 303 -571 0 1
rlabel polysilicon 303 -577 303 -577 0 3
rlabel polysilicon 310 -577 310 -577 0 3
rlabel polysilicon 324 -571 324 -571 0 1
rlabel polysilicon 324 -577 324 -577 0 3
rlabel polysilicon 355 -577 355 -577 0 4
rlabel polysilicon 359 -571 359 -571 0 1
rlabel polysilicon 359 -577 359 -577 0 3
rlabel polysilicon 23 -602 23 -602 0 1
rlabel polysilicon 26 -608 26 -608 0 4
rlabel polysilicon 30 -602 30 -602 0 1
rlabel polysilicon 30 -608 30 -608 0 3
rlabel polysilicon 40 -602 40 -602 0 2
rlabel polysilicon 37 -608 37 -608 0 3
rlabel polysilicon 44 -602 44 -602 0 1
rlabel polysilicon 44 -608 44 -608 0 3
rlabel polysilicon 51 -602 51 -602 0 1
rlabel polysilicon 51 -608 51 -608 0 3
rlabel polysilicon 58 -602 58 -602 0 1
rlabel polysilicon 58 -608 58 -608 0 3
rlabel polysilicon 65 -602 65 -602 0 1
rlabel polysilicon 65 -608 65 -608 0 3
rlabel polysilicon 75 -602 75 -602 0 2
rlabel polysilicon 75 -608 75 -608 0 4
rlabel polysilicon 79 -602 79 -602 0 1
rlabel polysilicon 79 -608 79 -608 0 3
rlabel polysilicon 82 -608 82 -608 0 4
rlabel polysilicon 86 -602 86 -602 0 1
rlabel polysilicon 86 -608 86 -608 0 3
rlabel polysilicon 93 -602 93 -602 0 1
rlabel polysilicon 96 -602 96 -602 0 2
rlabel polysilicon 100 -602 100 -602 0 1
rlabel polysilicon 100 -608 100 -608 0 3
rlabel polysilicon 107 -602 107 -602 0 1
rlabel polysilicon 107 -608 107 -608 0 3
rlabel polysilicon 114 -602 114 -602 0 1
rlabel polysilicon 114 -608 114 -608 0 3
rlabel polysilicon 117 -608 117 -608 0 4
rlabel polysilicon 121 -602 121 -602 0 1
rlabel polysilicon 121 -608 121 -608 0 3
rlabel polysilicon 128 -602 128 -602 0 1
rlabel polysilicon 131 -608 131 -608 0 4
rlabel polysilicon 135 -602 135 -602 0 1
rlabel polysilicon 138 -602 138 -602 0 2
rlabel polysilicon 135 -608 135 -608 0 3
rlabel polysilicon 138 -608 138 -608 0 4
rlabel polysilicon 142 -602 142 -602 0 1
rlabel polysilicon 142 -608 142 -608 0 3
rlabel polysilicon 149 -602 149 -602 0 1
rlabel polysilicon 152 -602 152 -602 0 2
rlabel polysilicon 149 -608 149 -608 0 3
rlabel polysilicon 152 -608 152 -608 0 4
rlabel polysilicon 156 -602 156 -602 0 1
rlabel polysilicon 159 -602 159 -602 0 2
rlabel polysilicon 156 -608 156 -608 0 3
rlabel polysilicon 159 -608 159 -608 0 4
rlabel polysilicon 163 -602 163 -602 0 1
rlabel polysilicon 163 -608 163 -608 0 3
rlabel polysilicon 170 -602 170 -602 0 1
rlabel polysilicon 170 -608 170 -608 0 3
rlabel polysilicon 177 -602 177 -602 0 1
rlabel polysilicon 177 -608 177 -608 0 3
rlabel polysilicon 180 -608 180 -608 0 4
rlabel polysilicon 184 -602 184 -602 0 1
rlabel polysilicon 187 -602 187 -602 0 2
rlabel polysilicon 191 -602 191 -602 0 1
rlabel polysilicon 191 -608 191 -608 0 3
rlabel polysilicon 198 -602 198 -602 0 1
rlabel polysilicon 198 -608 198 -608 0 3
rlabel polysilicon 205 -602 205 -602 0 1
rlabel polysilicon 205 -608 205 -608 0 3
rlabel polysilicon 212 -602 212 -602 0 1
rlabel polysilicon 212 -608 212 -608 0 3
rlabel polysilicon 219 -602 219 -602 0 1
rlabel polysilicon 219 -608 219 -608 0 3
rlabel polysilicon 229 -602 229 -602 0 2
rlabel polysilicon 226 -608 226 -608 0 3
rlabel polysilicon 233 -602 233 -602 0 1
rlabel polysilicon 233 -608 233 -608 0 3
rlabel polysilicon 243 -608 243 -608 0 4
rlabel polysilicon 247 -602 247 -602 0 1
rlabel polysilicon 247 -608 247 -608 0 3
rlabel polysilicon 254 -602 254 -602 0 1
rlabel polysilicon 254 -608 254 -608 0 3
rlabel polysilicon 261 -602 261 -602 0 1
rlabel polysilicon 261 -608 261 -608 0 3
rlabel polysilicon 268 -602 268 -602 0 1
rlabel polysilicon 268 -608 268 -608 0 3
rlabel polysilicon 278 -602 278 -602 0 2
rlabel polysilicon 275 -608 275 -608 0 3
rlabel polysilicon 282 -602 282 -602 0 1
rlabel polysilicon 282 -608 282 -608 0 3
rlabel polysilicon 289 -602 289 -602 0 1
rlabel polysilicon 289 -608 289 -608 0 3
rlabel polysilicon 303 -602 303 -602 0 1
rlabel polysilicon 306 -602 306 -602 0 2
rlabel polysilicon 324 -602 324 -602 0 1
rlabel polysilicon 324 -608 324 -608 0 3
rlabel polysilicon 26 -627 26 -627 0 2
rlabel polysilicon 51 -627 51 -627 0 1
rlabel polysilicon 51 -633 51 -633 0 3
rlabel polysilicon 65 -627 65 -627 0 1
rlabel polysilicon 65 -633 65 -633 0 3
rlabel polysilicon 72 -627 72 -627 0 1
rlabel polysilicon 75 -633 75 -633 0 4
rlabel polysilicon 79 -627 79 -627 0 1
rlabel polysilicon 82 -633 82 -633 0 4
rlabel polysilicon 86 -627 86 -627 0 1
rlabel polysilicon 93 -627 93 -627 0 1
rlabel polysilicon 93 -633 93 -633 0 3
rlabel polysilicon 103 -627 103 -627 0 2
rlabel polysilicon 100 -633 100 -633 0 3
rlabel polysilicon 107 -627 107 -627 0 1
rlabel polysilicon 107 -633 107 -633 0 3
rlabel polysilicon 114 -627 114 -627 0 1
rlabel polysilicon 117 -627 117 -627 0 2
rlabel polysilicon 121 -627 121 -627 0 1
rlabel polysilicon 121 -633 121 -633 0 3
rlabel polysilicon 128 -627 128 -627 0 1
rlabel polysilicon 128 -633 128 -633 0 3
rlabel polysilicon 135 -627 135 -627 0 1
rlabel polysilicon 135 -633 135 -633 0 3
rlabel polysilicon 142 -627 142 -627 0 1
rlabel polysilicon 145 -627 145 -627 0 2
rlabel polysilicon 145 -633 145 -633 0 4
rlabel polysilicon 149 -633 149 -633 0 3
rlabel polysilicon 152 -633 152 -633 0 4
rlabel polysilicon 156 -627 156 -627 0 1
rlabel polysilicon 156 -633 156 -633 0 3
rlabel polysilicon 163 -627 163 -627 0 1
rlabel polysilicon 163 -633 163 -633 0 3
rlabel polysilicon 173 -627 173 -627 0 2
rlabel polysilicon 180 -627 180 -627 0 2
rlabel polysilicon 184 -627 184 -627 0 1
rlabel polysilicon 187 -627 187 -627 0 2
rlabel polysilicon 187 -633 187 -633 0 4
rlabel polysilicon 191 -627 191 -627 0 1
rlabel polysilicon 191 -633 191 -633 0 3
rlabel polysilicon 198 -627 198 -627 0 1
rlabel polysilicon 198 -633 198 -633 0 3
rlabel polysilicon 205 -627 205 -627 0 1
rlabel polysilicon 205 -633 205 -633 0 3
rlabel polysilicon 212 -627 212 -627 0 1
rlabel polysilicon 212 -633 212 -633 0 3
rlabel polysilicon 219 -627 219 -627 0 1
rlabel polysilicon 219 -633 219 -633 0 3
rlabel polysilicon 226 -627 226 -627 0 1
rlabel polysilicon 226 -633 226 -633 0 3
rlabel polysilicon 233 -627 233 -627 0 1
rlabel polysilicon 233 -633 233 -633 0 3
rlabel polysilicon 236 -633 236 -633 0 4
rlabel polysilicon 240 -627 240 -627 0 1
rlabel polysilicon 240 -633 240 -633 0 3
rlabel polysilicon 247 -627 247 -627 0 1
rlabel polysilicon 247 -633 247 -633 0 3
rlabel polysilicon 254 -627 254 -627 0 1
rlabel polysilicon 257 -627 257 -627 0 2
rlabel polysilicon 257 -633 257 -633 0 4
rlabel polysilicon 261 -627 261 -627 0 1
rlabel polysilicon 264 -627 264 -627 0 2
rlabel polysilicon 324 -627 324 -627 0 1
rlabel polysilicon 30 -660 30 -660 0 1
rlabel polysilicon 30 -666 30 -666 0 3
rlabel polysilicon 37 -660 37 -660 0 1
rlabel polysilicon 37 -666 37 -666 0 3
rlabel polysilicon 44 -660 44 -660 0 1
rlabel polysilicon 44 -666 44 -666 0 3
rlabel polysilicon 51 -660 51 -660 0 1
rlabel polysilicon 51 -666 51 -666 0 3
rlabel polysilicon 58 -666 58 -666 0 3
rlabel polysilicon 61 -666 61 -666 0 4
rlabel polysilicon 68 -660 68 -660 0 2
rlabel polysilicon 68 -666 68 -666 0 4
rlabel polysilicon 72 -660 72 -660 0 1
rlabel polysilicon 75 -660 75 -660 0 2
rlabel polysilicon 79 -660 79 -660 0 1
rlabel polysilicon 79 -666 79 -666 0 3
rlabel polysilicon 86 -660 86 -660 0 1
rlabel polysilicon 86 -666 86 -666 0 3
rlabel polysilicon 96 -660 96 -660 0 2
rlabel polysilicon 93 -666 93 -666 0 3
rlabel polysilicon 96 -666 96 -666 0 4
rlabel polysilicon 100 -660 100 -660 0 1
rlabel polysilicon 100 -666 100 -666 0 3
rlabel polysilicon 107 -660 107 -660 0 1
rlabel polysilicon 107 -666 107 -666 0 3
rlabel polysilicon 117 -660 117 -660 0 2
rlabel polysilicon 114 -666 114 -666 0 3
rlabel polysilicon 117 -666 117 -666 0 4
rlabel polysilicon 121 -660 121 -660 0 1
rlabel polysilicon 124 -660 124 -660 0 2
rlabel polysilicon 128 -660 128 -660 0 1
rlabel polysilicon 128 -666 128 -666 0 3
rlabel polysilicon 135 -660 135 -660 0 1
rlabel polysilicon 138 -660 138 -660 0 2
rlabel polysilicon 138 -666 138 -666 0 4
rlabel polysilicon 142 -660 142 -660 0 1
rlabel polysilicon 145 -666 145 -666 0 4
rlabel polysilicon 149 -660 149 -660 0 1
rlabel polysilicon 149 -666 149 -666 0 3
rlabel polysilicon 156 -660 156 -660 0 1
rlabel polysilicon 156 -666 156 -666 0 3
rlabel polysilicon 159 -666 159 -666 0 4
rlabel polysilicon 163 -660 163 -660 0 1
rlabel polysilicon 163 -666 163 -666 0 3
rlabel polysilicon 170 -660 170 -660 0 1
rlabel polysilicon 173 -660 173 -660 0 2
rlabel polysilicon 173 -666 173 -666 0 4
rlabel polysilicon 177 -666 177 -666 0 3
rlabel polysilicon 180 -666 180 -666 0 4
rlabel polysilicon 184 -660 184 -660 0 1
rlabel polysilicon 187 -660 187 -660 0 2
rlabel polysilicon 184 -666 184 -666 0 3
rlabel polysilicon 191 -660 191 -660 0 1
rlabel polysilicon 191 -666 191 -666 0 3
rlabel polysilicon 201 -660 201 -660 0 2
rlabel polysilicon 201 -666 201 -666 0 4
rlabel polysilicon 205 -666 205 -666 0 3
rlabel polysilicon 208 -666 208 -666 0 4
rlabel polysilicon 212 -660 212 -660 0 1
rlabel polysilicon 212 -666 212 -666 0 3
rlabel polysilicon 219 -660 219 -660 0 1
rlabel polysilicon 219 -666 219 -666 0 3
rlabel polysilicon 226 -660 226 -660 0 1
rlabel polysilicon 226 -666 226 -666 0 3
rlabel polysilicon 233 -660 233 -660 0 1
rlabel polysilicon 233 -666 233 -666 0 3
rlabel polysilicon 240 -660 240 -660 0 1
rlabel polysilicon 240 -666 240 -666 0 3
rlabel polysilicon 247 -660 247 -660 0 1
rlabel polysilicon 247 -666 247 -666 0 3
rlabel polysilicon 254 -660 254 -660 0 1
rlabel polysilicon 254 -666 254 -666 0 3
rlabel polysilicon 261 -660 261 -660 0 1
rlabel polysilicon 261 -666 261 -666 0 3
rlabel polysilicon 268 -660 268 -660 0 1
rlabel polysilicon 268 -666 268 -666 0 3
rlabel polysilicon 275 -660 275 -660 0 1
rlabel polysilicon 275 -666 275 -666 0 3
rlabel polysilicon 282 -660 282 -660 0 1
rlabel polysilicon 282 -666 282 -666 0 3
rlabel polysilicon 289 -660 289 -660 0 1
rlabel polysilicon 289 -666 289 -666 0 3
rlabel polysilicon 296 -660 296 -660 0 1
rlabel polysilicon 61 -693 61 -693 0 2
rlabel polysilicon 61 -699 61 -699 0 4
rlabel polysilicon 72 -699 72 -699 0 3
rlabel polysilicon 75 -699 75 -699 0 4
rlabel polysilicon 79 -693 79 -693 0 1
rlabel polysilicon 79 -699 79 -699 0 3
rlabel polysilicon 89 -693 89 -693 0 2
rlabel polysilicon 93 -693 93 -693 0 1
rlabel polysilicon 93 -699 93 -699 0 3
rlabel polysilicon 100 -693 100 -693 0 1
rlabel polysilicon 100 -699 100 -699 0 3
rlabel polysilicon 107 -693 107 -693 0 1
rlabel polysilicon 110 -693 110 -693 0 2
rlabel polysilicon 114 -699 114 -699 0 3
rlabel polysilicon 117 -699 117 -699 0 4
rlabel polysilicon 121 -693 121 -693 0 1
rlabel polysilicon 121 -699 121 -699 0 3
rlabel polysilicon 128 -693 128 -693 0 1
rlabel polysilicon 128 -699 128 -699 0 3
rlabel polysilicon 138 -693 138 -693 0 2
rlabel polysilicon 142 -693 142 -693 0 1
rlabel polysilicon 142 -699 142 -699 0 3
rlabel polysilicon 152 -699 152 -699 0 4
rlabel polysilicon 156 -693 156 -693 0 1
rlabel polysilicon 163 -693 163 -693 0 1
rlabel polysilicon 163 -699 163 -699 0 3
rlabel polysilicon 170 -693 170 -693 0 1
rlabel polysilicon 170 -699 170 -699 0 3
rlabel polysilicon 177 -693 177 -693 0 1
rlabel polysilicon 180 -693 180 -693 0 2
rlabel polysilicon 177 -699 177 -699 0 3
rlabel polysilicon 187 -693 187 -693 0 2
rlabel polysilicon 187 -699 187 -699 0 4
rlabel polysilicon 191 -693 191 -693 0 1
rlabel polysilicon 194 -699 194 -699 0 4
rlabel polysilicon 198 -693 198 -693 0 1
rlabel polysilicon 198 -699 198 -699 0 3
rlabel polysilicon 205 -693 205 -693 0 1
rlabel polysilicon 205 -699 205 -699 0 3
rlabel polysilicon 212 -693 212 -693 0 1
rlabel polysilicon 219 -693 219 -693 0 1
rlabel polysilicon 219 -699 219 -699 0 3
rlabel polysilicon 226 -693 226 -693 0 1
rlabel polysilicon 226 -699 226 -699 0 3
rlabel polysilicon 233 -693 233 -693 0 1
rlabel polysilicon 233 -699 233 -699 0 3
rlabel polysilicon 240 -693 240 -693 0 1
rlabel polysilicon 240 -699 240 -699 0 3
rlabel polysilicon 247 -699 247 -699 0 3
rlabel polysilicon 254 -693 254 -693 0 1
rlabel polysilicon 254 -699 254 -699 0 3
rlabel polysilicon 261 -699 261 -699 0 3
rlabel polysilicon 268 -693 268 -693 0 1
rlabel polysilicon 268 -699 268 -699 0 3
rlabel polysilicon 278 -693 278 -693 0 2
rlabel polysilicon 114 -722 114 -722 0 3
rlabel polysilicon 121 -716 121 -716 0 1
rlabel polysilicon 121 -722 121 -722 0 3
rlabel polysilicon 131 -716 131 -716 0 2
rlabel polysilicon 131 -722 131 -722 0 4
rlabel polysilicon 135 -716 135 -716 0 1
rlabel polysilicon 142 -716 142 -716 0 1
rlabel polysilicon 142 -722 142 -722 0 3
rlabel polysilicon 149 -716 149 -716 0 1
rlabel polysilicon 163 -716 163 -716 0 1
rlabel polysilicon 163 -722 163 -722 0 3
rlabel polysilicon 170 -716 170 -716 0 1
rlabel polysilicon 173 -716 173 -716 0 2
rlabel polysilicon 173 -722 173 -722 0 4
rlabel polysilicon 180 -716 180 -716 0 2
rlabel polysilicon 177 -722 177 -722 0 3
rlabel polysilicon 180 -722 180 -722 0 4
rlabel polysilicon 184 -716 184 -716 0 1
rlabel polysilicon 184 -722 184 -722 0 3
rlabel polysilicon 194 -716 194 -716 0 2
rlabel polysilicon 191 -722 191 -722 0 3
rlabel polysilicon 194 -722 194 -722 0 4
rlabel polysilicon 198 -716 198 -716 0 1
rlabel polysilicon 198 -722 198 -722 0 3
rlabel polysilicon 205 -716 205 -716 0 1
rlabel polysilicon 205 -722 205 -722 0 3
rlabel polysilicon 215 -716 215 -716 0 2
rlabel polysilicon 229 -722 229 -722 0 4
rlabel polysilicon 240 -716 240 -716 0 1
rlabel polysilicon 240 -722 240 -722 0 3
rlabel polysilicon 117 -731 117 -731 0 2
rlabel polysilicon 121 -731 121 -731 0 1
rlabel polysilicon 121 -737 121 -737 0 3
rlabel polysilicon 131 -731 131 -731 0 2
rlabel polysilicon 128 -737 128 -737 0 3
rlabel polysilicon 135 -731 135 -731 0 1
rlabel polysilicon 135 -737 135 -737 0 3
rlabel polysilicon 159 -731 159 -731 0 2
rlabel polysilicon 156 -737 156 -737 0 3
rlabel polysilicon 166 -737 166 -737 0 4
rlabel polysilicon 170 -731 170 -731 0 1
rlabel polysilicon 170 -737 170 -737 0 3
rlabel polysilicon 177 -731 177 -731 0 1
rlabel polysilicon 177 -737 177 -737 0 3
rlabel polysilicon 184 -731 184 -731 0 1
rlabel polysilicon 187 -737 187 -737 0 4
rlabel polysilicon 191 -731 191 -731 0 1
rlabel polysilicon 191 -737 191 -737 0 3
rlabel polysilicon 124 -750 124 -750 0 4
rlabel polysilicon 128 -744 128 -744 0 1
rlabel polysilicon 128 -750 128 -750 0 3
rlabel polysilicon 149 -744 149 -744 0 1
rlabel polysilicon 156 -750 156 -750 0 3
rlabel polysilicon 159 -750 159 -750 0 4
rlabel polysilicon 163 -744 163 -744 0 1
rlabel polysilicon 163 -750 163 -750 0 3
rlabel polysilicon 170 -744 170 -744 0 1
rlabel polysilicon 170 -750 170 -750 0 3
rlabel polysilicon 184 -744 184 -744 0 1
rlabel polysilicon 184 -750 184 -750 0 3
rlabel polysilicon 191 -750 191 -750 0 3
rlabel metal2 103 1 103 1 0 net=200
rlabel metal2 128 1 128 1 0 net=539
rlabel metal2 142 1 142 1 0 net=757
rlabel metal2 177 1 177 1 0 net=969
rlabel metal2 194 1 194 1 0 net=781
rlabel metal2 198 -1 198 -1 0 net=737
rlabel metal2 79 -12 79 -12 0 net=407
rlabel metal2 100 -12 100 -12 0 net=106
rlabel metal2 110 -12 110 -12 0 net=1161
rlabel metal2 135 -12 135 -12 0 net=540
rlabel metal2 149 -12 149 -12 0 net=758
rlabel metal2 170 -12 170 -12 0 net=1031
rlabel metal2 208 -12 208 -12 0 net=1121
rlabel metal2 135 -14 135 -14 0 net=783
rlabel metal2 177 -14 177 -14 0 net=970
rlabel metal2 212 -14 212 -14 0 net=782
rlabel metal2 142 -16 142 -16 0 net=777
rlabel metal2 184 -16 184 -16 0 net=738
rlabel metal2 215 -16 215 -16 0 net=1111
rlabel metal2 149 -18 149 -18 0 net=263
rlabel metal2 152 -20 152 -20 0 net=719
rlabel metal2 65 -31 65 -31 0 net=533
rlabel metal2 93 -31 93 -31 0 net=787
rlabel metal2 114 -31 114 -31 0 net=457
rlabel metal2 184 -31 184 -31 0 net=1259
rlabel metal2 271 -31 271 -31 0 net=985
rlabel metal2 72 -33 72 -33 0 net=807
rlabel metal2 128 -33 128 -33 0 net=185
rlabel metal2 128 -33 128 -33 0 net=185
rlabel metal2 142 -33 142 -33 0 net=778
rlabel metal2 198 -33 198 -33 0 net=721
rlabel metal2 229 -33 229 -33 0 net=909
rlabel metal2 79 -35 79 -35 0 net=408
rlabel metal2 79 -35 79 -35 0 net=408
rlabel metal2 86 -35 86 -35 0 net=21
rlabel metal2 93 -35 93 -35 0 net=271
rlabel metal2 149 -35 149 -35 0 net=1032
rlabel metal2 180 -35 180 -35 0 net=1239
rlabel metal2 201 -35 201 -35 0 net=1373
rlabel metal2 86 -37 86 -37 0 net=293
rlabel metal2 135 -37 135 -37 0 net=784
rlabel metal2 152 -37 152 -37 0 net=1401
rlabel metal2 121 -39 121 -39 0 net=1163
rlabel metal2 156 -39 156 -39 0 net=503
rlabel metal2 215 -39 215 -39 0 net=1112
rlabel metal2 233 -39 233 -39 0 net=1123
rlabel metal2 156 -41 156 -41 0 net=817
rlabel metal2 191 -41 191 -41 0 net=1359
rlabel metal2 159 -43 159 -43 0 net=111
rlabel metal2 177 -43 177 -43 0 net=729
rlabel metal2 205 -43 205 -43 0 net=1393
rlabel metal2 30 -54 30 -54 0 net=1433
rlabel metal2 82 -54 82 -54 0 net=10
rlabel metal2 170 -54 170 -54 0 net=1124
rlabel metal2 44 -56 44 -56 0 net=459
rlabel metal2 117 -56 117 -56 0 net=1179
rlabel metal2 163 -56 163 -56 0 net=505
rlabel metal2 184 -56 184 -56 0 net=1241
rlabel metal2 51 -58 51 -58 0 net=1045
rlabel metal2 159 -58 159 -58 0 net=599
rlabel metal2 187 -58 187 -58 0 net=1385
rlabel metal2 58 -60 58 -60 0 net=819
rlabel metal2 191 -60 191 -60 0 net=730
rlabel metal2 201 -60 201 -60 0 net=1402
rlabel metal2 243 -60 243 -60 0 net=1387
rlabel metal2 61 -62 61 -62 0 net=180
rlabel metal2 93 -62 93 -62 0 net=479
rlabel metal2 198 -62 198 -62 0 net=722
rlabel metal2 233 -62 233 -62 0 net=1361
rlabel metal2 65 -64 65 -64 0 net=535
rlabel metal2 100 -64 100 -64 0 net=788
rlabel metal2 121 -64 121 -64 0 net=1164
rlabel metal2 142 -64 142 -64 0 net=685
rlabel metal2 219 -64 219 -64 0 net=987
rlabel metal2 65 -66 65 -66 0 net=523
rlabel metal2 100 -66 100 -66 0 net=218
rlabel metal2 180 -66 180 -66 0 net=663
rlabel metal2 254 -66 254 -66 0 net=1375
rlabel metal2 72 -68 72 -68 0 net=808
rlabel metal2 184 -68 184 -68 0 net=701
rlabel metal2 72 -70 72 -70 0 net=753
rlabel metal2 103 -70 103 -70 0 net=647
rlabel metal2 212 -70 212 -70 0 net=1053
rlabel metal2 110 -72 110 -72 0 net=78
rlabel metal2 205 -72 205 -72 0 net=1394
rlabel metal2 222 -72 222 -72 0 net=910
rlabel metal2 121 -74 121 -74 0 net=507
rlabel metal2 247 -74 247 -74 0 net=1261
rlabel metal2 16 -85 16 -85 0 net=755
rlabel metal2 86 -85 86 -85 0 net=536
rlabel metal2 103 -85 103 -85 0 net=341
rlabel metal2 114 -85 114 -85 0 net=149
rlabel metal2 170 -85 170 -85 0 net=506
rlabel metal2 184 -85 184 -85 0 net=228
rlabel metal2 201 -85 201 -85 0 net=38
rlabel metal2 243 -85 243 -85 0 net=1262
rlabel metal2 299 -85 299 -85 0 net=1251
rlabel metal2 30 -87 30 -87 0 net=1435
rlabel metal2 26 -89 26 -89 0 net=485
rlabel metal2 37 -89 37 -89 0 net=72
rlabel metal2 100 -89 100 -89 0 net=365
rlabel metal2 250 -89 250 -89 0 net=1386
rlabel metal2 37 -91 37 -91 0 net=481
rlabel metal2 107 -91 107 -91 0 net=491
rlabel metal2 131 -91 131 -91 0 net=664
rlabel metal2 254 -91 254 -91 0 net=1055
rlabel metal2 254 -91 254 -91 0 net=1055
rlabel metal2 268 -91 268 -91 0 net=1363
rlabel metal2 44 -93 44 -93 0 net=460
rlabel metal2 138 -93 138 -93 0 net=1093
rlabel metal2 51 -95 51 -95 0 net=1046
rlabel metal2 191 -95 191 -95 0 net=687
rlabel metal2 275 -95 275 -95 0 net=1377
rlabel metal2 58 -97 58 -97 0 net=820
rlabel metal2 142 -97 142 -97 0 net=649
rlabel metal2 65 -99 65 -99 0 net=525
rlabel metal2 93 -99 93 -99 0 net=475
rlabel metal2 163 -99 163 -99 0 net=601
rlabel metal2 177 -99 177 -99 0 net=1242
rlabel metal2 51 -101 51 -101 0 net=437
rlabel metal2 68 -101 68 -101 0 net=18
rlabel metal2 180 -101 180 -101 0 net=615
rlabel metal2 219 -101 219 -101 0 net=989
rlabel metal2 72 -103 72 -103 0 net=665
rlabel metal2 128 -103 128 -103 0 net=120
rlabel metal2 187 -103 187 -103 0 net=927
rlabel metal2 117 -105 117 -105 0 net=653
rlabel metal2 198 -107 198 -107 0 net=1113
rlabel metal2 198 -109 198 -109 0 net=1388
rlabel metal2 149 -111 149 -111 0 net=1181
rlabel metal2 121 -113 121 -113 0 net=508
rlabel metal2 201 -113 201 -113 0 net=702
rlabel metal2 205 -115 205 -115 0 net=1153
rlabel metal2 205 -117 205 -117 0 net=723
rlabel metal2 208 -119 208 -119 0 net=1231
rlabel metal2 23 -130 23 -130 0 net=119
rlabel metal2 159 -130 159 -130 0 net=688
rlabel metal2 275 -130 275 -130 0 net=1115
rlabel metal2 275 -130 275 -130 0 net=1115
rlabel metal2 26 -132 26 -132 0 net=486
rlabel metal2 37 -132 37 -132 0 net=482
rlabel metal2 198 -132 198 -132 0 net=724
rlabel metal2 23 -134 23 -134 0 net=1193
rlabel metal2 44 -134 44 -134 0 net=439
rlabel metal2 61 -134 61 -134 0 net=309
rlabel metal2 100 -134 100 -134 0 net=1094
rlabel metal2 37 -136 37 -136 0 net=213
rlabel metal2 65 -136 65 -136 0 net=1436
rlabel metal2 47 -138 47 -138 0 net=759
rlabel metal2 72 -138 72 -138 0 net=666
rlabel metal2 86 -138 86 -138 0 net=526
rlabel metal2 128 -138 128 -138 0 net=85
rlabel metal2 72 -140 72 -140 0 net=477
rlabel metal2 100 -140 100 -140 0 net=493
rlabel metal2 110 -140 110 -140 0 net=346
rlabel metal2 117 -140 117 -140 0 net=27
rlabel metal2 128 -140 128 -140 0 net=657
rlabel metal2 166 -140 166 -140 0 net=357
rlabel metal2 205 -140 205 -140 0 net=654
rlabel metal2 16 -142 16 -142 0 net=756
rlabel metal2 135 -142 135 -142 0 net=650
rlabel metal2 79 -144 79 -144 0 net=957
rlabel metal2 142 -144 142 -144 0 net=1182
rlabel metal2 79 -146 79 -146 0 net=939
rlabel metal2 170 -146 170 -146 0 net=602
rlabel metal2 205 -146 205 -146 0 net=1364
rlabel metal2 131 -148 131 -148 0 net=593
rlabel metal2 177 -148 177 -148 0 net=42
rlabel metal2 201 -148 201 -148 0 net=1297
rlabel metal2 103 -150 103 -150 0 net=821
rlabel metal2 201 -150 201 -150 0 net=1219
rlabel metal2 303 -150 303 -150 0 net=1253
rlabel metal2 142 -152 142 -152 0 net=433
rlabel metal2 215 -152 215 -152 0 net=1154
rlabel metal2 156 -154 156 -154 0 net=1029
rlabel metal2 219 -154 219 -154 0 net=1233
rlabel metal2 219 -154 219 -154 0 net=1233
rlabel metal2 226 -154 226 -154 0 net=991
rlabel metal2 233 -154 233 -154 0 net=1307
rlabel metal2 212 -156 212 -156 0 net=616
rlabel metal2 236 -156 236 -156 0 net=1378
rlabel metal2 212 -158 212 -158 0 net=1019
rlabel metal2 226 -160 226 -160 0 net=929
rlabel metal2 236 -162 236 -162 0 net=1171
rlabel metal2 254 -164 254 -164 0 net=1057
rlabel metal2 16 -177 16 -177 0 net=995
rlabel metal2 37 -177 37 -177 0 net=411
rlabel metal2 72 -177 72 -177 0 net=478
rlabel metal2 89 -177 89 -177 0 net=339
rlabel metal2 121 -177 121 -177 0 net=659
rlabel metal2 135 -177 135 -177 0 net=434
rlabel metal2 145 -177 145 -177 0 net=1449
rlabel metal2 9 -179 9 -179 0 net=1001
rlabel metal2 100 -179 100 -179 0 net=495
rlabel metal2 100 -179 100 -179 0 net=495
rlabel metal2 149 -179 149 -179 0 net=877
rlabel metal2 222 -179 222 -179 0 net=1308
rlabel metal2 303 -179 303 -179 0 net=1255
rlabel metal2 19 -181 19 -181 0 net=352
rlabel metal2 72 -181 72 -181 0 net=901
rlabel metal2 149 -181 149 -181 0 net=1030
rlabel metal2 191 -181 191 -181 0 net=555
rlabel metal2 240 -181 240 -181 0 net=1058
rlabel metal2 268 -181 268 -181 0 net=1167
rlabel metal2 23 -183 23 -183 0 net=1194
rlabel metal2 44 -183 44 -183 0 net=440
rlabel metal2 54 -183 54 -183 0 net=873
rlabel metal2 79 -183 79 -183 0 net=940
rlabel metal2 117 -183 117 -183 0 net=1095
rlabel metal2 243 -183 243 -183 0 net=1151
rlabel metal2 44 -185 44 -185 0 net=575
rlabel metal2 194 -185 194 -185 0 net=930
rlabel metal2 247 -185 247 -185 0 net=1021
rlabel metal2 271 -185 271 -185 0 net=1075
rlabel metal2 310 -185 310 -185 0 net=1299
rlabel metal2 51 -187 51 -187 0 net=958
rlabel metal2 107 -187 107 -187 0 net=319
rlabel metal2 247 -187 247 -187 0 net=895
rlabel metal2 65 -189 65 -189 0 net=761
rlabel metal2 93 -189 93 -189 0 net=839
rlabel metal2 212 -189 212 -189 0 net=1211
rlabel metal2 117 -191 117 -191 0 net=186
rlabel metal2 156 -191 156 -191 0 net=405
rlabel metal2 170 -191 170 -191 0 net=594
rlabel metal2 275 -191 275 -191 0 net=1117
rlabel metal2 114 -193 114 -193 0 net=861
rlabel metal2 282 -193 282 -193 0 net=1173
rlabel metal2 128 -195 128 -195 0 net=445
rlabel metal2 159 -195 159 -195 0 net=1234
rlabel metal2 285 -195 285 -195 0 net=1315
rlabel metal2 170 -197 170 -197 0 net=567
rlabel metal2 219 -197 219 -197 0 net=1407
rlabel metal2 177 -199 177 -199 0 net=823
rlabel metal2 289 -199 289 -199 0 net=1221
rlabel metal2 177 -201 177 -201 0 net=993
rlabel metal2 289 -201 289 -201 0 net=1223
rlabel metal2 201 -203 201 -203 0 net=905
rlabel metal2 292 -203 292 -203 0 net=1429
rlabel metal2 9 -214 9 -214 0 net=1002
rlabel metal2 149 -214 149 -214 0 net=775
rlabel metal2 187 -214 187 -214 0 net=1222
rlabel metal2 352 -214 352 -214 0 net=1317
rlabel metal2 352 -214 352 -214 0 net=1317
rlabel metal2 9 -216 9 -216 0 net=667
rlabel metal2 86 -216 86 -216 0 net=497
rlabel metal2 114 -216 114 -216 0 net=902
rlabel metal2 156 -216 156 -216 0 net=568
rlabel metal2 177 -216 177 -216 0 net=994
rlabel metal2 222 -216 222 -216 0 net=1300
rlabel metal2 16 -218 16 -218 0 net=996
rlabel metal2 72 -218 72 -218 0 net=762
rlabel metal2 93 -218 93 -218 0 net=840
rlabel metal2 163 -218 163 -218 0 net=406
rlabel metal2 261 -218 261 -218 0 net=1023
rlabel metal2 289 -218 289 -218 0 net=1152
rlabel metal2 16 -220 16 -220 0 net=537
rlabel metal2 128 -220 128 -220 0 net=447
rlabel metal2 170 -220 170 -220 0 net=625
rlabel metal2 229 -220 229 -220 0 net=1256
rlabel metal2 26 -222 26 -222 0 net=253
rlabel metal2 117 -222 117 -222 0 net=1408
rlabel metal2 30 -224 30 -224 0 net=557
rlabel metal2 215 -224 215 -224 0 net=1118
rlabel metal2 366 -224 366 -224 0 net=1431
rlabel metal2 37 -226 37 -226 0 net=413
rlabel metal2 191 -226 191 -226 0 net=907
rlabel metal2 268 -226 268 -226 0 net=1174
rlabel metal2 37 -228 37 -228 0 net=661
rlabel metal2 128 -228 128 -228 0 net=705
rlabel metal2 219 -228 219 -228 0 net=825
rlabel metal2 233 -228 233 -228 0 net=897
rlabel metal2 254 -228 254 -228 0 net=933
rlabel metal2 292 -228 292 -228 0 net=1423
rlabel metal2 44 -230 44 -230 0 net=577
rlabel metal2 198 -230 198 -230 0 net=879
rlabel metal2 296 -230 296 -230 0 net=1077
rlabel metal2 44 -232 44 -232 0 net=623
rlabel metal2 89 -232 89 -232 0 net=1439
rlabel metal2 51 -234 51 -234 0 net=875
rlabel metal2 72 -234 72 -234 0 net=252
rlabel metal2 93 -234 93 -234 0 net=613
rlabel metal2 114 -234 114 -234 0 net=427
rlabel metal2 240 -234 240 -234 0 net=1097
rlabel metal2 58 -236 58 -236 0 net=997
rlabel metal2 156 -236 156 -236 0 net=827
rlabel metal2 303 -236 303 -236 0 net=1213
rlabel metal2 121 -238 121 -238 0 net=1450
rlabel metal2 198 -240 198 -240 0 net=1168
rlabel metal2 208 -242 208 -242 0 net=1279
rlabel metal2 208 -244 208 -244 0 net=862
rlabel metal2 310 -244 310 -244 0 net=1225
rlabel metal2 331 -244 331 -244 0 net=1143
rlabel metal2 201 -246 201 -246 0 net=1059
rlabel metal2 240 -248 240 -248 0 net=955
rlabel metal2 2 -259 2 -259 0 net=1125
rlabel metal2 138 -259 138 -259 0 net=934
rlabel metal2 264 -259 264 -259 0 net=1078
rlabel metal2 345 -259 345 -259 0 net=1425
rlabel metal2 345 -259 345 -259 0 net=1425
rlabel metal2 359 -259 359 -259 0 net=1440
rlabel metal2 376 -259 376 -259 0 net=1432
rlabel metal2 9 -261 9 -261 0 net=668
rlabel metal2 79 -261 79 -261 0 net=331
rlabel metal2 121 -261 121 -261 0 net=9
rlabel metal2 166 -261 166 -261 0 net=731
rlabel metal2 275 -261 275 -261 0 net=1144
rlabel metal2 366 -261 366 -261 0 net=400
rlabel metal2 9 -263 9 -263 0 net=999
rlabel metal2 65 -263 65 -263 0 net=707
rlabel metal2 149 -263 149 -263 0 net=579
rlabel metal2 184 -263 184 -263 0 net=776
rlabel metal2 275 -263 275 -263 0 net=1025
rlabel metal2 289 -263 289 -263 0 net=1318
rlabel metal2 366 -263 366 -263 0 net=1367
rlabel metal2 16 -265 16 -265 0 net=538
rlabel metal2 107 -265 107 -265 0 net=735
rlabel metal2 212 -265 212 -265 0 net=826
rlabel metal2 247 -265 247 -265 0 net=829
rlabel metal2 289 -265 289 -265 0 net=1061
rlabel metal2 16 -267 16 -267 0 net=973
rlabel metal2 152 -267 152 -267 0 net=908
rlabel metal2 205 -267 205 -267 0 net=956
rlabel metal2 250 -267 250 -267 0 net=1287
rlabel metal2 37 -269 37 -269 0 net=662
rlabel metal2 215 -269 215 -269 0 net=1413
rlabel metal2 23 -271 23 -271 0 net=1105
rlabel metal2 233 -271 233 -271 0 net=898
rlabel metal2 296 -271 296 -271 0 net=1280
rlabel metal2 44 -273 44 -273 0 net=624
rlabel metal2 163 -273 163 -273 0 net=415
rlabel metal2 191 -273 191 -273 0 net=483
rlabel metal2 303 -273 303 -273 0 net=1215
rlabel metal2 51 -275 51 -275 0 net=876
rlabel metal2 68 -275 68 -275 0 net=375
rlabel metal2 86 -275 86 -275 0 net=499
rlabel metal2 170 -275 170 -275 0 net=627
rlabel metal2 303 -275 303 -275 0 net=1099
rlabel metal2 37 -277 37 -277 0 net=845
rlabel metal2 72 -277 72 -277 0 net=709
rlabel metal2 93 -277 93 -277 0 net=614
rlabel metal2 170 -277 170 -277 0 net=923
rlabel metal2 198 -277 198 -277 0 net=419
rlabel metal2 268 -277 268 -277 0 net=881
rlabel metal2 30 -279 30 -279 0 net=558
rlabel metal2 201 -279 201 -279 0 net=1281
rlabel metal2 30 -281 30 -281 0 net=739
rlabel metal2 205 -281 205 -281 0 net=1275
rlabel metal2 310 -281 310 -281 0 net=1227
rlabel metal2 44 -283 44 -283 0 net=655
rlabel metal2 61 -285 61 -285 0 net=1145
rlabel metal2 72 -287 72 -287 0 net=703
rlabel metal2 93 -289 93 -289 0 net=429
rlabel metal2 100 -291 100 -291 0 net=637
rlabel metal2 114 -293 114 -293 0 net=449
rlabel metal2 142 -295 142 -295 0 net=527
rlabel metal2 9 -306 9 -306 0 net=1000
rlabel metal2 68 -306 68 -306 0 net=704
rlabel metal2 79 -306 79 -306 0 net=587
rlabel metal2 107 -306 107 -306 0 net=736
rlabel metal2 240 -306 240 -306 0 net=1216
rlabel metal2 373 -306 373 -306 0 net=241
rlabel metal2 380 -306 380 -306 0 net=1369
rlabel metal2 9 -308 9 -308 0 net=847
rlabel metal2 72 -308 72 -308 0 net=711
rlabel metal2 110 -308 110 -308 0 net=924
rlabel metal2 173 -308 173 -308 0 net=484
rlabel metal2 198 -308 198 -308 0 net=645
rlabel metal2 250 -308 250 -308 0 net=1228
rlabel metal2 2 -310 2 -310 0 net=1126
rlabel metal2 124 -310 124 -310 0 net=580
rlabel metal2 152 -310 152 -310 0 net=420
rlabel metal2 296 -310 296 -310 0 net=1323
rlabel metal2 310 -310 310 -310 0 net=1146
rlabel metal2 2 -312 2 -312 0 net=893
rlabel metal2 159 -312 159 -312 0 net=1100
rlabel metal2 16 -314 16 -314 0 net=974
rlabel metal2 177 -314 177 -314 0 net=417
rlabel metal2 177 -314 177 -314 0 net=417
rlabel metal2 187 -314 187 -314 0 net=1414
rlabel metal2 23 -316 23 -316 0 net=1106
rlabel metal2 128 -316 128 -316 0 net=501
rlabel metal2 205 -316 205 -316 0 net=882
rlabel metal2 345 -316 345 -316 0 net=1427
rlabel metal2 23 -318 23 -318 0 net=651
rlabel metal2 93 -318 93 -318 0 net=430
rlabel metal2 208 -318 208 -318 0 net=1282
rlabel metal2 30 -320 30 -320 0 net=740
rlabel metal2 138 -320 138 -320 0 net=305
rlabel metal2 236 -320 236 -320 0 net=947
rlabel metal2 324 -320 324 -320 0 net=1289
rlabel metal2 338 -320 338 -320 0 net=797
rlabel metal2 30 -322 30 -322 0 net=529
rlabel metal2 145 -322 145 -322 0 net=1301
rlabel metal2 254 -322 254 -322 0 net=1283
rlabel metal2 37 -324 37 -324 0 net=451
rlabel metal2 135 -324 135 -324 0 net=441
rlabel metal2 268 -324 268 -324 0 net=1277
rlabel metal2 44 -326 44 -326 0 net=656
rlabel metal2 159 -326 159 -326 0 net=889
rlabel metal2 261 -326 261 -326 0 net=733
rlabel metal2 275 -326 275 -326 0 net=1027
rlabel metal2 44 -328 44 -328 0 net=617
rlabel metal2 93 -328 93 -328 0 net=551
rlabel metal2 163 -328 163 -328 0 net=1187
rlabel metal2 275 -328 275 -328 0 net=1063
rlabel metal2 100 -330 100 -330 0 net=639
rlabel metal2 163 -330 163 -330 0 net=401
rlabel metal2 212 -330 212 -330 0 net=1191
rlabel metal2 65 -332 65 -332 0 net=708
rlabel metal2 219 -332 219 -332 0 net=629
rlabel metal2 282 -332 282 -332 0 net=831
rlabel metal2 16 -334 16 -334 0 net=763
rlabel metal2 114 -334 114 -334 0 net=689
rlabel metal2 194 -336 194 -336 0 net=1415
rlabel metal2 2 -347 2 -347 0 net=894
rlabel metal2 170 -347 170 -347 0 net=1333
rlabel metal2 387 -347 387 -347 0 net=1371
rlabel metal2 387 -347 387 -347 0 net=1371
rlabel metal2 397 -347 397 -347 0 net=1229
rlabel metal2 9 -349 9 -349 0 net=848
rlabel metal2 51 -349 51 -349 0 net=619
rlabel metal2 51 -349 51 -349 0 net=619
rlabel metal2 61 -349 61 -349 0 net=204
rlabel metal2 194 -349 194 -349 0 net=832
rlabel metal2 324 -349 324 -349 0 net=1291
rlabel metal2 324 -349 324 -349 0 net=1291
rlabel metal2 331 -349 331 -349 0 net=1285
rlabel metal2 16 -351 16 -351 0 net=764
rlabel metal2 107 -351 107 -351 0 net=467
rlabel metal2 107 -351 107 -351 0 net=467
rlabel metal2 110 -351 110 -351 0 net=630
rlabel metal2 236 -351 236 -351 0 net=734
rlabel metal2 275 -351 275 -351 0 net=1065
rlabel metal2 275 -351 275 -351 0 net=1065
rlabel metal2 282 -351 282 -351 0 net=1417
rlabel metal2 16 -353 16 -353 0 net=713
rlabel metal2 86 -353 86 -353 0 net=91
rlabel metal2 142 -353 142 -353 0 net=361
rlabel metal2 142 -353 142 -353 0 net=361
rlabel metal2 170 -353 170 -353 0 net=1345
rlabel metal2 23 -355 23 -355 0 net=652
rlabel metal2 177 -355 177 -355 0 net=418
rlabel metal2 198 -355 198 -355 0 net=646
rlabel metal2 215 -355 215 -355 0 net=849
rlabel metal2 240 -355 240 -355 0 net=1278
rlabel metal2 23 -357 23 -357 0 net=1159
rlabel metal2 114 -357 114 -357 0 net=502
rlabel metal2 191 -357 191 -357 0 net=238
rlabel metal2 285 -357 285 -357 0 net=1428
rlabel metal2 30 -359 30 -359 0 net=530
rlabel metal2 163 -359 163 -359 0 net=403
rlabel metal2 198 -359 198 -359 0 net=549
rlabel metal2 247 -359 247 -359 0 net=1303
rlabel metal2 30 -361 30 -361 0 net=959
rlabel metal2 68 -361 68 -361 0 net=130
rlabel metal2 93 -361 93 -361 0 net=552
rlabel metal2 128 -361 128 -361 0 net=641
rlabel metal2 205 -361 205 -361 0 net=1137
rlabel metal2 296 -361 296 -361 0 net=1325
rlabel metal2 9 -363 9 -363 0 net=1349
rlabel metal2 100 -363 100 -363 0 net=857
rlabel metal2 208 -363 208 -363 0 net=867
rlabel metal2 37 -365 37 -365 0 net=452
rlabel metal2 212 -365 212 -365 0 net=1192
rlabel metal2 37 -367 37 -367 0 net=443
rlabel metal2 149 -367 149 -367 0 net=798
rlabel metal2 58 -369 58 -369 0 net=741
rlabel metal2 135 -369 135 -369 0 net=541
rlabel metal2 219 -369 219 -369 0 net=691
rlabel metal2 240 -369 240 -369 0 net=1271
rlabel metal2 72 -371 72 -371 0 net=435
rlabel metal2 121 -371 121 -371 0 net=863
rlabel metal2 219 -371 219 -371 0 net=1131
rlabel metal2 79 -373 79 -373 0 net=589
rlabel metal2 222 -373 222 -373 0 net=1028
rlabel metal2 44 -375 44 -375 0 net=1309
rlabel metal2 173 -375 173 -375 0 net=1155
rlabel metal2 243 -377 243 -377 0 net=948
rlabel metal2 247 -379 247 -379 0 net=891
rlabel metal2 261 -379 261 -379 0 net=1189
rlabel metal2 159 -381 159 -381 0 net=1047
rlabel metal2 271 -381 271 -381 0 net=1319
rlabel metal2 9 -392 9 -392 0 net=1350
rlabel metal2 170 -392 170 -392 0 net=590
rlabel metal2 240 -392 240 -392 0 net=1066
rlabel metal2 282 -392 282 -392 0 net=1292
rlabel metal2 373 -392 373 -392 0 net=1347
rlabel metal2 373 -392 373 -392 0 net=1347
rlabel metal2 387 -392 387 -392 0 net=1372
rlabel metal2 401 -392 401 -392 0 net=1230
rlabel metal2 16 -394 16 -394 0 net=714
rlabel metal2 131 -394 131 -394 0 net=324
rlabel metal2 184 -394 184 -394 0 net=56
rlabel metal2 243 -394 243 -394 0 net=40
rlabel metal2 243 -394 243 -394 0 net=40
rlabel metal2 268 -394 268 -394 0 net=1190
rlabel metal2 324 -394 324 -394 0 net=1335
rlabel metal2 23 -396 23 -396 0 net=1160
rlabel metal2 156 -396 156 -396 0 net=404
rlabel metal2 194 -396 194 -396 0 net=550
rlabel metal2 201 -396 201 -396 0 net=318
rlabel metal2 261 -396 261 -396 0 net=1049
rlabel metal2 296 -396 296 -396 0 net=1133
rlabel metal2 23 -398 23 -398 0 net=971
rlabel metal2 110 -398 110 -398 0 net=785
rlabel metal2 198 -398 198 -398 0 net=692
rlabel metal2 250 -398 250 -398 0 net=1293
rlabel metal2 296 -398 296 -398 0 net=1419
rlabel metal2 37 -400 37 -400 0 net=444
rlabel metal2 142 -400 142 -400 0 net=892
rlabel metal2 310 -400 310 -400 0 net=1321
rlabel metal2 30 -402 30 -402 0 net=960
rlabel metal2 58 -402 58 -402 0 net=743
rlabel metal2 58 -402 58 -402 0 net=743
rlabel metal2 65 -402 65 -402 0 net=112
rlabel metal2 128 -402 128 -402 0 net=543
rlabel metal2 149 -402 149 -402 0 net=425
rlabel metal2 226 -402 226 -402 0 net=981
rlabel metal2 331 -402 331 -402 0 net=869
rlabel metal2 30 -404 30 -404 0 net=621
rlabel metal2 65 -404 65 -404 0 net=850
rlabel metal2 285 -404 285 -404 0 net=843
rlabel metal2 338 -404 338 -404 0 net=1286
rlabel metal2 68 -406 68 -406 0 net=1267
rlabel metal2 72 -408 72 -408 0 net=436
rlabel metal2 233 -408 233 -408 0 net=1157
rlabel metal2 72 -410 72 -410 0 net=865
rlabel metal2 135 -410 135 -410 0 net=921
rlabel metal2 247 -410 247 -410 0 net=1399
rlabel metal2 79 -412 79 -412 0 net=20
rlabel metal2 107 -412 107 -412 0 net=469
rlabel metal2 156 -412 156 -412 0 net=841
rlabel metal2 303 -412 303 -412 0 net=1305
rlabel metal2 44 -414 44 -414 0 net=1311
rlabel metal2 86 -414 86 -414 0 net=859
rlabel metal2 114 -414 114 -414 0 net=358
rlabel metal2 317 -414 317 -414 0 net=1273
rlabel metal2 100 -416 100 -416 0 net=264
rlabel metal2 163 -416 163 -416 0 net=643
rlabel metal2 317 -416 317 -416 0 net=1327
rlabel metal2 121 -418 121 -418 0 net=699
rlabel metal2 163 -418 163 -418 0 net=269
rlabel metal2 289 -418 289 -418 0 net=1138
rlabel metal2 205 -420 205 -420 0 net=1329
rlabel metal2 23 -431 23 -431 0 net=972
rlabel metal2 58 -431 58 -431 0 net=745
rlabel metal2 58 -431 58 -431 0 net=745
rlabel metal2 65 -431 65 -431 0 net=396
rlabel metal2 107 -431 107 -431 0 net=545
rlabel metal2 142 -431 142 -431 0 net=471
rlabel metal2 159 -431 159 -431 0 net=644
rlabel metal2 191 -431 191 -431 0 net=1158
rlabel metal2 240 -431 240 -431 0 net=1051
rlabel metal2 282 -431 282 -431 0 net=1403
rlabel metal2 282 -431 282 -431 0 net=1403
rlabel metal2 306 -431 306 -431 0 net=1322
rlabel metal2 313 -431 313 -431 0 net=1400
rlabel metal2 352 -431 352 -431 0 net=1348
rlabel metal2 30 -433 30 -433 0 net=622
rlabel metal2 72 -433 72 -433 0 net=866
rlabel metal2 142 -433 142 -433 0 net=426
rlabel metal2 163 -433 163 -433 0 net=513
rlabel metal2 215 -433 215 -433 0 net=1328
rlabel metal2 320 -433 320 -433 0 net=1274
rlabel metal2 352 -433 352 -433 0 net=1135
rlabel metal2 37 -435 37 -435 0 net=1451
rlabel metal2 170 -435 170 -435 0 net=922
rlabel metal2 215 -435 215 -435 0 net=844
rlabel metal2 359 -435 359 -435 0 net=871
rlabel metal2 44 -437 44 -437 0 net=547
rlabel metal2 79 -437 79 -437 0 net=1313
rlabel metal2 79 -437 79 -437 0 net=1313
rlabel metal2 86 -437 86 -437 0 net=860
rlabel metal2 114 -437 114 -437 0 net=700
rlabel metal2 170 -437 170 -437 0 net=669
rlabel metal2 226 -437 226 -437 0 net=983
rlabel metal2 247 -437 247 -437 0 net=1306
rlabel metal2 362 -437 362 -437 0 net=793
rlabel metal2 51 -439 51 -439 0 net=561
rlabel metal2 229 -439 229 -439 0 net=1336
rlabel metal2 65 -441 65 -441 0 net=461
rlabel metal2 93 -441 93 -441 0 net=573
rlabel metal2 177 -441 177 -441 0 net=786
rlabel metal2 254 -441 254 -441 0 net=1294
rlabel metal2 268 -441 268 -441 0 net=1269
rlabel metal2 303 -441 303 -441 0 net=931
rlabel metal2 75 -443 75 -443 0 net=209
rlabel metal2 117 -443 117 -443 0 net=1013
rlabel metal2 275 -443 275 -443 0 net=1331
rlabel metal2 93 -445 93 -445 0 net=465
rlabel metal2 198 -445 198 -445 0 net=1205
rlabel metal2 289 -445 289 -445 0 net=1421
rlabel metal2 135 -447 135 -447 0 net=1107
rlabel metal2 191 -447 191 -447 0 net=1445
rlabel metal2 194 -449 194 -449 0 net=795
rlabel metal2 205 -449 205 -449 0 net=581
rlabel metal2 194 -451 194 -451 0 net=842
rlabel metal2 156 -453 156 -453 0 net=977
rlabel metal2 26 -464 26 -464 0 net=219
rlabel metal2 121 -464 121 -464 0 net=796
rlabel metal2 212 -464 212 -464 0 net=47
rlabel metal2 250 -464 250 -464 0 net=1332
rlabel metal2 296 -464 296 -464 0 net=1447
rlabel metal2 338 -464 338 -464 0 net=1136
rlabel metal2 366 -464 366 -464 0 net=794
rlabel metal2 33 -466 33 -466 0 net=332
rlabel metal2 79 -466 79 -466 0 net=1314
rlabel metal2 121 -466 121 -466 0 net=715
rlabel metal2 215 -466 215 -466 0 net=1052
rlabel metal2 254 -466 254 -466 0 net=1015
rlabel metal2 37 -468 37 -468 0 net=1452
rlabel metal2 142 -468 142 -468 0 net=583
rlabel metal2 240 -468 240 -468 0 net=1422
rlabel metal2 317 -468 317 -468 0 net=872
rlabel metal2 37 -470 37 -470 0 net=487
rlabel metal2 149 -470 149 -470 0 net=473
rlabel metal2 177 -470 177 -470 0 net=1109
rlabel metal2 261 -470 261 -470 0 net=1207
rlabel metal2 331 -470 331 -470 0 net=932
rlabel metal2 44 -472 44 -472 0 net=548
rlabel metal2 72 -472 72 -472 0 net=463
rlabel metal2 93 -472 93 -472 0 net=466
rlabel metal2 177 -472 177 -472 0 net=979
rlabel metal2 275 -472 275 -472 0 net=1343
rlabel metal2 331 -472 331 -472 0 net=1337
rlabel metal2 44 -474 44 -474 0 net=765
rlabel metal2 86 -474 86 -474 0 net=409
rlabel metal2 135 -474 135 -474 0 net=515
rlabel metal2 184 -474 184 -474 0 net=693
rlabel metal2 282 -474 282 -474 0 net=1405
rlabel metal2 58 -476 58 -476 0 net=747
rlabel metal2 107 -476 107 -476 0 net=546
rlabel metal2 163 -476 163 -476 0 net=671
rlabel metal2 187 -476 187 -476 0 net=1270
rlabel metal2 51 -478 51 -478 0 net=563
rlabel metal2 128 -478 128 -478 0 net=1355
rlabel metal2 170 -478 170 -478 0 net=1195
rlabel metal2 51 -480 51 -480 0 net=1397
rlabel metal2 173 -480 173 -480 0 net=975
rlabel metal2 100 -482 100 -482 0 net=574
rlabel metal2 191 -482 191 -482 0 net=984
rlabel metal2 100 -484 100 -484 0 net=519
rlabel metal2 194 -484 194 -484 0 net=941
rlabel metal2 198 -486 198 -486 0 net=1147
rlabel metal2 205 -488 205 -488 0 net=246
rlabel metal2 233 -490 233 -490 0 net=885
rlabel metal2 16 -501 16 -501 0 net=803
rlabel metal2 156 -501 156 -501 0 net=474
rlabel metal2 177 -501 177 -501 0 net=980
rlabel metal2 201 -501 201 -501 0 net=353
rlabel metal2 212 -501 212 -501 0 net=633
rlabel metal2 212 -501 212 -501 0 net=633
rlabel metal2 222 -501 222 -501 0 net=266
rlabel metal2 338 -501 338 -501 0 net=1441
rlabel metal2 30 -503 30 -503 0 net=767
rlabel metal2 51 -503 51 -503 0 net=1398
rlabel metal2 254 -503 254 -503 0 net=943
rlabel metal2 254 -503 254 -503 0 net=943
rlabel metal2 268 -503 268 -503 0 net=976
rlabel metal2 345 -503 345 -503 0 net=314
rlabel metal2 352 -503 352 -503 0 net=1017
rlabel metal2 65 -505 65 -505 0 net=748
rlabel metal2 86 -505 86 -505 0 net=410
rlabel metal2 110 -505 110 -505 0 net=232
rlabel metal2 159 -505 159 -505 0 net=1110
rlabel metal2 275 -505 275 -505 0 net=1344
rlabel metal2 317 -505 317 -505 0 net=1007
rlabel metal2 51 -507 51 -507 0 net=609
rlabel metal2 163 -507 163 -507 0 net=672
rlabel metal2 226 -507 226 -507 0 net=1406
rlabel metal2 296 -507 296 -507 0 net=1339
rlabel metal2 341 -507 341 -507 0 net=899
rlabel metal2 44 -509 44 -509 0 net=489
rlabel metal2 208 -509 208 -509 0 net=1237
rlabel metal2 341 -509 341 -509 0 net=815
rlabel metal2 65 -511 65 -511 0 net=585
rlabel metal2 149 -511 149 -511 0 net=1356
rlabel metal2 166 -511 166 -511 0 net=949
rlabel metal2 68 -513 68 -513 0 net=81
rlabel metal2 170 -513 170 -513 0 net=603
rlabel metal2 282 -513 282 -513 0 net=1448
rlabel metal2 72 -515 72 -515 0 net=464
rlabel metal2 191 -515 191 -515 0 net=93
rlabel metal2 233 -515 233 -515 0 net=887
rlabel metal2 247 -515 247 -515 0 net=1149
rlabel metal2 289 -515 289 -515 0 net=1209
rlabel metal2 37 -517 37 -517 0 net=488
rlabel metal2 79 -517 79 -517 0 net=851
rlabel metal2 194 -517 194 -517 0 net=883
rlabel metal2 261 -517 261 -517 0 net=1197
rlabel metal2 37 -519 37 -519 0 net=565
rlabel metal2 86 -519 86 -519 0 net=521
rlabel metal2 114 -519 114 -519 0 net=398
rlabel metal2 229 -519 229 -519 0 net=911
rlabel metal2 58 -521 58 -521 0 net=717
rlabel metal2 142 -521 142 -521 0 net=725
rlabel metal2 100 -523 100 -523 0 net=1033
rlabel metal2 114 -525 114 -525 0 net=517
rlabel metal2 201 -525 201 -525 0 net=809
rlabel metal2 135 -527 135 -527 0 net=695
rlabel metal2 177 -529 177 -529 0 net=749
rlabel metal2 9 -540 9 -540 0 net=1257
rlabel metal2 121 -540 121 -540 0 net=53
rlabel metal2 156 -540 156 -540 0 net=1035
rlabel metal2 222 -540 222 -540 0 net=1238
rlabel metal2 338 -540 338 -540 0 net=1018
rlabel metal2 16 -542 16 -542 0 net=804
rlabel metal2 275 -542 275 -542 0 net=1210
rlabel metal2 296 -542 296 -542 0 net=1341
rlabel metal2 296 -542 296 -542 0 net=1341
rlabel metal2 348 -542 348 -542 0 net=900
rlabel metal2 359 -542 359 -542 0 net=1443
rlabel metal2 359 -542 359 -542 0 net=1443
rlabel metal2 16 -544 16 -544 0 net=611
rlabel metal2 58 -544 58 -544 0 net=718
rlabel metal2 177 -544 177 -544 0 net=750
rlabel metal2 208 -544 208 -544 0 net=35
rlabel metal2 23 -546 23 -546 0 net=28
rlabel metal2 37 -546 37 -546 0 net=566
rlabel metal2 86 -546 86 -546 0 net=522
rlabel metal2 131 -546 131 -546 0 net=368
rlabel metal2 44 -548 44 -548 0 net=490
rlabel metal2 142 -548 142 -548 0 net=1263
rlabel metal2 226 -548 226 -548 0 net=811
rlabel metal2 275 -548 275 -548 0 net=816
rlabel metal2 30 -550 30 -550 0 net=768
rlabel metal2 58 -550 58 -550 0 net=853
rlabel metal2 86 -550 86 -550 0 net=607
rlabel metal2 114 -550 114 -550 0 net=518
rlabel metal2 145 -550 145 -550 0 net=884
rlabel metal2 254 -550 254 -550 0 net=945
rlabel metal2 65 -552 65 -552 0 net=586
rlabel metal2 177 -552 177 -552 0 net=1175
rlabel metal2 247 -552 247 -552 0 net=1183
rlabel metal2 65 -554 65 -554 0 net=1437
rlabel metal2 191 -554 191 -554 0 net=727
rlabel metal2 268 -554 268 -554 0 net=1034
rlabel metal2 72 -556 72 -556 0 net=697
rlabel metal2 201 -556 201 -556 0 net=1150
rlabel metal2 93 -558 93 -558 0 net=888
rlabel metal2 268 -558 268 -558 0 net=1199
rlabel metal2 93 -560 93 -560 0 net=1379
rlabel metal2 240 -560 240 -560 0 net=913
rlabel metal2 317 -560 317 -560 0 net=1009
rlabel metal2 100 -562 100 -562 0 net=5
rlabel metal2 282 -562 282 -562 0 net=1357
rlabel metal2 303 -562 303 -562 0 net=951
rlabel metal2 100 -564 100 -564 0 net=1081
rlabel metal2 135 -564 135 -564 0 net=679
rlabel metal2 198 -564 198 -564 0 net=635
rlabel metal2 114 -566 114 -566 0 net=569
rlabel metal2 170 -566 170 -566 0 net=605
rlabel metal2 163 -568 163 -568 0 net=769
rlabel metal2 9 -579 9 -579 0 net=1258
rlabel metal2 159 -579 159 -579 0 net=636
rlabel metal2 205 -579 205 -579 0 net=1265
rlabel metal2 257 -579 257 -579 0 net=946
rlabel metal2 282 -579 282 -579 0 net=1358
rlabel metal2 324 -579 324 -579 0 net=1011
rlabel metal2 324 -579 324 -579 0 net=1011
rlabel metal2 355 -579 355 -579 0 net=1444
rlabel metal2 16 -581 16 -581 0 net=612
rlabel metal2 65 -581 65 -581 0 net=1438
rlabel metal2 100 -581 100 -581 0 net=1082
rlabel metal2 135 -581 135 -581 0 net=681
rlabel metal2 187 -581 187 -581 0 net=728
rlabel metal2 198 -581 198 -581 0 net=1037
rlabel metal2 226 -581 226 -581 0 net=813
rlabel metal2 261 -581 261 -581 0 net=1201
rlabel metal2 282 -581 282 -581 0 net=1083
rlabel metal2 23 -583 23 -583 0 net=98
rlabel metal2 23 -583 23 -583 0 net=98
rlabel metal2 30 -583 30 -583 0 net=1365
rlabel metal2 86 -583 86 -583 0 net=608
rlabel metal2 163 -583 163 -583 0 net=771
rlabel metal2 205 -583 205 -583 0 net=1087
rlabel metal2 268 -583 268 -583 0 net=1139
rlabel metal2 289 -583 289 -583 0 net=953
rlabel metal2 40 -585 40 -585 0 net=150
rlabel metal2 40 -585 40 -585 0 net=150
rlabel metal2 44 -585 44 -585 0 net=1249
rlabel metal2 44 -585 44 -585 0 net=1249
rlabel metal2 51 -585 51 -585 0 net=773
rlabel metal2 135 -585 135 -585 0 net=141
rlabel metal2 163 -585 163 -585 0 net=509
rlabel metal2 219 -585 219 -585 0 net=915
rlabel metal2 296 -585 296 -585 0 net=1342
rlabel metal2 58 -587 58 -587 0 net=855
rlabel metal2 72 -587 72 -587 0 net=698
rlabel metal2 177 -587 177 -587 0 net=1176
rlabel metal2 58 -589 58 -589 0 net=1119
rlabel metal2 152 -589 152 -589 0 net=606
rlabel metal2 75 -591 75 -591 0 net=340
rlabel metal2 170 -591 170 -591 0 net=1067
rlabel metal2 212 -591 212 -591 0 net=1185
rlabel metal2 86 -593 86 -593 0 net=571
rlabel metal2 159 -593 159 -593 0 net=1409
rlabel metal2 93 -595 93 -595 0 net=1380
rlabel metal2 114 -595 114 -595 0 net=1389
rlabel metal2 79 -597 79 -597 0 net=110
rlabel metal2 107 -597 107 -597 0 net=935
rlabel metal2 33 -599 33 -599 0 net=171
rlabel metal2 26 -610 26 -610 0 net=202
rlabel metal2 26 -610 26 -610 0 net=202
rlabel metal2 30 -610 30 -610 0 net=1366
rlabel metal2 100 -610 100 -610 0 net=225
rlabel metal2 114 -610 114 -610 0 net=925
rlabel metal2 131 -610 131 -610 0 net=104
rlabel metal2 156 -610 156 -610 0 net=51
rlabel metal2 184 -610 184 -610 0 net=1186
rlabel metal2 226 -610 226 -610 0 net=814
rlabel metal2 257 -610 257 -610 0 net=1084
rlabel metal2 324 -610 324 -610 0 net=1012
rlabel metal2 324 -610 324 -610 0 net=1012
rlabel metal2 37 -612 37 -612 0 net=1250
rlabel metal2 51 -612 51 -612 0 net=774
rlabel metal2 135 -612 135 -612 0 net=772
rlabel metal2 205 -612 205 -612 0 net=1089
rlabel metal2 233 -612 233 -612 0 net=1266
rlabel metal2 275 -612 275 -612 0 net=954
rlabel metal2 51 -614 51 -614 0 net=1381
rlabel metal2 86 -614 86 -614 0 net=572
rlabel metal2 135 -614 135 -614 0 net=683
rlabel metal2 159 -614 159 -614 0 net=1038
rlabel metal2 205 -614 205 -614 0 net=917
rlabel metal2 233 -614 233 -614 0 net=1202
rlabel metal2 58 -616 58 -616 0 net=1120
rlabel metal2 142 -616 142 -616 0 net=779
rlabel metal2 163 -616 163 -616 0 net=510
rlabel metal2 177 -616 177 -616 0 net=257
rlabel metal2 187 -616 187 -616 0 net=965
rlabel metal2 240 -616 240 -616 0 net=1411
rlabel metal2 261 -616 261 -616 0 net=1140
rlabel metal2 65 -618 65 -618 0 net=856
rlabel metal2 114 -618 114 -618 0 net=304
rlabel metal2 152 -618 152 -618 0 net=1101
rlabel metal2 243 -618 243 -618 0 net=356
rlabel metal2 65 -620 65 -620 0 net=937
rlabel metal2 121 -620 121 -620 0 net=1391
rlabel metal2 170 -620 170 -620 0 net=1069
rlabel metal2 79 -622 79 -622 0 net=553
rlabel metal2 191 -622 191 -622 0 net=1295
rlabel metal2 75 -624 75 -624 0 net=247
rlabel metal2 93 -624 93 -624 0 net=675
rlabel metal2 30 -635 30 -635 0 net=1383
rlabel metal2 65 -635 65 -635 0 net=938
rlabel metal2 121 -635 121 -635 0 net=554
rlabel metal2 152 -635 152 -635 0 net=1296
rlabel metal2 201 -635 201 -635 0 net=1079
rlabel metal2 37 -637 37 -637 0 net=1085
rlabel metal2 82 -637 82 -637 0 net=32
rlabel metal2 107 -637 107 -637 0 net=1003
rlabel metal2 124 -637 124 -637 0 net=1392
rlabel metal2 184 -637 184 -637 0 net=1412
rlabel metal2 247 -637 247 -637 0 net=1235
rlabel metal2 44 -639 44 -639 0 net=591
rlabel metal2 96 -639 96 -639 0 net=87
rlabel metal2 254 -639 254 -639 0 net=1043
rlabel metal2 51 -641 51 -641 0 net=677
rlabel metal2 100 -641 100 -641 0 net=511
rlabel metal2 135 -641 135 -641 0 net=684
rlabel metal2 149 -641 149 -641 0 net=421
rlabel metal2 205 -641 205 -641 0 net=919
rlabel metal2 68 -643 68 -643 0 net=453
rlabel metal2 128 -643 128 -643 0 net=926
rlabel metal2 142 -643 142 -643 0 net=1351
rlabel metal2 75 -645 75 -645 0 net=631
rlabel metal2 128 -645 128 -645 0 net=595
rlabel metal2 156 -645 156 -645 0 net=780
rlabel metal2 187 -645 187 -645 0 net=214
rlabel metal2 156 -647 156 -647 0 net=673
rlabel metal2 170 -647 170 -647 0 net=1243
rlabel metal2 212 -649 212 -649 0 net=967
rlabel metal2 198 -651 198 -651 0 net=1071
rlabel metal2 219 -651 219 -651 0 net=1103
rlabel metal2 219 -653 219 -653 0 net=833
rlabel metal2 226 -655 226 -655 0 net=1091
rlabel metal2 191 -657 191 -657 0 net=903
rlabel metal2 37 -668 37 -668 0 net=1086
rlabel metal2 114 -668 114 -668 0 net=531
rlabel metal2 156 -668 156 -668 0 net=904
rlabel metal2 254 -668 254 -668 0 net=1044
rlabel metal2 44 -670 44 -670 0 net=592
rlabel metal2 156 -670 156 -670 0 net=674
rlabel metal2 173 -670 173 -670 0 net=1080
rlabel metal2 51 -672 51 -672 0 net=678
rlabel metal2 121 -672 121 -672 0 net=559
rlabel metal2 198 -672 198 -672 0 net=1073
rlabel metal2 247 -672 247 -672 0 net=1245
rlabel metal2 261 -672 261 -672 0 net=1353
rlabel metal2 58 -674 58 -674 0 net=632
rlabel metal2 89 -674 89 -674 0 net=250
rlabel metal2 159 -674 159 -674 0 net=342
rlabel metal2 205 -674 205 -674 0 net=1141
rlabel metal2 205 -674 205 -674 0 net=1141
rlabel metal2 208 -674 208 -674 0 net=1092
rlabel metal2 61 -676 61 -676 0 net=67
rlabel metal2 79 -676 79 -676 0 net=455
rlabel metal2 79 -676 79 -676 0 net=455
rlabel metal2 93 -676 93 -676 0 net=276
rlabel metal2 187 -676 187 -676 0 net=920
rlabel metal2 30 -678 30 -678 0 net=1384
rlabel metal2 93 -678 93 -678 0 net=423
rlabel metal2 180 -678 180 -678 0 net=1104
rlabel metal2 96 -680 96 -680 0 net=512
rlabel metal2 128 -680 128 -680 0 net=597
rlabel metal2 128 -680 128 -680 0 net=597
rlabel metal2 138 -680 138 -680 0 net=805
rlabel metal2 180 -680 180 -680 0 net=1236
rlabel metal2 100 -682 100 -682 0 net=1005
rlabel metal2 191 -682 191 -682 0 net=1127
rlabel metal2 107 -684 107 -684 0 net=1165
rlabel metal2 212 -684 212 -684 0 net=968
rlabel metal2 177 -686 177 -686 0 net=1217
rlabel metal2 219 -688 219 -688 0 net=835
rlabel metal2 177 -690 177 -690 0 net=1169
rlabel metal2 61 -701 61 -701 0 net=290
rlabel metal2 75 -701 75 -701 0 net=456
rlabel metal2 100 -701 100 -701 0 net=1006
rlabel metal2 121 -701 121 -701 0 net=560
rlabel metal2 184 -701 184 -701 0 net=1129
rlabel metal2 240 -701 240 -701 0 net=1218
rlabel metal2 114 -703 114 -703 0 net=751
rlabel metal2 128 -703 128 -703 0 net=598
rlabel metal2 142 -703 142 -703 0 net=532
rlabel metal2 194 -703 194 -703 0 net=1074
rlabel metal2 240 -703 240 -703 0 net=1247
rlabel metal2 131 -705 131 -705 0 net=789
rlabel metal2 149 -705 149 -705 0 net=1166
rlabel metal2 194 -705 194 -705 0 net=1170
rlabel metal2 247 -705 247 -705 0 net=1354
rlabel metal2 93 -707 93 -707 0 net=424
rlabel metal2 198 -707 198 -707 0 net=837
rlabel metal2 152 -709 152 -709 0 net=1142
rlabel metal2 163 -711 163 -711 0 net=806
rlabel metal2 205 -711 205 -711 0 net=1203
rlabel metal2 163 -713 163 -713 0 net=961
rlabel metal2 114 -724 114 -724 0 net=239
rlabel metal2 135 -724 135 -724 0 net=791
rlabel metal2 159 -724 159 -724 0 net=343
rlabel metal2 180 -724 180 -724 0 net=1130
rlabel metal2 191 -724 191 -724 0 net=1204
rlabel metal2 229 -724 229 -724 0 net=1248
rlabel metal2 121 -726 121 -726 0 net=752
rlabel metal2 163 -726 163 -726 0 net=963
rlabel metal2 173 -726 173 -726 0 net=838
rlabel metal2 117 -728 117 -728 0 net=1039
rlabel metal2 177 -728 177 -728 0 net=799
rlabel metal2 191 -728 191 -728 0 net=1177
rlabel metal2 128 -739 128 -739 0 net=792
rlabel metal2 149 -739 149 -739 0 net=1395
rlabel metal2 166 -739 166 -739 0 net=964
rlabel metal2 177 -739 177 -739 0 net=801
rlabel metal2 187 -739 187 -739 0 net=1178
rlabel metal2 121 -741 121 -741 0 net=1041
rlabel metal2 156 -741 156 -741 0 net=431
rlabel metal2 124 -752 124 -752 0 net=1042
rlabel metal2 156 -752 156 -752 0 net=432
rlabel metal2 184 -752 184 -752 0 net=802
rlabel metal2 159 -754 159 -754 0 net=1396
<< end >>
