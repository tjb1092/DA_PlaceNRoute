magic
tech scmos
timestamp 1555071782 
<< pdiffusion >>
rect 148 -12 154 -6
rect 204 -12 210 -6
rect 337 -12 343 -6
rect 344 -12 347 -6
rect 351 -12 354 -6
rect 358 -12 361 -6
rect 365 -12 368 -6
rect 372 -12 378 -6
rect 393 -12 396 -6
rect 400 -12 406 -6
rect 407 -12 413 -6
rect 428 -12 434 -6
rect 435 -12 441 -6
rect 449 -12 452 -6
rect 463 -12 466 -6
rect 470 -12 476 -6
rect 477 -12 483 -6
rect 491 -12 497 -6
rect 512 -12 515 -6
rect 575 -12 578 -6
rect 127 -43 130 -37
rect 197 -43 200 -37
rect 218 -43 221 -37
rect 239 -43 245 -37
rect 253 -43 256 -37
rect 281 -43 284 -37
rect 288 -43 294 -37
rect 295 -43 298 -37
rect 302 -43 305 -37
rect 309 -43 312 -37
rect 316 -43 322 -37
rect 323 -43 329 -37
rect 330 -43 333 -37
rect 337 -43 340 -37
rect 344 -43 347 -37
rect 351 -43 354 -37
rect 358 -43 361 -37
rect 365 -43 368 -37
rect 372 -43 378 -37
rect 379 -43 382 -37
rect 386 -43 389 -37
rect 393 -43 399 -37
rect 400 -43 403 -37
rect 407 -43 410 -37
rect 414 -43 417 -37
rect 421 -43 424 -37
rect 428 -43 434 -37
rect 435 -43 438 -37
rect 442 -43 448 -37
rect 449 -43 452 -37
rect 456 -43 459 -37
rect 463 -43 466 -37
rect 470 -43 473 -37
rect 477 -43 480 -37
rect 484 -43 487 -37
rect 491 -43 497 -37
rect 498 -43 504 -37
rect 505 -43 508 -37
rect 512 -43 515 -37
rect 526 -43 529 -37
rect 533 -43 539 -37
rect 540 -43 543 -37
rect 547 -43 550 -37
rect 589 -43 595 -37
rect 617 -43 620 -37
rect 624 -43 627 -37
rect 113 -96 119 -90
rect 141 -96 144 -90
rect 162 -96 165 -90
rect 169 -96 172 -90
rect 176 -96 179 -90
rect 183 -96 186 -90
rect 190 -96 193 -90
rect 197 -96 200 -90
rect 204 -96 207 -90
rect 211 -96 214 -90
rect 218 -96 221 -90
rect 225 -96 228 -90
rect 232 -96 235 -90
rect 239 -96 242 -90
rect 246 -96 249 -90
rect 253 -96 256 -90
rect 260 -96 263 -90
rect 267 -96 270 -90
rect 274 -96 280 -90
rect 281 -96 284 -90
rect 288 -96 291 -90
rect 295 -96 298 -90
rect 302 -96 305 -90
rect 309 -96 312 -90
rect 316 -96 319 -90
rect 323 -96 326 -90
rect 330 -96 336 -90
rect 337 -96 340 -90
rect 344 -96 350 -90
rect 351 -96 354 -90
rect 358 -96 361 -90
rect 365 -96 371 -90
rect 372 -96 378 -90
rect 379 -96 385 -90
rect 386 -96 392 -90
rect 393 -96 399 -90
rect 400 -96 403 -90
rect 407 -96 410 -90
rect 414 -96 417 -90
rect 421 -96 424 -90
rect 428 -96 431 -90
rect 435 -96 438 -90
rect 442 -96 445 -90
rect 449 -96 455 -90
rect 456 -96 459 -90
rect 463 -96 466 -90
rect 470 -96 476 -90
rect 477 -96 483 -90
rect 484 -96 487 -90
rect 491 -96 494 -90
rect 498 -96 501 -90
rect 505 -96 508 -90
rect 512 -96 515 -90
rect 519 -96 522 -90
rect 526 -96 529 -90
rect 533 -96 536 -90
rect 540 -96 543 -90
rect 547 -96 550 -90
rect 554 -96 557 -90
rect 561 -96 564 -90
rect 568 -96 571 -90
rect 575 -96 578 -90
rect 582 -96 585 -90
rect 589 -96 595 -90
rect 596 -96 599 -90
rect 603 -96 606 -90
rect 610 -96 613 -90
rect 617 -96 620 -90
rect 624 -96 627 -90
rect 631 -96 634 -90
rect 638 -96 641 -90
rect 645 -96 648 -90
rect 652 -96 655 -90
rect 659 -96 662 -90
rect 666 -96 669 -90
rect 673 -96 676 -90
rect 680 -96 683 -90
rect 687 -96 693 -90
rect 50 -163 53 -157
rect 57 -163 60 -157
rect 64 -163 67 -157
rect 71 -163 74 -157
rect 78 -163 84 -157
rect 85 -163 88 -157
rect 92 -163 95 -157
rect 99 -163 105 -157
rect 106 -163 109 -157
rect 113 -163 116 -157
rect 120 -163 123 -157
rect 127 -163 130 -157
rect 134 -163 137 -157
rect 141 -163 147 -157
rect 148 -163 154 -157
rect 155 -163 158 -157
rect 162 -163 165 -157
rect 169 -163 172 -157
rect 176 -163 179 -157
rect 183 -163 189 -157
rect 190 -163 196 -157
rect 197 -163 203 -157
rect 204 -163 207 -157
rect 211 -163 214 -157
rect 218 -163 221 -157
rect 225 -163 228 -157
rect 232 -163 235 -157
rect 239 -163 242 -157
rect 246 -163 249 -157
rect 253 -163 256 -157
rect 260 -163 263 -157
rect 267 -163 270 -157
rect 274 -163 277 -157
rect 281 -163 284 -157
rect 288 -163 291 -157
rect 295 -163 298 -157
rect 302 -163 305 -157
rect 309 -163 312 -157
rect 316 -163 319 -157
rect 323 -163 326 -157
rect 330 -163 333 -157
rect 337 -163 340 -157
rect 344 -163 347 -157
rect 351 -163 357 -157
rect 358 -163 361 -157
rect 365 -163 368 -157
rect 372 -163 375 -157
rect 379 -163 382 -157
rect 386 -163 389 -157
rect 393 -163 396 -157
rect 400 -163 403 -157
rect 407 -163 413 -157
rect 414 -163 420 -157
rect 421 -163 424 -157
rect 428 -163 431 -157
rect 435 -163 438 -157
rect 442 -163 445 -157
rect 449 -163 455 -157
rect 456 -163 459 -157
rect 463 -163 469 -157
rect 470 -163 476 -157
rect 477 -163 483 -157
rect 484 -163 487 -157
rect 491 -163 497 -157
rect 498 -163 501 -157
rect 505 -163 508 -157
rect 512 -163 515 -157
rect 519 -163 522 -157
rect 526 -163 529 -157
rect 533 -163 536 -157
rect 540 -163 543 -157
rect 547 -163 550 -157
rect 554 -163 557 -157
rect 561 -163 564 -157
rect 568 -163 571 -157
rect 575 -163 581 -157
rect 582 -163 585 -157
rect 589 -163 592 -157
rect 596 -163 599 -157
rect 603 -163 606 -157
rect 610 -163 613 -157
rect 617 -163 620 -157
rect 624 -163 627 -157
rect 631 -163 634 -157
rect 638 -163 641 -157
rect 645 -163 648 -157
rect 652 -163 655 -157
rect 659 -163 662 -157
rect 666 -163 669 -157
rect 673 -163 676 -157
rect 680 -163 683 -157
rect 687 -163 690 -157
rect 694 -163 697 -157
rect 701 -163 704 -157
rect 708 -163 711 -157
rect 715 -163 718 -157
rect 722 -163 725 -157
rect 729 -163 732 -157
rect 736 -163 739 -157
rect 743 -163 746 -157
rect 750 -163 753 -157
rect 757 -163 760 -157
rect 764 -163 767 -157
rect 771 -163 774 -157
rect 778 -163 781 -157
rect 785 -163 788 -157
rect 792 -163 795 -157
rect 799 -163 802 -157
rect 806 -163 809 -157
rect 813 -163 816 -157
rect 820 -163 823 -157
rect 43 -244 46 -238
rect 50 -244 53 -238
rect 57 -244 60 -238
rect 64 -244 67 -238
rect 71 -244 74 -238
rect 78 -244 81 -238
rect 85 -244 88 -238
rect 92 -244 95 -238
rect 99 -244 105 -238
rect 106 -244 109 -238
rect 113 -244 119 -238
rect 120 -244 126 -238
rect 127 -244 130 -238
rect 134 -244 140 -238
rect 141 -244 144 -238
rect 148 -244 151 -238
rect 155 -244 158 -238
rect 162 -244 168 -238
rect 169 -244 172 -238
rect 176 -244 179 -238
rect 183 -244 186 -238
rect 190 -244 193 -238
rect 197 -244 200 -238
rect 204 -244 207 -238
rect 211 -244 214 -238
rect 218 -244 221 -238
rect 225 -244 228 -238
rect 232 -244 235 -238
rect 239 -244 242 -238
rect 246 -244 249 -238
rect 253 -244 259 -238
rect 260 -244 263 -238
rect 267 -244 270 -238
rect 274 -244 277 -238
rect 281 -244 287 -238
rect 288 -244 294 -238
rect 295 -244 298 -238
rect 302 -244 305 -238
rect 309 -244 312 -238
rect 316 -244 319 -238
rect 323 -244 326 -238
rect 330 -244 333 -238
rect 337 -244 340 -238
rect 344 -244 350 -238
rect 351 -244 357 -238
rect 358 -244 364 -238
rect 365 -244 368 -238
rect 372 -244 378 -238
rect 379 -244 382 -238
rect 386 -244 389 -238
rect 393 -244 396 -238
rect 400 -244 406 -238
rect 407 -244 410 -238
rect 414 -244 417 -238
rect 421 -244 427 -238
rect 428 -244 431 -238
rect 435 -244 441 -238
rect 442 -244 445 -238
rect 449 -244 452 -238
rect 456 -244 462 -238
rect 463 -244 466 -238
rect 470 -244 476 -238
rect 477 -244 480 -238
rect 484 -244 487 -238
rect 491 -244 497 -238
rect 498 -244 501 -238
rect 505 -244 508 -238
rect 512 -244 515 -238
rect 519 -244 522 -238
rect 526 -244 529 -238
rect 533 -244 536 -238
rect 540 -244 543 -238
rect 547 -244 550 -238
rect 554 -244 557 -238
rect 561 -244 564 -238
rect 568 -244 571 -238
rect 575 -244 578 -238
rect 582 -244 585 -238
rect 589 -244 592 -238
rect 596 -244 599 -238
rect 603 -244 606 -238
rect 610 -244 613 -238
rect 617 -244 620 -238
rect 624 -244 627 -238
rect 631 -244 634 -238
rect 638 -244 641 -238
rect 645 -244 648 -238
rect 652 -244 655 -238
rect 659 -244 662 -238
rect 666 -244 669 -238
rect 673 -244 676 -238
rect 680 -244 683 -238
rect 687 -244 690 -238
rect 694 -244 697 -238
rect 701 -244 704 -238
rect 708 -244 711 -238
rect 715 -244 718 -238
rect 722 -244 725 -238
rect 729 -244 732 -238
rect 736 -244 739 -238
rect 743 -244 746 -238
rect 750 -244 753 -238
rect 757 -244 760 -238
rect 764 -244 767 -238
rect 771 -244 774 -238
rect 778 -244 781 -238
rect 785 -244 788 -238
rect 792 -244 795 -238
rect 799 -244 802 -238
rect 806 -244 809 -238
rect 813 -244 816 -238
rect 820 -244 823 -238
rect 827 -244 830 -238
rect 834 -244 837 -238
rect 841 -244 844 -238
rect 848 -244 851 -238
rect 855 -244 861 -238
rect 862 -244 865 -238
rect 1 -333 4 -327
rect 8 -333 11 -327
rect 15 -333 18 -327
rect 22 -333 25 -327
rect 29 -333 32 -327
rect 36 -333 39 -327
rect 43 -333 46 -327
rect 50 -333 53 -327
rect 57 -333 60 -327
rect 64 -333 70 -327
rect 71 -333 74 -327
rect 78 -333 81 -327
rect 85 -333 88 -327
rect 92 -333 95 -327
rect 99 -333 102 -327
rect 106 -333 109 -327
rect 113 -333 116 -327
rect 120 -333 123 -327
rect 127 -333 133 -327
rect 134 -333 137 -327
rect 141 -333 144 -327
rect 148 -333 151 -327
rect 155 -333 158 -327
rect 162 -333 165 -327
rect 169 -333 172 -327
rect 176 -333 179 -327
rect 183 -333 186 -327
rect 190 -333 196 -327
rect 197 -333 200 -327
rect 204 -333 207 -327
rect 211 -333 214 -327
rect 218 -333 221 -327
rect 225 -333 228 -327
rect 232 -333 235 -327
rect 239 -333 242 -327
rect 246 -333 249 -327
rect 253 -333 256 -327
rect 260 -333 263 -327
rect 267 -333 270 -327
rect 274 -333 277 -327
rect 281 -333 284 -327
rect 288 -333 291 -327
rect 295 -333 298 -327
rect 302 -333 308 -327
rect 309 -333 312 -327
rect 316 -333 319 -327
rect 323 -333 326 -327
rect 330 -333 333 -327
rect 337 -333 340 -327
rect 344 -333 347 -327
rect 351 -333 354 -327
rect 358 -333 361 -327
rect 365 -333 368 -327
rect 372 -333 378 -327
rect 379 -333 385 -327
rect 386 -333 389 -327
rect 393 -333 399 -327
rect 400 -333 406 -327
rect 407 -333 410 -327
rect 414 -333 420 -327
rect 421 -333 427 -327
rect 428 -333 431 -327
rect 435 -333 441 -327
rect 442 -333 448 -327
rect 449 -333 455 -327
rect 456 -333 462 -327
rect 463 -333 469 -327
rect 470 -333 476 -327
rect 477 -333 480 -327
rect 484 -333 490 -327
rect 491 -333 494 -327
rect 498 -333 501 -327
rect 505 -333 508 -327
rect 512 -333 515 -327
rect 519 -333 522 -327
rect 526 -333 529 -327
rect 533 -333 536 -327
rect 540 -333 543 -327
rect 547 -333 553 -327
rect 554 -333 557 -327
rect 561 -333 564 -327
rect 568 -333 574 -327
rect 575 -333 578 -327
rect 582 -333 585 -327
rect 589 -333 592 -327
rect 596 -333 599 -327
rect 603 -333 606 -327
rect 610 -333 613 -327
rect 617 -333 620 -327
rect 624 -333 627 -327
rect 631 -333 634 -327
rect 638 -333 641 -327
rect 645 -333 648 -327
rect 652 -333 655 -327
rect 659 -333 662 -327
rect 666 -333 669 -327
rect 673 -333 676 -327
rect 680 -333 683 -327
rect 687 -333 693 -327
rect 694 -333 697 -327
rect 701 -333 704 -327
rect 708 -333 711 -327
rect 715 -333 718 -327
rect 722 -333 725 -327
rect 729 -333 732 -327
rect 736 -333 739 -327
rect 743 -333 746 -327
rect 750 -333 753 -327
rect 757 -333 760 -327
rect 764 -333 767 -327
rect 771 -333 774 -327
rect 778 -333 781 -327
rect 785 -333 788 -327
rect 792 -333 795 -327
rect 799 -333 802 -327
rect 806 -333 809 -327
rect 813 -333 816 -327
rect 820 -333 823 -327
rect 827 -333 830 -327
rect 834 -333 837 -327
rect 841 -333 844 -327
rect 848 -333 851 -327
rect 855 -333 858 -327
rect 862 -333 865 -327
rect 869 -333 872 -327
rect 876 -333 879 -327
rect 883 -333 886 -327
rect 890 -333 893 -327
rect 897 -333 900 -327
rect 904 -333 907 -327
rect 911 -333 914 -327
rect 918 -333 921 -327
rect 925 -333 928 -327
rect 932 -333 935 -327
rect 939 -333 942 -327
rect 946 -333 949 -327
rect 953 -333 956 -327
rect 1 -420 4 -414
rect 8 -420 11 -414
rect 15 -420 18 -414
rect 22 -420 25 -414
rect 29 -420 32 -414
rect 36 -420 39 -414
rect 43 -420 46 -414
rect 50 -420 53 -414
rect 57 -420 60 -414
rect 64 -420 70 -414
rect 71 -420 77 -414
rect 78 -420 84 -414
rect 85 -420 91 -414
rect 92 -420 98 -414
rect 99 -420 102 -414
rect 106 -420 109 -414
rect 113 -420 116 -414
rect 120 -420 126 -414
rect 127 -420 130 -414
rect 134 -420 137 -414
rect 141 -420 144 -414
rect 148 -420 151 -414
rect 155 -420 161 -414
rect 162 -420 165 -414
rect 169 -420 172 -414
rect 176 -420 179 -414
rect 183 -420 189 -414
rect 190 -420 196 -414
rect 197 -420 200 -414
rect 204 -420 207 -414
rect 211 -420 214 -414
rect 218 -420 221 -414
rect 225 -420 228 -414
rect 232 -420 235 -414
rect 239 -420 245 -414
rect 246 -420 249 -414
rect 253 -420 256 -414
rect 260 -420 263 -414
rect 267 -420 270 -414
rect 274 -420 277 -414
rect 281 -420 284 -414
rect 288 -420 291 -414
rect 295 -420 298 -414
rect 302 -420 305 -414
rect 309 -420 312 -414
rect 316 -420 319 -414
rect 323 -420 326 -414
rect 330 -420 333 -414
rect 337 -420 340 -414
rect 344 -420 347 -414
rect 351 -420 357 -414
rect 358 -420 364 -414
rect 365 -420 368 -414
rect 372 -420 375 -414
rect 379 -420 382 -414
rect 386 -420 389 -414
rect 393 -420 399 -414
rect 400 -420 403 -414
rect 407 -420 413 -414
rect 414 -420 417 -414
rect 421 -420 424 -414
rect 428 -420 434 -414
rect 435 -420 438 -414
rect 442 -420 445 -414
rect 449 -420 452 -414
rect 456 -420 462 -414
rect 463 -420 469 -414
rect 470 -420 473 -414
rect 477 -420 480 -414
rect 484 -420 487 -414
rect 491 -420 494 -414
rect 498 -420 501 -414
rect 505 -420 508 -414
rect 512 -420 518 -414
rect 519 -420 522 -414
rect 526 -420 532 -414
rect 533 -420 536 -414
rect 540 -420 543 -414
rect 547 -420 553 -414
rect 554 -420 557 -414
rect 561 -420 564 -414
rect 568 -420 571 -414
rect 575 -420 578 -414
rect 582 -420 585 -414
rect 589 -420 592 -414
rect 596 -420 599 -414
rect 603 -420 606 -414
rect 610 -420 613 -414
rect 617 -420 623 -414
rect 624 -420 627 -414
rect 631 -420 634 -414
rect 638 -420 641 -414
rect 645 -420 648 -414
rect 652 -420 655 -414
rect 659 -420 662 -414
rect 666 -420 669 -414
rect 673 -420 676 -414
rect 680 -420 683 -414
rect 687 -420 690 -414
rect 694 -420 697 -414
rect 701 -420 704 -414
rect 708 -420 711 -414
rect 715 -420 718 -414
rect 722 -420 725 -414
rect 729 -420 732 -414
rect 736 -420 739 -414
rect 743 -420 746 -414
rect 750 -420 753 -414
rect 757 -420 760 -414
rect 764 -420 767 -414
rect 771 -420 774 -414
rect 778 -420 781 -414
rect 785 -420 788 -414
rect 792 -420 795 -414
rect 799 -420 802 -414
rect 806 -420 809 -414
rect 813 -420 816 -414
rect 820 -420 823 -414
rect 827 -420 830 -414
rect 834 -420 837 -414
rect 841 -420 844 -414
rect 848 -420 851 -414
rect 855 -420 858 -414
rect 862 -420 865 -414
rect 869 -420 872 -414
rect 876 -420 879 -414
rect 883 -420 886 -414
rect 890 -420 893 -414
rect 897 -420 900 -414
rect 904 -420 907 -414
rect 911 -420 914 -414
rect 918 -420 921 -414
rect 925 -420 928 -414
rect 932 -420 935 -414
rect 939 -420 942 -414
rect 946 -420 949 -414
rect 953 -420 956 -414
rect 960 -420 963 -414
rect 967 -420 970 -414
rect 974 -420 977 -414
rect 981 -420 984 -414
rect 988 -420 991 -414
rect 995 -420 998 -414
rect 1002 -420 1005 -414
rect 1023 -420 1026 -414
rect 1 -515 4 -509
rect 8 -515 11 -509
rect 15 -515 18 -509
rect 22 -515 25 -509
rect 29 -515 32 -509
rect 36 -515 39 -509
rect 43 -515 46 -509
rect 50 -515 53 -509
rect 57 -515 60 -509
rect 64 -515 67 -509
rect 71 -515 74 -509
rect 78 -515 81 -509
rect 85 -515 88 -509
rect 92 -515 98 -509
rect 99 -515 102 -509
rect 106 -515 109 -509
rect 113 -515 116 -509
rect 120 -515 123 -509
rect 127 -515 133 -509
rect 134 -515 140 -509
rect 141 -515 147 -509
rect 148 -515 154 -509
rect 155 -515 161 -509
rect 162 -515 165 -509
rect 169 -515 172 -509
rect 176 -515 179 -509
rect 183 -515 186 -509
rect 190 -515 193 -509
rect 197 -515 200 -509
rect 204 -515 207 -509
rect 211 -515 214 -509
rect 218 -515 221 -509
rect 225 -515 228 -509
rect 232 -515 235 -509
rect 239 -515 242 -509
rect 246 -515 252 -509
rect 253 -515 256 -509
rect 260 -515 263 -509
rect 267 -515 270 -509
rect 274 -515 277 -509
rect 281 -515 284 -509
rect 288 -515 291 -509
rect 295 -515 298 -509
rect 302 -515 305 -509
rect 309 -515 312 -509
rect 316 -515 319 -509
rect 323 -515 329 -509
rect 330 -515 333 -509
rect 337 -515 340 -509
rect 344 -515 347 -509
rect 351 -515 354 -509
rect 358 -515 361 -509
rect 365 -515 368 -509
rect 372 -515 375 -509
rect 379 -515 382 -509
rect 386 -515 392 -509
rect 393 -515 399 -509
rect 400 -515 403 -509
rect 407 -515 413 -509
rect 414 -515 417 -509
rect 421 -515 424 -509
rect 428 -515 431 -509
rect 435 -515 438 -509
rect 442 -515 448 -509
rect 449 -515 452 -509
rect 456 -515 459 -509
rect 463 -515 466 -509
rect 470 -515 473 -509
rect 477 -515 483 -509
rect 484 -515 487 -509
rect 491 -515 494 -509
rect 498 -515 501 -509
rect 505 -515 511 -509
rect 512 -515 515 -509
rect 519 -515 525 -509
rect 526 -515 529 -509
rect 533 -515 536 -509
rect 540 -515 543 -509
rect 547 -515 550 -509
rect 554 -515 557 -509
rect 561 -515 567 -509
rect 568 -515 574 -509
rect 575 -515 581 -509
rect 582 -515 585 -509
rect 589 -515 592 -509
rect 596 -515 599 -509
rect 603 -515 609 -509
rect 610 -515 613 -509
rect 617 -515 620 -509
rect 624 -515 627 -509
rect 631 -515 634 -509
rect 638 -515 641 -509
rect 645 -515 651 -509
rect 652 -515 655 -509
rect 659 -515 662 -509
rect 666 -515 672 -509
rect 673 -515 676 -509
rect 680 -515 683 -509
rect 687 -515 690 -509
rect 694 -515 697 -509
rect 701 -515 704 -509
rect 708 -515 711 -509
rect 715 -515 718 -509
rect 722 -515 725 -509
rect 729 -515 732 -509
rect 736 -515 739 -509
rect 743 -515 746 -509
rect 750 -515 756 -509
rect 757 -515 760 -509
rect 764 -515 767 -509
rect 771 -515 774 -509
rect 778 -515 781 -509
rect 785 -515 788 -509
rect 792 -515 795 -509
rect 799 -515 802 -509
rect 806 -515 809 -509
rect 813 -515 816 -509
rect 820 -515 823 -509
rect 827 -515 830 -509
rect 834 -515 837 -509
rect 841 -515 844 -509
rect 848 -515 851 -509
rect 855 -515 858 -509
rect 862 -515 865 -509
rect 869 -515 872 -509
rect 876 -515 879 -509
rect 883 -515 886 -509
rect 890 -515 893 -509
rect 897 -515 900 -509
rect 904 -515 907 -509
rect 911 -515 914 -509
rect 918 -515 921 -509
rect 925 -515 928 -509
rect 932 -515 935 -509
rect 939 -515 942 -509
rect 946 -515 949 -509
rect 953 -515 956 -509
rect 960 -515 963 -509
rect 967 -515 970 -509
rect 974 -515 977 -509
rect 981 -515 984 -509
rect 988 -515 991 -509
rect 995 -515 998 -509
rect 1002 -515 1005 -509
rect 1009 -515 1012 -509
rect 1016 -515 1019 -509
rect 1023 -515 1026 -509
rect 1030 -515 1033 -509
rect 1037 -515 1040 -509
rect 1044 -515 1047 -509
rect 1051 -515 1054 -509
rect 1058 -515 1061 -509
rect 1065 -515 1068 -509
rect 1072 -515 1075 -509
rect 1079 -515 1082 -509
rect 1086 -515 1089 -509
rect 1093 -515 1096 -509
rect 1100 -515 1103 -509
rect 1107 -515 1110 -509
rect 1114 -515 1117 -509
rect 1121 -515 1124 -509
rect 1 -614 4 -608
rect 8 -614 11 -608
rect 15 -614 18 -608
rect 22 -614 25 -608
rect 29 -614 32 -608
rect 36 -614 42 -608
rect 43 -614 46 -608
rect 50 -614 53 -608
rect 57 -614 63 -608
rect 64 -614 70 -608
rect 71 -614 77 -608
rect 78 -614 81 -608
rect 85 -614 88 -608
rect 92 -614 95 -608
rect 99 -614 102 -608
rect 106 -614 109 -608
rect 113 -614 116 -608
rect 120 -614 123 -608
rect 127 -614 130 -608
rect 134 -614 137 -608
rect 141 -614 147 -608
rect 148 -614 151 -608
rect 155 -614 158 -608
rect 162 -614 165 -608
rect 169 -614 172 -608
rect 176 -614 179 -608
rect 183 -614 189 -608
rect 190 -614 193 -608
rect 197 -614 200 -608
rect 204 -614 207 -608
rect 211 -614 214 -608
rect 218 -614 221 -608
rect 225 -614 228 -608
rect 232 -614 235 -608
rect 239 -614 242 -608
rect 246 -614 249 -608
rect 253 -614 256 -608
rect 260 -614 263 -608
rect 267 -614 270 -608
rect 274 -614 280 -608
rect 281 -614 284 -608
rect 288 -614 291 -608
rect 295 -614 298 -608
rect 302 -614 305 -608
rect 309 -614 312 -608
rect 316 -614 319 -608
rect 323 -614 326 -608
rect 330 -614 336 -608
rect 337 -614 340 -608
rect 344 -614 347 -608
rect 351 -614 354 -608
rect 358 -614 361 -608
rect 365 -614 368 -608
rect 372 -614 375 -608
rect 379 -614 385 -608
rect 386 -614 392 -608
rect 393 -614 396 -608
rect 400 -614 406 -608
rect 407 -614 410 -608
rect 414 -614 420 -608
rect 421 -614 427 -608
rect 428 -614 431 -608
rect 435 -614 438 -608
rect 442 -614 445 -608
rect 449 -614 455 -608
rect 456 -614 462 -608
rect 463 -614 469 -608
rect 470 -614 473 -608
rect 477 -614 480 -608
rect 484 -614 487 -608
rect 491 -614 494 -608
rect 498 -614 501 -608
rect 505 -614 508 -608
rect 512 -614 515 -608
rect 519 -614 525 -608
rect 526 -614 529 -608
rect 533 -614 536 -608
rect 540 -614 546 -608
rect 547 -614 553 -608
rect 554 -614 557 -608
rect 561 -614 567 -608
rect 568 -614 571 -608
rect 575 -614 578 -608
rect 582 -614 588 -608
rect 589 -614 592 -608
rect 596 -614 599 -608
rect 603 -614 606 -608
rect 610 -614 613 -608
rect 617 -614 623 -608
rect 624 -614 630 -608
rect 631 -614 634 -608
rect 638 -614 641 -608
rect 645 -614 648 -608
rect 652 -614 655 -608
rect 659 -614 662 -608
rect 666 -614 669 -608
rect 673 -614 676 -608
rect 680 -614 683 -608
rect 687 -614 690 -608
rect 694 -614 697 -608
rect 701 -614 704 -608
rect 708 -614 711 -608
rect 715 -614 718 -608
rect 722 -614 725 -608
rect 729 -614 732 -608
rect 736 -614 739 -608
rect 743 -614 746 -608
rect 750 -614 753 -608
rect 757 -614 760 -608
rect 764 -614 767 -608
rect 771 -614 774 -608
rect 778 -614 781 -608
rect 785 -614 788 -608
rect 792 -614 795 -608
rect 799 -614 802 -608
rect 806 -614 809 -608
rect 813 -614 816 -608
rect 820 -614 823 -608
rect 827 -614 830 -608
rect 834 -614 837 -608
rect 841 -614 844 -608
rect 848 -614 851 -608
rect 855 -614 858 -608
rect 862 -614 865 -608
rect 869 -614 872 -608
rect 876 -614 879 -608
rect 883 -614 886 -608
rect 890 -614 893 -608
rect 897 -614 900 -608
rect 904 -614 907 -608
rect 911 -614 914 -608
rect 918 -614 921 -608
rect 925 -614 928 -608
rect 932 -614 935 -608
rect 939 -614 942 -608
rect 946 -614 949 -608
rect 953 -614 956 -608
rect 960 -614 963 -608
rect 967 -614 970 -608
rect 974 -614 977 -608
rect 981 -614 984 -608
rect 988 -614 991 -608
rect 995 -614 998 -608
rect 1002 -614 1005 -608
rect 1009 -614 1012 -608
rect 1016 -614 1019 -608
rect 1023 -614 1026 -608
rect 1030 -614 1033 -608
rect 1037 -614 1040 -608
rect 1044 -614 1047 -608
rect 1051 -614 1054 -608
rect 1058 -614 1061 -608
rect 1065 -614 1068 -608
rect 1072 -614 1075 -608
rect 1079 -614 1085 -608
rect 1086 -614 1089 -608
rect 1 -723 4 -717
rect 8 -723 11 -717
rect 15 -723 18 -717
rect 22 -723 25 -717
rect 29 -723 32 -717
rect 36 -723 39 -717
rect 43 -723 49 -717
rect 50 -723 53 -717
rect 57 -723 63 -717
rect 64 -723 67 -717
rect 71 -723 74 -717
rect 78 -723 81 -717
rect 85 -723 91 -717
rect 92 -723 95 -717
rect 99 -723 102 -717
rect 106 -723 112 -717
rect 113 -723 116 -717
rect 120 -723 123 -717
rect 127 -723 130 -717
rect 134 -723 137 -717
rect 141 -723 144 -717
rect 148 -723 151 -717
rect 155 -723 158 -717
rect 162 -723 165 -717
rect 169 -723 172 -717
rect 176 -723 179 -717
rect 183 -723 186 -717
rect 190 -723 196 -717
rect 197 -723 200 -717
rect 204 -723 207 -717
rect 211 -723 214 -717
rect 218 -723 221 -717
rect 225 -723 231 -717
rect 232 -723 238 -717
rect 239 -723 242 -717
rect 246 -723 249 -717
rect 253 -723 256 -717
rect 260 -723 263 -717
rect 267 -723 270 -717
rect 274 -723 277 -717
rect 281 -723 284 -717
rect 288 -723 291 -717
rect 295 -723 298 -717
rect 302 -723 305 -717
rect 309 -723 312 -717
rect 316 -723 319 -717
rect 323 -723 326 -717
rect 330 -723 333 -717
rect 337 -723 340 -717
rect 344 -723 347 -717
rect 351 -723 354 -717
rect 358 -723 361 -717
rect 365 -723 371 -717
rect 372 -723 375 -717
rect 379 -723 385 -717
rect 386 -723 392 -717
rect 393 -723 396 -717
rect 400 -723 406 -717
rect 407 -723 410 -717
rect 414 -723 420 -717
rect 421 -723 424 -717
rect 428 -723 434 -717
rect 435 -723 438 -717
rect 442 -723 448 -717
rect 449 -723 452 -717
rect 456 -723 459 -717
rect 463 -723 466 -717
rect 470 -723 473 -717
rect 477 -723 480 -717
rect 484 -723 487 -717
rect 491 -723 494 -717
rect 498 -723 504 -717
rect 505 -723 508 -717
rect 512 -723 515 -717
rect 519 -723 522 -717
rect 526 -723 529 -717
rect 533 -723 536 -717
rect 540 -723 543 -717
rect 547 -723 550 -717
rect 554 -723 560 -717
rect 561 -723 567 -717
rect 568 -723 571 -717
rect 575 -723 578 -717
rect 582 -723 588 -717
rect 589 -723 592 -717
rect 596 -723 599 -717
rect 603 -723 606 -717
rect 610 -723 613 -717
rect 617 -723 620 -717
rect 624 -723 627 -717
rect 631 -723 637 -717
rect 638 -723 641 -717
rect 645 -723 651 -717
rect 652 -723 658 -717
rect 659 -723 662 -717
rect 666 -723 669 -717
rect 673 -723 676 -717
rect 680 -723 683 -717
rect 687 -723 690 -717
rect 694 -723 697 -717
rect 701 -723 704 -717
rect 708 -723 711 -717
rect 715 -723 718 -717
rect 722 -723 728 -717
rect 729 -723 735 -717
rect 736 -723 739 -717
rect 743 -723 746 -717
rect 750 -723 753 -717
rect 757 -723 760 -717
rect 764 -723 767 -717
rect 771 -723 774 -717
rect 778 -723 781 -717
rect 785 -723 788 -717
rect 792 -723 795 -717
rect 799 -723 802 -717
rect 806 -723 812 -717
rect 813 -723 816 -717
rect 820 -723 823 -717
rect 827 -723 830 -717
rect 834 -723 837 -717
rect 841 -723 844 -717
rect 848 -723 851 -717
rect 855 -723 858 -717
rect 862 -723 865 -717
rect 869 -723 872 -717
rect 876 -723 879 -717
rect 883 -723 886 -717
rect 890 -723 893 -717
rect 897 -723 900 -717
rect 904 -723 907 -717
rect 911 -723 914 -717
rect 918 -723 921 -717
rect 925 -723 928 -717
rect 932 -723 935 -717
rect 939 -723 942 -717
rect 946 -723 949 -717
rect 953 -723 956 -717
rect 960 -723 963 -717
rect 967 -723 970 -717
rect 974 -723 977 -717
rect 981 -723 984 -717
rect 988 -723 991 -717
rect 995 -723 998 -717
rect 1002 -723 1005 -717
rect 1009 -723 1012 -717
rect 1016 -723 1019 -717
rect 1023 -723 1026 -717
rect 1030 -723 1033 -717
rect 1037 -723 1040 -717
rect 1044 -723 1047 -717
rect 1051 -723 1054 -717
rect 1058 -723 1061 -717
rect 1065 -723 1068 -717
rect 1072 -723 1075 -717
rect 1079 -723 1082 -717
rect 1086 -723 1089 -717
rect 1093 -723 1096 -717
rect 1100 -723 1103 -717
rect 1107 -723 1110 -717
rect 1114 -723 1117 -717
rect 1121 -723 1124 -717
rect 1128 -723 1131 -717
rect 1135 -723 1138 -717
rect 1142 -723 1145 -717
rect 1149 -723 1152 -717
rect 1156 -723 1159 -717
rect 1163 -723 1166 -717
rect 1170 -723 1173 -717
rect 1177 -723 1180 -717
rect 1184 -723 1187 -717
rect 1191 -723 1194 -717
rect 1198 -723 1201 -717
rect 1205 -723 1208 -717
rect 1212 -723 1218 -717
rect 1359 -723 1362 -717
rect 1 -840 4 -834
rect 8 -840 11 -834
rect 15 -840 18 -834
rect 22 -840 28 -834
rect 29 -840 35 -834
rect 36 -840 39 -834
rect 43 -840 46 -834
rect 50 -840 53 -834
rect 57 -840 60 -834
rect 64 -840 67 -834
rect 71 -840 77 -834
rect 78 -840 81 -834
rect 85 -840 91 -834
rect 92 -840 95 -834
rect 99 -840 102 -834
rect 106 -840 109 -834
rect 113 -840 116 -834
rect 120 -840 123 -834
rect 127 -840 133 -834
rect 134 -840 137 -834
rect 141 -840 144 -834
rect 148 -840 151 -834
rect 155 -840 158 -834
rect 162 -840 165 -834
rect 169 -840 172 -834
rect 176 -840 182 -834
rect 183 -840 186 -834
rect 190 -840 193 -834
rect 197 -840 200 -834
rect 204 -840 207 -834
rect 211 -840 214 -834
rect 218 -840 221 -834
rect 225 -840 228 -834
rect 232 -840 235 -834
rect 239 -840 242 -834
rect 246 -840 249 -834
rect 253 -840 256 -834
rect 260 -840 263 -834
rect 267 -840 270 -834
rect 274 -840 277 -834
rect 281 -840 284 -834
rect 288 -840 291 -834
rect 295 -840 301 -834
rect 302 -840 305 -834
rect 309 -840 312 -834
rect 316 -840 319 -834
rect 323 -840 326 -834
rect 330 -840 333 -834
rect 337 -840 340 -834
rect 344 -840 347 -834
rect 351 -840 354 -834
rect 358 -840 361 -834
rect 365 -840 368 -834
rect 372 -840 375 -834
rect 379 -840 382 -834
rect 386 -840 392 -834
rect 393 -840 399 -834
rect 400 -840 406 -834
rect 407 -840 410 -834
rect 414 -840 417 -834
rect 421 -840 424 -834
rect 428 -840 434 -834
rect 435 -840 441 -834
rect 442 -840 445 -834
rect 449 -840 452 -834
rect 456 -840 459 -834
rect 463 -840 466 -834
rect 470 -840 473 -834
rect 477 -840 480 -834
rect 484 -840 487 -834
rect 491 -840 497 -834
rect 498 -840 501 -834
rect 505 -840 511 -834
rect 512 -840 518 -834
rect 519 -840 525 -834
rect 526 -840 529 -834
rect 533 -840 536 -834
rect 540 -840 543 -834
rect 547 -840 550 -834
rect 554 -840 557 -834
rect 561 -840 567 -834
rect 568 -840 574 -834
rect 575 -840 578 -834
rect 582 -840 588 -834
rect 589 -840 592 -834
rect 596 -840 599 -834
rect 603 -840 606 -834
rect 610 -840 613 -834
rect 617 -840 623 -834
rect 624 -840 627 -834
rect 631 -840 634 -834
rect 638 -840 641 -834
rect 645 -840 651 -834
rect 652 -840 658 -834
rect 659 -840 662 -834
rect 666 -840 669 -834
rect 673 -840 676 -834
rect 680 -840 683 -834
rect 687 -840 690 -834
rect 694 -840 697 -834
rect 701 -840 707 -834
rect 708 -840 711 -834
rect 715 -840 718 -834
rect 722 -840 725 -834
rect 729 -840 732 -834
rect 736 -840 739 -834
rect 743 -840 746 -834
rect 750 -840 753 -834
rect 757 -840 763 -834
rect 764 -840 767 -834
rect 771 -840 777 -834
rect 778 -840 781 -834
rect 785 -840 788 -834
rect 792 -840 795 -834
rect 799 -840 802 -834
rect 806 -840 809 -834
rect 813 -840 816 -834
rect 820 -840 823 -834
rect 827 -840 833 -834
rect 834 -840 837 -834
rect 841 -840 844 -834
rect 848 -840 851 -834
rect 855 -840 858 -834
rect 862 -840 865 -834
rect 869 -840 872 -834
rect 876 -840 879 -834
rect 883 -840 886 -834
rect 890 -840 893 -834
rect 897 -840 900 -834
rect 904 -840 907 -834
rect 911 -840 914 -834
rect 918 -840 921 -834
rect 925 -840 928 -834
rect 932 -840 935 -834
rect 939 -840 942 -834
rect 946 -840 949 -834
rect 953 -840 956 -834
rect 960 -840 963 -834
rect 967 -840 970 -834
rect 974 -840 977 -834
rect 981 -840 984 -834
rect 988 -840 991 -834
rect 995 -840 998 -834
rect 1002 -840 1005 -834
rect 1009 -840 1012 -834
rect 1016 -840 1019 -834
rect 1023 -840 1026 -834
rect 1030 -840 1033 -834
rect 1037 -840 1040 -834
rect 1044 -840 1047 -834
rect 1051 -840 1054 -834
rect 1058 -840 1061 -834
rect 1065 -840 1068 -834
rect 1072 -840 1075 -834
rect 1079 -840 1082 -834
rect 1086 -840 1089 -834
rect 1093 -840 1096 -834
rect 1100 -840 1103 -834
rect 1107 -840 1110 -834
rect 1114 -840 1117 -834
rect 1121 -840 1124 -834
rect 1128 -840 1131 -834
rect 1135 -840 1138 -834
rect 1142 -840 1145 -834
rect 1149 -840 1152 -834
rect 1156 -840 1159 -834
rect 1163 -840 1166 -834
rect 1170 -840 1173 -834
rect 1177 -840 1180 -834
rect 1184 -840 1187 -834
rect 1191 -840 1194 -834
rect 1198 -840 1201 -834
rect 1205 -840 1208 -834
rect 1212 -840 1215 -834
rect 1219 -840 1222 -834
rect 1226 -840 1229 -834
rect 1233 -840 1236 -834
rect 1240 -840 1243 -834
rect 1247 -840 1250 -834
rect 1254 -840 1257 -834
rect 1261 -840 1264 -834
rect 1415 -840 1418 -834
rect 1 -957 4 -951
rect 8 -957 11 -951
rect 15 -957 18 -951
rect 22 -957 25 -951
rect 29 -957 32 -951
rect 36 -957 39 -951
rect 43 -957 46 -951
rect 50 -957 53 -951
rect 57 -957 60 -951
rect 64 -957 70 -951
rect 71 -957 74 -951
rect 78 -957 81 -951
rect 85 -957 91 -951
rect 92 -957 95 -951
rect 99 -957 102 -951
rect 106 -957 109 -951
rect 113 -957 116 -951
rect 120 -957 126 -951
rect 127 -957 133 -951
rect 134 -957 137 -951
rect 141 -957 144 -951
rect 148 -957 154 -951
rect 155 -957 158 -951
rect 162 -957 165 -951
rect 169 -957 172 -951
rect 176 -957 179 -951
rect 183 -957 186 -951
rect 190 -957 193 -951
rect 197 -957 203 -951
rect 204 -957 207 -951
rect 211 -957 217 -951
rect 218 -957 221 -951
rect 225 -957 228 -951
rect 232 -957 235 -951
rect 239 -957 242 -951
rect 246 -957 249 -951
rect 253 -957 256 -951
rect 260 -957 263 -951
rect 267 -957 270 -951
rect 274 -957 277 -951
rect 281 -957 284 -951
rect 288 -957 291 -951
rect 295 -957 298 -951
rect 302 -957 305 -951
rect 309 -957 312 -951
rect 316 -957 322 -951
rect 323 -957 326 -951
rect 330 -957 333 -951
rect 337 -957 340 -951
rect 344 -957 347 -951
rect 351 -957 354 -951
rect 358 -957 361 -951
rect 365 -957 371 -951
rect 372 -957 375 -951
rect 379 -957 382 -951
rect 386 -957 389 -951
rect 393 -957 396 -951
rect 400 -957 403 -951
rect 407 -957 410 -951
rect 414 -957 417 -951
rect 421 -957 427 -951
rect 428 -957 431 -951
rect 435 -957 438 -951
rect 442 -957 445 -951
rect 449 -957 455 -951
rect 456 -957 459 -951
rect 463 -957 466 -951
rect 470 -957 473 -951
rect 477 -957 483 -951
rect 484 -957 487 -951
rect 491 -957 494 -951
rect 498 -957 504 -951
rect 505 -957 508 -951
rect 512 -957 515 -951
rect 519 -957 522 -951
rect 526 -957 532 -951
rect 533 -957 539 -951
rect 540 -957 546 -951
rect 547 -957 550 -951
rect 554 -957 557 -951
rect 561 -957 564 -951
rect 568 -957 571 -951
rect 575 -957 578 -951
rect 582 -957 585 -951
rect 589 -957 592 -951
rect 596 -957 599 -951
rect 603 -957 606 -951
rect 610 -957 616 -951
rect 617 -957 620 -951
rect 624 -957 630 -951
rect 631 -957 637 -951
rect 638 -957 641 -951
rect 645 -957 648 -951
rect 652 -957 658 -951
rect 659 -957 662 -951
rect 666 -957 669 -951
rect 673 -957 676 -951
rect 680 -957 683 -951
rect 687 -957 693 -951
rect 694 -957 697 -951
rect 701 -957 704 -951
rect 708 -957 714 -951
rect 715 -957 721 -951
rect 722 -957 725 -951
rect 729 -957 732 -951
rect 736 -957 739 -951
rect 743 -957 749 -951
rect 750 -957 753 -951
rect 757 -957 760 -951
rect 764 -957 767 -951
rect 771 -957 774 -951
rect 778 -957 781 -951
rect 785 -957 788 -951
rect 792 -957 795 -951
rect 799 -957 802 -951
rect 806 -957 809 -951
rect 813 -957 816 -951
rect 820 -957 826 -951
rect 827 -957 830 -951
rect 834 -957 837 -951
rect 841 -957 844 -951
rect 848 -957 851 -951
rect 855 -957 858 -951
rect 862 -957 865 -951
rect 869 -957 872 -951
rect 876 -957 879 -951
rect 883 -957 886 -951
rect 890 -957 893 -951
rect 897 -957 900 -951
rect 904 -957 907 -951
rect 911 -957 914 -951
rect 918 -957 921 -951
rect 925 -957 928 -951
rect 932 -957 935 -951
rect 939 -957 942 -951
rect 946 -957 949 -951
rect 953 -957 956 -951
rect 960 -957 963 -951
rect 967 -957 970 -951
rect 974 -957 977 -951
rect 981 -957 984 -951
rect 988 -957 991 -951
rect 995 -957 998 -951
rect 1002 -957 1005 -951
rect 1009 -957 1012 -951
rect 1016 -957 1019 -951
rect 1023 -957 1026 -951
rect 1030 -957 1033 -951
rect 1037 -957 1040 -951
rect 1044 -957 1047 -951
rect 1051 -957 1054 -951
rect 1058 -957 1061 -951
rect 1065 -957 1068 -951
rect 1072 -957 1075 -951
rect 1079 -957 1082 -951
rect 1086 -957 1089 -951
rect 1093 -957 1096 -951
rect 1100 -957 1103 -951
rect 1107 -957 1110 -951
rect 1114 -957 1117 -951
rect 1121 -957 1124 -951
rect 1128 -957 1131 -951
rect 1135 -957 1138 -951
rect 1142 -957 1145 -951
rect 1149 -957 1152 -951
rect 1156 -957 1159 -951
rect 1163 -957 1166 -951
rect 1170 -957 1173 -951
rect 1177 -957 1180 -951
rect 1184 -957 1187 -951
rect 1191 -957 1197 -951
rect 1198 -957 1204 -951
rect 1205 -957 1208 -951
rect 1436 -957 1439 -951
rect 1 -1086 7 -1080
rect 8 -1086 11 -1080
rect 15 -1086 18 -1080
rect 22 -1086 25 -1080
rect 29 -1086 35 -1080
rect 36 -1086 42 -1080
rect 43 -1086 46 -1080
rect 50 -1086 56 -1080
rect 57 -1086 60 -1080
rect 64 -1086 67 -1080
rect 71 -1086 77 -1080
rect 78 -1086 81 -1080
rect 85 -1086 88 -1080
rect 92 -1086 98 -1080
rect 99 -1086 105 -1080
rect 106 -1086 109 -1080
rect 113 -1086 116 -1080
rect 120 -1086 123 -1080
rect 127 -1086 130 -1080
rect 134 -1086 137 -1080
rect 141 -1086 144 -1080
rect 148 -1086 154 -1080
rect 155 -1086 158 -1080
rect 162 -1086 165 -1080
rect 169 -1086 172 -1080
rect 176 -1086 179 -1080
rect 183 -1086 186 -1080
rect 190 -1086 193 -1080
rect 197 -1086 200 -1080
rect 204 -1086 207 -1080
rect 211 -1086 214 -1080
rect 218 -1086 221 -1080
rect 225 -1086 228 -1080
rect 232 -1086 235 -1080
rect 239 -1086 242 -1080
rect 246 -1086 249 -1080
rect 253 -1086 256 -1080
rect 260 -1086 266 -1080
rect 267 -1086 270 -1080
rect 274 -1086 277 -1080
rect 281 -1086 284 -1080
rect 288 -1086 291 -1080
rect 295 -1086 298 -1080
rect 302 -1086 308 -1080
rect 309 -1086 312 -1080
rect 316 -1086 319 -1080
rect 323 -1086 326 -1080
rect 330 -1086 333 -1080
rect 337 -1086 343 -1080
rect 344 -1086 347 -1080
rect 351 -1086 354 -1080
rect 358 -1086 361 -1080
rect 365 -1086 368 -1080
rect 372 -1086 378 -1080
rect 379 -1086 382 -1080
rect 386 -1086 389 -1080
rect 393 -1086 396 -1080
rect 400 -1086 403 -1080
rect 407 -1086 410 -1080
rect 414 -1086 417 -1080
rect 421 -1086 424 -1080
rect 428 -1086 431 -1080
rect 435 -1086 441 -1080
rect 442 -1086 445 -1080
rect 449 -1086 452 -1080
rect 456 -1086 459 -1080
rect 463 -1086 466 -1080
rect 470 -1086 473 -1080
rect 477 -1086 483 -1080
rect 484 -1086 487 -1080
rect 491 -1086 497 -1080
rect 498 -1086 504 -1080
rect 505 -1086 508 -1080
rect 512 -1086 518 -1080
rect 519 -1086 522 -1080
rect 526 -1086 532 -1080
rect 533 -1086 536 -1080
rect 540 -1086 543 -1080
rect 547 -1086 550 -1080
rect 554 -1086 560 -1080
rect 561 -1086 567 -1080
rect 568 -1086 574 -1080
rect 575 -1086 578 -1080
rect 582 -1086 585 -1080
rect 589 -1086 592 -1080
rect 596 -1086 599 -1080
rect 603 -1086 606 -1080
rect 610 -1086 613 -1080
rect 617 -1086 620 -1080
rect 624 -1086 630 -1080
rect 631 -1086 637 -1080
rect 638 -1086 641 -1080
rect 645 -1086 648 -1080
rect 652 -1086 655 -1080
rect 659 -1086 662 -1080
rect 666 -1086 669 -1080
rect 673 -1086 679 -1080
rect 680 -1086 683 -1080
rect 687 -1086 690 -1080
rect 694 -1086 697 -1080
rect 701 -1086 704 -1080
rect 708 -1086 711 -1080
rect 715 -1086 718 -1080
rect 722 -1086 728 -1080
rect 729 -1086 732 -1080
rect 736 -1086 739 -1080
rect 743 -1086 749 -1080
rect 750 -1086 753 -1080
rect 757 -1086 760 -1080
rect 764 -1086 767 -1080
rect 771 -1086 774 -1080
rect 778 -1086 781 -1080
rect 785 -1086 788 -1080
rect 792 -1086 795 -1080
rect 799 -1086 802 -1080
rect 806 -1086 809 -1080
rect 813 -1086 816 -1080
rect 820 -1086 823 -1080
rect 827 -1086 830 -1080
rect 834 -1086 837 -1080
rect 841 -1086 844 -1080
rect 848 -1086 851 -1080
rect 855 -1086 858 -1080
rect 862 -1086 868 -1080
rect 869 -1086 872 -1080
rect 876 -1086 879 -1080
rect 883 -1086 886 -1080
rect 890 -1086 893 -1080
rect 897 -1086 900 -1080
rect 904 -1086 907 -1080
rect 911 -1086 914 -1080
rect 918 -1086 921 -1080
rect 925 -1086 931 -1080
rect 932 -1086 935 -1080
rect 939 -1086 942 -1080
rect 946 -1086 949 -1080
rect 953 -1086 956 -1080
rect 960 -1086 963 -1080
rect 967 -1086 970 -1080
rect 974 -1086 977 -1080
rect 981 -1086 984 -1080
rect 988 -1086 991 -1080
rect 995 -1086 998 -1080
rect 1002 -1086 1005 -1080
rect 1009 -1086 1012 -1080
rect 1016 -1086 1019 -1080
rect 1023 -1086 1026 -1080
rect 1030 -1086 1033 -1080
rect 1037 -1086 1040 -1080
rect 1044 -1086 1047 -1080
rect 1051 -1086 1054 -1080
rect 1058 -1086 1061 -1080
rect 1065 -1086 1068 -1080
rect 1072 -1086 1075 -1080
rect 1079 -1086 1082 -1080
rect 1086 -1086 1089 -1080
rect 1093 -1086 1096 -1080
rect 1100 -1086 1103 -1080
rect 1107 -1086 1110 -1080
rect 1114 -1086 1117 -1080
rect 1121 -1086 1124 -1080
rect 1128 -1086 1131 -1080
rect 1135 -1086 1138 -1080
rect 1142 -1086 1145 -1080
rect 1149 -1086 1152 -1080
rect 1156 -1086 1159 -1080
rect 1163 -1086 1166 -1080
rect 1170 -1086 1173 -1080
rect 1177 -1086 1180 -1080
rect 1184 -1086 1187 -1080
rect 1191 -1086 1194 -1080
rect 1198 -1086 1201 -1080
rect 1205 -1086 1208 -1080
rect 1212 -1086 1215 -1080
rect 1219 -1086 1222 -1080
rect 1226 -1086 1229 -1080
rect 1233 -1086 1236 -1080
rect 1240 -1086 1243 -1080
rect 1247 -1086 1250 -1080
rect 1254 -1086 1257 -1080
rect 1261 -1086 1264 -1080
rect 1268 -1086 1271 -1080
rect 1275 -1086 1278 -1080
rect 1282 -1086 1285 -1080
rect 1289 -1086 1292 -1080
rect 1296 -1086 1299 -1080
rect 1303 -1086 1306 -1080
rect 1310 -1086 1313 -1080
rect 1317 -1086 1320 -1080
rect 1324 -1086 1327 -1080
rect 1331 -1086 1334 -1080
rect 1338 -1086 1341 -1080
rect 1345 -1086 1348 -1080
rect 1443 -1086 1446 -1080
rect 1 -1211 7 -1205
rect 8 -1211 11 -1205
rect 15 -1211 18 -1205
rect 22 -1211 25 -1205
rect 29 -1211 32 -1205
rect 36 -1211 39 -1205
rect 43 -1211 46 -1205
rect 50 -1211 53 -1205
rect 57 -1211 60 -1205
rect 64 -1211 67 -1205
rect 71 -1211 77 -1205
rect 78 -1211 81 -1205
rect 85 -1211 88 -1205
rect 92 -1211 95 -1205
rect 99 -1211 105 -1205
rect 106 -1211 109 -1205
rect 113 -1211 119 -1205
rect 120 -1211 123 -1205
rect 127 -1211 130 -1205
rect 134 -1211 137 -1205
rect 141 -1211 144 -1205
rect 148 -1211 151 -1205
rect 155 -1211 158 -1205
rect 162 -1211 165 -1205
rect 169 -1211 172 -1205
rect 176 -1211 182 -1205
rect 183 -1211 186 -1205
rect 190 -1211 193 -1205
rect 197 -1211 200 -1205
rect 204 -1211 207 -1205
rect 211 -1211 217 -1205
rect 218 -1211 221 -1205
rect 225 -1211 228 -1205
rect 232 -1211 235 -1205
rect 239 -1211 242 -1205
rect 246 -1211 249 -1205
rect 253 -1211 256 -1205
rect 260 -1211 263 -1205
rect 267 -1211 270 -1205
rect 274 -1211 277 -1205
rect 281 -1211 284 -1205
rect 288 -1211 291 -1205
rect 295 -1211 298 -1205
rect 302 -1211 305 -1205
rect 309 -1211 312 -1205
rect 316 -1211 319 -1205
rect 323 -1211 326 -1205
rect 330 -1211 333 -1205
rect 337 -1211 340 -1205
rect 344 -1211 347 -1205
rect 351 -1211 354 -1205
rect 358 -1211 361 -1205
rect 365 -1211 368 -1205
rect 372 -1211 375 -1205
rect 379 -1211 382 -1205
rect 386 -1211 389 -1205
rect 393 -1211 396 -1205
rect 400 -1211 406 -1205
rect 407 -1211 410 -1205
rect 414 -1211 417 -1205
rect 421 -1211 424 -1205
rect 428 -1211 431 -1205
rect 435 -1211 438 -1205
rect 442 -1211 445 -1205
rect 449 -1211 452 -1205
rect 456 -1211 459 -1205
rect 463 -1211 469 -1205
rect 470 -1211 473 -1205
rect 477 -1211 480 -1205
rect 484 -1211 487 -1205
rect 491 -1211 497 -1205
rect 498 -1211 501 -1205
rect 505 -1211 508 -1205
rect 512 -1211 515 -1205
rect 519 -1211 525 -1205
rect 526 -1211 532 -1205
rect 533 -1211 536 -1205
rect 540 -1211 546 -1205
rect 547 -1211 553 -1205
rect 554 -1211 560 -1205
rect 561 -1211 564 -1205
rect 568 -1211 571 -1205
rect 575 -1211 578 -1205
rect 582 -1211 585 -1205
rect 589 -1211 592 -1205
rect 596 -1211 602 -1205
rect 603 -1211 609 -1205
rect 610 -1211 613 -1205
rect 617 -1211 620 -1205
rect 624 -1211 630 -1205
rect 631 -1211 637 -1205
rect 638 -1211 641 -1205
rect 645 -1211 651 -1205
rect 652 -1211 655 -1205
rect 659 -1211 662 -1205
rect 666 -1211 669 -1205
rect 673 -1211 676 -1205
rect 680 -1211 686 -1205
rect 687 -1211 690 -1205
rect 694 -1211 697 -1205
rect 701 -1211 704 -1205
rect 708 -1211 714 -1205
rect 715 -1211 718 -1205
rect 722 -1211 725 -1205
rect 729 -1211 735 -1205
rect 736 -1211 739 -1205
rect 743 -1211 749 -1205
rect 750 -1211 756 -1205
rect 757 -1211 763 -1205
rect 764 -1211 770 -1205
rect 771 -1211 774 -1205
rect 778 -1211 781 -1205
rect 785 -1211 788 -1205
rect 792 -1211 798 -1205
rect 799 -1211 802 -1205
rect 806 -1211 809 -1205
rect 813 -1211 816 -1205
rect 820 -1211 823 -1205
rect 827 -1211 830 -1205
rect 834 -1211 837 -1205
rect 841 -1211 847 -1205
rect 848 -1211 851 -1205
rect 855 -1211 858 -1205
rect 862 -1211 865 -1205
rect 869 -1211 872 -1205
rect 876 -1211 879 -1205
rect 883 -1211 886 -1205
rect 890 -1211 893 -1205
rect 897 -1211 900 -1205
rect 904 -1211 907 -1205
rect 911 -1211 914 -1205
rect 918 -1211 921 -1205
rect 925 -1211 928 -1205
rect 932 -1211 935 -1205
rect 939 -1211 942 -1205
rect 946 -1211 949 -1205
rect 953 -1211 956 -1205
rect 960 -1211 963 -1205
rect 967 -1211 970 -1205
rect 974 -1211 977 -1205
rect 981 -1211 984 -1205
rect 988 -1211 991 -1205
rect 995 -1211 998 -1205
rect 1002 -1211 1005 -1205
rect 1009 -1211 1012 -1205
rect 1016 -1211 1019 -1205
rect 1023 -1211 1026 -1205
rect 1030 -1211 1033 -1205
rect 1037 -1211 1040 -1205
rect 1044 -1211 1047 -1205
rect 1051 -1211 1054 -1205
rect 1058 -1211 1061 -1205
rect 1065 -1211 1068 -1205
rect 1072 -1211 1075 -1205
rect 1079 -1211 1082 -1205
rect 1086 -1211 1089 -1205
rect 1093 -1211 1096 -1205
rect 1100 -1211 1103 -1205
rect 1107 -1211 1110 -1205
rect 1114 -1211 1117 -1205
rect 1121 -1211 1124 -1205
rect 1128 -1211 1131 -1205
rect 1135 -1211 1138 -1205
rect 1142 -1211 1145 -1205
rect 1149 -1211 1152 -1205
rect 1156 -1211 1159 -1205
rect 1163 -1211 1166 -1205
rect 1170 -1211 1173 -1205
rect 1177 -1211 1180 -1205
rect 1184 -1211 1187 -1205
rect 1191 -1211 1194 -1205
rect 1198 -1211 1201 -1205
rect 1205 -1211 1208 -1205
rect 1212 -1211 1215 -1205
rect 1219 -1211 1222 -1205
rect 1226 -1211 1229 -1205
rect 1233 -1211 1236 -1205
rect 1240 -1211 1243 -1205
rect 1247 -1211 1250 -1205
rect 1254 -1211 1257 -1205
rect 1261 -1211 1264 -1205
rect 1268 -1211 1271 -1205
rect 1275 -1211 1278 -1205
rect 1282 -1211 1285 -1205
rect 1289 -1211 1292 -1205
rect 1296 -1211 1299 -1205
rect 1303 -1211 1306 -1205
rect 1310 -1211 1313 -1205
rect 1317 -1211 1320 -1205
rect 1324 -1211 1327 -1205
rect 1331 -1211 1334 -1205
rect 1338 -1211 1341 -1205
rect 1345 -1211 1348 -1205
rect 1352 -1211 1355 -1205
rect 1359 -1211 1362 -1205
rect 1366 -1211 1369 -1205
rect 1373 -1211 1376 -1205
rect 1450 -1211 1453 -1205
rect 1 -1332 4 -1326
rect 8 -1332 11 -1326
rect 15 -1332 18 -1326
rect 22 -1332 25 -1326
rect 29 -1332 32 -1326
rect 36 -1332 39 -1326
rect 43 -1332 46 -1326
rect 50 -1332 53 -1326
rect 57 -1332 63 -1326
rect 64 -1332 70 -1326
rect 71 -1332 74 -1326
rect 78 -1332 84 -1326
rect 85 -1332 91 -1326
rect 92 -1332 95 -1326
rect 99 -1332 102 -1326
rect 106 -1332 109 -1326
rect 113 -1332 116 -1326
rect 120 -1332 126 -1326
rect 127 -1332 130 -1326
rect 134 -1332 140 -1326
rect 141 -1332 144 -1326
rect 148 -1332 151 -1326
rect 155 -1332 158 -1326
rect 162 -1332 168 -1326
rect 169 -1332 175 -1326
rect 176 -1332 179 -1326
rect 183 -1332 186 -1326
rect 190 -1332 193 -1326
rect 197 -1332 200 -1326
rect 204 -1332 207 -1326
rect 211 -1332 214 -1326
rect 218 -1332 221 -1326
rect 225 -1332 228 -1326
rect 232 -1332 235 -1326
rect 239 -1332 242 -1326
rect 246 -1332 249 -1326
rect 253 -1332 256 -1326
rect 260 -1332 263 -1326
rect 267 -1332 270 -1326
rect 274 -1332 277 -1326
rect 281 -1332 284 -1326
rect 288 -1332 291 -1326
rect 295 -1332 298 -1326
rect 302 -1332 305 -1326
rect 309 -1332 312 -1326
rect 316 -1332 319 -1326
rect 323 -1332 326 -1326
rect 330 -1332 333 -1326
rect 337 -1332 340 -1326
rect 344 -1332 347 -1326
rect 351 -1332 354 -1326
rect 358 -1332 361 -1326
rect 365 -1332 371 -1326
rect 372 -1332 378 -1326
rect 379 -1332 382 -1326
rect 386 -1332 392 -1326
rect 393 -1332 396 -1326
rect 400 -1332 403 -1326
rect 407 -1332 410 -1326
rect 414 -1332 420 -1326
rect 421 -1332 424 -1326
rect 428 -1332 434 -1326
rect 435 -1332 438 -1326
rect 442 -1332 448 -1326
rect 449 -1332 452 -1326
rect 456 -1332 459 -1326
rect 463 -1332 466 -1326
rect 470 -1332 473 -1326
rect 477 -1332 480 -1326
rect 484 -1332 487 -1326
rect 491 -1332 494 -1326
rect 498 -1332 501 -1326
rect 505 -1332 508 -1326
rect 512 -1332 515 -1326
rect 519 -1332 522 -1326
rect 526 -1332 529 -1326
rect 533 -1332 536 -1326
rect 540 -1332 546 -1326
rect 547 -1332 550 -1326
rect 554 -1332 557 -1326
rect 561 -1332 564 -1326
rect 568 -1332 574 -1326
rect 575 -1332 578 -1326
rect 582 -1332 585 -1326
rect 589 -1332 592 -1326
rect 596 -1332 599 -1326
rect 603 -1332 606 -1326
rect 610 -1332 616 -1326
rect 617 -1332 623 -1326
rect 624 -1332 627 -1326
rect 631 -1332 637 -1326
rect 638 -1332 641 -1326
rect 645 -1332 648 -1326
rect 652 -1332 655 -1326
rect 659 -1332 662 -1326
rect 666 -1332 669 -1326
rect 673 -1332 676 -1326
rect 680 -1332 686 -1326
rect 687 -1332 690 -1326
rect 694 -1332 700 -1326
rect 701 -1332 707 -1326
rect 708 -1332 711 -1326
rect 715 -1332 721 -1326
rect 722 -1332 725 -1326
rect 729 -1332 735 -1326
rect 736 -1332 739 -1326
rect 743 -1332 746 -1326
rect 750 -1332 753 -1326
rect 757 -1332 760 -1326
rect 764 -1332 767 -1326
rect 771 -1332 774 -1326
rect 778 -1332 781 -1326
rect 785 -1332 788 -1326
rect 792 -1332 795 -1326
rect 799 -1332 802 -1326
rect 806 -1332 809 -1326
rect 813 -1332 819 -1326
rect 820 -1332 823 -1326
rect 827 -1332 830 -1326
rect 834 -1332 837 -1326
rect 841 -1332 844 -1326
rect 848 -1332 851 -1326
rect 855 -1332 858 -1326
rect 862 -1332 868 -1326
rect 869 -1332 872 -1326
rect 876 -1332 879 -1326
rect 883 -1332 886 -1326
rect 890 -1332 893 -1326
rect 897 -1332 903 -1326
rect 904 -1332 907 -1326
rect 911 -1332 917 -1326
rect 918 -1332 921 -1326
rect 925 -1332 928 -1326
rect 932 -1332 935 -1326
rect 939 -1332 942 -1326
rect 946 -1332 949 -1326
rect 953 -1332 956 -1326
rect 960 -1332 963 -1326
rect 967 -1332 970 -1326
rect 974 -1332 977 -1326
rect 981 -1332 984 -1326
rect 988 -1332 991 -1326
rect 995 -1332 998 -1326
rect 1002 -1332 1005 -1326
rect 1009 -1332 1012 -1326
rect 1016 -1332 1019 -1326
rect 1023 -1332 1026 -1326
rect 1030 -1332 1033 -1326
rect 1037 -1332 1040 -1326
rect 1044 -1332 1047 -1326
rect 1051 -1332 1054 -1326
rect 1058 -1332 1061 -1326
rect 1065 -1332 1068 -1326
rect 1072 -1332 1075 -1326
rect 1079 -1332 1082 -1326
rect 1086 -1332 1089 -1326
rect 1093 -1332 1096 -1326
rect 1100 -1332 1103 -1326
rect 1107 -1332 1110 -1326
rect 1114 -1332 1117 -1326
rect 1121 -1332 1124 -1326
rect 1128 -1332 1131 -1326
rect 1135 -1332 1138 -1326
rect 1142 -1332 1145 -1326
rect 1149 -1332 1152 -1326
rect 1156 -1332 1159 -1326
rect 1163 -1332 1166 -1326
rect 1170 -1332 1173 -1326
rect 1177 -1332 1180 -1326
rect 1184 -1332 1187 -1326
rect 1191 -1332 1194 -1326
rect 1198 -1332 1201 -1326
rect 1205 -1332 1208 -1326
rect 1212 -1332 1215 -1326
rect 1219 -1332 1222 -1326
rect 1226 -1332 1229 -1326
rect 1233 -1332 1236 -1326
rect 1240 -1332 1243 -1326
rect 1247 -1332 1250 -1326
rect 1254 -1332 1257 -1326
rect 1261 -1332 1264 -1326
rect 1268 -1332 1271 -1326
rect 1275 -1332 1278 -1326
rect 1282 -1332 1285 -1326
rect 1289 -1332 1292 -1326
rect 1296 -1332 1299 -1326
rect 1303 -1332 1306 -1326
rect 1310 -1332 1313 -1326
rect 1317 -1332 1320 -1326
rect 1324 -1332 1327 -1326
rect 1331 -1332 1334 -1326
rect 1338 -1332 1341 -1326
rect 1345 -1332 1348 -1326
rect 1352 -1332 1355 -1326
rect 1359 -1332 1362 -1326
rect 1366 -1332 1369 -1326
rect 1373 -1332 1376 -1326
rect 1380 -1332 1383 -1326
rect 1387 -1332 1390 -1326
rect 1457 -1332 1460 -1326
rect 1 -1457 4 -1451
rect 8 -1457 11 -1451
rect 15 -1457 18 -1451
rect 22 -1457 25 -1451
rect 29 -1457 35 -1451
rect 36 -1457 39 -1451
rect 43 -1457 46 -1451
rect 50 -1457 53 -1451
rect 57 -1457 60 -1451
rect 64 -1457 67 -1451
rect 71 -1457 74 -1451
rect 78 -1457 84 -1451
rect 85 -1457 88 -1451
rect 92 -1457 95 -1451
rect 99 -1457 102 -1451
rect 106 -1457 109 -1451
rect 113 -1457 116 -1451
rect 120 -1457 123 -1451
rect 127 -1457 133 -1451
rect 134 -1457 137 -1451
rect 141 -1457 144 -1451
rect 148 -1457 154 -1451
rect 155 -1457 158 -1451
rect 162 -1457 165 -1451
rect 169 -1457 172 -1451
rect 176 -1457 179 -1451
rect 183 -1457 186 -1451
rect 190 -1457 193 -1451
rect 197 -1457 200 -1451
rect 204 -1457 207 -1451
rect 211 -1457 214 -1451
rect 218 -1457 221 -1451
rect 225 -1457 228 -1451
rect 232 -1457 235 -1451
rect 239 -1457 242 -1451
rect 246 -1457 249 -1451
rect 253 -1457 256 -1451
rect 260 -1457 263 -1451
rect 267 -1457 270 -1451
rect 274 -1457 277 -1451
rect 281 -1457 284 -1451
rect 288 -1457 291 -1451
rect 295 -1457 298 -1451
rect 302 -1457 305 -1451
rect 309 -1457 312 -1451
rect 316 -1457 322 -1451
rect 323 -1457 326 -1451
rect 330 -1457 333 -1451
rect 337 -1457 340 -1451
rect 344 -1457 347 -1451
rect 351 -1457 354 -1451
rect 358 -1457 361 -1451
rect 365 -1457 368 -1451
rect 372 -1457 375 -1451
rect 379 -1457 382 -1451
rect 386 -1457 389 -1451
rect 393 -1457 399 -1451
rect 400 -1457 403 -1451
rect 407 -1457 413 -1451
rect 414 -1457 417 -1451
rect 421 -1457 424 -1451
rect 428 -1457 431 -1451
rect 435 -1457 438 -1451
rect 442 -1457 448 -1451
rect 449 -1457 452 -1451
rect 456 -1457 462 -1451
rect 463 -1457 466 -1451
rect 470 -1457 473 -1451
rect 477 -1457 480 -1451
rect 484 -1457 487 -1451
rect 491 -1457 494 -1451
rect 498 -1457 501 -1451
rect 505 -1457 511 -1451
rect 512 -1457 515 -1451
rect 519 -1457 525 -1451
rect 526 -1457 529 -1451
rect 533 -1457 539 -1451
rect 540 -1457 543 -1451
rect 547 -1457 553 -1451
rect 554 -1457 557 -1451
rect 561 -1457 567 -1451
rect 568 -1457 571 -1451
rect 575 -1457 578 -1451
rect 582 -1457 585 -1451
rect 589 -1457 592 -1451
rect 596 -1457 599 -1451
rect 603 -1457 606 -1451
rect 610 -1457 613 -1451
rect 617 -1457 620 -1451
rect 624 -1457 627 -1451
rect 631 -1457 634 -1451
rect 638 -1457 644 -1451
rect 645 -1457 651 -1451
rect 652 -1457 655 -1451
rect 659 -1457 662 -1451
rect 666 -1457 669 -1451
rect 673 -1457 676 -1451
rect 680 -1457 683 -1451
rect 687 -1457 690 -1451
rect 694 -1457 697 -1451
rect 701 -1457 704 -1451
rect 708 -1457 711 -1451
rect 715 -1457 718 -1451
rect 722 -1457 728 -1451
rect 729 -1457 732 -1451
rect 736 -1457 739 -1451
rect 743 -1457 749 -1451
rect 750 -1457 753 -1451
rect 757 -1457 760 -1451
rect 764 -1457 767 -1451
rect 771 -1457 774 -1451
rect 778 -1457 784 -1451
rect 785 -1457 788 -1451
rect 792 -1457 798 -1451
rect 799 -1457 802 -1451
rect 806 -1457 809 -1451
rect 813 -1457 819 -1451
rect 820 -1457 826 -1451
rect 827 -1457 833 -1451
rect 834 -1457 837 -1451
rect 841 -1457 844 -1451
rect 848 -1457 854 -1451
rect 855 -1457 861 -1451
rect 862 -1457 868 -1451
rect 869 -1457 872 -1451
rect 876 -1457 879 -1451
rect 883 -1457 889 -1451
rect 890 -1457 893 -1451
rect 897 -1457 900 -1451
rect 904 -1457 907 -1451
rect 911 -1457 914 -1451
rect 918 -1457 921 -1451
rect 925 -1457 928 -1451
rect 932 -1457 935 -1451
rect 939 -1457 942 -1451
rect 946 -1457 949 -1451
rect 953 -1457 956 -1451
rect 960 -1457 963 -1451
rect 967 -1457 970 -1451
rect 974 -1457 977 -1451
rect 981 -1457 984 -1451
rect 988 -1457 991 -1451
rect 995 -1457 998 -1451
rect 1002 -1457 1005 -1451
rect 1009 -1457 1012 -1451
rect 1016 -1457 1019 -1451
rect 1023 -1457 1026 -1451
rect 1030 -1457 1033 -1451
rect 1037 -1457 1040 -1451
rect 1044 -1457 1047 -1451
rect 1051 -1457 1054 -1451
rect 1058 -1457 1061 -1451
rect 1065 -1457 1068 -1451
rect 1072 -1457 1075 -1451
rect 1079 -1457 1082 -1451
rect 1086 -1457 1089 -1451
rect 1093 -1457 1096 -1451
rect 1100 -1457 1103 -1451
rect 1107 -1457 1110 -1451
rect 1114 -1457 1117 -1451
rect 1121 -1457 1124 -1451
rect 1128 -1457 1131 -1451
rect 1135 -1457 1138 -1451
rect 1142 -1457 1145 -1451
rect 1149 -1457 1152 -1451
rect 1156 -1457 1159 -1451
rect 1163 -1457 1166 -1451
rect 1170 -1457 1173 -1451
rect 1177 -1457 1180 -1451
rect 1184 -1457 1187 -1451
rect 1191 -1457 1194 -1451
rect 1198 -1457 1201 -1451
rect 1205 -1457 1208 -1451
rect 1212 -1457 1215 -1451
rect 1219 -1457 1222 -1451
rect 1226 -1457 1229 -1451
rect 1233 -1457 1236 -1451
rect 1240 -1457 1243 -1451
rect 1247 -1457 1250 -1451
rect 1254 -1457 1257 -1451
rect 1261 -1457 1264 -1451
rect 1268 -1457 1271 -1451
rect 1275 -1457 1278 -1451
rect 1282 -1457 1285 -1451
rect 1289 -1457 1292 -1451
rect 1296 -1457 1299 -1451
rect 1303 -1457 1306 -1451
rect 1310 -1457 1313 -1451
rect 1317 -1457 1320 -1451
rect 1324 -1457 1327 -1451
rect 1331 -1457 1334 -1451
rect 1338 -1457 1341 -1451
rect 1345 -1457 1348 -1451
rect 1352 -1457 1355 -1451
rect 1359 -1457 1362 -1451
rect 1366 -1457 1369 -1451
rect 1373 -1457 1376 -1451
rect 1380 -1457 1383 -1451
rect 1387 -1457 1390 -1451
rect 1394 -1457 1397 -1451
rect 1401 -1457 1404 -1451
rect 1408 -1457 1411 -1451
rect 1415 -1457 1418 -1451
rect 1422 -1457 1425 -1451
rect 1429 -1457 1432 -1451
rect 1436 -1457 1439 -1451
rect 1443 -1457 1446 -1451
rect 1450 -1457 1456 -1451
rect 1457 -1457 1460 -1451
rect 1464 -1457 1467 -1451
rect 1 -1594 4 -1588
rect 8 -1594 14 -1588
rect 15 -1594 21 -1588
rect 22 -1594 25 -1588
rect 29 -1594 32 -1588
rect 36 -1594 42 -1588
rect 43 -1594 46 -1588
rect 50 -1594 56 -1588
rect 57 -1594 60 -1588
rect 64 -1594 67 -1588
rect 71 -1594 74 -1588
rect 78 -1594 81 -1588
rect 85 -1594 91 -1588
rect 92 -1594 95 -1588
rect 99 -1594 105 -1588
rect 106 -1594 109 -1588
rect 113 -1594 119 -1588
rect 120 -1594 123 -1588
rect 127 -1594 130 -1588
rect 134 -1594 140 -1588
rect 141 -1594 147 -1588
rect 148 -1594 151 -1588
rect 155 -1594 158 -1588
rect 162 -1594 165 -1588
rect 169 -1594 172 -1588
rect 176 -1594 182 -1588
rect 183 -1594 186 -1588
rect 190 -1594 193 -1588
rect 197 -1594 200 -1588
rect 204 -1594 207 -1588
rect 211 -1594 214 -1588
rect 218 -1594 224 -1588
rect 225 -1594 228 -1588
rect 232 -1594 235 -1588
rect 239 -1594 242 -1588
rect 246 -1594 249 -1588
rect 253 -1594 256 -1588
rect 260 -1594 263 -1588
rect 267 -1594 270 -1588
rect 274 -1594 277 -1588
rect 281 -1594 284 -1588
rect 288 -1594 291 -1588
rect 295 -1594 298 -1588
rect 302 -1594 305 -1588
rect 309 -1594 312 -1588
rect 316 -1594 319 -1588
rect 323 -1594 326 -1588
rect 330 -1594 333 -1588
rect 337 -1594 340 -1588
rect 344 -1594 347 -1588
rect 351 -1594 354 -1588
rect 358 -1594 361 -1588
rect 365 -1594 368 -1588
rect 372 -1594 375 -1588
rect 379 -1594 382 -1588
rect 386 -1594 389 -1588
rect 393 -1594 396 -1588
rect 400 -1594 406 -1588
rect 407 -1594 410 -1588
rect 414 -1594 417 -1588
rect 421 -1594 424 -1588
rect 428 -1594 434 -1588
rect 435 -1594 438 -1588
rect 442 -1594 445 -1588
rect 449 -1594 452 -1588
rect 456 -1594 462 -1588
rect 463 -1594 466 -1588
rect 470 -1594 473 -1588
rect 477 -1594 480 -1588
rect 484 -1594 490 -1588
rect 491 -1594 497 -1588
rect 498 -1594 501 -1588
rect 505 -1594 508 -1588
rect 512 -1594 515 -1588
rect 519 -1594 525 -1588
rect 526 -1594 529 -1588
rect 533 -1594 539 -1588
rect 540 -1594 543 -1588
rect 547 -1594 550 -1588
rect 554 -1594 560 -1588
rect 561 -1594 564 -1588
rect 568 -1594 574 -1588
rect 575 -1594 578 -1588
rect 582 -1594 585 -1588
rect 589 -1594 592 -1588
rect 596 -1594 599 -1588
rect 603 -1594 606 -1588
rect 610 -1594 613 -1588
rect 617 -1594 623 -1588
rect 624 -1594 627 -1588
rect 631 -1594 634 -1588
rect 638 -1594 641 -1588
rect 645 -1594 648 -1588
rect 652 -1594 655 -1588
rect 659 -1594 665 -1588
rect 666 -1594 669 -1588
rect 673 -1594 676 -1588
rect 680 -1594 683 -1588
rect 687 -1594 690 -1588
rect 694 -1594 697 -1588
rect 701 -1594 707 -1588
rect 708 -1594 711 -1588
rect 715 -1594 718 -1588
rect 722 -1594 725 -1588
rect 729 -1594 732 -1588
rect 736 -1594 739 -1588
rect 743 -1594 746 -1588
rect 750 -1594 753 -1588
rect 757 -1594 760 -1588
rect 764 -1594 767 -1588
rect 771 -1594 774 -1588
rect 778 -1594 781 -1588
rect 785 -1594 788 -1588
rect 792 -1594 795 -1588
rect 799 -1594 805 -1588
rect 806 -1594 809 -1588
rect 813 -1594 816 -1588
rect 820 -1594 823 -1588
rect 827 -1594 833 -1588
rect 834 -1594 837 -1588
rect 841 -1594 844 -1588
rect 848 -1594 851 -1588
rect 855 -1594 861 -1588
rect 862 -1594 865 -1588
rect 869 -1594 872 -1588
rect 876 -1594 879 -1588
rect 883 -1594 886 -1588
rect 890 -1594 896 -1588
rect 897 -1594 900 -1588
rect 904 -1594 907 -1588
rect 911 -1594 914 -1588
rect 918 -1594 921 -1588
rect 925 -1594 928 -1588
rect 932 -1594 935 -1588
rect 939 -1594 942 -1588
rect 946 -1594 949 -1588
rect 953 -1594 956 -1588
rect 960 -1594 963 -1588
rect 967 -1594 970 -1588
rect 974 -1594 977 -1588
rect 981 -1594 984 -1588
rect 988 -1594 991 -1588
rect 995 -1594 998 -1588
rect 1002 -1594 1005 -1588
rect 1009 -1594 1012 -1588
rect 1016 -1594 1019 -1588
rect 1023 -1594 1026 -1588
rect 1030 -1594 1033 -1588
rect 1037 -1594 1040 -1588
rect 1044 -1594 1050 -1588
rect 1051 -1594 1054 -1588
rect 1058 -1594 1061 -1588
rect 1065 -1594 1068 -1588
rect 1072 -1594 1075 -1588
rect 1079 -1594 1082 -1588
rect 1086 -1594 1089 -1588
rect 1093 -1594 1096 -1588
rect 1100 -1594 1103 -1588
rect 1107 -1594 1110 -1588
rect 1114 -1594 1117 -1588
rect 1121 -1594 1124 -1588
rect 1128 -1594 1131 -1588
rect 1135 -1594 1138 -1588
rect 1142 -1594 1145 -1588
rect 1149 -1594 1152 -1588
rect 1156 -1594 1159 -1588
rect 1163 -1594 1166 -1588
rect 1170 -1594 1173 -1588
rect 1177 -1594 1180 -1588
rect 1184 -1594 1187 -1588
rect 1191 -1594 1194 -1588
rect 1198 -1594 1201 -1588
rect 1205 -1594 1208 -1588
rect 1212 -1594 1215 -1588
rect 1219 -1594 1222 -1588
rect 1226 -1594 1229 -1588
rect 1233 -1594 1236 -1588
rect 1240 -1594 1243 -1588
rect 1247 -1594 1250 -1588
rect 1254 -1594 1257 -1588
rect 1261 -1594 1264 -1588
rect 1268 -1594 1271 -1588
rect 1275 -1594 1278 -1588
rect 1282 -1594 1285 -1588
rect 1289 -1594 1292 -1588
rect 1296 -1594 1299 -1588
rect 1303 -1594 1306 -1588
rect 1310 -1594 1313 -1588
rect 1317 -1594 1320 -1588
rect 1324 -1594 1327 -1588
rect 1331 -1594 1334 -1588
rect 1338 -1594 1341 -1588
rect 1345 -1594 1348 -1588
rect 1352 -1594 1355 -1588
rect 1 -1725 4 -1719
rect 8 -1725 11 -1719
rect 15 -1725 21 -1719
rect 22 -1725 28 -1719
rect 29 -1725 35 -1719
rect 36 -1725 39 -1719
rect 43 -1725 49 -1719
rect 50 -1725 56 -1719
rect 57 -1725 60 -1719
rect 64 -1725 67 -1719
rect 71 -1725 74 -1719
rect 78 -1725 81 -1719
rect 85 -1725 88 -1719
rect 92 -1725 98 -1719
rect 99 -1725 102 -1719
rect 106 -1725 112 -1719
rect 113 -1725 116 -1719
rect 120 -1725 123 -1719
rect 127 -1725 130 -1719
rect 134 -1725 137 -1719
rect 141 -1725 144 -1719
rect 148 -1725 154 -1719
rect 155 -1725 161 -1719
rect 162 -1725 165 -1719
rect 169 -1725 172 -1719
rect 176 -1725 179 -1719
rect 183 -1725 186 -1719
rect 190 -1725 196 -1719
rect 197 -1725 200 -1719
rect 204 -1725 207 -1719
rect 211 -1725 214 -1719
rect 218 -1725 221 -1719
rect 225 -1725 228 -1719
rect 232 -1725 235 -1719
rect 239 -1725 242 -1719
rect 246 -1725 249 -1719
rect 253 -1725 256 -1719
rect 260 -1725 263 -1719
rect 267 -1725 270 -1719
rect 274 -1725 277 -1719
rect 281 -1725 284 -1719
rect 288 -1725 291 -1719
rect 295 -1725 298 -1719
rect 302 -1725 305 -1719
rect 309 -1725 312 -1719
rect 316 -1725 322 -1719
rect 323 -1725 326 -1719
rect 330 -1725 333 -1719
rect 337 -1725 340 -1719
rect 344 -1725 347 -1719
rect 351 -1725 354 -1719
rect 358 -1725 361 -1719
rect 365 -1725 368 -1719
rect 372 -1725 378 -1719
rect 379 -1725 382 -1719
rect 386 -1725 389 -1719
rect 393 -1725 396 -1719
rect 400 -1725 406 -1719
rect 407 -1725 410 -1719
rect 414 -1725 417 -1719
rect 421 -1725 424 -1719
rect 428 -1725 431 -1719
rect 435 -1725 438 -1719
rect 442 -1725 445 -1719
rect 449 -1725 452 -1719
rect 456 -1725 462 -1719
rect 463 -1725 466 -1719
rect 470 -1725 473 -1719
rect 477 -1725 480 -1719
rect 484 -1725 490 -1719
rect 491 -1725 494 -1719
rect 498 -1725 501 -1719
rect 505 -1725 508 -1719
rect 512 -1725 515 -1719
rect 519 -1725 525 -1719
rect 526 -1725 529 -1719
rect 533 -1725 536 -1719
rect 540 -1725 543 -1719
rect 547 -1725 553 -1719
rect 554 -1725 560 -1719
rect 561 -1725 564 -1719
rect 568 -1725 571 -1719
rect 575 -1725 578 -1719
rect 582 -1725 585 -1719
rect 589 -1725 592 -1719
rect 596 -1725 599 -1719
rect 603 -1725 606 -1719
rect 610 -1725 613 -1719
rect 617 -1725 620 -1719
rect 624 -1725 627 -1719
rect 631 -1725 634 -1719
rect 638 -1725 641 -1719
rect 645 -1725 648 -1719
rect 652 -1725 655 -1719
rect 659 -1725 662 -1719
rect 666 -1725 672 -1719
rect 673 -1725 676 -1719
rect 680 -1725 683 -1719
rect 687 -1725 690 -1719
rect 694 -1725 697 -1719
rect 701 -1725 704 -1719
rect 708 -1725 711 -1719
rect 715 -1725 718 -1719
rect 722 -1725 725 -1719
rect 729 -1725 732 -1719
rect 736 -1725 739 -1719
rect 743 -1725 749 -1719
rect 750 -1725 756 -1719
rect 757 -1725 760 -1719
rect 764 -1725 767 -1719
rect 771 -1725 777 -1719
rect 778 -1725 781 -1719
rect 785 -1725 788 -1719
rect 792 -1725 795 -1719
rect 799 -1725 802 -1719
rect 806 -1725 809 -1719
rect 813 -1725 816 -1719
rect 820 -1725 823 -1719
rect 827 -1725 830 -1719
rect 834 -1725 837 -1719
rect 841 -1725 844 -1719
rect 848 -1725 851 -1719
rect 855 -1725 858 -1719
rect 862 -1725 865 -1719
rect 869 -1725 872 -1719
rect 876 -1725 879 -1719
rect 883 -1725 886 -1719
rect 890 -1725 896 -1719
rect 897 -1725 903 -1719
rect 904 -1725 907 -1719
rect 911 -1725 914 -1719
rect 918 -1725 921 -1719
rect 925 -1725 928 -1719
rect 932 -1725 935 -1719
rect 939 -1725 945 -1719
rect 946 -1725 949 -1719
rect 953 -1725 956 -1719
rect 960 -1725 963 -1719
rect 967 -1725 970 -1719
rect 974 -1725 977 -1719
rect 981 -1725 984 -1719
rect 988 -1725 991 -1719
rect 995 -1725 998 -1719
rect 1002 -1725 1005 -1719
rect 1009 -1725 1012 -1719
rect 1016 -1725 1019 -1719
rect 1023 -1725 1026 -1719
rect 1030 -1725 1033 -1719
rect 1037 -1725 1040 -1719
rect 1044 -1725 1047 -1719
rect 1051 -1725 1054 -1719
rect 1058 -1725 1061 -1719
rect 1065 -1725 1071 -1719
rect 1072 -1725 1075 -1719
rect 1079 -1725 1082 -1719
rect 1086 -1725 1089 -1719
rect 1093 -1725 1096 -1719
rect 1100 -1725 1103 -1719
rect 1107 -1725 1110 -1719
rect 1114 -1725 1117 -1719
rect 1121 -1725 1127 -1719
rect 1128 -1725 1131 -1719
rect 1135 -1725 1138 -1719
rect 1142 -1725 1145 -1719
rect 1149 -1725 1152 -1719
rect 1156 -1725 1159 -1719
rect 1163 -1725 1166 -1719
rect 1170 -1725 1173 -1719
rect 1177 -1725 1180 -1719
rect 1184 -1725 1187 -1719
rect 1191 -1725 1194 -1719
rect 1198 -1725 1201 -1719
rect 1205 -1725 1208 -1719
rect 1212 -1725 1215 -1719
rect 1219 -1725 1222 -1719
rect 1226 -1725 1229 -1719
rect 1233 -1725 1236 -1719
rect 1240 -1725 1243 -1719
rect 1247 -1725 1250 -1719
rect 1254 -1725 1257 -1719
rect 1261 -1725 1264 -1719
rect 1268 -1725 1271 -1719
rect 1275 -1725 1278 -1719
rect 1282 -1725 1285 -1719
rect 1289 -1725 1292 -1719
rect 1296 -1725 1299 -1719
rect 1303 -1725 1306 -1719
rect 1310 -1725 1313 -1719
rect 1317 -1725 1320 -1719
rect 1324 -1725 1330 -1719
rect 1 -1844 4 -1838
rect 8 -1844 11 -1838
rect 15 -1844 18 -1838
rect 22 -1844 28 -1838
rect 29 -1844 32 -1838
rect 36 -1844 42 -1838
rect 43 -1844 49 -1838
rect 50 -1844 56 -1838
rect 57 -1844 60 -1838
rect 64 -1844 70 -1838
rect 71 -1844 74 -1838
rect 78 -1844 81 -1838
rect 85 -1844 88 -1838
rect 92 -1844 95 -1838
rect 99 -1844 102 -1838
rect 106 -1844 109 -1838
rect 113 -1844 119 -1838
rect 120 -1844 123 -1838
rect 127 -1844 130 -1838
rect 134 -1844 140 -1838
rect 141 -1844 144 -1838
rect 148 -1844 154 -1838
rect 155 -1844 158 -1838
rect 162 -1844 165 -1838
rect 169 -1844 172 -1838
rect 176 -1844 179 -1838
rect 183 -1844 186 -1838
rect 190 -1844 193 -1838
rect 197 -1844 200 -1838
rect 204 -1844 207 -1838
rect 211 -1844 214 -1838
rect 218 -1844 221 -1838
rect 225 -1844 228 -1838
rect 232 -1844 235 -1838
rect 239 -1844 242 -1838
rect 246 -1844 249 -1838
rect 253 -1844 256 -1838
rect 260 -1844 263 -1838
rect 267 -1844 270 -1838
rect 274 -1844 277 -1838
rect 281 -1844 284 -1838
rect 288 -1844 291 -1838
rect 295 -1844 301 -1838
rect 302 -1844 305 -1838
rect 309 -1844 312 -1838
rect 316 -1844 319 -1838
rect 323 -1844 326 -1838
rect 330 -1844 333 -1838
rect 337 -1844 340 -1838
rect 344 -1844 347 -1838
rect 351 -1844 357 -1838
rect 358 -1844 361 -1838
rect 365 -1844 371 -1838
rect 372 -1844 375 -1838
rect 379 -1844 382 -1838
rect 386 -1844 392 -1838
rect 393 -1844 396 -1838
rect 400 -1844 403 -1838
rect 407 -1844 410 -1838
rect 414 -1844 417 -1838
rect 421 -1844 424 -1838
rect 428 -1844 431 -1838
rect 435 -1844 438 -1838
rect 442 -1844 445 -1838
rect 449 -1844 452 -1838
rect 456 -1844 459 -1838
rect 463 -1844 469 -1838
rect 470 -1844 473 -1838
rect 477 -1844 483 -1838
rect 484 -1844 487 -1838
rect 491 -1844 494 -1838
rect 498 -1844 501 -1838
rect 505 -1844 508 -1838
rect 512 -1844 518 -1838
rect 519 -1844 522 -1838
rect 526 -1844 529 -1838
rect 533 -1844 536 -1838
rect 540 -1844 543 -1838
rect 547 -1844 550 -1838
rect 554 -1844 557 -1838
rect 561 -1844 564 -1838
rect 568 -1844 571 -1838
rect 575 -1844 578 -1838
rect 582 -1844 588 -1838
rect 589 -1844 592 -1838
rect 596 -1844 599 -1838
rect 603 -1844 609 -1838
rect 610 -1844 616 -1838
rect 617 -1844 620 -1838
rect 624 -1844 630 -1838
rect 631 -1844 634 -1838
rect 638 -1844 644 -1838
rect 645 -1844 648 -1838
rect 652 -1844 658 -1838
rect 659 -1844 662 -1838
rect 666 -1844 669 -1838
rect 673 -1844 676 -1838
rect 680 -1844 683 -1838
rect 687 -1844 690 -1838
rect 694 -1844 697 -1838
rect 701 -1844 704 -1838
rect 708 -1844 714 -1838
rect 715 -1844 721 -1838
rect 722 -1844 725 -1838
rect 729 -1844 735 -1838
rect 736 -1844 739 -1838
rect 743 -1844 746 -1838
rect 750 -1844 756 -1838
rect 757 -1844 763 -1838
rect 764 -1844 767 -1838
rect 771 -1844 774 -1838
rect 778 -1844 781 -1838
rect 785 -1844 788 -1838
rect 792 -1844 795 -1838
rect 799 -1844 802 -1838
rect 806 -1844 809 -1838
rect 813 -1844 816 -1838
rect 820 -1844 823 -1838
rect 827 -1844 830 -1838
rect 834 -1844 837 -1838
rect 841 -1844 844 -1838
rect 848 -1844 851 -1838
rect 855 -1844 858 -1838
rect 862 -1844 865 -1838
rect 869 -1844 872 -1838
rect 876 -1844 879 -1838
rect 883 -1844 886 -1838
rect 890 -1844 893 -1838
rect 897 -1844 900 -1838
rect 904 -1844 907 -1838
rect 911 -1844 914 -1838
rect 918 -1844 921 -1838
rect 925 -1844 928 -1838
rect 932 -1844 935 -1838
rect 939 -1844 942 -1838
rect 946 -1844 949 -1838
rect 953 -1844 956 -1838
rect 960 -1844 963 -1838
rect 967 -1844 970 -1838
rect 974 -1844 977 -1838
rect 981 -1844 984 -1838
rect 988 -1844 991 -1838
rect 995 -1844 998 -1838
rect 1002 -1844 1005 -1838
rect 1009 -1844 1012 -1838
rect 1016 -1844 1019 -1838
rect 1023 -1844 1026 -1838
rect 1030 -1844 1033 -1838
rect 1037 -1844 1040 -1838
rect 1044 -1844 1047 -1838
rect 1051 -1844 1054 -1838
rect 1058 -1844 1061 -1838
rect 1065 -1844 1068 -1838
rect 1072 -1844 1075 -1838
rect 1079 -1844 1082 -1838
rect 1086 -1844 1089 -1838
rect 1093 -1844 1096 -1838
rect 1100 -1844 1103 -1838
rect 1107 -1844 1110 -1838
rect 1114 -1844 1117 -1838
rect 1121 -1844 1124 -1838
rect 1128 -1844 1131 -1838
rect 1135 -1844 1138 -1838
rect 1142 -1844 1145 -1838
rect 1149 -1844 1152 -1838
rect 1156 -1844 1159 -1838
rect 1163 -1844 1166 -1838
rect 1170 -1844 1173 -1838
rect 1177 -1844 1180 -1838
rect 1184 -1844 1187 -1838
rect 1191 -1844 1194 -1838
rect 1198 -1844 1201 -1838
rect 1205 -1844 1208 -1838
rect 1212 -1844 1215 -1838
rect 1219 -1844 1222 -1838
rect 1226 -1844 1229 -1838
rect 1233 -1844 1236 -1838
rect 1240 -1844 1243 -1838
rect 1247 -1844 1250 -1838
rect 1254 -1844 1257 -1838
rect 1261 -1844 1264 -1838
rect 1268 -1844 1271 -1838
rect 1275 -1844 1278 -1838
rect 1282 -1844 1288 -1838
rect 8 -1967 11 -1961
rect 15 -1967 18 -1961
rect 22 -1967 25 -1961
rect 29 -1967 32 -1961
rect 36 -1967 39 -1961
rect 43 -1967 46 -1961
rect 50 -1967 56 -1961
rect 57 -1967 60 -1961
rect 64 -1967 70 -1961
rect 71 -1967 74 -1961
rect 78 -1967 81 -1961
rect 85 -1967 91 -1961
rect 92 -1967 98 -1961
rect 99 -1967 105 -1961
rect 106 -1967 109 -1961
rect 113 -1967 116 -1961
rect 120 -1967 123 -1961
rect 127 -1967 130 -1961
rect 134 -1967 140 -1961
rect 141 -1967 144 -1961
rect 148 -1967 151 -1961
rect 155 -1967 158 -1961
rect 162 -1967 165 -1961
rect 169 -1967 175 -1961
rect 176 -1967 179 -1961
rect 183 -1967 186 -1961
rect 190 -1967 193 -1961
rect 197 -1967 200 -1961
rect 204 -1967 207 -1961
rect 211 -1967 214 -1961
rect 218 -1967 221 -1961
rect 225 -1967 228 -1961
rect 232 -1967 235 -1961
rect 239 -1967 242 -1961
rect 246 -1967 249 -1961
rect 253 -1967 256 -1961
rect 260 -1967 266 -1961
rect 267 -1967 270 -1961
rect 274 -1967 277 -1961
rect 281 -1967 287 -1961
rect 288 -1967 291 -1961
rect 295 -1967 298 -1961
rect 302 -1967 305 -1961
rect 309 -1967 312 -1961
rect 316 -1967 322 -1961
rect 323 -1967 326 -1961
rect 330 -1967 333 -1961
rect 337 -1967 340 -1961
rect 344 -1967 347 -1961
rect 351 -1967 354 -1961
rect 358 -1967 361 -1961
rect 365 -1967 371 -1961
rect 372 -1967 375 -1961
rect 379 -1967 382 -1961
rect 386 -1967 389 -1961
rect 393 -1967 396 -1961
rect 400 -1967 403 -1961
rect 407 -1967 410 -1961
rect 414 -1967 417 -1961
rect 421 -1967 424 -1961
rect 428 -1967 434 -1961
rect 435 -1967 438 -1961
rect 442 -1967 445 -1961
rect 449 -1967 452 -1961
rect 456 -1967 462 -1961
rect 463 -1967 466 -1961
rect 470 -1967 473 -1961
rect 477 -1967 480 -1961
rect 484 -1967 487 -1961
rect 491 -1967 497 -1961
rect 498 -1967 501 -1961
rect 505 -1967 508 -1961
rect 512 -1967 515 -1961
rect 519 -1967 525 -1961
rect 526 -1967 529 -1961
rect 533 -1967 536 -1961
rect 540 -1967 543 -1961
rect 547 -1967 550 -1961
rect 554 -1967 560 -1961
rect 561 -1967 564 -1961
rect 568 -1967 574 -1961
rect 575 -1967 578 -1961
rect 582 -1967 585 -1961
rect 589 -1967 592 -1961
rect 596 -1967 599 -1961
rect 603 -1967 609 -1961
rect 610 -1967 613 -1961
rect 617 -1967 620 -1961
rect 624 -1967 627 -1961
rect 631 -1967 634 -1961
rect 638 -1967 641 -1961
rect 645 -1967 648 -1961
rect 652 -1967 655 -1961
rect 659 -1967 662 -1961
rect 666 -1967 669 -1961
rect 673 -1967 679 -1961
rect 680 -1967 683 -1961
rect 687 -1967 690 -1961
rect 694 -1967 697 -1961
rect 701 -1967 707 -1961
rect 708 -1967 711 -1961
rect 715 -1967 718 -1961
rect 722 -1967 725 -1961
rect 729 -1967 732 -1961
rect 736 -1967 739 -1961
rect 743 -1967 746 -1961
rect 750 -1967 753 -1961
rect 757 -1967 763 -1961
rect 764 -1967 767 -1961
rect 771 -1967 774 -1961
rect 778 -1967 781 -1961
rect 785 -1967 788 -1961
rect 792 -1967 795 -1961
rect 799 -1967 802 -1961
rect 806 -1967 809 -1961
rect 813 -1967 816 -1961
rect 820 -1967 823 -1961
rect 827 -1967 830 -1961
rect 834 -1967 840 -1961
rect 841 -1967 844 -1961
rect 848 -1967 851 -1961
rect 855 -1967 858 -1961
rect 862 -1967 865 -1961
rect 869 -1967 872 -1961
rect 876 -1967 879 -1961
rect 883 -1967 886 -1961
rect 890 -1967 893 -1961
rect 897 -1967 900 -1961
rect 904 -1967 907 -1961
rect 911 -1967 914 -1961
rect 918 -1967 924 -1961
rect 925 -1967 928 -1961
rect 932 -1967 935 -1961
rect 939 -1967 942 -1961
rect 946 -1967 949 -1961
rect 953 -1967 956 -1961
rect 960 -1967 966 -1961
rect 967 -1967 970 -1961
rect 974 -1967 977 -1961
rect 981 -1967 984 -1961
rect 988 -1967 991 -1961
rect 995 -1967 998 -1961
rect 1002 -1967 1005 -1961
rect 1009 -1967 1012 -1961
rect 1016 -1967 1019 -1961
rect 1023 -1967 1026 -1961
rect 1030 -1967 1033 -1961
rect 1037 -1967 1040 -1961
rect 1044 -1967 1047 -1961
rect 1051 -1967 1054 -1961
rect 1058 -1967 1061 -1961
rect 1065 -1967 1068 -1961
rect 1072 -1967 1075 -1961
rect 1079 -1967 1082 -1961
rect 1086 -1967 1089 -1961
rect 1093 -1967 1096 -1961
rect 1100 -1967 1103 -1961
rect 1107 -1967 1110 -1961
rect 1114 -1967 1117 -1961
rect 1121 -1967 1124 -1961
rect 1128 -1967 1131 -1961
rect 1135 -1967 1138 -1961
rect 1142 -1967 1145 -1961
rect 1149 -1967 1152 -1961
rect 1156 -1967 1159 -1961
rect 1163 -1967 1166 -1961
rect 1170 -1967 1173 -1961
rect 1177 -1967 1180 -1961
rect 1184 -1967 1187 -1961
rect 1191 -1967 1194 -1961
rect 1198 -1967 1201 -1961
rect 1205 -1967 1208 -1961
rect 1212 -1967 1215 -1961
rect 1219 -1967 1225 -1961
rect 1226 -1967 1229 -1961
rect 1233 -1967 1236 -1961
rect 1 -2070 4 -2064
rect 8 -2070 11 -2064
rect 15 -2070 18 -2064
rect 22 -2070 25 -2064
rect 29 -2070 32 -2064
rect 36 -2070 39 -2064
rect 43 -2070 46 -2064
rect 50 -2070 53 -2064
rect 57 -2070 60 -2064
rect 64 -2070 67 -2064
rect 71 -2070 74 -2064
rect 78 -2070 81 -2064
rect 85 -2070 91 -2064
rect 92 -2070 98 -2064
rect 99 -2070 102 -2064
rect 106 -2070 112 -2064
rect 113 -2070 119 -2064
rect 120 -2070 123 -2064
rect 127 -2070 130 -2064
rect 134 -2070 137 -2064
rect 141 -2070 144 -2064
rect 148 -2070 154 -2064
rect 155 -2070 158 -2064
rect 162 -2070 168 -2064
rect 169 -2070 172 -2064
rect 176 -2070 179 -2064
rect 183 -2070 186 -2064
rect 190 -2070 193 -2064
rect 197 -2070 200 -2064
rect 204 -2070 207 -2064
rect 211 -2070 214 -2064
rect 218 -2070 221 -2064
rect 225 -2070 228 -2064
rect 232 -2070 235 -2064
rect 239 -2070 245 -2064
rect 246 -2070 249 -2064
rect 253 -2070 256 -2064
rect 260 -2070 263 -2064
rect 267 -2070 270 -2064
rect 274 -2070 280 -2064
rect 281 -2070 284 -2064
rect 288 -2070 291 -2064
rect 295 -2070 298 -2064
rect 302 -2070 305 -2064
rect 309 -2070 312 -2064
rect 316 -2070 319 -2064
rect 323 -2070 329 -2064
rect 330 -2070 336 -2064
rect 337 -2070 340 -2064
rect 344 -2070 347 -2064
rect 351 -2070 354 -2064
rect 358 -2070 361 -2064
rect 365 -2070 368 -2064
rect 372 -2070 375 -2064
rect 379 -2070 382 -2064
rect 386 -2070 389 -2064
rect 393 -2070 396 -2064
rect 400 -2070 403 -2064
rect 407 -2070 413 -2064
rect 414 -2070 417 -2064
rect 421 -2070 424 -2064
rect 428 -2070 431 -2064
rect 435 -2070 438 -2064
rect 442 -2070 445 -2064
rect 449 -2070 452 -2064
rect 456 -2070 459 -2064
rect 463 -2070 466 -2064
rect 470 -2070 473 -2064
rect 477 -2070 483 -2064
rect 484 -2070 490 -2064
rect 491 -2070 494 -2064
rect 498 -2070 504 -2064
rect 505 -2070 508 -2064
rect 512 -2070 515 -2064
rect 519 -2070 522 -2064
rect 526 -2070 529 -2064
rect 533 -2070 536 -2064
rect 540 -2070 543 -2064
rect 547 -2070 550 -2064
rect 554 -2070 557 -2064
rect 561 -2070 564 -2064
rect 568 -2070 571 -2064
rect 575 -2070 581 -2064
rect 582 -2070 588 -2064
rect 589 -2070 592 -2064
rect 596 -2070 599 -2064
rect 603 -2070 606 -2064
rect 610 -2070 613 -2064
rect 617 -2070 623 -2064
rect 624 -2070 627 -2064
rect 631 -2070 634 -2064
rect 638 -2070 641 -2064
rect 645 -2070 648 -2064
rect 652 -2070 658 -2064
rect 659 -2070 665 -2064
rect 666 -2070 669 -2064
rect 673 -2070 676 -2064
rect 680 -2070 683 -2064
rect 687 -2070 690 -2064
rect 694 -2070 700 -2064
rect 701 -2070 704 -2064
rect 708 -2070 711 -2064
rect 715 -2070 718 -2064
rect 722 -2070 725 -2064
rect 729 -2070 732 -2064
rect 736 -2070 739 -2064
rect 743 -2070 746 -2064
rect 750 -2070 753 -2064
rect 757 -2070 760 -2064
rect 764 -2070 767 -2064
rect 771 -2070 774 -2064
rect 778 -2070 781 -2064
rect 785 -2070 788 -2064
rect 792 -2070 795 -2064
rect 799 -2070 802 -2064
rect 806 -2070 809 -2064
rect 813 -2070 819 -2064
rect 820 -2070 823 -2064
rect 827 -2070 830 -2064
rect 834 -2070 837 -2064
rect 841 -2070 844 -2064
rect 848 -2070 851 -2064
rect 855 -2070 858 -2064
rect 862 -2070 868 -2064
rect 869 -2070 872 -2064
rect 876 -2070 879 -2064
rect 883 -2070 886 -2064
rect 890 -2070 893 -2064
rect 897 -2070 900 -2064
rect 904 -2070 907 -2064
rect 911 -2070 914 -2064
rect 918 -2070 921 -2064
rect 925 -2070 928 -2064
rect 932 -2070 935 -2064
rect 939 -2070 942 -2064
rect 946 -2070 949 -2064
rect 953 -2070 956 -2064
rect 960 -2070 963 -2064
rect 967 -2070 970 -2064
rect 974 -2070 977 -2064
rect 981 -2070 984 -2064
rect 988 -2070 991 -2064
rect 995 -2070 998 -2064
rect 1002 -2070 1005 -2064
rect 1009 -2070 1012 -2064
rect 1016 -2070 1019 -2064
rect 1023 -2070 1029 -2064
rect 1030 -2070 1033 -2064
rect 1037 -2070 1040 -2064
rect 1044 -2070 1047 -2064
rect 1051 -2070 1054 -2064
rect 1058 -2070 1061 -2064
rect 1065 -2070 1068 -2064
rect 1072 -2070 1075 -2064
rect 1079 -2070 1082 -2064
rect 1086 -2070 1089 -2064
rect 1093 -2070 1096 -2064
rect 1100 -2070 1103 -2064
rect 1107 -2070 1110 -2064
rect 1114 -2070 1117 -2064
rect 1121 -2070 1124 -2064
rect 1128 -2070 1131 -2064
rect 1135 -2070 1141 -2064
rect 1142 -2070 1145 -2064
rect 1149 -2070 1152 -2064
rect 1156 -2070 1159 -2064
rect 1184 -2070 1187 -2064
rect 22 -2155 25 -2149
rect 29 -2155 32 -2149
rect 36 -2155 39 -2149
rect 43 -2155 46 -2149
rect 50 -2155 53 -2149
rect 57 -2155 60 -2149
rect 64 -2155 67 -2149
rect 71 -2155 74 -2149
rect 78 -2155 81 -2149
rect 85 -2155 88 -2149
rect 92 -2155 98 -2149
rect 99 -2155 105 -2149
rect 106 -2155 109 -2149
rect 113 -2155 119 -2149
rect 120 -2155 123 -2149
rect 127 -2155 130 -2149
rect 134 -2155 140 -2149
rect 141 -2155 144 -2149
rect 148 -2155 151 -2149
rect 155 -2155 158 -2149
rect 162 -2155 165 -2149
rect 169 -2155 175 -2149
rect 176 -2155 179 -2149
rect 183 -2155 186 -2149
rect 190 -2155 193 -2149
rect 197 -2155 200 -2149
rect 204 -2155 207 -2149
rect 211 -2155 214 -2149
rect 218 -2155 221 -2149
rect 225 -2155 228 -2149
rect 232 -2155 235 -2149
rect 239 -2155 242 -2149
rect 246 -2155 249 -2149
rect 253 -2155 256 -2149
rect 260 -2155 263 -2149
rect 267 -2155 270 -2149
rect 274 -2155 277 -2149
rect 281 -2155 284 -2149
rect 288 -2155 291 -2149
rect 295 -2155 301 -2149
rect 302 -2155 305 -2149
rect 309 -2155 312 -2149
rect 316 -2155 322 -2149
rect 323 -2155 326 -2149
rect 330 -2155 333 -2149
rect 337 -2155 340 -2149
rect 344 -2155 347 -2149
rect 351 -2155 354 -2149
rect 358 -2155 361 -2149
rect 365 -2155 368 -2149
rect 372 -2155 375 -2149
rect 379 -2155 382 -2149
rect 386 -2155 389 -2149
rect 393 -2155 396 -2149
rect 400 -2155 403 -2149
rect 407 -2155 410 -2149
rect 414 -2155 417 -2149
rect 421 -2155 424 -2149
rect 428 -2155 431 -2149
rect 435 -2155 438 -2149
rect 442 -2155 445 -2149
rect 449 -2155 452 -2149
rect 456 -2155 459 -2149
rect 463 -2155 469 -2149
rect 470 -2155 473 -2149
rect 477 -2155 483 -2149
rect 484 -2155 490 -2149
rect 491 -2155 494 -2149
rect 498 -2155 501 -2149
rect 505 -2155 511 -2149
rect 512 -2155 518 -2149
rect 519 -2155 522 -2149
rect 526 -2155 532 -2149
rect 533 -2155 536 -2149
rect 540 -2155 543 -2149
rect 547 -2155 550 -2149
rect 554 -2155 557 -2149
rect 561 -2155 564 -2149
rect 568 -2155 571 -2149
rect 575 -2155 578 -2149
rect 582 -2155 585 -2149
rect 589 -2155 592 -2149
rect 596 -2155 602 -2149
rect 603 -2155 606 -2149
rect 610 -2155 616 -2149
rect 617 -2155 620 -2149
rect 624 -2155 627 -2149
rect 631 -2155 634 -2149
rect 638 -2155 644 -2149
rect 645 -2155 648 -2149
rect 652 -2155 658 -2149
rect 659 -2155 662 -2149
rect 666 -2155 669 -2149
rect 673 -2155 676 -2149
rect 680 -2155 683 -2149
rect 687 -2155 693 -2149
rect 694 -2155 697 -2149
rect 701 -2155 704 -2149
rect 708 -2155 711 -2149
rect 715 -2155 718 -2149
rect 722 -2155 725 -2149
rect 729 -2155 732 -2149
rect 736 -2155 739 -2149
rect 743 -2155 746 -2149
rect 750 -2155 753 -2149
rect 757 -2155 760 -2149
rect 764 -2155 767 -2149
rect 771 -2155 774 -2149
rect 778 -2155 781 -2149
rect 785 -2155 791 -2149
rect 792 -2155 795 -2149
rect 799 -2155 802 -2149
rect 806 -2155 809 -2149
rect 813 -2155 816 -2149
rect 820 -2155 823 -2149
rect 827 -2155 830 -2149
rect 834 -2155 837 -2149
rect 841 -2155 844 -2149
rect 848 -2155 851 -2149
rect 855 -2155 858 -2149
rect 862 -2155 865 -2149
rect 869 -2155 872 -2149
rect 876 -2155 879 -2149
rect 883 -2155 886 -2149
rect 890 -2155 893 -2149
rect 897 -2155 900 -2149
rect 904 -2155 907 -2149
rect 911 -2155 914 -2149
rect 918 -2155 921 -2149
rect 925 -2155 928 -2149
rect 932 -2155 935 -2149
rect 939 -2155 942 -2149
rect 946 -2155 949 -2149
rect 953 -2155 956 -2149
rect 960 -2155 963 -2149
rect 967 -2155 973 -2149
rect 974 -2155 977 -2149
rect 981 -2155 984 -2149
rect 988 -2155 991 -2149
rect 995 -2155 1001 -2149
rect 1002 -2155 1005 -2149
rect 1009 -2155 1012 -2149
rect 1016 -2155 1019 -2149
rect 1023 -2155 1026 -2149
rect 1030 -2155 1033 -2149
rect 1037 -2155 1040 -2149
rect 1044 -2155 1047 -2149
rect 1051 -2155 1054 -2149
rect 1058 -2155 1061 -2149
rect 1065 -2155 1068 -2149
rect 1100 -2155 1106 -2149
rect 1107 -2155 1110 -2149
rect 1121 -2155 1124 -2149
rect 29 -2236 32 -2230
rect 36 -2236 39 -2230
rect 43 -2236 46 -2230
rect 50 -2236 53 -2230
rect 57 -2236 60 -2230
rect 64 -2236 67 -2230
rect 71 -2236 74 -2230
rect 78 -2236 84 -2230
rect 85 -2236 91 -2230
rect 92 -2236 98 -2230
rect 99 -2236 102 -2230
rect 106 -2236 109 -2230
rect 113 -2236 116 -2230
rect 120 -2236 126 -2230
rect 127 -2236 133 -2230
rect 134 -2236 137 -2230
rect 141 -2236 144 -2230
rect 148 -2236 151 -2230
rect 155 -2236 158 -2230
rect 162 -2236 165 -2230
rect 169 -2236 172 -2230
rect 176 -2236 182 -2230
rect 183 -2236 186 -2230
rect 190 -2236 193 -2230
rect 197 -2236 200 -2230
rect 204 -2236 207 -2230
rect 211 -2236 214 -2230
rect 218 -2236 221 -2230
rect 225 -2236 228 -2230
rect 232 -2236 235 -2230
rect 239 -2236 242 -2230
rect 246 -2236 249 -2230
rect 253 -2236 256 -2230
rect 260 -2236 263 -2230
rect 267 -2236 270 -2230
rect 274 -2236 277 -2230
rect 281 -2236 284 -2230
rect 288 -2236 291 -2230
rect 295 -2236 298 -2230
rect 302 -2236 305 -2230
rect 309 -2236 312 -2230
rect 316 -2236 319 -2230
rect 323 -2236 326 -2230
rect 330 -2236 333 -2230
rect 337 -2236 340 -2230
rect 344 -2236 347 -2230
rect 351 -2236 357 -2230
rect 358 -2236 361 -2230
rect 365 -2236 368 -2230
rect 372 -2236 375 -2230
rect 379 -2236 382 -2230
rect 386 -2236 389 -2230
rect 393 -2236 399 -2230
rect 400 -2236 403 -2230
rect 407 -2236 410 -2230
rect 414 -2236 417 -2230
rect 421 -2236 424 -2230
rect 428 -2236 431 -2230
rect 435 -2236 438 -2230
rect 442 -2236 448 -2230
rect 449 -2236 455 -2230
rect 456 -2236 459 -2230
rect 463 -2236 466 -2230
rect 470 -2236 473 -2230
rect 477 -2236 483 -2230
rect 484 -2236 490 -2230
rect 491 -2236 494 -2230
rect 498 -2236 501 -2230
rect 505 -2236 508 -2230
rect 512 -2236 515 -2230
rect 519 -2236 522 -2230
rect 526 -2236 532 -2230
rect 533 -2236 536 -2230
rect 540 -2236 543 -2230
rect 547 -2236 550 -2230
rect 554 -2236 557 -2230
rect 561 -2236 564 -2230
rect 568 -2236 571 -2230
rect 575 -2236 578 -2230
rect 582 -2236 585 -2230
rect 589 -2236 592 -2230
rect 596 -2236 599 -2230
rect 603 -2236 606 -2230
rect 610 -2236 613 -2230
rect 617 -2236 620 -2230
rect 624 -2236 627 -2230
rect 631 -2236 634 -2230
rect 638 -2236 641 -2230
rect 645 -2236 648 -2230
rect 652 -2236 658 -2230
rect 659 -2236 662 -2230
rect 666 -2236 672 -2230
rect 673 -2236 676 -2230
rect 680 -2236 683 -2230
rect 687 -2236 690 -2230
rect 694 -2236 700 -2230
rect 701 -2236 704 -2230
rect 708 -2236 711 -2230
rect 715 -2236 718 -2230
rect 722 -2236 725 -2230
rect 729 -2236 732 -2230
rect 736 -2236 742 -2230
rect 743 -2236 749 -2230
rect 750 -2236 753 -2230
rect 757 -2236 760 -2230
rect 764 -2236 767 -2230
rect 771 -2236 774 -2230
rect 778 -2236 781 -2230
rect 785 -2236 788 -2230
rect 792 -2236 795 -2230
rect 799 -2236 802 -2230
rect 806 -2236 809 -2230
rect 813 -2236 816 -2230
rect 820 -2236 823 -2230
rect 827 -2236 830 -2230
rect 834 -2236 837 -2230
rect 841 -2236 844 -2230
rect 848 -2236 851 -2230
rect 855 -2236 858 -2230
rect 862 -2236 865 -2230
rect 869 -2236 872 -2230
rect 876 -2236 879 -2230
rect 883 -2236 886 -2230
rect 890 -2236 893 -2230
rect 897 -2236 900 -2230
rect 904 -2236 907 -2230
rect 911 -2236 914 -2230
rect 918 -2236 921 -2230
rect 925 -2236 928 -2230
rect 932 -2236 935 -2230
rect 939 -2236 945 -2230
rect 946 -2236 949 -2230
rect 953 -2236 959 -2230
rect 960 -2236 963 -2230
rect 967 -2236 970 -2230
rect 974 -2236 977 -2230
rect 981 -2236 984 -2230
rect 995 -2236 998 -2230
rect 1002 -2236 1005 -2230
rect 1016 -2236 1019 -2230
rect 1065 -2236 1068 -2230
rect 43 -2319 46 -2313
rect 50 -2319 53 -2313
rect 57 -2319 60 -2313
rect 64 -2319 67 -2313
rect 71 -2319 74 -2313
rect 78 -2319 81 -2313
rect 85 -2319 91 -2313
rect 92 -2319 95 -2313
rect 99 -2319 102 -2313
rect 106 -2319 109 -2313
rect 113 -2319 116 -2313
rect 120 -2319 123 -2313
rect 127 -2319 130 -2313
rect 134 -2319 140 -2313
rect 141 -2319 144 -2313
rect 148 -2319 151 -2313
rect 155 -2319 158 -2313
rect 162 -2319 165 -2313
rect 169 -2319 172 -2313
rect 176 -2319 179 -2313
rect 183 -2319 189 -2313
rect 190 -2319 193 -2313
rect 197 -2319 200 -2313
rect 204 -2319 207 -2313
rect 211 -2319 214 -2313
rect 218 -2319 221 -2313
rect 225 -2319 228 -2313
rect 232 -2319 235 -2313
rect 239 -2319 242 -2313
rect 246 -2319 249 -2313
rect 253 -2319 256 -2313
rect 260 -2319 263 -2313
rect 267 -2319 270 -2313
rect 274 -2319 277 -2313
rect 281 -2319 284 -2313
rect 288 -2319 294 -2313
rect 295 -2319 298 -2313
rect 302 -2319 305 -2313
rect 309 -2319 312 -2313
rect 316 -2319 319 -2313
rect 323 -2319 326 -2313
rect 330 -2319 333 -2313
rect 337 -2319 340 -2313
rect 344 -2319 350 -2313
rect 351 -2319 354 -2313
rect 358 -2319 361 -2313
rect 365 -2319 368 -2313
rect 372 -2319 378 -2313
rect 379 -2319 382 -2313
rect 386 -2319 389 -2313
rect 393 -2319 396 -2313
rect 400 -2319 403 -2313
rect 407 -2319 410 -2313
rect 414 -2319 417 -2313
rect 421 -2319 427 -2313
rect 428 -2319 431 -2313
rect 435 -2319 438 -2313
rect 442 -2319 448 -2313
rect 449 -2319 455 -2313
rect 456 -2319 459 -2313
rect 463 -2319 466 -2313
rect 470 -2319 473 -2313
rect 477 -2319 480 -2313
rect 484 -2319 487 -2313
rect 491 -2319 497 -2313
rect 498 -2319 501 -2313
rect 505 -2319 508 -2313
rect 512 -2319 515 -2313
rect 519 -2319 522 -2313
rect 526 -2319 529 -2313
rect 533 -2319 539 -2313
rect 540 -2319 543 -2313
rect 547 -2319 550 -2313
rect 554 -2319 557 -2313
rect 561 -2319 567 -2313
rect 568 -2319 574 -2313
rect 575 -2319 581 -2313
rect 582 -2319 585 -2313
rect 589 -2319 592 -2313
rect 596 -2319 599 -2313
rect 603 -2319 606 -2313
rect 610 -2319 613 -2313
rect 617 -2319 623 -2313
rect 624 -2319 627 -2313
rect 631 -2319 634 -2313
rect 638 -2319 641 -2313
rect 645 -2319 648 -2313
rect 652 -2319 658 -2313
rect 659 -2319 662 -2313
rect 666 -2319 669 -2313
rect 673 -2319 676 -2313
rect 680 -2319 683 -2313
rect 687 -2319 690 -2313
rect 694 -2319 697 -2313
rect 701 -2319 704 -2313
rect 708 -2319 711 -2313
rect 715 -2319 718 -2313
rect 722 -2319 725 -2313
rect 729 -2319 732 -2313
rect 736 -2319 739 -2313
rect 743 -2319 746 -2313
rect 750 -2319 753 -2313
rect 757 -2319 760 -2313
rect 764 -2319 767 -2313
rect 771 -2319 774 -2313
rect 778 -2319 781 -2313
rect 785 -2319 788 -2313
rect 792 -2319 795 -2313
rect 799 -2319 805 -2313
rect 806 -2319 809 -2313
rect 813 -2319 816 -2313
rect 820 -2319 823 -2313
rect 827 -2319 830 -2313
rect 834 -2319 837 -2313
rect 841 -2319 844 -2313
rect 848 -2319 851 -2313
rect 855 -2319 858 -2313
rect 862 -2319 865 -2313
rect 869 -2319 872 -2313
rect 876 -2319 879 -2313
rect 883 -2319 886 -2313
rect 890 -2319 893 -2313
rect 897 -2319 900 -2313
rect 967 -2319 970 -2313
rect 988 -2319 991 -2313
rect 995 -2319 998 -2313
rect 1037 -2319 1040 -2313
rect 1058 -2319 1064 -2313
rect 71 -2384 74 -2378
rect 78 -2384 81 -2378
rect 85 -2384 88 -2378
rect 92 -2384 95 -2378
rect 99 -2384 102 -2378
rect 106 -2384 109 -2378
rect 113 -2384 116 -2378
rect 120 -2384 123 -2378
rect 127 -2384 130 -2378
rect 134 -2384 137 -2378
rect 141 -2384 144 -2378
rect 148 -2384 154 -2378
rect 155 -2384 158 -2378
rect 162 -2384 168 -2378
rect 169 -2384 175 -2378
rect 176 -2384 182 -2378
rect 183 -2384 189 -2378
rect 190 -2384 193 -2378
rect 197 -2384 200 -2378
rect 204 -2384 207 -2378
rect 211 -2384 214 -2378
rect 218 -2384 221 -2378
rect 225 -2384 228 -2378
rect 232 -2384 238 -2378
rect 239 -2384 242 -2378
rect 246 -2384 249 -2378
rect 253 -2384 256 -2378
rect 260 -2384 263 -2378
rect 267 -2384 273 -2378
rect 274 -2384 277 -2378
rect 281 -2384 284 -2378
rect 288 -2384 291 -2378
rect 295 -2384 298 -2378
rect 302 -2384 308 -2378
rect 309 -2384 312 -2378
rect 316 -2384 319 -2378
rect 323 -2384 326 -2378
rect 330 -2384 333 -2378
rect 337 -2384 340 -2378
rect 344 -2384 347 -2378
rect 351 -2384 354 -2378
rect 358 -2384 361 -2378
rect 365 -2384 368 -2378
rect 372 -2384 375 -2378
rect 379 -2384 385 -2378
rect 386 -2384 389 -2378
rect 393 -2384 396 -2378
rect 400 -2384 403 -2378
rect 407 -2384 410 -2378
rect 414 -2384 417 -2378
rect 421 -2384 424 -2378
rect 428 -2384 431 -2378
rect 435 -2384 438 -2378
rect 442 -2384 445 -2378
rect 449 -2384 455 -2378
rect 456 -2384 459 -2378
rect 463 -2384 466 -2378
rect 470 -2384 473 -2378
rect 477 -2384 480 -2378
rect 484 -2384 487 -2378
rect 491 -2384 494 -2378
rect 498 -2384 501 -2378
rect 505 -2384 508 -2378
rect 512 -2384 518 -2378
rect 519 -2384 522 -2378
rect 526 -2384 532 -2378
rect 533 -2384 536 -2378
rect 540 -2384 543 -2378
rect 547 -2384 550 -2378
rect 554 -2384 560 -2378
rect 561 -2384 564 -2378
rect 568 -2384 571 -2378
rect 575 -2384 578 -2378
rect 582 -2384 585 -2378
rect 589 -2384 592 -2378
rect 596 -2384 599 -2378
rect 603 -2384 606 -2378
rect 610 -2384 616 -2378
rect 617 -2384 620 -2378
rect 624 -2384 627 -2378
rect 631 -2384 634 -2378
rect 638 -2384 641 -2378
rect 645 -2384 648 -2378
rect 652 -2384 655 -2378
rect 659 -2384 662 -2378
rect 666 -2384 669 -2378
rect 673 -2384 676 -2378
rect 680 -2384 683 -2378
rect 687 -2384 690 -2378
rect 694 -2384 700 -2378
rect 701 -2384 704 -2378
rect 708 -2384 711 -2378
rect 715 -2384 718 -2378
rect 729 -2384 732 -2378
rect 736 -2384 739 -2378
rect 743 -2384 746 -2378
rect 750 -2384 753 -2378
rect 757 -2384 760 -2378
rect 764 -2384 767 -2378
rect 771 -2384 774 -2378
rect 778 -2384 781 -2378
rect 792 -2384 795 -2378
rect 799 -2384 802 -2378
rect 813 -2384 816 -2378
rect 897 -2384 900 -2378
rect 904 -2384 907 -2378
rect 939 -2384 942 -2378
rect 974 -2384 980 -2378
rect 981 -2384 984 -2378
rect 988 -2384 991 -2378
rect 1002 -2384 1008 -2378
rect 197 -2435 200 -2429
rect 218 -2435 221 -2429
rect 225 -2435 228 -2429
rect 232 -2435 235 -2429
rect 239 -2435 242 -2429
rect 246 -2435 249 -2429
rect 253 -2435 256 -2429
rect 260 -2435 263 -2429
rect 267 -2435 270 -2429
rect 274 -2435 277 -2429
rect 281 -2435 284 -2429
rect 288 -2435 291 -2429
rect 295 -2435 298 -2429
rect 302 -2435 305 -2429
rect 309 -2435 312 -2429
rect 316 -2435 319 -2429
rect 323 -2435 329 -2429
rect 330 -2435 333 -2429
rect 337 -2435 340 -2429
rect 344 -2435 347 -2429
rect 351 -2435 357 -2429
rect 358 -2435 361 -2429
rect 365 -2435 371 -2429
rect 372 -2435 375 -2429
rect 379 -2435 385 -2429
rect 386 -2435 389 -2429
rect 393 -2435 396 -2429
rect 400 -2435 403 -2429
rect 407 -2435 410 -2429
rect 414 -2435 420 -2429
rect 421 -2435 424 -2429
rect 428 -2435 431 -2429
rect 435 -2435 438 -2429
rect 442 -2435 445 -2429
rect 449 -2435 455 -2429
rect 456 -2435 462 -2429
rect 463 -2435 466 -2429
rect 470 -2435 473 -2429
rect 477 -2435 480 -2429
rect 484 -2435 490 -2429
rect 491 -2435 494 -2429
rect 498 -2435 501 -2429
rect 505 -2435 511 -2429
rect 512 -2435 518 -2429
rect 519 -2435 525 -2429
rect 526 -2435 529 -2429
rect 533 -2435 536 -2429
rect 540 -2435 543 -2429
rect 547 -2435 550 -2429
rect 554 -2435 557 -2429
rect 561 -2435 564 -2429
rect 568 -2435 574 -2429
rect 575 -2435 578 -2429
rect 582 -2435 585 -2429
rect 589 -2435 592 -2429
rect 596 -2435 599 -2429
rect 603 -2435 606 -2429
rect 610 -2435 613 -2429
rect 617 -2435 620 -2429
rect 624 -2435 627 -2429
rect 631 -2435 634 -2429
rect 645 -2435 648 -2429
rect 652 -2435 655 -2429
rect 659 -2435 662 -2429
rect 666 -2435 669 -2429
rect 673 -2435 676 -2429
rect 680 -2435 686 -2429
rect 687 -2435 693 -2429
rect 715 -2435 718 -2429
rect 722 -2435 725 -2429
rect 729 -2435 732 -2429
rect 736 -2435 739 -2429
rect 743 -2435 749 -2429
rect 750 -2435 753 -2429
rect 757 -2435 760 -2429
rect 764 -2435 767 -2429
rect 771 -2435 774 -2429
rect 799 -2435 802 -2429
rect 806 -2435 809 -2429
rect 827 -2435 830 -2429
rect 890 -2435 893 -2429
rect 897 -2435 900 -2429
rect 904 -2435 910 -2429
rect 225 -2476 228 -2470
rect 232 -2476 238 -2470
rect 239 -2476 242 -2470
rect 246 -2476 249 -2470
rect 253 -2476 259 -2470
rect 295 -2476 298 -2470
rect 309 -2476 312 -2470
rect 330 -2476 333 -2470
rect 337 -2476 343 -2470
rect 344 -2476 350 -2470
rect 351 -2476 354 -2470
rect 358 -2476 361 -2470
rect 365 -2476 368 -2470
rect 372 -2476 375 -2470
rect 386 -2476 389 -2470
rect 393 -2476 396 -2470
rect 400 -2476 403 -2470
rect 407 -2476 410 -2470
rect 421 -2476 424 -2470
rect 428 -2476 434 -2470
rect 435 -2476 438 -2470
rect 442 -2476 448 -2470
rect 449 -2476 455 -2470
rect 456 -2476 459 -2470
rect 463 -2476 466 -2470
rect 470 -2476 473 -2470
rect 477 -2476 480 -2470
rect 484 -2476 487 -2470
rect 491 -2476 494 -2470
rect 498 -2476 501 -2470
rect 505 -2476 511 -2470
rect 512 -2476 515 -2470
rect 526 -2476 529 -2470
rect 540 -2476 543 -2470
rect 547 -2476 550 -2470
rect 575 -2476 578 -2470
rect 596 -2476 599 -2470
rect 603 -2476 609 -2470
rect 610 -2476 616 -2470
rect 617 -2476 620 -2470
rect 624 -2476 627 -2470
rect 631 -2476 634 -2470
rect 638 -2476 641 -2470
rect 645 -2476 651 -2470
rect 652 -2476 655 -2470
rect 659 -2476 662 -2470
rect 673 -2476 676 -2470
rect 687 -2476 690 -2470
rect 701 -2476 704 -2470
rect 722 -2476 725 -2470
rect 743 -2476 746 -2470
rect 750 -2476 756 -2470
rect 806 -2476 809 -2470
rect 813 -2476 819 -2470
rect 827 -2476 830 -2470
rect 834 -2476 840 -2470
rect 897 -2476 900 -2470
rect 225 -2497 228 -2491
rect 232 -2497 238 -2491
rect 239 -2497 242 -2491
rect 358 -2497 361 -2491
rect 365 -2497 371 -2491
rect 372 -2497 375 -2491
rect 379 -2497 382 -2491
rect 386 -2497 392 -2491
rect 393 -2497 399 -2491
rect 400 -2497 406 -2491
rect 407 -2497 410 -2491
rect 533 -2497 536 -2491
rect 547 -2497 553 -2491
rect 554 -2497 560 -2491
rect 603 -2497 606 -2491
rect 610 -2497 616 -2491
rect 631 -2497 634 -2491
rect 652 -2497 658 -2491
rect 659 -2497 662 -2491
rect 687 -2497 693 -2491
rect 701 -2497 704 -2491
rect 722 -2497 728 -2491
rect 897 -2497 903 -2491
rect 904 -2497 907 -2491
<< polysilicon >>
rect 152 -7 153 -5
rect 149 -13 150 -11
rect 205 -7 206 -5
rect 208 -13 209 -11
rect 338 -7 339 -5
rect 341 -7 342 -5
rect 341 -13 342 -11
rect 345 -7 346 -5
rect 345 -13 346 -11
rect 352 -7 353 -5
rect 352 -13 353 -11
rect 359 -7 360 -5
rect 359 -13 360 -11
rect 366 -7 367 -5
rect 366 -13 367 -11
rect 376 -7 377 -5
rect 373 -13 374 -11
rect 394 -7 395 -5
rect 394 -13 395 -11
rect 401 -13 402 -11
rect 404 -13 405 -11
rect 408 -7 409 -5
rect 411 -7 412 -5
rect 432 -7 433 -5
rect 429 -13 430 -11
rect 432 -13 433 -11
rect 436 -13 437 -11
rect 439 -13 440 -11
rect 450 -7 451 -5
rect 450 -13 451 -11
rect 464 -7 465 -5
rect 464 -13 465 -11
rect 471 -7 472 -5
rect 474 -13 475 -11
rect 481 -7 482 -5
rect 478 -13 479 -11
rect 492 -7 493 -5
rect 492 -13 493 -11
rect 513 -7 514 -5
rect 513 -13 514 -11
rect 576 -7 577 -5
rect 576 -13 577 -11
rect 128 -38 129 -36
rect 128 -44 129 -42
rect 198 -38 199 -36
rect 198 -44 199 -42
rect 219 -38 220 -36
rect 219 -44 220 -42
rect 243 -38 244 -36
rect 240 -44 241 -42
rect 243 -44 244 -42
rect 254 -38 255 -36
rect 254 -44 255 -42
rect 282 -38 283 -36
rect 282 -44 283 -42
rect 289 -38 290 -36
rect 292 -38 293 -36
rect 289 -44 290 -42
rect 296 -38 297 -36
rect 296 -44 297 -42
rect 303 -38 304 -36
rect 303 -44 304 -42
rect 310 -38 311 -36
rect 310 -44 311 -42
rect 320 -38 321 -36
rect 320 -44 321 -42
rect 324 -38 325 -36
rect 327 -38 328 -36
rect 324 -44 325 -42
rect 331 -38 332 -36
rect 331 -44 332 -42
rect 338 -38 339 -36
rect 338 -44 339 -42
rect 345 -38 346 -36
rect 345 -44 346 -42
rect 352 -38 353 -36
rect 352 -44 353 -42
rect 359 -38 360 -36
rect 359 -44 360 -42
rect 366 -38 367 -36
rect 366 -44 367 -42
rect 373 -38 374 -36
rect 376 -38 377 -36
rect 373 -44 374 -42
rect 380 -38 381 -36
rect 380 -44 381 -42
rect 387 -38 388 -36
rect 387 -44 388 -42
rect 394 -38 395 -36
rect 394 -44 395 -42
rect 397 -44 398 -42
rect 401 -38 402 -36
rect 401 -44 402 -42
rect 408 -38 409 -36
rect 408 -44 409 -42
rect 415 -38 416 -36
rect 415 -44 416 -42
rect 422 -38 423 -36
rect 422 -44 423 -42
rect 432 -38 433 -36
rect 432 -44 433 -42
rect 436 -38 437 -36
rect 436 -44 437 -42
rect 446 -38 447 -36
rect 443 -44 444 -42
rect 446 -44 447 -42
rect 450 -38 451 -36
rect 450 -44 451 -42
rect 457 -38 458 -36
rect 457 -44 458 -42
rect 464 -38 465 -36
rect 464 -44 465 -42
rect 471 -38 472 -36
rect 471 -44 472 -42
rect 478 -38 479 -36
rect 478 -44 479 -42
rect 485 -38 486 -36
rect 485 -44 486 -42
rect 492 -44 493 -42
rect 495 -44 496 -42
rect 502 -38 503 -36
rect 499 -44 500 -42
rect 502 -44 503 -42
rect 506 -38 507 -36
rect 506 -44 507 -42
rect 513 -38 514 -36
rect 513 -44 514 -42
rect 527 -38 528 -36
rect 527 -44 528 -42
rect 534 -38 535 -36
rect 534 -44 535 -42
rect 541 -38 542 -36
rect 541 -44 542 -42
rect 548 -38 549 -36
rect 548 -44 549 -42
rect 593 -38 594 -36
rect 590 -44 591 -42
rect 593 -44 594 -42
rect 618 -38 619 -36
rect 618 -44 619 -42
rect 625 -38 626 -36
rect 625 -44 626 -42
rect 114 -91 115 -89
rect 114 -97 115 -95
rect 117 -97 118 -95
rect 142 -91 143 -89
rect 142 -97 143 -95
rect 163 -91 164 -89
rect 163 -97 164 -95
rect 170 -91 171 -89
rect 170 -97 171 -95
rect 177 -91 178 -89
rect 177 -97 178 -95
rect 184 -91 185 -89
rect 184 -97 185 -95
rect 191 -91 192 -89
rect 191 -97 192 -95
rect 198 -91 199 -89
rect 198 -97 199 -95
rect 205 -91 206 -89
rect 205 -97 206 -95
rect 212 -91 213 -89
rect 212 -97 213 -95
rect 219 -91 220 -89
rect 219 -97 220 -95
rect 226 -91 227 -89
rect 226 -97 227 -95
rect 233 -91 234 -89
rect 233 -97 234 -95
rect 240 -91 241 -89
rect 240 -97 241 -95
rect 247 -91 248 -89
rect 247 -97 248 -95
rect 254 -91 255 -89
rect 254 -97 255 -95
rect 261 -91 262 -89
rect 261 -97 262 -95
rect 268 -91 269 -89
rect 268 -97 269 -95
rect 275 -91 276 -89
rect 275 -97 276 -95
rect 278 -97 279 -95
rect 282 -91 283 -89
rect 282 -97 283 -95
rect 289 -91 290 -89
rect 289 -97 290 -95
rect 296 -91 297 -89
rect 296 -97 297 -95
rect 303 -91 304 -89
rect 303 -97 304 -95
rect 310 -91 311 -89
rect 310 -97 311 -95
rect 317 -91 318 -89
rect 317 -97 318 -95
rect 324 -91 325 -89
rect 324 -97 325 -95
rect 334 -91 335 -89
rect 331 -97 332 -95
rect 334 -97 335 -95
rect 338 -91 339 -89
rect 338 -97 339 -95
rect 345 -91 346 -89
rect 348 -91 349 -89
rect 345 -97 346 -95
rect 352 -91 353 -89
rect 352 -97 353 -95
rect 359 -91 360 -89
rect 359 -97 360 -95
rect 366 -91 367 -89
rect 369 -91 370 -89
rect 369 -97 370 -95
rect 373 -91 374 -89
rect 373 -97 374 -95
rect 376 -97 377 -95
rect 380 -91 381 -89
rect 380 -97 381 -95
rect 383 -97 384 -95
rect 387 -91 388 -89
rect 390 -91 391 -89
rect 387 -97 388 -95
rect 397 -91 398 -89
rect 394 -97 395 -95
rect 401 -91 402 -89
rect 401 -97 402 -95
rect 408 -91 409 -89
rect 408 -97 409 -95
rect 415 -91 416 -89
rect 415 -97 416 -95
rect 422 -91 423 -89
rect 422 -97 423 -95
rect 429 -91 430 -89
rect 429 -97 430 -95
rect 436 -91 437 -89
rect 436 -97 437 -95
rect 443 -91 444 -89
rect 443 -97 444 -95
rect 450 -91 451 -89
rect 450 -97 451 -95
rect 453 -97 454 -95
rect 457 -91 458 -89
rect 457 -97 458 -95
rect 464 -91 465 -89
rect 464 -97 465 -95
rect 474 -91 475 -89
rect 471 -97 472 -95
rect 474 -97 475 -95
rect 478 -91 479 -89
rect 481 -91 482 -89
rect 481 -97 482 -95
rect 485 -91 486 -89
rect 485 -97 486 -95
rect 492 -91 493 -89
rect 492 -97 493 -95
rect 499 -91 500 -89
rect 499 -97 500 -95
rect 506 -91 507 -89
rect 506 -97 507 -95
rect 513 -91 514 -89
rect 513 -97 514 -95
rect 520 -91 521 -89
rect 520 -97 521 -95
rect 527 -91 528 -89
rect 527 -97 528 -95
rect 534 -91 535 -89
rect 534 -97 535 -95
rect 541 -91 542 -89
rect 541 -97 542 -95
rect 548 -91 549 -89
rect 548 -97 549 -95
rect 555 -91 556 -89
rect 555 -97 556 -95
rect 562 -91 563 -89
rect 562 -97 563 -95
rect 569 -91 570 -89
rect 569 -97 570 -95
rect 576 -91 577 -89
rect 576 -97 577 -95
rect 583 -91 584 -89
rect 583 -97 584 -95
rect 590 -91 591 -89
rect 593 -91 594 -89
rect 593 -97 594 -95
rect 597 -91 598 -89
rect 597 -97 598 -95
rect 604 -91 605 -89
rect 604 -97 605 -95
rect 611 -91 612 -89
rect 611 -97 612 -95
rect 618 -91 619 -89
rect 618 -97 619 -95
rect 625 -91 626 -89
rect 625 -97 626 -95
rect 632 -91 633 -89
rect 632 -97 633 -95
rect 639 -91 640 -89
rect 639 -97 640 -95
rect 646 -91 647 -89
rect 646 -97 647 -95
rect 653 -91 654 -89
rect 653 -97 654 -95
rect 660 -91 661 -89
rect 660 -97 661 -95
rect 667 -91 668 -89
rect 667 -97 668 -95
rect 674 -91 675 -89
rect 674 -97 675 -95
rect 681 -91 682 -89
rect 681 -97 682 -95
rect 688 -91 689 -89
rect 691 -91 692 -89
rect 688 -97 689 -95
rect 51 -158 52 -156
rect 51 -164 52 -162
rect 58 -158 59 -156
rect 58 -164 59 -162
rect 65 -158 66 -156
rect 65 -164 66 -162
rect 72 -158 73 -156
rect 72 -164 73 -162
rect 82 -158 83 -156
rect 86 -158 87 -156
rect 86 -164 87 -162
rect 93 -158 94 -156
rect 93 -164 94 -162
rect 100 -158 101 -156
rect 100 -164 101 -162
rect 103 -164 104 -162
rect 107 -158 108 -156
rect 107 -164 108 -162
rect 114 -158 115 -156
rect 114 -164 115 -162
rect 121 -158 122 -156
rect 121 -164 122 -162
rect 128 -158 129 -156
rect 128 -164 129 -162
rect 135 -158 136 -156
rect 135 -164 136 -162
rect 145 -158 146 -156
rect 142 -164 143 -162
rect 145 -164 146 -162
rect 152 -158 153 -156
rect 149 -164 150 -162
rect 152 -164 153 -162
rect 156 -158 157 -156
rect 156 -164 157 -162
rect 163 -158 164 -156
rect 163 -164 164 -162
rect 170 -158 171 -156
rect 170 -164 171 -162
rect 177 -158 178 -156
rect 177 -164 178 -162
rect 184 -158 185 -156
rect 187 -158 188 -156
rect 184 -164 185 -162
rect 194 -158 195 -156
rect 191 -164 192 -162
rect 194 -164 195 -162
rect 198 -158 199 -156
rect 201 -158 202 -156
rect 201 -164 202 -162
rect 205 -158 206 -156
rect 205 -164 206 -162
rect 212 -158 213 -156
rect 212 -164 213 -162
rect 219 -158 220 -156
rect 219 -164 220 -162
rect 226 -158 227 -156
rect 226 -164 227 -162
rect 233 -158 234 -156
rect 233 -164 234 -162
rect 240 -158 241 -156
rect 240 -164 241 -162
rect 247 -158 248 -156
rect 247 -164 248 -162
rect 254 -158 255 -156
rect 254 -164 255 -162
rect 261 -158 262 -156
rect 261 -164 262 -162
rect 268 -158 269 -156
rect 268 -164 269 -162
rect 275 -158 276 -156
rect 275 -164 276 -162
rect 282 -158 283 -156
rect 282 -164 283 -162
rect 289 -158 290 -156
rect 289 -164 290 -162
rect 296 -158 297 -156
rect 296 -164 297 -162
rect 303 -158 304 -156
rect 303 -164 304 -162
rect 310 -158 311 -156
rect 310 -164 311 -162
rect 317 -158 318 -156
rect 317 -164 318 -162
rect 324 -158 325 -156
rect 324 -164 325 -162
rect 331 -158 332 -156
rect 331 -164 332 -162
rect 338 -158 339 -156
rect 338 -164 339 -162
rect 345 -158 346 -156
rect 345 -164 346 -162
rect 352 -158 353 -156
rect 352 -164 353 -162
rect 359 -158 360 -156
rect 359 -164 360 -162
rect 366 -158 367 -156
rect 366 -164 367 -162
rect 373 -158 374 -156
rect 373 -164 374 -162
rect 380 -158 381 -156
rect 380 -164 381 -162
rect 387 -158 388 -156
rect 387 -164 388 -162
rect 394 -158 395 -156
rect 394 -164 395 -162
rect 401 -158 402 -156
rect 401 -164 402 -162
rect 411 -158 412 -156
rect 408 -164 409 -162
rect 411 -164 412 -162
rect 415 -158 416 -156
rect 418 -158 419 -156
rect 415 -164 416 -162
rect 422 -158 423 -156
rect 422 -164 423 -162
rect 429 -158 430 -156
rect 429 -164 430 -162
rect 436 -158 437 -156
rect 436 -164 437 -162
rect 443 -158 444 -156
rect 443 -164 444 -162
rect 453 -158 454 -156
rect 450 -164 451 -162
rect 453 -164 454 -162
rect 457 -158 458 -156
rect 457 -164 458 -162
rect 464 -158 465 -156
rect 467 -158 468 -156
rect 464 -164 465 -162
rect 471 -158 472 -156
rect 474 -158 475 -156
rect 474 -164 475 -162
rect 478 -158 479 -156
rect 478 -164 479 -162
rect 481 -164 482 -162
rect 485 -158 486 -156
rect 485 -164 486 -162
rect 495 -158 496 -156
rect 492 -164 493 -162
rect 495 -164 496 -162
rect 499 -158 500 -156
rect 499 -164 500 -162
rect 506 -158 507 -156
rect 506 -164 507 -162
rect 513 -158 514 -156
rect 513 -164 514 -162
rect 520 -158 521 -156
rect 520 -164 521 -162
rect 527 -158 528 -156
rect 527 -164 528 -162
rect 534 -158 535 -156
rect 534 -164 535 -162
rect 541 -158 542 -156
rect 541 -164 542 -162
rect 548 -158 549 -156
rect 548 -164 549 -162
rect 555 -158 556 -156
rect 555 -164 556 -162
rect 562 -158 563 -156
rect 562 -164 563 -162
rect 569 -158 570 -156
rect 569 -164 570 -162
rect 576 -158 577 -156
rect 579 -158 580 -156
rect 576 -164 577 -162
rect 583 -158 584 -156
rect 583 -164 584 -162
rect 590 -158 591 -156
rect 590 -164 591 -162
rect 597 -158 598 -156
rect 597 -164 598 -162
rect 604 -158 605 -156
rect 604 -164 605 -162
rect 611 -158 612 -156
rect 611 -164 612 -162
rect 618 -158 619 -156
rect 618 -164 619 -162
rect 625 -158 626 -156
rect 625 -164 626 -162
rect 632 -158 633 -156
rect 632 -164 633 -162
rect 639 -158 640 -156
rect 639 -164 640 -162
rect 646 -158 647 -156
rect 646 -164 647 -162
rect 653 -158 654 -156
rect 653 -164 654 -162
rect 660 -158 661 -156
rect 660 -164 661 -162
rect 667 -158 668 -156
rect 667 -164 668 -162
rect 674 -158 675 -156
rect 674 -164 675 -162
rect 681 -158 682 -156
rect 681 -164 682 -162
rect 688 -158 689 -156
rect 688 -164 689 -162
rect 695 -158 696 -156
rect 695 -164 696 -162
rect 702 -158 703 -156
rect 702 -164 703 -162
rect 709 -158 710 -156
rect 709 -164 710 -162
rect 716 -158 717 -156
rect 716 -164 717 -162
rect 723 -158 724 -156
rect 723 -164 724 -162
rect 730 -158 731 -156
rect 730 -164 731 -162
rect 737 -158 738 -156
rect 737 -164 738 -162
rect 744 -158 745 -156
rect 744 -164 745 -162
rect 751 -158 752 -156
rect 751 -164 752 -162
rect 758 -158 759 -156
rect 758 -164 759 -162
rect 765 -158 766 -156
rect 765 -164 766 -162
rect 772 -158 773 -156
rect 772 -164 773 -162
rect 779 -158 780 -156
rect 779 -164 780 -162
rect 786 -158 787 -156
rect 786 -164 787 -162
rect 793 -158 794 -156
rect 793 -164 794 -162
rect 800 -158 801 -156
rect 800 -164 801 -162
rect 807 -158 808 -156
rect 807 -164 808 -162
rect 814 -158 815 -156
rect 814 -164 815 -162
rect 821 -158 822 -156
rect 821 -164 822 -162
rect 44 -239 45 -237
rect 44 -245 45 -243
rect 51 -239 52 -237
rect 51 -245 52 -243
rect 58 -239 59 -237
rect 58 -245 59 -243
rect 65 -239 66 -237
rect 65 -245 66 -243
rect 72 -239 73 -237
rect 72 -245 73 -243
rect 79 -239 80 -237
rect 79 -245 80 -243
rect 86 -239 87 -237
rect 86 -245 87 -243
rect 93 -239 94 -237
rect 93 -245 94 -243
rect 100 -245 101 -243
rect 103 -245 104 -243
rect 107 -239 108 -237
rect 107 -245 108 -243
rect 117 -239 118 -237
rect 114 -245 115 -243
rect 117 -245 118 -243
rect 121 -239 122 -237
rect 124 -239 125 -237
rect 121 -245 122 -243
rect 124 -245 125 -243
rect 128 -239 129 -237
rect 128 -245 129 -243
rect 135 -239 136 -237
rect 138 -239 139 -237
rect 135 -245 136 -243
rect 142 -239 143 -237
rect 142 -245 143 -243
rect 149 -239 150 -237
rect 149 -245 150 -243
rect 156 -239 157 -237
rect 156 -245 157 -243
rect 163 -239 164 -237
rect 166 -239 167 -237
rect 163 -245 164 -243
rect 166 -245 167 -243
rect 170 -239 171 -237
rect 170 -245 171 -243
rect 177 -239 178 -237
rect 177 -245 178 -243
rect 184 -239 185 -237
rect 184 -245 185 -243
rect 191 -239 192 -237
rect 191 -245 192 -243
rect 198 -239 199 -237
rect 198 -245 199 -243
rect 205 -239 206 -237
rect 205 -245 206 -243
rect 212 -239 213 -237
rect 212 -245 213 -243
rect 219 -239 220 -237
rect 219 -245 220 -243
rect 226 -239 227 -237
rect 226 -245 227 -243
rect 233 -239 234 -237
rect 233 -245 234 -243
rect 240 -239 241 -237
rect 240 -245 241 -243
rect 247 -239 248 -237
rect 247 -245 248 -243
rect 254 -239 255 -237
rect 257 -239 258 -237
rect 254 -245 255 -243
rect 257 -245 258 -243
rect 261 -239 262 -237
rect 261 -245 262 -243
rect 268 -239 269 -237
rect 268 -245 269 -243
rect 275 -239 276 -237
rect 275 -245 276 -243
rect 282 -239 283 -237
rect 285 -239 286 -237
rect 282 -245 283 -243
rect 285 -245 286 -243
rect 289 -239 290 -237
rect 292 -239 293 -237
rect 289 -245 290 -243
rect 292 -245 293 -243
rect 296 -239 297 -237
rect 296 -245 297 -243
rect 303 -239 304 -237
rect 303 -245 304 -243
rect 310 -239 311 -237
rect 310 -245 311 -243
rect 317 -239 318 -237
rect 317 -245 318 -243
rect 324 -239 325 -237
rect 324 -245 325 -243
rect 331 -239 332 -237
rect 331 -245 332 -243
rect 338 -239 339 -237
rect 338 -245 339 -243
rect 345 -239 346 -237
rect 348 -239 349 -237
rect 345 -245 346 -243
rect 348 -245 349 -243
rect 352 -239 353 -237
rect 355 -239 356 -237
rect 352 -245 353 -243
rect 355 -245 356 -243
rect 359 -239 360 -237
rect 362 -239 363 -237
rect 359 -245 360 -243
rect 362 -245 363 -243
rect 366 -239 367 -237
rect 366 -245 367 -243
rect 376 -239 377 -237
rect 376 -245 377 -243
rect 380 -239 381 -237
rect 380 -245 381 -243
rect 387 -239 388 -237
rect 387 -245 388 -243
rect 394 -239 395 -237
rect 394 -245 395 -243
rect 401 -239 402 -237
rect 404 -239 405 -237
rect 401 -245 402 -243
rect 408 -239 409 -237
rect 408 -245 409 -243
rect 415 -239 416 -237
rect 415 -245 416 -243
rect 422 -239 423 -237
rect 425 -239 426 -237
rect 422 -245 423 -243
rect 425 -245 426 -243
rect 429 -239 430 -237
rect 429 -245 430 -243
rect 436 -239 437 -237
rect 439 -239 440 -237
rect 436 -245 437 -243
rect 443 -239 444 -237
rect 443 -245 444 -243
rect 450 -239 451 -237
rect 450 -245 451 -243
rect 457 -239 458 -237
rect 460 -239 461 -237
rect 457 -245 458 -243
rect 464 -239 465 -237
rect 464 -245 465 -243
rect 471 -239 472 -237
rect 474 -239 475 -237
rect 474 -245 475 -243
rect 478 -239 479 -237
rect 478 -245 479 -243
rect 485 -239 486 -237
rect 485 -245 486 -243
rect 492 -239 493 -237
rect 495 -239 496 -237
rect 492 -245 493 -243
rect 495 -245 496 -243
rect 499 -239 500 -237
rect 499 -245 500 -243
rect 506 -239 507 -237
rect 506 -245 507 -243
rect 513 -239 514 -237
rect 513 -245 514 -243
rect 520 -239 521 -237
rect 520 -245 521 -243
rect 527 -239 528 -237
rect 534 -239 535 -237
rect 534 -245 535 -243
rect 541 -239 542 -237
rect 541 -245 542 -243
rect 548 -239 549 -237
rect 548 -245 549 -243
rect 555 -239 556 -237
rect 555 -245 556 -243
rect 562 -239 563 -237
rect 562 -245 563 -243
rect 569 -239 570 -237
rect 569 -245 570 -243
rect 576 -239 577 -237
rect 576 -245 577 -243
rect 579 -245 580 -243
rect 583 -239 584 -237
rect 583 -245 584 -243
rect 590 -239 591 -237
rect 590 -245 591 -243
rect 597 -239 598 -237
rect 597 -245 598 -243
rect 604 -239 605 -237
rect 604 -245 605 -243
rect 611 -239 612 -237
rect 611 -245 612 -243
rect 618 -239 619 -237
rect 618 -245 619 -243
rect 625 -239 626 -237
rect 625 -245 626 -243
rect 632 -239 633 -237
rect 632 -245 633 -243
rect 639 -239 640 -237
rect 639 -245 640 -243
rect 646 -239 647 -237
rect 646 -245 647 -243
rect 653 -239 654 -237
rect 653 -245 654 -243
rect 660 -239 661 -237
rect 660 -245 661 -243
rect 667 -239 668 -237
rect 667 -245 668 -243
rect 674 -239 675 -237
rect 674 -245 675 -243
rect 681 -239 682 -237
rect 681 -245 682 -243
rect 688 -239 689 -237
rect 688 -245 689 -243
rect 695 -239 696 -237
rect 695 -245 696 -243
rect 702 -239 703 -237
rect 702 -245 703 -243
rect 709 -239 710 -237
rect 709 -245 710 -243
rect 716 -239 717 -237
rect 716 -245 717 -243
rect 723 -239 724 -237
rect 723 -245 724 -243
rect 730 -239 731 -237
rect 730 -245 731 -243
rect 737 -239 738 -237
rect 737 -245 738 -243
rect 744 -239 745 -237
rect 744 -245 745 -243
rect 751 -239 752 -237
rect 751 -245 752 -243
rect 758 -239 759 -237
rect 758 -245 759 -243
rect 765 -239 766 -237
rect 765 -245 766 -243
rect 772 -239 773 -237
rect 772 -245 773 -243
rect 779 -239 780 -237
rect 779 -245 780 -243
rect 786 -239 787 -237
rect 786 -245 787 -243
rect 793 -239 794 -237
rect 793 -245 794 -243
rect 800 -239 801 -237
rect 800 -245 801 -243
rect 807 -239 808 -237
rect 807 -245 808 -243
rect 814 -239 815 -237
rect 814 -245 815 -243
rect 821 -239 822 -237
rect 821 -245 822 -243
rect 828 -239 829 -237
rect 828 -245 829 -243
rect 835 -239 836 -237
rect 835 -245 836 -243
rect 842 -239 843 -237
rect 842 -245 843 -243
rect 849 -239 850 -237
rect 849 -245 850 -243
rect 859 -239 860 -237
rect 863 -239 864 -237
rect 863 -245 864 -243
rect 2 -328 3 -326
rect 2 -334 3 -332
rect 9 -328 10 -326
rect 9 -334 10 -332
rect 16 -328 17 -326
rect 16 -334 17 -332
rect 23 -328 24 -326
rect 23 -334 24 -332
rect 30 -328 31 -326
rect 30 -334 31 -332
rect 37 -328 38 -326
rect 37 -334 38 -332
rect 44 -328 45 -326
rect 44 -334 45 -332
rect 51 -328 52 -326
rect 51 -334 52 -332
rect 58 -328 59 -326
rect 58 -334 59 -332
rect 65 -328 66 -326
rect 68 -328 69 -326
rect 68 -334 69 -332
rect 72 -328 73 -326
rect 72 -334 73 -332
rect 79 -328 80 -326
rect 79 -334 80 -332
rect 86 -328 87 -326
rect 86 -334 87 -332
rect 93 -328 94 -326
rect 93 -334 94 -332
rect 100 -328 101 -326
rect 100 -334 101 -332
rect 107 -328 108 -326
rect 107 -334 108 -332
rect 114 -328 115 -326
rect 114 -334 115 -332
rect 121 -328 122 -326
rect 121 -334 122 -332
rect 128 -334 129 -332
rect 131 -334 132 -332
rect 135 -328 136 -326
rect 135 -334 136 -332
rect 142 -328 143 -326
rect 142 -334 143 -332
rect 149 -328 150 -326
rect 149 -334 150 -332
rect 156 -328 157 -326
rect 156 -334 157 -332
rect 163 -328 164 -326
rect 163 -334 164 -332
rect 170 -328 171 -326
rect 170 -334 171 -332
rect 177 -328 178 -326
rect 177 -334 178 -332
rect 184 -328 185 -326
rect 184 -334 185 -332
rect 191 -328 192 -326
rect 198 -328 199 -326
rect 198 -334 199 -332
rect 205 -328 206 -326
rect 205 -334 206 -332
rect 212 -328 213 -326
rect 212 -334 213 -332
rect 219 -328 220 -326
rect 219 -334 220 -332
rect 226 -328 227 -326
rect 226 -334 227 -332
rect 233 -328 234 -326
rect 233 -334 234 -332
rect 240 -328 241 -326
rect 240 -334 241 -332
rect 247 -328 248 -326
rect 247 -334 248 -332
rect 254 -328 255 -326
rect 254 -334 255 -332
rect 261 -328 262 -326
rect 261 -334 262 -332
rect 268 -328 269 -326
rect 268 -334 269 -332
rect 275 -328 276 -326
rect 275 -334 276 -332
rect 282 -328 283 -326
rect 282 -334 283 -332
rect 289 -328 290 -326
rect 289 -334 290 -332
rect 296 -328 297 -326
rect 296 -334 297 -332
rect 303 -328 304 -326
rect 306 -328 307 -326
rect 306 -334 307 -332
rect 310 -328 311 -326
rect 310 -334 311 -332
rect 317 -328 318 -326
rect 317 -334 318 -332
rect 324 -328 325 -326
rect 324 -334 325 -332
rect 331 -328 332 -326
rect 331 -334 332 -332
rect 338 -328 339 -326
rect 338 -334 339 -332
rect 345 -328 346 -326
rect 345 -334 346 -332
rect 352 -328 353 -326
rect 352 -334 353 -332
rect 359 -328 360 -326
rect 359 -334 360 -332
rect 366 -328 367 -326
rect 366 -334 367 -332
rect 376 -328 377 -326
rect 373 -334 374 -332
rect 376 -334 377 -332
rect 380 -328 381 -326
rect 383 -328 384 -326
rect 383 -334 384 -332
rect 387 -328 388 -326
rect 387 -334 388 -332
rect 394 -328 395 -326
rect 397 -328 398 -326
rect 394 -334 395 -332
rect 397 -334 398 -332
rect 404 -328 405 -326
rect 401 -334 402 -332
rect 404 -334 405 -332
rect 408 -328 409 -326
rect 408 -334 409 -332
rect 418 -328 419 -326
rect 415 -334 416 -332
rect 418 -334 419 -332
rect 422 -328 423 -326
rect 425 -328 426 -326
rect 422 -334 423 -332
rect 425 -334 426 -332
rect 429 -328 430 -326
rect 429 -334 430 -332
rect 436 -328 437 -326
rect 439 -328 440 -326
rect 436 -334 437 -332
rect 439 -334 440 -332
rect 443 -328 444 -326
rect 446 -328 447 -326
rect 443 -334 444 -332
rect 446 -334 447 -332
rect 450 -328 451 -326
rect 453 -328 454 -326
rect 453 -334 454 -332
rect 457 -328 458 -326
rect 457 -334 458 -332
rect 460 -334 461 -332
rect 467 -328 468 -326
rect 464 -334 465 -332
rect 467 -334 468 -332
rect 471 -328 472 -326
rect 474 -328 475 -326
rect 471 -334 472 -332
rect 474 -334 475 -332
rect 478 -328 479 -326
rect 478 -334 479 -332
rect 485 -328 486 -326
rect 488 -328 489 -326
rect 485 -334 486 -332
rect 488 -334 489 -332
rect 492 -328 493 -326
rect 492 -334 493 -332
rect 499 -328 500 -326
rect 499 -334 500 -332
rect 506 -328 507 -326
rect 506 -334 507 -332
rect 513 -328 514 -326
rect 513 -334 514 -332
rect 520 -328 521 -326
rect 520 -334 521 -332
rect 527 -334 528 -332
rect 534 -328 535 -326
rect 534 -334 535 -332
rect 541 -328 542 -326
rect 541 -334 542 -332
rect 548 -328 549 -326
rect 551 -328 552 -326
rect 548 -334 549 -332
rect 551 -334 552 -332
rect 555 -328 556 -326
rect 555 -334 556 -332
rect 562 -328 563 -326
rect 562 -334 563 -332
rect 569 -328 570 -326
rect 569 -334 570 -332
rect 572 -334 573 -332
rect 576 -328 577 -326
rect 579 -328 580 -326
rect 576 -334 577 -332
rect 583 -328 584 -326
rect 583 -334 584 -332
rect 590 -328 591 -326
rect 590 -334 591 -332
rect 597 -328 598 -326
rect 597 -334 598 -332
rect 604 -328 605 -326
rect 604 -334 605 -332
rect 611 -328 612 -326
rect 611 -334 612 -332
rect 618 -328 619 -326
rect 618 -334 619 -332
rect 625 -328 626 -326
rect 625 -334 626 -332
rect 632 -328 633 -326
rect 632 -334 633 -332
rect 639 -328 640 -326
rect 639 -334 640 -332
rect 646 -328 647 -326
rect 646 -334 647 -332
rect 653 -328 654 -326
rect 653 -334 654 -332
rect 660 -328 661 -326
rect 660 -334 661 -332
rect 667 -328 668 -326
rect 667 -334 668 -332
rect 674 -328 675 -326
rect 674 -334 675 -332
rect 681 -328 682 -326
rect 681 -334 682 -332
rect 688 -328 689 -326
rect 688 -334 689 -332
rect 695 -328 696 -326
rect 695 -334 696 -332
rect 702 -328 703 -326
rect 702 -334 703 -332
rect 709 -328 710 -326
rect 709 -334 710 -332
rect 716 -328 717 -326
rect 716 -334 717 -332
rect 723 -328 724 -326
rect 723 -334 724 -332
rect 730 -328 731 -326
rect 730 -334 731 -332
rect 737 -328 738 -326
rect 737 -334 738 -332
rect 744 -328 745 -326
rect 744 -334 745 -332
rect 751 -328 752 -326
rect 751 -334 752 -332
rect 758 -328 759 -326
rect 758 -334 759 -332
rect 765 -328 766 -326
rect 765 -334 766 -332
rect 772 -328 773 -326
rect 772 -334 773 -332
rect 779 -328 780 -326
rect 779 -334 780 -332
rect 786 -328 787 -326
rect 786 -334 787 -332
rect 793 -328 794 -326
rect 793 -334 794 -332
rect 800 -328 801 -326
rect 800 -334 801 -332
rect 807 -328 808 -326
rect 807 -334 808 -332
rect 814 -328 815 -326
rect 814 -334 815 -332
rect 821 -328 822 -326
rect 821 -334 822 -332
rect 828 -328 829 -326
rect 828 -334 829 -332
rect 835 -328 836 -326
rect 835 -334 836 -332
rect 842 -328 843 -326
rect 842 -334 843 -332
rect 849 -328 850 -326
rect 849 -334 850 -332
rect 856 -328 857 -326
rect 856 -334 857 -332
rect 863 -328 864 -326
rect 863 -334 864 -332
rect 870 -328 871 -326
rect 870 -334 871 -332
rect 877 -328 878 -326
rect 877 -334 878 -332
rect 884 -328 885 -326
rect 884 -334 885 -332
rect 891 -328 892 -326
rect 891 -334 892 -332
rect 898 -328 899 -326
rect 898 -334 899 -332
rect 905 -328 906 -326
rect 905 -334 906 -332
rect 912 -328 913 -326
rect 912 -334 913 -332
rect 919 -328 920 -326
rect 919 -334 920 -332
rect 926 -328 927 -326
rect 926 -334 927 -332
rect 933 -328 934 -326
rect 933 -334 934 -332
rect 940 -328 941 -326
rect 940 -334 941 -332
rect 947 -328 948 -326
rect 947 -334 948 -332
rect 954 -328 955 -326
rect 954 -334 955 -332
rect 2 -415 3 -413
rect 2 -421 3 -419
rect 9 -415 10 -413
rect 9 -421 10 -419
rect 16 -415 17 -413
rect 16 -421 17 -419
rect 23 -415 24 -413
rect 23 -421 24 -419
rect 30 -415 31 -413
rect 30 -421 31 -419
rect 37 -415 38 -413
rect 37 -421 38 -419
rect 44 -415 45 -413
rect 44 -421 45 -419
rect 51 -415 52 -413
rect 51 -421 52 -419
rect 58 -415 59 -413
rect 58 -421 59 -419
rect 65 -415 66 -413
rect 68 -415 69 -413
rect 65 -421 66 -419
rect 68 -421 69 -419
rect 72 -415 73 -413
rect 75 -415 76 -413
rect 72 -421 73 -419
rect 75 -421 76 -419
rect 79 -415 80 -413
rect 82 -415 83 -413
rect 79 -421 80 -419
rect 82 -421 83 -419
rect 86 -415 87 -413
rect 89 -415 90 -413
rect 93 -415 94 -413
rect 96 -415 97 -413
rect 93 -421 94 -419
rect 96 -421 97 -419
rect 100 -415 101 -413
rect 100 -421 101 -419
rect 107 -415 108 -413
rect 107 -421 108 -419
rect 114 -415 115 -413
rect 114 -421 115 -419
rect 121 -415 122 -413
rect 124 -415 125 -413
rect 121 -421 122 -419
rect 124 -421 125 -419
rect 128 -415 129 -413
rect 128 -421 129 -419
rect 135 -415 136 -413
rect 135 -421 136 -419
rect 142 -415 143 -413
rect 142 -421 143 -419
rect 149 -415 150 -413
rect 149 -421 150 -419
rect 156 -415 157 -413
rect 159 -415 160 -413
rect 156 -421 157 -419
rect 159 -421 160 -419
rect 163 -415 164 -413
rect 163 -421 164 -419
rect 170 -415 171 -413
rect 170 -421 171 -419
rect 177 -415 178 -413
rect 177 -421 178 -419
rect 184 -415 185 -413
rect 184 -421 185 -419
rect 187 -421 188 -419
rect 191 -415 192 -413
rect 194 -415 195 -413
rect 191 -421 192 -419
rect 198 -415 199 -413
rect 198 -421 199 -419
rect 205 -415 206 -413
rect 205 -421 206 -419
rect 212 -415 213 -413
rect 212 -421 213 -419
rect 219 -415 220 -413
rect 219 -421 220 -419
rect 226 -415 227 -413
rect 226 -421 227 -419
rect 233 -415 234 -413
rect 233 -421 234 -419
rect 240 -415 241 -413
rect 243 -415 244 -413
rect 240 -421 241 -419
rect 243 -421 244 -419
rect 247 -415 248 -413
rect 247 -421 248 -419
rect 254 -415 255 -413
rect 254 -421 255 -419
rect 261 -415 262 -413
rect 261 -421 262 -419
rect 268 -415 269 -413
rect 268 -421 269 -419
rect 275 -415 276 -413
rect 275 -421 276 -419
rect 282 -415 283 -413
rect 282 -421 283 -419
rect 289 -415 290 -413
rect 289 -421 290 -419
rect 296 -415 297 -413
rect 296 -421 297 -419
rect 303 -415 304 -413
rect 303 -421 304 -419
rect 310 -415 311 -413
rect 310 -421 311 -419
rect 317 -415 318 -413
rect 317 -421 318 -419
rect 324 -415 325 -413
rect 324 -421 325 -419
rect 331 -415 332 -413
rect 331 -421 332 -419
rect 338 -415 339 -413
rect 338 -421 339 -419
rect 345 -415 346 -413
rect 345 -421 346 -419
rect 352 -415 353 -413
rect 355 -415 356 -413
rect 359 -415 360 -413
rect 362 -415 363 -413
rect 359 -421 360 -419
rect 362 -421 363 -419
rect 366 -415 367 -413
rect 366 -421 367 -419
rect 373 -415 374 -413
rect 373 -421 374 -419
rect 380 -415 381 -413
rect 380 -421 381 -419
rect 387 -415 388 -413
rect 387 -421 388 -419
rect 394 -415 395 -413
rect 397 -415 398 -413
rect 394 -421 395 -419
rect 397 -421 398 -419
rect 401 -415 402 -413
rect 401 -421 402 -419
rect 408 -415 409 -413
rect 411 -415 412 -413
rect 408 -421 409 -419
rect 411 -421 412 -419
rect 415 -415 416 -413
rect 415 -421 416 -419
rect 422 -415 423 -413
rect 422 -421 423 -419
rect 429 -415 430 -413
rect 432 -415 433 -413
rect 429 -421 430 -419
rect 432 -421 433 -419
rect 436 -415 437 -413
rect 436 -421 437 -419
rect 443 -415 444 -413
rect 443 -421 444 -419
rect 450 -415 451 -413
rect 450 -421 451 -419
rect 457 -415 458 -413
rect 460 -415 461 -413
rect 457 -421 458 -419
rect 460 -421 461 -419
rect 464 -415 465 -413
rect 467 -415 468 -413
rect 464 -421 465 -419
rect 467 -421 468 -419
rect 471 -415 472 -413
rect 471 -421 472 -419
rect 478 -415 479 -413
rect 478 -421 479 -419
rect 485 -415 486 -413
rect 485 -421 486 -419
rect 492 -415 493 -413
rect 492 -421 493 -419
rect 499 -415 500 -413
rect 499 -421 500 -419
rect 506 -415 507 -413
rect 506 -421 507 -419
rect 513 -415 514 -413
rect 516 -415 517 -413
rect 516 -421 517 -419
rect 520 -415 521 -413
rect 520 -421 521 -419
rect 527 -415 528 -413
rect 530 -415 531 -413
rect 527 -421 528 -419
rect 530 -421 531 -419
rect 534 -415 535 -413
rect 534 -421 535 -419
rect 541 -415 542 -413
rect 541 -421 542 -419
rect 551 -415 552 -413
rect 548 -421 549 -419
rect 551 -421 552 -419
rect 555 -415 556 -413
rect 555 -421 556 -419
rect 562 -415 563 -413
rect 562 -421 563 -419
rect 569 -415 570 -413
rect 569 -421 570 -419
rect 576 -415 577 -413
rect 576 -421 577 -419
rect 583 -415 584 -413
rect 583 -421 584 -419
rect 590 -415 591 -413
rect 590 -421 591 -419
rect 597 -415 598 -413
rect 597 -421 598 -419
rect 604 -415 605 -413
rect 604 -421 605 -419
rect 611 -415 612 -413
rect 611 -421 612 -419
rect 618 -415 619 -413
rect 621 -415 622 -413
rect 618 -421 619 -419
rect 621 -421 622 -419
rect 625 -415 626 -413
rect 625 -421 626 -419
rect 632 -415 633 -413
rect 632 -421 633 -419
rect 639 -415 640 -413
rect 639 -421 640 -419
rect 646 -415 647 -413
rect 646 -421 647 -419
rect 653 -415 654 -413
rect 653 -421 654 -419
rect 660 -415 661 -413
rect 660 -421 661 -419
rect 667 -415 668 -413
rect 667 -421 668 -419
rect 674 -415 675 -413
rect 674 -421 675 -419
rect 681 -415 682 -413
rect 681 -421 682 -419
rect 688 -415 689 -413
rect 688 -421 689 -419
rect 695 -415 696 -413
rect 695 -421 696 -419
rect 702 -415 703 -413
rect 702 -421 703 -419
rect 709 -415 710 -413
rect 709 -421 710 -419
rect 716 -415 717 -413
rect 716 -421 717 -419
rect 723 -415 724 -413
rect 723 -421 724 -419
rect 730 -415 731 -413
rect 730 -421 731 -419
rect 737 -415 738 -413
rect 737 -421 738 -419
rect 744 -415 745 -413
rect 744 -421 745 -419
rect 751 -415 752 -413
rect 751 -421 752 -419
rect 758 -415 759 -413
rect 758 -421 759 -419
rect 765 -415 766 -413
rect 765 -421 766 -419
rect 772 -415 773 -413
rect 772 -421 773 -419
rect 779 -415 780 -413
rect 779 -421 780 -419
rect 786 -415 787 -413
rect 786 -421 787 -419
rect 793 -415 794 -413
rect 793 -421 794 -419
rect 800 -415 801 -413
rect 800 -421 801 -419
rect 807 -415 808 -413
rect 807 -421 808 -419
rect 814 -415 815 -413
rect 814 -421 815 -419
rect 821 -415 822 -413
rect 821 -421 822 -419
rect 828 -415 829 -413
rect 828 -421 829 -419
rect 835 -415 836 -413
rect 835 -421 836 -419
rect 842 -415 843 -413
rect 842 -421 843 -419
rect 849 -415 850 -413
rect 849 -421 850 -419
rect 856 -415 857 -413
rect 856 -421 857 -419
rect 863 -415 864 -413
rect 863 -421 864 -419
rect 870 -415 871 -413
rect 870 -421 871 -419
rect 877 -415 878 -413
rect 877 -421 878 -419
rect 884 -415 885 -413
rect 884 -421 885 -419
rect 891 -415 892 -413
rect 891 -421 892 -419
rect 898 -415 899 -413
rect 898 -421 899 -419
rect 905 -415 906 -413
rect 905 -421 906 -419
rect 912 -415 913 -413
rect 912 -421 913 -419
rect 919 -415 920 -413
rect 919 -421 920 -419
rect 926 -415 927 -413
rect 926 -421 927 -419
rect 933 -415 934 -413
rect 933 -421 934 -419
rect 940 -415 941 -413
rect 940 -421 941 -419
rect 947 -415 948 -413
rect 947 -421 948 -419
rect 954 -415 955 -413
rect 954 -421 955 -419
rect 961 -415 962 -413
rect 961 -421 962 -419
rect 968 -415 969 -413
rect 968 -421 969 -419
rect 975 -415 976 -413
rect 975 -421 976 -419
rect 982 -415 983 -413
rect 982 -421 983 -419
rect 989 -415 990 -413
rect 989 -421 990 -419
rect 996 -415 997 -413
rect 996 -421 997 -419
rect 1003 -415 1004 -413
rect 1003 -421 1004 -419
rect 1024 -415 1025 -413
rect 1024 -421 1025 -419
rect 2 -510 3 -508
rect 2 -516 3 -514
rect 9 -510 10 -508
rect 9 -516 10 -514
rect 16 -510 17 -508
rect 16 -516 17 -514
rect 23 -510 24 -508
rect 23 -516 24 -514
rect 30 -510 31 -508
rect 30 -516 31 -514
rect 37 -510 38 -508
rect 37 -516 38 -514
rect 44 -510 45 -508
rect 44 -516 45 -514
rect 51 -510 52 -508
rect 51 -516 52 -514
rect 58 -510 59 -508
rect 58 -516 59 -514
rect 65 -510 66 -508
rect 65 -516 66 -514
rect 72 -510 73 -508
rect 72 -516 73 -514
rect 79 -510 80 -508
rect 79 -516 80 -514
rect 86 -510 87 -508
rect 86 -516 87 -514
rect 93 -510 94 -508
rect 96 -510 97 -508
rect 93 -516 94 -514
rect 100 -510 101 -508
rect 100 -516 101 -514
rect 107 -510 108 -508
rect 107 -516 108 -514
rect 114 -510 115 -508
rect 114 -516 115 -514
rect 121 -510 122 -508
rect 121 -516 122 -514
rect 128 -510 129 -508
rect 131 -510 132 -508
rect 128 -516 129 -514
rect 131 -516 132 -514
rect 138 -510 139 -508
rect 135 -516 136 -514
rect 138 -516 139 -514
rect 145 -516 146 -514
rect 152 -510 153 -508
rect 152 -516 153 -514
rect 156 -510 157 -508
rect 156 -516 157 -514
rect 159 -516 160 -514
rect 163 -510 164 -508
rect 163 -516 164 -514
rect 170 -510 171 -508
rect 170 -516 171 -514
rect 177 -510 178 -508
rect 177 -516 178 -514
rect 184 -510 185 -508
rect 184 -516 185 -514
rect 191 -510 192 -508
rect 191 -516 192 -514
rect 198 -510 199 -508
rect 198 -516 199 -514
rect 205 -510 206 -508
rect 205 -516 206 -514
rect 212 -510 213 -508
rect 212 -516 213 -514
rect 219 -510 220 -508
rect 219 -516 220 -514
rect 226 -510 227 -508
rect 226 -516 227 -514
rect 233 -510 234 -508
rect 233 -516 234 -514
rect 240 -510 241 -508
rect 240 -516 241 -514
rect 247 -510 248 -508
rect 250 -510 251 -508
rect 247 -516 248 -514
rect 250 -516 251 -514
rect 254 -510 255 -508
rect 254 -516 255 -514
rect 261 -510 262 -508
rect 261 -516 262 -514
rect 268 -510 269 -508
rect 268 -516 269 -514
rect 275 -510 276 -508
rect 275 -516 276 -514
rect 282 -510 283 -508
rect 282 -516 283 -514
rect 289 -510 290 -508
rect 289 -516 290 -514
rect 296 -510 297 -508
rect 296 -516 297 -514
rect 303 -510 304 -508
rect 303 -516 304 -514
rect 310 -510 311 -508
rect 310 -516 311 -514
rect 317 -510 318 -508
rect 317 -516 318 -514
rect 324 -510 325 -508
rect 327 -510 328 -508
rect 331 -510 332 -508
rect 331 -516 332 -514
rect 338 -510 339 -508
rect 338 -516 339 -514
rect 345 -510 346 -508
rect 345 -516 346 -514
rect 352 -510 353 -508
rect 352 -516 353 -514
rect 359 -510 360 -508
rect 359 -516 360 -514
rect 366 -510 367 -508
rect 366 -516 367 -514
rect 373 -510 374 -508
rect 373 -516 374 -514
rect 380 -510 381 -508
rect 380 -516 381 -514
rect 387 -510 388 -508
rect 390 -510 391 -508
rect 387 -516 388 -514
rect 394 -510 395 -508
rect 397 -510 398 -508
rect 394 -516 395 -514
rect 401 -510 402 -508
rect 401 -516 402 -514
rect 408 -510 409 -508
rect 411 -510 412 -508
rect 411 -516 412 -514
rect 415 -510 416 -508
rect 415 -516 416 -514
rect 422 -510 423 -508
rect 422 -516 423 -514
rect 429 -510 430 -508
rect 429 -516 430 -514
rect 436 -510 437 -508
rect 436 -516 437 -514
rect 443 -510 444 -508
rect 446 -510 447 -508
rect 446 -516 447 -514
rect 450 -510 451 -508
rect 450 -516 451 -514
rect 457 -510 458 -508
rect 457 -516 458 -514
rect 464 -510 465 -508
rect 464 -516 465 -514
rect 471 -510 472 -508
rect 471 -516 472 -514
rect 478 -510 479 -508
rect 481 -510 482 -508
rect 478 -516 479 -514
rect 481 -516 482 -514
rect 485 -510 486 -508
rect 485 -516 486 -514
rect 492 -510 493 -508
rect 492 -516 493 -514
rect 499 -510 500 -508
rect 499 -516 500 -514
rect 506 -510 507 -508
rect 509 -510 510 -508
rect 506 -516 507 -514
rect 509 -516 510 -514
rect 513 -510 514 -508
rect 513 -516 514 -514
rect 520 -510 521 -508
rect 523 -510 524 -508
rect 520 -516 521 -514
rect 523 -516 524 -514
rect 527 -510 528 -508
rect 527 -516 528 -514
rect 534 -510 535 -508
rect 534 -516 535 -514
rect 541 -510 542 -508
rect 541 -516 542 -514
rect 548 -510 549 -508
rect 548 -516 549 -514
rect 555 -510 556 -508
rect 555 -516 556 -514
rect 562 -510 563 -508
rect 565 -510 566 -508
rect 562 -516 563 -514
rect 565 -516 566 -514
rect 569 -510 570 -508
rect 572 -510 573 -508
rect 569 -516 570 -514
rect 572 -516 573 -514
rect 576 -510 577 -508
rect 579 -510 580 -508
rect 576 -516 577 -514
rect 579 -516 580 -514
rect 583 -510 584 -508
rect 583 -516 584 -514
rect 590 -510 591 -508
rect 590 -516 591 -514
rect 597 -510 598 -508
rect 597 -516 598 -514
rect 604 -510 605 -508
rect 607 -510 608 -508
rect 604 -516 605 -514
rect 607 -516 608 -514
rect 611 -510 612 -508
rect 611 -516 612 -514
rect 618 -510 619 -508
rect 618 -516 619 -514
rect 625 -510 626 -508
rect 625 -516 626 -514
rect 632 -510 633 -508
rect 632 -516 633 -514
rect 639 -510 640 -508
rect 639 -516 640 -514
rect 649 -510 650 -508
rect 646 -516 647 -514
rect 649 -516 650 -514
rect 653 -510 654 -508
rect 653 -516 654 -514
rect 660 -510 661 -508
rect 660 -516 661 -514
rect 667 -510 668 -508
rect 670 -510 671 -508
rect 667 -516 668 -514
rect 670 -516 671 -514
rect 674 -510 675 -508
rect 674 -516 675 -514
rect 681 -510 682 -508
rect 681 -516 682 -514
rect 688 -510 689 -508
rect 688 -516 689 -514
rect 695 -510 696 -508
rect 695 -516 696 -514
rect 702 -510 703 -508
rect 702 -516 703 -514
rect 709 -510 710 -508
rect 709 -516 710 -514
rect 716 -510 717 -508
rect 716 -516 717 -514
rect 723 -510 724 -508
rect 723 -516 724 -514
rect 730 -510 731 -508
rect 730 -516 731 -514
rect 737 -510 738 -508
rect 737 -516 738 -514
rect 744 -510 745 -508
rect 744 -516 745 -514
rect 751 -510 752 -508
rect 751 -516 752 -514
rect 754 -516 755 -514
rect 758 -510 759 -508
rect 758 -516 759 -514
rect 765 -510 766 -508
rect 765 -516 766 -514
rect 772 -510 773 -508
rect 772 -516 773 -514
rect 779 -510 780 -508
rect 779 -516 780 -514
rect 786 -510 787 -508
rect 786 -516 787 -514
rect 793 -510 794 -508
rect 793 -516 794 -514
rect 800 -510 801 -508
rect 800 -516 801 -514
rect 807 -510 808 -508
rect 807 -516 808 -514
rect 814 -510 815 -508
rect 814 -516 815 -514
rect 821 -510 822 -508
rect 821 -516 822 -514
rect 828 -510 829 -508
rect 828 -516 829 -514
rect 835 -510 836 -508
rect 835 -516 836 -514
rect 842 -510 843 -508
rect 842 -516 843 -514
rect 849 -510 850 -508
rect 849 -516 850 -514
rect 856 -510 857 -508
rect 856 -516 857 -514
rect 863 -510 864 -508
rect 863 -516 864 -514
rect 870 -510 871 -508
rect 870 -516 871 -514
rect 877 -510 878 -508
rect 877 -516 878 -514
rect 884 -510 885 -508
rect 884 -516 885 -514
rect 891 -510 892 -508
rect 891 -516 892 -514
rect 898 -510 899 -508
rect 898 -516 899 -514
rect 905 -510 906 -508
rect 905 -516 906 -514
rect 912 -510 913 -508
rect 912 -516 913 -514
rect 919 -510 920 -508
rect 919 -516 920 -514
rect 926 -510 927 -508
rect 926 -516 927 -514
rect 933 -510 934 -508
rect 933 -516 934 -514
rect 940 -510 941 -508
rect 940 -516 941 -514
rect 947 -510 948 -508
rect 947 -516 948 -514
rect 954 -510 955 -508
rect 954 -516 955 -514
rect 961 -510 962 -508
rect 961 -516 962 -514
rect 968 -510 969 -508
rect 968 -516 969 -514
rect 975 -510 976 -508
rect 975 -516 976 -514
rect 982 -510 983 -508
rect 982 -516 983 -514
rect 989 -510 990 -508
rect 989 -516 990 -514
rect 996 -510 997 -508
rect 996 -516 997 -514
rect 1003 -510 1004 -508
rect 1003 -516 1004 -514
rect 1010 -510 1011 -508
rect 1010 -516 1011 -514
rect 1017 -510 1018 -508
rect 1017 -516 1018 -514
rect 1024 -510 1025 -508
rect 1024 -516 1025 -514
rect 1031 -510 1032 -508
rect 1031 -516 1032 -514
rect 1038 -510 1039 -508
rect 1038 -516 1039 -514
rect 1045 -510 1046 -508
rect 1045 -516 1046 -514
rect 1052 -510 1053 -508
rect 1052 -516 1053 -514
rect 1059 -510 1060 -508
rect 1059 -516 1060 -514
rect 1066 -510 1067 -508
rect 1066 -516 1067 -514
rect 1073 -510 1074 -508
rect 1073 -516 1074 -514
rect 1080 -510 1081 -508
rect 1080 -516 1081 -514
rect 1087 -510 1088 -508
rect 1087 -516 1088 -514
rect 1094 -510 1095 -508
rect 1094 -516 1095 -514
rect 1101 -510 1102 -508
rect 1101 -516 1102 -514
rect 1108 -510 1109 -508
rect 1108 -516 1109 -514
rect 1115 -510 1116 -508
rect 1115 -516 1116 -514
rect 1122 -510 1123 -508
rect 1122 -516 1123 -514
rect 2 -609 3 -607
rect 2 -615 3 -613
rect 9 -609 10 -607
rect 9 -615 10 -613
rect 16 -609 17 -607
rect 16 -615 17 -613
rect 23 -609 24 -607
rect 23 -615 24 -613
rect 30 -609 31 -607
rect 30 -615 31 -613
rect 37 -609 38 -607
rect 40 -615 41 -613
rect 44 -609 45 -607
rect 44 -615 45 -613
rect 51 -609 52 -607
rect 51 -615 52 -613
rect 58 -609 59 -607
rect 58 -615 59 -613
rect 61 -615 62 -613
rect 65 -609 66 -607
rect 65 -615 66 -613
rect 68 -615 69 -613
rect 72 -609 73 -607
rect 75 -609 76 -607
rect 72 -615 73 -613
rect 75 -615 76 -613
rect 79 -609 80 -607
rect 79 -615 80 -613
rect 86 -609 87 -607
rect 86 -615 87 -613
rect 93 -609 94 -607
rect 93 -615 94 -613
rect 100 -609 101 -607
rect 100 -615 101 -613
rect 107 -609 108 -607
rect 107 -615 108 -613
rect 114 -609 115 -607
rect 114 -615 115 -613
rect 121 -609 122 -607
rect 121 -615 122 -613
rect 128 -609 129 -607
rect 128 -615 129 -613
rect 135 -609 136 -607
rect 135 -615 136 -613
rect 142 -609 143 -607
rect 145 -609 146 -607
rect 142 -615 143 -613
rect 145 -615 146 -613
rect 149 -609 150 -607
rect 149 -615 150 -613
rect 156 -609 157 -607
rect 156 -615 157 -613
rect 163 -609 164 -607
rect 163 -615 164 -613
rect 170 -609 171 -607
rect 170 -615 171 -613
rect 177 -609 178 -607
rect 177 -615 178 -613
rect 184 -609 185 -607
rect 187 -609 188 -607
rect 184 -615 185 -613
rect 187 -615 188 -613
rect 191 -609 192 -607
rect 191 -615 192 -613
rect 198 -609 199 -607
rect 198 -615 199 -613
rect 205 -609 206 -607
rect 205 -615 206 -613
rect 212 -609 213 -607
rect 212 -615 213 -613
rect 219 -609 220 -607
rect 219 -615 220 -613
rect 226 -609 227 -607
rect 226 -615 227 -613
rect 233 -609 234 -607
rect 233 -615 234 -613
rect 240 -609 241 -607
rect 240 -615 241 -613
rect 247 -609 248 -607
rect 247 -615 248 -613
rect 254 -609 255 -607
rect 254 -615 255 -613
rect 261 -609 262 -607
rect 261 -615 262 -613
rect 268 -609 269 -607
rect 268 -615 269 -613
rect 275 -609 276 -607
rect 278 -609 279 -607
rect 275 -615 276 -613
rect 278 -615 279 -613
rect 282 -609 283 -607
rect 282 -615 283 -613
rect 289 -609 290 -607
rect 289 -615 290 -613
rect 296 -609 297 -607
rect 296 -615 297 -613
rect 303 -609 304 -607
rect 303 -615 304 -613
rect 310 -609 311 -607
rect 310 -615 311 -613
rect 317 -609 318 -607
rect 317 -615 318 -613
rect 324 -609 325 -607
rect 324 -615 325 -613
rect 331 -609 332 -607
rect 334 -609 335 -607
rect 331 -615 332 -613
rect 334 -615 335 -613
rect 338 -609 339 -607
rect 338 -615 339 -613
rect 345 -609 346 -607
rect 345 -615 346 -613
rect 352 -609 353 -607
rect 352 -615 353 -613
rect 359 -609 360 -607
rect 359 -615 360 -613
rect 366 -609 367 -607
rect 366 -615 367 -613
rect 373 -609 374 -607
rect 373 -615 374 -613
rect 380 -609 381 -607
rect 383 -609 384 -607
rect 380 -615 381 -613
rect 383 -615 384 -613
rect 387 -609 388 -607
rect 390 -609 391 -607
rect 387 -615 388 -613
rect 390 -615 391 -613
rect 394 -609 395 -607
rect 394 -615 395 -613
rect 401 -609 402 -607
rect 404 -609 405 -607
rect 404 -615 405 -613
rect 408 -609 409 -607
rect 408 -615 409 -613
rect 415 -609 416 -607
rect 418 -615 419 -613
rect 422 -609 423 -607
rect 425 -609 426 -607
rect 422 -615 423 -613
rect 425 -615 426 -613
rect 429 -609 430 -607
rect 429 -615 430 -613
rect 436 -609 437 -607
rect 436 -615 437 -613
rect 443 -609 444 -607
rect 443 -615 444 -613
rect 450 -609 451 -607
rect 453 -609 454 -607
rect 450 -615 451 -613
rect 453 -615 454 -613
rect 457 -609 458 -607
rect 460 -609 461 -607
rect 457 -615 458 -613
rect 460 -615 461 -613
rect 464 -609 465 -607
rect 467 -609 468 -607
rect 464 -615 465 -613
rect 467 -615 468 -613
rect 471 -609 472 -607
rect 471 -615 472 -613
rect 478 -609 479 -607
rect 478 -615 479 -613
rect 485 -609 486 -607
rect 485 -615 486 -613
rect 492 -609 493 -607
rect 492 -615 493 -613
rect 499 -609 500 -607
rect 499 -615 500 -613
rect 506 -609 507 -607
rect 506 -615 507 -613
rect 513 -609 514 -607
rect 513 -615 514 -613
rect 520 -609 521 -607
rect 523 -609 524 -607
rect 520 -615 521 -613
rect 523 -615 524 -613
rect 527 -609 528 -607
rect 527 -615 528 -613
rect 534 -609 535 -607
rect 534 -615 535 -613
rect 541 -609 542 -607
rect 544 -609 545 -607
rect 541 -615 542 -613
rect 544 -615 545 -613
rect 548 -609 549 -607
rect 551 -609 552 -607
rect 548 -615 549 -613
rect 551 -615 552 -613
rect 555 -609 556 -607
rect 555 -615 556 -613
rect 562 -609 563 -607
rect 565 -609 566 -607
rect 562 -615 563 -613
rect 565 -615 566 -613
rect 569 -609 570 -607
rect 569 -615 570 -613
rect 576 -609 577 -607
rect 576 -615 577 -613
rect 583 -609 584 -607
rect 583 -615 584 -613
rect 586 -615 587 -613
rect 590 -609 591 -607
rect 590 -615 591 -613
rect 597 -609 598 -607
rect 597 -615 598 -613
rect 604 -609 605 -607
rect 604 -615 605 -613
rect 611 -609 612 -607
rect 611 -615 612 -613
rect 618 -609 619 -607
rect 621 -609 622 -607
rect 618 -615 619 -613
rect 621 -615 622 -613
rect 625 -609 626 -607
rect 628 -609 629 -607
rect 625 -615 626 -613
rect 628 -615 629 -613
rect 632 -609 633 -607
rect 632 -615 633 -613
rect 639 -609 640 -607
rect 639 -615 640 -613
rect 646 -609 647 -607
rect 646 -615 647 -613
rect 653 -609 654 -607
rect 653 -615 654 -613
rect 660 -609 661 -607
rect 660 -615 661 -613
rect 667 -609 668 -607
rect 667 -615 668 -613
rect 674 -609 675 -607
rect 674 -615 675 -613
rect 681 -609 682 -607
rect 681 -615 682 -613
rect 688 -609 689 -607
rect 688 -615 689 -613
rect 695 -609 696 -607
rect 695 -615 696 -613
rect 702 -609 703 -607
rect 702 -615 703 -613
rect 709 -609 710 -607
rect 709 -615 710 -613
rect 716 -609 717 -607
rect 716 -615 717 -613
rect 723 -609 724 -607
rect 723 -615 724 -613
rect 730 -609 731 -607
rect 730 -615 731 -613
rect 737 -609 738 -607
rect 737 -615 738 -613
rect 744 -609 745 -607
rect 744 -615 745 -613
rect 751 -609 752 -607
rect 751 -615 752 -613
rect 758 -609 759 -607
rect 758 -615 759 -613
rect 765 -609 766 -607
rect 765 -615 766 -613
rect 772 -609 773 -607
rect 772 -615 773 -613
rect 779 -609 780 -607
rect 779 -615 780 -613
rect 786 -609 787 -607
rect 786 -615 787 -613
rect 793 -609 794 -607
rect 793 -615 794 -613
rect 800 -609 801 -607
rect 800 -615 801 -613
rect 807 -609 808 -607
rect 807 -615 808 -613
rect 814 -609 815 -607
rect 814 -615 815 -613
rect 821 -609 822 -607
rect 821 -615 822 -613
rect 828 -609 829 -607
rect 828 -615 829 -613
rect 835 -609 836 -607
rect 835 -615 836 -613
rect 842 -609 843 -607
rect 842 -615 843 -613
rect 849 -609 850 -607
rect 849 -615 850 -613
rect 856 -609 857 -607
rect 856 -615 857 -613
rect 863 -609 864 -607
rect 863 -615 864 -613
rect 870 -609 871 -607
rect 870 -615 871 -613
rect 877 -609 878 -607
rect 877 -615 878 -613
rect 884 -609 885 -607
rect 884 -615 885 -613
rect 891 -609 892 -607
rect 891 -615 892 -613
rect 898 -609 899 -607
rect 898 -615 899 -613
rect 905 -609 906 -607
rect 905 -615 906 -613
rect 912 -609 913 -607
rect 912 -615 913 -613
rect 919 -609 920 -607
rect 919 -615 920 -613
rect 926 -609 927 -607
rect 926 -615 927 -613
rect 933 -609 934 -607
rect 933 -615 934 -613
rect 940 -609 941 -607
rect 940 -615 941 -613
rect 947 -609 948 -607
rect 947 -615 948 -613
rect 954 -609 955 -607
rect 954 -615 955 -613
rect 961 -609 962 -607
rect 961 -615 962 -613
rect 968 -609 969 -607
rect 968 -615 969 -613
rect 975 -609 976 -607
rect 975 -615 976 -613
rect 982 -609 983 -607
rect 982 -615 983 -613
rect 989 -609 990 -607
rect 989 -615 990 -613
rect 996 -609 997 -607
rect 996 -615 997 -613
rect 1003 -609 1004 -607
rect 1003 -615 1004 -613
rect 1010 -609 1011 -607
rect 1010 -615 1011 -613
rect 1017 -609 1018 -607
rect 1017 -615 1018 -613
rect 1024 -609 1025 -607
rect 1024 -615 1025 -613
rect 1031 -609 1032 -607
rect 1031 -615 1032 -613
rect 1038 -609 1039 -607
rect 1038 -615 1039 -613
rect 1045 -609 1046 -607
rect 1045 -615 1046 -613
rect 1052 -609 1053 -607
rect 1052 -615 1053 -613
rect 1059 -609 1060 -607
rect 1059 -615 1060 -613
rect 1066 -609 1067 -607
rect 1066 -615 1067 -613
rect 1073 -609 1074 -607
rect 1073 -615 1074 -613
rect 1080 -609 1081 -607
rect 1083 -615 1084 -613
rect 1087 -609 1088 -607
rect 1087 -615 1088 -613
rect 2 -718 3 -716
rect 2 -724 3 -722
rect 9 -718 10 -716
rect 9 -724 10 -722
rect 16 -718 17 -716
rect 16 -724 17 -722
rect 23 -718 24 -716
rect 23 -724 24 -722
rect 30 -718 31 -716
rect 30 -724 31 -722
rect 37 -718 38 -716
rect 37 -724 38 -722
rect 44 -718 45 -716
rect 47 -718 48 -716
rect 44 -724 45 -722
rect 51 -718 52 -716
rect 51 -724 52 -722
rect 58 -718 59 -716
rect 61 -718 62 -716
rect 58 -724 59 -722
rect 61 -724 62 -722
rect 65 -718 66 -716
rect 65 -724 66 -722
rect 72 -718 73 -716
rect 72 -724 73 -722
rect 79 -718 80 -716
rect 79 -724 80 -722
rect 86 -718 87 -716
rect 89 -718 90 -716
rect 89 -724 90 -722
rect 93 -718 94 -716
rect 93 -724 94 -722
rect 100 -718 101 -716
rect 100 -724 101 -722
rect 107 -718 108 -716
rect 110 -718 111 -716
rect 107 -724 108 -722
rect 110 -724 111 -722
rect 114 -718 115 -716
rect 114 -724 115 -722
rect 121 -718 122 -716
rect 121 -724 122 -722
rect 128 -718 129 -716
rect 128 -724 129 -722
rect 135 -718 136 -716
rect 135 -724 136 -722
rect 142 -718 143 -716
rect 142 -724 143 -722
rect 149 -718 150 -716
rect 149 -724 150 -722
rect 156 -718 157 -716
rect 156 -724 157 -722
rect 163 -718 164 -716
rect 163 -724 164 -722
rect 170 -718 171 -716
rect 170 -724 171 -722
rect 177 -718 178 -716
rect 177 -724 178 -722
rect 184 -718 185 -716
rect 184 -724 185 -722
rect 191 -718 192 -716
rect 191 -724 192 -722
rect 194 -724 195 -722
rect 198 -718 199 -716
rect 198 -724 199 -722
rect 205 -718 206 -716
rect 205 -724 206 -722
rect 212 -718 213 -716
rect 212 -724 213 -722
rect 219 -718 220 -716
rect 219 -724 220 -722
rect 226 -718 227 -716
rect 229 -718 230 -716
rect 226 -724 227 -722
rect 233 -718 234 -716
rect 236 -718 237 -716
rect 233 -724 234 -722
rect 240 -718 241 -716
rect 240 -724 241 -722
rect 247 -718 248 -716
rect 247 -724 248 -722
rect 254 -718 255 -716
rect 254 -724 255 -722
rect 261 -718 262 -716
rect 261 -724 262 -722
rect 268 -718 269 -716
rect 268 -724 269 -722
rect 275 -718 276 -716
rect 275 -724 276 -722
rect 282 -718 283 -716
rect 282 -724 283 -722
rect 289 -718 290 -716
rect 289 -724 290 -722
rect 296 -718 297 -716
rect 296 -724 297 -722
rect 303 -718 304 -716
rect 303 -724 304 -722
rect 310 -718 311 -716
rect 310 -724 311 -722
rect 317 -718 318 -716
rect 317 -724 318 -722
rect 324 -718 325 -716
rect 324 -724 325 -722
rect 331 -718 332 -716
rect 331 -724 332 -722
rect 338 -718 339 -716
rect 338 -724 339 -722
rect 345 -718 346 -716
rect 345 -724 346 -722
rect 352 -718 353 -716
rect 352 -724 353 -722
rect 359 -718 360 -716
rect 359 -724 360 -722
rect 366 -718 367 -716
rect 369 -718 370 -716
rect 366 -724 367 -722
rect 369 -724 370 -722
rect 373 -718 374 -716
rect 373 -724 374 -722
rect 380 -718 381 -716
rect 383 -718 384 -716
rect 380 -724 381 -722
rect 383 -724 384 -722
rect 387 -718 388 -716
rect 387 -724 388 -722
rect 390 -724 391 -722
rect 394 -718 395 -716
rect 394 -724 395 -722
rect 404 -718 405 -716
rect 404 -724 405 -722
rect 408 -718 409 -716
rect 408 -724 409 -722
rect 415 -718 416 -716
rect 418 -718 419 -716
rect 415 -724 416 -722
rect 422 -718 423 -716
rect 422 -724 423 -722
rect 429 -718 430 -716
rect 432 -718 433 -716
rect 429 -724 430 -722
rect 432 -724 433 -722
rect 436 -718 437 -716
rect 436 -724 437 -722
rect 443 -718 444 -716
rect 446 -718 447 -716
rect 443 -724 444 -722
rect 446 -724 447 -722
rect 450 -718 451 -716
rect 450 -724 451 -722
rect 457 -718 458 -716
rect 457 -724 458 -722
rect 464 -718 465 -716
rect 464 -724 465 -722
rect 471 -718 472 -716
rect 471 -724 472 -722
rect 478 -718 479 -716
rect 478 -724 479 -722
rect 485 -718 486 -716
rect 485 -724 486 -722
rect 492 -718 493 -716
rect 492 -724 493 -722
rect 499 -718 500 -716
rect 502 -718 503 -716
rect 499 -724 500 -722
rect 502 -724 503 -722
rect 506 -718 507 -716
rect 506 -724 507 -722
rect 513 -718 514 -716
rect 513 -724 514 -722
rect 520 -718 521 -716
rect 520 -724 521 -722
rect 527 -718 528 -716
rect 527 -724 528 -722
rect 534 -718 535 -716
rect 534 -724 535 -722
rect 541 -718 542 -716
rect 541 -724 542 -722
rect 548 -718 549 -716
rect 548 -724 549 -722
rect 555 -718 556 -716
rect 558 -718 559 -716
rect 558 -724 559 -722
rect 562 -718 563 -716
rect 565 -718 566 -716
rect 562 -724 563 -722
rect 565 -724 566 -722
rect 569 -718 570 -716
rect 569 -724 570 -722
rect 576 -718 577 -716
rect 576 -724 577 -722
rect 583 -718 584 -716
rect 586 -718 587 -716
rect 583 -724 584 -722
rect 586 -724 587 -722
rect 590 -718 591 -716
rect 590 -724 591 -722
rect 597 -718 598 -716
rect 597 -724 598 -722
rect 604 -718 605 -716
rect 604 -724 605 -722
rect 611 -718 612 -716
rect 611 -724 612 -722
rect 618 -718 619 -716
rect 618 -724 619 -722
rect 625 -718 626 -716
rect 625 -724 626 -722
rect 632 -718 633 -716
rect 635 -718 636 -716
rect 632 -724 633 -722
rect 635 -724 636 -722
rect 639 -718 640 -716
rect 639 -724 640 -722
rect 646 -718 647 -716
rect 649 -718 650 -716
rect 649 -724 650 -722
rect 653 -718 654 -716
rect 656 -718 657 -716
rect 653 -724 654 -722
rect 656 -724 657 -722
rect 660 -718 661 -716
rect 660 -724 661 -722
rect 667 -718 668 -716
rect 667 -724 668 -722
rect 674 -718 675 -716
rect 674 -724 675 -722
rect 681 -718 682 -716
rect 681 -724 682 -722
rect 688 -718 689 -716
rect 688 -724 689 -722
rect 695 -718 696 -716
rect 695 -724 696 -722
rect 702 -718 703 -716
rect 702 -724 703 -722
rect 709 -718 710 -716
rect 709 -724 710 -722
rect 716 -718 717 -716
rect 716 -724 717 -722
rect 723 -718 724 -716
rect 726 -718 727 -716
rect 723 -724 724 -722
rect 726 -724 727 -722
rect 730 -718 731 -716
rect 733 -718 734 -716
rect 730 -724 731 -722
rect 733 -724 734 -722
rect 737 -718 738 -716
rect 737 -724 738 -722
rect 744 -718 745 -716
rect 744 -724 745 -722
rect 751 -718 752 -716
rect 751 -724 752 -722
rect 758 -718 759 -716
rect 758 -724 759 -722
rect 765 -718 766 -716
rect 765 -724 766 -722
rect 772 -718 773 -716
rect 772 -724 773 -722
rect 779 -718 780 -716
rect 779 -724 780 -722
rect 786 -718 787 -716
rect 786 -724 787 -722
rect 793 -718 794 -716
rect 793 -724 794 -722
rect 800 -718 801 -716
rect 800 -724 801 -722
rect 810 -718 811 -716
rect 807 -724 808 -722
rect 814 -718 815 -716
rect 814 -724 815 -722
rect 821 -718 822 -716
rect 821 -724 822 -722
rect 828 -718 829 -716
rect 828 -724 829 -722
rect 835 -718 836 -716
rect 835 -724 836 -722
rect 842 -718 843 -716
rect 842 -724 843 -722
rect 849 -718 850 -716
rect 849 -724 850 -722
rect 856 -718 857 -716
rect 856 -724 857 -722
rect 863 -718 864 -716
rect 863 -724 864 -722
rect 870 -718 871 -716
rect 870 -724 871 -722
rect 877 -718 878 -716
rect 877 -724 878 -722
rect 884 -718 885 -716
rect 884 -724 885 -722
rect 891 -718 892 -716
rect 891 -724 892 -722
rect 898 -718 899 -716
rect 898 -724 899 -722
rect 905 -718 906 -716
rect 905 -724 906 -722
rect 912 -718 913 -716
rect 912 -724 913 -722
rect 919 -718 920 -716
rect 919 -724 920 -722
rect 926 -718 927 -716
rect 926 -724 927 -722
rect 933 -718 934 -716
rect 933 -724 934 -722
rect 940 -718 941 -716
rect 940 -724 941 -722
rect 947 -718 948 -716
rect 947 -724 948 -722
rect 954 -718 955 -716
rect 954 -724 955 -722
rect 961 -718 962 -716
rect 961 -724 962 -722
rect 968 -718 969 -716
rect 968 -724 969 -722
rect 975 -718 976 -716
rect 975 -724 976 -722
rect 982 -718 983 -716
rect 982 -724 983 -722
rect 989 -718 990 -716
rect 989 -724 990 -722
rect 996 -718 997 -716
rect 996 -724 997 -722
rect 1003 -718 1004 -716
rect 1003 -724 1004 -722
rect 1010 -718 1011 -716
rect 1010 -724 1011 -722
rect 1017 -718 1018 -716
rect 1017 -724 1018 -722
rect 1024 -718 1025 -716
rect 1024 -724 1025 -722
rect 1031 -718 1032 -716
rect 1031 -724 1032 -722
rect 1038 -718 1039 -716
rect 1038 -724 1039 -722
rect 1045 -718 1046 -716
rect 1045 -724 1046 -722
rect 1052 -718 1053 -716
rect 1052 -724 1053 -722
rect 1059 -718 1060 -716
rect 1059 -724 1060 -722
rect 1066 -718 1067 -716
rect 1066 -724 1067 -722
rect 1073 -718 1074 -716
rect 1073 -724 1074 -722
rect 1080 -718 1081 -716
rect 1080 -724 1081 -722
rect 1087 -718 1088 -716
rect 1087 -724 1088 -722
rect 1094 -718 1095 -716
rect 1094 -724 1095 -722
rect 1101 -718 1102 -716
rect 1101 -724 1102 -722
rect 1108 -718 1109 -716
rect 1108 -724 1109 -722
rect 1115 -718 1116 -716
rect 1115 -724 1116 -722
rect 1122 -718 1123 -716
rect 1122 -724 1123 -722
rect 1129 -718 1130 -716
rect 1129 -724 1130 -722
rect 1136 -718 1137 -716
rect 1136 -724 1137 -722
rect 1143 -718 1144 -716
rect 1143 -724 1144 -722
rect 1150 -718 1151 -716
rect 1150 -724 1151 -722
rect 1157 -718 1158 -716
rect 1157 -724 1158 -722
rect 1164 -718 1165 -716
rect 1164 -724 1165 -722
rect 1171 -718 1172 -716
rect 1171 -724 1172 -722
rect 1178 -718 1179 -716
rect 1178 -724 1179 -722
rect 1185 -718 1186 -716
rect 1185 -724 1186 -722
rect 1192 -718 1193 -716
rect 1192 -724 1193 -722
rect 1199 -718 1200 -716
rect 1199 -724 1200 -722
rect 1206 -718 1207 -716
rect 1206 -724 1207 -722
rect 1213 -718 1214 -716
rect 1216 -718 1217 -716
rect 1213 -724 1214 -722
rect 1360 -718 1361 -716
rect 1360 -724 1361 -722
rect 2 -835 3 -833
rect 2 -841 3 -839
rect 9 -835 10 -833
rect 9 -841 10 -839
rect 16 -835 17 -833
rect 16 -841 17 -839
rect 23 -841 24 -839
rect 26 -841 27 -839
rect 33 -835 34 -833
rect 30 -841 31 -839
rect 33 -841 34 -839
rect 37 -835 38 -833
rect 37 -841 38 -839
rect 44 -835 45 -833
rect 44 -841 45 -839
rect 51 -835 52 -833
rect 51 -841 52 -839
rect 58 -835 59 -833
rect 58 -841 59 -839
rect 65 -835 66 -833
rect 65 -841 66 -839
rect 72 -835 73 -833
rect 75 -835 76 -833
rect 72 -841 73 -839
rect 75 -841 76 -839
rect 79 -835 80 -833
rect 79 -841 80 -839
rect 86 -835 87 -833
rect 89 -835 90 -833
rect 86 -841 87 -839
rect 89 -841 90 -839
rect 93 -835 94 -833
rect 93 -841 94 -839
rect 100 -835 101 -833
rect 100 -841 101 -839
rect 107 -835 108 -833
rect 107 -841 108 -839
rect 114 -835 115 -833
rect 114 -841 115 -839
rect 121 -835 122 -833
rect 121 -841 122 -839
rect 128 -835 129 -833
rect 131 -835 132 -833
rect 131 -841 132 -839
rect 135 -835 136 -833
rect 135 -841 136 -839
rect 142 -835 143 -833
rect 142 -841 143 -839
rect 149 -835 150 -833
rect 149 -841 150 -839
rect 156 -835 157 -833
rect 156 -841 157 -839
rect 163 -835 164 -833
rect 163 -841 164 -839
rect 170 -835 171 -833
rect 170 -841 171 -839
rect 177 -835 178 -833
rect 180 -841 181 -839
rect 184 -835 185 -833
rect 184 -841 185 -839
rect 191 -835 192 -833
rect 191 -841 192 -839
rect 198 -835 199 -833
rect 198 -841 199 -839
rect 205 -835 206 -833
rect 205 -841 206 -839
rect 212 -835 213 -833
rect 212 -841 213 -839
rect 219 -835 220 -833
rect 219 -841 220 -839
rect 226 -835 227 -833
rect 226 -841 227 -839
rect 233 -835 234 -833
rect 233 -841 234 -839
rect 240 -835 241 -833
rect 240 -841 241 -839
rect 247 -835 248 -833
rect 247 -841 248 -839
rect 254 -835 255 -833
rect 254 -841 255 -839
rect 261 -835 262 -833
rect 261 -841 262 -839
rect 268 -835 269 -833
rect 268 -841 269 -839
rect 275 -835 276 -833
rect 275 -841 276 -839
rect 282 -835 283 -833
rect 282 -841 283 -839
rect 289 -835 290 -833
rect 289 -841 290 -839
rect 296 -835 297 -833
rect 299 -835 300 -833
rect 296 -841 297 -839
rect 299 -841 300 -839
rect 303 -835 304 -833
rect 303 -841 304 -839
rect 310 -835 311 -833
rect 310 -841 311 -839
rect 317 -835 318 -833
rect 317 -841 318 -839
rect 324 -835 325 -833
rect 324 -841 325 -839
rect 331 -835 332 -833
rect 331 -841 332 -839
rect 338 -835 339 -833
rect 338 -841 339 -839
rect 345 -835 346 -833
rect 345 -841 346 -839
rect 352 -835 353 -833
rect 352 -841 353 -839
rect 359 -835 360 -833
rect 359 -841 360 -839
rect 366 -835 367 -833
rect 366 -841 367 -839
rect 373 -835 374 -833
rect 373 -841 374 -839
rect 380 -835 381 -833
rect 380 -841 381 -839
rect 387 -835 388 -833
rect 390 -835 391 -833
rect 387 -841 388 -839
rect 390 -841 391 -839
rect 394 -835 395 -833
rect 397 -835 398 -833
rect 394 -841 395 -839
rect 397 -841 398 -839
rect 401 -835 402 -833
rect 404 -835 405 -833
rect 401 -841 402 -839
rect 404 -841 405 -839
rect 408 -835 409 -833
rect 408 -841 409 -839
rect 415 -835 416 -833
rect 415 -841 416 -839
rect 422 -835 423 -833
rect 422 -841 423 -839
rect 429 -835 430 -833
rect 432 -835 433 -833
rect 429 -841 430 -839
rect 432 -841 433 -839
rect 436 -841 437 -839
rect 439 -841 440 -839
rect 443 -835 444 -833
rect 443 -841 444 -839
rect 450 -835 451 -833
rect 450 -841 451 -839
rect 457 -835 458 -833
rect 457 -841 458 -839
rect 464 -835 465 -833
rect 464 -841 465 -839
rect 471 -835 472 -833
rect 471 -841 472 -839
rect 478 -835 479 -833
rect 478 -841 479 -839
rect 485 -835 486 -833
rect 485 -841 486 -839
rect 492 -835 493 -833
rect 495 -835 496 -833
rect 492 -841 493 -839
rect 495 -841 496 -839
rect 499 -835 500 -833
rect 499 -841 500 -839
rect 506 -835 507 -833
rect 509 -835 510 -833
rect 506 -841 507 -839
rect 509 -841 510 -839
rect 513 -835 514 -833
rect 516 -835 517 -833
rect 513 -841 514 -839
rect 516 -841 517 -839
rect 520 -835 521 -833
rect 523 -835 524 -833
rect 520 -841 521 -839
rect 523 -841 524 -839
rect 527 -835 528 -833
rect 527 -841 528 -839
rect 534 -835 535 -833
rect 534 -841 535 -839
rect 541 -835 542 -833
rect 541 -841 542 -839
rect 548 -835 549 -833
rect 548 -841 549 -839
rect 555 -835 556 -833
rect 555 -841 556 -839
rect 562 -835 563 -833
rect 565 -835 566 -833
rect 562 -841 563 -839
rect 565 -841 566 -839
rect 569 -835 570 -833
rect 572 -835 573 -833
rect 569 -841 570 -839
rect 572 -841 573 -839
rect 576 -835 577 -833
rect 576 -841 577 -839
rect 583 -835 584 -833
rect 586 -835 587 -833
rect 583 -841 584 -839
rect 586 -841 587 -839
rect 590 -835 591 -833
rect 590 -841 591 -839
rect 597 -835 598 -833
rect 597 -841 598 -839
rect 604 -835 605 -833
rect 604 -841 605 -839
rect 611 -835 612 -833
rect 611 -841 612 -839
rect 618 -835 619 -833
rect 621 -835 622 -833
rect 618 -841 619 -839
rect 625 -835 626 -833
rect 625 -841 626 -839
rect 632 -835 633 -833
rect 632 -841 633 -839
rect 639 -835 640 -833
rect 639 -841 640 -839
rect 646 -835 647 -833
rect 649 -835 650 -833
rect 646 -841 647 -839
rect 649 -841 650 -839
rect 653 -835 654 -833
rect 656 -835 657 -833
rect 653 -841 654 -839
rect 656 -841 657 -839
rect 660 -835 661 -833
rect 660 -841 661 -839
rect 667 -835 668 -833
rect 667 -841 668 -839
rect 674 -835 675 -833
rect 674 -841 675 -839
rect 681 -835 682 -833
rect 681 -841 682 -839
rect 688 -835 689 -833
rect 688 -841 689 -839
rect 695 -835 696 -833
rect 695 -841 696 -839
rect 702 -835 703 -833
rect 705 -835 706 -833
rect 702 -841 703 -839
rect 705 -841 706 -839
rect 709 -835 710 -833
rect 709 -841 710 -839
rect 716 -835 717 -833
rect 716 -841 717 -839
rect 723 -835 724 -833
rect 723 -841 724 -839
rect 730 -835 731 -833
rect 730 -841 731 -839
rect 737 -835 738 -833
rect 737 -841 738 -839
rect 744 -835 745 -833
rect 744 -841 745 -839
rect 751 -835 752 -833
rect 751 -841 752 -839
rect 758 -835 759 -833
rect 761 -835 762 -833
rect 758 -841 759 -839
rect 761 -841 762 -839
rect 765 -835 766 -833
rect 765 -841 766 -839
rect 772 -835 773 -833
rect 772 -841 773 -839
rect 775 -841 776 -839
rect 779 -835 780 -833
rect 779 -841 780 -839
rect 786 -835 787 -833
rect 786 -841 787 -839
rect 793 -835 794 -833
rect 793 -841 794 -839
rect 800 -835 801 -833
rect 800 -841 801 -839
rect 807 -835 808 -833
rect 807 -841 808 -839
rect 814 -835 815 -833
rect 814 -841 815 -839
rect 821 -835 822 -833
rect 821 -841 822 -839
rect 828 -835 829 -833
rect 828 -841 829 -839
rect 831 -841 832 -839
rect 835 -835 836 -833
rect 835 -841 836 -839
rect 842 -835 843 -833
rect 842 -841 843 -839
rect 849 -835 850 -833
rect 849 -841 850 -839
rect 856 -835 857 -833
rect 856 -841 857 -839
rect 863 -835 864 -833
rect 863 -841 864 -839
rect 870 -835 871 -833
rect 870 -841 871 -839
rect 877 -835 878 -833
rect 877 -841 878 -839
rect 884 -835 885 -833
rect 884 -841 885 -839
rect 891 -835 892 -833
rect 891 -841 892 -839
rect 898 -835 899 -833
rect 898 -841 899 -839
rect 905 -835 906 -833
rect 905 -841 906 -839
rect 912 -835 913 -833
rect 912 -841 913 -839
rect 919 -835 920 -833
rect 919 -841 920 -839
rect 926 -835 927 -833
rect 926 -841 927 -839
rect 933 -835 934 -833
rect 933 -841 934 -839
rect 940 -835 941 -833
rect 940 -841 941 -839
rect 947 -835 948 -833
rect 947 -841 948 -839
rect 954 -835 955 -833
rect 954 -841 955 -839
rect 961 -835 962 -833
rect 961 -841 962 -839
rect 968 -835 969 -833
rect 968 -841 969 -839
rect 975 -835 976 -833
rect 975 -841 976 -839
rect 982 -835 983 -833
rect 982 -841 983 -839
rect 989 -835 990 -833
rect 989 -841 990 -839
rect 996 -835 997 -833
rect 996 -841 997 -839
rect 1003 -835 1004 -833
rect 1003 -841 1004 -839
rect 1010 -835 1011 -833
rect 1010 -841 1011 -839
rect 1017 -835 1018 -833
rect 1017 -841 1018 -839
rect 1024 -835 1025 -833
rect 1024 -841 1025 -839
rect 1031 -835 1032 -833
rect 1031 -841 1032 -839
rect 1038 -835 1039 -833
rect 1038 -841 1039 -839
rect 1045 -835 1046 -833
rect 1045 -841 1046 -839
rect 1052 -835 1053 -833
rect 1052 -841 1053 -839
rect 1059 -835 1060 -833
rect 1059 -841 1060 -839
rect 1066 -835 1067 -833
rect 1066 -841 1067 -839
rect 1073 -835 1074 -833
rect 1073 -841 1074 -839
rect 1080 -835 1081 -833
rect 1080 -841 1081 -839
rect 1087 -835 1088 -833
rect 1087 -841 1088 -839
rect 1094 -835 1095 -833
rect 1094 -841 1095 -839
rect 1101 -835 1102 -833
rect 1101 -841 1102 -839
rect 1108 -835 1109 -833
rect 1108 -841 1109 -839
rect 1115 -835 1116 -833
rect 1115 -841 1116 -839
rect 1122 -835 1123 -833
rect 1122 -841 1123 -839
rect 1129 -835 1130 -833
rect 1129 -841 1130 -839
rect 1136 -835 1137 -833
rect 1136 -841 1137 -839
rect 1143 -835 1144 -833
rect 1143 -841 1144 -839
rect 1150 -835 1151 -833
rect 1150 -841 1151 -839
rect 1157 -835 1158 -833
rect 1157 -841 1158 -839
rect 1164 -835 1165 -833
rect 1164 -841 1165 -839
rect 1171 -835 1172 -833
rect 1171 -841 1172 -839
rect 1178 -835 1179 -833
rect 1178 -841 1179 -839
rect 1185 -835 1186 -833
rect 1185 -841 1186 -839
rect 1192 -835 1193 -833
rect 1192 -841 1193 -839
rect 1199 -835 1200 -833
rect 1199 -841 1200 -839
rect 1206 -835 1207 -833
rect 1206 -841 1207 -839
rect 1213 -835 1214 -833
rect 1213 -841 1214 -839
rect 1220 -835 1221 -833
rect 1220 -841 1221 -839
rect 1227 -835 1228 -833
rect 1227 -841 1228 -839
rect 1234 -835 1235 -833
rect 1234 -841 1235 -839
rect 1241 -835 1242 -833
rect 1241 -841 1242 -839
rect 1248 -835 1249 -833
rect 1248 -841 1249 -839
rect 1255 -835 1256 -833
rect 1255 -841 1256 -839
rect 1262 -835 1263 -833
rect 1262 -841 1263 -839
rect 1416 -835 1417 -833
rect 1416 -841 1417 -839
rect 2 -952 3 -950
rect 2 -958 3 -956
rect 9 -952 10 -950
rect 9 -958 10 -956
rect 16 -952 17 -950
rect 16 -958 17 -956
rect 23 -952 24 -950
rect 23 -958 24 -956
rect 30 -952 31 -950
rect 30 -958 31 -956
rect 37 -952 38 -950
rect 37 -958 38 -956
rect 44 -952 45 -950
rect 44 -958 45 -956
rect 51 -952 52 -950
rect 51 -958 52 -956
rect 58 -952 59 -950
rect 58 -958 59 -956
rect 65 -952 66 -950
rect 68 -952 69 -950
rect 65 -958 66 -956
rect 68 -958 69 -956
rect 72 -952 73 -950
rect 72 -958 73 -956
rect 79 -952 80 -950
rect 79 -958 80 -956
rect 86 -952 87 -950
rect 89 -952 90 -950
rect 86 -958 87 -956
rect 89 -958 90 -956
rect 93 -952 94 -950
rect 93 -958 94 -956
rect 100 -952 101 -950
rect 100 -958 101 -956
rect 107 -952 108 -950
rect 107 -958 108 -956
rect 114 -952 115 -950
rect 114 -958 115 -956
rect 121 -952 122 -950
rect 124 -952 125 -950
rect 121 -958 122 -956
rect 124 -958 125 -956
rect 128 -952 129 -950
rect 131 -952 132 -950
rect 128 -958 129 -956
rect 131 -958 132 -956
rect 135 -952 136 -950
rect 135 -958 136 -956
rect 142 -952 143 -950
rect 142 -958 143 -956
rect 152 -952 153 -950
rect 149 -958 150 -956
rect 152 -958 153 -956
rect 156 -952 157 -950
rect 156 -958 157 -956
rect 163 -952 164 -950
rect 163 -958 164 -956
rect 170 -952 171 -950
rect 170 -958 171 -956
rect 177 -952 178 -950
rect 177 -958 178 -956
rect 184 -952 185 -950
rect 184 -958 185 -956
rect 191 -952 192 -950
rect 191 -958 192 -956
rect 198 -952 199 -950
rect 201 -952 202 -950
rect 198 -958 199 -956
rect 201 -958 202 -956
rect 205 -952 206 -950
rect 205 -958 206 -956
rect 212 -952 213 -950
rect 215 -952 216 -950
rect 212 -958 213 -956
rect 219 -952 220 -950
rect 219 -958 220 -956
rect 226 -952 227 -950
rect 226 -958 227 -956
rect 233 -952 234 -950
rect 233 -958 234 -956
rect 240 -952 241 -950
rect 240 -958 241 -956
rect 247 -952 248 -950
rect 247 -958 248 -956
rect 254 -952 255 -950
rect 254 -958 255 -956
rect 261 -952 262 -950
rect 261 -958 262 -956
rect 268 -952 269 -950
rect 268 -958 269 -956
rect 275 -952 276 -950
rect 275 -958 276 -956
rect 282 -952 283 -950
rect 282 -958 283 -956
rect 289 -952 290 -950
rect 289 -958 290 -956
rect 296 -952 297 -950
rect 296 -958 297 -956
rect 303 -952 304 -950
rect 303 -958 304 -956
rect 310 -952 311 -950
rect 310 -958 311 -956
rect 317 -952 318 -950
rect 320 -952 321 -950
rect 317 -958 318 -956
rect 320 -958 321 -956
rect 324 -952 325 -950
rect 324 -958 325 -956
rect 331 -952 332 -950
rect 331 -958 332 -956
rect 338 -952 339 -950
rect 338 -958 339 -956
rect 345 -952 346 -950
rect 345 -958 346 -956
rect 352 -952 353 -950
rect 352 -958 353 -956
rect 359 -952 360 -950
rect 359 -958 360 -956
rect 366 -952 367 -950
rect 369 -952 370 -950
rect 366 -958 367 -956
rect 369 -958 370 -956
rect 373 -952 374 -950
rect 373 -958 374 -956
rect 380 -952 381 -950
rect 380 -958 381 -956
rect 387 -952 388 -950
rect 387 -958 388 -956
rect 394 -952 395 -950
rect 394 -958 395 -956
rect 401 -952 402 -950
rect 401 -958 402 -956
rect 408 -952 409 -950
rect 408 -958 409 -956
rect 415 -952 416 -950
rect 415 -958 416 -956
rect 422 -952 423 -950
rect 425 -952 426 -950
rect 422 -958 423 -956
rect 425 -958 426 -956
rect 429 -952 430 -950
rect 429 -958 430 -956
rect 436 -952 437 -950
rect 436 -958 437 -956
rect 443 -952 444 -950
rect 443 -958 444 -956
rect 450 -952 451 -950
rect 450 -958 451 -956
rect 453 -958 454 -956
rect 457 -952 458 -950
rect 457 -958 458 -956
rect 464 -952 465 -950
rect 464 -958 465 -956
rect 471 -952 472 -950
rect 471 -958 472 -956
rect 478 -952 479 -950
rect 481 -952 482 -950
rect 478 -958 479 -956
rect 481 -958 482 -956
rect 485 -952 486 -950
rect 485 -958 486 -956
rect 492 -952 493 -950
rect 492 -958 493 -956
rect 499 -952 500 -950
rect 502 -952 503 -950
rect 499 -958 500 -956
rect 502 -958 503 -956
rect 506 -952 507 -950
rect 506 -958 507 -956
rect 513 -952 514 -950
rect 513 -958 514 -956
rect 520 -952 521 -950
rect 520 -958 521 -956
rect 527 -958 528 -956
rect 530 -958 531 -956
rect 534 -952 535 -950
rect 537 -952 538 -950
rect 534 -958 535 -956
rect 537 -958 538 -956
rect 541 -952 542 -950
rect 544 -952 545 -950
rect 541 -958 542 -956
rect 544 -958 545 -956
rect 548 -952 549 -950
rect 548 -958 549 -956
rect 555 -952 556 -950
rect 555 -958 556 -956
rect 562 -952 563 -950
rect 562 -958 563 -956
rect 569 -952 570 -950
rect 569 -958 570 -956
rect 576 -952 577 -950
rect 576 -958 577 -956
rect 583 -952 584 -950
rect 583 -958 584 -956
rect 590 -952 591 -950
rect 590 -958 591 -956
rect 597 -952 598 -950
rect 597 -958 598 -956
rect 604 -952 605 -950
rect 604 -958 605 -956
rect 611 -952 612 -950
rect 614 -952 615 -950
rect 611 -958 612 -956
rect 614 -958 615 -956
rect 618 -952 619 -950
rect 618 -958 619 -956
rect 625 -952 626 -950
rect 628 -952 629 -950
rect 625 -958 626 -956
rect 632 -952 633 -950
rect 635 -952 636 -950
rect 632 -958 633 -956
rect 635 -958 636 -956
rect 639 -952 640 -950
rect 639 -958 640 -956
rect 646 -952 647 -950
rect 646 -958 647 -956
rect 653 -952 654 -950
rect 656 -952 657 -950
rect 653 -958 654 -956
rect 656 -958 657 -956
rect 660 -952 661 -950
rect 660 -958 661 -956
rect 667 -952 668 -950
rect 667 -958 668 -956
rect 674 -952 675 -950
rect 674 -958 675 -956
rect 681 -952 682 -950
rect 681 -958 682 -956
rect 688 -952 689 -950
rect 691 -952 692 -950
rect 688 -958 689 -956
rect 695 -952 696 -950
rect 695 -958 696 -956
rect 702 -952 703 -950
rect 702 -958 703 -956
rect 709 -952 710 -950
rect 712 -952 713 -950
rect 709 -958 710 -956
rect 712 -958 713 -956
rect 716 -952 717 -950
rect 719 -952 720 -950
rect 719 -958 720 -956
rect 723 -952 724 -950
rect 723 -958 724 -956
rect 730 -952 731 -950
rect 730 -958 731 -956
rect 737 -952 738 -950
rect 737 -958 738 -956
rect 747 -952 748 -950
rect 744 -958 745 -956
rect 747 -958 748 -956
rect 751 -952 752 -950
rect 751 -958 752 -956
rect 758 -952 759 -950
rect 758 -958 759 -956
rect 765 -952 766 -950
rect 765 -958 766 -956
rect 772 -952 773 -950
rect 772 -958 773 -956
rect 779 -952 780 -950
rect 779 -958 780 -956
rect 786 -952 787 -950
rect 786 -958 787 -956
rect 793 -952 794 -950
rect 793 -958 794 -956
rect 800 -952 801 -950
rect 800 -958 801 -956
rect 807 -952 808 -950
rect 807 -958 808 -956
rect 814 -952 815 -950
rect 814 -958 815 -956
rect 821 -952 822 -950
rect 824 -952 825 -950
rect 821 -958 822 -956
rect 824 -958 825 -956
rect 828 -952 829 -950
rect 828 -958 829 -956
rect 835 -952 836 -950
rect 835 -958 836 -956
rect 842 -952 843 -950
rect 842 -958 843 -956
rect 849 -952 850 -950
rect 849 -958 850 -956
rect 856 -952 857 -950
rect 856 -958 857 -956
rect 863 -952 864 -950
rect 863 -958 864 -956
rect 870 -952 871 -950
rect 870 -958 871 -956
rect 877 -952 878 -950
rect 877 -958 878 -956
rect 884 -952 885 -950
rect 884 -958 885 -956
rect 891 -952 892 -950
rect 891 -958 892 -956
rect 898 -952 899 -950
rect 898 -958 899 -956
rect 905 -952 906 -950
rect 905 -958 906 -956
rect 912 -952 913 -950
rect 912 -958 913 -956
rect 919 -952 920 -950
rect 919 -958 920 -956
rect 926 -952 927 -950
rect 926 -958 927 -956
rect 933 -952 934 -950
rect 933 -958 934 -956
rect 940 -952 941 -950
rect 940 -958 941 -956
rect 947 -952 948 -950
rect 947 -958 948 -956
rect 954 -952 955 -950
rect 954 -958 955 -956
rect 961 -952 962 -950
rect 961 -958 962 -956
rect 968 -952 969 -950
rect 968 -958 969 -956
rect 975 -952 976 -950
rect 975 -958 976 -956
rect 982 -952 983 -950
rect 982 -958 983 -956
rect 989 -952 990 -950
rect 989 -958 990 -956
rect 996 -952 997 -950
rect 996 -958 997 -956
rect 1003 -952 1004 -950
rect 1003 -958 1004 -956
rect 1010 -952 1011 -950
rect 1010 -958 1011 -956
rect 1017 -952 1018 -950
rect 1017 -958 1018 -956
rect 1024 -952 1025 -950
rect 1024 -958 1025 -956
rect 1031 -952 1032 -950
rect 1031 -958 1032 -956
rect 1038 -952 1039 -950
rect 1038 -958 1039 -956
rect 1045 -952 1046 -950
rect 1045 -958 1046 -956
rect 1052 -952 1053 -950
rect 1052 -958 1053 -956
rect 1059 -952 1060 -950
rect 1059 -958 1060 -956
rect 1066 -952 1067 -950
rect 1066 -958 1067 -956
rect 1073 -952 1074 -950
rect 1073 -958 1074 -956
rect 1080 -952 1081 -950
rect 1080 -958 1081 -956
rect 1087 -952 1088 -950
rect 1087 -958 1088 -956
rect 1094 -952 1095 -950
rect 1094 -958 1095 -956
rect 1101 -952 1102 -950
rect 1101 -958 1102 -956
rect 1108 -952 1109 -950
rect 1108 -958 1109 -956
rect 1115 -952 1116 -950
rect 1115 -958 1116 -956
rect 1122 -952 1123 -950
rect 1122 -958 1123 -956
rect 1129 -952 1130 -950
rect 1129 -958 1130 -956
rect 1136 -952 1137 -950
rect 1136 -958 1137 -956
rect 1143 -952 1144 -950
rect 1143 -958 1144 -956
rect 1150 -952 1151 -950
rect 1150 -958 1151 -956
rect 1157 -952 1158 -950
rect 1157 -958 1158 -956
rect 1164 -952 1165 -950
rect 1164 -958 1165 -956
rect 1171 -952 1172 -950
rect 1171 -958 1172 -956
rect 1178 -952 1179 -950
rect 1178 -958 1179 -956
rect 1185 -952 1186 -950
rect 1185 -958 1186 -956
rect 1192 -952 1193 -950
rect 1192 -958 1193 -956
rect 1195 -958 1196 -956
rect 1199 -952 1200 -950
rect 1202 -952 1203 -950
rect 1199 -958 1200 -956
rect 1206 -952 1207 -950
rect 1206 -958 1207 -956
rect 1437 -952 1438 -950
rect 1437 -958 1438 -956
rect 2 -1081 3 -1079
rect 5 -1081 6 -1079
rect 5 -1087 6 -1085
rect 9 -1081 10 -1079
rect 9 -1087 10 -1085
rect 16 -1081 17 -1079
rect 16 -1087 17 -1085
rect 23 -1081 24 -1079
rect 23 -1087 24 -1085
rect 30 -1081 31 -1079
rect 33 -1081 34 -1079
rect 33 -1087 34 -1085
rect 37 -1081 38 -1079
rect 40 -1081 41 -1079
rect 40 -1087 41 -1085
rect 44 -1081 45 -1079
rect 44 -1087 45 -1085
rect 51 -1081 52 -1079
rect 54 -1081 55 -1079
rect 51 -1087 52 -1085
rect 54 -1087 55 -1085
rect 58 -1081 59 -1079
rect 58 -1087 59 -1085
rect 65 -1081 66 -1079
rect 65 -1087 66 -1085
rect 72 -1081 73 -1079
rect 75 -1081 76 -1079
rect 72 -1087 73 -1085
rect 75 -1087 76 -1085
rect 79 -1081 80 -1079
rect 79 -1087 80 -1085
rect 86 -1081 87 -1079
rect 86 -1087 87 -1085
rect 93 -1081 94 -1079
rect 96 -1081 97 -1079
rect 93 -1087 94 -1085
rect 96 -1087 97 -1085
rect 100 -1081 101 -1079
rect 103 -1081 104 -1079
rect 100 -1087 101 -1085
rect 103 -1087 104 -1085
rect 107 -1081 108 -1079
rect 107 -1087 108 -1085
rect 114 -1081 115 -1079
rect 114 -1087 115 -1085
rect 121 -1081 122 -1079
rect 121 -1087 122 -1085
rect 128 -1081 129 -1079
rect 128 -1087 129 -1085
rect 135 -1081 136 -1079
rect 135 -1087 136 -1085
rect 142 -1081 143 -1079
rect 142 -1087 143 -1085
rect 149 -1081 150 -1079
rect 149 -1087 150 -1085
rect 152 -1087 153 -1085
rect 156 -1081 157 -1079
rect 156 -1087 157 -1085
rect 163 -1081 164 -1079
rect 163 -1087 164 -1085
rect 170 -1081 171 -1079
rect 170 -1087 171 -1085
rect 177 -1081 178 -1079
rect 177 -1087 178 -1085
rect 184 -1081 185 -1079
rect 184 -1087 185 -1085
rect 191 -1081 192 -1079
rect 191 -1087 192 -1085
rect 198 -1081 199 -1079
rect 198 -1087 199 -1085
rect 205 -1081 206 -1079
rect 205 -1087 206 -1085
rect 212 -1081 213 -1079
rect 212 -1087 213 -1085
rect 219 -1081 220 -1079
rect 219 -1087 220 -1085
rect 226 -1081 227 -1079
rect 226 -1087 227 -1085
rect 233 -1081 234 -1079
rect 233 -1087 234 -1085
rect 240 -1081 241 -1079
rect 240 -1087 241 -1085
rect 247 -1081 248 -1079
rect 247 -1087 248 -1085
rect 254 -1081 255 -1079
rect 254 -1087 255 -1085
rect 261 -1081 262 -1079
rect 264 -1081 265 -1079
rect 261 -1087 262 -1085
rect 264 -1087 265 -1085
rect 268 -1081 269 -1079
rect 268 -1087 269 -1085
rect 275 -1081 276 -1079
rect 275 -1087 276 -1085
rect 282 -1081 283 -1079
rect 282 -1087 283 -1085
rect 289 -1081 290 -1079
rect 289 -1087 290 -1085
rect 296 -1081 297 -1079
rect 296 -1087 297 -1085
rect 303 -1081 304 -1079
rect 306 -1081 307 -1079
rect 303 -1087 304 -1085
rect 310 -1081 311 -1079
rect 310 -1087 311 -1085
rect 317 -1081 318 -1079
rect 317 -1087 318 -1085
rect 324 -1081 325 -1079
rect 324 -1087 325 -1085
rect 331 -1081 332 -1079
rect 331 -1087 332 -1085
rect 338 -1081 339 -1079
rect 341 -1081 342 -1079
rect 341 -1087 342 -1085
rect 345 -1081 346 -1079
rect 345 -1087 346 -1085
rect 352 -1081 353 -1079
rect 352 -1087 353 -1085
rect 359 -1081 360 -1079
rect 359 -1087 360 -1085
rect 366 -1081 367 -1079
rect 366 -1087 367 -1085
rect 373 -1081 374 -1079
rect 376 -1081 377 -1079
rect 373 -1087 374 -1085
rect 376 -1087 377 -1085
rect 380 -1081 381 -1079
rect 380 -1087 381 -1085
rect 387 -1081 388 -1079
rect 387 -1087 388 -1085
rect 394 -1081 395 -1079
rect 394 -1087 395 -1085
rect 401 -1081 402 -1079
rect 401 -1087 402 -1085
rect 408 -1081 409 -1079
rect 408 -1087 409 -1085
rect 415 -1081 416 -1079
rect 415 -1087 416 -1085
rect 422 -1081 423 -1079
rect 422 -1087 423 -1085
rect 429 -1081 430 -1079
rect 429 -1087 430 -1085
rect 436 -1081 437 -1079
rect 439 -1081 440 -1079
rect 436 -1087 437 -1085
rect 439 -1087 440 -1085
rect 443 -1081 444 -1079
rect 443 -1087 444 -1085
rect 450 -1081 451 -1079
rect 450 -1087 451 -1085
rect 457 -1081 458 -1079
rect 457 -1087 458 -1085
rect 464 -1081 465 -1079
rect 464 -1087 465 -1085
rect 471 -1081 472 -1079
rect 471 -1087 472 -1085
rect 478 -1081 479 -1079
rect 481 -1081 482 -1079
rect 478 -1087 479 -1085
rect 481 -1087 482 -1085
rect 485 -1081 486 -1079
rect 485 -1087 486 -1085
rect 492 -1081 493 -1079
rect 495 -1081 496 -1079
rect 492 -1087 493 -1085
rect 495 -1087 496 -1085
rect 499 -1081 500 -1079
rect 502 -1081 503 -1079
rect 499 -1087 500 -1085
rect 502 -1087 503 -1085
rect 506 -1081 507 -1079
rect 506 -1087 507 -1085
rect 513 -1081 514 -1079
rect 516 -1081 517 -1079
rect 513 -1087 514 -1085
rect 516 -1087 517 -1085
rect 520 -1081 521 -1079
rect 520 -1087 521 -1085
rect 527 -1081 528 -1079
rect 530 -1081 531 -1079
rect 527 -1087 528 -1085
rect 530 -1087 531 -1085
rect 534 -1081 535 -1079
rect 534 -1087 535 -1085
rect 541 -1081 542 -1079
rect 541 -1087 542 -1085
rect 548 -1081 549 -1079
rect 548 -1087 549 -1085
rect 558 -1081 559 -1079
rect 555 -1087 556 -1085
rect 558 -1087 559 -1085
rect 565 -1081 566 -1079
rect 562 -1087 563 -1085
rect 565 -1087 566 -1085
rect 569 -1081 570 -1079
rect 572 -1081 573 -1079
rect 569 -1087 570 -1085
rect 572 -1087 573 -1085
rect 576 -1081 577 -1079
rect 576 -1087 577 -1085
rect 583 -1081 584 -1079
rect 583 -1087 584 -1085
rect 590 -1081 591 -1079
rect 590 -1087 591 -1085
rect 597 -1081 598 -1079
rect 597 -1087 598 -1085
rect 604 -1081 605 -1079
rect 604 -1087 605 -1085
rect 611 -1081 612 -1079
rect 611 -1087 612 -1085
rect 618 -1081 619 -1079
rect 618 -1087 619 -1085
rect 625 -1081 626 -1079
rect 628 -1081 629 -1079
rect 625 -1087 626 -1085
rect 635 -1081 636 -1079
rect 632 -1087 633 -1085
rect 635 -1087 636 -1085
rect 639 -1081 640 -1079
rect 639 -1087 640 -1085
rect 646 -1081 647 -1079
rect 646 -1087 647 -1085
rect 653 -1081 654 -1079
rect 653 -1087 654 -1085
rect 660 -1081 661 -1079
rect 660 -1087 661 -1085
rect 667 -1081 668 -1079
rect 667 -1087 668 -1085
rect 674 -1081 675 -1079
rect 677 -1081 678 -1079
rect 674 -1087 675 -1085
rect 677 -1087 678 -1085
rect 681 -1081 682 -1079
rect 681 -1087 682 -1085
rect 688 -1081 689 -1079
rect 688 -1087 689 -1085
rect 695 -1081 696 -1079
rect 695 -1087 696 -1085
rect 702 -1081 703 -1079
rect 702 -1087 703 -1085
rect 709 -1081 710 -1079
rect 709 -1087 710 -1085
rect 716 -1081 717 -1079
rect 716 -1087 717 -1085
rect 723 -1081 724 -1079
rect 726 -1081 727 -1079
rect 723 -1087 724 -1085
rect 726 -1087 727 -1085
rect 730 -1081 731 -1079
rect 730 -1087 731 -1085
rect 737 -1081 738 -1079
rect 737 -1087 738 -1085
rect 744 -1081 745 -1079
rect 747 -1081 748 -1079
rect 744 -1087 745 -1085
rect 747 -1087 748 -1085
rect 751 -1081 752 -1079
rect 751 -1087 752 -1085
rect 758 -1081 759 -1079
rect 758 -1087 759 -1085
rect 765 -1081 766 -1079
rect 765 -1087 766 -1085
rect 772 -1081 773 -1079
rect 772 -1087 773 -1085
rect 779 -1081 780 -1079
rect 779 -1087 780 -1085
rect 786 -1081 787 -1079
rect 786 -1087 787 -1085
rect 793 -1081 794 -1079
rect 793 -1087 794 -1085
rect 800 -1081 801 -1079
rect 800 -1087 801 -1085
rect 807 -1081 808 -1079
rect 807 -1087 808 -1085
rect 814 -1081 815 -1079
rect 814 -1087 815 -1085
rect 821 -1081 822 -1079
rect 821 -1087 822 -1085
rect 828 -1081 829 -1079
rect 828 -1087 829 -1085
rect 835 -1081 836 -1079
rect 835 -1087 836 -1085
rect 842 -1081 843 -1079
rect 842 -1087 843 -1085
rect 849 -1081 850 -1079
rect 849 -1087 850 -1085
rect 856 -1081 857 -1079
rect 856 -1087 857 -1085
rect 863 -1081 864 -1079
rect 866 -1081 867 -1079
rect 863 -1087 864 -1085
rect 866 -1087 867 -1085
rect 870 -1081 871 -1079
rect 870 -1087 871 -1085
rect 877 -1081 878 -1079
rect 877 -1087 878 -1085
rect 884 -1081 885 -1079
rect 884 -1087 885 -1085
rect 891 -1081 892 -1079
rect 891 -1087 892 -1085
rect 898 -1081 899 -1079
rect 898 -1087 899 -1085
rect 905 -1081 906 -1079
rect 905 -1087 906 -1085
rect 912 -1081 913 -1079
rect 912 -1087 913 -1085
rect 919 -1081 920 -1079
rect 919 -1087 920 -1085
rect 926 -1081 927 -1079
rect 929 -1081 930 -1079
rect 929 -1087 930 -1085
rect 933 -1081 934 -1079
rect 933 -1087 934 -1085
rect 940 -1081 941 -1079
rect 940 -1087 941 -1085
rect 947 -1081 948 -1079
rect 947 -1087 948 -1085
rect 954 -1081 955 -1079
rect 954 -1087 955 -1085
rect 961 -1081 962 -1079
rect 961 -1087 962 -1085
rect 968 -1081 969 -1079
rect 968 -1087 969 -1085
rect 975 -1081 976 -1079
rect 975 -1087 976 -1085
rect 982 -1081 983 -1079
rect 982 -1087 983 -1085
rect 989 -1081 990 -1079
rect 989 -1087 990 -1085
rect 996 -1081 997 -1079
rect 996 -1087 997 -1085
rect 1003 -1081 1004 -1079
rect 1003 -1087 1004 -1085
rect 1010 -1081 1011 -1079
rect 1010 -1087 1011 -1085
rect 1017 -1081 1018 -1079
rect 1017 -1087 1018 -1085
rect 1024 -1081 1025 -1079
rect 1024 -1087 1025 -1085
rect 1031 -1081 1032 -1079
rect 1031 -1087 1032 -1085
rect 1038 -1081 1039 -1079
rect 1038 -1087 1039 -1085
rect 1045 -1081 1046 -1079
rect 1045 -1087 1046 -1085
rect 1052 -1081 1053 -1079
rect 1052 -1087 1053 -1085
rect 1059 -1081 1060 -1079
rect 1059 -1087 1060 -1085
rect 1066 -1081 1067 -1079
rect 1066 -1087 1067 -1085
rect 1073 -1081 1074 -1079
rect 1073 -1087 1074 -1085
rect 1080 -1081 1081 -1079
rect 1080 -1087 1081 -1085
rect 1087 -1081 1088 -1079
rect 1087 -1087 1088 -1085
rect 1094 -1081 1095 -1079
rect 1094 -1087 1095 -1085
rect 1101 -1081 1102 -1079
rect 1101 -1087 1102 -1085
rect 1108 -1081 1109 -1079
rect 1108 -1087 1109 -1085
rect 1115 -1081 1116 -1079
rect 1115 -1087 1116 -1085
rect 1122 -1081 1123 -1079
rect 1122 -1087 1123 -1085
rect 1129 -1081 1130 -1079
rect 1129 -1087 1130 -1085
rect 1136 -1081 1137 -1079
rect 1136 -1087 1137 -1085
rect 1143 -1081 1144 -1079
rect 1143 -1087 1144 -1085
rect 1150 -1081 1151 -1079
rect 1150 -1087 1151 -1085
rect 1157 -1081 1158 -1079
rect 1157 -1087 1158 -1085
rect 1164 -1081 1165 -1079
rect 1164 -1087 1165 -1085
rect 1171 -1081 1172 -1079
rect 1171 -1087 1172 -1085
rect 1178 -1081 1179 -1079
rect 1178 -1087 1179 -1085
rect 1185 -1081 1186 -1079
rect 1185 -1087 1186 -1085
rect 1192 -1081 1193 -1079
rect 1192 -1087 1193 -1085
rect 1199 -1081 1200 -1079
rect 1199 -1087 1200 -1085
rect 1206 -1081 1207 -1079
rect 1206 -1087 1207 -1085
rect 1213 -1081 1214 -1079
rect 1213 -1087 1214 -1085
rect 1220 -1081 1221 -1079
rect 1220 -1087 1221 -1085
rect 1227 -1081 1228 -1079
rect 1227 -1087 1228 -1085
rect 1234 -1081 1235 -1079
rect 1234 -1087 1235 -1085
rect 1241 -1081 1242 -1079
rect 1241 -1087 1242 -1085
rect 1248 -1081 1249 -1079
rect 1248 -1087 1249 -1085
rect 1255 -1081 1256 -1079
rect 1255 -1087 1256 -1085
rect 1262 -1081 1263 -1079
rect 1262 -1087 1263 -1085
rect 1269 -1081 1270 -1079
rect 1269 -1087 1270 -1085
rect 1276 -1081 1277 -1079
rect 1276 -1087 1277 -1085
rect 1283 -1081 1284 -1079
rect 1283 -1087 1284 -1085
rect 1290 -1081 1291 -1079
rect 1290 -1087 1291 -1085
rect 1297 -1081 1298 -1079
rect 1297 -1087 1298 -1085
rect 1304 -1081 1305 -1079
rect 1304 -1087 1305 -1085
rect 1311 -1081 1312 -1079
rect 1311 -1087 1312 -1085
rect 1318 -1081 1319 -1079
rect 1318 -1087 1319 -1085
rect 1325 -1081 1326 -1079
rect 1325 -1087 1326 -1085
rect 1332 -1081 1333 -1079
rect 1332 -1087 1333 -1085
rect 1339 -1081 1340 -1079
rect 1339 -1087 1340 -1085
rect 1346 -1081 1347 -1079
rect 1346 -1087 1347 -1085
rect 1444 -1081 1445 -1079
rect 1444 -1087 1445 -1085
rect 2 -1206 3 -1204
rect 5 -1206 6 -1204
rect 5 -1212 6 -1210
rect 9 -1206 10 -1204
rect 9 -1212 10 -1210
rect 16 -1206 17 -1204
rect 16 -1212 17 -1210
rect 23 -1206 24 -1204
rect 23 -1212 24 -1210
rect 30 -1206 31 -1204
rect 30 -1212 31 -1210
rect 37 -1206 38 -1204
rect 37 -1212 38 -1210
rect 44 -1206 45 -1204
rect 44 -1212 45 -1210
rect 51 -1206 52 -1204
rect 51 -1212 52 -1210
rect 58 -1206 59 -1204
rect 58 -1212 59 -1210
rect 65 -1206 66 -1204
rect 65 -1212 66 -1210
rect 72 -1206 73 -1204
rect 75 -1206 76 -1204
rect 75 -1212 76 -1210
rect 79 -1206 80 -1204
rect 79 -1212 80 -1210
rect 86 -1206 87 -1204
rect 86 -1212 87 -1210
rect 93 -1206 94 -1204
rect 93 -1212 94 -1210
rect 100 -1206 101 -1204
rect 103 -1206 104 -1204
rect 103 -1212 104 -1210
rect 107 -1206 108 -1204
rect 107 -1212 108 -1210
rect 114 -1206 115 -1204
rect 117 -1206 118 -1204
rect 114 -1212 115 -1210
rect 117 -1212 118 -1210
rect 121 -1206 122 -1204
rect 121 -1212 122 -1210
rect 128 -1206 129 -1204
rect 128 -1212 129 -1210
rect 135 -1206 136 -1204
rect 135 -1212 136 -1210
rect 142 -1206 143 -1204
rect 142 -1212 143 -1210
rect 149 -1206 150 -1204
rect 149 -1212 150 -1210
rect 156 -1206 157 -1204
rect 156 -1212 157 -1210
rect 163 -1206 164 -1204
rect 163 -1212 164 -1210
rect 170 -1206 171 -1204
rect 170 -1212 171 -1210
rect 177 -1206 178 -1204
rect 180 -1206 181 -1204
rect 184 -1206 185 -1204
rect 184 -1212 185 -1210
rect 191 -1206 192 -1204
rect 191 -1212 192 -1210
rect 198 -1206 199 -1204
rect 198 -1212 199 -1210
rect 205 -1206 206 -1204
rect 205 -1212 206 -1210
rect 212 -1206 213 -1204
rect 215 -1206 216 -1204
rect 212 -1212 213 -1210
rect 219 -1206 220 -1204
rect 219 -1212 220 -1210
rect 226 -1206 227 -1204
rect 226 -1212 227 -1210
rect 233 -1206 234 -1204
rect 233 -1212 234 -1210
rect 240 -1206 241 -1204
rect 240 -1212 241 -1210
rect 247 -1206 248 -1204
rect 247 -1212 248 -1210
rect 254 -1206 255 -1204
rect 254 -1212 255 -1210
rect 261 -1206 262 -1204
rect 261 -1212 262 -1210
rect 268 -1206 269 -1204
rect 268 -1212 269 -1210
rect 275 -1206 276 -1204
rect 275 -1212 276 -1210
rect 282 -1206 283 -1204
rect 282 -1212 283 -1210
rect 289 -1206 290 -1204
rect 289 -1212 290 -1210
rect 296 -1206 297 -1204
rect 296 -1212 297 -1210
rect 303 -1206 304 -1204
rect 303 -1212 304 -1210
rect 310 -1206 311 -1204
rect 310 -1212 311 -1210
rect 317 -1206 318 -1204
rect 317 -1212 318 -1210
rect 324 -1206 325 -1204
rect 324 -1212 325 -1210
rect 331 -1206 332 -1204
rect 331 -1212 332 -1210
rect 338 -1206 339 -1204
rect 338 -1212 339 -1210
rect 345 -1206 346 -1204
rect 345 -1212 346 -1210
rect 352 -1206 353 -1204
rect 352 -1212 353 -1210
rect 359 -1206 360 -1204
rect 359 -1212 360 -1210
rect 366 -1206 367 -1204
rect 366 -1212 367 -1210
rect 373 -1206 374 -1204
rect 373 -1212 374 -1210
rect 380 -1206 381 -1204
rect 380 -1212 381 -1210
rect 387 -1206 388 -1204
rect 387 -1212 388 -1210
rect 394 -1206 395 -1204
rect 394 -1212 395 -1210
rect 401 -1206 402 -1204
rect 404 -1206 405 -1204
rect 401 -1212 402 -1210
rect 404 -1212 405 -1210
rect 408 -1206 409 -1204
rect 408 -1212 409 -1210
rect 415 -1206 416 -1204
rect 415 -1212 416 -1210
rect 422 -1206 423 -1204
rect 422 -1212 423 -1210
rect 429 -1206 430 -1204
rect 429 -1212 430 -1210
rect 436 -1206 437 -1204
rect 436 -1212 437 -1210
rect 443 -1206 444 -1204
rect 443 -1212 444 -1210
rect 450 -1206 451 -1204
rect 450 -1212 451 -1210
rect 457 -1206 458 -1204
rect 457 -1212 458 -1210
rect 464 -1206 465 -1204
rect 467 -1206 468 -1204
rect 464 -1212 465 -1210
rect 467 -1212 468 -1210
rect 471 -1206 472 -1204
rect 471 -1212 472 -1210
rect 478 -1206 479 -1204
rect 478 -1212 479 -1210
rect 485 -1206 486 -1204
rect 485 -1212 486 -1210
rect 492 -1206 493 -1204
rect 495 -1206 496 -1204
rect 492 -1212 493 -1210
rect 495 -1212 496 -1210
rect 499 -1206 500 -1204
rect 499 -1212 500 -1210
rect 506 -1206 507 -1204
rect 506 -1212 507 -1210
rect 513 -1206 514 -1204
rect 513 -1212 514 -1210
rect 523 -1206 524 -1204
rect 520 -1212 521 -1210
rect 523 -1212 524 -1210
rect 527 -1206 528 -1204
rect 530 -1206 531 -1204
rect 527 -1212 528 -1210
rect 530 -1212 531 -1210
rect 534 -1206 535 -1204
rect 534 -1212 535 -1210
rect 541 -1206 542 -1204
rect 544 -1206 545 -1204
rect 541 -1212 542 -1210
rect 544 -1212 545 -1210
rect 551 -1206 552 -1204
rect 548 -1212 549 -1210
rect 551 -1212 552 -1210
rect 555 -1206 556 -1204
rect 558 -1206 559 -1204
rect 555 -1212 556 -1210
rect 558 -1212 559 -1210
rect 562 -1206 563 -1204
rect 562 -1212 563 -1210
rect 569 -1206 570 -1204
rect 569 -1212 570 -1210
rect 576 -1206 577 -1204
rect 576 -1212 577 -1210
rect 583 -1206 584 -1204
rect 583 -1212 584 -1210
rect 590 -1206 591 -1204
rect 590 -1212 591 -1210
rect 597 -1206 598 -1204
rect 600 -1206 601 -1204
rect 597 -1212 598 -1210
rect 600 -1212 601 -1210
rect 607 -1206 608 -1204
rect 604 -1212 605 -1210
rect 607 -1212 608 -1210
rect 611 -1206 612 -1204
rect 611 -1212 612 -1210
rect 618 -1206 619 -1204
rect 618 -1212 619 -1210
rect 625 -1206 626 -1204
rect 628 -1206 629 -1204
rect 625 -1212 626 -1210
rect 628 -1212 629 -1210
rect 632 -1206 633 -1204
rect 635 -1206 636 -1204
rect 632 -1212 633 -1210
rect 639 -1206 640 -1204
rect 639 -1212 640 -1210
rect 646 -1206 647 -1204
rect 649 -1206 650 -1204
rect 646 -1212 647 -1210
rect 649 -1212 650 -1210
rect 653 -1206 654 -1204
rect 653 -1212 654 -1210
rect 660 -1206 661 -1204
rect 660 -1212 661 -1210
rect 667 -1206 668 -1204
rect 667 -1212 668 -1210
rect 674 -1206 675 -1204
rect 674 -1212 675 -1210
rect 681 -1206 682 -1204
rect 684 -1206 685 -1204
rect 681 -1212 682 -1210
rect 688 -1206 689 -1204
rect 688 -1212 689 -1210
rect 695 -1206 696 -1204
rect 695 -1212 696 -1210
rect 702 -1206 703 -1204
rect 702 -1212 703 -1210
rect 709 -1206 710 -1204
rect 712 -1206 713 -1204
rect 709 -1212 710 -1210
rect 712 -1212 713 -1210
rect 716 -1206 717 -1204
rect 716 -1212 717 -1210
rect 723 -1206 724 -1204
rect 723 -1212 724 -1210
rect 730 -1206 731 -1204
rect 733 -1206 734 -1204
rect 730 -1212 731 -1210
rect 733 -1212 734 -1210
rect 737 -1206 738 -1204
rect 737 -1212 738 -1210
rect 744 -1206 745 -1204
rect 747 -1206 748 -1204
rect 744 -1212 745 -1210
rect 747 -1212 748 -1210
rect 751 -1206 752 -1204
rect 754 -1206 755 -1204
rect 751 -1212 752 -1210
rect 754 -1212 755 -1210
rect 758 -1206 759 -1204
rect 761 -1206 762 -1204
rect 758 -1212 759 -1210
rect 761 -1212 762 -1210
rect 765 -1206 766 -1204
rect 765 -1212 766 -1210
rect 768 -1212 769 -1210
rect 772 -1206 773 -1204
rect 772 -1212 773 -1210
rect 779 -1206 780 -1204
rect 779 -1212 780 -1210
rect 786 -1206 787 -1204
rect 786 -1212 787 -1210
rect 793 -1206 794 -1204
rect 796 -1206 797 -1204
rect 796 -1212 797 -1210
rect 800 -1206 801 -1204
rect 800 -1212 801 -1210
rect 807 -1206 808 -1204
rect 807 -1212 808 -1210
rect 814 -1206 815 -1204
rect 814 -1212 815 -1210
rect 821 -1206 822 -1204
rect 821 -1212 822 -1210
rect 828 -1206 829 -1204
rect 828 -1212 829 -1210
rect 835 -1206 836 -1204
rect 835 -1212 836 -1210
rect 845 -1206 846 -1204
rect 842 -1212 843 -1210
rect 845 -1212 846 -1210
rect 849 -1206 850 -1204
rect 849 -1212 850 -1210
rect 856 -1206 857 -1204
rect 856 -1212 857 -1210
rect 863 -1206 864 -1204
rect 863 -1212 864 -1210
rect 870 -1206 871 -1204
rect 870 -1212 871 -1210
rect 877 -1206 878 -1204
rect 877 -1212 878 -1210
rect 884 -1206 885 -1204
rect 884 -1212 885 -1210
rect 891 -1206 892 -1204
rect 891 -1212 892 -1210
rect 898 -1206 899 -1204
rect 898 -1212 899 -1210
rect 905 -1206 906 -1204
rect 905 -1212 906 -1210
rect 912 -1206 913 -1204
rect 912 -1212 913 -1210
rect 919 -1206 920 -1204
rect 919 -1212 920 -1210
rect 926 -1206 927 -1204
rect 926 -1212 927 -1210
rect 933 -1206 934 -1204
rect 933 -1212 934 -1210
rect 940 -1206 941 -1204
rect 940 -1212 941 -1210
rect 947 -1206 948 -1204
rect 947 -1212 948 -1210
rect 954 -1206 955 -1204
rect 954 -1212 955 -1210
rect 961 -1206 962 -1204
rect 961 -1212 962 -1210
rect 968 -1206 969 -1204
rect 968 -1212 969 -1210
rect 975 -1206 976 -1204
rect 975 -1212 976 -1210
rect 982 -1206 983 -1204
rect 982 -1212 983 -1210
rect 989 -1206 990 -1204
rect 989 -1212 990 -1210
rect 996 -1206 997 -1204
rect 996 -1212 997 -1210
rect 1003 -1206 1004 -1204
rect 1003 -1212 1004 -1210
rect 1010 -1206 1011 -1204
rect 1010 -1212 1011 -1210
rect 1017 -1206 1018 -1204
rect 1017 -1212 1018 -1210
rect 1024 -1206 1025 -1204
rect 1024 -1212 1025 -1210
rect 1031 -1206 1032 -1204
rect 1031 -1212 1032 -1210
rect 1038 -1206 1039 -1204
rect 1038 -1212 1039 -1210
rect 1045 -1206 1046 -1204
rect 1045 -1212 1046 -1210
rect 1052 -1206 1053 -1204
rect 1052 -1212 1053 -1210
rect 1059 -1206 1060 -1204
rect 1059 -1212 1060 -1210
rect 1066 -1206 1067 -1204
rect 1066 -1212 1067 -1210
rect 1073 -1206 1074 -1204
rect 1073 -1212 1074 -1210
rect 1080 -1206 1081 -1204
rect 1080 -1212 1081 -1210
rect 1087 -1206 1088 -1204
rect 1087 -1212 1088 -1210
rect 1094 -1206 1095 -1204
rect 1094 -1212 1095 -1210
rect 1101 -1206 1102 -1204
rect 1101 -1212 1102 -1210
rect 1108 -1206 1109 -1204
rect 1108 -1212 1109 -1210
rect 1115 -1206 1116 -1204
rect 1122 -1206 1123 -1204
rect 1122 -1212 1123 -1210
rect 1129 -1206 1130 -1204
rect 1129 -1212 1130 -1210
rect 1136 -1206 1137 -1204
rect 1136 -1212 1137 -1210
rect 1143 -1206 1144 -1204
rect 1143 -1212 1144 -1210
rect 1150 -1206 1151 -1204
rect 1150 -1212 1151 -1210
rect 1157 -1206 1158 -1204
rect 1157 -1212 1158 -1210
rect 1164 -1206 1165 -1204
rect 1164 -1212 1165 -1210
rect 1171 -1206 1172 -1204
rect 1171 -1212 1172 -1210
rect 1178 -1206 1179 -1204
rect 1178 -1212 1179 -1210
rect 1185 -1206 1186 -1204
rect 1185 -1212 1186 -1210
rect 1192 -1206 1193 -1204
rect 1192 -1212 1193 -1210
rect 1199 -1206 1200 -1204
rect 1199 -1212 1200 -1210
rect 1206 -1206 1207 -1204
rect 1206 -1212 1207 -1210
rect 1213 -1206 1214 -1204
rect 1213 -1212 1214 -1210
rect 1220 -1206 1221 -1204
rect 1220 -1212 1221 -1210
rect 1227 -1206 1228 -1204
rect 1227 -1212 1228 -1210
rect 1234 -1206 1235 -1204
rect 1234 -1212 1235 -1210
rect 1241 -1206 1242 -1204
rect 1241 -1212 1242 -1210
rect 1248 -1206 1249 -1204
rect 1248 -1212 1249 -1210
rect 1255 -1206 1256 -1204
rect 1255 -1212 1256 -1210
rect 1262 -1206 1263 -1204
rect 1262 -1212 1263 -1210
rect 1269 -1206 1270 -1204
rect 1269 -1212 1270 -1210
rect 1272 -1212 1273 -1210
rect 1276 -1206 1277 -1204
rect 1276 -1212 1277 -1210
rect 1283 -1206 1284 -1204
rect 1283 -1212 1284 -1210
rect 1290 -1206 1291 -1204
rect 1290 -1212 1291 -1210
rect 1297 -1206 1298 -1204
rect 1297 -1212 1298 -1210
rect 1304 -1206 1305 -1204
rect 1304 -1212 1305 -1210
rect 1311 -1206 1312 -1204
rect 1311 -1212 1312 -1210
rect 1318 -1206 1319 -1204
rect 1318 -1212 1319 -1210
rect 1325 -1206 1326 -1204
rect 1325 -1212 1326 -1210
rect 1332 -1206 1333 -1204
rect 1332 -1212 1333 -1210
rect 1339 -1206 1340 -1204
rect 1339 -1212 1340 -1210
rect 1346 -1206 1347 -1204
rect 1346 -1212 1347 -1210
rect 1353 -1206 1354 -1204
rect 1353 -1212 1354 -1210
rect 1360 -1206 1361 -1204
rect 1360 -1212 1361 -1210
rect 1367 -1206 1368 -1204
rect 1367 -1212 1368 -1210
rect 1374 -1206 1375 -1204
rect 1374 -1212 1375 -1210
rect 1451 -1206 1452 -1204
rect 1451 -1212 1452 -1210
rect 2 -1327 3 -1325
rect 2 -1333 3 -1331
rect 9 -1327 10 -1325
rect 9 -1333 10 -1331
rect 16 -1327 17 -1325
rect 16 -1333 17 -1331
rect 23 -1327 24 -1325
rect 23 -1333 24 -1331
rect 30 -1327 31 -1325
rect 30 -1333 31 -1331
rect 37 -1327 38 -1325
rect 37 -1333 38 -1331
rect 44 -1327 45 -1325
rect 44 -1333 45 -1331
rect 51 -1327 52 -1325
rect 51 -1333 52 -1331
rect 58 -1327 59 -1325
rect 61 -1327 62 -1325
rect 58 -1333 59 -1331
rect 61 -1333 62 -1331
rect 68 -1327 69 -1325
rect 65 -1333 66 -1331
rect 68 -1333 69 -1331
rect 72 -1327 73 -1325
rect 72 -1333 73 -1331
rect 79 -1327 80 -1325
rect 79 -1333 80 -1331
rect 82 -1333 83 -1331
rect 86 -1327 87 -1325
rect 89 -1327 90 -1325
rect 86 -1333 87 -1331
rect 89 -1333 90 -1331
rect 93 -1327 94 -1325
rect 93 -1333 94 -1331
rect 100 -1327 101 -1325
rect 100 -1333 101 -1331
rect 107 -1327 108 -1325
rect 107 -1333 108 -1331
rect 114 -1327 115 -1325
rect 114 -1333 115 -1331
rect 121 -1327 122 -1325
rect 124 -1327 125 -1325
rect 121 -1333 122 -1331
rect 124 -1333 125 -1331
rect 128 -1327 129 -1325
rect 128 -1333 129 -1331
rect 135 -1327 136 -1325
rect 138 -1327 139 -1325
rect 135 -1333 136 -1331
rect 138 -1333 139 -1331
rect 142 -1327 143 -1325
rect 142 -1333 143 -1331
rect 149 -1327 150 -1325
rect 149 -1333 150 -1331
rect 156 -1327 157 -1325
rect 156 -1333 157 -1331
rect 163 -1327 164 -1325
rect 163 -1333 164 -1331
rect 166 -1333 167 -1331
rect 170 -1327 171 -1325
rect 173 -1327 174 -1325
rect 170 -1333 171 -1331
rect 173 -1333 174 -1331
rect 177 -1327 178 -1325
rect 177 -1333 178 -1331
rect 184 -1327 185 -1325
rect 184 -1333 185 -1331
rect 191 -1327 192 -1325
rect 191 -1333 192 -1331
rect 198 -1327 199 -1325
rect 198 -1333 199 -1331
rect 205 -1327 206 -1325
rect 205 -1333 206 -1331
rect 212 -1327 213 -1325
rect 212 -1333 213 -1331
rect 219 -1327 220 -1325
rect 219 -1333 220 -1331
rect 226 -1327 227 -1325
rect 226 -1333 227 -1331
rect 233 -1327 234 -1325
rect 233 -1333 234 -1331
rect 240 -1327 241 -1325
rect 240 -1333 241 -1331
rect 247 -1327 248 -1325
rect 247 -1333 248 -1331
rect 254 -1327 255 -1325
rect 254 -1333 255 -1331
rect 261 -1327 262 -1325
rect 261 -1333 262 -1331
rect 268 -1327 269 -1325
rect 268 -1333 269 -1331
rect 275 -1327 276 -1325
rect 275 -1333 276 -1331
rect 282 -1327 283 -1325
rect 282 -1333 283 -1331
rect 289 -1327 290 -1325
rect 289 -1333 290 -1331
rect 296 -1327 297 -1325
rect 296 -1333 297 -1331
rect 303 -1327 304 -1325
rect 303 -1333 304 -1331
rect 310 -1327 311 -1325
rect 310 -1333 311 -1331
rect 317 -1327 318 -1325
rect 317 -1333 318 -1331
rect 324 -1327 325 -1325
rect 324 -1333 325 -1331
rect 331 -1327 332 -1325
rect 331 -1333 332 -1331
rect 338 -1327 339 -1325
rect 338 -1333 339 -1331
rect 345 -1327 346 -1325
rect 345 -1333 346 -1331
rect 352 -1327 353 -1325
rect 352 -1333 353 -1331
rect 359 -1327 360 -1325
rect 359 -1333 360 -1331
rect 366 -1327 367 -1325
rect 369 -1327 370 -1325
rect 366 -1333 367 -1331
rect 369 -1333 370 -1331
rect 376 -1327 377 -1325
rect 373 -1333 374 -1331
rect 376 -1333 377 -1331
rect 380 -1327 381 -1325
rect 380 -1333 381 -1331
rect 387 -1327 388 -1325
rect 390 -1327 391 -1325
rect 387 -1333 388 -1331
rect 390 -1333 391 -1331
rect 394 -1327 395 -1325
rect 394 -1333 395 -1331
rect 401 -1327 402 -1325
rect 401 -1333 402 -1331
rect 408 -1327 409 -1325
rect 408 -1333 409 -1331
rect 415 -1327 416 -1325
rect 418 -1327 419 -1325
rect 415 -1333 416 -1331
rect 418 -1333 419 -1331
rect 422 -1327 423 -1325
rect 422 -1333 423 -1331
rect 432 -1327 433 -1325
rect 429 -1333 430 -1331
rect 436 -1327 437 -1325
rect 436 -1333 437 -1331
rect 443 -1327 444 -1325
rect 446 -1327 447 -1325
rect 443 -1333 444 -1331
rect 446 -1333 447 -1331
rect 450 -1327 451 -1325
rect 450 -1333 451 -1331
rect 457 -1327 458 -1325
rect 457 -1333 458 -1331
rect 464 -1327 465 -1325
rect 464 -1333 465 -1331
rect 471 -1327 472 -1325
rect 471 -1333 472 -1331
rect 478 -1327 479 -1325
rect 478 -1333 479 -1331
rect 485 -1327 486 -1325
rect 485 -1333 486 -1331
rect 492 -1327 493 -1325
rect 492 -1333 493 -1331
rect 499 -1327 500 -1325
rect 499 -1333 500 -1331
rect 506 -1327 507 -1325
rect 506 -1333 507 -1331
rect 513 -1327 514 -1325
rect 513 -1333 514 -1331
rect 520 -1327 521 -1325
rect 520 -1333 521 -1331
rect 527 -1327 528 -1325
rect 527 -1333 528 -1331
rect 534 -1327 535 -1325
rect 534 -1333 535 -1331
rect 541 -1327 542 -1325
rect 544 -1327 545 -1325
rect 541 -1333 542 -1331
rect 544 -1333 545 -1331
rect 548 -1327 549 -1325
rect 548 -1333 549 -1331
rect 555 -1327 556 -1325
rect 555 -1333 556 -1331
rect 562 -1327 563 -1325
rect 562 -1333 563 -1331
rect 569 -1327 570 -1325
rect 572 -1327 573 -1325
rect 569 -1333 570 -1331
rect 572 -1333 573 -1331
rect 576 -1327 577 -1325
rect 576 -1333 577 -1331
rect 583 -1327 584 -1325
rect 583 -1333 584 -1331
rect 590 -1327 591 -1325
rect 590 -1333 591 -1331
rect 597 -1327 598 -1325
rect 597 -1333 598 -1331
rect 604 -1327 605 -1325
rect 604 -1333 605 -1331
rect 611 -1327 612 -1325
rect 614 -1327 615 -1325
rect 611 -1333 612 -1331
rect 614 -1333 615 -1331
rect 618 -1327 619 -1325
rect 621 -1327 622 -1325
rect 625 -1327 626 -1325
rect 625 -1333 626 -1331
rect 632 -1327 633 -1325
rect 635 -1327 636 -1325
rect 632 -1333 633 -1331
rect 635 -1333 636 -1331
rect 639 -1327 640 -1325
rect 639 -1333 640 -1331
rect 646 -1327 647 -1325
rect 646 -1333 647 -1331
rect 653 -1327 654 -1325
rect 653 -1333 654 -1331
rect 660 -1327 661 -1325
rect 660 -1333 661 -1331
rect 667 -1327 668 -1325
rect 667 -1333 668 -1331
rect 674 -1327 675 -1325
rect 674 -1333 675 -1331
rect 681 -1327 682 -1325
rect 684 -1327 685 -1325
rect 681 -1333 682 -1331
rect 684 -1333 685 -1331
rect 688 -1327 689 -1325
rect 688 -1333 689 -1331
rect 695 -1327 696 -1325
rect 698 -1327 699 -1325
rect 695 -1333 696 -1331
rect 698 -1333 699 -1331
rect 702 -1327 703 -1325
rect 705 -1327 706 -1325
rect 702 -1333 703 -1331
rect 705 -1333 706 -1331
rect 709 -1327 710 -1325
rect 709 -1333 710 -1331
rect 719 -1327 720 -1325
rect 716 -1333 717 -1331
rect 719 -1333 720 -1331
rect 723 -1327 724 -1325
rect 723 -1333 724 -1331
rect 730 -1327 731 -1325
rect 733 -1327 734 -1325
rect 730 -1333 731 -1331
rect 737 -1327 738 -1325
rect 737 -1333 738 -1331
rect 744 -1327 745 -1325
rect 744 -1333 745 -1331
rect 751 -1327 752 -1325
rect 751 -1333 752 -1331
rect 758 -1327 759 -1325
rect 758 -1333 759 -1331
rect 765 -1327 766 -1325
rect 765 -1333 766 -1331
rect 772 -1327 773 -1325
rect 772 -1333 773 -1331
rect 779 -1327 780 -1325
rect 779 -1333 780 -1331
rect 786 -1327 787 -1325
rect 786 -1333 787 -1331
rect 793 -1327 794 -1325
rect 793 -1333 794 -1331
rect 800 -1327 801 -1325
rect 800 -1333 801 -1331
rect 807 -1327 808 -1325
rect 807 -1333 808 -1331
rect 814 -1327 815 -1325
rect 817 -1327 818 -1325
rect 814 -1333 815 -1331
rect 821 -1327 822 -1325
rect 821 -1333 822 -1331
rect 828 -1327 829 -1325
rect 828 -1333 829 -1331
rect 835 -1327 836 -1325
rect 835 -1333 836 -1331
rect 842 -1327 843 -1325
rect 842 -1333 843 -1331
rect 849 -1327 850 -1325
rect 849 -1333 850 -1331
rect 856 -1327 857 -1325
rect 856 -1333 857 -1331
rect 863 -1327 864 -1325
rect 866 -1327 867 -1325
rect 866 -1333 867 -1331
rect 870 -1327 871 -1325
rect 870 -1333 871 -1331
rect 877 -1327 878 -1325
rect 877 -1333 878 -1331
rect 884 -1327 885 -1325
rect 884 -1333 885 -1331
rect 891 -1327 892 -1325
rect 891 -1333 892 -1331
rect 898 -1327 899 -1325
rect 898 -1333 899 -1331
rect 905 -1327 906 -1325
rect 905 -1333 906 -1331
rect 912 -1327 913 -1325
rect 915 -1327 916 -1325
rect 912 -1333 913 -1331
rect 915 -1333 916 -1331
rect 919 -1327 920 -1325
rect 919 -1333 920 -1331
rect 926 -1327 927 -1325
rect 926 -1333 927 -1331
rect 933 -1327 934 -1325
rect 933 -1333 934 -1331
rect 940 -1327 941 -1325
rect 940 -1333 941 -1331
rect 947 -1327 948 -1325
rect 947 -1333 948 -1331
rect 954 -1327 955 -1325
rect 954 -1333 955 -1331
rect 961 -1327 962 -1325
rect 961 -1333 962 -1331
rect 968 -1327 969 -1325
rect 968 -1333 969 -1331
rect 975 -1327 976 -1325
rect 975 -1333 976 -1331
rect 982 -1327 983 -1325
rect 982 -1333 983 -1331
rect 989 -1327 990 -1325
rect 989 -1333 990 -1331
rect 996 -1327 997 -1325
rect 996 -1333 997 -1331
rect 1003 -1327 1004 -1325
rect 1003 -1333 1004 -1331
rect 1010 -1327 1011 -1325
rect 1010 -1333 1011 -1331
rect 1017 -1327 1018 -1325
rect 1017 -1333 1018 -1331
rect 1024 -1327 1025 -1325
rect 1024 -1333 1025 -1331
rect 1031 -1327 1032 -1325
rect 1031 -1333 1032 -1331
rect 1038 -1327 1039 -1325
rect 1038 -1333 1039 -1331
rect 1045 -1327 1046 -1325
rect 1045 -1333 1046 -1331
rect 1052 -1327 1053 -1325
rect 1052 -1333 1053 -1331
rect 1059 -1327 1060 -1325
rect 1059 -1333 1060 -1331
rect 1066 -1327 1067 -1325
rect 1066 -1333 1067 -1331
rect 1073 -1327 1074 -1325
rect 1073 -1333 1074 -1331
rect 1080 -1327 1081 -1325
rect 1080 -1333 1081 -1331
rect 1087 -1327 1088 -1325
rect 1087 -1333 1088 -1331
rect 1094 -1327 1095 -1325
rect 1094 -1333 1095 -1331
rect 1101 -1327 1102 -1325
rect 1101 -1333 1102 -1331
rect 1108 -1327 1109 -1325
rect 1108 -1333 1109 -1331
rect 1115 -1333 1116 -1331
rect 1122 -1327 1123 -1325
rect 1122 -1333 1123 -1331
rect 1129 -1327 1130 -1325
rect 1129 -1333 1130 -1331
rect 1136 -1327 1137 -1325
rect 1136 -1333 1137 -1331
rect 1143 -1327 1144 -1325
rect 1143 -1333 1144 -1331
rect 1150 -1327 1151 -1325
rect 1150 -1333 1151 -1331
rect 1157 -1327 1158 -1325
rect 1157 -1333 1158 -1331
rect 1164 -1327 1165 -1325
rect 1164 -1333 1165 -1331
rect 1171 -1327 1172 -1325
rect 1171 -1333 1172 -1331
rect 1178 -1327 1179 -1325
rect 1178 -1333 1179 -1331
rect 1185 -1327 1186 -1325
rect 1185 -1333 1186 -1331
rect 1192 -1327 1193 -1325
rect 1192 -1333 1193 -1331
rect 1199 -1327 1200 -1325
rect 1199 -1333 1200 -1331
rect 1206 -1327 1207 -1325
rect 1206 -1333 1207 -1331
rect 1213 -1327 1214 -1325
rect 1213 -1333 1214 -1331
rect 1220 -1327 1221 -1325
rect 1220 -1333 1221 -1331
rect 1227 -1327 1228 -1325
rect 1227 -1333 1228 -1331
rect 1234 -1327 1235 -1325
rect 1234 -1333 1235 -1331
rect 1241 -1327 1242 -1325
rect 1241 -1333 1242 -1331
rect 1248 -1327 1249 -1325
rect 1248 -1333 1249 -1331
rect 1255 -1327 1256 -1325
rect 1255 -1333 1256 -1331
rect 1262 -1327 1263 -1325
rect 1262 -1333 1263 -1331
rect 1269 -1327 1270 -1325
rect 1272 -1327 1273 -1325
rect 1269 -1333 1270 -1331
rect 1276 -1327 1277 -1325
rect 1276 -1333 1277 -1331
rect 1283 -1327 1284 -1325
rect 1283 -1333 1284 -1331
rect 1290 -1327 1291 -1325
rect 1290 -1333 1291 -1331
rect 1297 -1327 1298 -1325
rect 1297 -1333 1298 -1331
rect 1304 -1327 1305 -1325
rect 1304 -1333 1305 -1331
rect 1311 -1327 1312 -1325
rect 1311 -1333 1312 -1331
rect 1318 -1327 1319 -1325
rect 1318 -1333 1319 -1331
rect 1325 -1327 1326 -1325
rect 1325 -1333 1326 -1331
rect 1332 -1327 1333 -1325
rect 1332 -1333 1333 -1331
rect 1339 -1327 1340 -1325
rect 1339 -1333 1340 -1331
rect 1346 -1327 1347 -1325
rect 1346 -1333 1347 -1331
rect 1353 -1327 1354 -1325
rect 1353 -1333 1354 -1331
rect 1360 -1327 1361 -1325
rect 1360 -1333 1361 -1331
rect 1367 -1327 1368 -1325
rect 1367 -1333 1368 -1331
rect 1374 -1327 1375 -1325
rect 1374 -1333 1375 -1331
rect 1381 -1327 1382 -1325
rect 1381 -1333 1382 -1331
rect 1388 -1327 1389 -1325
rect 1388 -1333 1389 -1331
rect 1458 -1327 1459 -1325
rect 1458 -1333 1459 -1331
rect 2 -1452 3 -1450
rect 2 -1458 3 -1456
rect 9 -1452 10 -1450
rect 9 -1458 10 -1456
rect 16 -1452 17 -1450
rect 16 -1458 17 -1456
rect 23 -1452 24 -1450
rect 23 -1458 24 -1456
rect 33 -1452 34 -1450
rect 30 -1458 31 -1456
rect 33 -1458 34 -1456
rect 37 -1452 38 -1450
rect 37 -1458 38 -1456
rect 44 -1452 45 -1450
rect 44 -1458 45 -1456
rect 51 -1452 52 -1450
rect 51 -1458 52 -1456
rect 58 -1452 59 -1450
rect 58 -1458 59 -1456
rect 65 -1452 66 -1450
rect 65 -1458 66 -1456
rect 72 -1452 73 -1450
rect 72 -1458 73 -1456
rect 79 -1452 80 -1450
rect 82 -1452 83 -1450
rect 79 -1458 80 -1456
rect 82 -1458 83 -1456
rect 86 -1452 87 -1450
rect 86 -1458 87 -1456
rect 93 -1452 94 -1450
rect 93 -1458 94 -1456
rect 100 -1452 101 -1450
rect 100 -1458 101 -1456
rect 107 -1452 108 -1450
rect 107 -1458 108 -1456
rect 114 -1452 115 -1450
rect 114 -1458 115 -1456
rect 121 -1452 122 -1450
rect 121 -1458 122 -1456
rect 128 -1452 129 -1450
rect 131 -1452 132 -1450
rect 128 -1458 129 -1456
rect 131 -1458 132 -1456
rect 135 -1452 136 -1450
rect 135 -1458 136 -1456
rect 142 -1452 143 -1450
rect 142 -1458 143 -1456
rect 149 -1452 150 -1450
rect 152 -1452 153 -1450
rect 149 -1458 150 -1456
rect 152 -1458 153 -1456
rect 156 -1452 157 -1450
rect 156 -1458 157 -1456
rect 163 -1452 164 -1450
rect 163 -1458 164 -1456
rect 170 -1452 171 -1450
rect 170 -1458 171 -1456
rect 177 -1452 178 -1450
rect 177 -1458 178 -1456
rect 184 -1452 185 -1450
rect 184 -1458 185 -1456
rect 191 -1452 192 -1450
rect 191 -1458 192 -1456
rect 198 -1452 199 -1450
rect 198 -1458 199 -1456
rect 205 -1452 206 -1450
rect 205 -1458 206 -1456
rect 212 -1452 213 -1450
rect 212 -1458 213 -1456
rect 219 -1452 220 -1450
rect 219 -1458 220 -1456
rect 226 -1452 227 -1450
rect 226 -1458 227 -1456
rect 233 -1452 234 -1450
rect 233 -1458 234 -1456
rect 240 -1452 241 -1450
rect 240 -1458 241 -1456
rect 247 -1452 248 -1450
rect 247 -1458 248 -1456
rect 254 -1452 255 -1450
rect 254 -1458 255 -1456
rect 261 -1452 262 -1450
rect 261 -1458 262 -1456
rect 268 -1452 269 -1450
rect 268 -1458 269 -1456
rect 275 -1452 276 -1450
rect 275 -1458 276 -1456
rect 282 -1452 283 -1450
rect 282 -1458 283 -1456
rect 289 -1452 290 -1450
rect 289 -1458 290 -1456
rect 296 -1452 297 -1450
rect 296 -1458 297 -1456
rect 303 -1452 304 -1450
rect 303 -1458 304 -1456
rect 310 -1452 311 -1450
rect 310 -1458 311 -1456
rect 317 -1452 318 -1450
rect 320 -1452 321 -1450
rect 317 -1458 318 -1456
rect 324 -1452 325 -1450
rect 324 -1458 325 -1456
rect 331 -1452 332 -1450
rect 331 -1458 332 -1456
rect 338 -1452 339 -1450
rect 338 -1458 339 -1456
rect 345 -1452 346 -1450
rect 345 -1458 346 -1456
rect 352 -1452 353 -1450
rect 352 -1458 353 -1456
rect 359 -1452 360 -1450
rect 359 -1458 360 -1456
rect 366 -1452 367 -1450
rect 366 -1458 367 -1456
rect 373 -1452 374 -1450
rect 373 -1458 374 -1456
rect 380 -1452 381 -1450
rect 380 -1458 381 -1456
rect 387 -1452 388 -1450
rect 387 -1458 388 -1456
rect 394 -1452 395 -1450
rect 397 -1452 398 -1450
rect 394 -1458 395 -1456
rect 397 -1458 398 -1456
rect 401 -1452 402 -1450
rect 401 -1458 402 -1456
rect 408 -1452 409 -1450
rect 411 -1452 412 -1450
rect 408 -1458 409 -1456
rect 415 -1452 416 -1450
rect 415 -1458 416 -1456
rect 422 -1452 423 -1450
rect 422 -1458 423 -1456
rect 429 -1452 430 -1450
rect 429 -1458 430 -1456
rect 436 -1452 437 -1450
rect 436 -1458 437 -1456
rect 446 -1452 447 -1450
rect 443 -1458 444 -1456
rect 446 -1458 447 -1456
rect 450 -1452 451 -1450
rect 450 -1458 451 -1456
rect 457 -1452 458 -1450
rect 460 -1452 461 -1450
rect 457 -1458 458 -1456
rect 464 -1452 465 -1450
rect 464 -1458 465 -1456
rect 471 -1452 472 -1450
rect 471 -1458 472 -1456
rect 478 -1452 479 -1450
rect 478 -1458 479 -1456
rect 485 -1452 486 -1450
rect 485 -1458 486 -1456
rect 492 -1452 493 -1450
rect 492 -1458 493 -1456
rect 499 -1452 500 -1450
rect 499 -1458 500 -1456
rect 506 -1452 507 -1450
rect 509 -1452 510 -1450
rect 506 -1458 507 -1456
rect 509 -1458 510 -1456
rect 513 -1452 514 -1450
rect 513 -1458 514 -1456
rect 520 -1452 521 -1450
rect 520 -1458 521 -1456
rect 527 -1452 528 -1450
rect 527 -1458 528 -1456
rect 534 -1452 535 -1450
rect 534 -1458 535 -1456
rect 537 -1458 538 -1456
rect 541 -1452 542 -1450
rect 541 -1458 542 -1456
rect 548 -1452 549 -1450
rect 551 -1452 552 -1450
rect 548 -1458 549 -1456
rect 551 -1458 552 -1456
rect 555 -1452 556 -1450
rect 555 -1458 556 -1456
rect 562 -1452 563 -1450
rect 565 -1452 566 -1450
rect 562 -1458 563 -1456
rect 565 -1458 566 -1456
rect 569 -1452 570 -1450
rect 569 -1458 570 -1456
rect 576 -1452 577 -1450
rect 576 -1458 577 -1456
rect 583 -1452 584 -1450
rect 583 -1458 584 -1456
rect 590 -1452 591 -1450
rect 590 -1458 591 -1456
rect 597 -1452 598 -1450
rect 597 -1458 598 -1456
rect 604 -1452 605 -1450
rect 604 -1458 605 -1456
rect 611 -1452 612 -1450
rect 611 -1458 612 -1456
rect 618 -1452 619 -1450
rect 618 -1458 619 -1456
rect 625 -1452 626 -1450
rect 625 -1458 626 -1456
rect 632 -1452 633 -1450
rect 632 -1458 633 -1456
rect 639 -1452 640 -1450
rect 642 -1452 643 -1450
rect 639 -1458 640 -1456
rect 642 -1458 643 -1456
rect 646 -1452 647 -1450
rect 649 -1452 650 -1450
rect 646 -1458 647 -1456
rect 649 -1458 650 -1456
rect 653 -1452 654 -1450
rect 653 -1458 654 -1456
rect 660 -1452 661 -1450
rect 660 -1458 661 -1456
rect 667 -1452 668 -1450
rect 667 -1458 668 -1456
rect 674 -1452 675 -1450
rect 674 -1458 675 -1456
rect 681 -1452 682 -1450
rect 681 -1458 682 -1456
rect 688 -1452 689 -1450
rect 688 -1458 689 -1456
rect 695 -1452 696 -1450
rect 695 -1458 696 -1456
rect 702 -1452 703 -1450
rect 702 -1458 703 -1456
rect 709 -1452 710 -1450
rect 709 -1458 710 -1456
rect 716 -1452 717 -1450
rect 716 -1458 717 -1456
rect 723 -1452 724 -1450
rect 726 -1452 727 -1450
rect 723 -1458 724 -1456
rect 730 -1452 731 -1450
rect 730 -1458 731 -1456
rect 737 -1452 738 -1450
rect 737 -1458 738 -1456
rect 744 -1452 745 -1450
rect 747 -1452 748 -1450
rect 744 -1458 745 -1456
rect 747 -1458 748 -1456
rect 751 -1452 752 -1450
rect 751 -1458 752 -1456
rect 758 -1452 759 -1450
rect 758 -1458 759 -1456
rect 765 -1452 766 -1450
rect 765 -1458 766 -1456
rect 772 -1452 773 -1450
rect 772 -1458 773 -1456
rect 779 -1452 780 -1450
rect 782 -1452 783 -1450
rect 779 -1458 780 -1456
rect 782 -1458 783 -1456
rect 786 -1452 787 -1450
rect 786 -1458 787 -1456
rect 793 -1452 794 -1450
rect 796 -1452 797 -1450
rect 793 -1458 794 -1456
rect 796 -1458 797 -1456
rect 800 -1452 801 -1450
rect 800 -1458 801 -1456
rect 807 -1452 808 -1450
rect 807 -1458 808 -1456
rect 814 -1452 815 -1450
rect 817 -1452 818 -1450
rect 814 -1458 815 -1456
rect 817 -1458 818 -1456
rect 821 -1452 822 -1450
rect 824 -1452 825 -1450
rect 824 -1458 825 -1456
rect 828 -1452 829 -1450
rect 831 -1452 832 -1450
rect 831 -1458 832 -1456
rect 835 -1452 836 -1450
rect 835 -1458 836 -1456
rect 842 -1452 843 -1450
rect 842 -1458 843 -1456
rect 849 -1452 850 -1450
rect 852 -1452 853 -1450
rect 849 -1458 850 -1456
rect 852 -1458 853 -1456
rect 856 -1452 857 -1450
rect 859 -1452 860 -1450
rect 856 -1458 857 -1456
rect 859 -1458 860 -1456
rect 866 -1452 867 -1450
rect 863 -1458 864 -1456
rect 866 -1458 867 -1456
rect 870 -1452 871 -1450
rect 870 -1458 871 -1456
rect 877 -1452 878 -1450
rect 877 -1458 878 -1456
rect 887 -1452 888 -1450
rect 887 -1458 888 -1456
rect 891 -1452 892 -1450
rect 891 -1458 892 -1456
rect 898 -1452 899 -1450
rect 898 -1458 899 -1456
rect 905 -1452 906 -1450
rect 905 -1458 906 -1456
rect 912 -1452 913 -1450
rect 912 -1458 913 -1456
rect 919 -1452 920 -1450
rect 919 -1458 920 -1456
rect 926 -1452 927 -1450
rect 926 -1458 927 -1456
rect 933 -1452 934 -1450
rect 933 -1458 934 -1456
rect 940 -1452 941 -1450
rect 940 -1458 941 -1456
rect 947 -1452 948 -1450
rect 947 -1458 948 -1456
rect 954 -1452 955 -1450
rect 954 -1458 955 -1456
rect 961 -1452 962 -1450
rect 961 -1458 962 -1456
rect 968 -1452 969 -1450
rect 968 -1458 969 -1456
rect 975 -1452 976 -1450
rect 975 -1458 976 -1456
rect 982 -1452 983 -1450
rect 982 -1458 983 -1456
rect 989 -1452 990 -1450
rect 989 -1458 990 -1456
rect 996 -1452 997 -1450
rect 996 -1458 997 -1456
rect 1003 -1452 1004 -1450
rect 1003 -1458 1004 -1456
rect 1010 -1452 1011 -1450
rect 1010 -1458 1011 -1456
rect 1017 -1452 1018 -1450
rect 1017 -1458 1018 -1456
rect 1024 -1452 1025 -1450
rect 1024 -1458 1025 -1456
rect 1031 -1452 1032 -1450
rect 1031 -1458 1032 -1456
rect 1038 -1452 1039 -1450
rect 1038 -1458 1039 -1456
rect 1045 -1452 1046 -1450
rect 1045 -1458 1046 -1456
rect 1052 -1452 1053 -1450
rect 1052 -1458 1053 -1456
rect 1059 -1452 1060 -1450
rect 1059 -1458 1060 -1456
rect 1066 -1452 1067 -1450
rect 1066 -1458 1067 -1456
rect 1073 -1452 1074 -1450
rect 1073 -1458 1074 -1456
rect 1080 -1452 1081 -1450
rect 1080 -1458 1081 -1456
rect 1087 -1452 1088 -1450
rect 1087 -1458 1088 -1456
rect 1094 -1452 1095 -1450
rect 1094 -1458 1095 -1456
rect 1101 -1452 1102 -1450
rect 1101 -1458 1102 -1456
rect 1108 -1452 1109 -1450
rect 1108 -1458 1109 -1456
rect 1115 -1452 1116 -1450
rect 1115 -1458 1116 -1456
rect 1122 -1452 1123 -1450
rect 1122 -1458 1123 -1456
rect 1129 -1452 1130 -1450
rect 1129 -1458 1130 -1456
rect 1136 -1452 1137 -1450
rect 1136 -1458 1137 -1456
rect 1143 -1452 1144 -1450
rect 1143 -1458 1144 -1456
rect 1150 -1452 1151 -1450
rect 1150 -1458 1151 -1456
rect 1157 -1452 1158 -1450
rect 1157 -1458 1158 -1456
rect 1164 -1452 1165 -1450
rect 1164 -1458 1165 -1456
rect 1171 -1452 1172 -1450
rect 1171 -1458 1172 -1456
rect 1178 -1452 1179 -1450
rect 1178 -1458 1179 -1456
rect 1185 -1452 1186 -1450
rect 1185 -1458 1186 -1456
rect 1192 -1452 1193 -1450
rect 1192 -1458 1193 -1456
rect 1199 -1452 1200 -1450
rect 1199 -1458 1200 -1456
rect 1206 -1452 1207 -1450
rect 1206 -1458 1207 -1456
rect 1213 -1452 1214 -1450
rect 1213 -1458 1214 -1456
rect 1220 -1452 1221 -1450
rect 1220 -1458 1221 -1456
rect 1227 -1452 1228 -1450
rect 1227 -1458 1228 -1456
rect 1234 -1452 1235 -1450
rect 1234 -1458 1235 -1456
rect 1241 -1452 1242 -1450
rect 1241 -1458 1242 -1456
rect 1248 -1452 1249 -1450
rect 1248 -1458 1249 -1456
rect 1255 -1452 1256 -1450
rect 1255 -1458 1256 -1456
rect 1262 -1452 1263 -1450
rect 1262 -1458 1263 -1456
rect 1269 -1452 1270 -1450
rect 1269 -1458 1270 -1456
rect 1276 -1452 1277 -1450
rect 1276 -1458 1277 -1456
rect 1283 -1452 1284 -1450
rect 1283 -1458 1284 -1456
rect 1290 -1452 1291 -1450
rect 1290 -1458 1291 -1456
rect 1297 -1452 1298 -1450
rect 1297 -1458 1298 -1456
rect 1304 -1452 1305 -1450
rect 1304 -1458 1305 -1456
rect 1311 -1452 1312 -1450
rect 1311 -1458 1312 -1456
rect 1318 -1452 1319 -1450
rect 1318 -1458 1319 -1456
rect 1325 -1452 1326 -1450
rect 1325 -1458 1326 -1456
rect 1332 -1452 1333 -1450
rect 1332 -1458 1333 -1456
rect 1339 -1452 1340 -1450
rect 1339 -1458 1340 -1456
rect 1346 -1452 1347 -1450
rect 1346 -1458 1347 -1456
rect 1353 -1452 1354 -1450
rect 1353 -1458 1354 -1456
rect 1360 -1452 1361 -1450
rect 1360 -1458 1361 -1456
rect 1367 -1452 1368 -1450
rect 1367 -1458 1368 -1456
rect 1374 -1452 1375 -1450
rect 1374 -1458 1375 -1456
rect 1381 -1452 1382 -1450
rect 1381 -1458 1382 -1456
rect 1388 -1452 1389 -1450
rect 1388 -1458 1389 -1456
rect 1395 -1452 1396 -1450
rect 1395 -1458 1396 -1456
rect 1402 -1452 1403 -1450
rect 1402 -1458 1403 -1456
rect 1409 -1452 1410 -1450
rect 1409 -1458 1410 -1456
rect 1416 -1452 1417 -1450
rect 1416 -1458 1417 -1456
rect 1423 -1452 1424 -1450
rect 1423 -1458 1424 -1456
rect 1430 -1452 1431 -1450
rect 1430 -1458 1431 -1456
rect 1437 -1452 1438 -1450
rect 1437 -1458 1438 -1456
rect 1444 -1452 1445 -1450
rect 1444 -1458 1445 -1456
rect 1451 -1452 1452 -1450
rect 1451 -1458 1452 -1456
rect 1454 -1458 1455 -1456
rect 1458 -1452 1459 -1450
rect 1458 -1458 1459 -1456
rect 1465 -1452 1466 -1450
rect 1465 -1458 1466 -1456
rect 2 -1589 3 -1587
rect 2 -1595 3 -1593
rect 9 -1589 10 -1587
rect 12 -1589 13 -1587
rect 12 -1595 13 -1593
rect 16 -1589 17 -1587
rect 19 -1589 20 -1587
rect 16 -1595 17 -1593
rect 23 -1589 24 -1587
rect 23 -1595 24 -1593
rect 30 -1589 31 -1587
rect 30 -1595 31 -1593
rect 37 -1589 38 -1587
rect 40 -1589 41 -1587
rect 37 -1595 38 -1593
rect 40 -1595 41 -1593
rect 44 -1589 45 -1587
rect 44 -1595 45 -1593
rect 51 -1589 52 -1587
rect 54 -1589 55 -1587
rect 51 -1595 52 -1593
rect 54 -1595 55 -1593
rect 58 -1589 59 -1587
rect 58 -1595 59 -1593
rect 65 -1589 66 -1587
rect 65 -1595 66 -1593
rect 72 -1589 73 -1587
rect 72 -1595 73 -1593
rect 79 -1589 80 -1587
rect 79 -1595 80 -1593
rect 86 -1589 87 -1587
rect 89 -1589 90 -1587
rect 86 -1595 87 -1593
rect 89 -1595 90 -1593
rect 93 -1589 94 -1587
rect 93 -1595 94 -1593
rect 100 -1589 101 -1587
rect 103 -1589 104 -1587
rect 100 -1595 101 -1593
rect 103 -1595 104 -1593
rect 107 -1589 108 -1587
rect 107 -1595 108 -1593
rect 114 -1589 115 -1587
rect 117 -1589 118 -1587
rect 114 -1595 115 -1593
rect 117 -1595 118 -1593
rect 121 -1589 122 -1587
rect 121 -1595 122 -1593
rect 128 -1589 129 -1587
rect 128 -1595 129 -1593
rect 135 -1589 136 -1587
rect 138 -1589 139 -1587
rect 135 -1595 136 -1593
rect 138 -1595 139 -1593
rect 142 -1589 143 -1587
rect 145 -1589 146 -1587
rect 142 -1595 143 -1593
rect 145 -1595 146 -1593
rect 149 -1589 150 -1587
rect 149 -1595 150 -1593
rect 156 -1589 157 -1587
rect 156 -1595 157 -1593
rect 163 -1589 164 -1587
rect 163 -1595 164 -1593
rect 170 -1589 171 -1587
rect 170 -1595 171 -1593
rect 180 -1589 181 -1587
rect 177 -1595 178 -1593
rect 180 -1595 181 -1593
rect 184 -1589 185 -1587
rect 184 -1595 185 -1593
rect 191 -1589 192 -1587
rect 191 -1595 192 -1593
rect 198 -1589 199 -1587
rect 198 -1595 199 -1593
rect 205 -1589 206 -1587
rect 205 -1595 206 -1593
rect 212 -1589 213 -1587
rect 212 -1595 213 -1593
rect 219 -1589 220 -1587
rect 219 -1595 220 -1593
rect 226 -1589 227 -1587
rect 226 -1595 227 -1593
rect 233 -1589 234 -1587
rect 233 -1595 234 -1593
rect 240 -1589 241 -1587
rect 240 -1595 241 -1593
rect 247 -1589 248 -1587
rect 247 -1595 248 -1593
rect 254 -1589 255 -1587
rect 254 -1595 255 -1593
rect 261 -1589 262 -1587
rect 261 -1595 262 -1593
rect 268 -1589 269 -1587
rect 268 -1595 269 -1593
rect 275 -1589 276 -1587
rect 275 -1595 276 -1593
rect 282 -1589 283 -1587
rect 282 -1595 283 -1593
rect 289 -1589 290 -1587
rect 289 -1595 290 -1593
rect 296 -1589 297 -1587
rect 296 -1595 297 -1593
rect 303 -1589 304 -1587
rect 303 -1595 304 -1593
rect 310 -1589 311 -1587
rect 310 -1595 311 -1593
rect 317 -1589 318 -1587
rect 317 -1595 318 -1593
rect 324 -1589 325 -1587
rect 324 -1595 325 -1593
rect 331 -1589 332 -1587
rect 331 -1595 332 -1593
rect 338 -1589 339 -1587
rect 338 -1595 339 -1593
rect 345 -1589 346 -1587
rect 345 -1595 346 -1593
rect 352 -1589 353 -1587
rect 352 -1595 353 -1593
rect 359 -1589 360 -1587
rect 359 -1595 360 -1593
rect 366 -1589 367 -1587
rect 366 -1595 367 -1593
rect 373 -1589 374 -1587
rect 373 -1595 374 -1593
rect 380 -1589 381 -1587
rect 380 -1595 381 -1593
rect 387 -1589 388 -1587
rect 387 -1595 388 -1593
rect 394 -1589 395 -1587
rect 394 -1595 395 -1593
rect 401 -1589 402 -1587
rect 404 -1589 405 -1587
rect 404 -1595 405 -1593
rect 408 -1589 409 -1587
rect 408 -1595 409 -1593
rect 415 -1589 416 -1587
rect 415 -1595 416 -1593
rect 422 -1589 423 -1587
rect 422 -1595 423 -1593
rect 429 -1589 430 -1587
rect 432 -1589 433 -1587
rect 429 -1595 430 -1593
rect 432 -1595 433 -1593
rect 436 -1589 437 -1587
rect 436 -1595 437 -1593
rect 443 -1589 444 -1587
rect 443 -1595 444 -1593
rect 450 -1589 451 -1587
rect 450 -1595 451 -1593
rect 457 -1589 458 -1587
rect 460 -1589 461 -1587
rect 457 -1595 458 -1593
rect 460 -1595 461 -1593
rect 464 -1589 465 -1587
rect 464 -1595 465 -1593
rect 471 -1589 472 -1587
rect 471 -1595 472 -1593
rect 478 -1589 479 -1587
rect 478 -1595 479 -1593
rect 485 -1589 486 -1587
rect 488 -1589 489 -1587
rect 485 -1595 486 -1593
rect 492 -1589 493 -1587
rect 492 -1595 493 -1593
rect 495 -1595 496 -1593
rect 499 -1589 500 -1587
rect 499 -1595 500 -1593
rect 506 -1589 507 -1587
rect 506 -1595 507 -1593
rect 513 -1589 514 -1587
rect 513 -1595 514 -1593
rect 520 -1589 521 -1587
rect 523 -1589 524 -1587
rect 520 -1595 521 -1593
rect 523 -1595 524 -1593
rect 527 -1589 528 -1587
rect 527 -1595 528 -1593
rect 534 -1589 535 -1587
rect 537 -1589 538 -1587
rect 534 -1595 535 -1593
rect 537 -1595 538 -1593
rect 541 -1589 542 -1587
rect 541 -1595 542 -1593
rect 548 -1589 549 -1587
rect 548 -1595 549 -1593
rect 555 -1589 556 -1587
rect 558 -1589 559 -1587
rect 555 -1595 556 -1593
rect 558 -1595 559 -1593
rect 562 -1589 563 -1587
rect 562 -1595 563 -1593
rect 569 -1589 570 -1587
rect 572 -1589 573 -1587
rect 569 -1595 570 -1593
rect 572 -1595 573 -1593
rect 576 -1589 577 -1587
rect 576 -1595 577 -1593
rect 583 -1589 584 -1587
rect 583 -1595 584 -1593
rect 590 -1589 591 -1587
rect 590 -1595 591 -1593
rect 597 -1589 598 -1587
rect 597 -1595 598 -1593
rect 604 -1589 605 -1587
rect 604 -1595 605 -1593
rect 611 -1589 612 -1587
rect 611 -1595 612 -1593
rect 618 -1589 619 -1587
rect 621 -1589 622 -1587
rect 618 -1595 619 -1593
rect 621 -1595 622 -1593
rect 625 -1589 626 -1587
rect 625 -1595 626 -1593
rect 632 -1589 633 -1587
rect 632 -1595 633 -1593
rect 639 -1589 640 -1587
rect 639 -1595 640 -1593
rect 646 -1589 647 -1587
rect 646 -1595 647 -1593
rect 653 -1589 654 -1587
rect 653 -1595 654 -1593
rect 663 -1589 664 -1587
rect 660 -1595 661 -1593
rect 663 -1595 664 -1593
rect 667 -1589 668 -1587
rect 667 -1595 668 -1593
rect 674 -1589 675 -1587
rect 674 -1595 675 -1593
rect 681 -1589 682 -1587
rect 681 -1595 682 -1593
rect 688 -1589 689 -1587
rect 688 -1595 689 -1593
rect 695 -1589 696 -1587
rect 695 -1595 696 -1593
rect 702 -1589 703 -1587
rect 705 -1589 706 -1587
rect 702 -1595 703 -1593
rect 705 -1595 706 -1593
rect 709 -1589 710 -1587
rect 709 -1595 710 -1593
rect 716 -1589 717 -1587
rect 716 -1595 717 -1593
rect 723 -1589 724 -1587
rect 723 -1595 724 -1593
rect 730 -1589 731 -1587
rect 730 -1595 731 -1593
rect 737 -1589 738 -1587
rect 737 -1595 738 -1593
rect 744 -1589 745 -1587
rect 744 -1595 745 -1593
rect 751 -1589 752 -1587
rect 751 -1595 752 -1593
rect 758 -1589 759 -1587
rect 758 -1595 759 -1593
rect 765 -1589 766 -1587
rect 765 -1595 766 -1593
rect 772 -1589 773 -1587
rect 772 -1595 773 -1593
rect 779 -1589 780 -1587
rect 779 -1595 780 -1593
rect 786 -1589 787 -1587
rect 786 -1595 787 -1593
rect 793 -1589 794 -1587
rect 793 -1595 794 -1593
rect 800 -1589 801 -1587
rect 803 -1589 804 -1587
rect 800 -1595 801 -1593
rect 803 -1595 804 -1593
rect 807 -1589 808 -1587
rect 807 -1595 808 -1593
rect 814 -1589 815 -1587
rect 814 -1595 815 -1593
rect 821 -1589 822 -1587
rect 821 -1595 822 -1593
rect 828 -1589 829 -1587
rect 831 -1589 832 -1587
rect 828 -1595 829 -1593
rect 831 -1595 832 -1593
rect 835 -1589 836 -1587
rect 835 -1595 836 -1593
rect 842 -1589 843 -1587
rect 842 -1595 843 -1593
rect 849 -1589 850 -1587
rect 849 -1595 850 -1593
rect 856 -1589 857 -1587
rect 859 -1589 860 -1587
rect 856 -1595 857 -1593
rect 859 -1595 860 -1593
rect 863 -1589 864 -1587
rect 863 -1595 864 -1593
rect 870 -1589 871 -1587
rect 870 -1595 871 -1593
rect 877 -1589 878 -1587
rect 877 -1595 878 -1593
rect 884 -1589 885 -1587
rect 884 -1595 885 -1593
rect 891 -1589 892 -1587
rect 894 -1589 895 -1587
rect 898 -1589 899 -1587
rect 898 -1595 899 -1593
rect 905 -1589 906 -1587
rect 905 -1595 906 -1593
rect 912 -1589 913 -1587
rect 912 -1595 913 -1593
rect 919 -1589 920 -1587
rect 919 -1595 920 -1593
rect 926 -1589 927 -1587
rect 926 -1595 927 -1593
rect 933 -1589 934 -1587
rect 933 -1595 934 -1593
rect 940 -1589 941 -1587
rect 940 -1595 941 -1593
rect 947 -1589 948 -1587
rect 947 -1595 948 -1593
rect 954 -1589 955 -1587
rect 954 -1595 955 -1593
rect 961 -1589 962 -1587
rect 961 -1595 962 -1593
rect 968 -1589 969 -1587
rect 968 -1595 969 -1593
rect 975 -1589 976 -1587
rect 975 -1595 976 -1593
rect 982 -1589 983 -1587
rect 982 -1595 983 -1593
rect 989 -1589 990 -1587
rect 989 -1595 990 -1593
rect 996 -1589 997 -1587
rect 996 -1595 997 -1593
rect 1003 -1589 1004 -1587
rect 1003 -1595 1004 -1593
rect 1010 -1589 1011 -1587
rect 1010 -1595 1011 -1593
rect 1017 -1589 1018 -1587
rect 1017 -1595 1018 -1593
rect 1024 -1589 1025 -1587
rect 1024 -1595 1025 -1593
rect 1031 -1589 1032 -1587
rect 1031 -1595 1032 -1593
rect 1038 -1589 1039 -1587
rect 1038 -1595 1039 -1593
rect 1045 -1589 1046 -1587
rect 1048 -1589 1049 -1587
rect 1045 -1595 1046 -1593
rect 1052 -1589 1053 -1587
rect 1052 -1595 1053 -1593
rect 1059 -1589 1060 -1587
rect 1059 -1595 1060 -1593
rect 1066 -1589 1067 -1587
rect 1066 -1595 1067 -1593
rect 1073 -1589 1074 -1587
rect 1073 -1595 1074 -1593
rect 1080 -1589 1081 -1587
rect 1080 -1595 1081 -1593
rect 1087 -1589 1088 -1587
rect 1087 -1595 1088 -1593
rect 1094 -1589 1095 -1587
rect 1094 -1595 1095 -1593
rect 1101 -1589 1102 -1587
rect 1101 -1595 1102 -1593
rect 1108 -1589 1109 -1587
rect 1108 -1595 1109 -1593
rect 1115 -1589 1116 -1587
rect 1115 -1595 1116 -1593
rect 1122 -1589 1123 -1587
rect 1122 -1595 1123 -1593
rect 1129 -1589 1130 -1587
rect 1129 -1595 1130 -1593
rect 1136 -1589 1137 -1587
rect 1136 -1595 1137 -1593
rect 1143 -1589 1144 -1587
rect 1143 -1595 1144 -1593
rect 1150 -1589 1151 -1587
rect 1157 -1589 1158 -1587
rect 1157 -1595 1158 -1593
rect 1164 -1589 1165 -1587
rect 1164 -1595 1165 -1593
rect 1171 -1589 1172 -1587
rect 1171 -1595 1172 -1593
rect 1178 -1589 1179 -1587
rect 1178 -1595 1179 -1593
rect 1185 -1589 1186 -1587
rect 1185 -1595 1186 -1593
rect 1192 -1589 1193 -1587
rect 1192 -1595 1193 -1593
rect 1199 -1589 1200 -1587
rect 1199 -1595 1200 -1593
rect 1206 -1589 1207 -1587
rect 1206 -1595 1207 -1593
rect 1213 -1589 1214 -1587
rect 1213 -1595 1214 -1593
rect 1220 -1589 1221 -1587
rect 1220 -1595 1221 -1593
rect 1227 -1589 1228 -1587
rect 1227 -1595 1228 -1593
rect 1234 -1589 1235 -1587
rect 1234 -1595 1235 -1593
rect 1241 -1589 1242 -1587
rect 1241 -1595 1242 -1593
rect 1248 -1589 1249 -1587
rect 1248 -1595 1249 -1593
rect 1255 -1589 1256 -1587
rect 1255 -1595 1256 -1593
rect 1258 -1595 1259 -1593
rect 1262 -1589 1263 -1587
rect 1262 -1595 1263 -1593
rect 1269 -1589 1270 -1587
rect 1269 -1595 1270 -1593
rect 1276 -1589 1277 -1587
rect 1276 -1595 1277 -1593
rect 1283 -1589 1284 -1587
rect 1283 -1595 1284 -1593
rect 1290 -1589 1291 -1587
rect 1290 -1595 1291 -1593
rect 1297 -1589 1298 -1587
rect 1297 -1595 1298 -1593
rect 1304 -1589 1305 -1587
rect 1304 -1595 1305 -1593
rect 1311 -1589 1312 -1587
rect 1311 -1595 1312 -1593
rect 1318 -1589 1319 -1587
rect 1318 -1595 1319 -1593
rect 1325 -1589 1326 -1587
rect 1325 -1595 1326 -1593
rect 1332 -1589 1333 -1587
rect 1332 -1595 1333 -1593
rect 1339 -1589 1340 -1587
rect 1339 -1595 1340 -1593
rect 1346 -1589 1347 -1587
rect 1346 -1595 1347 -1593
rect 1353 -1589 1354 -1587
rect 1353 -1595 1354 -1593
rect 2 -1720 3 -1718
rect 2 -1726 3 -1724
rect 9 -1720 10 -1718
rect 9 -1726 10 -1724
rect 16 -1726 17 -1724
rect 19 -1726 20 -1724
rect 23 -1726 24 -1724
rect 26 -1726 27 -1724
rect 30 -1720 31 -1718
rect 30 -1726 31 -1724
rect 33 -1726 34 -1724
rect 37 -1720 38 -1718
rect 37 -1726 38 -1724
rect 44 -1720 45 -1718
rect 47 -1720 48 -1718
rect 44 -1726 45 -1724
rect 51 -1720 52 -1718
rect 54 -1720 55 -1718
rect 51 -1726 52 -1724
rect 54 -1726 55 -1724
rect 58 -1720 59 -1718
rect 58 -1726 59 -1724
rect 65 -1720 66 -1718
rect 65 -1726 66 -1724
rect 72 -1720 73 -1718
rect 72 -1726 73 -1724
rect 79 -1720 80 -1718
rect 79 -1726 80 -1724
rect 86 -1720 87 -1718
rect 86 -1726 87 -1724
rect 93 -1720 94 -1718
rect 96 -1720 97 -1718
rect 93 -1726 94 -1724
rect 96 -1726 97 -1724
rect 100 -1720 101 -1718
rect 100 -1726 101 -1724
rect 107 -1720 108 -1718
rect 110 -1720 111 -1718
rect 107 -1726 108 -1724
rect 110 -1726 111 -1724
rect 114 -1720 115 -1718
rect 114 -1726 115 -1724
rect 121 -1720 122 -1718
rect 121 -1726 122 -1724
rect 128 -1720 129 -1718
rect 128 -1726 129 -1724
rect 135 -1720 136 -1718
rect 135 -1726 136 -1724
rect 142 -1720 143 -1718
rect 142 -1726 143 -1724
rect 149 -1720 150 -1718
rect 152 -1720 153 -1718
rect 149 -1726 150 -1724
rect 152 -1726 153 -1724
rect 159 -1720 160 -1718
rect 156 -1726 157 -1724
rect 159 -1726 160 -1724
rect 163 -1720 164 -1718
rect 163 -1726 164 -1724
rect 170 -1720 171 -1718
rect 170 -1726 171 -1724
rect 177 -1720 178 -1718
rect 177 -1726 178 -1724
rect 184 -1720 185 -1718
rect 184 -1726 185 -1724
rect 191 -1720 192 -1718
rect 194 -1720 195 -1718
rect 191 -1726 192 -1724
rect 194 -1726 195 -1724
rect 198 -1720 199 -1718
rect 198 -1726 199 -1724
rect 205 -1720 206 -1718
rect 205 -1726 206 -1724
rect 212 -1720 213 -1718
rect 212 -1726 213 -1724
rect 219 -1720 220 -1718
rect 219 -1726 220 -1724
rect 226 -1720 227 -1718
rect 226 -1726 227 -1724
rect 233 -1720 234 -1718
rect 233 -1726 234 -1724
rect 240 -1720 241 -1718
rect 240 -1726 241 -1724
rect 247 -1720 248 -1718
rect 247 -1726 248 -1724
rect 254 -1720 255 -1718
rect 254 -1726 255 -1724
rect 261 -1720 262 -1718
rect 261 -1726 262 -1724
rect 268 -1720 269 -1718
rect 268 -1726 269 -1724
rect 275 -1720 276 -1718
rect 275 -1726 276 -1724
rect 282 -1720 283 -1718
rect 282 -1726 283 -1724
rect 289 -1720 290 -1718
rect 289 -1726 290 -1724
rect 296 -1720 297 -1718
rect 296 -1726 297 -1724
rect 303 -1720 304 -1718
rect 303 -1726 304 -1724
rect 310 -1720 311 -1718
rect 310 -1726 311 -1724
rect 317 -1720 318 -1718
rect 320 -1720 321 -1718
rect 317 -1726 318 -1724
rect 320 -1726 321 -1724
rect 324 -1720 325 -1718
rect 324 -1726 325 -1724
rect 331 -1720 332 -1718
rect 331 -1726 332 -1724
rect 338 -1720 339 -1718
rect 338 -1726 339 -1724
rect 345 -1720 346 -1718
rect 345 -1726 346 -1724
rect 352 -1720 353 -1718
rect 352 -1726 353 -1724
rect 359 -1720 360 -1718
rect 359 -1726 360 -1724
rect 366 -1720 367 -1718
rect 366 -1726 367 -1724
rect 373 -1720 374 -1718
rect 376 -1720 377 -1718
rect 373 -1726 374 -1724
rect 376 -1726 377 -1724
rect 380 -1720 381 -1718
rect 380 -1726 381 -1724
rect 387 -1720 388 -1718
rect 387 -1726 388 -1724
rect 394 -1720 395 -1718
rect 394 -1726 395 -1724
rect 401 -1720 402 -1718
rect 404 -1720 405 -1718
rect 401 -1726 402 -1724
rect 404 -1726 405 -1724
rect 408 -1720 409 -1718
rect 408 -1726 409 -1724
rect 415 -1720 416 -1718
rect 415 -1726 416 -1724
rect 422 -1720 423 -1718
rect 422 -1726 423 -1724
rect 429 -1720 430 -1718
rect 429 -1726 430 -1724
rect 436 -1720 437 -1718
rect 436 -1726 437 -1724
rect 443 -1720 444 -1718
rect 443 -1726 444 -1724
rect 450 -1720 451 -1718
rect 450 -1726 451 -1724
rect 457 -1720 458 -1718
rect 460 -1720 461 -1718
rect 457 -1726 458 -1724
rect 460 -1726 461 -1724
rect 464 -1720 465 -1718
rect 464 -1726 465 -1724
rect 471 -1720 472 -1718
rect 471 -1726 472 -1724
rect 478 -1720 479 -1718
rect 478 -1726 479 -1724
rect 485 -1720 486 -1718
rect 488 -1720 489 -1718
rect 485 -1726 486 -1724
rect 488 -1726 489 -1724
rect 492 -1720 493 -1718
rect 492 -1726 493 -1724
rect 499 -1720 500 -1718
rect 499 -1726 500 -1724
rect 506 -1720 507 -1718
rect 506 -1726 507 -1724
rect 513 -1720 514 -1718
rect 513 -1726 514 -1724
rect 520 -1720 521 -1718
rect 523 -1720 524 -1718
rect 520 -1726 521 -1724
rect 523 -1726 524 -1724
rect 527 -1720 528 -1718
rect 527 -1726 528 -1724
rect 534 -1720 535 -1718
rect 534 -1726 535 -1724
rect 541 -1720 542 -1718
rect 541 -1726 542 -1724
rect 551 -1720 552 -1718
rect 548 -1726 549 -1724
rect 551 -1726 552 -1724
rect 555 -1720 556 -1718
rect 555 -1726 556 -1724
rect 558 -1726 559 -1724
rect 562 -1720 563 -1718
rect 562 -1726 563 -1724
rect 569 -1720 570 -1718
rect 569 -1726 570 -1724
rect 576 -1720 577 -1718
rect 576 -1726 577 -1724
rect 583 -1720 584 -1718
rect 583 -1726 584 -1724
rect 590 -1720 591 -1718
rect 590 -1726 591 -1724
rect 597 -1720 598 -1718
rect 597 -1726 598 -1724
rect 604 -1720 605 -1718
rect 604 -1726 605 -1724
rect 611 -1720 612 -1718
rect 611 -1726 612 -1724
rect 618 -1720 619 -1718
rect 618 -1726 619 -1724
rect 625 -1720 626 -1718
rect 625 -1726 626 -1724
rect 632 -1720 633 -1718
rect 632 -1726 633 -1724
rect 639 -1720 640 -1718
rect 639 -1726 640 -1724
rect 646 -1720 647 -1718
rect 646 -1726 647 -1724
rect 653 -1720 654 -1718
rect 653 -1726 654 -1724
rect 660 -1720 661 -1718
rect 660 -1726 661 -1724
rect 667 -1720 668 -1718
rect 670 -1720 671 -1718
rect 667 -1726 668 -1724
rect 674 -1720 675 -1718
rect 674 -1726 675 -1724
rect 681 -1720 682 -1718
rect 681 -1726 682 -1724
rect 688 -1720 689 -1718
rect 688 -1726 689 -1724
rect 695 -1720 696 -1718
rect 695 -1726 696 -1724
rect 702 -1720 703 -1718
rect 702 -1726 703 -1724
rect 709 -1720 710 -1718
rect 709 -1726 710 -1724
rect 716 -1720 717 -1718
rect 716 -1726 717 -1724
rect 723 -1720 724 -1718
rect 723 -1726 724 -1724
rect 730 -1720 731 -1718
rect 730 -1726 731 -1724
rect 737 -1720 738 -1718
rect 737 -1726 738 -1724
rect 744 -1720 745 -1718
rect 747 -1720 748 -1718
rect 744 -1726 745 -1724
rect 747 -1726 748 -1724
rect 751 -1720 752 -1718
rect 754 -1720 755 -1718
rect 751 -1726 752 -1724
rect 754 -1726 755 -1724
rect 758 -1720 759 -1718
rect 758 -1726 759 -1724
rect 765 -1720 766 -1718
rect 765 -1726 766 -1724
rect 772 -1720 773 -1718
rect 775 -1720 776 -1718
rect 772 -1726 773 -1724
rect 775 -1726 776 -1724
rect 779 -1720 780 -1718
rect 779 -1726 780 -1724
rect 786 -1720 787 -1718
rect 786 -1726 787 -1724
rect 793 -1720 794 -1718
rect 793 -1726 794 -1724
rect 800 -1720 801 -1718
rect 800 -1726 801 -1724
rect 807 -1720 808 -1718
rect 807 -1726 808 -1724
rect 814 -1720 815 -1718
rect 814 -1726 815 -1724
rect 821 -1720 822 -1718
rect 821 -1726 822 -1724
rect 828 -1720 829 -1718
rect 828 -1726 829 -1724
rect 835 -1720 836 -1718
rect 835 -1726 836 -1724
rect 842 -1720 843 -1718
rect 842 -1726 843 -1724
rect 849 -1720 850 -1718
rect 849 -1726 850 -1724
rect 856 -1720 857 -1718
rect 856 -1726 857 -1724
rect 863 -1720 864 -1718
rect 863 -1726 864 -1724
rect 870 -1720 871 -1718
rect 870 -1726 871 -1724
rect 877 -1720 878 -1718
rect 877 -1726 878 -1724
rect 884 -1720 885 -1718
rect 884 -1726 885 -1724
rect 891 -1720 892 -1718
rect 894 -1720 895 -1718
rect 894 -1726 895 -1724
rect 898 -1720 899 -1718
rect 901 -1720 902 -1718
rect 898 -1726 899 -1724
rect 901 -1726 902 -1724
rect 905 -1720 906 -1718
rect 905 -1726 906 -1724
rect 912 -1720 913 -1718
rect 912 -1726 913 -1724
rect 919 -1720 920 -1718
rect 919 -1726 920 -1724
rect 926 -1720 927 -1718
rect 926 -1726 927 -1724
rect 933 -1720 934 -1718
rect 933 -1726 934 -1724
rect 940 -1720 941 -1718
rect 940 -1726 941 -1724
rect 943 -1726 944 -1724
rect 947 -1720 948 -1718
rect 947 -1726 948 -1724
rect 954 -1720 955 -1718
rect 954 -1726 955 -1724
rect 961 -1720 962 -1718
rect 961 -1726 962 -1724
rect 968 -1720 969 -1718
rect 968 -1726 969 -1724
rect 975 -1720 976 -1718
rect 975 -1726 976 -1724
rect 982 -1720 983 -1718
rect 982 -1726 983 -1724
rect 989 -1720 990 -1718
rect 989 -1726 990 -1724
rect 996 -1720 997 -1718
rect 996 -1726 997 -1724
rect 1003 -1720 1004 -1718
rect 1003 -1726 1004 -1724
rect 1010 -1720 1011 -1718
rect 1010 -1726 1011 -1724
rect 1017 -1720 1018 -1718
rect 1017 -1726 1018 -1724
rect 1024 -1720 1025 -1718
rect 1024 -1726 1025 -1724
rect 1031 -1720 1032 -1718
rect 1031 -1726 1032 -1724
rect 1038 -1720 1039 -1718
rect 1038 -1726 1039 -1724
rect 1045 -1720 1046 -1718
rect 1045 -1726 1046 -1724
rect 1052 -1720 1053 -1718
rect 1052 -1726 1053 -1724
rect 1059 -1720 1060 -1718
rect 1059 -1726 1060 -1724
rect 1066 -1720 1067 -1718
rect 1066 -1726 1067 -1724
rect 1069 -1726 1070 -1724
rect 1073 -1720 1074 -1718
rect 1073 -1726 1074 -1724
rect 1080 -1720 1081 -1718
rect 1080 -1726 1081 -1724
rect 1087 -1720 1088 -1718
rect 1087 -1726 1088 -1724
rect 1094 -1720 1095 -1718
rect 1094 -1726 1095 -1724
rect 1101 -1720 1102 -1718
rect 1101 -1726 1102 -1724
rect 1108 -1720 1109 -1718
rect 1108 -1726 1109 -1724
rect 1115 -1720 1116 -1718
rect 1115 -1726 1116 -1724
rect 1122 -1726 1123 -1724
rect 1125 -1726 1126 -1724
rect 1129 -1720 1130 -1718
rect 1129 -1726 1130 -1724
rect 1136 -1720 1137 -1718
rect 1136 -1726 1137 -1724
rect 1143 -1720 1144 -1718
rect 1143 -1726 1144 -1724
rect 1150 -1726 1151 -1724
rect 1157 -1720 1158 -1718
rect 1157 -1726 1158 -1724
rect 1164 -1720 1165 -1718
rect 1164 -1726 1165 -1724
rect 1171 -1720 1172 -1718
rect 1171 -1726 1172 -1724
rect 1178 -1720 1179 -1718
rect 1178 -1726 1179 -1724
rect 1185 -1720 1186 -1718
rect 1185 -1726 1186 -1724
rect 1192 -1720 1193 -1718
rect 1192 -1726 1193 -1724
rect 1199 -1720 1200 -1718
rect 1199 -1726 1200 -1724
rect 1206 -1720 1207 -1718
rect 1206 -1726 1207 -1724
rect 1213 -1720 1214 -1718
rect 1213 -1726 1214 -1724
rect 1220 -1720 1221 -1718
rect 1220 -1726 1221 -1724
rect 1227 -1720 1228 -1718
rect 1227 -1726 1228 -1724
rect 1234 -1720 1235 -1718
rect 1234 -1726 1235 -1724
rect 1241 -1720 1242 -1718
rect 1241 -1726 1242 -1724
rect 1248 -1720 1249 -1718
rect 1248 -1726 1249 -1724
rect 1255 -1720 1256 -1718
rect 1258 -1720 1259 -1718
rect 1255 -1726 1256 -1724
rect 1262 -1720 1263 -1718
rect 1262 -1726 1263 -1724
rect 1269 -1720 1270 -1718
rect 1269 -1726 1270 -1724
rect 1276 -1720 1277 -1718
rect 1276 -1726 1277 -1724
rect 1283 -1720 1284 -1718
rect 1283 -1726 1284 -1724
rect 1290 -1720 1291 -1718
rect 1290 -1726 1291 -1724
rect 1297 -1720 1298 -1718
rect 1297 -1726 1298 -1724
rect 1304 -1720 1305 -1718
rect 1304 -1726 1305 -1724
rect 1311 -1720 1312 -1718
rect 1311 -1726 1312 -1724
rect 1318 -1720 1319 -1718
rect 1318 -1726 1319 -1724
rect 1325 -1720 1326 -1718
rect 1328 -1720 1329 -1718
rect 1328 -1726 1329 -1724
rect 2 -1839 3 -1837
rect 2 -1845 3 -1843
rect 9 -1839 10 -1837
rect 9 -1845 10 -1843
rect 16 -1839 17 -1837
rect 16 -1845 17 -1843
rect 23 -1839 24 -1837
rect 26 -1839 27 -1837
rect 23 -1845 24 -1843
rect 30 -1839 31 -1837
rect 30 -1845 31 -1843
rect 40 -1839 41 -1837
rect 37 -1845 38 -1843
rect 40 -1845 41 -1843
rect 44 -1839 45 -1837
rect 47 -1839 48 -1837
rect 44 -1845 45 -1843
rect 47 -1845 48 -1843
rect 51 -1839 52 -1837
rect 54 -1839 55 -1837
rect 51 -1845 52 -1843
rect 54 -1845 55 -1843
rect 58 -1839 59 -1837
rect 58 -1845 59 -1843
rect 65 -1839 66 -1837
rect 68 -1839 69 -1837
rect 68 -1845 69 -1843
rect 72 -1839 73 -1837
rect 72 -1845 73 -1843
rect 79 -1839 80 -1837
rect 79 -1845 80 -1843
rect 86 -1839 87 -1837
rect 86 -1845 87 -1843
rect 93 -1839 94 -1837
rect 93 -1845 94 -1843
rect 100 -1839 101 -1837
rect 100 -1845 101 -1843
rect 107 -1839 108 -1837
rect 107 -1845 108 -1843
rect 114 -1839 115 -1837
rect 117 -1839 118 -1837
rect 114 -1845 115 -1843
rect 121 -1839 122 -1837
rect 121 -1845 122 -1843
rect 128 -1839 129 -1837
rect 128 -1845 129 -1843
rect 135 -1839 136 -1837
rect 138 -1839 139 -1837
rect 135 -1845 136 -1843
rect 138 -1845 139 -1843
rect 142 -1839 143 -1837
rect 142 -1845 143 -1843
rect 149 -1839 150 -1837
rect 152 -1839 153 -1837
rect 149 -1845 150 -1843
rect 152 -1845 153 -1843
rect 156 -1839 157 -1837
rect 156 -1845 157 -1843
rect 163 -1839 164 -1837
rect 163 -1845 164 -1843
rect 170 -1839 171 -1837
rect 170 -1845 171 -1843
rect 177 -1839 178 -1837
rect 177 -1845 178 -1843
rect 184 -1839 185 -1837
rect 184 -1845 185 -1843
rect 191 -1839 192 -1837
rect 191 -1845 192 -1843
rect 198 -1839 199 -1837
rect 198 -1845 199 -1843
rect 205 -1839 206 -1837
rect 205 -1845 206 -1843
rect 212 -1839 213 -1837
rect 212 -1845 213 -1843
rect 219 -1839 220 -1837
rect 219 -1845 220 -1843
rect 226 -1839 227 -1837
rect 226 -1845 227 -1843
rect 233 -1839 234 -1837
rect 233 -1845 234 -1843
rect 240 -1839 241 -1837
rect 240 -1845 241 -1843
rect 247 -1839 248 -1837
rect 247 -1845 248 -1843
rect 254 -1839 255 -1837
rect 254 -1845 255 -1843
rect 261 -1839 262 -1837
rect 261 -1845 262 -1843
rect 268 -1839 269 -1837
rect 268 -1845 269 -1843
rect 275 -1839 276 -1837
rect 275 -1845 276 -1843
rect 282 -1839 283 -1837
rect 282 -1845 283 -1843
rect 289 -1839 290 -1837
rect 289 -1845 290 -1843
rect 296 -1839 297 -1837
rect 299 -1839 300 -1837
rect 296 -1845 297 -1843
rect 299 -1845 300 -1843
rect 303 -1839 304 -1837
rect 303 -1845 304 -1843
rect 310 -1839 311 -1837
rect 310 -1845 311 -1843
rect 317 -1839 318 -1837
rect 317 -1845 318 -1843
rect 324 -1839 325 -1837
rect 324 -1845 325 -1843
rect 331 -1839 332 -1837
rect 331 -1845 332 -1843
rect 338 -1839 339 -1837
rect 338 -1845 339 -1843
rect 345 -1839 346 -1837
rect 345 -1845 346 -1843
rect 352 -1839 353 -1837
rect 355 -1839 356 -1837
rect 352 -1845 353 -1843
rect 355 -1845 356 -1843
rect 359 -1839 360 -1837
rect 359 -1845 360 -1843
rect 366 -1839 367 -1837
rect 369 -1839 370 -1837
rect 366 -1845 367 -1843
rect 369 -1845 370 -1843
rect 373 -1839 374 -1837
rect 373 -1845 374 -1843
rect 380 -1839 381 -1837
rect 380 -1845 381 -1843
rect 387 -1839 388 -1837
rect 390 -1839 391 -1837
rect 387 -1845 388 -1843
rect 394 -1839 395 -1837
rect 394 -1845 395 -1843
rect 401 -1839 402 -1837
rect 401 -1845 402 -1843
rect 408 -1839 409 -1837
rect 408 -1845 409 -1843
rect 415 -1839 416 -1837
rect 415 -1845 416 -1843
rect 422 -1839 423 -1837
rect 422 -1845 423 -1843
rect 429 -1839 430 -1837
rect 429 -1845 430 -1843
rect 436 -1839 437 -1837
rect 436 -1845 437 -1843
rect 443 -1839 444 -1837
rect 443 -1845 444 -1843
rect 450 -1839 451 -1837
rect 450 -1845 451 -1843
rect 457 -1839 458 -1837
rect 457 -1845 458 -1843
rect 464 -1839 465 -1837
rect 467 -1839 468 -1837
rect 464 -1845 465 -1843
rect 467 -1845 468 -1843
rect 471 -1839 472 -1837
rect 471 -1845 472 -1843
rect 478 -1839 479 -1837
rect 481 -1839 482 -1837
rect 478 -1845 479 -1843
rect 481 -1845 482 -1843
rect 485 -1839 486 -1837
rect 485 -1845 486 -1843
rect 492 -1839 493 -1837
rect 492 -1845 493 -1843
rect 499 -1839 500 -1837
rect 499 -1845 500 -1843
rect 506 -1839 507 -1837
rect 506 -1845 507 -1843
rect 513 -1839 514 -1837
rect 516 -1845 517 -1843
rect 520 -1839 521 -1837
rect 520 -1845 521 -1843
rect 527 -1839 528 -1837
rect 527 -1845 528 -1843
rect 534 -1839 535 -1837
rect 534 -1845 535 -1843
rect 541 -1839 542 -1837
rect 541 -1845 542 -1843
rect 548 -1839 549 -1837
rect 548 -1845 549 -1843
rect 555 -1839 556 -1837
rect 555 -1845 556 -1843
rect 562 -1839 563 -1837
rect 562 -1845 563 -1843
rect 569 -1839 570 -1837
rect 569 -1845 570 -1843
rect 576 -1839 577 -1837
rect 576 -1845 577 -1843
rect 583 -1839 584 -1837
rect 586 -1839 587 -1837
rect 583 -1845 584 -1843
rect 586 -1845 587 -1843
rect 590 -1839 591 -1837
rect 590 -1845 591 -1843
rect 597 -1839 598 -1837
rect 597 -1845 598 -1843
rect 604 -1839 605 -1837
rect 607 -1839 608 -1837
rect 604 -1845 605 -1843
rect 607 -1845 608 -1843
rect 611 -1839 612 -1837
rect 614 -1839 615 -1837
rect 611 -1845 612 -1843
rect 614 -1845 615 -1843
rect 618 -1839 619 -1837
rect 618 -1845 619 -1843
rect 625 -1839 626 -1837
rect 628 -1839 629 -1837
rect 625 -1845 626 -1843
rect 628 -1845 629 -1843
rect 632 -1839 633 -1837
rect 632 -1845 633 -1843
rect 639 -1839 640 -1837
rect 642 -1839 643 -1837
rect 639 -1845 640 -1843
rect 642 -1845 643 -1843
rect 646 -1839 647 -1837
rect 646 -1845 647 -1843
rect 653 -1839 654 -1837
rect 653 -1845 654 -1843
rect 656 -1845 657 -1843
rect 660 -1839 661 -1837
rect 660 -1845 661 -1843
rect 667 -1839 668 -1837
rect 667 -1845 668 -1843
rect 674 -1839 675 -1837
rect 674 -1845 675 -1843
rect 681 -1839 682 -1837
rect 681 -1845 682 -1843
rect 688 -1839 689 -1837
rect 688 -1845 689 -1843
rect 695 -1839 696 -1837
rect 695 -1845 696 -1843
rect 702 -1839 703 -1837
rect 702 -1845 703 -1843
rect 709 -1839 710 -1837
rect 712 -1839 713 -1837
rect 709 -1845 710 -1843
rect 712 -1845 713 -1843
rect 716 -1839 717 -1837
rect 719 -1839 720 -1837
rect 716 -1845 717 -1843
rect 719 -1845 720 -1843
rect 723 -1839 724 -1837
rect 723 -1845 724 -1843
rect 730 -1839 731 -1837
rect 733 -1839 734 -1837
rect 737 -1839 738 -1837
rect 737 -1845 738 -1843
rect 744 -1839 745 -1837
rect 744 -1845 745 -1843
rect 751 -1839 752 -1837
rect 754 -1839 755 -1837
rect 751 -1845 752 -1843
rect 754 -1845 755 -1843
rect 758 -1839 759 -1837
rect 761 -1839 762 -1837
rect 758 -1845 759 -1843
rect 761 -1845 762 -1843
rect 765 -1839 766 -1837
rect 765 -1845 766 -1843
rect 772 -1839 773 -1837
rect 772 -1845 773 -1843
rect 779 -1839 780 -1837
rect 779 -1845 780 -1843
rect 786 -1839 787 -1837
rect 786 -1845 787 -1843
rect 793 -1839 794 -1837
rect 793 -1845 794 -1843
rect 800 -1839 801 -1837
rect 800 -1845 801 -1843
rect 807 -1839 808 -1837
rect 807 -1845 808 -1843
rect 814 -1839 815 -1837
rect 814 -1845 815 -1843
rect 821 -1839 822 -1837
rect 821 -1845 822 -1843
rect 828 -1839 829 -1837
rect 828 -1845 829 -1843
rect 835 -1839 836 -1837
rect 835 -1845 836 -1843
rect 842 -1839 843 -1837
rect 842 -1845 843 -1843
rect 849 -1839 850 -1837
rect 849 -1845 850 -1843
rect 856 -1839 857 -1837
rect 856 -1845 857 -1843
rect 863 -1839 864 -1837
rect 863 -1845 864 -1843
rect 870 -1839 871 -1837
rect 870 -1845 871 -1843
rect 877 -1839 878 -1837
rect 877 -1845 878 -1843
rect 884 -1839 885 -1837
rect 884 -1845 885 -1843
rect 891 -1839 892 -1837
rect 891 -1845 892 -1843
rect 898 -1839 899 -1837
rect 898 -1845 899 -1843
rect 905 -1839 906 -1837
rect 905 -1845 906 -1843
rect 912 -1839 913 -1837
rect 912 -1845 913 -1843
rect 919 -1839 920 -1837
rect 919 -1845 920 -1843
rect 926 -1839 927 -1837
rect 926 -1845 927 -1843
rect 933 -1839 934 -1837
rect 933 -1845 934 -1843
rect 940 -1839 941 -1837
rect 940 -1845 941 -1843
rect 947 -1839 948 -1837
rect 947 -1845 948 -1843
rect 954 -1839 955 -1837
rect 954 -1845 955 -1843
rect 961 -1839 962 -1837
rect 961 -1845 962 -1843
rect 968 -1839 969 -1837
rect 968 -1845 969 -1843
rect 975 -1839 976 -1837
rect 975 -1845 976 -1843
rect 982 -1839 983 -1837
rect 982 -1845 983 -1843
rect 989 -1839 990 -1837
rect 989 -1845 990 -1843
rect 996 -1839 997 -1837
rect 996 -1845 997 -1843
rect 1003 -1839 1004 -1837
rect 1003 -1845 1004 -1843
rect 1010 -1839 1011 -1837
rect 1010 -1845 1011 -1843
rect 1017 -1839 1018 -1837
rect 1017 -1845 1018 -1843
rect 1024 -1839 1025 -1837
rect 1024 -1845 1025 -1843
rect 1031 -1839 1032 -1837
rect 1031 -1845 1032 -1843
rect 1038 -1839 1039 -1837
rect 1038 -1845 1039 -1843
rect 1045 -1839 1046 -1837
rect 1045 -1845 1046 -1843
rect 1052 -1839 1053 -1837
rect 1052 -1845 1053 -1843
rect 1059 -1839 1060 -1837
rect 1059 -1845 1060 -1843
rect 1066 -1839 1067 -1837
rect 1066 -1845 1067 -1843
rect 1073 -1839 1074 -1837
rect 1073 -1845 1074 -1843
rect 1080 -1839 1081 -1837
rect 1080 -1845 1081 -1843
rect 1087 -1839 1088 -1837
rect 1087 -1845 1088 -1843
rect 1094 -1839 1095 -1837
rect 1094 -1845 1095 -1843
rect 1101 -1839 1102 -1837
rect 1101 -1845 1102 -1843
rect 1108 -1839 1109 -1837
rect 1108 -1845 1109 -1843
rect 1115 -1839 1116 -1837
rect 1115 -1845 1116 -1843
rect 1122 -1839 1123 -1837
rect 1122 -1845 1123 -1843
rect 1129 -1839 1130 -1837
rect 1129 -1845 1130 -1843
rect 1136 -1839 1137 -1837
rect 1136 -1845 1137 -1843
rect 1143 -1839 1144 -1837
rect 1143 -1845 1144 -1843
rect 1150 -1839 1151 -1837
rect 1150 -1845 1151 -1843
rect 1157 -1839 1158 -1837
rect 1157 -1845 1158 -1843
rect 1164 -1839 1165 -1837
rect 1164 -1845 1165 -1843
rect 1171 -1839 1172 -1837
rect 1171 -1845 1172 -1843
rect 1178 -1839 1179 -1837
rect 1178 -1845 1179 -1843
rect 1185 -1839 1186 -1837
rect 1185 -1845 1186 -1843
rect 1192 -1839 1193 -1837
rect 1192 -1845 1193 -1843
rect 1199 -1839 1200 -1837
rect 1199 -1845 1200 -1843
rect 1206 -1839 1207 -1837
rect 1206 -1845 1207 -1843
rect 1213 -1839 1214 -1837
rect 1213 -1845 1214 -1843
rect 1220 -1839 1221 -1837
rect 1220 -1845 1221 -1843
rect 1227 -1839 1228 -1837
rect 1227 -1845 1228 -1843
rect 1234 -1839 1235 -1837
rect 1234 -1845 1235 -1843
rect 1241 -1839 1242 -1837
rect 1241 -1845 1242 -1843
rect 1248 -1839 1249 -1837
rect 1248 -1845 1249 -1843
rect 1255 -1839 1256 -1837
rect 1255 -1845 1256 -1843
rect 1262 -1839 1263 -1837
rect 1262 -1845 1263 -1843
rect 1269 -1839 1270 -1837
rect 1269 -1845 1270 -1843
rect 1276 -1839 1277 -1837
rect 1276 -1845 1277 -1843
rect 1283 -1839 1284 -1837
rect 1286 -1839 1287 -1837
rect 9 -1962 10 -1960
rect 9 -1968 10 -1966
rect 16 -1962 17 -1960
rect 16 -1968 17 -1966
rect 23 -1962 24 -1960
rect 23 -1968 24 -1966
rect 30 -1962 31 -1960
rect 30 -1968 31 -1966
rect 37 -1962 38 -1960
rect 37 -1968 38 -1966
rect 44 -1962 45 -1960
rect 44 -1968 45 -1966
rect 51 -1962 52 -1960
rect 51 -1968 52 -1966
rect 54 -1968 55 -1966
rect 58 -1962 59 -1960
rect 58 -1968 59 -1966
rect 65 -1962 66 -1960
rect 68 -1962 69 -1960
rect 65 -1968 66 -1966
rect 68 -1968 69 -1966
rect 72 -1962 73 -1960
rect 72 -1968 73 -1966
rect 79 -1962 80 -1960
rect 79 -1968 80 -1966
rect 86 -1962 87 -1960
rect 89 -1962 90 -1960
rect 86 -1968 87 -1966
rect 89 -1968 90 -1966
rect 93 -1962 94 -1960
rect 96 -1962 97 -1960
rect 93 -1968 94 -1966
rect 96 -1968 97 -1966
rect 100 -1962 101 -1960
rect 103 -1962 104 -1960
rect 103 -1968 104 -1966
rect 107 -1962 108 -1960
rect 107 -1968 108 -1966
rect 114 -1962 115 -1960
rect 114 -1968 115 -1966
rect 121 -1962 122 -1960
rect 121 -1968 122 -1966
rect 128 -1962 129 -1960
rect 128 -1968 129 -1966
rect 135 -1962 136 -1960
rect 138 -1962 139 -1960
rect 135 -1968 136 -1966
rect 138 -1968 139 -1966
rect 142 -1962 143 -1960
rect 142 -1968 143 -1966
rect 149 -1962 150 -1960
rect 149 -1968 150 -1966
rect 156 -1962 157 -1960
rect 156 -1968 157 -1966
rect 163 -1962 164 -1960
rect 163 -1968 164 -1966
rect 170 -1962 171 -1960
rect 170 -1968 171 -1966
rect 173 -1968 174 -1966
rect 177 -1962 178 -1960
rect 177 -1968 178 -1966
rect 184 -1962 185 -1960
rect 184 -1968 185 -1966
rect 191 -1962 192 -1960
rect 191 -1968 192 -1966
rect 198 -1962 199 -1960
rect 198 -1968 199 -1966
rect 205 -1962 206 -1960
rect 205 -1968 206 -1966
rect 212 -1962 213 -1960
rect 212 -1968 213 -1966
rect 219 -1962 220 -1960
rect 219 -1968 220 -1966
rect 226 -1962 227 -1960
rect 226 -1968 227 -1966
rect 233 -1962 234 -1960
rect 233 -1968 234 -1966
rect 240 -1962 241 -1960
rect 240 -1968 241 -1966
rect 247 -1962 248 -1960
rect 247 -1968 248 -1966
rect 254 -1962 255 -1960
rect 254 -1968 255 -1966
rect 261 -1962 262 -1960
rect 264 -1962 265 -1960
rect 261 -1968 262 -1966
rect 268 -1962 269 -1960
rect 268 -1968 269 -1966
rect 275 -1962 276 -1960
rect 275 -1968 276 -1966
rect 282 -1962 283 -1960
rect 285 -1962 286 -1960
rect 282 -1968 283 -1966
rect 285 -1968 286 -1966
rect 289 -1962 290 -1960
rect 289 -1968 290 -1966
rect 296 -1962 297 -1960
rect 296 -1968 297 -1966
rect 303 -1962 304 -1960
rect 303 -1968 304 -1966
rect 310 -1962 311 -1960
rect 310 -1968 311 -1966
rect 317 -1962 318 -1960
rect 320 -1962 321 -1960
rect 317 -1968 318 -1966
rect 320 -1968 321 -1966
rect 324 -1962 325 -1960
rect 324 -1968 325 -1966
rect 331 -1962 332 -1960
rect 331 -1968 332 -1966
rect 338 -1962 339 -1960
rect 338 -1968 339 -1966
rect 345 -1962 346 -1960
rect 345 -1968 346 -1966
rect 352 -1962 353 -1960
rect 352 -1968 353 -1966
rect 359 -1962 360 -1960
rect 359 -1968 360 -1966
rect 366 -1962 367 -1960
rect 369 -1962 370 -1960
rect 366 -1968 367 -1966
rect 369 -1968 370 -1966
rect 373 -1962 374 -1960
rect 373 -1968 374 -1966
rect 380 -1962 381 -1960
rect 387 -1962 388 -1960
rect 387 -1968 388 -1966
rect 394 -1962 395 -1960
rect 394 -1968 395 -1966
rect 401 -1962 402 -1960
rect 401 -1968 402 -1966
rect 408 -1962 409 -1960
rect 408 -1968 409 -1966
rect 415 -1962 416 -1960
rect 415 -1968 416 -1966
rect 422 -1962 423 -1960
rect 422 -1968 423 -1966
rect 429 -1962 430 -1960
rect 432 -1962 433 -1960
rect 429 -1968 430 -1966
rect 432 -1968 433 -1966
rect 436 -1962 437 -1960
rect 436 -1968 437 -1966
rect 443 -1962 444 -1960
rect 443 -1968 444 -1966
rect 450 -1962 451 -1960
rect 450 -1968 451 -1966
rect 457 -1962 458 -1960
rect 460 -1962 461 -1960
rect 457 -1968 458 -1966
rect 460 -1968 461 -1966
rect 464 -1962 465 -1960
rect 464 -1968 465 -1966
rect 471 -1962 472 -1960
rect 471 -1968 472 -1966
rect 478 -1962 479 -1960
rect 478 -1968 479 -1966
rect 485 -1962 486 -1960
rect 485 -1968 486 -1966
rect 492 -1962 493 -1960
rect 495 -1962 496 -1960
rect 492 -1968 493 -1966
rect 499 -1962 500 -1960
rect 499 -1968 500 -1966
rect 506 -1962 507 -1960
rect 506 -1968 507 -1966
rect 513 -1962 514 -1960
rect 513 -1968 514 -1966
rect 520 -1962 521 -1960
rect 523 -1962 524 -1960
rect 520 -1968 521 -1966
rect 523 -1968 524 -1966
rect 527 -1962 528 -1960
rect 527 -1968 528 -1966
rect 534 -1962 535 -1960
rect 534 -1968 535 -1966
rect 541 -1962 542 -1960
rect 541 -1968 542 -1966
rect 548 -1962 549 -1960
rect 548 -1968 549 -1966
rect 555 -1962 556 -1960
rect 558 -1962 559 -1960
rect 555 -1968 556 -1966
rect 558 -1968 559 -1966
rect 562 -1962 563 -1960
rect 562 -1968 563 -1966
rect 569 -1962 570 -1960
rect 572 -1962 573 -1960
rect 569 -1968 570 -1966
rect 572 -1968 573 -1966
rect 576 -1962 577 -1960
rect 576 -1968 577 -1966
rect 583 -1962 584 -1960
rect 583 -1968 584 -1966
rect 590 -1962 591 -1960
rect 590 -1968 591 -1966
rect 597 -1962 598 -1960
rect 597 -1968 598 -1966
rect 604 -1962 605 -1960
rect 607 -1962 608 -1960
rect 604 -1968 605 -1966
rect 607 -1968 608 -1966
rect 611 -1962 612 -1960
rect 611 -1968 612 -1966
rect 618 -1962 619 -1960
rect 618 -1968 619 -1966
rect 625 -1962 626 -1960
rect 625 -1968 626 -1966
rect 632 -1962 633 -1960
rect 632 -1968 633 -1966
rect 639 -1962 640 -1960
rect 639 -1968 640 -1966
rect 646 -1962 647 -1960
rect 646 -1968 647 -1966
rect 653 -1962 654 -1960
rect 653 -1968 654 -1966
rect 660 -1962 661 -1960
rect 660 -1968 661 -1966
rect 667 -1962 668 -1960
rect 667 -1968 668 -1966
rect 677 -1962 678 -1960
rect 674 -1968 675 -1966
rect 677 -1968 678 -1966
rect 681 -1962 682 -1960
rect 681 -1968 682 -1966
rect 688 -1962 689 -1960
rect 688 -1968 689 -1966
rect 695 -1962 696 -1960
rect 695 -1968 696 -1966
rect 702 -1962 703 -1960
rect 705 -1962 706 -1960
rect 702 -1968 703 -1966
rect 709 -1962 710 -1960
rect 709 -1968 710 -1966
rect 716 -1962 717 -1960
rect 716 -1968 717 -1966
rect 723 -1962 724 -1960
rect 723 -1968 724 -1966
rect 730 -1962 731 -1960
rect 730 -1968 731 -1966
rect 737 -1962 738 -1960
rect 737 -1968 738 -1966
rect 744 -1962 745 -1960
rect 744 -1968 745 -1966
rect 751 -1962 752 -1960
rect 751 -1968 752 -1966
rect 758 -1962 759 -1960
rect 761 -1962 762 -1960
rect 758 -1968 759 -1966
rect 761 -1968 762 -1966
rect 765 -1962 766 -1960
rect 765 -1968 766 -1966
rect 772 -1962 773 -1960
rect 772 -1968 773 -1966
rect 779 -1962 780 -1960
rect 779 -1968 780 -1966
rect 786 -1962 787 -1960
rect 786 -1968 787 -1966
rect 793 -1962 794 -1960
rect 793 -1968 794 -1966
rect 800 -1962 801 -1960
rect 800 -1968 801 -1966
rect 807 -1962 808 -1960
rect 807 -1968 808 -1966
rect 814 -1962 815 -1960
rect 814 -1968 815 -1966
rect 821 -1962 822 -1960
rect 821 -1968 822 -1966
rect 828 -1962 829 -1960
rect 828 -1968 829 -1966
rect 835 -1962 836 -1960
rect 838 -1962 839 -1960
rect 835 -1968 836 -1966
rect 838 -1968 839 -1966
rect 842 -1962 843 -1960
rect 842 -1968 843 -1966
rect 849 -1962 850 -1960
rect 849 -1968 850 -1966
rect 856 -1962 857 -1960
rect 856 -1968 857 -1966
rect 863 -1962 864 -1960
rect 863 -1968 864 -1966
rect 870 -1962 871 -1960
rect 870 -1968 871 -1966
rect 877 -1962 878 -1960
rect 877 -1968 878 -1966
rect 884 -1962 885 -1960
rect 884 -1968 885 -1966
rect 891 -1962 892 -1960
rect 891 -1968 892 -1966
rect 898 -1962 899 -1960
rect 898 -1968 899 -1966
rect 905 -1962 906 -1960
rect 905 -1968 906 -1966
rect 912 -1962 913 -1960
rect 912 -1968 913 -1966
rect 919 -1962 920 -1960
rect 922 -1962 923 -1960
rect 919 -1968 920 -1966
rect 926 -1962 927 -1960
rect 926 -1968 927 -1966
rect 933 -1962 934 -1960
rect 933 -1968 934 -1966
rect 940 -1962 941 -1960
rect 940 -1968 941 -1966
rect 947 -1962 948 -1960
rect 947 -1968 948 -1966
rect 954 -1962 955 -1960
rect 954 -1968 955 -1966
rect 961 -1962 962 -1960
rect 961 -1968 962 -1966
rect 964 -1968 965 -1966
rect 968 -1962 969 -1960
rect 968 -1968 969 -1966
rect 971 -1968 972 -1966
rect 975 -1962 976 -1960
rect 975 -1968 976 -1966
rect 982 -1962 983 -1960
rect 982 -1968 983 -1966
rect 989 -1962 990 -1960
rect 989 -1968 990 -1966
rect 996 -1962 997 -1960
rect 996 -1968 997 -1966
rect 1003 -1962 1004 -1960
rect 1003 -1968 1004 -1966
rect 1010 -1962 1011 -1960
rect 1010 -1968 1011 -1966
rect 1017 -1962 1018 -1960
rect 1017 -1968 1018 -1966
rect 1024 -1962 1025 -1960
rect 1024 -1968 1025 -1966
rect 1031 -1962 1032 -1960
rect 1031 -1968 1032 -1966
rect 1038 -1962 1039 -1960
rect 1038 -1968 1039 -1966
rect 1045 -1962 1046 -1960
rect 1045 -1968 1046 -1966
rect 1052 -1962 1053 -1960
rect 1052 -1968 1053 -1966
rect 1059 -1962 1060 -1960
rect 1059 -1968 1060 -1966
rect 1066 -1962 1067 -1960
rect 1066 -1968 1067 -1966
rect 1073 -1962 1074 -1960
rect 1073 -1968 1074 -1966
rect 1080 -1962 1081 -1960
rect 1080 -1968 1081 -1966
rect 1087 -1962 1088 -1960
rect 1087 -1968 1088 -1966
rect 1094 -1962 1095 -1960
rect 1094 -1968 1095 -1966
rect 1101 -1962 1102 -1960
rect 1101 -1968 1102 -1966
rect 1108 -1962 1109 -1960
rect 1108 -1968 1109 -1966
rect 1115 -1962 1116 -1960
rect 1115 -1968 1116 -1966
rect 1122 -1962 1123 -1960
rect 1122 -1968 1123 -1966
rect 1129 -1962 1130 -1960
rect 1129 -1968 1130 -1966
rect 1136 -1962 1137 -1960
rect 1136 -1968 1137 -1966
rect 1143 -1962 1144 -1960
rect 1143 -1968 1144 -1966
rect 1150 -1962 1151 -1960
rect 1150 -1968 1151 -1966
rect 1157 -1962 1158 -1960
rect 1157 -1968 1158 -1966
rect 1164 -1962 1165 -1960
rect 1164 -1968 1165 -1966
rect 1171 -1962 1172 -1960
rect 1171 -1968 1172 -1966
rect 1178 -1962 1179 -1960
rect 1178 -1968 1179 -1966
rect 1185 -1962 1186 -1960
rect 1185 -1968 1186 -1966
rect 1192 -1962 1193 -1960
rect 1192 -1968 1193 -1966
rect 1199 -1962 1200 -1960
rect 1199 -1968 1200 -1966
rect 1206 -1962 1207 -1960
rect 1206 -1968 1207 -1966
rect 1213 -1962 1214 -1960
rect 1213 -1968 1214 -1966
rect 1223 -1962 1224 -1960
rect 1220 -1968 1221 -1966
rect 1223 -1968 1224 -1966
rect 1227 -1962 1228 -1960
rect 1227 -1968 1228 -1966
rect 1234 -1962 1235 -1960
rect 1234 -1968 1235 -1966
rect 2 -2065 3 -2063
rect 2 -2071 3 -2069
rect 9 -2065 10 -2063
rect 9 -2071 10 -2069
rect 16 -2065 17 -2063
rect 16 -2071 17 -2069
rect 23 -2065 24 -2063
rect 23 -2071 24 -2069
rect 30 -2065 31 -2063
rect 30 -2071 31 -2069
rect 37 -2065 38 -2063
rect 37 -2071 38 -2069
rect 44 -2065 45 -2063
rect 44 -2071 45 -2069
rect 51 -2065 52 -2063
rect 51 -2071 52 -2069
rect 58 -2065 59 -2063
rect 58 -2071 59 -2069
rect 65 -2065 66 -2063
rect 65 -2071 66 -2069
rect 72 -2065 73 -2063
rect 72 -2071 73 -2069
rect 79 -2065 80 -2063
rect 79 -2071 80 -2069
rect 86 -2065 87 -2063
rect 89 -2065 90 -2063
rect 86 -2071 87 -2069
rect 89 -2071 90 -2069
rect 93 -2065 94 -2063
rect 96 -2065 97 -2063
rect 93 -2071 94 -2069
rect 100 -2065 101 -2063
rect 100 -2071 101 -2069
rect 107 -2065 108 -2063
rect 110 -2065 111 -2063
rect 107 -2071 108 -2069
rect 110 -2071 111 -2069
rect 114 -2065 115 -2063
rect 117 -2065 118 -2063
rect 114 -2071 115 -2069
rect 117 -2071 118 -2069
rect 121 -2065 122 -2063
rect 121 -2071 122 -2069
rect 128 -2065 129 -2063
rect 128 -2071 129 -2069
rect 135 -2065 136 -2063
rect 135 -2071 136 -2069
rect 142 -2065 143 -2063
rect 142 -2071 143 -2069
rect 149 -2065 150 -2063
rect 152 -2065 153 -2063
rect 149 -2071 150 -2069
rect 152 -2071 153 -2069
rect 156 -2065 157 -2063
rect 156 -2071 157 -2069
rect 163 -2065 164 -2063
rect 166 -2065 167 -2063
rect 163 -2071 164 -2069
rect 166 -2071 167 -2069
rect 170 -2065 171 -2063
rect 170 -2071 171 -2069
rect 177 -2065 178 -2063
rect 177 -2071 178 -2069
rect 184 -2065 185 -2063
rect 184 -2071 185 -2069
rect 191 -2065 192 -2063
rect 191 -2071 192 -2069
rect 198 -2065 199 -2063
rect 198 -2071 199 -2069
rect 205 -2065 206 -2063
rect 205 -2071 206 -2069
rect 212 -2065 213 -2063
rect 212 -2071 213 -2069
rect 219 -2065 220 -2063
rect 219 -2071 220 -2069
rect 226 -2065 227 -2063
rect 226 -2071 227 -2069
rect 233 -2065 234 -2063
rect 233 -2071 234 -2069
rect 240 -2065 241 -2063
rect 243 -2065 244 -2063
rect 240 -2071 241 -2069
rect 243 -2071 244 -2069
rect 247 -2065 248 -2063
rect 247 -2071 248 -2069
rect 254 -2065 255 -2063
rect 254 -2071 255 -2069
rect 261 -2065 262 -2063
rect 261 -2071 262 -2069
rect 268 -2065 269 -2063
rect 268 -2071 269 -2069
rect 275 -2065 276 -2063
rect 278 -2065 279 -2063
rect 278 -2071 279 -2069
rect 282 -2065 283 -2063
rect 282 -2071 283 -2069
rect 289 -2065 290 -2063
rect 289 -2071 290 -2069
rect 296 -2065 297 -2063
rect 296 -2071 297 -2069
rect 303 -2065 304 -2063
rect 303 -2071 304 -2069
rect 310 -2065 311 -2063
rect 310 -2071 311 -2069
rect 317 -2065 318 -2063
rect 317 -2071 318 -2069
rect 324 -2071 325 -2069
rect 327 -2071 328 -2069
rect 331 -2065 332 -2063
rect 334 -2065 335 -2063
rect 331 -2071 332 -2069
rect 334 -2071 335 -2069
rect 338 -2065 339 -2063
rect 338 -2071 339 -2069
rect 345 -2065 346 -2063
rect 345 -2071 346 -2069
rect 352 -2065 353 -2063
rect 352 -2071 353 -2069
rect 359 -2065 360 -2063
rect 359 -2071 360 -2069
rect 366 -2065 367 -2063
rect 366 -2071 367 -2069
rect 373 -2065 374 -2063
rect 373 -2071 374 -2069
rect 380 -2071 381 -2069
rect 387 -2065 388 -2063
rect 387 -2071 388 -2069
rect 394 -2065 395 -2063
rect 394 -2071 395 -2069
rect 401 -2065 402 -2063
rect 401 -2071 402 -2069
rect 408 -2065 409 -2063
rect 408 -2071 409 -2069
rect 415 -2065 416 -2063
rect 415 -2071 416 -2069
rect 422 -2065 423 -2063
rect 422 -2071 423 -2069
rect 429 -2065 430 -2063
rect 429 -2071 430 -2069
rect 436 -2065 437 -2063
rect 436 -2071 437 -2069
rect 443 -2065 444 -2063
rect 443 -2071 444 -2069
rect 450 -2065 451 -2063
rect 450 -2071 451 -2069
rect 457 -2065 458 -2063
rect 457 -2071 458 -2069
rect 464 -2065 465 -2063
rect 464 -2071 465 -2069
rect 471 -2065 472 -2063
rect 471 -2071 472 -2069
rect 478 -2065 479 -2063
rect 481 -2065 482 -2063
rect 478 -2071 479 -2069
rect 481 -2071 482 -2069
rect 488 -2065 489 -2063
rect 485 -2071 486 -2069
rect 488 -2071 489 -2069
rect 492 -2065 493 -2063
rect 492 -2071 493 -2069
rect 499 -2065 500 -2063
rect 502 -2065 503 -2063
rect 499 -2071 500 -2069
rect 502 -2071 503 -2069
rect 506 -2065 507 -2063
rect 506 -2071 507 -2069
rect 513 -2065 514 -2063
rect 513 -2071 514 -2069
rect 520 -2065 521 -2063
rect 520 -2071 521 -2069
rect 527 -2065 528 -2063
rect 527 -2071 528 -2069
rect 534 -2065 535 -2063
rect 534 -2071 535 -2069
rect 541 -2065 542 -2063
rect 541 -2071 542 -2069
rect 548 -2065 549 -2063
rect 548 -2071 549 -2069
rect 555 -2065 556 -2063
rect 555 -2071 556 -2069
rect 562 -2065 563 -2063
rect 562 -2071 563 -2069
rect 569 -2065 570 -2063
rect 569 -2071 570 -2069
rect 576 -2065 577 -2063
rect 579 -2065 580 -2063
rect 576 -2071 577 -2069
rect 579 -2071 580 -2069
rect 583 -2065 584 -2063
rect 583 -2071 584 -2069
rect 590 -2065 591 -2063
rect 590 -2071 591 -2069
rect 597 -2065 598 -2063
rect 597 -2071 598 -2069
rect 604 -2065 605 -2063
rect 604 -2071 605 -2069
rect 611 -2065 612 -2063
rect 611 -2071 612 -2069
rect 618 -2065 619 -2063
rect 621 -2065 622 -2063
rect 618 -2071 619 -2069
rect 621 -2071 622 -2069
rect 625 -2065 626 -2063
rect 625 -2071 626 -2069
rect 632 -2065 633 -2063
rect 632 -2071 633 -2069
rect 639 -2065 640 -2063
rect 639 -2071 640 -2069
rect 646 -2065 647 -2063
rect 646 -2071 647 -2069
rect 653 -2065 654 -2063
rect 660 -2065 661 -2063
rect 663 -2065 664 -2063
rect 660 -2071 661 -2069
rect 663 -2071 664 -2069
rect 667 -2065 668 -2063
rect 667 -2071 668 -2069
rect 674 -2065 675 -2063
rect 674 -2071 675 -2069
rect 681 -2065 682 -2063
rect 681 -2071 682 -2069
rect 688 -2065 689 -2063
rect 688 -2071 689 -2069
rect 695 -2065 696 -2063
rect 698 -2065 699 -2063
rect 695 -2071 696 -2069
rect 698 -2071 699 -2069
rect 702 -2065 703 -2063
rect 702 -2071 703 -2069
rect 709 -2065 710 -2063
rect 709 -2071 710 -2069
rect 716 -2065 717 -2063
rect 716 -2071 717 -2069
rect 723 -2065 724 -2063
rect 723 -2071 724 -2069
rect 730 -2065 731 -2063
rect 730 -2071 731 -2069
rect 737 -2065 738 -2063
rect 737 -2071 738 -2069
rect 744 -2065 745 -2063
rect 744 -2071 745 -2069
rect 751 -2065 752 -2063
rect 751 -2071 752 -2069
rect 758 -2065 759 -2063
rect 758 -2071 759 -2069
rect 765 -2065 766 -2063
rect 765 -2071 766 -2069
rect 772 -2065 773 -2063
rect 772 -2071 773 -2069
rect 779 -2065 780 -2063
rect 779 -2071 780 -2069
rect 786 -2065 787 -2063
rect 786 -2071 787 -2069
rect 793 -2065 794 -2063
rect 793 -2071 794 -2069
rect 800 -2065 801 -2063
rect 800 -2071 801 -2069
rect 807 -2065 808 -2063
rect 807 -2071 808 -2069
rect 814 -2065 815 -2063
rect 814 -2071 815 -2069
rect 817 -2071 818 -2069
rect 821 -2065 822 -2063
rect 821 -2071 822 -2069
rect 828 -2065 829 -2063
rect 828 -2071 829 -2069
rect 835 -2065 836 -2063
rect 835 -2071 836 -2069
rect 842 -2065 843 -2063
rect 842 -2071 843 -2069
rect 849 -2065 850 -2063
rect 849 -2071 850 -2069
rect 856 -2065 857 -2063
rect 856 -2071 857 -2069
rect 863 -2065 864 -2063
rect 863 -2071 864 -2069
rect 866 -2071 867 -2069
rect 870 -2065 871 -2063
rect 870 -2071 871 -2069
rect 877 -2065 878 -2063
rect 877 -2071 878 -2069
rect 884 -2065 885 -2063
rect 884 -2071 885 -2069
rect 891 -2065 892 -2063
rect 891 -2071 892 -2069
rect 898 -2065 899 -2063
rect 898 -2071 899 -2069
rect 905 -2065 906 -2063
rect 905 -2071 906 -2069
rect 912 -2065 913 -2063
rect 912 -2071 913 -2069
rect 919 -2065 920 -2063
rect 919 -2071 920 -2069
rect 926 -2065 927 -2063
rect 926 -2071 927 -2069
rect 933 -2065 934 -2063
rect 933 -2071 934 -2069
rect 940 -2065 941 -2063
rect 940 -2071 941 -2069
rect 947 -2065 948 -2063
rect 947 -2071 948 -2069
rect 954 -2065 955 -2063
rect 954 -2071 955 -2069
rect 961 -2065 962 -2063
rect 961 -2071 962 -2069
rect 968 -2065 969 -2063
rect 971 -2065 972 -2063
rect 968 -2071 969 -2069
rect 975 -2065 976 -2063
rect 975 -2071 976 -2069
rect 982 -2065 983 -2063
rect 982 -2071 983 -2069
rect 989 -2065 990 -2063
rect 989 -2071 990 -2069
rect 996 -2065 997 -2063
rect 996 -2071 997 -2069
rect 1003 -2065 1004 -2063
rect 1003 -2071 1004 -2069
rect 1010 -2065 1011 -2063
rect 1010 -2071 1011 -2069
rect 1017 -2065 1018 -2063
rect 1017 -2071 1018 -2069
rect 1024 -2065 1025 -2063
rect 1027 -2065 1028 -2063
rect 1031 -2065 1032 -2063
rect 1031 -2071 1032 -2069
rect 1038 -2065 1039 -2063
rect 1038 -2071 1039 -2069
rect 1045 -2065 1046 -2063
rect 1045 -2071 1046 -2069
rect 1052 -2065 1053 -2063
rect 1052 -2071 1053 -2069
rect 1059 -2065 1060 -2063
rect 1059 -2071 1060 -2069
rect 1066 -2065 1067 -2063
rect 1066 -2071 1067 -2069
rect 1073 -2065 1074 -2063
rect 1073 -2071 1074 -2069
rect 1080 -2065 1081 -2063
rect 1080 -2071 1081 -2069
rect 1087 -2065 1088 -2063
rect 1087 -2071 1088 -2069
rect 1094 -2065 1095 -2063
rect 1094 -2071 1095 -2069
rect 1101 -2065 1102 -2063
rect 1101 -2071 1102 -2069
rect 1108 -2065 1109 -2063
rect 1108 -2071 1109 -2069
rect 1115 -2065 1116 -2063
rect 1115 -2071 1116 -2069
rect 1122 -2065 1123 -2063
rect 1122 -2071 1123 -2069
rect 1129 -2065 1130 -2063
rect 1129 -2071 1130 -2069
rect 1136 -2065 1137 -2063
rect 1136 -2071 1137 -2069
rect 1139 -2071 1140 -2069
rect 1143 -2065 1144 -2063
rect 1143 -2071 1144 -2069
rect 1150 -2065 1151 -2063
rect 1150 -2071 1151 -2069
rect 1157 -2065 1158 -2063
rect 1157 -2071 1158 -2069
rect 1185 -2065 1186 -2063
rect 1185 -2071 1186 -2069
rect 23 -2150 24 -2148
rect 23 -2156 24 -2154
rect 30 -2150 31 -2148
rect 30 -2156 31 -2154
rect 37 -2150 38 -2148
rect 37 -2156 38 -2154
rect 44 -2150 45 -2148
rect 44 -2156 45 -2154
rect 51 -2150 52 -2148
rect 51 -2156 52 -2154
rect 58 -2150 59 -2148
rect 58 -2156 59 -2154
rect 65 -2150 66 -2148
rect 65 -2156 66 -2154
rect 72 -2150 73 -2148
rect 72 -2156 73 -2154
rect 79 -2150 80 -2148
rect 79 -2156 80 -2154
rect 86 -2150 87 -2148
rect 86 -2156 87 -2154
rect 93 -2150 94 -2148
rect 96 -2150 97 -2148
rect 93 -2156 94 -2154
rect 96 -2156 97 -2154
rect 100 -2150 101 -2148
rect 103 -2150 104 -2148
rect 100 -2156 101 -2154
rect 103 -2156 104 -2154
rect 107 -2150 108 -2148
rect 107 -2156 108 -2154
rect 114 -2150 115 -2148
rect 117 -2150 118 -2148
rect 114 -2156 115 -2154
rect 117 -2156 118 -2154
rect 121 -2150 122 -2148
rect 121 -2156 122 -2154
rect 128 -2150 129 -2148
rect 128 -2156 129 -2154
rect 135 -2150 136 -2148
rect 138 -2150 139 -2148
rect 135 -2156 136 -2154
rect 138 -2156 139 -2154
rect 142 -2150 143 -2148
rect 142 -2156 143 -2154
rect 149 -2150 150 -2148
rect 149 -2156 150 -2154
rect 156 -2150 157 -2148
rect 156 -2156 157 -2154
rect 163 -2150 164 -2148
rect 163 -2156 164 -2154
rect 173 -2150 174 -2148
rect 170 -2156 171 -2154
rect 177 -2150 178 -2148
rect 177 -2156 178 -2154
rect 184 -2150 185 -2148
rect 184 -2156 185 -2154
rect 191 -2150 192 -2148
rect 191 -2156 192 -2154
rect 198 -2150 199 -2148
rect 198 -2156 199 -2154
rect 205 -2150 206 -2148
rect 205 -2156 206 -2154
rect 212 -2150 213 -2148
rect 212 -2156 213 -2154
rect 219 -2150 220 -2148
rect 219 -2156 220 -2154
rect 226 -2150 227 -2148
rect 226 -2156 227 -2154
rect 233 -2150 234 -2148
rect 233 -2156 234 -2154
rect 240 -2150 241 -2148
rect 240 -2156 241 -2154
rect 247 -2150 248 -2148
rect 247 -2156 248 -2154
rect 254 -2150 255 -2148
rect 254 -2156 255 -2154
rect 261 -2150 262 -2148
rect 261 -2156 262 -2154
rect 268 -2150 269 -2148
rect 268 -2156 269 -2154
rect 275 -2150 276 -2148
rect 275 -2156 276 -2154
rect 282 -2150 283 -2148
rect 282 -2156 283 -2154
rect 289 -2150 290 -2148
rect 289 -2156 290 -2154
rect 299 -2150 300 -2148
rect 296 -2156 297 -2154
rect 299 -2156 300 -2154
rect 303 -2150 304 -2148
rect 303 -2156 304 -2154
rect 310 -2150 311 -2148
rect 310 -2156 311 -2154
rect 317 -2150 318 -2148
rect 320 -2150 321 -2148
rect 320 -2156 321 -2154
rect 324 -2150 325 -2148
rect 324 -2156 325 -2154
rect 331 -2150 332 -2148
rect 331 -2156 332 -2154
rect 338 -2150 339 -2148
rect 338 -2156 339 -2154
rect 345 -2150 346 -2148
rect 345 -2156 346 -2154
rect 352 -2150 353 -2148
rect 352 -2156 353 -2154
rect 359 -2150 360 -2148
rect 359 -2156 360 -2154
rect 366 -2150 367 -2148
rect 366 -2156 367 -2154
rect 373 -2150 374 -2148
rect 373 -2156 374 -2154
rect 380 -2150 381 -2148
rect 380 -2156 381 -2154
rect 387 -2150 388 -2148
rect 387 -2156 388 -2154
rect 394 -2150 395 -2148
rect 394 -2156 395 -2154
rect 401 -2150 402 -2148
rect 401 -2156 402 -2154
rect 408 -2150 409 -2148
rect 408 -2156 409 -2154
rect 415 -2150 416 -2148
rect 415 -2156 416 -2154
rect 422 -2150 423 -2148
rect 422 -2156 423 -2154
rect 429 -2150 430 -2148
rect 429 -2156 430 -2154
rect 436 -2150 437 -2148
rect 436 -2156 437 -2154
rect 443 -2150 444 -2148
rect 443 -2156 444 -2154
rect 450 -2150 451 -2148
rect 450 -2156 451 -2154
rect 457 -2150 458 -2148
rect 457 -2156 458 -2154
rect 464 -2150 465 -2148
rect 467 -2150 468 -2148
rect 464 -2156 465 -2154
rect 467 -2156 468 -2154
rect 471 -2150 472 -2148
rect 471 -2156 472 -2154
rect 478 -2150 479 -2148
rect 481 -2150 482 -2148
rect 478 -2156 479 -2154
rect 485 -2150 486 -2148
rect 485 -2156 486 -2154
rect 488 -2156 489 -2154
rect 492 -2150 493 -2148
rect 492 -2156 493 -2154
rect 499 -2150 500 -2148
rect 499 -2156 500 -2154
rect 509 -2150 510 -2148
rect 506 -2156 507 -2154
rect 509 -2156 510 -2154
rect 513 -2150 514 -2148
rect 516 -2150 517 -2148
rect 513 -2156 514 -2154
rect 516 -2156 517 -2154
rect 520 -2150 521 -2148
rect 520 -2156 521 -2154
rect 527 -2150 528 -2148
rect 530 -2150 531 -2148
rect 527 -2156 528 -2154
rect 534 -2150 535 -2148
rect 534 -2156 535 -2154
rect 541 -2150 542 -2148
rect 541 -2156 542 -2154
rect 548 -2150 549 -2148
rect 548 -2156 549 -2154
rect 555 -2150 556 -2148
rect 555 -2156 556 -2154
rect 562 -2150 563 -2148
rect 562 -2156 563 -2154
rect 569 -2150 570 -2148
rect 569 -2156 570 -2154
rect 576 -2150 577 -2148
rect 576 -2156 577 -2154
rect 583 -2150 584 -2148
rect 583 -2156 584 -2154
rect 590 -2150 591 -2148
rect 590 -2156 591 -2154
rect 597 -2150 598 -2148
rect 600 -2150 601 -2148
rect 597 -2156 598 -2154
rect 600 -2156 601 -2154
rect 604 -2150 605 -2148
rect 604 -2156 605 -2154
rect 611 -2150 612 -2148
rect 614 -2150 615 -2148
rect 611 -2156 612 -2154
rect 614 -2156 615 -2154
rect 618 -2150 619 -2148
rect 618 -2156 619 -2154
rect 625 -2150 626 -2148
rect 625 -2156 626 -2154
rect 632 -2150 633 -2148
rect 632 -2156 633 -2154
rect 639 -2150 640 -2148
rect 642 -2150 643 -2148
rect 646 -2150 647 -2148
rect 646 -2156 647 -2154
rect 653 -2150 654 -2148
rect 656 -2150 657 -2148
rect 653 -2156 654 -2154
rect 656 -2156 657 -2154
rect 660 -2150 661 -2148
rect 660 -2156 661 -2154
rect 667 -2150 668 -2148
rect 667 -2156 668 -2154
rect 674 -2150 675 -2148
rect 674 -2156 675 -2154
rect 681 -2150 682 -2148
rect 681 -2156 682 -2154
rect 688 -2150 689 -2148
rect 691 -2150 692 -2148
rect 688 -2156 689 -2154
rect 691 -2156 692 -2154
rect 695 -2150 696 -2148
rect 695 -2156 696 -2154
rect 702 -2150 703 -2148
rect 702 -2156 703 -2154
rect 709 -2150 710 -2148
rect 709 -2156 710 -2154
rect 716 -2150 717 -2148
rect 716 -2156 717 -2154
rect 723 -2150 724 -2148
rect 723 -2156 724 -2154
rect 730 -2150 731 -2148
rect 730 -2156 731 -2154
rect 737 -2150 738 -2148
rect 737 -2156 738 -2154
rect 744 -2150 745 -2148
rect 744 -2156 745 -2154
rect 751 -2150 752 -2148
rect 751 -2156 752 -2154
rect 758 -2150 759 -2148
rect 758 -2156 759 -2154
rect 765 -2150 766 -2148
rect 765 -2156 766 -2154
rect 772 -2150 773 -2148
rect 772 -2156 773 -2154
rect 779 -2150 780 -2148
rect 779 -2156 780 -2154
rect 786 -2150 787 -2148
rect 789 -2150 790 -2148
rect 786 -2156 787 -2154
rect 789 -2156 790 -2154
rect 793 -2150 794 -2148
rect 793 -2156 794 -2154
rect 800 -2150 801 -2148
rect 800 -2156 801 -2154
rect 807 -2150 808 -2148
rect 807 -2156 808 -2154
rect 814 -2150 815 -2148
rect 814 -2156 815 -2154
rect 821 -2150 822 -2148
rect 821 -2156 822 -2154
rect 828 -2150 829 -2148
rect 828 -2156 829 -2154
rect 835 -2150 836 -2148
rect 835 -2156 836 -2154
rect 842 -2150 843 -2148
rect 842 -2156 843 -2154
rect 849 -2150 850 -2148
rect 849 -2156 850 -2154
rect 856 -2150 857 -2148
rect 856 -2156 857 -2154
rect 863 -2150 864 -2148
rect 863 -2156 864 -2154
rect 870 -2150 871 -2148
rect 870 -2156 871 -2154
rect 877 -2150 878 -2148
rect 877 -2156 878 -2154
rect 884 -2150 885 -2148
rect 884 -2156 885 -2154
rect 891 -2150 892 -2148
rect 891 -2156 892 -2154
rect 898 -2150 899 -2148
rect 898 -2156 899 -2154
rect 905 -2150 906 -2148
rect 905 -2156 906 -2154
rect 912 -2150 913 -2148
rect 912 -2156 913 -2154
rect 919 -2150 920 -2148
rect 919 -2156 920 -2154
rect 926 -2150 927 -2148
rect 926 -2156 927 -2154
rect 933 -2150 934 -2148
rect 933 -2156 934 -2154
rect 940 -2150 941 -2148
rect 940 -2156 941 -2154
rect 947 -2150 948 -2148
rect 947 -2156 948 -2154
rect 954 -2150 955 -2148
rect 954 -2156 955 -2154
rect 961 -2150 962 -2148
rect 961 -2156 962 -2154
rect 968 -2150 969 -2148
rect 971 -2156 972 -2154
rect 975 -2150 976 -2148
rect 975 -2156 976 -2154
rect 982 -2150 983 -2148
rect 982 -2156 983 -2154
rect 989 -2150 990 -2148
rect 989 -2156 990 -2154
rect 996 -2150 997 -2148
rect 996 -2156 997 -2154
rect 1003 -2150 1004 -2148
rect 1003 -2156 1004 -2154
rect 1010 -2150 1011 -2148
rect 1010 -2156 1011 -2154
rect 1017 -2150 1018 -2148
rect 1017 -2156 1018 -2154
rect 1024 -2150 1025 -2148
rect 1024 -2156 1025 -2154
rect 1031 -2150 1032 -2148
rect 1031 -2156 1032 -2154
rect 1038 -2150 1039 -2148
rect 1038 -2156 1039 -2154
rect 1045 -2150 1046 -2148
rect 1045 -2156 1046 -2154
rect 1052 -2150 1053 -2148
rect 1052 -2156 1053 -2154
rect 1059 -2150 1060 -2148
rect 1059 -2156 1060 -2154
rect 1066 -2150 1067 -2148
rect 1066 -2156 1067 -2154
rect 1101 -2150 1102 -2148
rect 1104 -2150 1105 -2148
rect 1101 -2156 1102 -2154
rect 1104 -2156 1105 -2154
rect 1108 -2150 1109 -2148
rect 1108 -2156 1109 -2154
rect 1122 -2150 1123 -2148
rect 1122 -2156 1123 -2154
rect 30 -2231 31 -2229
rect 30 -2237 31 -2235
rect 37 -2231 38 -2229
rect 37 -2237 38 -2235
rect 44 -2231 45 -2229
rect 44 -2237 45 -2235
rect 51 -2231 52 -2229
rect 51 -2237 52 -2235
rect 58 -2231 59 -2229
rect 65 -2231 66 -2229
rect 65 -2237 66 -2235
rect 72 -2231 73 -2229
rect 72 -2237 73 -2235
rect 79 -2231 80 -2229
rect 86 -2231 87 -2229
rect 89 -2237 90 -2235
rect 93 -2231 94 -2229
rect 96 -2231 97 -2229
rect 93 -2237 94 -2235
rect 96 -2237 97 -2235
rect 100 -2231 101 -2229
rect 100 -2237 101 -2235
rect 107 -2231 108 -2229
rect 107 -2237 108 -2235
rect 114 -2231 115 -2229
rect 114 -2237 115 -2235
rect 121 -2231 122 -2229
rect 124 -2231 125 -2229
rect 121 -2237 122 -2235
rect 124 -2237 125 -2235
rect 128 -2231 129 -2229
rect 131 -2231 132 -2229
rect 128 -2237 129 -2235
rect 131 -2237 132 -2235
rect 135 -2231 136 -2229
rect 135 -2237 136 -2235
rect 142 -2231 143 -2229
rect 142 -2237 143 -2235
rect 149 -2231 150 -2229
rect 149 -2237 150 -2235
rect 156 -2231 157 -2229
rect 156 -2237 157 -2235
rect 163 -2231 164 -2229
rect 163 -2237 164 -2235
rect 170 -2231 171 -2229
rect 170 -2237 171 -2235
rect 177 -2231 178 -2229
rect 180 -2231 181 -2229
rect 177 -2237 178 -2235
rect 180 -2237 181 -2235
rect 184 -2231 185 -2229
rect 184 -2237 185 -2235
rect 191 -2231 192 -2229
rect 191 -2237 192 -2235
rect 198 -2231 199 -2229
rect 198 -2237 199 -2235
rect 205 -2231 206 -2229
rect 205 -2237 206 -2235
rect 212 -2231 213 -2229
rect 212 -2237 213 -2235
rect 219 -2231 220 -2229
rect 219 -2237 220 -2235
rect 226 -2231 227 -2229
rect 226 -2237 227 -2235
rect 233 -2231 234 -2229
rect 233 -2237 234 -2235
rect 240 -2231 241 -2229
rect 240 -2237 241 -2235
rect 247 -2231 248 -2229
rect 247 -2237 248 -2235
rect 254 -2231 255 -2229
rect 254 -2237 255 -2235
rect 261 -2231 262 -2229
rect 261 -2237 262 -2235
rect 268 -2231 269 -2229
rect 268 -2237 269 -2235
rect 275 -2231 276 -2229
rect 275 -2237 276 -2235
rect 282 -2231 283 -2229
rect 282 -2237 283 -2235
rect 289 -2231 290 -2229
rect 289 -2237 290 -2235
rect 296 -2231 297 -2229
rect 296 -2237 297 -2235
rect 303 -2231 304 -2229
rect 303 -2237 304 -2235
rect 310 -2231 311 -2229
rect 310 -2237 311 -2235
rect 317 -2231 318 -2229
rect 317 -2237 318 -2235
rect 324 -2231 325 -2229
rect 324 -2237 325 -2235
rect 331 -2231 332 -2229
rect 331 -2237 332 -2235
rect 338 -2231 339 -2229
rect 338 -2237 339 -2235
rect 345 -2231 346 -2229
rect 345 -2237 346 -2235
rect 355 -2231 356 -2229
rect 352 -2237 353 -2235
rect 355 -2237 356 -2235
rect 359 -2231 360 -2229
rect 359 -2237 360 -2235
rect 366 -2231 367 -2229
rect 366 -2237 367 -2235
rect 373 -2231 374 -2229
rect 373 -2237 374 -2235
rect 380 -2231 381 -2229
rect 380 -2237 381 -2235
rect 387 -2231 388 -2229
rect 387 -2237 388 -2235
rect 394 -2231 395 -2229
rect 397 -2231 398 -2229
rect 394 -2237 395 -2235
rect 397 -2237 398 -2235
rect 401 -2231 402 -2229
rect 401 -2237 402 -2235
rect 408 -2231 409 -2229
rect 408 -2237 409 -2235
rect 415 -2231 416 -2229
rect 415 -2237 416 -2235
rect 422 -2231 423 -2229
rect 422 -2237 423 -2235
rect 429 -2231 430 -2229
rect 429 -2237 430 -2235
rect 436 -2231 437 -2229
rect 436 -2237 437 -2235
rect 443 -2231 444 -2229
rect 443 -2237 444 -2235
rect 446 -2237 447 -2235
rect 450 -2231 451 -2229
rect 453 -2231 454 -2229
rect 450 -2237 451 -2235
rect 453 -2237 454 -2235
rect 457 -2231 458 -2229
rect 457 -2237 458 -2235
rect 464 -2231 465 -2229
rect 464 -2237 465 -2235
rect 471 -2231 472 -2229
rect 471 -2237 472 -2235
rect 481 -2231 482 -2229
rect 478 -2237 479 -2235
rect 481 -2237 482 -2235
rect 485 -2231 486 -2229
rect 488 -2231 489 -2229
rect 485 -2237 486 -2235
rect 492 -2231 493 -2229
rect 492 -2237 493 -2235
rect 499 -2231 500 -2229
rect 499 -2237 500 -2235
rect 506 -2231 507 -2229
rect 506 -2237 507 -2235
rect 513 -2231 514 -2229
rect 513 -2237 514 -2235
rect 520 -2231 521 -2229
rect 520 -2237 521 -2235
rect 527 -2231 528 -2229
rect 530 -2231 531 -2229
rect 527 -2237 528 -2235
rect 530 -2237 531 -2235
rect 534 -2231 535 -2229
rect 534 -2237 535 -2235
rect 541 -2231 542 -2229
rect 541 -2237 542 -2235
rect 548 -2231 549 -2229
rect 548 -2237 549 -2235
rect 555 -2231 556 -2229
rect 555 -2237 556 -2235
rect 562 -2231 563 -2229
rect 562 -2237 563 -2235
rect 569 -2231 570 -2229
rect 569 -2237 570 -2235
rect 576 -2231 577 -2229
rect 576 -2237 577 -2235
rect 583 -2231 584 -2229
rect 583 -2237 584 -2235
rect 590 -2231 591 -2229
rect 590 -2237 591 -2235
rect 597 -2231 598 -2229
rect 604 -2231 605 -2229
rect 604 -2237 605 -2235
rect 611 -2231 612 -2229
rect 611 -2237 612 -2235
rect 618 -2231 619 -2229
rect 618 -2237 619 -2235
rect 625 -2231 626 -2229
rect 625 -2237 626 -2235
rect 632 -2231 633 -2229
rect 632 -2237 633 -2235
rect 639 -2231 640 -2229
rect 639 -2237 640 -2235
rect 646 -2231 647 -2229
rect 646 -2237 647 -2235
rect 653 -2231 654 -2229
rect 656 -2231 657 -2229
rect 653 -2237 654 -2235
rect 656 -2237 657 -2235
rect 660 -2231 661 -2229
rect 660 -2237 661 -2235
rect 667 -2231 668 -2229
rect 670 -2231 671 -2229
rect 667 -2237 668 -2235
rect 670 -2237 671 -2235
rect 674 -2231 675 -2229
rect 674 -2237 675 -2235
rect 681 -2231 682 -2229
rect 681 -2237 682 -2235
rect 684 -2237 685 -2235
rect 688 -2231 689 -2229
rect 688 -2237 689 -2235
rect 695 -2231 696 -2229
rect 698 -2231 699 -2229
rect 698 -2237 699 -2235
rect 702 -2231 703 -2229
rect 702 -2237 703 -2235
rect 709 -2231 710 -2229
rect 709 -2237 710 -2235
rect 716 -2231 717 -2229
rect 716 -2237 717 -2235
rect 723 -2231 724 -2229
rect 723 -2237 724 -2235
rect 730 -2231 731 -2229
rect 730 -2237 731 -2235
rect 740 -2231 741 -2229
rect 737 -2237 738 -2235
rect 740 -2237 741 -2235
rect 747 -2231 748 -2229
rect 744 -2237 745 -2235
rect 747 -2237 748 -2235
rect 751 -2231 752 -2229
rect 751 -2237 752 -2235
rect 758 -2231 759 -2229
rect 758 -2237 759 -2235
rect 765 -2231 766 -2229
rect 765 -2237 766 -2235
rect 772 -2231 773 -2229
rect 772 -2237 773 -2235
rect 779 -2231 780 -2229
rect 779 -2237 780 -2235
rect 786 -2231 787 -2229
rect 786 -2237 787 -2235
rect 793 -2231 794 -2229
rect 793 -2237 794 -2235
rect 800 -2231 801 -2229
rect 800 -2237 801 -2235
rect 807 -2231 808 -2229
rect 807 -2237 808 -2235
rect 810 -2237 811 -2235
rect 814 -2231 815 -2229
rect 814 -2237 815 -2235
rect 821 -2231 822 -2229
rect 821 -2237 822 -2235
rect 828 -2231 829 -2229
rect 828 -2237 829 -2235
rect 835 -2231 836 -2229
rect 835 -2237 836 -2235
rect 842 -2231 843 -2229
rect 842 -2237 843 -2235
rect 849 -2231 850 -2229
rect 849 -2237 850 -2235
rect 856 -2231 857 -2229
rect 856 -2237 857 -2235
rect 863 -2231 864 -2229
rect 863 -2237 864 -2235
rect 870 -2231 871 -2229
rect 870 -2237 871 -2235
rect 877 -2231 878 -2229
rect 877 -2237 878 -2235
rect 884 -2231 885 -2229
rect 884 -2237 885 -2235
rect 891 -2231 892 -2229
rect 891 -2237 892 -2235
rect 898 -2231 899 -2229
rect 898 -2237 899 -2235
rect 905 -2231 906 -2229
rect 905 -2237 906 -2235
rect 912 -2231 913 -2229
rect 912 -2237 913 -2235
rect 919 -2231 920 -2229
rect 919 -2237 920 -2235
rect 926 -2231 927 -2229
rect 926 -2237 927 -2235
rect 933 -2231 934 -2229
rect 933 -2237 934 -2235
rect 940 -2231 941 -2229
rect 943 -2231 944 -2229
rect 940 -2237 941 -2235
rect 943 -2237 944 -2235
rect 947 -2231 948 -2229
rect 947 -2237 948 -2235
rect 954 -2231 955 -2229
rect 954 -2237 955 -2235
rect 957 -2237 958 -2235
rect 961 -2231 962 -2229
rect 961 -2237 962 -2235
rect 968 -2231 969 -2229
rect 968 -2237 969 -2235
rect 975 -2231 976 -2229
rect 975 -2237 976 -2235
rect 982 -2231 983 -2229
rect 982 -2237 983 -2235
rect 996 -2231 997 -2229
rect 996 -2237 997 -2235
rect 1003 -2231 1004 -2229
rect 1003 -2237 1004 -2235
rect 1017 -2231 1018 -2229
rect 1017 -2237 1018 -2235
rect 1066 -2231 1067 -2229
rect 1066 -2237 1067 -2235
rect 44 -2314 45 -2312
rect 44 -2320 45 -2318
rect 51 -2314 52 -2312
rect 51 -2320 52 -2318
rect 58 -2320 59 -2318
rect 65 -2314 66 -2312
rect 65 -2320 66 -2318
rect 72 -2314 73 -2312
rect 72 -2320 73 -2318
rect 79 -2314 80 -2312
rect 79 -2320 80 -2318
rect 89 -2314 90 -2312
rect 86 -2320 87 -2318
rect 89 -2320 90 -2318
rect 93 -2314 94 -2312
rect 93 -2320 94 -2318
rect 100 -2314 101 -2312
rect 100 -2320 101 -2318
rect 107 -2314 108 -2312
rect 107 -2320 108 -2318
rect 114 -2314 115 -2312
rect 114 -2320 115 -2318
rect 121 -2314 122 -2312
rect 121 -2320 122 -2318
rect 128 -2314 129 -2312
rect 128 -2320 129 -2318
rect 135 -2314 136 -2312
rect 138 -2314 139 -2312
rect 138 -2320 139 -2318
rect 142 -2314 143 -2312
rect 142 -2320 143 -2318
rect 149 -2314 150 -2312
rect 149 -2320 150 -2318
rect 156 -2314 157 -2312
rect 156 -2320 157 -2318
rect 163 -2314 164 -2312
rect 163 -2320 164 -2318
rect 170 -2314 171 -2312
rect 170 -2320 171 -2318
rect 177 -2314 178 -2312
rect 177 -2320 178 -2318
rect 184 -2314 185 -2312
rect 187 -2314 188 -2312
rect 184 -2320 185 -2318
rect 191 -2314 192 -2312
rect 191 -2320 192 -2318
rect 198 -2314 199 -2312
rect 198 -2320 199 -2318
rect 205 -2314 206 -2312
rect 205 -2320 206 -2318
rect 212 -2314 213 -2312
rect 212 -2320 213 -2318
rect 219 -2314 220 -2312
rect 219 -2320 220 -2318
rect 226 -2314 227 -2312
rect 226 -2320 227 -2318
rect 233 -2314 234 -2312
rect 233 -2320 234 -2318
rect 240 -2314 241 -2312
rect 240 -2320 241 -2318
rect 247 -2314 248 -2312
rect 247 -2320 248 -2318
rect 254 -2314 255 -2312
rect 254 -2320 255 -2318
rect 261 -2314 262 -2312
rect 261 -2320 262 -2318
rect 268 -2314 269 -2312
rect 268 -2320 269 -2318
rect 275 -2314 276 -2312
rect 275 -2320 276 -2318
rect 282 -2314 283 -2312
rect 282 -2320 283 -2318
rect 292 -2314 293 -2312
rect 289 -2320 290 -2318
rect 292 -2320 293 -2318
rect 296 -2314 297 -2312
rect 296 -2320 297 -2318
rect 303 -2314 304 -2312
rect 303 -2320 304 -2318
rect 310 -2314 311 -2312
rect 310 -2320 311 -2318
rect 317 -2314 318 -2312
rect 317 -2320 318 -2318
rect 324 -2314 325 -2312
rect 324 -2320 325 -2318
rect 331 -2314 332 -2312
rect 331 -2320 332 -2318
rect 338 -2314 339 -2312
rect 338 -2320 339 -2318
rect 345 -2314 346 -2312
rect 348 -2314 349 -2312
rect 345 -2320 346 -2318
rect 348 -2320 349 -2318
rect 352 -2314 353 -2312
rect 352 -2320 353 -2318
rect 359 -2314 360 -2312
rect 359 -2320 360 -2318
rect 366 -2314 367 -2312
rect 366 -2320 367 -2318
rect 373 -2314 374 -2312
rect 376 -2314 377 -2312
rect 373 -2320 374 -2318
rect 376 -2320 377 -2318
rect 380 -2314 381 -2312
rect 380 -2320 381 -2318
rect 387 -2314 388 -2312
rect 387 -2320 388 -2318
rect 394 -2314 395 -2312
rect 394 -2320 395 -2318
rect 401 -2314 402 -2312
rect 401 -2320 402 -2318
rect 408 -2314 409 -2312
rect 408 -2320 409 -2318
rect 415 -2314 416 -2312
rect 415 -2320 416 -2318
rect 422 -2314 423 -2312
rect 422 -2320 423 -2318
rect 425 -2320 426 -2318
rect 429 -2314 430 -2312
rect 429 -2320 430 -2318
rect 436 -2314 437 -2312
rect 436 -2320 437 -2318
rect 443 -2314 444 -2312
rect 446 -2314 447 -2312
rect 443 -2320 444 -2318
rect 446 -2320 447 -2318
rect 453 -2314 454 -2312
rect 450 -2320 451 -2318
rect 453 -2320 454 -2318
rect 457 -2314 458 -2312
rect 457 -2320 458 -2318
rect 464 -2314 465 -2312
rect 464 -2320 465 -2318
rect 471 -2314 472 -2312
rect 471 -2320 472 -2318
rect 478 -2314 479 -2312
rect 478 -2320 479 -2318
rect 485 -2314 486 -2312
rect 485 -2320 486 -2318
rect 492 -2314 493 -2312
rect 492 -2320 493 -2318
rect 495 -2320 496 -2318
rect 499 -2314 500 -2312
rect 499 -2320 500 -2318
rect 506 -2314 507 -2312
rect 506 -2320 507 -2318
rect 513 -2314 514 -2312
rect 513 -2320 514 -2318
rect 520 -2314 521 -2312
rect 520 -2320 521 -2318
rect 527 -2314 528 -2312
rect 527 -2320 528 -2318
rect 534 -2314 535 -2312
rect 537 -2314 538 -2312
rect 534 -2320 535 -2318
rect 541 -2314 542 -2312
rect 541 -2320 542 -2318
rect 548 -2314 549 -2312
rect 548 -2320 549 -2318
rect 555 -2314 556 -2312
rect 555 -2320 556 -2318
rect 562 -2314 563 -2312
rect 565 -2314 566 -2312
rect 562 -2320 563 -2318
rect 565 -2320 566 -2318
rect 569 -2314 570 -2312
rect 572 -2314 573 -2312
rect 569 -2320 570 -2318
rect 572 -2320 573 -2318
rect 576 -2314 577 -2312
rect 579 -2314 580 -2312
rect 576 -2320 577 -2318
rect 583 -2314 584 -2312
rect 583 -2320 584 -2318
rect 590 -2314 591 -2312
rect 590 -2320 591 -2318
rect 597 -2320 598 -2318
rect 604 -2314 605 -2312
rect 604 -2320 605 -2318
rect 611 -2314 612 -2312
rect 611 -2320 612 -2318
rect 618 -2314 619 -2312
rect 621 -2314 622 -2312
rect 618 -2320 619 -2318
rect 621 -2320 622 -2318
rect 625 -2314 626 -2312
rect 625 -2320 626 -2318
rect 632 -2314 633 -2312
rect 632 -2320 633 -2318
rect 639 -2314 640 -2312
rect 639 -2320 640 -2318
rect 646 -2314 647 -2312
rect 653 -2314 654 -2312
rect 656 -2314 657 -2312
rect 653 -2320 654 -2318
rect 656 -2320 657 -2318
rect 660 -2314 661 -2312
rect 660 -2320 661 -2318
rect 667 -2314 668 -2312
rect 667 -2320 668 -2318
rect 674 -2314 675 -2312
rect 674 -2320 675 -2318
rect 681 -2314 682 -2312
rect 684 -2314 685 -2312
rect 681 -2320 682 -2318
rect 688 -2314 689 -2312
rect 688 -2320 689 -2318
rect 695 -2314 696 -2312
rect 695 -2320 696 -2318
rect 702 -2314 703 -2312
rect 702 -2320 703 -2318
rect 709 -2314 710 -2312
rect 709 -2320 710 -2318
rect 716 -2314 717 -2312
rect 716 -2320 717 -2318
rect 719 -2320 720 -2318
rect 723 -2314 724 -2312
rect 723 -2320 724 -2318
rect 730 -2314 731 -2312
rect 730 -2320 731 -2318
rect 737 -2314 738 -2312
rect 737 -2320 738 -2318
rect 744 -2314 745 -2312
rect 744 -2320 745 -2318
rect 751 -2314 752 -2312
rect 751 -2320 752 -2318
rect 758 -2314 759 -2312
rect 758 -2320 759 -2318
rect 765 -2314 766 -2312
rect 765 -2320 766 -2318
rect 772 -2314 773 -2312
rect 772 -2320 773 -2318
rect 779 -2314 780 -2312
rect 779 -2320 780 -2318
rect 786 -2314 787 -2312
rect 786 -2320 787 -2318
rect 793 -2314 794 -2312
rect 793 -2320 794 -2318
rect 800 -2314 801 -2312
rect 803 -2314 804 -2312
rect 803 -2320 804 -2318
rect 807 -2314 808 -2312
rect 810 -2314 811 -2312
rect 807 -2320 808 -2318
rect 814 -2314 815 -2312
rect 814 -2320 815 -2318
rect 821 -2314 822 -2312
rect 821 -2320 822 -2318
rect 828 -2314 829 -2312
rect 828 -2320 829 -2318
rect 835 -2314 836 -2312
rect 835 -2320 836 -2318
rect 842 -2314 843 -2312
rect 842 -2320 843 -2318
rect 849 -2314 850 -2312
rect 849 -2320 850 -2318
rect 856 -2314 857 -2312
rect 856 -2320 857 -2318
rect 863 -2314 864 -2312
rect 863 -2320 864 -2318
rect 870 -2314 871 -2312
rect 870 -2320 871 -2318
rect 877 -2314 878 -2312
rect 877 -2320 878 -2318
rect 884 -2314 885 -2312
rect 884 -2320 885 -2318
rect 891 -2314 892 -2312
rect 891 -2320 892 -2318
rect 898 -2314 899 -2312
rect 898 -2320 899 -2318
rect 968 -2314 969 -2312
rect 968 -2320 969 -2318
rect 989 -2314 990 -2312
rect 989 -2320 990 -2318
rect 996 -2314 997 -2312
rect 996 -2320 997 -2318
rect 1038 -2314 1039 -2312
rect 1038 -2320 1039 -2318
rect 1059 -2314 1060 -2312
rect 1059 -2320 1060 -2318
rect 72 -2379 73 -2377
rect 72 -2385 73 -2383
rect 79 -2379 80 -2377
rect 79 -2385 80 -2383
rect 86 -2379 87 -2377
rect 86 -2385 87 -2383
rect 93 -2379 94 -2377
rect 93 -2385 94 -2383
rect 100 -2379 101 -2377
rect 100 -2385 101 -2383
rect 107 -2379 108 -2377
rect 107 -2385 108 -2383
rect 114 -2379 115 -2377
rect 114 -2385 115 -2383
rect 121 -2379 122 -2377
rect 121 -2385 122 -2383
rect 128 -2379 129 -2377
rect 128 -2385 129 -2383
rect 135 -2379 136 -2377
rect 135 -2385 136 -2383
rect 142 -2379 143 -2377
rect 142 -2385 143 -2383
rect 149 -2379 150 -2377
rect 152 -2379 153 -2377
rect 149 -2385 150 -2383
rect 156 -2379 157 -2377
rect 156 -2385 157 -2383
rect 163 -2379 164 -2377
rect 163 -2385 164 -2383
rect 166 -2385 167 -2383
rect 170 -2379 171 -2377
rect 173 -2385 174 -2383
rect 177 -2385 178 -2383
rect 184 -2379 185 -2377
rect 187 -2379 188 -2377
rect 184 -2385 185 -2383
rect 187 -2385 188 -2383
rect 191 -2379 192 -2377
rect 191 -2385 192 -2383
rect 198 -2379 199 -2377
rect 198 -2385 199 -2383
rect 205 -2379 206 -2377
rect 205 -2385 206 -2383
rect 212 -2379 213 -2377
rect 212 -2385 213 -2383
rect 219 -2379 220 -2377
rect 219 -2385 220 -2383
rect 226 -2379 227 -2377
rect 226 -2385 227 -2383
rect 233 -2379 234 -2377
rect 236 -2379 237 -2377
rect 233 -2385 234 -2383
rect 236 -2385 237 -2383
rect 240 -2379 241 -2377
rect 240 -2385 241 -2383
rect 247 -2379 248 -2377
rect 247 -2385 248 -2383
rect 254 -2379 255 -2377
rect 254 -2385 255 -2383
rect 261 -2379 262 -2377
rect 261 -2385 262 -2383
rect 271 -2379 272 -2377
rect 268 -2385 269 -2383
rect 275 -2379 276 -2377
rect 275 -2385 276 -2383
rect 282 -2379 283 -2377
rect 282 -2385 283 -2383
rect 289 -2379 290 -2377
rect 289 -2385 290 -2383
rect 296 -2379 297 -2377
rect 296 -2385 297 -2383
rect 303 -2379 304 -2377
rect 306 -2379 307 -2377
rect 303 -2385 304 -2383
rect 306 -2385 307 -2383
rect 310 -2379 311 -2377
rect 310 -2385 311 -2383
rect 317 -2379 318 -2377
rect 317 -2385 318 -2383
rect 324 -2379 325 -2377
rect 324 -2385 325 -2383
rect 331 -2379 332 -2377
rect 331 -2385 332 -2383
rect 338 -2379 339 -2377
rect 338 -2385 339 -2383
rect 345 -2379 346 -2377
rect 345 -2385 346 -2383
rect 352 -2379 353 -2377
rect 352 -2385 353 -2383
rect 359 -2379 360 -2377
rect 359 -2385 360 -2383
rect 366 -2379 367 -2377
rect 366 -2385 367 -2383
rect 373 -2379 374 -2377
rect 373 -2385 374 -2383
rect 383 -2379 384 -2377
rect 380 -2385 381 -2383
rect 383 -2385 384 -2383
rect 387 -2379 388 -2377
rect 387 -2385 388 -2383
rect 394 -2379 395 -2377
rect 394 -2385 395 -2383
rect 401 -2379 402 -2377
rect 401 -2385 402 -2383
rect 408 -2379 409 -2377
rect 408 -2385 409 -2383
rect 415 -2379 416 -2377
rect 415 -2385 416 -2383
rect 422 -2379 423 -2377
rect 422 -2385 423 -2383
rect 429 -2379 430 -2377
rect 429 -2385 430 -2383
rect 436 -2379 437 -2377
rect 436 -2385 437 -2383
rect 443 -2379 444 -2377
rect 443 -2385 444 -2383
rect 450 -2379 451 -2377
rect 450 -2385 451 -2383
rect 453 -2385 454 -2383
rect 457 -2379 458 -2377
rect 457 -2385 458 -2383
rect 464 -2379 465 -2377
rect 464 -2385 465 -2383
rect 471 -2379 472 -2377
rect 471 -2385 472 -2383
rect 478 -2379 479 -2377
rect 478 -2385 479 -2383
rect 485 -2379 486 -2377
rect 485 -2385 486 -2383
rect 492 -2379 493 -2377
rect 492 -2385 493 -2383
rect 499 -2379 500 -2377
rect 499 -2385 500 -2383
rect 506 -2379 507 -2377
rect 506 -2385 507 -2383
rect 513 -2379 514 -2377
rect 516 -2379 517 -2377
rect 513 -2385 514 -2383
rect 516 -2385 517 -2383
rect 520 -2379 521 -2377
rect 520 -2385 521 -2383
rect 527 -2379 528 -2377
rect 530 -2379 531 -2377
rect 530 -2385 531 -2383
rect 534 -2379 535 -2377
rect 534 -2385 535 -2383
rect 541 -2379 542 -2377
rect 541 -2385 542 -2383
rect 548 -2379 549 -2377
rect 548 -2385 549 -2383
rect 555 -2379 556 -2377
rect 558 -2379 559 -2377
rect 555 -2385 556 -2383
rect 558 -2385 559 -2383
rect 562 -2379 563 -2377
rect 562 -2385 563 -2383
rect 569 -2379 570 -2377
rect 569 -2385 570 -2383
rect 576 -2379 577 -2377
rect 576 -2385 577 -2383
rect 583 -2379 584 -2377
rect 583 -2385 584 -2383
rect 590 -2379 591 -2377
rect 590 -2385 591 -2383
rect 597 -2379 598 -2377
rect 597 -2385 598 -2383
rect 604 -2379 605 -2377
rect 604 -2385 605 -2383
rect 611 -2379 612 -2377
rect 614 -2379 615 -2377
rect 611 -2385 612 -2383
rect 614 -2385 615 -2383
rect 618 -2379 619 -2377
rect 618 -2385 619 -2383
rect 625 -2379 626 -2377
rect 625 -2385 626 -2383
rect 632 -2379 633 -2377
rect 632 -2385 633 -2383
rect 639 -2379 640 -2377
rect 639 -2385 640 -2383
rect 646 -2385 647 -2383
rect 653 -2379 654 -2377
rect 653 -2385 654 -2383
rect 660 -2379 661 -2377
rect 660 -2385 661 -2383
rect 667 -2379 668 -2377
rect 667 -2385 668 -2383
rect 674 -2379 675 -2377
rect 674 -2385 675 -2383
rect 681 -2379 682 -2377
rect 681 -2385 682 -2383
rect 688 -2379 689 -2377
rect 688 -2385 689 -2383
rect 695 -2379 696 -2377
rect 698 -2379 699 -2377
rect 698 -2385 699 -2383
rect 702 -2379 703 -2377
rect 702 -2385 703 -2383
rect 709 -2379 710 -2377
rect 709 -2385 710 -2383
rect 716 -2379 717 -2377
rect 719 -2379 720 -2377
rect 716 -2385 717 -2383
rect 730 -2379 731 -2377
rect 730 -2385 731 -2383
rect 737 -2379 738 -2377
rect 737 -2385 738 -2383
rect 744 -2379 745 -2377
rect 744 -2385 745 -2383
rect 751 -2379 752 -2377
rect 751 -2385 752 -2383
rect 758 -2379 759 -2377
rect 758 -2385 759 -2383
rect 765 -2379 766 -2377
rect 765 -2385 766 -2383
rect 772 -2379 773 -2377
rect 772 -2385 773 -2383
rect 779 -2379 780 -2377
rect 779 -2385 780 -2383
rect 793 -2379 794 -2377
rect 793 -2385 794 -2383
rect 800 -2379 801 -2377
rect 800 -2385 801 -2383
rect 814 -2379 815 -2377
rect 814 -2385 815 -2383
rect 898 -2379 899 -2377
rect 898 -2385 899 -2383
rect 905 -2379 906 -2377
rect 905 -2385 906 -2383
rect 940 -2379 941 -2377
rect 940 -2385 941 -2383
rect 978 -2379 979 -2377
rect 975 -2385 976 -2383
rect 978 -2385 979 -2383
rect 982 -2379 983 -2377
rect 982 -2385 983 -2383
rect 989 -2379 990 -2377
rect 989 -2385 990 -2383
rect 1003 -2379 1004 -2377
rect 1006 -2379 1007 -2377
rect 1006 -2385 1007 -2383
rect 198 -2430 199 -2428
rect 198 -2436 199 -2434
rect 219 -2430 220 -2428
rect 219 -2436 220 -2434
rect 226 -2430 227 -2428
rect 226 -2436 227 -2434
rect 233 -2430 234 -2428
rect 233 -2436 234 -2434
rect 240 -2430 241 -2428
rect 240 -2436 241 -2434
rect 247 -2430 248 -2428
rect 254 -2430 255 -2428
rect 254 -2436 255 -2434
rect 261 -2430 262 -2428
rect 261 -2436 262 -2434
rect 268 -2430 269 -2428
rect 268 -2436 269 -2434
rect 275 -2430 276 -2428
rect 275 -2436 276 -2434
rect 282 -2430 283 -2428
rect 282 -2436 283 -2434
rect 289 -2430 290 -2428
rect 289 -2436 290 -2434
rect 296 -2430 297 -2428
rect 296 -2436 297 -2434
rect 303 -2430 304 -2428
rect 303 -2436 304 -2434
rect 310 -2430 311 -2428
rect 310 -2436 311 -2434
rect 317 -2430 318 -2428
rect 317 -2436 318 -2434
rect 324 -2430 325 -2428
rect 327 -2436 328 -2434
rect 331 -2430 332 -2428
rect 331 -2436 332 -2434
rect 338 -2430 339 -2428
rect 338 -2436 339 -2434
rect 345 -2430 346 -2428
rect 345 -2436 346 -2434
rect 355 -2430 356 -2428
rect 352 -2436 353 -2434
rect 359 -2430 360 -2428
rect 359 -2436 360 -2434
rect 369 -2430 370 -2428
rect 366 -2436 367 -2434
rect 369 -2436 370 -2434
rect 373 -2430 374 -2428
rect 373 -2436 374 -2434
rect 380 -2430 381 -2428
rect 383 -2430 384 -2428
rect 380 -2436 381 -2434
rect 387 -2430 388 -2428
rect 387 -2436 388 -2434
rect 394 -2430 395 -2428
rect 394 -2436 395 -2434
rect 401 -2430 402 -2428
rect 401 -2436 402 -2434
rect 408 -2430 409 -2428
rect 408 -2436 409 -2434
rect 418 -2430 419 -2428
rect 415 -2436 416 -2434
rect 418 -2436 419 -2434
rect 422 -2430 423 -2428
rect 422 -2436 423 -2434
rect 429 -2430 430 -2428
rect 429 -2436 430 -2434
rect 436 -2430 437 -2428
rect 436 -2436 437 -2434
rect 443 -2430 444 -2428
rect 443 -2436 444 -2434
rect 450 -2430 451 -2428
rect 450 -2436 451 -2434
rect 453 -2436 454 -2434
rect 460 -2430 461 -2428
rect 457 -2436 458 -2434
rect 460 -2436 461 -2434
rect 464 -2430 465 -2428
rect 464 -2436 465 -2434
rect 471 -2430 472 -2428
rect 471 -2436 472 -2434
rect 478 -2430 479 -2428
rect 478 -2436 479 -2434
rect 488 -2430 489 -2428
rect 485 -2436 486 -2434
rect 492 -2430 493 -2428
rect 492 -2436 493 -2434
rect 499 -2430 500 -2428
rect 499 -2436 500 -2434
rect 506 -2430 507 -2428
rect 509 -2430 510 -2428
rect 506 -2436 507 -2434
rect 509 -2436 510 -2434
rect 513 -2430 514 -2428
rect 516 -2430 517 -2428
rect 516 -2436 517 -2434
rect 520 -2430 521 -2428
rect 523 -2430 524 -2428
rect 523 -2436 524 -2434
rect 527 -2430 528 -2428
rect 527 -2436 528 -2434
rect 534 -2430 535 -2428
rect 534 -2436 535 -2434
rect 541 -2430 542 -2428
rect 541 -2436 542 -2434
rect 548 -2430 549 -2428
rect 548 -2436 549 -2434
rect 555 -2430 556 -2428
rect 555 -2436 556 -2434
rect 562 -2430 563 -2428
rect 562 -2436 563 -2434
rect 569 -2430 570 -2428
rect 569 -2436 570 -2434
rect 572 -2436 573 -2434
rect 576 -2430 577 -2428
rect 576 -2436 577 -2434
rect 583 -2430 584 -2428
rect 583 -2436 584 -2434
rect 590 -2430 591 -2428
rect 590 -2436 591 -2434
rect 597 -2430 598 -2428
rect 597 -2436 598 -2434
rect 604 -2430 605 -2428
rect 604 -2436 605 -2434
rect 611 -2430 612 -2428
rect 611 -2436 612 -2434
rect 618 -2430 619 -2428
rect 618 -2436 619 -2434
rect 625 -2430 626 -2428
rect 625 -2436 626 -2434
rect 632 -2430 633 -2428
rect 632 -2436 633 -2434
rect 646 -2430 647 -2428
rect 646 -2436 647 -2434
rect 653 -2430 654 -2428
rect 653 -2436 654 -2434
rect 660 -2430 661 -2428
rect 660 -2436 661 -2434
rect 663 -2436 664 -2434
rect 667 -2430 668 -2428
rect 667 -2436 668 -2434
rect 674 -2430 675 -2428
rect 674 -2436 675 -2434
rect 681 -2430 682 -2428
rect 684 -2430 685 -2428
rect 688 -2430 689 -2428
rect 691 -2430 692 -2428
rect 688 -2436 689 -2434
rect 691 -2436 692 -2434
rect 716 -2430 717 -2428
rect 716 -2436 717 -2434
rect 723 -2430 724 -2428
rect 723 -2436 724 -2434
rect 730 -2430 731 -2428
rect 730 -2436 731 -2434
rect 737 -2430 738 -2428
rect 737 -2436 738 -2434
rect 744 -2430 745 -2428
rect 744 -2436 745 -2434
rect 747 -2436 748 -2434
rect 751 -2430 752 -2428
rect 751 -2436 752 -2434
rect 758 -2430 759 -2428
rect 758 -2436 759 -2434
rect 765 -2430 766 -2428
rect 765 -2436 766 -2434
rect 772 -2430 773 -2428
rect 772 -2436 773 -2434
rect 800 -2430 801 -2428
rect 800 -2436 801 -2434
rect 807 -2430 808 -2428
rect 807 -2436 808 -2434
rect 828 -2430 829 -2428
rect 828 -2436 829 -2434
rect 891 -2430 892 -2428
rect 891 -2436 892 -2434
rect 898 -2430 899 -2428
rect 898 -2436 899 -2434
rect 905 -2430 906 -2428
rect 905 -2436 906 -2434
rect 908 -2436 909 -2434
rect 226 -2471 227 -2469
rect 226 -2477 227 -2475
rect 233 -2471 234 -2469
rect 236 -2471 237 -2469
rect 240 -2471 241 -2469
rect 240 -2477 241 -2475
rect 247 -2477 248 -2475
rect 254 -2471 255 -2469
rect 254 -2477 255 -2475
rect 296 -2471 297 -2469
rect 296 -2477 297 -2475
rect 310 -2471 311 -2469
rect 310 -2477 311 -2475
rect 331 -2471 332 -2469
rect 331 -2477 332 -2475
rect 341 -2471 342 -2469
rect 341 -2477 342 -2475
rect 345 -2471 346 -2469
rect 348 -2471 349 -2469
rect 348 -2477 349 -2475
rect 352 -2471 353 -2469
rect 352 -2477 353 -2475
rect 359 -2471 360 -2469
rect 359 -2477 360 -2475
rect 366 -2471 367 -2469
rect 366 -2477 367 -2475
rect 373 -2471 374 -2469
rect 373 -2477 374 -2475
rect 387 -2471 388 -2469
rect 387 -2477 388 -2475
rect 394 -2471 395 -2469
rect 394 -2477 395 -2475
rect 401 -2471 402 -2469
rect 401 -2477 402 -2475
rect 408 -2471 409 -2469
rect 408 -2477 409 -2475
rect 422 -2471 423 -2469
rect 422 -2477 423 -2475
rect 432 -2471 433 -2469
rect 429 -2477 430 -2475
rect 432 -2477 433 -2475
rect 436 -2471 437 -2469
rect 436 -2477 437 -2475
rect 443 -2471 444 -2469
rect 443 -2477 444 -2475
rect 446 -2477 447 -2475
rect 450 -2471 451 -2469
rect 453 -2471 454 -2469
rect 453 -2477 454 -2475
rect 457 -2471 458 -2469
rect 457 -2477 458 -2475
rect 464 -2471 465 -2469
rect 464 -2477 465 -2475
rect 471 -2471 472 -2469
rect 471 -2477 472 -2475
rect 478 -2471 479 -2469
rect 478 -2477 479 -2475
rect 485 -2471 486 -2469
rect 485 -2477 486 -2475
rect 492 -2471 493 -2469
rect 492 -2477 493 -2475
rect 499 -2471 500 -2469
rect 499 -2477 500 -2475
rect 509 -2471 510 -2469
rect 509 -2477 510 -2475
rect 513 -2471 514 -2469
rect 513 -2477 514 -2475
rect 527 -2471 528 -2469
rect 527 -2477 528 -2475
rect 541 -2471 542 -2469
rect 541 -2477 542 -2475
rect 548 -2471 549 -2469
rect 548 -2477 549 -2475
rect 576 -2471 577 -2469
rect 576 -2477 577 -2475
rect 597 -2471 598 -2469
rect 597 -2477 598 -2475
rect 607 -2471 608 -2469
rect 604 -2477 605 -2475
rect 611 -2471 612 -2469
rect 614 -2471 615 -2469
rect 614 -2477 615 -2475
rect 618 -2471 619 -2469
rect 618 -2477 619 -2475
rect 625 -2471 626 -2469
rect 625 -2477 626 -2475
rect 632 -2471 633 -2469
rect 632 -2477 633 -2475
rect 639 -2471 640 -2469
rect 639 -2477 640 -2475
rect 646 -2471 647 -2469
rect 649 -2471 650 -2469
rect 649 -2477 650 -2475
rect 653 -2471 654 -2469
rect 653 -2477 654 -2475
rect 660 -2471 661 -2469
rect 663 -2471 664 -2469
rect 660 -2477 661 -2475
rect 674 -2471 675 -2469
rect 674 -2477 675 -2475
rect 688 -2471 689 -2469
rect 688 -2477 689 -2475
rect 702 -2471 703 -2469
rect 702 -2477 703 -2475
rect 723 -2471 724 -2469
rect 723 -2477 724 -2475
rect 744 -2471 745 -2469
rect 744 -2477 745 -2475
rect 751 -2471 752 -2469
rect 754 -2471 755 -2469
rect 751 -2477 752 -2475
rect 807 -2471 808 -2469
rect 807 -2477 808 -2475
rect 817 -2471 818 -2469
rect 817 -2477 818 -2475
rect 828 -2471 829 -2469
rect 828 -2477 829 -2475
rect 838 -2471 839 -2469
rect 835 -2477 836 -2475
rect 898 -2471 899 -2469
rect 898 -2477 899 -2475
rect 226 -2492 227 -2490
rect 226 -2498 227 -2496
rect 233 -2498 234 -2496
rect 236 -2498 237 -2496
rect 240 -2492 241 -2490
rect 240 -2498 241 -2496
rect 359 -2492 360 -2490
rect 359 -2498 360 -2496
rect 366 -2492 367 -2490
rect 369 -2492 370 -2490
rect 366 -2498 367 -2496
rect 373 -2492 374 -2490
rect 373 -2498 374 -2496
rect 380 -2492 381 -2490
rect 380 -2498 381 -2496
rect 387 -2492 388 -2490
rect 390 -2492 391 -2490
rect 394 -2492 395 -2490
rect 394 -2498 395 -2496
rect 397 -2498 398 -2496
rect 401 -2492 402 -2490
rect 404 -2492 405 -2490
rect 401 -2498 402 -2496
rect 408 -2492 409 -2490
rect 408 -2498 409 -2496
rect 534 -2492 535 -2490
rect 534 -2498 535 -2496
rect 548 -2492 549 -2490
rect 551 -2492 552 -2490
rect 548 -2498 549 -2496
rect 555 -2492 556 -2490
rect 558 -2498 559 -2496
rect 604 -2492 605 -2490
rect 604 -2498 605 -2496
rect 611 -2492 612 -2490
rect 614 -2492 615 -2490
rect 611 -2498 612 -2496
rect 632 -2492 633 -2490
rect 632 -2498 633 -2496
rect 653 -2492 654 -2490
rect 653 -2498 654 -2496
rect 660 -2492 661 -2490
rect 660 -2498 661 -2496
rect 688 -2492 689 -2490
rect 691 -2492 692 -2490
rect 691 -2498 692 -2496
rect 702 -2492 703 -2490
rect 702 -2498 703 -2496
rect 723 -2492 724 -2490
rect 726 -2492 727 -2490
rect 726 -2498 727 -2496
rect 901 -2492 902 -2490
rect 898 -2498 899 -2496
rect 901 -2498 902 -2496
rect 905 -2492 906 -2490
rect 905 -2498 906 -2496
<< metal1 >>
rect 152 0 206 1
rect 338 0 353 1
rect 366 0 412 1
rect 432 0 514 1
rect 341 -2 360 -1
rect 394 -2 472 -1
rect 492 -2 577 -1
rect 345 -4 377 -3
rect 408 -4 451 -3
rect 464 -4 482 -3
rect 128 -15 150 -14
rect 198 -15 290 -14
rect 292 -15 311 -14
rect 320 -15 458 -14
rect 464 -15 486 -14
rect 502 -15 549 -14
rect 576 -15 626 -14
rect 208 -17 220 -16
rect 243 -17 255 -16
rect 282 -17 342 -16
rect 352 -17 381 -16
rect 415 -17 493 -16
rect 513 -17 542 -16
rect 593 -17 619 -16
rect 296 -19 447 -18
rect 450 -19 472 -18
rect 474 -19 528 -18
rect 303 -21 433 -20
rect 450 -21 479 -20
rect 324 -23 346 -22
rect 352 -23 433 -22
rect 436 -23 479 -22
rect 327 -25 409 -24
rect 429 -25 514 -24
rect 331 -27 367 -26
rect 376 -27 388 -26
rect 401 -27 437 -26
rect 464 -27 535 -26
rect 338 -29 395 -28
rect 401 -29 440 -28
rect 345 -31 405 -30
rect 366 -33 374 -32
rect 394 -33 423 -32
rect 373 -35 507 -34
rect 114 -46 129 -45
rect 142 -46 199 -45
rect 205 -46 220 -45
rect 233 -46 244 -45
rect 247 -46 391 -45
rect 415 -46 430 -45
rect 432 -46 570 -45
rect 593 -46 682 -45
rect 170 -48 241 -47
rect 254 -48 276 -47
rect 317 -48 388 -47
rect 443 -48 556 -47
rect 593 -48 598 -47
rect 618 -48 647 -47
rect 653 -48 692 -47
rect 191 -50 297 -49
rect 331 -50 416 -49
rect 443 -50 493 -49
rect 495 -50 619 -49
rect 625 -50 661 -49
rect 674 -50 689 -49
rect 198 -52 335 -51
rect 338 -52 374 -51
rect 394 -52 493 -51
rect 502 -52 584 -51
rect 212 -54 304 -53
rect 338 -54 381 -53
rect 478 -54 640 -53
rect 219 -56 311 -55
rect 369 -56 521 -55
rect 527 -56 531 -55
rect 534 -56 668 -55
rect 240 -58 325 -57
rect 380 -58 577 -57
rect 254 -60 451 -59
rect 478 -60 626 -59
rect 177 -62 451 -61
rect 485 -62 563 -61
rect 261 -64 367 -63
rect 408 -64 486 -63
rect 499 -64 535 -63
rect 548 -64 633 -63
rect 226 -66 367 -65
rect 387 -66 549 -65
rect 268 -68 321 -67
rect 408 -68 458 -67
rect 506 -68 605 -67
rect 282 -70 311 -69
rect 436 -70 458 -69
rect 474 -70 507 -69
rect 513 -70 612 -69
rect 282 -72 346 -71
rect 422 -72 437 -71
rect 446 -72 500 -71
rect 527 -72 591 -71
rect 163 -74 346 -73
rect 422 -74 472 -73
rect 530 -74 591 -73
rect 289 -76 325 -75
rect 464 -76 514 -75
rect 289 -78 402 -77
rect 296 -80 398 -79
rect 184 -82 398 -81
rect 303 -84 353 -83
rect 373 -84 402 -83
rect 348 -86 465 -85
rect 352 -88 482 -87
rect 51 -99 412 -98
rect 464 -99 724 -98
rect 58 -101 454 -100
rect 471 -101 815 -100
rect 65 -103 143 -102
rect 145 -103 185 -102
rect 198 -103 209 -102
rect 275 -103 377 -102
rect 394 -103 773 -102
rect 72 -105 83 -104
rect 86 -105 118 -104
rect 121 -105 195 -104
rect 198 -105 269 -104
rect 275 -105 475 -104
rect 485 -105 808 -104
rect 93 -107 297 -106
rect 331 -107 384 -106
rect 485 -107 612 -106
rect 632 -107 780 -106
rect 107 -109 248 -108
rect 268 -109 339 -108
rect 345 -109 430 -108
rect 492 -109 696 -108
rect 114 -111 136 -110
rect 156 -111 290 -110
rect 359 -111 395 -110
rect 418 -111 612 -110
rect 639 -111 787 -110
rect 114 -113 279 -112
rect 324 -113 360 -112
rect 366 -113 388 -112
rect 450 -113 640 -112
rect 653 -113 738 -112
rect 128 -115 255 -114
rect 261 -115 290 -114
rect 310 -115 325 -114
rect 369 -115 430 -114
rect 495 -115 710 -114
rect 152 -117 262 -116
rect 303 -117 311 -116
rect 387 -117 402 -116
rect 520 -117 654 -116
rect 660 -117 717 -116
rect 170 -119 297 -118
rect 303 -119 465 -118
rect 478 -119 661 -118
rect 667 -119 752 -118
rect 170 -121 227 -120
rect 247 -121 381 -120
rect 534 -121 766 -120
rect 100 -123 227 -122
rect 254 -123 472 -122
rect 534 -123 580 -122
rect 583 -123 633 -122
rect 646 -123 668 -122
rect 674 -123 731 -122
rect 184 -125 188 -124
rect 201 -125 332 -124
rect 380 -125 475 -124
rect 499 -125 647 -124
rect 681 -125 822 -124
rect 219 -127 339 -126
rect 436 -127 500 -126
rect 513 -127 682 -126
rect 688 -127 794 -126
rect 191 -129 437 -128
rect 467 -129 584 -128
rect 590 -129 619 -128
rect 625 -129 689 -128
rect 219 -131 241 -130
rect 317 -131 402 -130
rect 453 -131 619 -130
rect 205 -133 241 -132
rect 282 -133 318 -132
rect 481 -133 514 -132
rect 527 -133 675 -132
rect 177 -135 283 -134
rect 506 -135 528 -134
rect 548 -135 745 -134
rect 177 -137 213 -136
rect 373 -137 549 -136
rect 562 -137 801 -136
rect 163 -139 213 -138
rect 334 -139 563 -138
rect 569 -139 759 -138
rect 163 -141 353 -140
rect 373 -141 598 -140
rect 205 -143 234 -142
rect 352 -143 626 -142
rect 208 -145 234 -144
rect 415 -145 507 -144
rect 541 -145 570 -144
rect 576 -145 703 -144
rect 345 -147 416 -146
rect 422 -147 542 -146
rect 555 -147 598 -146
rect 422 -149 458 -148
rect 520 -149 577 -148
rect 443 -151 556 -150
rect 408 -153 444 -152
rect 457 -153 605 -152
rect 593 -155 605 -154
rect 44 -166 185 -165
rect 191 -166 213 -165
rect 268 -166 353 -165
rect 362 -166 766 -165
rect 793 -166 850 -165
rect 65 -168 167 -167
rect 184 -168 311 -167
rect 348 -168 696 -167
rect 751 -168 794 -167
rect 800 -168 864 -167
rect 65 -170 73 -169
rect 79 -170 87 -169
rect 100 -170 258 -169
rect 310 -170 325 -169
rect 352 -170 454 -169
rect 464 -170 808 -169
rect 814 -170 836 -169
rect 72 -172 360 -171
rect 408 -172 787 -171
rect 821 -172 843 -171
rect 86 -174 195 -173
rect 198 -174 234 -173
rect 324 -174 423 -173
rect 471 -174 808 -173
rect 103 -176 356 -175
rect 411 -176 724 -175
rect 730 -176 787 -175
rect 117 -178 766 -177
rect 772 -178 815 -177
rect 121 -180 202 -179
rect 212 -180 276 -179
rect 285 -180 423 -179
rect 492 -180 549 -179
rect 576 -180 829 -179
rect 121 -182 125 -181
rect 128 -182 465 -181
rect 495 -182 745 -181
rect 779 -182 822 -181
rect 128 -184 227 -183
rect 275 -184 318 -183
rect 415 -184 759 -183
rect 138 -186 426 -185
rect 460 -186 759 -185
rect 145 -188 367 -187
rect 415 -188 479 -187
rect 495 -188 738 -187
rect 163 -190 409 -189
rect 443 -190 479 -189
rect 499 -190 577 -189
rect 632 -190 801 -189
rect 58 -192 164 -191
rect 177 -192 234 -191
rect 296 -192 318 -191
rect 359 -192 738 -191
rect 51 -194 59 -193
rect 177 -194 248 -193
rect 282 -194 297 -193
rect 366 -194 402 -193
rect 443 -194 482 -193
rect 520 -194 524 -193
rect 548 -194 563 -193
rect 660 -194 724 -193
rect 730 -194 860 -193
rect 51 -196 388 -195
rect 450 -196 633 -195
rect 667 -196 696 -195
rect 709 -196 752 -195
rect 191 -198 220 -197
rect 247 -198 381 -197
rect 429 -198 451 -197
rect 457 -198 500 -197
rect 520 -198 535 -197
rect 618 -198 661 -197
rect 681 -198 780 -197
rect 205 -200 220 -199
rect 226 -200 458 -199
rect 474 -200 668 -199
rect 688 -200 745 -199
rect 205 -202 255 -201
rect 303 -202 381 -201
rect 394 -202 430 -201
rect 439 -202 619 -201
rect 646 -202 689 -201
rect 702 -202 710 -201
rect 716 -202 773 -201
rect 156 -204 395 -203
rect 474 -204 542 -203
rect 653 -204 682 -203
rect 114 -206 157 -205
rect 254 -206 269 -205
rect 289 -206 304 -205
rect 331 -206 402 -205
rect 404 -206 542 -205
rect 639 -206 654 -205
rect 674 -206 703 -205
rect 289 -208 647 -207
rect 331 -210 437 -209
rect 492 -210 717 -209
rect 338 -212 437 -211
rect 523 -212 535 -211
rect 569 -212 640 -211
rect 261 -214 339 -213
rect 373 -214 388 -213
rect 527 -214 563 -213
rect 611 -214 675 -213
rect 261 -216 346 -215
rect 506 -216 528 -215
rect 555 -216 570 -215
rect 583 -216 612 -215
rect 107 -218 584 -217
rect 107 -220 283 -219
rect 345 -220 626 -219
rect 142 -222 507 -221
rect 597 -222 626 -221
rect 142 -224 377 -223
rect 597 -224 605 -223
rect 149 -226 556 -225
rect 590 -226 605 -225
rect 149 -228 171 -227
rect 513 -228 591 -227
rect 135 -230 171 -229
rect 485 -230 514 -229
rect 93 -232 486 -231
rect 93 -234 153 -233
rect 135 -236 293 -235
rect 2 -247 69 -246
rect 72 -247 349 -246
rect 352 -247 780 -246
rect 807 -247 906 -246
rect 9 -249 286 -248
rect 289 -249 311 -248
rect 352 -249 535 -248
rect 569 -249 941 -248
rect 16 -251 360 -250
rect 383 -251 675 -250
rect 681 -251 892 -250
rect 23 -253 59 -252
rect 72 -253 269 -252
rect 289 -253 451 -252
rect 471 -253 857 -252
rect 30 -255 454 -254
rect 492 -255 612 -254
rect 730 -255 885 -254
rect 37 -257 66 -256
rect 86 -257 293 -256
rect 303 -257 311 -256
rect 359 -257 496 -256
rect 520 -257 524 -256
rect 548 -257 612 -256
rect 667 -257 731 -256
rect 744 -257 780 -256
rect 814 -257 955 -256
rect 51 -259 255 -258
rect 268 -259 339 -258
rect 401 -259 591 -258
rect 597 -259 682 -258
rect 758 -259 871 -258
rect 51 -261 395 -260
rect 418 -261 808 -260
rect 821 -261 920 -260
rect 58 -263 500 -262
rect 506 -263 745 -262
rect 758 -263 801 -262
rect 828 -263 927 -262
rect 65 -265 913 -264
rect 79 -267 87 -266
rect 93 -267 283 -266
rect 303 -267 307 -266
rect 376 -267 500 -266
rect 520 -267 528 -266
rect 555 -267 675 -266
rect 751 -267 801 -266
rect 835 -267 934 -266
rect 79 -269 444 -268
rect 464 -269 507 -268
rect 541 -269 556 -268
rect 569 -269 598 -268
rect 653 -269 668 -268
rect 723 -269 752 -268
rect 765 -269 829 -268
rect 842 -269 948 -268
rect 93 -271 101 -270
rect 103 -271 591 -270
rect 632 -271 654 -270
rect 709 -271 724 -270
rect 793 -271 815 -270
rect 849 -271 878 -270
rect 100 -273 416 -272
rect 425 -273 864 -272
rect 121 -275 164 -274
rect 170 -275 283 -274
rect 338 -275 377 -274
rect 387 -275 444 -274
rect 450 -275 843 -274
rect 121 -277 367 -276
rect 394 -277 689 -276
rect 702 -277 864 -276
rect 142 -279 258 -278
rect 366 -279 549 -278
rect 576 -279 580 -278
rect 583 -279 633 -278
rect 646 -279 703 -278
rect 772 -279 850 -278
rect 142 -281 468 -280
rect 474 -281 542 -280
rect 576 -281 605 -280
rect 625 -281 647 -280
rect 660 -281 710 -280
rect 716 -281 773 -280
rect 786 -281 794 -280
rect 156 -283 388 -282
rect 397 -283 822 -282
rect 156 -285 276 -284
rect 425 -285 535 -284
rect 551 -285 717 -284
rect 737 -285 787 -284
rect 163 -287 262 -286
rect 275 -287 346 -286
rect 436 -287 836 -286
rect 44 -289 437 -288
rect 439 -289 766 -288
rect 170 -291 332 -290
rect 457 -291 584 -290
rect 639 -291 661 -290
rect 688 -291 899 -290
rect 128 -293 332 -292
rect 457 -293 640 -292
rect 695 -293 738 -292
rect 184 -295 363 -294
rect 478 -295 493 -294
rect 579 -295 605 -294
rect 618 -295 696 -294
rect 166 -297 619 -296
rect 184 -299 192 -298
rect 205 -299 405 -298
rect 478 -299 486 -298
rect 488 -299 626 -298
rect 107 -301 192 -300
rect 205 -301 220 -300
rect 254 -301 475 -300
rect 485 -301 563 -300
rect 107 -303 125 -302
rect 219 -303 234 -302
rect 261 -303 423 -302
rect 446 -303 563 -302
rect 198 -305 234 -304
rect 247 -305 423 -304
rect 114 -307 248 -306
rect 317 -307 346 -306
rect 114 -309 430 -308
rect 198 -311 297 -310
rect 380 -311 430 -310
rect 44 -313 381 -312
rect 135 -315 297 -314
rect 135 -317 213 -316
rect 226 -317 318 -316
rect 212 -319 325 -318
rect 226 -321 409 -320
rect 117 -323 409 -322
rect 324 -325 356 -324
rect 16 -336 416 -335
rect 436 -336 682 -335
rect 905 -336 962 -335
rect 16 -338 108 -337
rect 124 -338 283 -337
rect 289 -338 398 -337
rect 401 -338 696 -337
rect 758 -338 906 -337
rect 912 -338 1025 -337
rect 44 -340 76 -339
rect 79 -340 416 -339
rect 439 -340 573 -339
rect 618 -340 1004 -339
rect 37 -342 80 -341
rect 96 -342 682 -341
rect 730 -342 759 -341
rect 779 -342 913 -341
rect 919 -342 983 -341
rect 2 -344 38 -343
rect 44 -344 94 -343
rect 100 -344 283 -343
rect 296 -344 304 -343
rect 310 -344 461 -343
rect 467 -344 885 -343
rect 926 -344 990 -343
rect 2 -346 346 -345
rect 355 -346 437 -345
rect 443 -346 997 -345
rect 51 -348 461 -347
rect 467 -348 899 -347
rect 933 -348 976 -347
rect 51 -350 489 -349
rect 548 -350 969 -349
rect 65 -352 164 -351
rect 191 -352 311 -351
rect 331 -352 402 -351
rect 411 -352 941 -351
rect 93 -354 199 -353
rect 212 -354 454 -353
rect 457 -354 955 -353
rect 100 -356 143 -355
rect 149 -356 164 -355
rect 198 -356 234 -355
rect 243 -356 290 -355
rect 296 -356 531 -355
rect 583 -356 619 -355
rect 621 -356 780 -355
rect 793 -356 934 -355
rect 107 -358 132 -357
rect 142 -358 220 -357
rect 226 -358 419 -357
rect 422 -358 885 -357
rect 72 -360 227 -359
rect 233 -360 377 -359
rect 380 -360 552 -359
rect 667 -360 696 -359
rect 751 -360 794 -359
rect 800 -360 920 -359
rect 114 -362 398 -361
rect 446 -362 633 -361
rect 744 -362 801 -361
rect 842 -362 899 -361
rect 86 -364 115 -363
rect 177 -364 220 -363
rect 254 -364 384 -363
rect 387 -364 423 -363
rect 457 -364 577 -363
rect 597 -364 668 -363
rect 702 -364 745 -363
rect 786 -364 843 -363
rect 849 -364 927 -363
rect 177 -366 185 -365
rect 194 -366 703 -365
rect 737 -366 787 -365
rect 814 -366 850 -365
rect 856 -366 941 -365
rect 128 -368 185 -367
rect 254 -368 276 -367
rect 338 -368 444 -367
rect 464 -368 857 -367
rect 877 -368 955 -367
rect 128 -370 136 -369
rect 156 -370 339 -369
rect 352 -370 598 -369
rect 632 -370 640 -369
rect 660 -370 738 -369
rect 835 -370 878 -369
rect 86 -372 136 -371
rect 156 -372 318 -371
rect 359 -372 475 -371
rect 485 -372 731 -371
rect 772 -372 836 -371
rect 170 -374 353 -373
rect 373 -374 871 -373
rect 82 -376 171 -375
rect 212 -376 360 -375
rect 387 -376 430 -375
rect 464 -376 486 -375
rect 516 -376 640 -375
rect 646 -376 661 -375
rect 709 -376 871 -375
rect 261 -378 346 -377
rect 425 -378 577 -377
rect 653 -378 710 -377
rect 723 -378 815 -377
rect 247 -380 262 -379
rect 268 -380 374 -379
rect 429 -380 451 -379
rect 471 -380 864 -379
rect 72 -382 472 -381
rect 541 -382 584 -381
rect 625 -382 654 -381
rect 674 -382 724 -381
rect 821 -382 864 -381
rect 121 -384 269 -383
rect 275 -384 395 -383
rect 506 -384 542 -383
rect 551 -384 773 -383
rect 23 -386 122 -385
rect 240 -386 248 -385
rect 306 -386 647 -385
rect 765 -386 822 -385
rect 23 -388 31 -387
rect 58 -388 507 -387
rect 520 -388 626 -387
rect 716 -388 766 -387
rect 30 -390 69 -389
rect 149 -390 241 -389
rect 317 -390 367 -389
rect 394 -390 808 -389
rect 58 -392 325 -391
rect 362 -392 675 -391
rect 688 -392 717 -391
rect 68 -394 332 -393
rect 366 -394 433 -393
rect 513 -394 521 -393
rect 562 -394 689 -393
rect 324 -396 556 -395
rect 569 -396 752 -395
rect 499 -398 563 -397
rect 569 -398 612 -397
rect 478 -400 500 -399
rect 513 -400 892 -399
rect 478 -402 493 -401
rect 527 -402 556 -401
rect 590 -402 612 -401
rect 828 -402 892 -401
rect 9 -404 528 -403
rect 534 -404 591 -403
rect 604 -404 808 -403
rect 9 -406 90 -405
rect 159 -406 829 -405
rect 404 -408 605 -407
rect 408 -410 535 -409
rect 408 -412 493 -411
rect 9 -423 132 -422
rect 142 -423 244 -422
rect 275 -423 353 -422
rect 362 -423 626 -422
rect 814 -423 1074 -422
rect 9 -425 640 -424
rect 849 -425 1046 -424
rect 16 -427 94 -426
rect 156 -427 283 -426
rect 324 -427 412 -426
rect 415 -427 815 -426
rect 912 -427 1032 -426
rect 16 -429 654 -428
rect 765 -429 850 -428
rect 926 -429 1053 -428
rect 23 -431 153 -430
rect 191 -431 423 -430
rect 429 -431 808 -430
rect 828 -431 927 -430
rect 933 -431 1011 -430
rect 1024 -431 1088 -430
rect 23 -433 391 -432
rect 394 -433 808 -432
rect 828 -433 892 -432
rect 940 -433 1039 -432
rect 30 -435 185 -434
rect 226 -435 328 -434
rect 373 -435 482 -434
rect 513 -435 535 -434
rect 548 -435 920 -434
rect 940 -435 1004 -434
rect 30 -437 59 -436
rect 65 -437 360 -436
rect 397 -437 668 -436
rect 670 -437 1004 -436
rect 37 -439 73 -438
rect 86 -439 101 -438
rect 163 -439 192 -438
rect 219 -439 227 -438
rect 275 -439 398 -438
rect 401 -439 416 -438
rect 432 -439 717 -438
rect 730 -439 1025 -438
rect 37 -441 94 -440
rect 100 -441 108 -440
rect 184 -441 318 -440
rect 324 -441 423 -440
rect 450 -441 454 -440
rect 467 -441 479 -440
rect 523 -441 1102 -440
rect 44 -443 80 -442
rect 187 -443 220 -442
rect 296 -443 430 -442
rect 450 -443 724 -442
rect 730 -443 752 -442
rect 786 -443 892 -442
rect 954 -443 1060 -442
rect 44 -445 251 -444
rect 310 -445 318 -444
rect 331 -445 374 -444
rect 401 -445 412 -444
rect 478 -445 906 -444
rect 961 -445 1095 -444
rect 51 -447 241 -446
rect 247 -447 297 -446
rect 331 -447 367 -446
rect 460 -447 962 -446
rect 968 -447 1109 -446
rect 51 -449 486 -448
rect 530 -449 871 -448
rect 975 -449 1081 -448
rect 58 -451 552 -450
rect 562 -451 640 -450
rect 649 -451 766 -450
rect 772 -451 871 -450
rect 884 -451 976 -450
rect 982 -451 1116 -450
rect 65 -453 388 -452
rect 408 -453 563 -452
rect 576 -453 626 -452
rect 674 -453 906 -452
rect 989 -453 1123 -452
rect 68 -455 717 -454
rect 737 -455 990 -454
rect 996 -455 1067 -454
rect 72 -457 668 -456
rect 709 -457 787 -456
rect 800 -457 913 -456
rect 75 -459 108 -458
rect 121 -459 885 -458
rect 79 -461 171 -460
rect 205 -461 248 -460
rect 261 -461 367 -460
rect 387 -461 1018 -460
rect 82 -463 773 -462
rect 779 -463 955 -462
rect 121 -465 178 -464
rect 233 -465 409 -464
rect 485 -465 577 -464
rect 597 -465 654 -464
rect 702 -465 710 -464
rect 744 -465 801 -464
rect 821 -465 920 -464
rect 128 -467 171 -466
rect 177 -467 381 -466
rect 520 -467 598 -466
rect 604 -467 675 -466
rect 681 -467 745 -466
rect 835 -467 934 -466
rect 96 -469 129 -468
rect 135 -469 311 -468
rect 338 -469 360 -468
rect 464 -469 836 -468
rect 856 -469 983 -468
rect 96 -471 164 -470
rect 212 -471 381 -470
rect 464 -471 528 -470
rect 534 -471 580 -470
rect 607 -471 703 -470
rect 793 -471 857 -470
rect 863 -471 969 -470
rect 156 -473 339 -472
rect 471 -473 528 -472
rect 548 -473 752 -472
rect 758 -473 864 -472
rect 877 -473 997 -472
rect 149 -475 472 -474
rect 509 -475 794 -474
rect 212 -477 304 -476
rect 516 -477 878 -476
rect 2 -479 304 -478
rect 520 -479 689 -478
rect 2 -481 139 -480
rect 233 -481 255 -480
rect 261 -481 269 -480
rect 572 -481 759 -480
rect 124 -483 269 -482
rect 604 -483 689 -482
rect 240 -485 290 -484
rect 611 -485 780 -484
rect 254 -487 444 -486
rect 618 -487 724 -486
rect 205 -489 444 -488
rect 569 -489 619 -488
rect 621 -489 948 -488
rect 289 -491 500 -490
rect 569 -491 899 -490
rect 345 -493 612 -492
rect 632 -493 738 -492
rect 842 -493 948 -492
rect 159 -495 346 -494
rect 436 -495 500 -494
rect 583 -495 843 -494
rect 394 -497 437 -496
rect 446 -497 633 -496
rect 646 -497 822 -496
rect 457 -499 899 -498
rect 457 -501 542 -500
rect 583 -501 591 -500
rect 660 -501 682 -500
rect 492 -503 542 -502
rect 565 -503 661 -502
rect 453 -505 493 -504
rect 506 -505 591 -504
rect 282 -507 507 -506
rect 2 -518 143 -517
rect 149 -518 384 -517
rect 390 -518 409 -517
rect 411 -518 822 -517
rect 2 -520 405 -519
rect 425 -520 479 -519
rect 509 -520 1116 -519
rect 9 -522 139 -521
rect 159 -522 451 -521
rect 544 -522 1109 -521
rect 9 -524 787 -523
rect 821 -524 850 -523
rect 16 -526 94 -525
rect 107 -526 129 -525
rect 177 -526 479 -525
rect 572 -526 990 -525
rect 58 -528 563 -527
rect 576 -528 843 -527
rect 989 -528 1018 -527
rect 72 -530 157 -529
rect 177 -530 188 -529
rect 212 -530 563 -529
rect 579 -530 1123 -529
rect 75 -532 381 -531
rect 429 -532 622 -531
rect 628 -532 1074 -531
rect 79 -534 388 -533
rect 415 -534 430 -533
rect 443 -534 465 -533
rect 555 -534 577 -533
rect 646 -534 1032 -533
rect 58 -536 80 -535
rect 86 -536 94 -535
rect 128 -536 304 -535
rect 317 -536 451 -535
rect 464 -536 780 -535
rect 786 -536 948 -535
rect 1017 -536 1039 -535
rect 86 -538 132 -537
rect 145 -538 213 -537
rect 240 -538 325 -537
rect 387 -538 591 -537
rect 667 -538 1095 -537
rect 51 -540 591 -539
rect 674 -540 850 -539
rect 947 -540 997 -539
rect 1031 -540 1046 -539
rect 51 -542 598 -541
rect 674 -542 731 -541
rect 754 -542 1102 -541
rect 121 -544 304 -543
rect 446 -544 815 -543
rect 828 -544 1074 -543
rect 72 -546 122 -545
rect 135 -546 241 -545
rect 247 -546 297 -545
rect 481 -546 668 -545
rect 695 -546 699 -545
rect 730 -546 773 -545
rect 807 -546 1046 -545
rect 135 -548 206 -547
rect 247 -548 416 -547
rect 520 -548 647 -547
rect 695 -548 703 -547
rect 772 -548 885 -547
rect 996 -548 1025 -547
rect 1038 -548 1060 -547
rect 145 -550 227 -549
rect 250 -550 318 -549
rect 471 -550 521 -549
rect 551 -550 885 -549
rect 1059 -550 1067 -549
rect 37 -552 227 -551
rect 261 -552 507 -551
rect 555 -552 570 -551
rect 597 -552 640 -551
rect 698 -552 703 -551
rect 723 -552 1025 -551
rect 44 -554 570 -553
rect 632 -554 808 -553
rect 814 -554 892 -553
rect 940 -554 1067 -553
rect 44 -556 423 -555
rect 436 -556 472 -555
rect 492 -556 507 -555
rect 583 -556 633 -555
rect 639 -556 654 -555
rect 723 -556 801 -555
rect 828 -556 857 -555
rect 940 -556 969 -555
rect 156 -558 192 -557
rect 205 -558 276 -557
rect 289 -558 381 -557
rect 422 -558 780 -557
rect 800 -558 864 -557
rect 114 -560 290 -559
rect 296 -560 402 -559
rect 492 -560 500 -559
rect 583 -560 608 -559
rect 653 -560 661 -559
rect 835 -560 969 -559
rect 100 -562 115 -561
rect 152 -562 276 -561
rect 338 -562 437 -561
rect 499 -562 528 -561
rect 604 -562 892 -561
rect 30 -564 339 -563
rect 401 -564 612 -563
rect 660 -564 689 -563
rect 835 -564 871 -563
rect 30 -566 486 -565
rect 513 -566 528 -565
rect 604 -566 626 -565
rect 842 -566 878 -565
rect 16 -568 626 -567
rect 856 -568 955 -567
rect 100 -570 220 -569
rect 261 -570 279 -569
rect 352 -570 486 -569
rect 513 -570 542 -569
rect 863 -570 899 -569
rect 954 -570 1004 -569
rect 37 -572 220 -571
rect 254 -572 353 -571
rect 394 -572 689 -571
rect 870 -572 906 -571
rect 975 -572 1004 -571
rect 191 -574 234 -573
rect 254 -574 283 -573
rect 394 -574 535 -573
rect 541 -574 717 -573
rect 877 -574 913 -573
rect 975 -574 1011 -573
rect 233 -576 671 -575
rect 716 -576 738 -575
rect 898 -576 920 -575
rect 1010 -576 1081 -575
rect 107 -578 1081 -577
rect 282 -580 367 -579
rect 457 -580 535 -579
rect 565 -580 913 -579
rect 919 -580 927 -579
rect 65 -582 367 -581
rect 457 -582 983 -581
rect 65 -584 311 -583
rect 523 -584 612 -583
rect 709 -584 738 -583
rect 751 -584 983 -583
rect 170 -586 311 -585
rect 373 -586 524 -585
rect 565 -586 906 -585
rect 170 -588 199 -587
rect 345 -588 374 -587
rect 681 -588 710 -587
rect 751 -588 766 -587
rect 198 -590 461 -589
rect 618 -590 766 -589
rect 345 -592 360 -591
rect 453 -592 682 -591
rect 758 -592 927 -591
rect 184 -594 360 -593
rect 618 -594 1053 -593
rect 23 -596 185 -595
rect 744 -596 759 -595
rect 933 -596 1053 -595
rect 23 -598 164 -597
rect 744 -598 794 -597
rect 933 -598 962 -597
rect 163 -600 549 -599
rect 334 -602 794 -601
rect 467 -604 962 -603
rect 548 -606 650 -605
rect 23 -617 381 -616
rect 415 -617 437 -616
rect 453 -617 766 -616
rect 905 -617 1214 -616
rect 1216 -617 1361 -616
rect 40 -619 587 -618
rect 618 -619 675 -618
rect 716 -619 766 -618
rect 814 -619 906 -618
rect 961 -619 1158 -618
rect 2 -621 675 -620
rect 702 -621 717 -620
rect 723 -621 815 -620
rect 961 -621 983 -620
rect 989 -621 1102 -620
rect 2 -623 941 -622
rect 975 -623 1095 -622
rect 44 -625 619 -624
rect 621 -625 983 -624
rect 996 -625 1109 -624
rect 44 -627 339 -626
rect 380 -627 612 -626
rect 635 -627 1053 -626
rect 1059 -627 1193 -626
rect 47 -629 206 -628
rect 229 -629 304 -628
rect 324 -629 339 -628
rect 387 -629 724 -628
rect 726 -629 857 -628
rect 884 -629 976 -628
rect 1010 -629 1186 -628
rect 51 -631 433 -630
rect 460 -631 626 -630
rect 649 -631 1172 -630
rect 58 -633 787 -632
rect 821 -633 857 -632
rect 870 -633 885 -632
rect 891 -633 990 -632
rect 1031 -633 1130 -632
rect 51 -635 59 -634
rect 65 -635 549 -634
rect 551 -635 850 -634
rect 898 -635 1011 -634
rect 1038 -635 1123 -634
rect 65 -637 108 -636
rect 121 -637 325 -636
rect 331 -637 346 -636
rect 404 -637 1053 -636
rect 1066 -637 1200 -636
rect 16 -639 108 -638
rect 121 -639 657 -638
rect 667 -639 703 -638
rect 730 -639 997 -638
rect 1045 -639 1081 -638
rect 1083 -639 1088 -638
rect 16 -641 188 -640
rect 226 -641 388 -640
rect 418 -641 426 -640
rect 464 -641 1165 -640
rect 75 -643 1004 -642
rect 86 -645 206 -644
rect 247 -645 346 -644
rect 422 -645 444 -644
rect 464 -645 514 -644
rect 523 -645 1025 -644
rect 37 -647 87 -646
rect 89 -647 1179 -646
rect 100 -649 468 -648
rect 492 -649 514 -648
rect 541 -649 787 -648
rect 800 -649 871 -648
rect 912 -649 1004 -648
rect 100 -651 391 -650
rect 408 -651 423 -650
rect 478 -651 542 -650
rect 544 -651 752 -650
rect 779 -651 941 -650
rect 947 -651 1067 -650
rect 128 -653 276 -652
rect 289 -653 409 -652
rect 492 -653 661 -652
rect 709 -653 752 -652
rect 807 -653 850 -652
rect 912 -653 927 -652
rect 947 -653 1018 -652
rect 93 -655 129 -654
rect 142 -655 1144 -654
rect 61 -657 143 -656
rect 240 -657 444 -656
rect 502 -657 1039 -656
rect 9 -659 62 -658
rect 93 -659 199 -658
rect 247 -659 283 -658
rect 289 -659 367 -658
rect 394 -659 479 -658
rect 520 -659 801 -658
rect 810 -659 1088 -658
rect 9 -661 370 -660
rect 418 -661 521 -660
rect 548 -661 570 -660
rect 590 -661 612 -660
rect 632 -661 661 -660
rect 709 -661 745 -660
rect 821 -661 920 -660
rect 933 -661 1018 -660
rect 23 -663 367 -662
rect 534 -663 570 -662
rect 576 -663 591 -662
rect 597 -663 626 -662
rect 632 -663 1116 -662
rect 110 -665 395 -664
rect 534 -665 556 -664
rect 558 -665 1032 -664
rect 145 -667 241 -666
rect 261 -667 283 -666
rect 296 -667 437 -666
rect 555 -667 577 -666
rect 597 -667 731 -666
rect 733 -667 1046 -666
rect 198 -669 237 -668
rect 254 -669 262 -668
rect 275 -669 405 -668
rect 562 -669 1074 -668
rect 278 -671 297 -670
rect 303 -671 311 -670
rect 317 -671 332 -670
rect 334 -671 892 -670
rect 954 -671 1060 -670
rect 163 -673 318 -672
rect 457 -673 1074 -672
rect 163 -675 213 -674
rect 268 -675 458 -674
rect 562 -675 759 -674
rect 772 -675 920 -674
rect 968 -675 1025 -674
rect 191 -677 213 -676
rect 219 -677 269 -676
rect 310 -677 486 -676
rect 565 -677 1137 -676
rect 177 -679 192 -678
rect 383 -679 969 -678
rect 177 -681 500 -680
rect 565 -681 1151 -680
rect 149 -683 500 -682
rect 583 -683 773 -682
rect 842 -683 899 -682
rect 149 -685 157 -684
rect 184 -685 220 -684
rect 485 -685 528 -684
rect 583 -685 1207 -684
rect 156 -687 430 -686
rect 506 -687 528 -686
rect 586 -687 759 -686
rect 863 -687 927 -686
rect 72 -689 507 -688
rect 628 -689 843 -688
rect 877 -689 955 -688
rect 72 -691 80 -690
rect 170 -691 185 -690
rect 429 -691 668 -690
rect 695 -691 745 -690
rect 828 -691 864 -690
rect 68 -693 80 -692
rect 114 -693 171 -692
rect 646 -693 934 -692
rect 114 -695 374 -694
rect 681 -695 696 -694
rect 737 -695 780 -694
rect 835 -695 878 -694
rect 373 -697 472 -696
rect 688 -697 829 -696
rect 233 -699 472 -698
rect 653 -699 689 -698
rect 793 -699 836 -698
rect 233 -701 360 -700
rect 383 -701 738 -700
rect 226 -703 360 -702
rect 446 -703 682 -702
rect 254 -705 654 -704
rect 639 -707 794 -706
rect 135 -709 640 -708
rect 135 -711 605 -710
rect 450 -713 605 -712
rect 450 -715 647 -714
rect 2 -726 108 -725
rect 131 -726 311 -725
rect 338 -726 447 -725
rect 464 -726 556 -725
rect 569 -726 573 -725
rect 586 -726 934 -725
rect 1136 -726 1221 -725
rect 1360 -726 1417 -725
rect 2 -728 80 -727
rect 89 -728 195 -727
rect 198 -728 202 -727
rect 254 -728 734 -727
rect 828 -728 1263 -727
rect 9 -730 724 -729
rect 726 -730 1088 -729
rect 1143 -730 1228 -729
rect 9 -732 52 -731
rect 79 -732 241 -731
rect 254 -732 374 -731
rect 390 -732 1207 -731
rect 16 -734 62 -733
rect 89 -734 696 -733
rect 705 -734 1200 -733
rect 16 -736 370 -735
rect 401 -736 990 -735
rect 1017 -736 1088 -735
rect 1164 -736 1242 -735
rect 30 -738 111 -737
rect 156 -738 241 -737
rect 338 -738 409 -737
rect 422 -738 465 -737
rect 485 -738 566 -737
rect 611 -738 633 -737
rect 635 -738 1151 -737
rect 1178 -738 1249 -737
rect 37 -740 381 -739
rect 390 -740 423 -739
rect 436 -740 486 -739
rect 495 -740 535 -739
rect 576 -740 612 -739
rect 646 -740 745 -739
rect 828 -740 1207 -739
rect 37 -742 94 -741
rect 100 -742 559 -741
rect 576 -742 626 -741
rect 649 -742 822 -741
rect 905 -742 934 -741
rect 975 -742 990 -741
rect 1017 -742 1046 -741
rect 1080 -742 1200 -741
rect 51 -744 1214 -743
rect 65 -746 94 -745
rect 100 -746 129 -745
rect 142 -746 157 -745
rect 163 -746 367 -745
rect 380 -746 416 -745
rect 443 -746 1235 -745
rect 65 -748 234 -747
rect 289 -748 444 -747
rect 457 -748 633 -747
rect 649 -748 1172 -747
rect 1185 -748 1256 -747
rect 86 -750 1081 -749
rect 1094 -750 1151 -749
rect 1157 -750 1186 -749
rect 107 -752 150 -751
rect 170 -752 174 -751
rect 177 -752 535 -751
rect 590 -752 976 -751
rect 1101 -752 1179 -751
rect 142 -754 388 -753
rect 408 -754 479 -753
rect 502 -754 997 -753
rect 1108 -754 1172 -753
rect 149 -756 514 -755
rect 516 -756 696 -755
rect 709 -756 745 -755
rect 856 -756 906 -755
rect 912 -756 1046 -755
rect 1115 -756 1165 -755
rect 170 -758 206 -757
rect 212 -758 234 -757
rect 299 -758 822 -757
rect 856 -758 969 -757
rect 1059 -758 1116 -757
rect 1122 -758 1214 -757
rect 44 -760 969 -759
rect 44 -762 384 -761
rect 415 -762 682 -761
rect 709 -762 717 -761
rect 723 -762 752 -761
rect 765 -762 913 -761
rect 961 -762 1095 -761
rect 33 -764 752 -763
rect 765 -764 1053 -763
rect 114 -766 682 -765
rect 702 -766 717 -765
rect 730 -766 1011 -765
rect 114 -768 500 -767
rect 506 -768 626 -767
rect 639 -768 1158 -767
rect 128 -770 1060 -769
rect 135 -772 640 -771
rect 653 -772 1144 -771
rect 75 -774 136 -773
rect 191 -774 213 -773
rect 352 -774 405 -773
rect 457 -774 507 -773
rect 513 -774 1193 -773
rect 121 -776 192 -775
rect 198 -776 220 -775
rect 359 -776 374 -775
rect 478 -776 598 -775
rect 656 -776 1130 -775
rect 121 -778 762 -777
rect 870 -778 997 -777
rect 1024 -778 1130 -777
rect 177 -780 353 -779
rect 359 -780 398 -779
rect 432 -780 1025 -779
rect 205 -782 346 -781
rect 366 -782 451 -781
rect 492 -782 1109 -781
rect 184 -784 346 -783
rect 492 -784 794 -783
rect 870 -784 941 -783
rect 947 -784 1193 -783
rect 184 -786 304 -785
rect 520 -786 566 -785
rect 569 -786 1102 -785
rect 23 -788 521 -787
rect 523 -788 920 -787
rect 926 -788 941 -787
rect 954 -788 1011 -787
rect 219 -790 262 -789
rect 275 -790 451 -789
rect 527 -790 955 -789
rect 961 -790 1004 -789
rect 261 -792 283 -791
rect 527 -792 787 -791
rect 877 -792 927 -791
rect 201 -794 283 -793
rect 583 -794 948 -793
rect 268 -796 276 -795
rect 499 -796 584 -795
rect 586 -796 1123 -795
rect 268 -798 395 -797
rect 590 -798 619 -797
rect 653 -798 794 -797
rect 849 -798 878 -797
rect 898 -798 1004 -797
rect 163 -800 619 -799
rect 656 -800 1053 -799
rect 387 -802 395 -801
rect 429 -802 899 -801
rect 919 -802 983 -801
rect 429 -804 1137 -803
rect 597 -806 675 -805
rect 688 -806 787 -805
rect 814 -806 850 -805
rect 884 -806 983 -805
rect 58 -808 689 -807
rect 702 -808 892 -807
rect 58 -810 73 -809
rect 404 -810 675 -809
rect 779 -810 892 -809
rect 72 -812 290 -811
rect 471 -812 780 -811
rect 800 -812 815 -811
rect 863 -812 885 -811
rect 317 -814 472 -813
rect 604 -814 801 -813
rect 842 -814 864 -813
rect 226 -816 318 -815
rect 548 -816 605 -815
rect 667 -816 731 -815
rect 835 -816 843 -815
rect 226 -818 248 -817
rect 541 -818 549 -817
rect 660 -818 668 -817
rect 807 -818 836 -817
rect 247 -820 325 -819
rect 509 -820 542 -819
rect 562 -820 661 -819
rect 758 -820 808 -819
rect 324 -822 332 -821
rect 562 -822 622 -821
rect 758 -822 1067 -821
rect 296 -824 332 -823
rect 1031 -824 1067 -823
rect 296 -826 1074 -825
rect 432 -828 1032 -827
rect 1038 -828 1074 -827
rect 772 -830 1039 -829
rect 310 -832 773 -831
rect 16 -843 636 -842
rect 649 -843 780 -842
rect 824 -843 1249 -842
rect 1416 -843 1438 -842
rect 16 -845 59 -844
rect 68 -845 339 -844
rect 390 -845 899 -844
rect 961 -845 965 -844
rect 26 -847 45 -846
rect 58 -847 164 -846
rect 170 -847 433 -846
rect 439 -847 1137 -846
rect 30 -849 94 -848
rect 124 -849 1144 -848
rect 30 -851 416 -850
rect 425 -851 787 -850
rect 828 -851 1221 -850
rect 33 -853 948 -852
rect 961 -853 990 -852
rect 1143 -853 1200 -852
rect 37 -855 521 -854
rect 537 -855 577 -854
rect 586 -855 1011 -854
rect 1129 -855 1200 -854
rect 37 -857 52 -856
rect 72 -857 185 -856
rect 198 -857 402 -856
rect 443 -857 517 -856
rect 544 -857 626 -856
rect 653 -857 892 -856
rect 898 -857 941 -856
rect 947 -857 969 -856
rect 1010 -857 1053 -856
rect 44 -859 738 -858
rect 758 -859 1228 -858
rect 51 -861 202 -860
rect 205 -861 584 -860
rect 618 -861 1004 -860
rect 1052 -861 1203 -860
rect 65 -863 73 -862
rect 79 -863 584 -862
rect 611 -863 619 -862
rect 625 -863 1172 -862
rect 65 -865 101 -864
rect 121 -865 416 -864
rect 443 -865 696 -864
rect 702 -865 1039 -864
rect 1164 -865 1172 -864
rect 79 -867 479 -866
rect 485 -867 521 -866
rect 565 -867 1088 -866
rect 86 -869 829 -868
rect 856 -869 941 -868
rect 964 -869 990 -868
rect 1003 -869 1046 -868
rect 1059 -869 1165 -868
rect 9 -871 87 -870
rect 89 -871 304 -870
rect 380 -871 402 -870
rect 471 -871 486 -870
rect 506 -871 955 -870
rect 968 -871 1074 -870
rect 1087 -871 1123 -870
rect 2 -873 304 -872
rect 331 -873 381 -872
rect 397 -873 1158 -872
rect 23 -875 857 -874
rect 982 -875 1123 -874
rect 23 -877 496 -876
rect 509 -877 661 -876
rect 674 -877 1060 -876
rect 93 -879 216 -878
rect 240 -879 395 -878
rect 408 -879 507 -878
rect 569 -879 1179 -878
rect 100 -881 500 -880
rect 572 -881 759 -880
rect 761 -881 955 -880
rect 1017 -881 1046 -880
rect 121 -883 675 -882
rect 688 -883 1130 -882
rect 131 -885 1179 -884
rect 152 -887 983 -886
rect 1017 -887 1067 -886
rect 156 -889 332 -888
rect 369 -889 395 -888
rect 422 -889 472 -888
rect 478 -889 913 -888
rect 1031 -889 1039 -888
rect 2 -891 423 -890
rect 499 -891 976 -890
rect 1031 -891 1081 -890
rect 156 -893 713 -892
rect 723 -893 738 -892
rect 765 -893 1067 -892
rect 1080 -893 1116 -892
rect 89 -895 1116 -894
rect 131 -897 724 -896
rect 730 -897 780 -896
rect 786 -897 864 -896
rect 919 -897 976 -896
rect 163 -899 192 -898
rect 198 -899 241 -898
rect 254 -899 388 -898
rect 611 -899 1193 -898
rect 114 -901 192 -900
rect 205 -901 290 -900
rect 296 -901 346 -900
rect 632 -901 661 -900
rect 695 -901 717 -900
rect 765 -901 801 -900
rect 807 -901 892 -900
rect 919 -901 927 -900
rect 1094 -901 1193 -900
rect 107 -903 115 -902
rect 170 -903 405 -902
rect 569 -903 633 -902
rect 646 -903 1074 -902
rect 1094 -903 1151 -902
rect 107 -905 360 -904
rect 590 -905 647 -904
rect 653 -905 997 -904
rect 1150 -905 1207 -904
rect 177 -907 276 -906
rect 282 -907 321 -906
rect 345 -907 563 -906
rect 614 -907 927 -906
rect 996 -907 1025 -906
rect 1185 -907 1207 -906
rect 180 -909 682 -908
rect 702 -909 843 -908
rect 863 -909 934 -908
rect 1024 -909 1102 -908
rect 1185 -909 1235 -908
rect 184 -911 692 -910
rect 709 -911 731 -910
rect 751 -911 801 -910
rect 807 -911 815 -910
rect 870 -911 934 -910
rect 212 -913 360 -912
rect 513 -913 815 -912
rect 870 -913 1263 -912
rect 212 -915 430 -914
rect 555 -915 591 -914
rect 656 -915 906 -914
rect 219 -917 297 -916
rect 299 -917 388 -916
rect 450 -917 556 -916
rect 562 -917 748 -916
rect 772 -917 1242 -916
rect 219 -919 503 -918
rect 527 -919 773 -918
rect 775 -919 843 -918
rect 247 -921 255 -920
rect 261 -921 276 -920
rect 282 -921 437 -920
rect 450 -921 1137 -920
rect 247 -923 832 -922
rect 261 -925 367 -924
rect 373 -925 514 -924
rect 576 -925 657 -924
rect 667 -925 682 -924
rect 709 -925 1256 -924
rect 226 -927 367 -926
rect 436 -927 542 -926
rect 597 -927 906 -926
rect 135 -929 227 -928
rect 268 -929 339 -928
rect 352 -929 430 -928
rect 541 -929 850 -928
rect 135 -931 493 -930
rect 548 -931 598 -930
rect 639 -931 668 -930
rect 716 -931 1109 -930
rect 142 -933 353 -932
rect 457 -933 549 -932
rect 604 -933 640 -932
rect 688 -933 1109 -932
rect 142 -935 706 -934
rect 719 -935 1102 -934
rect 149 -937 493 -936
rect 534 -937 605 -936
rect 744 -937 752 -936
rect 793 -937 913 -936
rect 268 -939 482 -938
rect 534 -939 1158 -938
rect 289 -941 325 -940
rect 457 -941 465 -940
rect 793 -941 836 -940
rect 849 -941 878 -940
rect 310 -943 374 -942
rect 464 -943 524 -942
rect 821 -943 836 -942
rect 877 -943 885 -942
rect 75 -945 311 -944
rect 317 -945 409 -944
rect 821 -945 1214 -944
rect 9 -947 318 -946
rect 324 -947 629 -946
rect 128 -949 885 -948
rect 2 -960 150 -959
rect 152 -960 440 -959
rect 502 -960 682 -959
rect 688 -960 920 -959
rect 929 -960 1326 -959
rect 1437 -960 1445 -959
rect 5 -962 409 -961
rect 541 -962 1263 -961
rect 9 -964 423 -963
rect 548 -964 713 -963
rect 719 -964 1291 -963
rect 16 -966 90 -965
rect 103 -966 717 -965
rect 744 -966 1123 -965
rect 1136 -966 1270 -965
rect 16 -968 535 -967
rect 558 -968 787 -967
rect 863 -968 1137 -967
rect 1143 -968 1305 -967
rect 30 -970 538 -969
rect 565 -970 1060 -969
rect 1073 -970 1221 -969
rect 2 -972 31 -971
rect 33 -972 773 -971
rect 866 -972 969 -971
rect 1087 -972 1214 -971
rect 44 -974 318 -973
rect 320 -974 423 -973
rect 502 -974 787 -973
rect 877 -974 1123 -973
rect 1157 -974 1312 -973
rect 44 -976 171 -975
rect 201 -976 388 -975
rect 611 -976 1277 -975
rect 37 -978 171 -977
rect 212 -978 727 -977
rect 744 -978 864 -977
rect 870 -978 878 -977
rect 912 -978 920 -977
rect 954 -978 1074 -977
rect 1094 -978 1249 -977
rect 75 -980 661 -979
rect 667 -980 773 -979
rect 849 -980 955 -979
rect 961 -980 1256 -979
rect 51 -982 661 -981
rect 695 -982 1298 -981
rect 51 -984 885 -983
rect 968 -984 1011 -983
rect 1052 -984 1095 -983
rect 1101 -984 1235 -983
rect 79 -986 451 -985
rect 572 -986 871 -985
rect 884 -986 941 -985
rect 975 -986 1088 -985
rect 1115 -986 1242 -985
rect 23 -988 451 -987
rect 576 -988 913 -987
rect 933 -988 1053 -987
rect 1150 -988 1158 -987
rect 1164 -988 1319 -987
rect 23 -990 269 -989
rect 282 -990 426 -989
rect 436 -990 696 -989
rect 702 -990 934 -989
rect 1003 -990 1116 -989
rect 1185 -990 1340 -989
rect 79 -992 220 -991
rect 254 -992 615 -991
rect 618 -992 689 -991
rect 709 -992 1060 -991
rect 1192 -992 1207 -991
rect 114 -994 132 -993
rect 149 -994 409 -993
rect 436 -994 577 -993
rect 611 -994 822 -993
rect 856 -994 1102 -993
rect 96 -996 115 -995
rect 124 -996 654 -995
rect 723 -996 941 -995
rect 1017 -996 1151 -995
rect 177 -998 255 -997
rect 264 -998 479 -997
rect 499 -998 857 -997
rect 891 -998 976 -997
rect 982 -998 1018 -997
rect 1045 -998 1186 -997
rect 177 -1000 241 -999
rect 268 -1000 454 -999
rect 471 -1000 983 -999
rect 1066 -1000 1193 -999
rect 205 -1002 213 -1001
rect 219 -1002 1196 -1001
rect 240 -1004 325 -1003
rect 338 -1004 388 -1003
rect 471 -1004 507 -1003
rect 513 -1004 654 -1003
rect 723 -1004 962 -1003
rect 1080 -1004 1207 -1003
rect 282 -1006 416 -1005
rect 478 -1006 1109 -1005
rect 289 -1008 325 -1007
rect 341 -1008 402 -1007
rect 499 -1008 549 -1007
rect 555 -1008 619 -1007
rect 628 -1008 738 -1007
rect 747 -1008 780 -1007
rect 800 -1008 822 -1007
rect 835 -1008 892 -1007
rect 926 -1008 1046 -1007
rect 1080 -1008 1130 -1007
rect 128 -1010 738 -1009
rect 747 -1010 1228 -1009
rect 37 -1012 129 -1011
rect 142 -1012 290 -1011
rect 303 -1012 416 -1011
rect 506 -1012 563 -1011
rect 632 -1012 1333 -1011
rect 86 -1014 304 -1013
rect 306 -1014 311 -1013
rect 317 -1014 482 -1013
rect 513 -1014 647 -1013
rect 656 -1014 801 -1013
rect 814 -1014 850 -1013
rect 996 -1014 1109 -1013
rect 86 -1016 545 -1015
rect 597 -1016 647 -1015
rect 751 -1016 780 -1015
rect 807 -1016 815 -1015
rect 989 -1016 997 -1015
rect 1031 -1016 1130 -1015
rect 40 -1018 598 -1017
rect 635 -1018 1347 -1017
rect 310 -1020 339 -1019
rect 345 -1020 703 -1019
rect 730 -1020 752 -1019
rect 758 -1020 1004 -1019
rect 345 -1022 374 -1021
rect 376 -1022 1179 -1021
rect 352 -1024 531 -1023
rect 569 -1024 759 -1023
rect 765 -1024 1144 -1023
rect 9 -1026 531 -1025
rect 569 -1026 605 -1025
rect 639 -1026 682 -1025
rect 793 -1026 990 -1025
rect 1024 -1026 1179 -1025
rect 261 -1028 353 -1027
rect 359 -1028 668 -1027
rect 677 -1028 766 -1027
rect 793 -1028 825 -1027
rect 898 -1028 1025 -1027
rect 68 -1030 899 -1029
rect 905 -1030 1032 -1029
rect 107 -1032 360 -1031
rect 366 -1032 1011 -1031
rect 107 -1034 626 -1033
rect 842 -1034 906 -1033
rect 100 -1036 843 -1035
rect 100 -1038 1039 -1037
rect 296 -1040 640 -1039
rect 947 -1040 1039 -1039
rect 135 -1042 297 -1041
rect 366 -1042 1200 -1041
rect 65 -1044 136 -1043
rect 369 -1044 1284 -1043
rect 65 -1046 496 -1045
rect 520 -1046 1067 -1045
rect 373 -1048 395 -1047
rect 401 -1048 458 -1047
rect 464 -1048 731 -1047
rect 828 -1048 948 -1047
rect 191 -1050 395 -1049
rect 429 -1050 458 -1049
rect 481 -1050 1200 -1049
rect 163 -1052 192 -1051
rect 261 -1052 465 -1051
rect 492 -1052 521 -1051
rect 527 -1052 1165 -1051
rect 163 -1054 927 -1053
rect 184 -1056 430 -1055
rect 492 -1056 836 -1055
rect 184 -1058 248 -1057
rect 380 -1058 542 -1057
rect 583 -1058 808 -1057
rect 233 -1060 248 -1059
rect 380 -1060 517 -1059
rect 527 -1060 710 -1059
rect 54 -1062 234 -1061
rect 534 -1062 626 -1061
rect 674 -1062 829 -1061
rect 443 -1064 675 -1063
rect 93 -1066 444 -1065
rect 583 -1066 636 -1065
rect 93 -1068 143 -1067
rect 590 -1068 605 -1067
rect 226 -1070 591 -1069
rect 226 -1072 276 -1071
rect 58 -1074 276 -1073
rect 58 -1076 73 -1075
rect 72 -1078 206 -1077
rect 2 -1089 983 -1088
rect 1241 -1089 1368 -1088
rect 1444 -1089 1452 -1088
rect 9 -1091 339 -1090
rect 404 -1091 668 -1090
rect 674 -1091 1270 -1090
rect 1318 -1091 1354 -1090
rect 9 -1093 34 -1092
rect 37 -1093 122 -1092
rect 149 -1093 227 -1092
rect 247 -1093 265 -1092
rect 439 -1093 521 -1092
rect 527 -1093 1144 -1092
rect 1213 -1093 1242 -1092
rect 1325 -1093 1361 -1092
rect 30 -1095 563 -1094
rect 569 -1095 1319 -1094
rect 1339 -1095 1375 -1094
rect 54 -1097 843 -1096
rect 845 -1097 983 -1096
rect 1220 -1097 1270 -1096
rect 1311 -1097 1340 -1096
rect 58 -1099 101 -1098
rect 121 -1099 290 -1098
rect 408 -1099 563 -1098
rect 572 -1099 773 -1098
rect 786 -1099 1312 -1098
rect 58 -1101 178 -1100
rect 212 -1101 524 -1100
rect 530 -1101 619 -1100
rect 628 -1101 1137 -1100
rect 1192 -1101 1221 -1100
rect 75 -1103 1102 -1102
rect 75 -1105 661 -1104
rect 667 -1105 731 -1104
rect 733 -1105 1137 -1104
rect 79 -1107 545 -1106
rect 558 -1107 766 -1106
rect 863 -1107 1326 -1106
rect 79 -1109 444 -1108
rect 471 -1109 636 -1108
rect 653 -1109 675 -1108
rect 684 -1109 1207 -1108
rect 93 -1111 517 -1110
rect 541 -1111 570 -1110
rect 576 -1111 724 -1110
rect 726 -1111 1151 -1110
rect 1178 -1111 1207 -1110
rect 93 -1113 171 -1112
rect 177 -1113 297 -1112
rect 310 -1113 444 -1112
rect 450 -1113 654 -1112
rect 660 -1113 762 -1112
rect 765 -1113 1235 -1112
rect 72 -1115 171 -1114
rect 205 -1115 472 -1114
rect 478 -1115 486 -1114
rect 492 -1115 990 -1114
rect 1087 -1115 1102 -1114
rect 1150 -1115 1158 -1114
rect 44 -1117 479 -1116
rect 499 -1117 878 -1116
rect 929 -1117 1305 -1116
rect 44 -1119 381 -1118
rect 408 -1119 423 -1118
rect 457 -1119 486 -1118
rect 499 -1119 612 -1118
rect 632 -1119 1249 -1118
rect 1290 -1119 1305 -1118
rect 23 -1121 381 -1120
rect 394 -1121 423 -1120
rect 457 -1121 507 -1120
rect 541 -1121 1298 -1120
rect 23 -1123 367 -1122
rect 464 -1123 612 -1122
rect 695 -1123 755 -1122
rect 828 -1123 878 -1122
rect 954 -1123 1144 -1122
rect 1227 -1123 1249 -1122
rect 1283 -1123 1298 -1122
rect 72 -1125 759 -1124
rect 821 -1125 829 -1124
rect 849 -1125 990 -1124
rect 1045 -1125 1088 -1124
rect 1171 -1125 1284 -1124
rect 96 -1127 640 -1126
rect 681 -1127 696 -1126
rect 712 -1127 1193 -1126
rect 1199 -1127 1228 -1126
rect 100 -1129 850 -1128
rect 866 -1129 1186 -1128
rect 117 -1131 1186 -1130
rect 128 -1133 395 -1132
rect 464 -1133 1277 -1132
rect 128 -1135 633 -1134
rect 716 -1135 724 -1134
rect 730 -1135 1116 -1134
rect 1262 -1135 1277 -1134
rect 149 -1137 647 -1136
rect 702 -1137 717 -1136
rect 744 -1137 836 -1136
rect 870 -1137 1179 -1136
rect 163 -1139 206 -1138
rect 212 -1139 678 -1138
rect 688 -1139 703 -1138
rect 744 -1139 1123 -1138
rect 163 -1141 496 -1140
rect 502 -1141 1067 -1140
rect 1073 -1141 1116 -1140
rect 226 -1143 276 -1142
rect 282 -1143 528 -1142
rect 548 -1143 577 -1142
rect 600 -1143 1256 -1142
rect 152 -1145 276 -1144
rect 289 -1145 468 -1144
rect 495 -1145 871 -1144
rect 905 -1145 955 -1144
rect 968 -1145 1158 -1144
rect 1255 -1145 1333 -1144
rect 184 -1147 283 -1146
rect 296 -1147 353 -1146
rect 373 -1147 640 -1146
rect 649 -1147 689 -1146
rect 747 -1147 941 -1146
rect 1010 -1147 1046 -1146
rect 1066 -1147 1130 -1146
rect 103 -1149 374 -1148
rect 506 -1149 797 -1148
rect 800 -1149 822 -1148
rect 856 -1149 906 -1148
rect 933 -1149 1074 -1148
rect 1080 -1149 1263 -1148
rect 5 -1151 857 -1150
rect 891 -1151 941 -1150
rect 961 -1151 1011 -1150
rect 1017 -1151 1172 -1150
rect 5 -1153 1291 -1152
rect 103 -1155 216 -1154
rect 233 -1155 451 -1154
rect 534 -1155 969 -1154
rect 1017 -1155 1095 -1154
rect 1108 -1155 1333 -1154
rect 135 -1157 234 -1156
rect 240 -1157 248 -1156
rect 254 -1157 377 -1156
rect 534 -1157 647 -1156
rect 709 -1157 892 -1156
rect 912 -1157 962 -1156
rect 1031 -1157 1200 -1156
rect 40 -1159 136 -1158
rect 156 -1159 185 -1158
rect 240 -1159 584 -1158
rect 604 -1159 619 -1158
rect 747 -1159 1081 -1158
rect 156 -1161 437 -1160
rect 481 -1161 584 -1160
rect 607 -1161 1165 -1160
rect 261 -1163 787 -1162
rect 814 -1163 934 -1162
rect 1052 -1163 1095 -1162
rect 191 -1165 262 -1164
rect 303 -1165 836 -1164
rect 884 -1165 1109 -1164
rect 142 -1167 192 -1166
rect 219 -1167 304 -1166
rect 310 -1167 598 -1166
rect 751 -1167 801 -1166
rect 807 -1167 885 -1166
rect 919 -1167 1032 -1166
rect 1059 -1167 1130 -1166
rect 107 -1169 143 -1168
rect 219 -1169 556 -1168
rect 558 -1169 1123 -1168
rect 107 -1171 199 -1170
rect 317 -1171 367 -1170
rect 401 -1171 437 -1170
rect 513 -1171 1053 -1170
rect 180 -1173 514 -1172
rect 530 -1173 1165 -1172
rect 198 -1175 269 -1174
rect 317 -1175 325 -1174
rect 341 -1175 353 -1174
rect 359 -1175 808 -1174
rect 1024 -1175 1060 -1174
rect 254 -1177 402 -1176
rect 555 -1177 1214 -1176
rect 268 -1179 430 -1178
rect 565 -1179 773 -1178
rect 779 -1179 913 -1178
rect 975 -1179 1025 -1178
rect 324 -1181 346 -1180
rect 359 -1181 682 -1180
rect 751 -1181 927 -1180
rect 975 -1181 1039 -1180
rect 331 -1183 780 -1182
rect 793 -1183 815 -1182
rect 1003 -1183 1039 -1182
rect 331 -1185 416 -1184
rect 429 -1185 636 -1184
rect 758 -1185 1347 -1184
rect 51 -1187 1347 -1186
rect 345 -1189 738 -1188
rect 793 -1189 864 -1188
rect 996 -1189 1004 -1188
rect 65 -1191 738 -1190
rect 947 -1191 997 -1190
rect 65 -1193 87 -1192
rect 387 -1193 416 -1192
rect 597 -1193 1235 -1192
rect 86 -1195 115 -1194
rect 387 -1195 493 -1194
rect 625 -1195 920 -1194
rect 51 -1197 626 -1196
rect 898 -1197 948 -1196
rect 114 -1199 591 -1198
rect 551 -1201 899 -1200
rect 590 -1203 710 -1202
rect 2 -1214 304 -1213
rect 366 -1214 559 -1213
rect 607 -1214 969 -1213
rect 1017 -1214 1021 -1213
rect 1269 -1214 1273 -1213
rect 1360 -1214 1382 -1213
rect 1451 -1214 1459 -1213
rect 5 -1216 780 -1215
rect 793 -1216 850 -1215
rect 870 -1216 969 -1215
rect 1017 -1216 1116 -1215
rect 1269 -1216 1284 -1215
rect 30 -1218 552 -1217
rect 614 -1218 619 -1217
rect 628 -1218 696 -1217
rect 698 -1218 1074 -1217
rect 1283 -1218 1319 -1217
rect 30 -1220 563 -1219
rect 632 -1220 1144 -1219
rect 1272 -1220 1319 -1219
rect 37 -1222 213 -1221
rect 289 -1222 563 -1221
rect 646 -1222 1375 -1221
rect 37 -1224 59 -1223
rect 72 -1224 122 -1223
rect 124 -1224 353 -1223
rect 366 -1224 636 -1223
rect 653 -1224 1389 -1223
rect 44 -1226 650 -1225
rect 653 -1226 717 -1225
rect 719 -1226 1144 -1225
rect 44 -1228 94 -1227
rect 100 -1228 118 -1227
rect 121 -1228 556 -1227
rect 600 -1228 647 -1227
rect 684 -1228 1298 -1227
rect 51 -1230 94 -1229
rect 138 -1230 570 -1229
rect 709 -1230 738 -1229
rect 751 -1230 1375 -1229
rect 51 -1232 419 -1231
rect 432 -1232 535 -1231
rect 544 -1232 1361 -1231
rect 58 -1234 479 -1233
rect 492 -1234 885 -1233
rect 915 -1234 1081 -1233
rect 1150 -1234 1298 -1233
rect 75 -1236 423 -1235
rect 436 -1236 465 -1235
rect 520 -1236 710 -1235
rect 712 -1236 1095 -1235
rect 1150 -1236 1158 -1235
rect 89 -1238 227 -1237
rect 289 -1238 374 -1237
rect 394 -1238 531 -1237
rect 534 -1238 706 -1237
rect 754 -1238 1340 -1237
rect 149 -1240 598 -1239
rect 604 -1240 885 -1239
rect 1010 -1240 1074 -1239
rect 1080 -1240 1109 -1239
rect 1157 -1240 1172 -1239
rect 149 -1242 346 -1241
rect 352 -1242 388 -1241
rect 436 -1242 542 -1241
rect 548 -1242 997 -1241
rect 1010 -1242 1039 -1241
rect 1094 -1242 1179 -1241
rect 173 -1244 1200 -1243
rect 177 -1246 255 -1245
rect 282 -1246 388 -1245
rect 446 -1246 1200 -1245
rect 191 -1248 304 -1247
rect 310 -1248 619 -1247
rect 660 -1248 752 -1247
rect 765 -1248 1025 -1247
rect 1038 -1248 1046 -1247
rect 1129 -1248 1172 -1247
rect 1178 -1248 1193 -1247
rect 170 -1250 192 -1249
rect 198 -1250 682 -1249
rect 695 -1250 738 -1249
rect 758 -1250 1046 -1249
rect 1164 -1250 1340 -1249
rect 198 -1252 297 -1251
rect 310 -1252 496 -1251
rect 520 -1252 573 -1251
rect 604 -1252 612 -1251
rect 660 -1252 703 -1251
rect 758 -1252 787 -1251
rect 796 -1252 1207 -1251
rect 205 -1254 395 -1253
rect 450 -1254 493 -1253
rect 527 -1254 1235 -1253
rect 135 -1256 206 -1255
rect 212 -1256 318 -1255
rect 331 -1256 423 -1255
rect 464 -1256 472 -1255
rect 527 -1256 545 -1255
rect 548 -1256 734 -1255
rect 765 -1256 808 -1255
rect 842 -1256 1263 -1255
rect 135 -1258 1221 -1257
rect 1234 -1258 1249 -1257
rect 219 -1260 598 -1259
rect 621 -1260 1249 -1259
rect 156 -1262 220 -1261
rect 226 -1262 468 -1261
rect 555 -1262 577 -1261
rect 681 -1262 1368 -1261
rect 103 -1264 157 -1263
rect 233 -1264 283 -1263
rect 296 -1264 409 -1263
rect 457 -1264 472 -1263
rect 569 -1264 1333 -1263
rect 1353 -1264 1368 -1263
rect 16 -1266 458 -1265
rect 576 -1266 591 -1265
rect 779 -1266 801 -1265
rect 807 -1266 822 -1265
rect 828 -1266 843 -1265
rect 845 -1266 955 -1265
rect 989 -1266 997 -1265
rect 1003 -1266 1130 -1265
rect 1164 -1266 1186 -1265
rect 1332 -1266 1347 -1265
rect 16 -1268 640 -1267
rect 786 -1268 836 -1267
rect 849 -1268 892 -1267
rect 961 -1268 990 -1267
rect 1003 -1268 1032 -1267
rect 1066 -1268 1207 -1267
rect 1255 -1268 1347 -1267
rect 61 -1270 1354 -1269
rect 170 -1272 1067 -1271
rect 1087 -1272 1221 -1271
rect 1255 -1272 1277 -1271
rect 233 -1274 507 -1273
rect 625 -1274 836 -1273
rect 866 -1274 1263 -1273
rect 1276 -1274 1291 -1273
rect 240 -1276 451 -1275
rect 485 -1276 507 -1275
rect 583 -1276 626 -1275
rect 639 -1276 675 -1275
rect 800 -1276 899 -1275
rect 933 -1276 962 -1275
rect 975 -1276 1032 -1275
rect 1087 -1276 1102 -1275
rect 1122 -1276 1186 -1275
rect 1290 -1276 1326 -1275
rect 68 -1278 1123 -1277
rect 1311 -1278 1326 -1277
rect 114 -1280 1102 -1279
rect 65 -1282 115 -1281
rect 240 -1282 633 -1281
rect 744 -1282 934 -1281
rect 1024 -1282 1053 -1281
rect 247 -1284 318 -1283
rect 324 -1284 486 -1283
rect 499 -1284 675 -1283
rect 730 -1284 1053 -1283
rect 79 -1286 500 -1285
rect 583 -1286 769 -1285
rect 821 -1286 857 -1285
rect 870 -1286 948 -1285
rect 79 -1288 255 -1287
rect 331 -1288 430 -1287
rect 443 -1288 591 -1287
rect 730 -1288 1060 -1287
rect 107 -1290 444 -1289
rect 513 -1290 948 -1289
rect 1059 -1290 1228 -1289
rect 86 -1292 108 -1291
rect 184 -1292 325 -1291
rect 338 -1292 479 -1291
rect 513 -1292 689 -1291
rect 744 -1292 818 -1291
rect 828 -1292 927 -1291
rect 1213 -1292 1228 -1291
rect 86 -1294 1109 -1293
rect 1213 -1294 1242 -1293
rect 184 -1296 734 -1295
rect 747 -1296 976 -1295
rect 247 -1298 612 -1297
rect 688 -1298 724 -1297
rect 856 -1298 864 -1297
rect 891 -1298 906 -1297
rect 338 -1300 402 -1299
rect 523 -1300 1242 -1299
rect 9 -1302 402 -1301
rect 702 -1302 927 -1301
rect 9 -1304 773 -1303
rect 863 -1304 1312 -1303
rect 345 -1306 416 -1305
rect 772 -1306 815 -1305
rect 898 -1306 955 -1305
rect 268 -1308 416 -1307
rect 814 -1308 1137 -1307
rect 268 -1310 360 -1309
rect 369 -1310 1193 -1309
rect 359 -1312 542 -1311
rect 905 -1312 920 -1311
rect 376 -1314 724 -1313
rect 912 -1314 920 -1313
rect 380 -1316 409 -1315
rect 761 -1316 913 -1315
rect 23 -1318 381 -1317
rect 404 -1318 1137 -1317
rect 23 -1320 129 -1319
rect 128 -1322 276 -1321
rect 275 -1324 391 -1323
rect 33 -1335 108 -1334
rect 121 -1335 1354 -1334
rect 1423 -1335 1452 -1334
rect 1458 -1335 1466 -1334
rect 44 -1337 374 -1336
rect 387 -1337 1067 -1336
rect 1122 -1337 1403 -1336
rect 44 -1339 752 -1338
rect 814 -1339 1228 -1338
rect 1255 -1339 1354 -1338
rect 1360 -1339 1459 -1338
rect 65 -1341 556 -1340
rect 583 -1341 619 -1340
rect 635 -1341 878 -1340
rect 887 -1341 1375 -1340
rect 65 -1343 125 -1342
rect 135 -1343 1431 -1342
rect 61 -1345 136 -1344
rect 163 -1345 783 -1344
rect 793 -1345 878 -1344
rect 898 -1345 1074 -1344
rect 1129 -1345 1410 -1344
rect 68 -1347 447 -1346
rect 464 -1347 570 -1346
rect 614 -1347 1081 -1346
rect 1150 -1347 1228 -1346
rect 1262 -1347 1361 -1346
rect 30 -1349 570 -1348
rect 646 -1349 818 -1348
rect 821 -1349 899 -1348
rect 912 -1349 1368 -1348
rect 79 -1351 325 -1350
rect 380 -1351 447 -1350
rect 509 -1351 1305 -1350
rect 1332 -1351 1438 -1350
rect 82 -1353 1221 -1352
rect 1234 -1353 1333 -1352
rect 1339 -1353 1375 -1352
rect 82 -1355 748 -1354
rect 821 -1355 1249 -1354
rect 1269 -1355 1368 -1354
rect 86 -1357 101 -1356
rect 107 -1357 367 -1356
rect 380 -1357 685 -1356
rect 695 -1357 724 -1356
rect 852 -1357 1053 -1356
rect 1094 -1357 1249 -1356
rect 1297 -1357 1417 -1356
rect 86 -1359 220 -1358
rect 254 -1359 367 -1358
rect 376 -1359 1053 -1358
rect 1059 -1359 1298 -1358
rect 1318 -1359 1340 -1358
rect 1346 -1359 1445 -1358
rect 100 -1361 297 -1360
rect 317 -1361 374 -1360
rect 415 -1361 1312 -1360
rect 23 -1363 297 -1362
rect 324 -1363 332 -1362
rect 418 -1363 857 -1362
rect 866 -1363 969 -1362
rect 982 -1363 1067 -1362
rect 1157 -1363 1221 -1362
rect 1241 -1363 1347 -1362
rect 23 -1365 248 -1364
rect 429 -1365 860 -1364
rect 968 -1365 976 -1364
rect 996 -1365 1074 -1364
rect 1164 -1365 1235 -1364
rect 37 -1367 318 -1366
rect 429 -1367 573 -1366
rect 583 -1367 647 -1366
rect 649 -1367 1039 -1366
rect 1045 -1367 1049 -1366
rect 1164 -1367 1172 -1366
rect 1178 -1367 1263 -1366
rect 37 -1369 535 -1368
rect 541 -1369 948 -1368
rect 954 -1369 1039 -1368
rect 1045 -1369 1389 -1368
rect 93 -1371 332 -1370
rect 436 -1371 696 -1370
rect 698 -1371 955 -1370
rect 1017 -1371 1130 -1370
rect 1192 -1371 1256 -1370
rect 1276 -1371 1389 -1370
rect 93 -1373 461 -1372
rect 534 -1373 556 -1372
rect 632 -1373 1312 -1372
rect 121 -1375 150 -1374
rect 152 -1375 416 -1374
rect 436 -1375 458 -1374
rect 541 -1375 787 -1374
rect 793 -1375 983 -1374
rect 1024 -1375 1095 -1374
rect 1101 -1375 1172 -1374
rect 1192 -1375 1284 -1374
rect 128 -1377 255 -1376
rect 443 -1377 1158 -1376
rect 1199 -1377 1284 -1376
rect 128 -1379 311 -1378
rect 457 -1379 1319 -1378
rect 131 -1381 1270 -1380
rect 149 -1383 591 -1382
rect 632 -1383 857 -1382
rect 870 -1383 1025 -1382
rect 1031 -1383 1123 -1382
rect 1199 -1383 1291 -1382
rect 163 -1385 412 -1384
rect 527 -1385 871 -1384
rect 884 -1385 948 -1384
rect 1010 -1385 1102 -1384
rect 1206 -1385 1277 -1384
rect 170 -1387 913 -1386
rect 933 -1387 997 -1386
rect 1143 -1387 1207 -1386
rect 170 -1389 682 -1388
rect 702 -1389 990 -1388
rect 1048 -1389 1144 -1388
rect 198 -1391 398 -1390
rect 513 -1391 682 -1390
rect 705 -1391 962 -1390
rect 184 -1393 199 -1392
rect 212 -1393 370 -1392
rect 394 -1393 528 -1392
rect 544 -1393 661 -1392
rect 667 -1393 752 -1392
rect 758 -1393 787 -1392
rect 814 -1393 1291 -1392
rect 184 -1395 241 -1394
rect 247 -1395 566 -1394
rect 590 -1395 654 -1394
rect 667 -1395 801 -1394
rect 828 -1395 1011 -1394
rect 191 -1397 213 -1396
rect 219 -1397 321 -1396
rect 401 -1397 514 -1396
rect 551 -1397 1081 -1396
rect 2 -1399 192 -1398
rect 240 -1399 486 -1398
rect 492 -1399 654 -1398
rect 716 -1399 780 -1398
rect 831 -1399 1179 -1398
rect 2 -1401 52 -1400
rect 275 -1401 801 -1400
rect 842 -1401 934 -1400
rect 940 -1401 1018 -1400
rect 51 -1403 262 -1402
rect 275 -1403 549 -1402
rect 625 -1403 703 -1402
rect 716 -1403 745 -1402
rect 758 -1403 773 -1402
rect 779 -1403 1151 -1402
rect 79 -1405 262 -1404
rect 303 -1405 395 -1404
rect 450 -1405 486 -1404
rect 492 -1405 521 -1404
rect 548 -1405 1326 -1404
rect 89 -1407 941 -1406
rect 1213 -1407 1326 -1406
rect 138 -1409 843 -1408
rect 866 -1409 1032 -1408
rect 1185 -1409 1214 -1408
rect 282 -1411 451 -1410
rect 464 -1411 745 -1410
rect 891 -1411 962 -1410
rect 1115 -1411 1186 -1410
rect 282 -1413 290 -1412
rect 303 -1413 353 -1412
rect 520 -1413 1396 -1412
rect 289 -1415 766 -1414
rect 796 -1415 1116 -1414
rect 310 -1417 727 -1416
rect 730 -1417 1060 -1416
rect 352 -1419 360 -1418
rect 562 -1419 766 -1418
rect 905 -1419 976 -1418
rect 338 -1421 563 -1420
rect 597 -1421 626 -1420
rect 639 -1421 661 -1420
rect 688 -1421 731 -1420
rect 737 -1421 773 -1420
rect 905 -1421 1109 -1420
rect 166 -1423 598 -1422
rect 604 -1423 689 -1422
rect 709 -1423 738 -1422
rect 926 -1423 990 -1422
rect 1087 -1423 1109 -1422
rect 268 -1425 339 -1424
rect 359 -1425 500 -1424
rect 576 -1425 605 -1424
rect 642 -1425 892 -1424
rect 915 -1425 927 -1424
rect 1003 -1425 1088 -1424
rect 58 -1427 1004 -1426
rect 58 -1429 73 -1428
rect 114 -1429 269 -1428
rect 387 -1429 640 -1428
rect 674 -1429 710 -1428
rect 719 -1429 1382 -1428
rect 72 -1431 227 -1430
rect 499 -1431 507 -1430
rect 611 -1431 675 -1430
rect 723 -1431 1305 -1430
rect 16 -1433 612 -1432
rect 919 -1433 1382 -1432
rect 16 -1435 409 -1434
rect 506 -1435 1242 -1434
rect 114 -1437 346 -1436
rect 408 -1437 808 -1436
rect 835 -1437 920 -1436
rect 173 -1439 577 -1438
rect 807 -1439 850 -1438
rect 226 -1441 234 -1440
rect 345 -1441 423 -1440
rect 828 -1441 836 -1440
rect 156 -1443 234 -1442
rect 401 -1443 850 -1442
rect 156 -1445 178 -1444
rect 422 -1445 472 -1444
rect 142 -1447 178 -1446
rect 390 -1447 472 -1446
rect 142 -1449 825 -1448
rect 9 -1460 34 -1459
rect 44 -1460 458 -1459
rect 460 -1460 941 -1459
rect 1454 -1460 1466 -1459
rect 12 -1462 269 -1461
rect 282 -1462 521 -1461
rect 523 -1462 710 -1461
rect 723 -1462 836 -1461
rect 852 -1462 1277 -1461
rect 19 -1464 1403 -1463
rect 44 -1466 486 -1465
rect 520 -1466 689 -1465
rect 702 -1466 783 -1465
rect 793 -1466 1270 -1465
rect 51 -1468 510 -1467
rect 534 -1468 591 -1467
rect 621 -1468 1298 -1467
rect 51 -1470 731 -1469
rect 744 -1470 1228 -1469
rect 1269 -1470 1368 -1469
rect 65 -1472 538 -1471
rect 558 -1472 1011 -1471
rect 1297 -1472 1396 -1471
rect 65 -1474 871 -1473
rect 884 -1474 1039 -1473
rect 93 -1476 489 -1475
rect 534 -1476 668 -1475
rect 688 -1476 696 -1475
rect 705 -1476 1053 -1475
rect 37 -1478 94 -1477
rect 100 -1478 549 -1477
rect 562 -1478 1235 -1477
rect 37 -1480 899 -1479
rect 940 -1480 997 -1479
rect 1010 -1480 1074 -1479
rect 1234 -1480 1319 -1479
rect 103 -1482 451 -1481
rect 548 -1482 605 -1481
rect 639 -1482 1382 -1481
rect 107 -1484 118 -1483
rect 121 -1484 153 -1483
rect 180 -1484 731 -1483
rect 779 -1484 1333 -1483
rect 100 -1486 108 -1485
rect 121 -1486 416 -1485
rect 443 -1486 766 -1485
rect 793 -1486 843 -1485
rect 859 -1486 1326 -1485
rect 1332 -1486 1431 -1485
rect 128 -1488 1172 -1487
rect 1318 -1488 1417 -1487
rect 128 -1490 423 -1489
rect 446 -1490 1228 -1489
rect 1325 -1490 1424 -1489
rect 131 -1492 433 -1491
rect 450 -1492 654 -1491
rect 663 -1492 1452 -1491
rect 138 -1494 801 -1493
rect 814 -1494 1158 -1493
rect 1171 -1494 1256 -1493
rect 149 -1496 850 -1495
rect 863 -1496 1410 -1495
rect 149 -1498 171 -1497
rect 240 -1498 538 -1497
rect 562 -1498 619 -1497
rect 639 -1498 661 -1497
rect 667 -1498 738 -1497
rect 758 -1498 780 -1497
rect 796 -1498 1046 -1497
rect 1052 -1498 1102 -1497
rect 1157 -1498 1214 -1497
rect 72 -1500 171 -1499
rect 191 -1500 241 -1499
rect 261 -1500 605 -1499
rect 653 -1500 682 -1499
rect 702 -1500 1214 -1499
rect 58 -1502 73 -1501
rect 86 -1502 192 -1501
rect 254 -1502 262 -1501
rect 268 -1502 409 -1501
rect 415 -1502 612 -1501
rect 709 -1502 748 -1501
rect 765 -1502 787 -1501
rect 800 -1502 1347 -1501
rect 23 -1504 787 -1503
rect 814 -1504 878 -1503
rect 898 -1504 1095 -1503
rect 1192 -1504 1256 -1503
rect 1346 -1504 1445 -1503
rect 23 -1506 55 -1505
rect 58 -1506 311 -1505
rect 331 -1506 696 -1505
rect 716 -1506 745 -1505
rect 817 -1506 1088 -1505
rect 1094 -1506 1312 -1505
rect 16 -1508 311 -1507
rect 338 -1508 423 -1507
rect 478 -1508 619 -1507
rect 716 -1508 752 -1507
rect 821 -1508 895 -1507
rect 982 -1508 1277 -1507
rect 16 -1510 682 -1509
rect 723 -1510 773 -1509
rect 824 -1510 1375 -1509
rect 219 -1512 332 -1511
rect 338 -1512 500 -1511
rect 565 -1512 752 -1511
rect 828 -1512 1186 -1511
rect 1192 -1512 1291 -1511
rect 2 -1514 220 -1513
rect 247 -1514 255 -1513
rect 282 -1514 346 -1513
rect 380 -1514 444 -1513
rect 478 -1514 493 -1513
rect 572 -1514 867 -1513
rect 870 -1514 1018 -1513
rect 1038 -1514 1081 -1513
rect 1185 -1514 1284 -1513
rect 2 -1516 276 -1515
rect 289 -1516 773 -1515
rect 831 -1516 1123 -1515
rect 1199 -1516 1312 -1515
rect 9 -1518 276 -1517
rect 289 -1518 458 -1517
rect 485 -1518 759 -1517
rect 831 -1518 1361 -1517
rect 114 -1520 500 -1519
rect 583 -1520 643 -1519
rect 835 -1520 892 -1519
rect 905 -1520 1123 -1519
rect 1129 -1520 1200 -1519
rect 1283 -1520 1389 -1519
rect 40 -1522 584 -1521
rect 590 -1522 675 -1521
rect 842 -1522 913 -1521
rect 954 -1522 983 -1521
rect 996 -1522 1151 -1521
rect 89 -1524 913 -1523
rect 1059 -1524 1102 -1523
rect 1129 -1524 1179 -1523
rect 30 -1526 1179 -1525
rect 30 -1528 360 -1527
rect 380 -1528 598 -1527
rect 611 -1528 647 -1527
rect 649 -1528 675 -1527
rect 807 -1528 955 -1527
rect 1073 -1528 1305 -1527
rect 114 -1530 738 -1529
rect 849 -1530 920 -1529
rect 1080 -1530 1221 -1529
rect 1304 -1530 1340 -1529
rect 142 -1532 1018 -1531
rect 1115 -1532 1221 -1531
rect 1339 -1532 1438 -1531
rect 142 -1534 234 -1533
rect 317 -1534 1060 -1533
rect 1108 -1534 1116 -1533
rect 1150 -1534 1242 -1533
rect 198 -1536 248 -1535
rect 324 -1536 906 -1535
rect 919 -1536 962 -1535
rect 82 -1538 325 -1537
rect 345 -1538 367 -1537
rect 397 -1538 1137 -1537
rect 198 -1540 213 -1539
rect 233 -1540 304 -1539
rect 352 -1540 360 -1539
rect 366 -1540 577 -1539
rect 625 -1540 647 -1539
rect 859 -1540 1137 -1539
rect 177 -1542 213 -1541
rect 296 -1542 304 -1541
rect 352 -1542 374 -1541
rect 404 -1542 633 -1541
rect 863 -1542 934 -1541
rect 961 -1542 1025 -1541
rect 135 -1544 297 -1543
rect 373 -1544 388 -1543
rect 408 -1544 493 -1543
rect 513 -1544 577 -1543
rect 625 -1544 927 -1543
rect 933 -1544 990 -1543
rect 1024 -1544 1207 -1543
rect 79 -1546 514 -1545
rect 541 -1546 808 -1545
rect 877 -1546 948 -1545
rect 968 -1546 990 -1545
rect 1143 -1546 1207 -1545
rect 79 -1548 87 -1547
rect 135 -1548 1242 -1547
rect 205 -1550 318 -1549
rect 387 -1550 465 -1549
rect 541 -1550 570 -1549
rect 891 -1550 1263 -1549
rect 205 -1552 552 -1551
rect 555 -1552 598 -1551
rect 926 -1552 976 -1551
rect 1143 -1552 1165 -1551
rect 1262 -1552 1354 -1551
rect 394 -1554 465 -1553
rect 555 -1554 1046 -1553
rect 1353 -1554 1459 -1553
rect 394 -1556 437 -1555
rect 569 -1556 1291 -1555
rect 401 -1558 437 -1557
rect 856 -1558 976 -1557
rect 163 -1560 402 -1559
rect 429 -1560 633 -1559
rect 856 -1560 1109 -1559
rect 163 -1562 1004 -1561
rect 429 -1564 1088 -1563
rect 887 -1566 1165 -1565
rect 947 -1568 1049 -1567
rect 968 -1570 1032 -1569
rect 145 -1572 1032 -1571
rect 1003 -1574 1067 -1573
rect 1066 -1576 1249 -1575
rect 506 -1578 1249 -1577
rect 471 -1580 507 -1579
rect 184 -1582 472 -1581
rect 156 -1584 185 -1583
rect 156 -1586 804 -1585
rect 2 -1597 559 -1596
rect 569 -1597 850 -1596
rect 856 -1597 1067 -1596
rect 1094 -1597 1098 -1596
rect 1255 -1597 1259 -1596
rect 2 -1599 402 -1598
rect 415 -1599 570 -1598
rect 572 -1599 577 -1598
rect 632 -1599 664 -1598
rect 705 -1599 955 -1598
rect 1045 -1599 1347 -1598
rect 9 -1601 941 -1600
rect 954 -1601 1130 -1600
rect 1255 -1601 1284 -1600
rect 12 -1603 164 -1602
rect 177 -1603 213 -1602
rect 320 -1603 906 -1602
rect 940 -1603 1319 -1602
rect 51 -1605 584 -1604
rect 632 -1605 717 -1604
rect 754 -1605 1137 -1604
rect 1304 -1605 1319 -1604
rect 58 -1607 416 -1606
rect 485 -1607 640 -1606
rect 660 -1607 689 -1606
rect 716 -1607 738 -1606
rect 775 -1607 864 -1606
rect 884 -1607 906 -1606
rect 975 -1607 1137 -1606
rect 1304 -1607 1333 -1606
rect 58 -1609 514 -1608
rect 534 -1609 983 -1608
rect 1045 -1609 1109 -1608
rect 1129 -1609 1172 -1608
rect 65 -1611 552 -1610
rect 639 -1611 675 -1610
rect 688 -1611 766 -1610
rect 800 -1611 1200 -1610
rect 65 -1613 703 -1612
rect 765 -1613 780 -1612
rect 803 -1613 1109 -1612
rect 1199 -1613 1235 -1612
rect 79 -1615 801 -1614
rect 849 -1615 871 -1614
rect 884 -1615 899 -1614
rect 975 -1615 1053 -1614
rect 1094 -1615 1151 -1614
rect 1234 -1615 1326 -1614
rect 86 -1617 489 -1616
rect 495 -1617 549 -1616
rect 625 -1617 675 -1616
rect 779 -1617 815 -1616
rect 856 -1617 1329 -1616
rect 86 -1619 108 -1618
rect 110 -1619 577 -1618
rect 621 -1619 626 -1618
rect 660 -1619 1004 -1618
rect 1052 -1619 1123 -1618
rect 1220 -1619 1326 -1618
rect 40 -1621 1004 -1620
rect 1220 -1621 1277 -1620
rect 89 -1623 710 -1622
rect 814 -1623 843 -1622
rect 859 -1623 1060 -1622
rect 1258 -1623 1284 -1622
rect 100 -1625 1186 -1624
rect 1276 -1625 1354 -1624
rect 23 -1627 101 -1626
rect 107 -1627 584 -1626
rect 709 -1627 745 -1626
rect 842 -1627 878 -1626
rect 891 -1627 1263 -1626
rect 117 -1629 185 -1628
rect 194 -1629 381 -1628
rect 499 -1629 535 -1628
rect 537 -1629 703 -1628
rect 737 -1629 745 -1628
rect 863 -1629 920 -1628
rect 947 -1629 1186 -1628
rect 1262 -1629 1291 -1628
rect 138 -1631 472 -1630
rect 485 -1631 500 -1630
rect 506 -1631 524 -1630
rect 730 -1631 948 -1630
rect 982 -1631 1039 -1630
rect 1290 -1631 1312 -1630
rect 142 -1633 1102 -1632
rect 1311 -1633 1340 -1632
rect 47 -1635 143 -1634
rect 145 -1635 255 -1634
rect 338 -1635 458 -1634
rect 471 -1635 612 -1634
rect 730 -1635 748 -1634
rect 870 -1635 969 -1634
rect 996 -1635 1039 -1634
rect 1080 -1635 1102 -1634
rect 93 -1637 339 -1636
rect 352 -1637 458 -1636
rect 506 -1637 962 -1636
rect 968 -1637 990 -1636
rect 996 -1637 1165 -1636
rect 93 -1639 1207 -1638
rect 103 -1641 990 -1640
rect 1164 -1641 1214 -1640
rect 135 -1643 1214 -1642
rect 135 -1645 199 -1644
rect 212 -1645 248 -1644
rect 254 -1645 430 -1644
rect 443 -1645 612 -1644
rect 877 -1645 934 -1644
rect 961 -1645 1032 -1644
rect 1206 -1645 1228 -1644
rect 121 -1647 444 -1646
rect 460 -1647 934 -1646
rect 1031 -1647 1088 -1646
rect 1157 -1647 1228 -1646
rect 114 -1649 1088 -1648
rect 96 -1651 115 -1650
rect 121 -1651 241 -1650
rect 247 -1651 276 -1650
rect 352 -1651 493 -1650
rect 513 -1651 759 -1650
rect 894 -1651 1179 -1650
rect 152 -1653 283 -1652
rect 366 -1653 433 -1652
rect 492 -1653 528 -1652
rect 758 -1653 773 -1652
rect 1066 -1653 1179 -1652
rect 159 -1655 1060 -1654
rect 1073 -1655 1158 -1654
rect 163 -1657 832 -1656
rect 1024 -1657 1074 -1656
rect 177 -1659 752 -1658
rect 772 -1659 1116 -1658
rect 180 -1661 360 -1660
rect 366 -1661 563 -1660
rect 751 -1661 920 -1660
rect 1024 -1661 1242 -1660
rect 44 -1663 360 -1662
rect 373 -1663 430 -1662
rect 523 -1663 1172 -1662
rect 1241 -1663 1270 -1662
rect 44 -1665 55 -1664
rect 184 -1665 206 -1664
rect 240 -1665 297 -1664
rect 376 -1665 1018 -1664
rect 1115 -1665 1144 -1664
rect 54 -1667 80 -1666
rect 198 -1667 332 -1666
rect 380 -1667 423 -1666
rect 450 -1667 1018 -1666
rect 1143 -1667 1193 -1666
rect 51 -1669 1193 -1668
rect 205 -1671 405 -1670
rect 422 -1671 437 -1670
rect 450 -1671 696 -1670
rect 828 -1671 1270 -1670
rect 226 -1673 297 -1672
rect 324 -1673 829 -1672
rect 226 -1675 311 -1674
rect 324 -1675 388 -1674
rect 394 -1675 437 -1674
rect 527 -1675 542 -1674
rect 562 -1675 671 -1674
rect 695 -1675 902 -1674
rect 128 -1677 388 -1676
rect 394 -1677 598 -1676
rect 72 -1679 129 -1678
rect 275 -1679 290 -1678
rect 303 -1679 311 -1678
rect 331 -1679 521 -1678
rect 541 -1679 787 -1678
rect 72 -1681 262 -1680
rect 282 -1681 619 -1680
rect 786 -1681 822 -1680
rect 156 -1683 262 -1682
rect 404 -1683 461 -1682
rect 555 -1683 619 -1682
rect 821 -1683 899 -1682
rect 30 -1685 556 -1684
rect 590 -1685 598 -1684
rect 16 -1687 31 -1686
rect 170 -1687 304 -1686
rect 408 -1687 591 -1686
rect 170 -1689 269 -1688
rect 408 -1689 605 -1688
rect 149 -1691 269 -1690
rect 604 -1691 647 -1690
rect 149 -1693 913 -1692
rect 219 -1695 290 -1694
rect 520 -1695 913 -1694
rect 191 -1697 220 -1696
rect 646 -1697 682 -1696
rect 191 -1699 654 -1698
rect 681 -1699 724 -1698
rect 653 -1701 668 -1700
rect 723 -1701 794 -1700
rect 667 -1703 1298 -1702
rect 793 -1705 808 -1704
rect 1248 -1705 1298 -1704
rect 37 -1707 1249 -1706
rect 37 -1709 318 -1708
rect 807 -1709 836 -1708
rect 317 -1711 1081 -1710
rect 835 -1713 927 -1712
rect 926 -1715 1011 -1714
rect 373 -1717 1011 -1716
rect 9 -1728 111 -1727
rect 117 -1728 647 -1727
rect 667 -1728 934 -1727
rect 940 -1728 969 -1727
rect 1069 -1728 1242 -1727
rect 1318 -1728 1329 -1727
rect 16 -1730 31 -1729
rect 33 -1730 69 -1729
rect 72 -1730 374 -1729
rect 390 -1730 857 -1729
rect 898 -1730 1102 -1729
rect 1122 -1730 1277 -1729
rect 16 -1732 150 -1731
rect 152 -1732 1102 -1731
rect 1122 -1732 1172 -1731
rect 1227 -1732 1287 -1731
rect 9 -1734 153 -1733
rect 205 -1734 356 -1733
rect 359 -1734 647 -1733
rect 667 -1734 703 -1733
rect 712 -1734 766 -1733
rect 814 -1734 892 -1733
rect 898 -1734 976 -1733
rect 1171 -1734 1214 -1733
rect 1241 -1734 1291 -1733
rect 19 -1736 794 -1735
rect 835 -1736 857 -1735
rect 901 -1736 1277 -1735
rect 23 -1738 612 -1737
rect 702 -1738 724 -1737
rect 744 -1738 850 -1737
rect 933 -1738 948 -1737
rect 968 -1738 1046 -1737
rect 1213 -1738 1256 -1737
rect 26 -1740 101 -1739
rect 107 -1740 1018 -1739
rect 1255 -1740 1305 -1739
rect 26 -1742 983 -1741
rect 1010 -1742 1046 -1741
rect 30 -1744 269 -1743
rect 324 -1744 377 -1743
rect 404 -1744 535 -1743
rect 548 -1744 794 -1743
rect 835 -1744 871 -1743
rect 940 -1744 997 -1743
rect 1017 -1744 1074 -1743
rect 37 -1746 160 -1745
rect 205 -1746 311 -1745
rect 359 -1746 388 -1745
rect 457 -1746 1298 -1745
rect 44 -1748 241 -1747
rect 268 -1748 416 -1747
rect 457 -1748 552 -1747
rect 555 -1748 633 -1747
rect 719 -1748 885 -1747
rect 975 -1748 1032 -1747
rect 1073 -1748 1116 -1747
rect 44 -1750 1060 -1749
rect 1115 -1750 1165 -1749
rect 47 -1752 997 -1751
rect 1031 -1752 1095 -1751
rect 1164 -1752 1193 -1751
rect 54 -1754 1249 -1753
rect 72 -1756 94 -1755
rect 100 -1756 468 -1755
rect 485 -1756 1228 -1755
rect 1234 -1756 1249 -1755
rect 51 -1758 94 -1757
rect 107 -1758 290 -1757
rect 369 -1758 745 -1757
rect 747 -1758 822 -1757
rect 849 -1758 913 -1757
rect 1059 -1758 1109 -1757
rect 1192 -1758 1221 -1757
rect 1234 -1758 1284 -1757
rect 51 -1760 843 -1759
rect 912 -1760 990 -1759
rect 1108 -1760 1151 -1759
rect 1220 -1760 1270 -1759
rect 58 -1762 843 -1761
rect 989 -1762 1053 -1761
rect 1269 -1762 1312 -1761
rect 58 -1764 185 -1763
rect 226 -1764 524 -1763
rect 534 -1764 808 -1763
rect 821 -1764 927 -1763
rect 1052 -1764 1088 -1763
rect 2 -1766 227 -1765
rect 233 -1766 241 -1765
rect 275 -1766 325 -1765
rect 373 -1766 615 -1765
rect 625 -1766 808 -1765
rect 926 -1766 1004 -1765
rect 1087 -1766 1144 -1765
rect 2 -1768 55 -1767
rect 79 -1768 587 -1767
rect 604 -1768 948 -1767
rect 1143 -1768 1186 -1767
rect 79 -1770 87 -1769
rect 121 -1770 318 -1769
rect 401 -1770 1186 -1769
rect 86 -1772 300 -1771
rect 317 -1772 332 -1771
rect 401 -1772 423 -1771
rect 488 -1772 895 -1771
rect 114 -1774 122 -1773
rect 128 -1774 290 -1773
rect 331 -1774 346 -1773
rect 415 -1774 437 -1773
rect 506 -1774 643 -1773
rect 660 -1774 885 -1773
rect 128 -1776 262 -1775
rect 345 -1776 381 -1775
rect 436 -1776 472 -1775
rect 506 -1776 542 -1775
rect 555 -1776 773 -1775
rect 138 -1778 304 -1777
rect 464 -1778 472 -1777
rect 513 -1778 549 -1777
rect 576 -1778 1095 -1777
rect 142 -1780 1284 -1779
rect 142 -1782 482 -1781
rect 513 -1782 528 -1781
rect 541 -1782 563 -1781
rect 576 -1782 598 -1781
rect 611 -1782 689 -1781
rect 723 -1782 776 -1781
rect 149 -1784 591 -1783
rect 597 -1784 640 -1783
rect 660 -1784 682 -1783
rect 730 -1784 1011 -1783
rect 156 -1786 591 -1785
rect 625 -1786 864 -1785
rect 156 -1788 171 -1787
rect 177 -1788 682 -1787
rect 730 -1788 920 -1787
rect 96 -1790 920 -1789
rect 163 -1792 381 -1791
rect 408 -1792 528 -1791
rect 562 -1792 619 -1791
rect 628 -1792 1004 -1791
rect 170 -1794 283 -1793
rect 394 -1794 409 -1793
rect 464 -1794 983 -1793
rect 177 -1796 297 -1795
rect 394 -1796 461 -1795
rect 520 -1796 1207 -1795
rect 184 -1798 220 -1797
rect 233 -1798 451 -1797
rect 520 -1798 944 -1797
rect 65 -1800 220 -1799
rect 247 -1800 276 -1799
rect 282 -1800 500 -1799
rect 569 -1800 689 -1799
rect 733 -1800 773 -1799
rect 863 -1800 955 -1799
rect 40 -1802 66 -1801
rect 191 -1802 1207 -1801
rect 114 -1804 192 -1803
rect 198 -1804 304 -1803
rect 338 -1804 451 -1803
rect 569 -1804 696 -1803
rect 737 -1804 871 -1803
rect 135 -1806 199 -1805
rect 247 -1806 255 -1805
rect 261 -1806 493 -1805
rect 583 -1806 955 -1805
rect 135 -1808 164 -1807
rect 254 -1808 388 -1807
rect 443 -1808 500 -1807
rect 583 -1808 759 -1807
rect 761 -1808 878 -1807
rect 296 -1810 717 -1809
rect 751 -1810 1158 -1809
rect 310 -1812 759 -1811
rect 765 -1812 801 -1811
rect 877 -1812 906 -1811
rect 1024 -1812 1158 -1811
rect 338 -1814 353 -1813
rect 366 -1814 493 -1813
rect 618 -1814 654 -1813
rect 674 -1814 801 -1813
rect 905 -1814 962 -1813
rect 1024 -1814 1081 -1813
rect 320 -1816 675 -1815
rect 695 -1816 710 -1815
rect 716 -1816 1151 -1815
rect 352 -1818 755 -1817
rect 961 -1818 1039 -1817
rect 1080 -1818 1137 -1817
rect 366 -1820 430 -1819
rect 443 -1820 605 -1819
rect 607 -1820 1137 -1819
rect 23 -1822 430 -1821
rect 485 -1822 755 -1821
rect 1038 -1822 1067 -1821
rect 422 -1824 710 -1823
rect 737 -1824 752 -1823
rect 1066 -1824 1130 -1823
rect 632 -1826 780 -1825
rect 1129 -1826 1179 -1825
rect 639 -1828 1126 -1827
rect 1178 -1828 1200 -1827
rect 653 -1830 815 -1829
rect 1199 -1830 1263 -1829
rect 558 -1832 1263 -1831
rect 779 -1834 787 -1833
rect 194 -1836 787 -1835
rect 2 -1847 524 -1846
rect 604 -1847 647 -1846
rect 653 -1847 696 -1846
rect 712 -1847 878 -1846
rect 16 -1849 388 -1848
rect 432 -1849 1011 -1848
rect 9 -1851 17 -1850
rect 23 -1851 31 -1850
rect 37 -1851 1179 -1850
rect 9 -1853 80 -1852
rect 89 -1853 248 -1852
rect 254 -1853 367 -1852
rect 387 -1853 556 -1852
rect 558 -1853 654 -1852
rect 656 -1853 892 -1852
rect 1178 -1853 1270 -1852
rect 23 -1855 94 -1854
rect 103 -1855 1095 -1854
rect 30 -1857 521 -1856
rect 555 -1857 1053 -1856
rect 1094 -1857 1242 -1856
rect 37 -1859 339 -1858
rect 366 -1859 437 -1858
rect 464 -1859 507 -1858
rect 513 -1859 542 -1858
rect 607 -1859 857 -1858
rect 877 -1859 997 -1858
rect 1052 -1859 1158 -1858
rect 40 -1861 290 -1860
rect 296 -1861 468 -1860
rect 478 -1861 633 -1860
rect 639 -1861 766 -1860
rect 856 -1861 1060 -1860
rect 1157 -1861 1235 -1860
rect 44 -1863 1004 -1862
rect 1115 -1863 1235 -1862
rect 44 -1865 97 -1864
rect 114 -1865 234 -1864
rect 254 -1865 325 -1864
rect 408 -1865 465 -1864
rect 471 -1865 479 -1864
rect 492 -1865 706 -1864
rect 719 -1865 948 -1864
rect 996 -1865 1081 -1864
rect 1115 -1865 1200 -1864
rect 47 -1867 920 -1866
rect 933 -1867 1060 -1866
rect 1080 -1867 1193 -1866
rect 79 -1869 416 -1868
rect 429 -1869 640 -1868
rect 646 -1869 927 -1868
rect 933 -1869 1032 -1868
rect 1143 -1869 1200 -1868
rect 93 -1871 101 -1870
rect 114 -1871 563 -1870
rect 597 -1871 608 -1870
rect 614 -1871 843 -1870
rect 891 -1871 923 -1870
rect 926 -1871 1186 -1870
rect 100 -1873 528 -1872
rect 534 -1873 563 -1872
rect 597 -1873 619 -1872
rect 628 -1873 1032 -1872
rect 1038 -1873 1186 -1872
rect 135 -1875 808 -1874
rect 842 -1875 969 -1874
rect 1164 -1875 1193 -1874
rect 135 -1877 1144 -1876
rect 149 -1879 234 -1878
rect 264 -1879 283 -1878
rect 289 -1879 311 -1878
rect 324 -1879 395 -1878
rect 408 -1879 675 -1878
rect 677 -1879 689 -1878
rect 695 -1879 787 -1878
rect 919 -1879 1011 -1878
rect 1073 -1879 1165 -1878
rect 86 -1881 283 -1880
rect 299 -1881 573 -1880
rect 688 -1881 773 -1880
rect 786 -1881 899 -1880
rect 947 -1881 1102 -1880
rect 86 -1883 1228 -1882
rect 149 -1885 199 -1884
rect 226 -1885 626 -1884
rect 730 -1885 829 -1884
rect 863 -1885 1102 -1884
rect 152 -1887 269 -1886
rect 275 -1887 416 -1886
rect 436 -1887 451 -1886
rect 457 -1887 626 -1886
rect 709 -1887 829 -1886
rect 863 -1887 962 -1886
rect 968 -1887 1109 -1886
rect 163 -1889 297 -1888
rect 303 -1889 311 -1888
rect 352 -1889 962 -1888
rect 1073 -1889 1256 -1888
rect 163 -1891 356 -1890
rect 422 -1891 451 -1890
rect 471 -1891 839 -1890
rect 898 -1891 1088 -1890
rect 177 -1893 269 -1892
rect 275 -1893 1224 -1892
rect 177 -1895 213 -1894
rect 285 -1895 1109 -1894
rect 184 -1897 227 -1896
rect 303 -1897 521 -1896
rect 527 -1897 577 -1896
rect 709 -1897 745 -1896
rect 751 -1897 976 -1896
rect 1066 -1897 1088 -1896
rect 128 -1899 185 -1898
rect 198 -1899 206 -1898
rect 212 -1899 220 -1898
rect 345 -1899 353 -1898
rect 380 -1899 423 -1898
rect 443 -1899 619 -1898
rect 737 -1899 808 -1898
rect 912 -1899 1228 -1898
rect 128 -1901 143 -1900
rect 205 -1901 241 -1900
rect 345 -1901 402 -1900
rect 495 -1901 794 -1900
rect 912 -1901 1046 -1900
rect 1066 -1901 1172 -1900
rect 51 -1903 402 -1902
rect 506 -1903 724 -1902
rect 737 -1903 850 -1902
rect 975 -1903 1137 -1902
rect 1171 -1903 1263 -1902
rect 51 -1905 458 -1904
rect 516 -1905 1004 -1904
rect 1045 -1905 1151 -1904
rect 58 -1907 143 -1906
rect 219 -1907 318 -1906
rect 359 -1907 444 -1906
rect 534 -1907 591 -1906
rect 744 -1907 836 -1906
rect 849 -1907 1025 -1906
rect 1150 -1907 1249 -1906
rect 58 -1909 500 -1908
rect 541 -1909 668 -1908
rect 751 -1909 762 -1908
rect 765 -1909 885 -1908
rect 1024 -1909 1130 -1908
rect 65 -1911 794 -1910
rect 835 -1911 1214 -1910
rect 138 -1913 724 -1912
rect 754 -1913 941 -1912
rect 1213 -1913 1277 -1912
rect 138 -1915 157 -1914
rect 191 -1915 500 -1914
rect 548 -1915 633 -1914
rect 667 -1915 703 -1914
rect 758 -1915 780 -1914
rect 156 -1917 482 -1916
rect 548 -1917 643 -1916
rect 702 -1917 1039 -1916
rect 191 -1919 370 -1918
rect 380 -1919 605 -1918
rect 761 -1919 885 -1918
rect 72 -1921 370 -1920
rect 429 -1921 1137 -1920
rect 68 -1923 73 -1922
rect 240 -1923 262 -1922
rect 317 -1923 339 -1922
rect 359 -1923 584 -1922
rect 590 -1923 661 -1922
rect 772 -1923 990 -1922
rect 54 -1925 69 -1924
rect 107 -1925 262 -1924
rect 320 -1925 661 -1924
rect 779 -1925 822 -1924
rect 107 -1927 122 -1926
rect 247 -1927 759 -1926
rect 821 -1927 955 -1926
rect 121 -1929 171 -1928
rect 460 -1929 1130 -1928
rect 170 -1931 395 -1930
rect 492 -1931 990 -1930
rect 569 -1933 584 -1932
rect 954 -1933 1221 -1932
rect 569 -1935 941 -1934
rect 576 -1937 815 -1936
rect 814 -1939 871 -1938
rect 870 -1941 983 -1940
rect 611 -1943 983 -1942
rect 611 -1945 682 -1944
rect 681 -1947 717 -1946
rect 716 -1949 801 -1948
rect 800 -1951 906 -1950
rect 905 -1953 1018 -1952
rect 1017 -1955 1123 -1954
rect 1122 -1957 1207 -1956
rect 586 -1959 1207 -1958
rect 2 -1970 647 -1969
rect 674 -1970 955 -1969
rect 964 -1970 1095 -1969
rect 1164 -1970 1221 -1969
rect 9 -1972 136 -1971
rect 142 -1972 286 -1971
rect 310 -1972 318 -1971
rect 320 -1972 332 -1971
rect 373 -1972 377 -1971
rect 401 -1972 675 -1971
rect 702 -1972 1102 -1971
rect 9 -1974 167 -1973
rect 184 -1974 493 -1973
rect 499 -1974 622 -1973
rect 702 -1974 738 -1973
rect 758 -1974 1088 -1973
rect 1094 -1974 1137 -1973
rect 16 -1976 262 -1975
rect 282 -1976 458 -1975
rect 464 -1976 493 -1975
rect 499 -1976 1214 -1975
rect 37 -1978 174 -1977
rect 184 -1978 325 -1977
rect 331 -1978 395 -1977
rect 408 -1978 412 -1977
rect 464 -1978 542 -1977
rect 569 -1978 717 -1977
rect 737 -1978 892 -1977
rect 919 -1978 997 -1977
rect 1027 -1978 1193 -1977
rect 37 -1980 164 -1979
rect 191 -1980 370 -1979
rect 373 -1980 381 -1979
rect 394 -1980 689 -1979
rect 716 -1980 801 -1979
rect 891 -1980 934 -1979
rect 954 -1980 962 -1979
rect 968 -1980 972 -1979
rect 996 -1980 1123 -1979
rect 16 -1982 164 -1981
rect 198 -1982 430 -1981
rect 481 -1982 1011 -1981
rect 1073 -1982 1123 -1981
rect 51 -1984 241 -1983
rect 243 -1984 689 -1983
rect 758 -1984 787 -1983
rect 800 -1984 843 -1983
rect 919 -1984 941 -1983
rect 968 -1984 976 -1983
rect 1010 -1984 1144 -1983
rect 54 -1986 745 -1985
rect 761 -1986 990 -1985
rect 1059 -1986 1144 -1985
rect 58 -1988 458 -1987
rect 488 -1988 773 -1987
rect 786 -1988 871 -1987
rect 940 -1988 948 -1987
rect 982 -1988 1060 -1987
rect 1073 -1988 1109 -1987
rect 58 -1990 367 -1989
rect 408 -1990 416 -1989
rect 429 -1990 479 -1989
rect 502 -1990 647 -1989
rect 677 -1990 962 -1989
rect 982 -1990 1046 -1989
rect 1087 -1990 1228 -1989
rect 65 -1992 97 -1991
rect 100 -1992 290 -1991
rect 310 -1992 598 -1991
rect 604 -1992 1200 -1991
rect 23 -1994 97 -1993
rect 110 -1994 486 -1993
rect 513 -1994 559 -1993
rect 569 -1994 612 -1993
rect 744 -1994 836 -1993
rect 842 -1994 1018 -1993
rect 1101 -1994 1172 -1993
rect 23 -1996 507 -1995
rect 520 -1996 899 -1995
rect 947 -1996 1004 -1995
rect 1017 -1996 1067 -1995
rect 1108 -1996 1179 -1995
rect 44 -1998 66 -1997
rect 68 -1998 731 -1997
rect 772 -1998 839 -1997
rect 849 -1998 871 -1997
rect 898 -1998 1039 -1997
rect 1066 -1998 1081 -1997
rect 72 -2000 664 -1999
rect 835 -2000 878 -1999
rect 971 -2000 976 -1999
rect 989 -2000 1025 -1999
rect 1031 -2000 1039 -1999
rect 1080 -2000 1116 -1999
rect 72 -2002 108 -2001
rect 114 -2002 367 -2001
rect 478 -2002 731 -2001
rect 877 -2002 885 -2001
rect 1003 -2002 1053 -2001
rect 1115 -2002 1207 -2001
rect 86 -2004 136 -2003
rect 142 -2004 269 -2003
rect 282 -2004 451 -2003
rect 506 -2004 699 -2003
rect 926 -2004 1053 -2003
rect 86 -2006 563 -2005
rect 576 -2006 885 -2005
rect 1031 -2006 1151 -2005
rect 44 -2008 577 -2007
rect 579 -2008 815 -2007
rect 856 -2008 927 -2007
rect 1136 -2008 1151 -2007
rect 51 -2010 815 -2009
rect 856 -2010 906 -2009
rect 89 -2012 108 -2011
rect 117 -2012 213 -2011
rect 226 -2012 279 -2011
rect 317 -2012 346 -2011
rect 450 -2012 472 -2011
rect 534 -2012 934 -2011
rect 93 -2014 710 -2013
rect 905 -2014 913 -2013
rect 93 -2016 304 -2015
rect 338 -2016 605 -2015
rect 611 -2016 626 -2015
rect 709 -2016 766 -2015
rect 30 -2018 304 -2017
rect 471 -2018 549 -2017
rect 562 -2018 682 -2017
rect 751 -2018 913 -2017
rect 30 -2020 360 -2019
rect 534 -2020 591 -2019
rect 597 -2020 633 -2019
rect 681 -2020 696 -2019
rect 751 -2020 780 -2019
rect 114 -2022 339 -2021
rect 432 -2022 591 -2021
rect 625 -2022 661 -2021
rect 765 -2022 822 -2021
rect 121 -2024 521 -2023
rect 541 -2024 584 -2023
rect 632 -2024 640 -2023
rect 660 -2024 668 -2023
rect 821 -2024 864 -2023
rect 103 -2026 668 -2025
rect 863 -2026 1186 -2025
rect 121 -2028 654 -2027
rect 1185 -2028 1235 -2027
rect 128 -2030 573 -2029
rect 583 -2030 780 -2029
rect 152 -2032 850 -2031
rect 170 -2034 346 -2033
rect 548 -2034 619 -2033
rect 639 -2034 1025 -2033
rect 149 -2036 171 -2035
rect 177 -2036 213 -2035
rect 226 -2036 276 -2035
rect 618 -2036 1046 -2035
rect 128 -2038 150 -2037
rect 177 -2038 696 -2037
rect 191 -2040 241 -2039
rect 247 -2040 514 -2039
rect 653 -2040 808 -2039
rect 198 -2042 388 -2041
rect 807 -2042 829 -2041
rect 205 -2044 262 -2043
rect 268 -2044 353 -2043
rect 828 -2044 1130 -2043
rect 156 -2046 206 -2045
rect 233 -2046 360 -2045
rect 723 -2046 1130 -2045
rect 79 -2048 157 -2047
rect 233 -2048 524 -2047
rect 723 -2048 794 -2047
rect 79 -2050 335 -2049
rect 352 -2050 423 -2049
rect 555 -2050 794 -2049
rect 247 -2052 461 -2051
rect 555 -2052 1224 -2051
rect 254 -2054 290 -2053
rect 296 -2054 388 -2053
rect 422 -2054 528 -2053
rect 138 -2056 297 -2055
rect 436 -2056 528 -2055
rect 219 -2058 255 -2057
rect 275 -2058 402 -2057
rect 436 -2058 444 -2057
rect 89 -2060 444 -2059
rect 219 -2062 608 -2061
rect 2 -2073 94 -2072
rect 103 -2073 745 -2072
rect 789 -2073 1123 -2072
rect 1136 -2073 1186 -2072
rect 30 -2075 244 -2074
rect 247 -2075 279 -2074
rect 394 -2075 619 -2074
rect 621 -2075 801 -2074
rect 817 -2075 976 -2074
rect 1122 -2075 1151 -2074
rect 30 -2077 87 -2076
rect 93 -2077 164 -2076
rect 166 -2077 997 -2076
rect 1139 -2077 1158 -2076
rect 37 -2079 325 -2078
rect 394 -2079 472 -2078
rect 481 -2079 528 -2078
rect 562 -2079 566 -2078
rect 576 -2079 878 -2078
rect 975 -2079 1039 -2078
rect 65 -2081 153 -2080
rect 156 -2081 500 -2080
rect 509 -2081 640 -2080
rect 653 -2081 1025 -2080
rect 65 -2083 297 -2082
rect 387 -2083 482 -2082
rect 492 -2083 531 -2082
rect 562 -2083 591 -2082
rect 600 -2083 633 -2082
rect 639 -2083 885 -2082
rect 86 -2085 136 -2084
rect 138 -2085 794 -2084
rect 863 -2085 1088 -2084
rect 37 -2087 136 -2086
rect 142 -2087 489 -2086
rect 565 -2087 591 -2086
rect 614 -2087 997 -2086
rect 100 -2089 248 -2088
rect 254 -2089 300 -2088
rect 387 -2089 451 -2088
rect 457 -2089 500 -2088
rect 576 -2089 626 -2088
rect 632 -2089 668 -2088
rect 695 -2089 759 -2088
rect 793 -2089 1130 -2088
rect 100 -2091 164 -2090
rect 170 -2091 241 -2090
rect 254 -2091 290 -2090
rect 401 -2091 493 -2090
rect 579 -2091 612 -2090
rect 618 -2091 675 -2090
rect 695 -2091 948 -2090
rect 107 -2093 115 -2092
rect 117 -2093 283 -2092
rect 289 -2093 304 -2092
rect 401 -2093 465 -2092
rect 467 -2093 1039 -2092
rect 58 -2095 108 -2094
rect 114 -2095 381 -2094
rect 429 -2095 451 -2094
rect 457 -2095 647 -2094
rect 656 -2095 710 -2094
rect 716 -2095 801 -2094
rect 863 -2095 927 -2094
rect 947 -2095 1102 -2094
rect 23 -2097 59 -2096
rect 142 -2097 234 -2096
rect 240 -2097 335 -2096
rect 373 -2097 381 -2096
rect 408 -2097 647 -2096
rect 660 -2097 843 -2096
rect 877 -2097 955 -2096
rect 23 -2099 90 -2098
rect 96 -2099 374 -2098
rect 429 -2099 437 -2098
rect 443 -2099 612 -2098
rect 625 -2099 689 -2098
rect 709 -2099 808 -2098
rect 842 -2099 892 -2098
rect 926 -2099 983 -2098
rect 149 -2101 486 -2100
rect 583 -2101 913 -2100
rect 933 -2101 955 -2100
rect 982 -2101 1067 -2100
rect 44 -2103 150 -2102
rect 156 -2103 220 -2102
rect 233 -2103 318 -2102
rect 345 -2103 409 -2102
rect 443 -2103 692 -2102
rect 716 -2103 773 -2102
rect 807 -2103 822 -2102
rect 884 -2103 962 -2102
rect 1066 -2103 1081 -2102
rect 44 -2105 699 -2104
rect 737 -2105 759 -2104
rect 772 -2105 787 -2104
rect 821 -2105 906 -2104
rect 933 -2105 1018 -2104
rect 51 -2107 220 -2106
rect 261 -2107 321 -2106
rect 338 -2107 962 -2106
rect 1017 -2107 1116 -2106
rect 16 -2109 52 -2108
rect 173 -2109 682 -2108
rect 737 -2109 766 -2108
rect 891 -2109 969 -2108
rect 110 -2111 766 -2110
rect 898 -2111 913 -2110
rect 968 -2111 1032 -2110
rect 184 -2113 283 -2112
rect 303 -2113 517 -2112
rect 583 -2113 598 -2112
rect 660 -2113 664 -2112
rect 667 -2113 703 -2112
rect 744 -2113 752 -2112
rect 814 -2113 899 -2112
rect 905 -2113 1060 -2112
rect 184 -2115 535 -2114
rect 674 -2115 724 -2114
rect 751 -2115 780 -2114
rect 814 -2115 857 -2114
rect 866 -2115 1060 -2114
rect 205 -2117 325 -2116
rect 338 -2117 503 -2116
rect 681 -2117 850 -2116
rect 856 -2117 1004 -2116
rect 1031 -2117 1105 -2116
rect 205 -2119 227 -2118
rect 261 -2119 528 -2118
rect 702 -2119 871 -2118
rect 1003 -2119 1144 -2118
rect 79 -2121 227 -2120
rect 268 -2121 332 -2120
rect 345 -2121 423 -2120
rect 471 -2121 549 -2120
rect 723 -2121 836 -2120
rect 849 -2121 1053 -2120
rect 79 -2123 479 -2122
rect 548 -2123 643 -2122
rect 730 -2123 780 -2122
rect 835 -2123 1046 -2122
rect 1052 -2123 1102 -2122
rect 128 -2125 332 -2124
rect 352 -2125 437 -2124
rect 478 -2125 990 -2124
rect 128 -2127 178 -2126
rect 212 -2127 328 -2126
rect 352 -2127 514 -2126
rect 597 -2127 1046 -2126
rect 9 -2129 514 -2128
rect 730 -2129 829 -2128
rect 870 -2129 941 -2128
rect 989 -2129 1074 -2128
rect 177 -2131 192 -2130
rect 212 -2131 360 -2130
rect 366 -2131 423 -2130
rect 485 -2131 941 -2130
rect 121 -2133 192 -2132
rect 268 -2133 507 -2132
rect 828 -2133 920 -2132
rect 117 -2135 122 -2134
rect 275 -2135 556 -2134
rect 919 -2135 1095 -2134
rect 310 -2137 535 -2136
rect 555 -2137 570 -2136
rect 198 -2139 311 -2138
rect 359 -2139 416 -2138
rect 464 -2139 570 -2138
rect 198 -2141 318 -2140
rect 366 -2141 521 -2140
rect 415 -2143 605 -2142
rect 520 -2145 542 -2144
rect 604 -2145 689 -2144
rect 541 -2147 787 -2146
rect 23 -2158 118 -2157
rect 124 -2158 304 -2157
rect 317 -2158 325 -2157
rect 331 -2158 972 -2157
rect 975 -2158 997 -2157
rect 1101 -2158 1109 -2157
rect 37 -2160 101 -2159
rect 103 -2160 157 -2159
rect 198 -2160 304 -2159
rect 324 -2160 381 -2159
rect 387 -2160 489 -2159
rect 509 -2160 850 -2159
rect 933 -2160 969 -2159
rect 982 -2160 997 -2159
rect 1104 -2160 1123 -2159
rect 37 -2162 87 -2161
rect 93 -2162 262 -2161
rect 275 -2162 465 -2161
rect 485 -2162 584 -2161
rect 597 -2162 703 -2161
rect 786 -2162 899 -2161
rect 933 -2162 1039 -2161
rect 30 -2164 94 -2163
rect 100 -2164 143 -2163
rect 198 -2164 248 -2163
rect 254 -2164 468 -2163
rect 513 -2164 696 -2163
rect 702 -2164 738 -2163
rect 786 -2164 885 -2163
rect 943 -2164 1060 -2163
rect 30 -2166 528 -2165
rect 597 -2166 633 -2165
rect 639 -2166 675 -2165
rect 688 -2166 920 -2165
rect 982 -2166 1004 -2165
rect 51 -2168 157 -2167
rect 233 -2168 479 -2167
rect 513 -2168 542 -2167
rect 611 -2168 955 -2167
rect 1003 -2168 1053 -2167
rect 44 -2170 52 -2169
rect 65 -2170 262 -2169
rect 289 -2170 489 -2169
rect 541 -2170 570 -2169
rect 611 -2170 699 -2169
rect 842 -2170 976 -2169
rect 58 -2172 66 -2171
rect 72 -2172 136 -2171
rect 138 -2172 584 -2171
rect 614 -2172 899 -2171
rect 919 -2172 1032 -2171
rect 58 -2174 398 -2173
rect 408 -2174 482 -2173
rect 632 -2174 710 -2173
rect 842 -2174 962 -2173
rect 72 -2176 185 -2175
rect 240 -2176 248 -2175
rect 254 -2176 269 -2175
rect 289 -2176 395 -2175
rect 401 -2176 409 -2175
rect 429 -2176 507 -2175
rect 646 -2176 885 -2175
rect 96 -2178 185 -2177
rect 205 -2178 241 -2177
rect 268 -2178 790 -2177
rect 96 -2180 657 -2179
rect 674 -2180 682 -2179
rect 688 -2180 766 -2179
rect 114 -2182 276 -2181
rect 296 -2182 332 -2181
rect 355 -2182 605 -2181
rect 646 -2182 668 -2181
rect 681 -2182 759 -2181
rect 114 -2184 122 -2183
rect 131 -2184 360 -2183
rect 366 -2184 395 -2183
rect 401 -2184 451 -2183
rect 464 -2184 500 -2183
rect 506 -2184 556 -2183
rect 604 -2184 748 -2183
rect 751 -2184 962 -2183
rect 121 -2186 444 -2185
rect 457 -2186 556 -2185
rect 656 -2186 857 -2185
rect 135 -2188 220 -2187
rect 282 -2188 297 -2187
rect 310 -2188 367 -2187
rect 373 -2188 430 -2187
rect 443 -2188 493 -2187
rect 499 -2188 531 -2187
rect 691 -2188 801 -2187
rect 856 -2188 906 -2187
rect 79 -2190 283 -2189
rect 310 -2190 353 -2189
rect 359 -2190 549 -2189
rect 695 -2190 1046 -2189
rect 79 -2192 129 -2191
rect 142 -2192 150 -2191
rect 163 -2192 570 -2191
rect 709 -2192 780 -2191
rect 800 -2192 808 -2191
rect 905 -2192 1025 -2191
rect 44 -2194 129 -2193
rect 163 -2194 654 -2193
rect 751 -2194 871 -2193
rect 86 -2196 150 -2195
rect 170 -2196 234 -2195
rect 320 -2196 850 -2195
rect 870 -2196 1018 -2195
rect 170 -2198 178 -2197
rect 180 -2198 493 -2197
rect 548 -2198 591 -2197
rect 653 -2198 773 -2197
rect 779 -2198 822 -2197
rect 954 -2198 1018 -2197
rect 177 -2200 213 -2199
rect 219 -2200 346 -2199
rect 373 -2200 472 -2199
rect 590 -2200 626 -2199
rect 758 -2200 878 -2199
rect 107 -2202 346 -2201
rect 380 -2202 577 -2201
rect 618 -2202 626 -2201
rect 772 -2202 829 -2201
rect 877 -2202 948 -2201
rect 107 -2204 300 -2203
rect 387 -2204 437 -2203
rect 450 -2204 577 -2203
rect 618 -2204 794 -2203
rect 807 -2204 815 -2203
rect 821 -2204 892 -2203
rect 191 -2206 668 -2205
rect 670 -2206 892 -2205
rect 191 -2208 563 -2207
rect 793 -2208 836 -2207
rect 205 -2210 661 -2209
rect 814 -2210 913 -2209
rect 212 -2212 454 -2211
rect 471 -2212 521 -2211
rect 660 -2212 717 -2211
rect 828 -2212 941 -2211
rect 338 -2214 717 -2213
rect 765 -2214 941 -2213
rect 338 -2216 741 -2215
rect 835 -2216 927 -2215
rect 422 -2218 458 -2217
rect 485 -2218 948 -2217
rect 415 -2220 423 -2219
rect 436 -2220 724 -2219
rect 912 -2220 990 -2219
rect 415 -2222 528 -2221
rect 723 -2222 864 -2221
rect 926 -2222 1011 -2221
rect 516 -2224 563 -2223
rect 730 -2224 864 -2223
rect 520 -2226 535 -2225
rect 730 -2226 745 -2225
rect 534 -2228 601 -2227
rect 30 -2239 129 -2238
rect 131 -2239 339 -2238
rect 345 -2239 349 -2238
rect 359 -2239 657 -2238
rect 667 -2239 836 -2238
rect 940 -2239 962 -2238
rect 989 -2239 1004 -2238
rect 1017 -2239 1039 -2238
rect 1059 -2239 1067 -2238
rect 44 -2241 48 -2240
rect 51 -2241 90 -2240
rect 93 -2241 451 -2240
rect 481 -2241 633 -2240
rect 667 -2241 689 -2240
rect 695 -2241 752 -2240
rect 800 -2241 804 -2240
rect 807 -2241 811 -2240
rect 835 -2241 871 -2240
rect 943 -2241 983 -2240
rect 37 -2243 90 -2242
rect 135 -2243 339 -2242
rect 359 -2243 374 -2242
rect 429 -2243 479 -2242
rect 527 -2243 661 -2242
rect 674 -2243 678 -2242
rect 681 -2243 685 -2242
rect 688 -2243 766 -2242
rect 800 -2243 927 -2242
rect 957 -2243 976 -2242
rect 44 -2245 59 -2244
rect 65 -2245 129 -2244
rect 135 -2245 157 -2244
rect 177 -2245 241 -2244
rect 261 -2245 356 -2244
rect 429 -2245 507 -2244
rect 527 -2245 549 -2244
rect 583 -2245 587 -2244
rect 632 -2245 647 -2244
rect 674 -2245 759 -2244
rect 765 -2245 815 -2244
rect 870 -2245 955 -2244
rect 51 -2247 115 -2246
rect 138 -2247 566 -2246
rect 583 -2247 598 -2246
rect 621 -2247 647 -2246
rect 681 -2247 717 -2246
rect 723 -2247 759 -2246
rect 807 -2247 843 -2246
rect 65 -2249 101 -2248
rect 114 -2249 143 -2248
rect 170 -2249 178 -2248
rect 180 -2249 241 -2248
rect 247 -2249 262 -2248
rect 303 -2249 353 -2248
rect 436 -2249 454 -2248
rect 478 -2249 573 -2248
rect 639 -2249 661 -2248
rect 698 -2249 913 -2248
rect 72 -2251 531 -2250
rect 534 -2251 549 -2250
rect 611 -2251 640 -2250
rect 702 -2251 717 -2250
rect 730 -2251 745 -2250
rect 747 -2251 885 -2250
rect 72 -2253 164 -2252
rect 184 -2253 395 -2252
rect 408 -2253 437 -2252
rect 446 -2253 458 -2252
rect 499 -2253 507 -2252
rect 604 -2253 612 -2252
rect 656 -2253 885 -2252
rect 79 -2255 213 -2254
rect 226 -2255 654 -2254
rect 709 -2255 724 -2254
rect 730 -2255 773 -2254
rect 814 -2255 864 -2254
rect 96 -2257 227 -2256
rect 247 -2257 388 -2256
rect 408 -2257 542 -2256
rect 576 -2257 605 -2256
rect 737 -2257 752 -2256
rect 772 -2257 780 -2256
rect 842 -2257 892 -2256
rect 100 -2259 290 -2258
rect 303 -2259 377 -2258
rect 387 -2259 538 -2258
rect 737 -2259 787 -2258
rect 810 -2259 892 -2258
rect 107 -2261 143 -2260
rect 156 -2261 447 -2260
rect 471 -2261 500 -2260
rect 740 -2261 857 -2260
rect 863 -2261 948 -2260
rect 107 -2263 192 -2262
rect 198 -2263 293 -2262
rect 310 -2263 353 -2262
rect 366 -2263 395 -2262
rect 492 -2263 542 -2262
rect 744 -2263 794 -2262
rect 856 -2263 920 -2262
rect 124 -2265 171 -2264
rect 198 -2265 269 -2264
rect 275 -2265 454 -2264
rect 779 -2265 822 -2264
rect 149 -2267 192 -2266
rect 212 -2267 234 -2266
rect 254 -2267 535 -2266
rect 653 -2267 822 -2266
rect 149 -2269 188 -2268
rect 219 -2269 577 -2268
rect 786 -2269 829 -2268
rect 163 -2271 398 -2270
rect 793 -2271 906 -2270
rect 184 -2273 255 -2272
rect 268 -2273 486 -2272
rect 828 -2273 850 -2272
rect 219 -2275 374 -2274
rect 443 -2275 486 -2274
rect 849 -2275 899 -2274
rect 93 -2277 444 -2276
rect 877 -2277 899 -2276
rect 233 -2279 297 -2278
rect 310 -2279 381 -2278
rect 877 -2279 934 -2278
rect 275 -2281 283 -2280
rect 296 -2281 493 -2280
rect 282 -2283 318 -2282
rect 324 -2283 381 -2282
rect 317 -2285 580 -2284
rect 324 -2287 402 -2286
rect 345 -2289 458 -2288
rect 366 -2291 416 -2290
rect 121 -2293 416 -2292
rect 121 -2295 514 -2294
rect 401 -2297 556 -2296
rect 422 -2299 514 -2298
rect 555 -2299 570 -2298
rect 422 -2301 626 -2300
rect 464 -2303 570 -2302
rect 590 -2303 626 -2302
rect 464 -2305 671 -2304
rect 590 -2307 619 -2306
rect 562 -2309 619 -2308
rect 471 -2311 563 -2310
rect 51 -2322 185 -2321
rect 187 -2322 377 -2321
rect 383 -2322 472 -2321
rect 492 -2322 794 -2321
rect 884 -2322 941 -2321
rect 968 -2322 979 -2321
rect 982 -2322 990 -2321
rect 996 -2322 1004 -2321
rect 1038 -2322 1060 -2321
rect 65 -2324 87 -2323
rect 89 -2324 752 -2323
rect 772 -2324 801 -2323
rect 898 -2324 906 -2323
rect 989 -2324 1007 -2323
rect 44 -2326 87 -2325
rect 135 -2326 283 -2325
rect 306 -2326 472 -2325
rect 492 -2326 622 -2325
rect 632 -2326 657 -2325
rect 698 -2326 871 -2325
rect 891 -2326 899 -2325
rect 138 -2328 297 -2327
rect 310 -2328 451 -2327
rect 457 -2328 804 -2327
rect 152 -2330 262 -2329
rect 275 -2330 496 -2329
rect 558 -2330 829 -2329
rect 114 -2332 262 -2331
rect 292 -2332 297 -2331
rect 338 -2332 349 -2331
rect 352 -2332 444 -2331
rect 446 -2332 710 -2331
rect 716 -2332 720 -2331
rect 751 -2332 836 -2331
rect 114 -2334 185 -2333
rect 205 -2334 276 -2333
rect 338 -2334 367 -2333
rect 387 -2334 531 -2333
rect 548 -2334 710 -2333
rect 716 -2334 815 -2333
rect 93 -2336 206 -2335
rect 233 -2336 283 -2335
rect 359 -2336 374 -2335
rect 387 -2336 423 -2335
rect 429 -2336 535 -2335
rect 562 -2336 703 -2335
rect 772 -2336 864 -2335
rect 93 -2338 150 -2337
rect 163 -2338 353 -2337
rect 359 -2338 486 -2337
rect 534 -2338 626 -2337
rect 632 -2338 668 -2337
rect 702 -2338 822 -2337
rect 121 -2340 367 -2339
rect 401 -2340 444 -2339
rect 453 -2340 549 -2339
rect 555 -2340 563 -2339
rect 569 -2340 591 -2339
rect 604 -2340 608 -2339
rect 614 -2340 759 -2339
rect 779 -2340 815 -2339
rect 121 -2342 213 -2341
rect 226 -2342 402 -2341
rect 415 -2342 566 -2341
rect 569 -2342 612 -2341
rect 618 -2342 878 -2341
rect 149 -2344 311 -2343
rect 324 -2344 423 -2343
rect 429 -2344 465 -2343
rect 485 -2344 514 -2343
rect 555 -2344 619 -2343
rect 667 -2344 850 -2343
rect 72 -2346 514 -2345
rect 572 -2346 696 -2345
rect 730 -2346 780 -2345
rect 793 -2346 857 -2345
rect 72 -2348 318 -2347
rect 457 -2348 507 -2347
rect 576 -2348 661 -2347
rect 730 -2348 738 -2347
rect 758 -2348 766 -2347
rect 107 -2350 325 -2349
rect 464 -2350 528 -2349
rect 576 -2350 584 -2349
rect 590 -2350 598 -2349
rect 604 -2350 647 -2349
rect 660 -2350 675 -2349
rect 765 -2350 843 -2349
rect 107 -2352 381 -2351
rect 478 -2352 507 -2351
rect 583 -2352 689 -2351
rect 719 -2352 738 -2351
rect 156 -2354 213 -2353
rect 226 -2354 234 -2353
rect 236 -2354 696 -2353
rect 128 -2356 157 -2355
rect 247 -2356 426 -2355
rect 478 -2356 542 -2355
rect 597 -2356 640 -2355
rect 674 -2356 787 -2355
rect 128 -2358 220 -2357
rect 254 -2358 374 -2357
rect 499 -2358 612 -2357
rect 639 -2358 682 -2357
rect 191 -2360 248 -2359
rect 254 -2360 451 -2359
rect 527 -2360 689 -2359
rect 170 -2362 192 -2361
rect 219 -2362 269 -2361
rect 271 -2362 416 -2361
rect 681 -2362 745 -2361
rect 142 -2364 171 -2363
rect 289 -2364 542 -2363
rect 723 -2364 745 -2363
rect 100 -2366 290 -2365
rect 303 -2366 626 -2365
rect 79 -2368 304 -2367
rect 317 -2368 346 -2367
rect 408 -2368 500 -2367
rect 58 -2370 80 -2369
rect 100 -2370 164 -2369
rect 331 -2370 346 -2369
rect 408 -2370 654 -2369
rect 142 -2372 517 -2371
rect 653 -2372 808 -2371
rect 198 -2374 332 -2373
rect 177 -2376 199 -2375
rect 72 -2387 164 -2386
rect 166 -2387 199 -2386
rect 303 -2387 346 -2386
rect 355 -2387 542 -2386
rect 646 -2387 685 -2386
rect 723 -2387 731 -2386
rect 800 -2387 808 -2386
rect 814 -2387 829 -2386
rect 891 -2387 906 -2386
rect 940 -2387 1007 -2386
rect 79 -2389 188 -2388
rect 191 -2389 237 -2388
rect 303 -2389 402 -2388
rect 418 -2389 699 -2388
rect 730 -2389 745 -2388
rect 779 -2389 801 -2388
rect 975 -2389 990 -2388
rect 86 -2391 150 -2390
rect 156 -2391 174 -2390
rect 177 -2391 248 -2390
rect 282 -2391 402 -2390
rect 422 -2391 615 -2390
rect 688 -2391 745 -2390
rect 978 -2391 983 -2390
rect 93 -2393 185 -2392
rect 219 -2393 423 -2392
rect 429 -2393 489 -2392
rect 499 -2393 528 -2392
rect 530 -2393 626 -2392
rect 691 -2393 906 -2392
rect 121 -2395 269 -2394
rect 310 -2395 384 -2394
rect 394 -2395 510 -2394
rect 516 -2395 703 -2394
rect 135 -2397 451 -2396
rect 453 -2397 654 -2396
rect 142 -2399 199 -2398
rect 205 -2399 220 -2398
rect 247 -2399 262 -2398
rect 268 -2399 307 -2398
rect 310 -2399 409 -2398
rect 443 -2399 559 -2398
rect 576 -2399 626 -2398
rect 653 -2399 675 -2398
rect 261 -2401 325 -2400
rect 345 -2401 384 -2400
rect 436 -2401 444 -2400
rect 450 -2401 465 -2400
rect 499 -2401 507 -2400
rect 516 -2401 584 -2400
rect 674 -2401 717 -2400
rect 254 -2403 325 -2402
rect 352 -2403 542 -2402
rect 548 -2403 647 -2402
rect 716 -2403 752 -2402
rect 128 -2405 255 -2404
rect 296 -2405 395 -2404
rect 415 -2405 465 -2404
rect 492 -2405 507 -2404
rect 513 -2405 584 -2404
rect 709 -2405 752 -2404
rect 212 -2407 297 -2406
rect 359 -2407 409 -2406
rect 436 -2407 458 -2406
rect 460 -2407 486 -2406
rect 492 -2407 535 -2406
rect 548 -2407 556 -2406
rect 576 -2407 598 -2406
rect 289 -2409 360 -2408
rect 366 -2409 612 -2408
rect 100 -2411 290 -2410
rect 369 -2411 388 -2410
rect 478 -2411 535 -2410
rect 555 -2411 689 -2410
rect 114 -2413 388 -2412
rect 523 -2413 570 -2412
rect 597 -2413 605 -2412
rect 611 -2413 633 -2412
rect 331 -2415 479 -2414
rect 604 -2415 668 -2414
rect 233 -2417 332 -2416
rect 373 -2417 514 -2416
rect 632 -2417 661 -2416
rect 667 -2417 682 -2416
rect 226 -2419 234 -2418
rect 338 -2419 374 -2418
rect 471 -2419 570 -2418
rect 618 -2419 661 -2418
rect 681 -2419 766 -2418
rect 107 -2421 227 -2420
rect 317 -2421 339 -2420
rect 471 -2421 563 -2420
rect 618 -2421 640 -2420
rect 758 -2421 766 -2420
rect 275 -2423 318 -2422
rect 562 -2423 591 -2422
rect 737 -2423 759 -2422
rect 275 -2425 381 -2424
rect 520 -2425 591 -2424
rect 737 -2425 773 -2424
rect 282 -2427 381 -2426
rect 429 -2427 521 -2426
rect 772 -2427 794 -2426
rect 226 -2438 353 -2437
rect 380 -2438 472 -2437
rect 509 -2438 577 -2437
rect 607 -2438 619 -2437
rect 639 -2438 692 -2437
rect 702 -2438 717 -2437
rect 744 -2438 759 -2437
rect 807 -2438 818 -2437
rect 898 -2438 906 -2437
rect 219 -2440 227 -2439
rect 233 -2440 244 -2439
rect 261 -2440 367 -2439
rect 387 -2440 514 -2439
rect 569 -2440 612 -2439
rect 614 -2440 909 -2439
rect 233 -2442 248 -2441
rect 275 -2442 370 -2441
rect 387 -2442 430 -2441
rect 432 -2442 563 -2441
rect 572 -2442 598 -2441
rect 611 -2442 654 -2441
rect 660 -2442 664 -2441
rect 688 -2442 738 -2441
rect 747 -2442 766 -2441
rect 800 -2442 808 -2441
rect 891 -2442 899 -2441
rect 236 -2444 328 -2443
rect 331 -2444 458 -2443
rect 460 -2444 839 -2443
rect 282 -2446 419 -2445
rect 450 -2446 507 -2445
rect 509 -2446 584 -2445
rect 590 -2446 619 -2445
rect 625 -2446 654 -2445
rect 660 -2446 675 -2445
rect 730 -2446 745 -2445
rect 751 -2446 755 -2445
rect 296 -2448 332 -2447
rect 338 -2448 367 -2447
rect 401 -2448 454 -2447
rect 457 -2448 524 -2447
rect 576 -2448 605 -2447
rect 625 -2448 650 -2447
rect 663 -2448 675 -2447
rect 751 -2448 773 -2447
rect 254 -2450 297 -2449
rect 310 -2450 353 -2449
rect 373 -2450 402 -2449
rect 453 -2450 500 -2449
rect 597 -2450 633 -2449
rect 646 -2450 689 -2449
rect 198 -2452 255 -2451
rect 268 -2452 311 -2451
rect 317 -2452 451 -2451
rect 464 -2452 472 -2451
rect 499 -2452 535 -2451
rect 541 -2452 633 -2451
rect 646 -2452 668 -2451
rect 341 -2454 549 -2453
rect 345 -2456 374 -2455
rect 443 -2456 465 -2455
rect 478 -2456 549 -2455
rect 303 -2458 346 -2457
rect 348 -2458 556 -2457
rect 394 -2460 444 -2459
rect 478 -2460 486 -2459
rect 527 -2460 542 -2459
rect 359 -2462 395 -2461
rect 422 -2462 486 -2461
rect 492 -2462 528 -2461
rect 289 -2464 360 -2463
rect 415 -2464 493 -2463
rect 422 -2466 437 -2465
rect 436 -2468 517 -2467
rect 247 -2479 255 -2478
rect 296 -2479 342 -2478
rect 359 -2479 381 -2478
rect 390 -2479 458 -2478
rect 492 -2479 510 -2478
rect 513 -2479 612 -2478
rect 649 -2479 654 -2478
rect 674 -2479 692 -2478
rect 726 -2479 902 -2478
rect 310 -2481 349 -2480
rect 359 -2481 388 -2480
rect 394 -2481 430 -2480
rect 432 -2481 500 -2480
rect 527 -2481 535 -2480
rect 541 -2481 556 -2480
rect 604 -2481 640 -2480
rect 653 -2481 661 -2480
rect 688 -2481 696 -2480
rect 744 -2481 752 -2480
rect 807 -2481 818 -2480
rect 828 -2481 836 -2480
rect 898 -2481 906 -2480
rect 331 -2483 370 -2482
rect 373 -2483 395 -2482
rect 401 -2483 409 -2482
rect 443 -2483 472 -2482
rect 548 -2483 615 -2482
rect 632 -2483 661 -2482
rect 688 -2483 703 -2482
rect 352 -2485 374 -2484
rect 404 -2485 423 -2484
rect 446 -2485 465 -2484
rect 485 -2485 549 -2484
rect 551 -2485 577 -2484
rect 597 -2485 605 -2484
rect 614 -2485 626 -2484
rect 695 -2485 703 -2484
rect 366 -2487 388 -2486
rect 453 -2487 479 -2486
rect 618 -2487 633 -2486
rect 366 -2489 437 -2488
rect 226 -2500 234 -2499
rect 236 -2500 241 -2499
rect 359 -2500 367 -2499
rect 373 -2500 395 -2499
rect 397 -2500 409 -2499
rect 534 -2500 549 -2499
rect 558 -2500 902 -2499
rect 380 -2502 402 -2501
rect 604 -2502 612 -2501
rect 632 -2502 654 -2501
rect 660 -2502 692 -2501
rect 702 -2502 727 -2501
rect 898 -2502 906 -2501
<< m2contact >>
rect 152 0 153 1
rect 205 0 206 1
rect 338 0 339 1
rect 352 0 353 1
rect 366 0 367 1
rect 411 0 412 1
rect 432 0 433 1
rect 513 0 514 1
rect 341 -2 342 -1
rect 359 -2 360 -1
rect 394 -2 395 -1
rect 471 -2 472 -1
rect 492 -2 493 -1
rect 576 -2 577 -1
rect 345 -4 346 -3
rect 376 -4 377 -3
rect 408 -4 409 -3
rect 450 -4 451 -3
rect 464 -4 465 -3
rect 481 -4 482 -3
rect 128 -15 129 -14
rect 149 -15 150 -14
rect 198 -15 199 -14
rect 289 -15 290 -14
rect 292 -15 293 -14
rect 310 -15 311 -14
rect 320 -15 321 -14
rect 457 -15 458 -14
rect 464 -15 465 -14
rect 485 -15 486 -14
rect 502 -15 503 -14
rect 548 -15 549 -14
rect 576 -15 577 -14
rect 625 -15 626 -14
rect 208 -17 209 -16
rect 219 -17 220 -16
rect 243 -17 244 -16
rect 254 -17 255 -16
rect 282 -17 283 -16
rect 341 -17 342 -16
rect 352 -17 353 -16
rect 380 -17 381 -16
rect 415 -17 416 -16
rect 492 -17 493 -16
rect 513 -17 514 -16
rect 541 -17 542 -16
rect 593 -17 594 -16
rect 618 -17 619 -16
rect 296 -19 297 -18
rect 446 -19 447 -18
rect 450 -19 451 -18
rect 471 -19 472 -18
rect 474 -19 475 -18
rect 527 -19 528 -18
rect 303 -21 304 -20
rect 432 -21 433 -20
rect 450 -21 451 -20
rect 478 -21 479 -20
rect 324 -23 325 -22
rect 345 -23 346 -22
rect 352 -23 353 -22
rect 432 -23 433 -22
rect 436 -23 437 -22
rect 478 -23 479 -22
rect 327 -25 328 -24
rect 408 -25 409 -24
rect 429 -25 430 -24
rect 513 -25 514 -24
rect 331 -27 332 -26
rect 366 -27 367 -26
rect 376 -27 377 -26
rect 387 -27 388 -26
rect 401 -27 402 -26
rect 436 -27 437 -26
rect 464 -27 465 -26
rect 534 -27 535 -26
rect 338 -29 339 -28
rect 394 -29 395 -28
rect 401 -29 402 -28
rect 439 -29 440 -28
rect 345 -31 346 -30
rect 404 -31 405 -30
rect 366 -33 367 -32
rect 373 -33 374 -32
rect 394 -33 395 -32
rect 422 -33 423 -32
rect 373 -35 374 -34
rect 506 -35 507 -34
rect 114 -46 115 -45
rect 128 -46 129 -45
rect 142 -46 143 -45
rect 198 -46 199 -45
rect 205 -46 206 -45
rect 219 -46 220 -45
rect 233 -46 234 -45
rect 243 -46 244 -45
rect 247 -46 248 -45
rect 390 -46 391 -45
rect 415 -46 416 -45
rect 429 -46 430 -45
rect 432 -46 433 -45
rect 569 -46 570 -45
rect 593 -46 594 -45
rect 681 -46 682 -45
rect 170 -48 171 -47
rect 240 -48 241 -47
rect 254 -48 255 -47
rect 275 -48 276 -47
rect 317 -48 318 -47
rect 387 -48 388 -47
rect 443 -48 444 -47
rect 555 -48 556 -47
rect 593 -48 594 -47
rect 597 -48 598 -47
rect 618 -48 619 -47
rect 646 -48 647 -47
rect 653 -48 654 -47
rect 691 -48 692 -47
rect 191 -50 192 -49
rect 296 -50 297 -49
rect 331 -50 332 -49
rect 415 -50 416 -49
rect 443 -50 444 -49
rect 492 -50 493 -49
rect 495 -50 496 -49
rect 618 -50 619 -49
rect 625 -50 626 -49
rect 660 -50 661 -49
rect 674 -50 675 -49
rect 688 -50 689 -49
rect 198 -52 199 -51
rect 334 -52 335 -51
rect 338 -52 339 -51
rect 373 -52 374 -51
rect 394 -52 395 -51
rect 492 -52 493 -51
rect 502 -52 503 -51
rect 583 -52 584 -51
rect 212 -54 213 -53
rect 303 -54 304 -53
rect 338 -54 339 -53
rect 380 -54 381 -53
rect 478 -54 479 -53
rect 639 -54 640 -53
rect 219 -56 220 -55
rect 310 -56 311 -55
rect 369 -56 370 -55
rect 520 -56 521 -55
rect 527 -56 528 -55
rect 530 -56 531 -55
rect 534 -56 535 -55
rect 667 -56 668 -55
rect 240 -58 241 -57
rect 324 -58 325 -57
rect 380 -58 381 -57
rect 576 -58 577 -57
rect 254 -60 255 -59
rect 450 -60 451 -59
rect 478 -60 479 -59
rect 625 -60 626 -59
rect 177 -62 178 -61
rect 450 -62 451 -61
rect 485 -62 486 -61
rect 562 -62 563 -61
rect 261 -64 262 -63
rect 366 -64 367 -63
rect 408 -64 409 -63
rect 485 -64 486 -63
rect 499 -64 500 -63
rect 534 -64 535 -63
rect 548 -64 549 -63
rect 632 -64 633 -63
rect 226 -66 227 -65
rect 366 -66 367 -65
rect 387 -66 388 -65
rect 548 -66 549 -65
rect 268 -68 269 -67
rect 320 -68 321 -67
rect 408 -68 409 -67
rect 457 -68 458 -67
rect 506 -68 507 -67
rect 604 -68 605 -67
rect 282 -70 283 -69
rect 310 -70 311 -69
rect 436 -70 437 -69
rect 457 -70 458 -69
rect 474 -70 475 -69
rect 506 -70 507 -69
rect 513 -70 514 -69
rect 611 -70 612 -69
rect 282 -72 283 -71
rect 345 -72 346 -71
rect 422 -72 423 -71
rect 436 -72 437 -71
rect 446 -72 447 -71
rect 499 -72 500 -71
rect 527 -72 528 -71
rect 590 -72 591 -71
rect 163 -74 164 -73
rect 345 -74 346 -73
rect 422 -74 423 -73
rect 471 -74 472 -73
rect 530 -74 531 -73
rect 590 -74 591 -73
rect 289 -76 290 -75
rect 324 -76 325 -75
rect 464 -76 465 -75
rect 513 -76 514 -75
rect 289 -78 290 -77
rect 401 -78 402 -77
rect 296 -80 297 -79
rect 397 -80 398 -79
rect 184 -82 185 -81
rect 397 -82 398 -81
rect 303 -84 304 -83
rect 352 -84 353 -83
rect 373 -84 374 -83
rect 401 -84 402 -83
rect 348 -86 349 -85
rect 464 -86 465 -85
rect 352 -88 353 -87
rect 481 -88 482 -87
rect 51 -99 52 -98
rect 411 -99 412 -98
rect 464 -99 465 -98
rect 723 -99 724 -98
rect 58 -101 59 -100
rect 453 -101 454 -100
rect 471 -101 472 -100
rect 814 -101 815 -100
rect 65 -103 66 -102
rect 142 -103 143 -102
rect 145 -103 146 -102
rect 184 -103 185 -102
rect 198 -103 199 -102
rect 208 -103 209 -102
rect 275 -103 276 -102
rect 376 -103 377 -102
rect 394 -103 395 -102
rect 772 -103 773 -102
rect 72 -105 73 -104
rect 82 -105 83 -104
rect 86 -105 87 -104
rect 117 -105 118 -104
rect 121 -105 122 -104
rect 194 -105 195 -104
rect 198 -105 199 -104
rect 268 -105 269 -104
rect 275 -105 276 -104
rect 474 -105 475 -104
rect 485 -105 486 -104
rect 807 -105 808 -104
rect 93 -107 94 -106
rect 296 -107 297 -106
rect 331 -107 332 -106
rect 383 -107 384 -106
rect 485 -107 486 -106
rect 611 -107 612 -106
rect 632 -107 633 -106
rect 779 -107 780 -106
rect 107 -109 108 -108
rect 247 -109 248 -108
rect 268 -109 269 -108
rect 338 -109 339 -108
rect 345 -109 346 -108
rect 429 -109 430 -108
rect 492 -109 493 -108
rect 695 -109 696 -108
rect 114 -111 115 -110
rect 135 -111 136 -110
rect 156 -111 157 -110
rect 289 -111 290 -110
rect 359 -111 360 -110
rect 394 -111 395 -110
rect 418 -111 419 -110
rect 611 -111 612 -110
rect 639 -111 640 -110
rect 786 -111 787 -110
rect 114 -113 115 -112
rect 278 -113 279 -112
rect 324 -113 325 -112
rect 359 -113 360 -112
rect 366 -113 367 -112
rect 387 -113 388 -112
rect 450 -113 451 -112
rect 639 -113 640 -112
rect 653 -113 654 -112
rect 737 -113 738 -112
rect 128 -115 129 -114
rect 254 -115 255 -114
rect 261 -115 262 -114
rect 289 -115 290 -114
rect 310 -115 311 -114
rect 324 -115 325 -114
rect 369 -115 370 -114
rect 429 -115 430 -114
rect 495 -115 496 -114
rect 709 -115 710 -114
rect 152 -117 153 -116
rect 261 -117 262 -116
rect 303 -117 304 -116
rect 310 -117 311 -116
rect 387 -117 388 -116
rect 401 -117 402 -116
rect 520 -117 521 -116
rect 653 -117 654 -116
rect 660 -117 661 -116
rect 716 -117 717 -116
rect 170 -119 171 -118
rect 296 -119 297 -118
rect 303 -119 304 -118
rect 464 -119 465 -118
rect 478 -119 479 -118
rect 660 -119 661 -118
rect 667 -119 668 -118
rect 751 -119 752 -118
rect 170 -121 171 -120
rect 226 -121 227 -120
rect 247 -121 248 -120
rect 380 -121 381 -120
rect 534 -121 535 -120
rect 765 -121 766 -120
rect 100 -123 101 -122
rect 226 -123 227 -122
rect 254 -123 255 -122
rect 471 -123 472 -122
rect 534 -123 535 -122
rect 579 -123 580 -122
rect 583 -123 584 -122
rect 632 -123 633 -122
rect 646 -123 647 -122
rect 667 -123 668 -122
rect 674 -123 675 -122
rect 730 -123 731 -122
rect 184 -125 185 -124
rect 187 -125 188 -124
rect 201 -125 202 -124
rect 331 -125 332 -124
rect 380 -125 381 -124
rect 474 -125 475 -124
rect 499 -125 500 -124
rect 646 -125 647 -124
rect 681 -125 682 -124
rect 821 -125 822 -124
rect 219 -127 220 -126
rect 338 -127 339 -126
rect 436 -127 437 -126
rect 499 -127 500 -126
rect 513 -127 514 -126
rect 681 -127 682 -126
rect 688 -127 689 -126
rect 793 -127 794 -126
rect 191 -129 192 -128
rect 436 -129 437 -128
rect 467 -129 468 -128
rect 583 -129 584 -128
rect 590 -129 591 -128
rect 618 -129 619 -128
rect 625 -129 626 -128
rect 688 -129 689 -128
rect 219 -131 220 -130
rect 240 -131 241 -130
rect 317 -131 318 -130
rect 401 -131 402 -130
rect 453 -131 454 -130
rect 618 -131 619 -130
rect 205 -133 206 -132
rect 240 -133 241 -132
rect 282 -133 283 -132
rect 317 -133 318 -132
rect 481 -133 482 -132
rect 513 -133 514 -132
rect 527 -133 528 -132
rect 674 -133 675 -132
rect 177 -135 178 -134
rect 282 -135 283 -134
rect 506 -135 507 -134
rect 527 -135 528 -134
rect 548 -135 549 -134
rect 744 -135 745 -134
rect 177 -137 178 -136
rect 212 -137 213 -136
rect 373 -137 374 -136
rect 548 -137 549 -136
rect 562 -137 563 -136
rect 800 -137 801 -136
rect 163 -139 164 -138
rect 212 -139 213 -138
rect 334 -139 335 -138
rect 562 -139 563 -138
rect 569 -139 570 -138
rect 758 -139 759 -138
rect 163 -141 164 -140
rect 352 -141 353 -140
rect 373 -141 374 -140
rect 597 -141 598 -140
rect 205 -143 206 -142
rect 233 -143 234 -142
rect 352 -143 353 -142
rect 625 -143 626 -142
rect 208 -145 209 -144
rect 233 -145 234 -144
rect 415 -145 416 -144
rect 506 -145 507 -144
rect 541 -145 542 -144
rect 569 -145 570 -144
rect 576 -145 577 -144
rect 702 -145 703 -144
rect 345 -147 346 -146
rect 415 -147 416 -146
rect 422 -147 423 -146
rect 541 -147 542 -146
rect 555 -147 556 -146
rect 597 -147 598 -146
rect 422 -149 423 -148
rect 457 -149 458 -148
rect 520 -149 521 -148
rect 576 -149 577 -148
rect 443 -151 444 -150
rect 555 -151 556 -150
rect 408 -153 409 -152
rect 443 -153 444 -152
rect 457 -153 458 -152
rect 604 -153 605 -152
rect 593 -155 594 -154
rect 604 -155 605 -154
rect 44 -166 45 -165
rect 184 -166 185 -165
rect 191 -166 192 -165
rect 212 -166 213 -165
rect 268 -166 269 -165
rect 352 -166 353 -165
rect 362 -166 363 -165
rect 765 -166 766 -165
rect 793 -166 794 -165
rect 849 -166 850 -165
rect 65 -168 66 -167
rect 166 -168 167 -167
rect 184 -168 185 -167
rect 310 -168 311 -167
rect 348 -168 349 -167
rect 695 -168 696 -167
rect 751 -168 752 -167
rect 793 -168 794 -167
rect 800 -168 801 -167
rect 863 -168 864 -167
rect 65 -170 66 -169
rect 72 -170 73 -169
rect 79 -170 80 -169
rect 86 -170 87 -169
rect 100 -170 101 -169
rect 257 -170 258 -169
rect 310 -170 311 -169
rect 324 -170 325 -169
rect 352 -170 353 -169
rect 453 -170 454 -169
rect 464 -170 465 -169
rect 807 -170 808 -169
rect 814 -170 815 -169
rect 835 -170 836 -169
rect 72 -172 73 -171
rect 359 -172 360 -171
rect 408 -172 409 -171
rect 786 -172 787 -171
rect 821 -172 822 -171
rect 842 -172 843 -171
rect 86 -174 87 -173
rect 194 -174 195 -173
rect 198 -174 199 -173
rect 233 -174 234 -173
rect 324 -174 325 -173
rect 422 -174 423 -173
rect 471 -174 472 -173
rect 807 -174 808 -173
rect 103 -176 104 -175
rect 355 -176 356 -175
rect 411 -176 412 -175
rect 723 -176 724 -175
rect 730 -176 731 -175
rect 786 -176 787 -175
rect 117 -178 118 -177
rect 765 -178 766 -177
rect 772 -178 773 -177
rect 814 -178 815 -177
rect 121 -180 122 -179
rect 201 -180 202 -179
rect 212 -180 213 -179
rect 275 -180 276 -179
rect 285 -180 286 -179
rect 422 -180 423 -179
rect 492 -180 493 -179
rect 548 -180 549 -179
rect 576 -180 577 -179
rect 828 -180 829 -179
rect 121 -182 122 -181
rect 124 -182 125 -181
rect 128 -182 129 -181
rect 464 -182 465 -181
rect 495 -182 496 -181
rect 744 -182 745 -181
rect 779 -182 780 -181
rect 821 -182 822 -181
rect 128 -184 129 -183
rect 226 -184 227 -183
rect 275 -184 276 -183
rect 317 -184 318 -183
rect 415 -184 416 -183
rect 758 -184 759 -183
rect 138 -186 139 -185
rect 425 -186 426 -185
rect 460 -186 461 -185
rect 758 -186 759 -185
rect 145 -188 146 -187
rect 366 -188 367 -187
rect 415 -188 416 -187
rect 478 -188 479 -187
rect 495 -188 496 -187
rect 737 -188 738 -187
rect 163 -190 164 -189
rect 408 -190 409 -189
rect 443 -190 444 -189
rect 478 -190 479 -189
rect 499 -190 500 -189
rect 576 -190 577 -189
rect 632 -190 633 -189
rect 800 -190 801 -189
rect 58 -192 59 -191
rect 163 -192 164 -191
rect 177 -192 178 -191
rect 233 -192 234 -191
rect 296 -192 297 -191
rect 317 -192 318 -191
rect 359 -192 360 -191
rect 737 -192 738 -191
rect 51 -194 52 -193
rect 58 -194 59 -193
rect 177 -194 178 -193
rect 247 -194 248 -193
rect 282 -194 283 -193
rect 296 -194 297 -193
rect 366 -194 367 -193
rect 401 -194 402 -193
rect 443 -194 444 -193
rect 481 -194 482 -193
rect 520 -194 521 -193
rect 523 -194 524 -193
rect 548 -194 549 -193
rect 562 -194 563 -193
rect 660 -194 661 -193
rect 723 -194 724 -193
rect 730 -194 731 -193
rect 859 -194 860 -193
rect 51 -196 52 -195
rect 387 -196 388 -195
rect 450 -196 451 -195
rect 632 -196 633 -195
rect 667 -196 668 -195
rect 695 -196 696 -195
rect 709 -196 710 -195
rect 751 -196 752 -195
rect 191 -198 192 -197
rect 219 -198 220 -197
rect 247 -198 248 -197
rect 380 -198 381 -197
rect 429 -198 430 -197
rect 450 -198 451 -197
rect 457 -198 458 -197
rect 499 -198 500 -197
rect 520 -198 521 -197
rect 534 -198 535 -197
rect 618 -198 619 -197
rect 660 -198 661 -197
rect 681 -198 682 -197
rect 779 -198 780 -197
rect 205 -200 206 -199
rect 219 -200 220 -199
rect 226 -200 227 -199
rect 457 -200 458 -199
rect 474 -200 475 -199
rect 667 -200 668 -199
rect 688 -200 689 -199
rect 744 -200 745 -199
rect 205 -202 206 -201
rect 254 -202 255 -201
rect 303 -202 304 -201
rect 380 -202 381 -201
rect 394 -202 395 -201
rect 429 -202 430 -201
rect 439 -202 440 -201
rect 618 -202 619 -201
rect 646 -202 647 -201
rect 688 -202 689 -201
rect 702 -202 703 -201
rect 709 -202 710 -201
rect 716 -202 717 -201
rect 772 -202 773 -201
rect 156 -204 157 -203
rect 394 -204 395 -203
rect 474 -204 475 -203
rect 541 -204 542 -203
rect 653 -204 654 -203
rect 681 -204 682 -203
rect 114 -206 115 -205
rect 156 -206 157 -205
rect 254 -206 255 -205
rect 268 -206 269 -205
rect 289 -206 290 -205
rect 303 -206 304 -205
rect 331 -206 332 -205
rect 401 -206 402 -205
rect 404 -206 405 -205
rect 541 -206 542 -205
rect 639 -206 640 -205
rect 653 -206 654 -205
rect 674 -206 675 -205
rect 702 -206 703 -205
rect 289 -208 290 -207
rect 646 -208 647 -207
rect 331 -210 332 -209
rect 436 -210 437 -209
rect 492 -210 493 -209
rect 716 -210 717 -209
rect 338 -212 339 -211
rect 436 -212 437 -211
rect 523 -212 524 -211
rect 534 -212 535 -211
rect 569 -212 570 -211
rect 639 -212 640 -211
rect 261 -214 262 -213
rect 338 -214 339 -213
rect 373 -214 374 -213
rect 387 -214 388 -213
rect 527 -214 528 -213
rect 562 -214 563 -213
rect 611 -214 612 -213
rect 674 -214 675 -213
rect 261 -216 262 -215
rect 345 -216 346 -215
rect 506 -216 507 -215
rect 527 -216 528 -215
rect 555 -216 556 -215
rect 569 -216 570 -215
rect 583 -216 584 -215
rect 611 -216 612 -215
rect 107 -218 108 -217
rect 583 -218 584 -217
rect 107 -220 108 -219
rect 282 -220 283 -219
rect 345 -220 346 -219
rect 625 -220 626 -219
rect 142 -222 143 -221
rect 506 -222 507 -221
rect 597 -222 598 -221
rect 625 -222 626 -221
rect 142 -224 143 -223
rect 376 -224 377 -223
rect 597 -224 598 -223
rect 604 -224 605 -223
rect 149 -226 150 -225
rect 555 -226 556 -225
rect 590 -226 591 -225
rect 604 -226 605 -225
rect 149 -228 150 -227
rect 170 -228 171 -227
rect 513 -228 514 -227
rect 590 -228 591 -227
rect 135 -230 136 -229
rect 170 -230 171 -229
rect 485 -230 486 -229
rect 513 -230 514 -229
rect 93 -232 94 -231
rect 485 -232 486 -231
rect 93 -234 94 -233
rect 152 -234 153 -233
rect 135 -236 136 -235
rect 292 -236 293 -235
rect 2 -247 3 -246
rect 68 -247 69 -246
rect 72 -247 73 -246
rect 348 -247 349 -246
rect 352 -247 353 -246
rect 779 -247 780 -246
rect 807 -247 808 -246
rect 905 -247 906 -246
rect 9 -249 10 -248
rect 285 -249 286 -248
rect 289 -249 290 -248
rect 310 -249 311 -248
rect 352 -249 353 -248
rect 534 -249 535 -248
rect 569 -249 570 -248
rect 940 -249 941 -248
rect 16 -251 17 -250
rect 359 -251 360 -250
rect 383 -251 384 -250
rect 674 -251 675 -250
rect 681 -251 682 -250
rect 891 -251 892 -250
rect 23 -253 24 -252
rect 58 -253 59 -252
rect 72 -253 73 -252
rect 268 -253 269 -252
rect 289 -253 290 -252
rect 450 -253 451 -252
rect 471 -253 472 -252
rect 856 -253 857 -252
rect 30 -255 31 -254
rect 453 -255 454 -254
rect 492 -255 493 -254
rect 611 -255 612 -254
rect 730 -255 731 -254
rect 884 -255 885 -254
rect 37 -257 38 -256
rect 65 -257 66 -256
rect 86 -257 87 -256
rect 292 -257 293 -256
rect 303 -257 304 -256
rect 310 -257 311 -256
rect 359 -257 360 -256
rect 495 -257 496 -256
rect 520 -257 521 -256
rect 523 -257 524 -256
rect 548 -257 549 -256
rect 611 -257 612 -256
rect 667 -257 668 -256
rect 730 -257 731 -256
rect 744 -257 745 -256
rect 779 -257 780 -256
rect 814 -257 815 -256
rect 954 -257 955 -256
rect 51 -259 52 -258
rect 254 -259 255 -258
rect 268 -259 269 -258
rect 338 -259 339 -258
rect 401 -259 402 -258
rect 590 -259 591 -258
rect 597 -259 598 -258
rect 681 -259 682 -258
rect 758 -259 759 -258
rect 870 -259 871 -258
rect 51 -261 52 -260
rect 394 -261 395 -260
rect 418 -261 419 -260
rect 807 -261 808 -260
rect 821 -261 822 -260
rect 919 -261 920 -260
rect 58 -263 59 -262
rect 499 -263 500 -262
rect 506 -263 507 -262
rect 744 -263 745 -262
rect 758 -263 759 -262
rect 800 -263 801 -262
rect 828 -263 829 -262
rect 926 -263 927 -262
rect 65 -265 66 -264
rect 912 -265 913 -264
rect 79 -267 80 -266
rect 86 -267 87 -266
rect 93 -267 94 -266
rect 282 -267 283 -266
rect 303 -267 304 -266
rect 306 -267 307 -266
rect 376 -267 377 -266
rect 499 -267 500 -266
rect 520 -267 521 -266
rect 527 -267 528 -266
rect 555 -267 556 -266
rect 674 -267 675 -266
rect 751 -267 752 -266
rect 800 -267 801 -266
rect 835 -267 836 -266
rect 933 -267 934 -266
rect 79 -269 80 -268
rect 443 -269 444 -268
rect 464 -269 465 -268
rect 506 -269 507 -268
rect 541 -269 542 -268
rect 555 -269 556 -268
rect 569 -269 570 -268
rect 597 -269 598 -268
rect 653 -269 654 -268
rect 667 -269 668 -268
rect 723 -269 724 -268
rect 751 -269 752 -268
rect 765 -269 766 -268
rect 828 -269 829 -268
rect 842 -269 843 -268
rect 947 -269 948 -268
rect 93 -271 94 -270
rect 100 -271 101 -270
rect 103 -271 104 -270
rect 590 -271 591 -270
rect 632 -271 633 -270
rect 653 -271 654 -270
rect 709 -271 710 -270
rect 723 -271 724 -270
rect 793 -271 794 -270
rect 814 -271 815 -270
rect 849 -271 850 -270
rect 877 -271 878 -270
rect 100 -273 101 -272
rect 415 -273 416 -272
rect 425 -273 426 -272
rect 863 -273 864 -272
rect 121 -275 122 -274
rect 163 -275 164 -274
rect 170 -275 171 -274
rect 282 -275 283 -274
rect 338 -275 339 -274
rect 376 -275 377 -274
rect 387 -275 388 -274
rect 443 -275 444 -274
rect 450 -275 451 -274
rect 842 -275 843 -274
rect 121 -277 122 -276
rect 366 -277 367 -276
rect 394 -277 395 -276
rect 688 -277 689 -276
rect 702 -277 703 -276
rect 863 -277 864 -276
rect 142 -279 143 -278
rect 257 -279 258 -278
rect 366 -279 367 -278
rect 548 -279 549 -278
rect 576 -279 577 -278
rect 579 -279 580 -278
rect 583 -279 584 -278
rect 632 -279 633 -278
rect 646 -279 647 -278
rect 702 -279 703 -278
rect 772 -279 773 -278
rect 849 -279 850 -278
rect 142 -281 143 -280
rect 467 -281 468 -280
rect 474 -281 475 -280
rect 541 -281 542 -280
rect 576 -281 577 -280
rect 604 -281 605 -280
rect 625 -281 626 -280
rect 646 -281 647 -280
rect 660 -281 661 -280
rect 709 -281 710 -280
rect 716 -281 717 -280
rect 772 -281 773 -280
rect 786 -281 787 -280
rect 793 -281 794 -280
rect 156 -283 157 -282
rect 387 -283 388 -282
rect 397 -283 398 -282
rect 821 -283 822 -282
rect 156 -285 157 -284
rect 275 -285 276 -284
rect 425 -285 426 -284
rect 534 -285 535 -284
rect 551 -285 552 -284
rect 716 -285 717 -284
rect 737 -285 738 -284
rect 786 -285 787 -284
rect 163 -287 164 -286
rect 261 -287 262 -286
rect 275 -287 276 -286
rect 345 -287 346 -286
rect 436 -287 437 -286
rect 835 -287 836 -286
rect 44 -289 45 -288
rect 436 -289 437 -288
rect 439 -289 440 -288
rect 765 -289 766 -288
rect 170 -291 171 -290
rect 331 -291 332 -290
rect 457 -291 458 -290
rect 583 -291 584 -290
rect 639 -291 640 -290
rect 660 -291 661 -290
rect 688 -291 689 -290
rect 898 -291 899 -290
rect 128 -293 129 -292
rect 331 -293 332 -292
rect 457 -293 458 -292
rect 639 -293 640 -292
rect 695 -293 696 -292
rect 737 -293 738 -292
rect 184 -295 185 -294
rect 362 -295 363 -294
rect 478 -295 479 -294
rect 492 -295 493 -294
rect 579 -295 580 -294
rect 604 -295 605 -294
rect 618 -295 619 -294
rect 695 -295 696 -294
rect 166 -297 167 -296
rect 618 -297 619 -296
rect 184 -299 185 -298
rect 191 -299 192 -298
rect 205 -299 206 -298
rect 404 -299 405 -298
rect 478 -299 479 -298
rect 485 -299 486 -298
rect 488 -299 489 -298
rect 625 -299 626 -298
rect 107 -301 108 -300
rect 191 -301 192 -300
rect 205 -301 206 -300
rect 219 -301 220 -300
rect 254 -301 255 -300
rect 474 -301 475 -300
rect 485 -301 486 -300
rect 562 -301 563 -300
rect 107 -303 108 -302
rect 124 -303 125 -302
rect 219 -303 220 -302
rect 233 -303 234 -302
rect 261 -303 262 -302
rect 422 -303 423 -302
rect 446 -303 447 -302
rect 562 -303 563 -302
rect 198 -305 199 -304
rect 233 -305 234 -304
rect 247 -305 248 -304
rect 422 -305 423 -304
rect 114 -307 115 -306
rect 247 -307 248 -306
rect 317 -307 318 -306
rect 345 -307 346 -306
rect 114 -309 115 -308
rect 429 -309 430 -308
rect 198 -311 199 -310
rect 296 -311 297 -310
rect 380 -311 381 -310
rect 429 -311 430 -310
rect 44 -313 45 -312
rect 380 -313 381 -312
rect 135 -315 136 -314
rect 296 -315 297 -314
rect 135 -317 136 -316
rect 212 -317 213 -316
rect 226 -317 227 -316
rect 317 -317 318 -316
rect 212 -319 213 -318
rect 324 -319 325 -318
rect 226 -321 227 -320
rect 408 -321 409 -320
rect 117 -323 118 -322
rect 408 -323 409 -322
rect 324 -325 325 -324
rect 355 -325 356 -324
rect 16 -336 17 -335
rect 415 -336 416 -335
rect 436 -336 437 -335
rect 681 -336 682 -335
rect 905 -336 906 -335
rect 961 -336 962 -335
rect 16 -338 17 -337
rect 107 -338 108 -337
rect 124 -338 125 -337
rect 282 -338 283 -337
rect 289 -338 290 -337
rect 397 -338 398 -337
rect 401 -338 402 -337
rect 695 -338 696 -337
rect 758 -338 759 -337
rect 905 -338 906 -337
rect 912 -338 913 -337
rect 1024 -338 1025 -337
rect 44 -340 45 -339
rect 75 -340 76 -339
rect 79 -340 80 -339
rect 415 -340 416 -339
rect 439 -340 440 -339
rect 572 -340 573 -339
rect 618 -340 619 -339
rect 1003 -340 1004 -339
rect 37 -342 38 -341
rect 79 -342 80 -341
rect 96 -342 97 -341
rect 681 -342 682 -341
rect 730 -342 731 -341
rect 758 -342 759 -341
rect 779 -342 780 -341
rect 912 -342 913 -341
rect 919 -342 920 -341
rect 982 -342 983 -341
rect 2 -344 3 -343
rect 37 -344 38 -343
rect 44 -344 45 -343
rect 93 -344 94 -343
rect 100 -344 101 -343
rect 282 -344 283 -343
rect 296 -344 297 -343
rect 303 -344 304 -343
rect 310 -344 311 -343
rect 460 -344 461 -343
rect 467 -344 468 -343
rect 884 -344 885 -343
rect 926 -344 927 -343
rect 989 -344 990 -343
rect 2 -346 3 -345
rect 345 -346 346 -345
rect 355 -346 356 -345
rect 436 -346 437 -345
rect 443 -346 444 -345
rect 996 -346 997 -345
rect 51 -348 52 -347
rect 460 -348 461 -347
rect 467 -348 468 -347
rect 898 -348 899 -347
rect 933 -348 934 -347
rect 975 -348 976 -347
rect 51 -350 52 -349
rect 488 -350 489 -349
rect 548 -350 549 -349
rect 968 -350 969 -349
rect 65 -352 66 -351
rect 163 -352 164 -351
rect 191 -352 192 -351
rect 310 -352 311 -351
rect 331 -352 332 -351
rect 401 -352 402 -351
rect 411 -352 412 -351
rect 940 -352 941 -351
rect 93 -354 94 -353
rect 198 -354 199 -353
rect 212 -354 213 -353
rect 453 -354 454 -353
rect 457 -354 458 -353
rect 954 -354 955 -353
rect 100 -356 101 -355
rect 142 -356 143 -355
rect 149 -356 150 -355
rect 163 -356 164 -355
rect 198 -356 199 -355
rect 233 -356 234 -355
rect 243 -356 244 -355
rect 289 -356 290 -355
rect 296 -356 297 -355
rect 530 -356 531 -355
rect 583 -356 584 -355
rect 618 -356 619 -355
rect 621 -356 622 -355
rect 779 -356 780 -355
rect 793 -356 794 -355
rect 933 -356 934 -355
rect 107 -358 108 -357
rect 131 -358 132 -357
rect 142 -358 143 -357
rect 219 -358 220 -357
rect 226 -358 227 -357
rect 418 -358 419 -357
rect 422 -358 423 -357
rect 884 -358 885 -357
rect 72 -360 73 -359
rect 226 -360 227 -359
rect 233 -360 234 -359
rect 376 -360 377 -359
rect 380 -360 381 -359
rect 551 -360 552 -359
rect 667 -360 668 -359
rect 695 -360 696 -359
rect 751 -360 752 -359
rect 793 -360 794 -359
rect 800 -360 801 -359
rect 919 -360 920 -359
rect 114 -362 115 -361
rect 397 -362 398 -361
rect 446 -362 447 -361
rect 632 -362 633 -361
rect 744 -362 745 -361
rect 800 -362 801 -361
rect 842 -362 843 -361
rect 898 -362 899 -361
rect 86 -364 87 -363
rect 114 -364 115 -363
rect 177 -364 178 -363
rect 219 -364 220 -363
rect 254 -364 255 -363
rect 383 -364 384 -363
rect 387 -364 388 -363
rect 422 -364 423 -363
rect 457 -364 458 -363
rect 576 -364 577 -363
rect 597 -364 598 -363
rect 667 -364 668 -363
rect 702 -364 703 -363
rect 744 -364 745 -363
rect 786 -364 787 -363
rect 842 -364 843 -363
rect 849 -364 850 -363
rect 926 -364 927 -363
rect 177 -366 178 -365
rect 184 -366 185 -365
rect 194 -366 195 -365
rect 702 -366 703 -365
rect 737 -366 738 -365
rect 786 -366 787 -365
rect 814 -366 815 -365
rect 849 -366 850 -365
rect 856 -366 857 -365
rect 940 -366 941 -365
rect 128 -368 129 -367
rect 184 -368 185 -367
rect 254 -368 255 -367
rect 275 -368 276 -367
rect 338 -368 339 -367
rect 443 -368 444 -367
rect 464 -368 465 -367
rect 856 -368 857 -367
rect 877 -368 878 -367
rect 954 -368 955 -367
rect 128 -370 129 -369
rect 135 -370 136 -369
rect 156 -370 157 -369
rect 338 -370 339 -369
rect 352 -370 353 -369
rect 597 -370 598 -369
rect 632 -370 633 -369
rect 639 -370 640 -369
rect 660 -370 661 -369
rect 737 -370 738 -369
rect 835 -370 836 -369
rect 877 -370 878 -369
rect 86 -372 87 -371
rect 135 -372 136 -371
rect 156 -372 157 -371
rect 317 -372 318 -371
rect 359 -372 360 -371
rect 474 -372 475 -371
rect 485 -372 486 -371
rect 730 -372 731 -371
rect 772 -372 773 -371
rect 835 -372 836 -371
rect 170 -374 171 -373
rect 352 -374 353 -373
rect 373 -374 374 -373
rect 870 -374 871 -373
rect 82 -376 83 -375
rect 170 -376 171 -375
rect 212 -376 213 -375
rect 359 -376 360 -375
rect 387 -376 388 -375
rect 429 -376 430 -375
rect 464 -376 465 -375
rect 485 -376 486 -375
rect 516 -376 517 -375
rect 639 -376 640 -375
rect 646 -376 647 -375
rect 660 -376 661 -375
rect 709 -376 710 -375
rect 870 -376 871 -375
rect 261 -378 262 -377
rect 345 -378 346 -377
rect 425 -378 426 -377
rect 576 -378 577 -377
rect 653 -378 654 -377
rect 709 -378 710 -377
rect 723 -378 724 -377
rect 814 -378 815 -377
rect 247 -380 248 -379
rect 261 -380 262 -379
rect 268 -380 269 -379
rect 373 -380 374 -379
rect 429 -380 430 -379
rect 450 -380 451 -379
rect 471 -380 472 -379
rect 863 -380 864 -379
rect 72 -382 73 -381
rect 471 -382 472 -381
rect 541 -382 542 -381
rect 583 -382 584 -381
rect 625 -382 626 -381
rect 653 -382 654 -381
rect 674 -382 675 -381
rect 723 -382 724 -381
rect 821 -382 822 -381
rect 863 -382 864 -381
rect 121 -384 122 -383
rect 268 -384 269 -383
rect 275 -384 276 -383
rect 394 -384 395 -383
rect 506 -384 507 -383
rect 541 -384 542 -383
rect 551 -384 552 -383
rect 772 -384 773 -383
rect 23 -386 24 -385
rect 121 -386 122 -385
rect 240 -386 241 -385
rect 247 -386 248 -385
rect 306 -386 307 -385
rect 646 -386 647 -385
rect 765 -386 766 -385
rect 821 -386 822 -385
rect 23 -388 24 -387
rect 30 -388 31 -387
rect 58 -388 59 -387
rect 506 -388 507 -387
rect 520 -388 521 -387
rect 625 -388 626 -387
rect 716 -388 717 -387
rect 765 -388 766 -387
rect 30 -390 31 -389
rect 68 -390 69 -389
rect 149 -390 150 -389
rect 240 -390 241 -389
rect 317 -390 318 -389
rect 366 -390 367 -389
rect 394 -390 395 -389
rect 807 -390 808 -389
rect 58 -392 59 -391
rect 324 -392 325 -391
rect 362 -392 363 -391
rect 674 -392 675 -391
rect 688 -392 689 -391
rect 716 -392 717 -391
rect 68 -394 69 -393
rect 331 -394 332 -393
rect 366 -394 367 -393
rect 432 -394 433 -393
rect 513 -394 514 -393
rect 520 -394 521 -393
rect 562 -394 563 -393
rect 688 -394 689 -393
rect 324 -396 325 -395
rect 555 -396 556 -395
rect 569 -396 570 -395
rect 751 -396 752 -395
rect 499 -398 500 -397
rect 562 -398 563 -397
rect 569 -398 570 -397
rect 611 -398 612 -397
rect 478 -400 479 -399
rect 499 -400 500 -399
rect 513 -400 514 -399
rect 891 -400 892 -399
rect 478 -402 479 -401
rect 492 -402 493 -401
rect 527 -402 528 -401
rect 555 -402 556 -401
rect 590 -402 591 -401
rect 611 -402 612 -401
rect 828 -402 829 -401
rect 891 -402 892 -401
rect 9 -404 10 -403
rect 527 -404 528 -403
rect 534 -404 535 -403
rect 590 -404 591 -403
rect 604 -404 605 -403
rect 807 -404 808 -403
rect 9 -406 10 -405
rect 89 -406 90 -405
rect 159 -406 160 -405
rect 828 -406 829 -405
rect 404 -408 405 -407
rect 604 -408 605 -407
rect 408 -410 409 -409
rect 534 -410 535 -409
rect 408 -412 409 -411
rect 492 -412 493 -411
rect 9 -423 10 -422
rect 131 -423 132 -422
rect 142 -423 143 -422
rect 243 -423 244 -422
rect 275 -423 276 -422
rect 352 -423 353 -422
rect 362 -423 363 -422
rect 625 -423 626 -422
rect 814 -423 815 -422
rect 1073 -423 1074 -422
rect 9 -425 10 -424
rect 639 -425 640 -424
rect 849 -425 850 -424
rect 1045 -425 1046 -424
rect 16 -427 17 -426
rect 93 -427 94 -426
rect 156 -427 157 -426
rect 282 -427 283 -426
rect 324 -427 325 -426
rect 411 -427 412 -426
rect 415 -427 416 -426
rect 814 -427 815 -426
rect 912 -427 913 -426
rect 1031 -427 1032 -426
rect 16 -429 17 -428
rect 653 -429 654 -428
rect 765 -429 766 -428
rect 849 -429 850 -428
rect 926 -429 927 -428
rect 1052 -429 1053 -428
rect 23 -431 24 -430
rect 152 -431 153 -430
rect 191 -431 192 -430
rect 422 -431 423 -430
rect 429 -431 430 -430
rect 807 -431 808 -430
rect 828 -431 829 -430
rect 926 -431 927 -430
rect 933 -431 934 -430
rect 1010 -431 1011 -430
rect 1024 -431 1025 -430
rect 1087 -431 1088 -430
rect 23 -433 24 -432
rect 390 -433 391 -432
rect 394 -433 395 -432
rect 807 -433 808 -432
rect 828 -433 829 -432
rect 891 -433 892 -432
rect 940 -433 941 -432
rect 1038 -433 1039 -432
rect 30 -435 31 -434
rect 184 -435 185 -434
rect 226 -435 227 -434
rect 327 -435 328 -434
rect 373 -435 374 -434
rect 481 -435 482 -434
rect 513 -435 514 -434
rect 534 -435 535 -434
rect 548 -435 549 -434
rect 919 -435 920 -434
rect 940 -435 941 -434
rect 1003 -435 1004 -434
rect 30 -437 31 -436
rect 58 -437 59 -436
rect 65 -437 66 -436
rect 359 -437 360 -436
rect 397 -437 398 -436
rect 667 -437 668 -436
rect 670 -437 671 -436
rect 1003 -437 1004 -436
rect 37 -439 38 -438
rect 72 -439 73 -438
rect 86 -439 87 -438
rect 100 -439 101 -438
rect 163 -439 164 -438
rect 191 -439 192 -438
rect 219 -439 220 -438
rect 226 -439 227 -438
rect 275 -439 276 -438
rect 397 -439 398 -438
rect 401 -439 402 -438
rect 415 -439 416 -438
rect 432 -439 433 -438
rect 716 -439 717 -438
rect 730 -439 731 -438
rect 1024 -439 1025 -438
rect 37 -441 38 -440
rect 93 -441 94 -440
rect 100 -441 101 -440
rect 107 -441 108 -440
rect 184 -441 185 -440
rect 317 -441 318 -440
rect 324 -441 325 -440
rect 422 -441 423 -440
rect 450 -441 451 -440
rect 453 -441 454 -440
rect 467 -441 468 -440
rect 478 -441 479 -440
rect 523 -441 524 -440
rect 1101 -441 1102 -440
rect 44 -443 45 -442
rect 79 -443 80 -442
rect 187 -443 188 -442
rect 219 -443 220 -442
rect 296 -443 297 -442
rect 429 -443 430 -442
rect 450 -443 451 -442
rect 723 -443 724 -442
rect 730 -443 731 -442
rect 751 -443 752 -442
rect 786 -443 787 -442
rect 891 -443 892 -442
rect 954 -443 955 -442
rect 1059 -443 1060 -442
rect 44 -445 45 -444
rect 250 -445 251 -444
rect 310 -445 311 -444
rect 317 -445 318 -444
rect 331 -445 332 -444
rect 373 -445 374 -444
rect 401 -445 402 -444
rect 411 -445 412 -444
rect 478 -445 479 -444
rect 905 -445 906 -444
rect 961 -445 962 -444
rect 1094 -445 1095 -444
rect 51 -447 52 -446
rect 240 -447 241 -446
rect 247 -447 248 -446
rect 296 -447 297 -446
rect 331 -447 332 -446
rect 366 -447 367 -446
rect 460 -447 461 -446
rect 961 -447 962 -446
rect 968 -447 969 -446
rect 1108 -447 1109 -446
rect 51 -449 52 -448
rect 485 -449 486 -448
rect 530 -449 531 -448
rect 870 -449 871 -448
rect 975 -449 976 -448
rect 1080 -449 1081 -448
rect 58 -451 59 -450
rect 551 -451 552 -450
rect 562 -451 563 -450
rect 639 -451 640 -450
rect 649 -451 650 -450
rect 765 -451 766 -450
rect 772 -451 773 -450
rect 870 -451 871 -450
rect 884 -451 885 -450
rect 975 -451 976 -450
rect 982 -451 983 -450
rect 1115 -451 1116 -450
rect 65 -453 66 -452
rect 387 -453 388 -452
rect 408 -453 409 -452
rect 562 -453 563 -452
rect 576 -453 577 -452
rect 625 -453 626 -452
rect 674 -453 675 -452
rect 905 -453 906 -452
rect 989 -453 990 -452
rect 1122 -453 1123 -452
rect 68 -455 69 -454
rect 716 -455 717 -454
rect 737 -455 738 -454
rect 989 -455 990 -454
rect 996 -455 997 -454
rect 1066 -455 1067 -454
rect 72 -457 73 -456
rect 667 -457 668 -456
rect 709 -457 710 -456
rect 786 -457 787 -456
rect 800 -457 801 -456
rect 912 -457 913 -456
rect 75 -459 76 -458
rect 107 -459 108 -458
rect 121 -459 122 -458
rect 884 -459 885 -458
rect 79 -461 80 -460
rect 170 -461 171 -460
rect 205 -461 206 -460
rect 247 -461 248 -460
rect 261 -461 262 -460
rect 366 -461 367 -460
rect 387 -461 388 -460
rect 1017 -461 1018 -460
rect 82 -463 83 -462
rect 772 -463 773 -462
rect 779 -463 780 -462
rect 954 -463 955 -462
rect 121 -465 122 -464
rect 177 -465 178 -464
rect 233 -465 234 -464
rect 408 -465 409 -464
rect 485 -465 486 -464
rect 576 -465 577 -464
rect 597 -465 598 -464
rect 653 -465 654 -464
rect 702 -465 703 -464
rect 709 -465 710 -464
rect 744 -465 745 -464
rect 800 -465 801 -464
rect 821 -465 822 -464
rect 919 -465 920 -464
rect 128 -467 129 -466
rect 170 -467 171 -466
rect 177 -467 178 -466
rect 380 -467 381 -466
rect 520 -467 521 -466
rect 597 -467 598 -466
rect 604 -467 605 -466
rect 674 -467 675 -466
rect 681 -467 682 -466
rect 744 -467 745 -466
rect 835 -467 836 -466
rect 933 -467 934 -466
rect 96 -469 97 -468
rect 128 -469 129 -468
rect 135 -469 136 -468
rect 310 -469 311 -468
rect 338 -469 339 -468
rect 359 -469 360 -468
rect 464 -469 465 -468
rect 835 -469 836 -468
rect 856 -469 857 -468
rect 982 -469 983 -468
rect 96 -471 97 -470
rect 163 -471 164 -470
rect 212 -471 213 -470
rect 380 -471 381 -470
rect 464 -471 465 -470
rect 527 -471 528 -470
rect 534 -471 535 -470
rect 579 -471 580 -470
rect 607 -471 608 -470
rect 702 -471 703 -470
rect 793 -471 794 -470
rect 856 -471 857 -470
rect 863 -471 864 -470
rect 968 -471 969 -470
rect 156 -473 157 -472
rect 338 -473 339 -472
rect 471 -473 472 -472
rect 527 -473 528 -472
rect 548 -473 549 -472
rect 751 -473 752 -472
rect 758 -473 759 -472
rect 863 -473 864 -472
rect 877 -473 878 -472
rect 996 -473 997 -472
rect 149 -475 150 -474
rect 471 -475 472 -474
rect 509 -475 510 -474
rect 793 -475 794 -474
rect 212 -477 213 -476
rect 303 -477 304 -476
rect 516 -477 517 -476
rect 877 -477 878 -476
rect 2 -479 3 -478
rect 303 -479 304 -478
rect 520 -479 521 -478
rect 688 -479 689 -478
rect 2 -481 3 -480
rect 138 -481 139 -480
rect 233 -481 234 -480
rect 254 -481 255 -480
rect 261 -481 262 -480
rect 268 -481 269 -480
rect 572 -481 573 -480
rect 758 -481 759 -480
rect 124 -483 125 -482
rect 268 -483 269 -482
rect 604 -483 605 -482
rect 688 -483 689 -482
rect 240 -485 241 -484
rect 289 -485 290 -484
rect 611 -485 612 -484
rect 779 -485 780 -484
rect 254 -487 255 -486
rect 443 -487 444 -486
rect 618 -487 619 -486
rect 723 -487 724 -486
rect 205 -489 206 -488
rect 443 -489 444 -488
rect 569 -489 570 -488
rect 618 -489 619 -488
rect 621 -489 622 -488
rect 947 -489 948 -488
rect 289 -491 290 -490
rect 499 -491 500 -490
rect 569 -491 570 -490
rect 898 -491 899 -490
rect 345 -493 346 -492
rect 611 -493 612 -492
rect 632 -493 633 -492
rect 737 -493 738 -492
rect 842 -493 843 -492
rect 947 -493 948 -492
rect 159 -495 160 -494
rect 345 -495 346 -494
rect 436 -495 437 -494
rect 499 -495 500 -494
rect 583 -495 584 -494
rect 842 -495 843 -494
rect 394 -497 395 -496
rect 436 -497 437 -496
rect 446 -497 447 -496
rect 632 -497 633 -496
rect 646 -497 647 -496
rect 821 -497 822 -496
rect 457 -499 458 -498
rect 898 -499 899 -498
rect 457 -501 458 -500
rect 541 -501 542 -500
rect 583 -501 584 -500
rect 590 -501 591 -500
rect 660 -501 661 -500
rect 681 -501 682 -500
rect 492 -503 493 -502
rect 541 -503 542 -502
rect 565 -503 566 -502
rect 660 -503 661 -502
rect 453 -505 454 -504
rect 492 -505 493 -504
rect 506 -505 507 -504
rect 590 -505 591 -504
rect 282 -507 283 -506
rect 506 -507 507 -506
rect 2 -518 3 -517
rect 142 -518 143 -517
rect 149 -518 150 -517
rect 383 -518 384 -517
rect 390 -518 391 -517
rect 408 -518 409 -517
rect 411 -518 412 -517
rect 821 -518 822 -517
rect 2 -520 3 -519
rect 404 -520 405 -519
rect 425 -520 426 -519
rect 478 -520 479 -519
rect 509 -520 510 -519
rect 1115 -520 1116 -519
rect 9 -522 10 -521
rect 138 -522 139 -521
rect 159 -522 160 -521
rect 450 -522 451 -521
rect 544 -522 545 -521
rect 1108 -522 1109 -521
rect 9 -524 10 -523
rect 786 -524 787 -523
rect 821 -524 822 -523
rect 849 -524 850 -523
rect 16 -526 17 -525
rect 93 -526 94 -525
rect 107 -526 108 -525
rect 128 -526 129 -525
rect 177 -526 178 -525
rect 478 -526 479 -525
rect 572 -526 573 -525
rect 989 -526 990 -525
rect 58 -528 59 -527
rect 562 -528 563 -527
rect 576 -528 577 -527
rect 842 -528 843 -527
rect 989 -528 990 -527
rect 1017 -528 1018 -527
rect 72 -530 73 -529
rect 156 -530 157 -529
rect 177 -530 178 -529
rect 187 -530 188 -529
rect 212 -530 213 -529
rect 562 -530 563 -529
rect 579 -530 580 -529
rect 1122 -530 1123 -529
rect 75 -532 76 -531
rect 380 -532 381 -531
rect 429 -532 430 -531
rect 621 -532 622 -531
rect 628 -532 629 -531
rect 1073 -532 1074 -531
rect 79 -534 80 -533
rect 387 -534 388 -533
rect 415 -534 416 -533
rect 429 -534 430 -533
rect 443 -534 444 -533
rect 464 -534 465 -533
rect 555 -534 556 -533
rect 576 -534 577 -533
rect 646 -534 647 -533
rect 1031 -534 1032 -533
rect 58 -536 59 -535
rect 79 -536 80 -535
rect 86 -536 87 -535
rect 93 -536 94 -535
rect 128 -536 129 -535
rect 303 -536 304 -535
rect 317 -536 318 -535
rect 450 -536 451 -535
rect 464 -536 465 -535
rect 779 -536 780 -535
rect 786 -536 787 -535
rect 947 -536 948 -535
rect 1017 -536 1018 -535
rect 1038 -536 1039 -535
rect 86 -538 87 -537
rect 131 -538 132 -537
rect 145 -538 146 -537
rect 212 -538 213 -537
rect 240 -538 241 -537
rect 324 -538 325 -537
rect 387 -538 388 -537
rect 590 -538 591 -537
rect 667 -538 668 -537
rect 1094 -538 1095 -537
rect 51 -540 52 -539
rect 590 -540 591 -539
rect 674 -540 675 -539
rect 849 -540 850 -539
rect 947 -540 948 -539
rect 996 -540 997 -539
rect 1031 -540 1032 -539
rect 1045 -540 1046 -539
rect 51 -542 52 -541
rect 597 -542 598 -541
rect 674 -542 675 -541
rect 730 -542 731 -541
rect 754 -542 755 -541
rect 1101 -542 1102 -541
rect 121 -544 122 -543
rect 303 -544 304 -543
rect 446 -544 447 -543
rect 814 -544 815 -543
rect 828 -544 829 -543
rect 1073 -544 1074 -543
rect 72 -546 73 -545
rect 121 -546 122 -545
rect 135 -546 136 -545
rect 240 -546 241 -545
rect 247 -546 248 -545
rect 296 -546 297 -545
rect 481 -546 482 -545
rect 667 -546 668 -545
rect 695 -546 696 -545
rect 698 -546 699 -545
rect 730 -546 731 -545
rect 772 -546 773 -545
rect 807 -546 808 -545
rect 1045 -546 1046 -545
rect 135 -548 136 -547
rect 205 -548 206 -547
rect 247 -548 248 -547
rect 415 -548 416 -547
rect 520 -548 521 -547
rect 646 -548 647 -547
rect 695 -548 696 -547
rect 702 -548 703 -547
rect 772 -548 773 -547
rect 884 -548 885 -547
rect 996 -548 997 -547
rect 1024 -548 1025 -547
rect 1038 -548 1039 -547
rect 1059 -548 1060 -547
rect 145 -550 146 -549
rect 226 -550 227 -549
rect 250 -550 251 -549
rect 317 -550 318 -549
rect 471 -550 472 -549
rect 520 -550 521 -549
rect 551 -550 552 -549
rect 884 -550 885 -549
rect 1059 -550 1060 -549
rect 1066 -550 1067 -549
rect 37 -552 38 -551
rect 226 -552 227 -551
rect 261 -552 262 -551
rect 506 -552 507 -551
rect 555 -552 556 -551
rect 569 -552 570 -551
rect 597 -552 598 -551
rect 639 -552 640 -551
rect 698 -552 699 -551
rect 702 -552 703 -551
rect 723 -552 724 -551
rect 1024 -552 1025 -551
rect 44 -554 45 -553
rect 569 -554 570 -553
rect 632 -554 633 -553
rect 807 -554 808 -553
rect 814 -554 815 -553
rect 891 -554 892 -553
rect 940 -554 941 -553
rect 1066 -554 1067 -553
rect 44 -556 45 -555
rect 422 -556 423 -555
rect 436 -556 437 -555
rect 471 -556 472 -555
rect 492 -556 493 -555
rect 506 -556 507 -555
rect 583 -556 584 -555
rect 632 -556 633 -555
rect 639 -556 640 -555
rect 653 -556 654 -555
rect 723 -556 724 -555
rect 800 -556 801 -555
rect 828 -556 829 -555
rect 856 -556 857 -555
rect 940 -556 941 -555
rect 968 -556 969 -555
rect 156 -558 157 -557
rect 191 -558 192 -557
rect 205 -558 206 -557
rect 275 -558 276 -557
rect 289 -558 290 -557
rect 380 -558 381 -557
rect 422 -558 423 -557
rect 779 -558 780 -557
rect 800 -558 801 -557
rect 863 -558 864 -557
rect 114 -560 115 -559
rect 289 -560 290 -559
rect 296 -560 297 -559
rect 401 -560 402 -559
rect 492 -560 493 -559
rect 499 -560 500 -559
rect 583 -560 584 -559
rect 607 -560 608 -559
rect 653 -560 654 -559
rect 660 -560 661 -559
rect 835 -560 836 -559
rect 968 -560 969 -559
rect 100 -562 101 -561
rect 114 -562 115 -561
rect 152 -562 153 -561
rect 275 -562 276 -561
rect 338 -562 339 -561
rect 436 -562 437 -561
rect 499 -562 500 -561
rect 527 -562 528 -561
rect 604 -562 605 -561
rect 891 -562 892 -561
rect 30 -564 31 -563
rect 338 -564 339 -563
rect 401 -564 402 -563
rect 611 -564 612 -563
rect 660 -564 661 -563
rect 688 -564 689 -563
rect 835 -564 836 -563
rect 870 -564 871 -563
rect 30 -566 31 -565
rect 485 -566 486 -565
rect 513 -566 514 -565
rect 527 -566 528 -565
rect 604 -566 605 -565
rect 625 -566 626 -565
rect 842 -566 843 -565
rect 877 -566 878 -565
rect 16 -568 17 -567
rect 625 -568 626 -567
rect 856 -568 857 -567
rect 954 -568 955 -567
rect 100 -570 101 -569
rect 219 -570 220 -569
rect 261 -570 262 -569
rect 278 -570 279 -569
rect 352 -570 353 -569
rect 485 -570 486 -569
rect 513 -570 514 -569
rect 541 -570 542 -569
rect 863 -570 864 -569
rect 898 -570 899 -569
rect 954 -570 955 -569
rect 1003 -570 1004 -569
rect 37 -572 38 -571
rect 219 -572 220 -571
rect 254 -572 255 -571
rect 352 -572 353 -571
rect 394 -572 395 -571
rect 688 -572 689 -571
rect 870 -572 871 -571
rect 905 -572 906 -571
rect 975 -572 976 -571
rect 1003 -572 1004 -571
rect 191 -574 192 -573
rect 233 -574 234 -573
rect 254 -574 255 -573
rect 282 -574 283 -573
rect 394 -574 395 -573
rect 534 -574 535 -573
rect 541 -574 542 -573
rect 716 -574 717 -573
rect 877 -574 878 -573
rect 912 -574 913 -573
rect 975 -574 976 -573
rect 1010 -574 1011 -573
rect 233 -576 234 -575
rect 670 -576 671 -575
rect 716 -576 717 -575
rect 737 -576 738 -575
rect 898 -576 899 -575
rect 919 -576 920 -575
rect 1010 -576 1011 -575
rect 1080 -576 1081 -575
rect 107 -578 108 -577
rect 1080 -578 1081 -577
rect 282 -580 283 -579
rect 366 -580 367 -579
rect 457 -580 458 -579
rect 534 -580 535 -579
rect 565 -580 566 -579
rect 912 -580 913 -579
rect 919 -580 920 -579
rect 926 -580 927 -579
rect 65 -582 66 -581
rect 366 -582 367 -581
rect 457 -582 458 -581
rect 982 -582 983 -581
rect 65 -584 66 -583
rect 310 -584 311 -583
rect 523 -584 524 -583
rect 611 -584 612 -583
rect 709 -584 710 -583
rect 737 -584 738 -583
rect 751 -584 752 -583
rect 982 -584 983 -583
rect 170 -586 171 -585
rect 310 -586 311 -585
rect 373 -586 374 -585
rect 523 -586 524 -585
rect 565 -586 566 -585
rect 905 -586 906 -585
rect 170 -588 171 -587
rect 198 -588 199 -587
rect 345 -588 346 -587
rect 373 -588 374 -587
rect 681 -588 682 -587
rect 709 -588 710 -587
rect 751 -588 752 -587
rect 765 -588 766 -587
rect 198 -590 199 -589
rect 460 -590 461 -589
rect 618 -590 619 -589
rect 765 -590 766 -589
rect 345 -592 346 -591
rect 359 -592 360 -591
rect 453 -592 454 -591
rect 681 -592 682 -591
rect 758 -592 759 -591
rect 926 -592 927 -591
rect 184 -594 185 -593
rect 359 -594 360 -593
rect 618 -594 619 -593
rect 1052 -594 1053 -593
rect 23 -596 24 -595
rect 184 -596 185 -595
rect 744 -596 745 -595
rect 758 -596 759 -595
rect 933 -596 934 -595
rect 1052 -596 1053 -595
rect 23 -598 24 -597
rect 163 -598 164 -597
rect 744 -598 745 -597
rect 793 -598 794 -597
rect 933 -598 934 -597
rect 961 -598 962 -597
rect 163 -600 164 -599
rect 548 -600 549 -599
rect 334 -602 335 -601
rect 793 -602 794 -601
rect 467 -604 468 -603
rect 961 -604 962 -603
rect 548 -606 549 -605
rect 649 -606 650 -605
rect 23 -617 24 -616
rect 380 -617 381 -616
rect 415 -617 416 -616
rect 436 -617 437 -616
rect 453 -617 454 -616
rect 765 -617 766 -616
rect 905 -617 906 -616
rect 1213 -617 1214 -616
rect 1216 -617 1217 -616
rect 1360 -617 1361 -616
rect 40 -619 41 -618
rect 586 -619 587 -618
rect 618 -619 619 -618
rect 674 -619 675 -618
rect 716 -619 717 -618
rect 765 -619 766 -618
rect 814 -619 815 -618
rect 905 -619 906 -618
rect 961 -619 962 -618
rect 1157 -619 1158 -618
rect 2 -621 3 -620
rect 674 -621 675 -620
rect 702 -621 703 -620
rect 716 -621 717 -620
rect 723 -621 724 -620
rect 814 -621 815 -620
rect 961 -621 962 -620
rect 982 -621 983 -620
rect 989 -621 990 -620
rect 1101 -621 1102 -620
rect 2 -623 3 -622
rect 940 -623 941 -622
rect 975 -623 976 -622
rect 1094 -623 1095 -622
rect 44 -625 45 -624
rect 618 -625 619 -624
rect 621 -625 622 -624
rect 982 -625 983 -624
rect 996 -625 997 -624
rect 1108 -625 1109 -624
rect 44 -627 45 -626
rect 338 -627 339 -626
rect 380 -627 381 -626
rect 611 -627 612 -626
rect 635 -627 636 -626
rect 1052 -627 1053 -626
rect 1059 -627 1060 -626
rect 1192 -627 1193 -626
rect 47 -629 48 -628
rect 205 -629 206 -628
rect 229 -629 230 -628
rect 303 -629 304 -628
rect 324 -629 325 -628
rect 338 -629 339 -628
rect 387 -629 388 -628
rect 723 -629 724 -628
rect 726 -629 727 -628
rect 856 -629 857 -628
rect 884 -629 885 -628
rect 975 -629 976 -628
rect 1010 -629 1011 -628
rect 1185 -629 1186 -628
rect 51 -631 52 -630
rect 432 -631 433 -630
rect 460 -631 461 -630
rect 625 -631 626 -630
rect 649 -631 650 -630
rect 1171 -631 1172 -630
rect 58 -633 59 -632
rect 786 -633 787 -632
rect 821 -633 822 -632
rect 856 -633 857 -632
rect 870 -633 871 -632
rect 884 -633 885 -632
rect 891 -633 892 -632
rect 989 -633 990 -632
rect 1031 -633 1032 -632
rect 1129 -633 1130 -632
rect 51 -635 52 -634
rect 58 -635 59 -634
rect 65 -635 66 -634
rect 548 -635 549 -634
rect 551 -635 552 -634
rect 849 -635 850 -634
rect 898 -635 899 -634
rect 1010 -635 1011 -634
rect 1038 -635 1039 -634
rect 1122 -635 1123 -634
rect 65 -637 66 -636
rect 107 -637 108 -636
rect 121 -637 122 -636
rect 324 -637 325 -636
rect 331 -637 332 -636
rect 345 -637 346 -636
rect 404 -637 405 -636
rect 1052 -637 1053 -636
rect 1066 -637 1067 -636
rect 1199 -637 1200 -636
rect 16 -639 17 -638
rect 107 -639 108 -638
rect 121 -639 122 -638
rect 656 -639 657 -638
rect 667 -639 668 -638
rect 702 -639 703 -638
rect 730 -639 731 -638
rect 996 -639 997 -638
rect 1045 -639 1046 -638
rect 1080 -639 1081 -638
rect 1083 -639 1084 -638
rect 1087 -639 1088 -638
rect 16 -641 17 -640
rect 187 -641 188 -640
rect 226 -641 227 -640
rect 387 -641 388 -640
rect 418 -641 419 -640
rect 425 -641 426 -640
rect 464 -641 465 -640
rect 1164 -641 1165 -640
rect 75 -643 76 -642
rect 1003 -643 1004 -642
rect 86 -645 87 -644
rect 205 -645 206 -644
rect 247 -645 248 -644
rect 345 -645 346 -644
rect 422 -645 423 -644
rect 443 -645 444 -644
rect 464 -645 465 -644
rect 513 -645 514 -644
rect 523 -645 524 -644
rect 1024 -645 1025 -644
rect 37 -647 38 -646
rect 86 -647 87 -646
rect 89 -647 90 -646
rect 1178 -647 1179 -646
rect 100 -649 101 -648
rect 467 -649 468 -648
rect 492 -649 493 -648
rect 513 -649 514 -648
rect 541 -649 542 -648
rect 786 -649 787 -648
rect 800 -649 801 -648
rect 870 -649 871 -648
rect 912 -649 913 -648
rect 1003 -649 1004 -648
rect 100 -651 101 -650
rect 390 -651 391 -650
rect 408 -651 409 -650
rect 422 -651 423 -650
rect 478 -651 479 -650
rect 541 -651 542 -650
rect 544 -651 545 -650
rect 751 -651 752 -650
rect 779 -651 780 -650
rect 940 -651 941 -650
rect 947 -651 948 -650
rect 1066 -651 1067 -650
rect 128 -653 129 -652
rect 275 -653 276 -652
rect 289 -653 290 -652
rect 408 -653 409 -652
rect 492 -653 493 -652
rect 660 -653 661 -652
rect 709 -653 710 -652
rect 751 -653 752 -652
rect 807 -653 808 -652
rect 849 -653 850 -652
rect 912 -653 913 -652
rect 926 -653 927 -652
rect 947 -653 948 -652
rect 1017 -653 1018 -652
rect 93 -655 94 -654
rect 128 -655 129 -654
rect 142 -655 143 -654
rect 1143 -655 1144 -654
rect 61 -657 62 -656
rect 142 -657 143 -656
rect 240 -657 241 -656
rect 443 -657 444 -656
rect 502 -657 503 -656
rect 1038 -657 1039 -656
rect 9 -659 10 -658
rect 61 -659 62 -658
rect 93 -659 94 -658
rect 198 -659 199 -658
rect 247 -659 248 -658
rect 282 -659 283 -658
rect 289 -659 290 -658
rect 366 -659 367 -658
rect 394 -659 395 -658
rect 478 -659 479 -658
rect 520 -659 521 -658
rect 800 -659 801 -658
rect 810 -659 811 -658
rect 1087 -659 1088 -658
rect 9 -661 10 -660
rect 369 -661 370 -660
rect 418 -661 419 -660
rect 520 -661 521 -660
rect 548 -661 549 -660
rect 569 -661 570 -660
rect 590 -661 591 -660
rect 611 -661 612 -660
rect 632 -661 633 -660
rect 660 -661 661 -660
rect 709 -661 710 -660
rect 744 -661 745 -660
rect 821 -661 822 -660
rect 919 -661 920 -660
rect 933 -661 934 -660
rect 1017 -661 1018 -660
rect 23 -663 24 -662
rect 366 -663 367 -662
rect 534 -663 535 -662
rect 569 -663 570 -662
rect 576 -663 577 -662
rect 590 -663 591 -662
rect 597 -663 598 -662
rect 625 -663 626 -662
rect 632 -663 633 -662
rect 1115 -663 1116 -662
rect 110 -665 111 -664
rect 394 -665 395 -664
rect 534 -665 535 -664
rect 555 -665 556 -664
rect 558 -665 559 -664
rect 1031 -665 1032 -664
rect 145 -667 146 -666
rect 240 -667 241 -666
rect 261 -667 262 -666
rect 282 -667 283 -666
rect 296 -667 297 -666
rect 436 -667 437 -666
rect 555 -667 556 -666
rect 576 -667 577 -666
rect 597 -667 598 -666
rect 730 -667 731 -666
rect 733 -667 734 -666
rect 1045 -667 1046 -666
rect 198 -669 199 -668
rect 236 -669 237 -668
rect 254 -669 255 -668
rect 261 -669 262 -668
rect 275 -669 276 -668
rect 404 -669 405 -668
rect 562 -669 563 -668
rect 1073 -669 1074 -668
rect 278 -671 279 -670
rect 296 -671 297 -670
rect 303 -671 304 -670
rect 310 -671 311 -670
rect 317 -671 318 -670
rect 331 -671 332 -670
rect 334 -671 335 -670
rect 891 -671 892 -670
rect 954 -671 955 -670
rect 1059 -671 1060 -670
rect 163 -673 164 -672
rect 317 -673 318 -672
rect 457 -673 458 -672
rect 1073 -673 1074 -672
rect 163 -675 164 -674
rect 212 -675 213 -674
rect 268 -675 269 -674
rect 457 -675 458 -674
rect 562 -675 563 -674
rect 758 -675 759 -674
rect 772 -675 773 -674
rect 919 -675 920 -674
rect 968 -675 969 -674
rect 1024 -675 1025 -674
rect 191 -677 192 -676
rect 212 -677 213 -676
rect 219 -677 220 -676
rect 268 -677 269 -676
rect 310 -677 311 -676
rect 485 -677 486 -676
rect 565 -677 566 -676
rect 1136 -677 1137 -676
rect 177 -679 178 -678
rect 191 -679 192 -678
rect 383 -679 384 -678
rect 968 -679 969 -678
rect 177 -681 178 -680
rect 499 -681 500 -680
rect 565 -681 566 -680
rect 1150 -681 1151 -680
rect 149 -683 150 -682
rect 499 -683 500 -682
rect 583 -683 584 -682
rect 772 -683 773 -682
rect 842 -683 843 -682
rect 898 -683 899 -682
rect 149 -685 150 -684
rect 156 -685 157 -684
rect 184 -685 185 -684
rect 219 -685 220 -684
rect 485 -685 486 -684
rect 527 -685 528 -684
rect 583 -685 584 -684
rect 1206 -685 1207 -684
rect 156 -687 157 -686
rect 429 -687 430 -686
rect 506 -687 507 -686
rect 527 -687 528 -686
rect 586 -687 587 -686
rect 758 -687 759 -686
rect 863 -687 864 -686
rect 926 -687 927 -686
rect 72 -689 73 -688
rect 506 -689 507 -688
rect 628 -689 629 -688
rect 842 -689 843 -688
rect 877 -689 878 -688
rect 954 -689 955 -688
rect 72 -691 73 -690
rect 79 -691 80 -690
rect 170 -691 171 -690
rect 184 -691 185 -690
rect 429 -691 430 -690
rect 667 -691 668 -690
rect 695 -691 696 -690
rect 744 -691 745 -690
rect 828 -691 829 -690
rect 863 -691 864 -690
rect 68 -693 69 -692
rect 79 -693 80 -692
rect 114 -693 115 -692
rect 170 -693 171 -692
rect 646 -693 647 -692
rect 933 -693 934 -692
rect 114 -695 115 -694
rect 373 -695 374 -694
rect 681 -695 682 -694
rect 695 -695 696 -694
rect 737 -695 738 -694
rect 779 -695 780 -694
rect 835 -695 836 -694
rect 877 -695 878 -694
rect 373 -697 374 -696
rect 471 -697 472 -696
rect 688 -697 689 -696
rect 828 -697 829 -696
rect 233 -699 234 -698
rect 471 -699 472 -698
rect 653 -699 654 -698
rect 688 -699 689 -698
rect 793 -699 794 -698
rect 835 -699 836 -698
rect 233 -701 234 -700
rect 359 -701 360 -700
rect 383 -701 384 -700
rect 737 -701 738 -700
rect 226 -703 227 -702
rect 359 -703 360 -702
rect 446 -703 447 -702
rect 681 -703 682 -702
rect 254 -705 255 -704
rect 653 -705 654 -704
rect 639 -707 640 -706
rect 793 -707 794 -706
rect 135 -709 136 -708
rect 639 -709 640 -708
rect 135 -711 136 -710
rect 604 -711 605 -710
rect 450 -713 451 -712
rect 604 -713 605 -712
rect 450 -715 451 -714
rect 646 -715 647 -714
rect 2 -726 3 -725
rect 107 -726 108 -725
rect 131 -726 132 -725
rect 310 -726 311 -725
rect 338 -726 339 -725
rect 446 -726 447 -725
rect 464 -726 465 -725
rect 555 -726 556 -725
rect 569 -726 570 -725
rect 572 -726 573 -725
rect 586 -726 587 -725
rect 933 -726 934 -725
rect 1136 -726 1137 -725
rect 1220 -726 1221 -725
rect 1360 -726 1361 -725
rect 1416 -726 1417 -725
rect 2 -728 3 -727
rect 79 -728 80 -727
rect 89 -728 90 -727
rect 194 -728 195 -727
rect 198 -728 199 -727
rect 201 -728 202 -727
rect 254 -728 255 -727
rect 733 -728 734 -727
rect 828 -728 829 -727
rect 1262 -728 1263 -727
rect 9 -730 10 -729
rect 723 -730 724 -729
rect 726 -730 727 -729
rect 1087 -730 1088 -729
rect 1143 -730 1144 -729
rect 1227 -730 1228 -729
rect 9 -732 10 -731
rect 51 -732 52 -731
rect 79 -732 80 -731
rect 240 -732 241 -731
rect 254 -732 255 -731
rect 373 -732 374 -731
rect 390 -732 391 -731
rect 1206 -732 1207 -731
rect 16 -734 17 -733
rect 61 -734 62 -733
rect 89 -734 90 -733
rect 695 -734 696 -733
rect 705 -734 706 -733
rect 1199 -734 1200 -733
rect 16 -736 17 -735
rect 369 -736 370 -735
rect 401 -736 402 -735
rect 989 -736 990 -735
rect 1017 -736 1018 -735
rect 1087 -736 1088 -735
rect 1164 -736 1165 -735
rect 1241 -736 1242 -735
rect 30 -738 31 -737
rect 110 -738 111 -737
rect 156 -738 157 -737
rect 240 -738 241 -737
rect 338 -738 339 -737
rect 408 -738 409 -737
rect 422 -738 423 -737
rect 464 -738 465 -737
rect 485 -738 486 -737
rect 565 -738 566 -737
rect 611 -738 612 -737
rect 632 -738 633 -737
rect 635 -738 636 -737
rect 1150 -738 1151 -737
rect 1178 -738 1179 -737
rect 1248 -738 1249 -737
rect 37 -740 38 -739
rect 380 -740 381 -739
rect 390 -740 391 -739
rect 422 -740 423 -739
rect 436 -740 437 -739
rect 485 -740 486 -739
rect 495 -740 496 -739
rect 534 -740 535 -739
rect 576 -740 577 -739
rect 611 -740 612 -739
rect 646 -740 647 -739
rect 744 -740 745 -739
rect 828 -740 829 -739
rect 1206 -740 1207 -739
rect 37 -742 38 -741
rect 93 -742 94 -741
rect 100 -742 101 -741
rect 558 -742 559 -741
rect 576 -742 577 -741
rect 625 -742 626 -741
rect 649 -742 650 -741
rect 821 -742 822 -741
rect 905 -742 906 -741
rect 933 -742 934 -741
rect 975 -742 976 -741
rect 989 -742 990 -741
rect 1017 -742 1018 -741
rect 1045 -742 1046 -741
rect 1080 -742 1081 -741
rect 1199 -742 1200 -741
rect 51 -744 52 -743
rect 1213 -744 1214 -743
rect 65 -746 66 -745
rect 93 -746 94 -745
rect 100 -746 101 -745
rect 128 -746 129 -745
rect 142 -746 143 -745
rect 156 -746 157 -745
rect 163 -746 164 -745
rect 366 -746 367 -745
rect 380 -746 381 -745
rect 415 -746 416 -745
rect 443 -746 444 -745
rect 1234 -746 1235 -745
rect 65 -748 66 -747
rect 233 -748 234 -747
rect 289 -748 290 -747
rect 443 -748 444 -747
rect 457 -748 458 -747
rect 632 -748 633 -747
rect 649 -748 650 -747
rect 1171 -748 1172 -747
rect 1185 -748 1186 -747
rect 1255 -748 1256 -747
rect 86 -750 87 -749
rect 1080 -750 1081 -749
rect 1094 -750 1095 -749
rect 1150 -750 1151 -749
rect 1157 -750 1158 -749
rect 1185 -750 1186 -749
rect 107 -752 108 -751
rect 149 -752 150 -751
rect 170 -752 171 -751
rect 173 -752 174 -751
rect 177 -752 178 -751
rect 534 -752 535 -751
rect 590 -752 591 -751
rect 975 -752 976 -751
rect 1101 -752 1102 -751
rect 1178 -752 1179 -751
rect 142 -754 143 -753
rect 387 -754 388 -753
rect 408 -754 409 -753
rect 478 -754 479 -753
rect 502 -754 503 -753
rect 996 -754 997 -753
rect 1108 -754 1109 -753
rect 1171 -754 1172 -753
rect 149 -756 150 -755
rect 513 -756 514 -755
rect 516 -756 517 -755
rect 695 -756 696 -755
rect 709 -756 710 -755
rect 744 -756 745 -755
rect 856 -756 857 -755
rect 905 -756 906 -755
rect 912 -756 913 -755
rect 1045 -756 1046 -755
rect 1115 -756 1116 -755
rect 1164 -756 1165 -755
rect 170 -758 171 -757
rect 205 -758 206 -757
rect 212 -758 213 -757
rect 233 -758 234 -757
rect 299 -758 300 -757
rect 821 -758 822 -757
rect 856 -758 857 -757
rect 968 -758 969 -757
rect 1059 -758 1060 -757
rect 1115 -758 1116 -757
rect 1122 -758 1123 -757
rect 1213 -758 1214 -757
rect 44 -760 45 -759
rect 968 -760 969 -759
rect 44 -762 45 -761
rect 383 -762 384 -761
rect 415 -762 416 -761
rect 681 -762 682 -761
rect 709 -762 710 -761
rect 716 -762 717 -761
rect 723 -762 724 -761
rect 751 -762 752 -761
rect 765 -762 766 -761
rect 912 -762 913 -761
rect 961 -762 962 -761
rect 1094 -762 1095 -761
rect 33 -764 34 -763
rect 751 -764 752 -763
rect 765 -764 766 -763
rect 1052 -764 1053 -763
rect 114 -766 115 -765
rect 681 -766 682 -765
rect 702 -766 703 -765
rect 716 -766 717 -765
rect 730 -766 731 -765
rect 1010 -766 1011 -765
rect 114 -768 115 -767
rect 499 -768 500 -767
rect 506 -768 507 -767
rect 625 -768 626 -767
rect 639 -768 640 -767
rect 1157 -768 1158 -767
rect 128 -770 129 -769
rect 1059 -770 1060 -769
rect 135 -772 136 -771
rect 639 -772 640 -771
rect 653 -772 654 -771
rect 1143 -772 1144 -771
rect 75 -774 76 -773
rect 135 -774 136 -773
rect 191 -774 192 -773
rect 212 -774 213 -773
rect 352 -774 353 -773
rect 404 -774 405 -773
rect 457 -774 458 -773
rect 506 -774 507 -773
rect 513 -774 514 -773
rect 1192 -774 1193 -773
rect 121 -776 122 -775
rect 191 -776 192 -775
rect 198 -776 199 -775
rect 219 -776 220 -775
rect 359 -776 360 -775
rect 373 -776 374 -775
rect 478 -776 479 -775
rect 597 -776 598 -775
rect 656 -776 657 -775
rect 1129 -776 1130 -775
rect 121 -778 122 -777
rect 761 -778 762 -777
rect 870 -778 871 -777
rect 996 -778 997 -777
rect 1024 -778 1025 -777
rect 1129 -778 1130 -777
rect 177 -780 178 -779
rect 352 -780 353 -779
rect 359 -780 360 -779
rect 397 -780 398 -779
rect 432 -780 433 -779
rect 1024 -780 1025 -779
rect 205 -782 206 -781
rect 345 -782 346 -781
rect 366 -782 367 -781
rect 450 -782 451 -781
rect 492 -782 493 -781
rect 1108 -782 1109 -781
rect 184 -784 185 -783
rect 345 -784 346 -783
rect 492 -784 493 -783
rect 793 -784 794 -783
rect 870 -784 871 -783
rect 940 -784 941 -783
rect 947 -784 948 -783
rect 1192 -784 1193 -783
rect 184 -786 185 -785
rect 303 -786 304 -785
rect 520 -786 521 -785
rect 565 -786 566 -785
rect 569 -786 570 -785
rect 1101 -786 1102 -785
rect 23 -788 24 -787
rect 520 -788 521 -787
rect 523 -788 524 -787
rect 919 -788 920 -787
rect 926 -788 927 -787
rect 940 -788 941 -787
rect 954 -788 955 -787
rect 1010 -788 1011 -787
rect 219 -790 220 -789
rect 261 -790 262 -789
rect 275 -790 276 -789
rect 450 -790 451 -789
rect 527 -790 528 -789
rect 954 -790 955 -789
rect 961 -790 962 -789
rect 1003 -790 1004 -789
rect 261 -792 262 -791
rect 282 -792 283 -791
rect 527 -792 528 -791
rect 786 -792 787 -791
rect 877 -792 878 -791
rect 926 -792 927 -791
rect 201 -794 202 -793
rect 282 -794 283 -793
rect 583 -794 584 -793
rect 947 -794 948 -793
rect 268 -796 269 -795
rect 275 -796 276 -795
rect 499 -796 500 -795
rect 583 -796 584 -795
rect 586 -796 587 -795
rect 1122 -796 1123 -795
rect 268 -798 269 -797
rect 394 -798 395 -797
rect 590 -798 591 -797
rect 618 -798 619 -797
rect 653 -798 654 -797
rect 793 -798 794 -797
rect 849 -798 850 -797
rect 877 -798 878 -797
rect 898 -798 899 -797
rect 1003 -798 1004 -797
rect 163 -800 164 -799
rect 618 -800 619 -799
rect 656 -800 657 -799
rect 1052 -800 1053 -799
rect 387 -802 388 -801
rect 394 -802 395 -801
rect 429 -802 430 -801
rect 898 -802 899 -801
rect 919 -802 920 -801
rect 982 -802 983 -801
rect 429 -804 430 -803
rect 1136 -804 1137 -803
rect 597 -806 598 -805
rect 674 -806 675 -805
rect 688 -806 689 -805
rect 786 -806 787 -805
rect 814 -806 815 -805
rect 849 -806 850 -805
rect 884 -806 885 -805
rect 982 -806 983 -805
rect 58 -808 59 -807
rect 688 -808 689 -807
rect 702 -808 703 -807
rect 891 -808 892 -807
rect 58 -810 59 -809
rect 72 -810 73 -809
rect 404 -810 405 -809
rect 674 -810 675 -809
rect 779 -810 780 -809
rect 891 -810 892 -809
rect 72 -812 73 -811
rect 289 -812 290 -811
rect 471 -812 472 -811
rect 779 -812 780 -811
rect 800 -812 801 -811
rect 814 -812 815 -811
rect 863 -812 864 -811
rect 884 -812 885 -811
rect 317 -814 318 -813
rect 471 -814 472 -813
rect 604 -814 605 -813
rect 800 -814 801 -813
rect 842 -814 843 -813
rect 863 -814 864 -813
rect 226 -816 227 -815
rect 317 -816 318 -815
rect 548 -816 549 -815
rect 604 -816 605 -815
rect 667 -816 668 -815
rect 730 -816 731 -815
rect 835 -816 836 -815
rect 842 -816 843 -815
rect 226 -818 227 -817
rect 247 -818 248 -817
rect 541 -818 542 -817
rect 548 -818 549 -817
rect 660 -818 661 -817
rect 667 -818 668 -817
rect 807 -818 808 -817
rect 835 -818 836 -817
rect 247 -820 248 -819
rect 324 -820 325 -819
rect 509 -820 510 -819
rect 541 -820 542 -819
rect 562 -820 563 -819
rect 660 -820 661 -819
rect 758 -820 759 -819
rect 807 -820 808 -819
rect 324 -822 325 -821
rect 331 -822 332 -821
rect 562 -822 563 -821
rect 621 -822 622 -821
rect 758 -822 759 -821
rect 1066 -822 1067 -821
rect 296 -824 297 -823
rect 331 -824 332 -823
rect 1031 -824 1032 -823
rect 1066 -824 1067 -823
rect 296 -826 297 -825
rect 1073 -826 1074 -825
rect 432 -828 433 -827
rect 1031 -828 1032 -827
rect 1038 -828 1039 -827
rect 1073 -828 1074 -827
rect 772 -830 773 -829
rect 1038 -830 1039 -829
rect 310 -832 311 -831
rect 772 -832 773 -831
rect 16 -843 17 -842
rect 635 -843 636 -842
rect 649 -843 650 -842
rect 779 -843 780 -842
rect 824 -843 825 -842
rect 1248 -843 1249 -842
rect 1416 -843 1417 -842
rect 1437 -843 1438 -842
rect 16 -845 17 -844
rect 58 -845 59 -844
rect 68 -845 69 -844
rect 338 -845 339 -844
rect 390 -845 391 -844
rect 898 -845 899 -844
rect 961 -845 962 -844
rect 964 -845 965 -844
rect 26 -847 27 -846
rect 44 -847 45 -846
rect 58 -847 59 -846
rect 163 -847 164 -846
rect 170 -847 171 -846
rect 432 -847 433 -846
rect 439 -847 440 -846
rect 1136 -847 1137 -846
rect 30 -849 31 -848
rect 93 -849 94 -848
rect 124 -849 125 -848
rect 1143 -849 1144 -848
rect 30 -851 31 -850
rect 415 -851 416 -850
rect 425 -851 426 -850
rect 786 -851 787 -850
rect 828 -851 829 -850
rect 1220 -851 1221 -850
rect 33 -853 34 -852
rect 947 -853 948 -852
rect 961 -853 962 -852
rect 989 -853 990 -852
rect 1143 -853 1144 -852
rect 1199 -853 1200 -852
rect 37 -855 38 -854
rect 520 -855 521 -854
rect 537 -855 538 -854
rect 576 -855 577 -854
rect 586 -855 587 -854
rect 1010 -855 1011 -854
rect 1129 -855 1130 -854
rect 1199 -855 1200 -854
rect 37 -857 38 -856
rect 51 -857 52 -856
rect 72 -857 73 -856
rect 184 -857 185 -856
rect 198 -857 199 -856
rect 401 -857 402 -856
rect 443 -857 444 -856
rect 516 -857 517 -856
rect 544 -857 545 -856
rect 625 -857 626 -856
rect 653 -857 654 -856
rect 891 -857 892 -856
rect 898 -857 899 -856
rect 940 -857 941 -856
rect 947 -857 948 -856
rect 968 -857 969 -856
rect 1010 -857 1011 -856
rect 1052 -857 1053 -856
rect 44 -859 45 -858
rect 737 -859 738 -858
rect 758 -859 759 -858
rect 1227 -859 1228 -858
rect 51 -861 52 -860
rect 201 -861 202 -860
rect 205 -861 206 -860
rect 583 -861 584 -860
rect 618 -861 619 -860
rect 1003 -861 1004 -860
rect 1052 -861 1053 -860
rect 1202 -861 1203 -860
rect 65 -863 66 -862
rect 72 -863 73 -862
rect 79 -863 80 -862
rect 583 -863 584 -862
rect 611 -863 612 -862
rect 618 -863 619 -862
rect 625 -863 626 -862
rect 1171 -863 1172 -862
rect 65 -865 66 -864
rect 100 -865 101 -864
rect 121 -865 122 -864
rect 415 -865 416 -864
rect 443 -865 444 -864
rect 695 -865 696 -864
rect 702 -865 703 -864
rect 1038 -865 1039 -864
rect 1164 -865 1165 -864
rect 1171 -865 1172 -864
rect 79 -867 80 -866
rect 478 -867 479 -866
rect 485 -867 486 -866
rect 520 -867 521 -866
rect 565 -867 566 -866
rect 1087 -867 1088 -866
rect 86 -869 87 -868
rect 828 -869 829 -868
rect 856 -869 857 -868
rect 940 -869 941 -868
rect 964 -869 965 -868
rect 989 -869 990 -868
rect 1003 -869 1004 -868
rect 1045 -869 1046 -868
rect 1059 -869 1060 -868
rect 1164 -869 1165 -868
rect 9 -871 10 -870
rect 86 -871 87 -870
rect 89 -871 90 -870
rect 303 -871 304 -870
rect 380 -871 381 -870
rect 401 -871 402 -870
rect 471 -871 472 -870
rect 485 -871 486 -870
rect 506 -871 507 -870
rect 954 -871 955 -870
rect 968 -871 969 -870
rect 1073 -871 1074 -870
rect 1087 -871 1088 -870
rect 1122 -871 1123 -870
rect 2 -873 3 -872
rect 303 -873 304 -872
rect 331 -873 332 -872
rect 380 -873 381 -872
rect 397 -873 398 -872
rect 1157 -873 1158 -872
rect 23 -875 24 -874
rect 856 -875 857 -874
rect 982 -875 983 -874
rect 1122 -875 1123 -874
rect 23 -877 24 -876
rect 495 -877 496 -876
rect 509 -877 510 -876
rect 660 -877 661 -876
rect 674 -877 675 -876
rect 1059 -877 1060 -876
rect 93 -879 94 -878
rect 215 -879 216 -878
rect 240 -879 241 -878
rect 394 -879 395 -878
rect 408 -879 409 -878
rect 506 -879 507 -878
rect 569 -879 570 -878
rect 1178 -879 1179 -878
rect 100 -881 101 -880
rect 499 -881 500 -880
rect 572 -881 573 -880
rect 758 -881 759 -880
rect 761 -881 762 -880
rect 954 -881 955 -880
rect 1017 -881 1018 -880
rect 1045 -881 1046 -880
rect 121 -883 122 -882
rect 674 -883 675 -882
rect 688 -883 689 -882
rect 1129 -883 1130 -882
rect 131 -885 132 -884
rect 1178 -885 1179 -884
rect 152 -887 153 -886
rect 982 -887 983 -886
rect 1017 -887 1018 -886
rect 1066 -887 1067 -886
rect 156 -889 157 -888
rect 331 -889 332 -888
rect 369 -889 370 -888
rect 394 -889 395 -888
rect 422 -889 423 -888
rect 471 -889 472 -888
rect 478 -889 479 -888
rect 912 -889 913 -888
rect 1031 -889 1032 -888
rect 1038 -889 1039 -888
rect 2 -891 3 -890
rect 422 -891 423 -890
rect 499 -891 500 -890
rect 975 -891 976 -890
rect 1031 -891 1032 -890
rect 1080 -891 1081 -890
rect 156 -893 157 -892
rect 712 -893 713 -892
rect 723 -893 724 -892
rect 737 -893 738 -892
rect 765 -893 766 -892
rect 1066 -893 1067 -892
rect 1080 -893 1081 -892
rect 1115 -893 1116 -892
rect 89 -895 90 -894
rect 1115 -895 1116 -894
rect 131 -897 132 -896
rect 723 -897 724 -896
rect 730 -897 731 -896
rect 779 -897 780 -896
rect 786 -897 787 -896
rect 863 -897 864 -896
rect 919 -897 920 -896
rect 975 -897 976 -896
rect 163 -899 164 -898
rect 191 -899 192 -898
rect 198 -899 199 -898
rect 240 -899 241 -898
rect 254 -899 255 -898
rect 387 -899 388 -898
rect 611 -899 612 -898
rect 1192 -899 1193 -898
rect 114 -901 115 -900
rect 191 -901 192 -900
rect 205 -901 206 -900
rect 289 -901 290 -900
rect 296 -901 297 -900
rect 345 -901 346 -900
rect 632 -901 633 -900
rect 660 -901 661 -900
rect 695 -901 696 -900
rect 716 -901 717 -900
rect 765 -901 766 -900
rect 800 -901 801 -900
rect 807 -901 808 -900
rect 891 -901 892 -900
rect 919 -901 920 -900
rect 926 -901 927 -900
rect 1094 -901 1095 -900
rect 1192 -901 1193 -900
rect 107 -903 108 -902
rect 114 -903 115 -902
rect 170 -903 171 -902
rect 404 -903 405 -902
rect 569 -903 570 -902
rect 632 -903 633 -902
rect 646 -903 647 -902
rect 1073 -903 1074 -902
rect 1094 -903 1095 -902
rect 1150 -903 1151 -902
rect 107 -905 108 -904
rect 359 -905 360 -904
rect 590 -905 591 -904
rect 646 -905 647 -904
rect 653 -905 654 -904
rect 996 -905 997 -904
rect 1150 -905 1151 -904
rect 1206 -905 1207 -904
rect 177 -907 178 -906
rect 275 -907 276 -906
rect 282 -907 283 -906
rect 320 -907 321 -906
rect 345 -907 346 -906
rect 562 -907 563 -906
rect 614 -907 615 -906
rect 926 -907 927 -906
rect 996 -907 997 -906
rect 1024 -907 1025 -906
rect 1185 -907 1186 -906
rect 1206 -907 1207 -906
rect 180 -909 181 -908
rect 681 -909 682 -908
rect 702 -909 703 -908
rect 842 -909 843 -908
rect 863 -909 864 -908
rect 933 -909 934 -908
rect 1024 -909 1025 -908
rect 1101 -909 1102 -908
rect 1185 -909 1186 -908
rect 1234 -909 1235 -908
rect 184 -911 185 -910
rect 691 -911 692 -910
rect 709 -911 710 -910
rect 730 -911 731 -910
rect 751 -911 752 -910
rect 800 -911 801 -910
rect 807 -911 808 -910
rect 814 -911 815 -910
rect 870 -911 871 -910
rect 933 -911 934 -910
rect 212 -913 213 -912
rect 359 -913 360 -912
rect 513 -913 514 -912
rect 814 -913 815 -912
rect 870 -913 871 -912
rect 1262 -913 1263 -912
rect 212 -915 213 -914
rect 429 -915 430 -914
rect 555 -915 556 -914
rect 590 -915 591 -914
rect 656 -915 657 -914
rect 905 -915 906 -914
rect 219 -917 220 -916
rect 296 -917 297 -916
rect 299 -917 300 -916
rect 387 -917 388 -916
rect 450 -917 451 -916
rect 555 -917 556 -916
rect 562 -917 563 -916
rect 747 -917 748 -916
rect 772 -917 773 -916
rect 1241 -917 1242 -916
rect 219 -919 220 -918
rect 502 -919 503 -918
rect 527 -919 528 -918
rect 772 -919 773 -918
rect 775 -919 776 -918
rect 842 -919 843 -918
rect 247 -921 248 -920
rect 254 -921 255 -920
rect 261 -921 262 -920
rect 275 -921 276 -920
rect 282 -921 283 -920
rect 436 -921 437 -920
rect 450 -921 451 -920
rect 1136 -921 1137 -920
rect 247 -923 248 -922
rect 831 -923 832 -922
rect 261 -925 262 -924
rect 366 -925 367 -924
rect 373 -925 374 -924
rect 513 -925 514 -924
rect 576 -925 577 -924
rect 656 -925 657 -924
rect 667 -925 668 -924
rect 681 -925 682 -924
rect 709 -925 710 -924
rect 1255 -925 1256 -924
rect 226 -927 227 -926
rect 366 -927 367 -926
rect 436 -927 437 -926
rect 541 -927 542 -926
rect 597 -927 598 -926
rect 905 -927 906 -926
rect 135 -929 136 -928
rect 226 -929 227 -928
rect 268 -929 269 -928
rect 338 -929 339 -928
rect 352 -929 353 -928
rect 429 -929 430 -928
rect 541 -929 542 -928
rect 849 -929 850 -928
rect 135 -931 136 -930
rect 492 -931 493 -930
rect 548 -931 549 -930
rect 597 -931 598 -930
rect 639 -931 640 -930
rect 667 -931 668 -930
rect 716 -931 717 -930
rect 1108 -931 1109 -930
rect 142 -933 143 -932
rect 352 -933 353 -932
rect 457 -933 458 -932
rect 548 -933 549 -932
rect 604 -933 605 -932
rect 639 -933 640 -932
rect 688 -933 689 -932
rect 1108 -933 1109 -932
rect 142 -935 143 -934
rect 705 -935 706 -934
rect 719 -935 720 -934
rect 1101 -935 1102 -934
rect 149 -937 150 -936
rect 492 -937 493 -936
rect 534 -937 535 -936
rect 604 -937 605 -936
rect 744 -937 745 -936
rect 751 -937 752 -936
rect 793 -937 794 -936
rect 912 -937 913 -936
rect 268 -939 269 -938
rect 481 -939 482 -938
rect 534 -939 535 -938
rect 1157 -939 1158 -938
rect 289 -941 290 -940
rect 324 -941 325 -940
rect 457 -941 458 -940
rect 464 -941 465 -940
rect 793 -941 794 -940
rect 835 -941 836 -940
rect 849 -941 850 -940
rect 877 -941 878 -940
rect 310 -943 311 -942
rect 373 -943 374 -942
rect 464 -943 465 -942
rect 523 -943 524 -942
rect 821 -943 822 -942
rect 835 -943 836 -942
rect 877 -943 878 -942
rect 884 -943 885 -942
rect 75 -945 76 -944
rect 310 -945 311 -944
rect 317 -945 318 -944
rect 408 -945 409 -944
rect 821 -945 822 -944
rect 1213 -945 1214 -944
rect 9 -947 10 -946
rect 317 -947 318 -946
rect 324 -947 325 -946
rect 628 -947 629 -946
rect 128 -949 129 -948
rect 884 -949 885 -948
rect 2 -960 3 -959
rect 149 -960 150 -959
rect 152 -960 153 -959
rect 439 -960 440 -959
rect 502 -960 503 -959
rect 681 -960 682 -959
rect 688 -960 689 -959
rect 919 -960 920 -959
rect 929 -960 930 -959
rect 1325 -960 1326 -959
rect 1437 -960 1438 -959
rect 1444 -960 1445 -959
rect 5 -962 6 -961
rect 408 -962 409 -961
rect 541 -962 542 -961
rect 1262 -962 1263 -961
rect 9 -964 10 -963
rect 422 -964 423 -963
rect 548 -964 549 -963
rect 712 -964 713 -963
rect 719 -964 720 -963
rect 1290 -964 1291 -963
rect 16 -966 17 -965
rect 89 -966 90 -965
rect 103 -966 104 -965
rect 716 -966 717 -965
rect 744 -966 745 -965
rect 1122 -966 1123 -965
rect 1136 -966 1137 -965
rect 1269 -966 1270 -965
rect 16 -968 17 -967
rect 534 -968 535 -967
rect 558 -968 559 -967
rect 786 -968 787 -967
rect 863 -968 864 -967
rect 1136 -968 1137 -967
rect 1143 -968 1144 -967
rect 1304 -968 1305 -967
rect 30 -970 31 -969
rect 537 -970 538 -969
rect 565 -970 566 -969
rect 1059 -970 1060 -969
rect 1073 -970 1074 -969
rect 1220 -970 1221 -969
rect 2 -972 3 -971
rect 30 -972 31 -971
rect 33 -972 34 -971
rect 772 -972 773 -971
rect 866 -972 867 -971
rect 968 -972 969 -971
rect 1087 -972 1088 -971
rect 1213 -972 1214 -971
rect 44 -974 45 -973
rect 317 -974 318 -973
rect 320 -974 321 -973
rect 422 -974 423 -973
rect 502 -974 503 -973
rect 786 -974 787 -973
rect 877 -974 878 -973
rect 1122 -974 1123 -973
rect 1157 -974 1158 -973
rect 1311 -974 1312 -973
rect 44 -976 45 -975
rect 170 -976 171 -975
rect 201 -976 202 -975
rect 387 -976 388 -975
rect 611 -976 612 -975
rect 1276 -976 1277 -975
rect 37 -978 38 -977
rect 170 -978 171 -977
rect 212 -978 213 -977
rect 726 -978 727 -977
rect 744 -978 745 -977
rect 863 -978 864 -977
rect 870 -978 871 -977
rect 877 -978 878 -977
rect 912 -978 913 -977
rect 919 -978 920 -977
rect 954 -978 955 -977
rect 1073 -978 1074 -977
rect 1094 -978 1095 -977
rect 1248 -978 1249 -977
rect 75 -980 76 -979
rect 660 -980 661 -979
rect 667 -980 668 -979
rect 772 -980 773 -979
rect 849 -980 850 -979
rect 954 -980 955 -979
rect 961 -980 962 -979
rect 1255 -980 1256 -979
rect 51 -982 52 -981
rect 660 -982 661 -981
rect 695 -982 696 -981
rect 1297 -982 1298 -981
rect 51 -984 52 -983
rect 884 -984 885 -983
rect 968 -984 969 -983
rect 1010 -984 1011 -983
rect 1052 -984 1053 -983
rect 1094 -984 1095 -983
rect 1101 -984 1102 -983
rect 1234 -984 1235 -983
rect 79 -986 80 -985
rect 450 -986 451 -985
rect 572 -986 573 -985
rect 870 -986 871 -985
rect 884 -986 885 -985
rect 940 -986 941 -985
rect 975 -986 976 -985
rect 1087 -986 1088 -985
rect 1115 -986 1116 -985
rect 1241 -986 1242 -985
rect 23 -988 24 -987
rect 450 -988 451 -987
rect 576 -988 577 -987
rect 912 -988 913 -987
rect 933 -988 934 -987
rect 1052 -988 1053 -987
rect 1150 -988 1151 -987
rect 1157 -988 1158 -987
rect 1164 -988 1165 -987
rect 1318 -988 1319 -987
rect 23 -990 24 -989
rect 268 -990 269 -989
rect 282 -990 283 -989
rect 425 -990 426 -989
rect 436 -990 437 -989
rect 695 -990 696 -989
rect 702 -990 703 -989
rect 933 -990 934 -989
rect 1003 -990 1004 -989
rect 1115 -990 1116 -989
rect 1185 -990 1186 -989
rect 1339 -990 1340 -989
rect 79 -992 80 -991
rect 219 -992 220 -991
rect 254 -992 255 -991
rect 614 -992 615 -991
rect 618 -992 619 -991
rect 688 -992 689 -991
rect 709 -992 710 -991
rect 1059 -992 1060 -991
rect 1192 -992 1193 -991
rect 1206 -992 1207 -991
rect 114 -994 115 -993
rect 131 -994 132 -993
rect 149 -994 150 -993
rect 408 -994 409 -993
rect 436 -994 437 -993
rect 576 -994 577 -993
rect 611 -994 612 -993
rect 821 -994 822 -993
rect 856 -994 857 -993
rect 1101 -994 1102 -993
rect 96 -996 97 -995
rect 114 -996 115 -995
rect 124 -996 125 -995
rect 653 -996 654 -995
rect 723 -996 724 -995
rect 940 -996 941 -995
rect 1017 -996 1018 -995
rect 1150 -996 1151 -995
rect 177 -998 178 -997
rect 254 -998 255 -997
rect 264 -998 265 -997
rect 478 -998 479 -997
rect 499 -998 500 -997
rect 856 -998 857 -997
rect 891 -998 892 -997
rect 975 -998 976 -997
rect 982 -998 983 -997
rect 1017 -998 1018 -997
rect 1045 -998 1046 -997
rect 1185 -998 1186 -997
rect 177 -1000 178 -999
rect 240 -1000 241 -999
rect 268 -1000 269 -999
rect 453 -1000 454 -999
rect 471 -1000 472 -999
rect 982 -1000 983 -999
rect 1066 -1000 1067 -999
rect 1192 -1000 1193 -999
rect 205 -1002 206 -1001
rect 212 -1002 213 -1001
rect 219 -1002 220 -1001
rect 1195 -1002 1196 -1001
rect 240 -1004 241 -1003
rect 324 -1004 325 -1003
rect 338 -1004 339 -1003
rect 387 -1004 388 -1003
rect 471 -1004 472 -1003
rect 506 -1004 507 -1003
rect 513 -1004 514 -1003
rect 653 -1004 654 -1003
rect 723 -1004 724 -1003
rect 961 -1004 962 -1003
rect 1080 -1004 1081 -1003
rect 1206 -1004 1207 -1003
rect 282 -1006 283 -1005
rect 415 -1006 416 -1005
rect 478 -1006 479 -1005
rect 1108 -1006 1109 -1005
rect 289 -1008 290 -1007
rect 324 -1008 325 -1007
rect 341 -1008 342 -1007
rect 401 -1008 402 -1007
rect 499 -1008 500 -1007
rect 548 -1008 549 -1007
rect 555 -1008 556 -1007
rect 618 -1008 619 -1007
rect 628 -1008 629 -1007
rect 737 -1008 738 -1007
rect 747 -1008 748 -1007
rect 779 -1008 780 -1007
rect 800 -1008 801 -1007
rect 821 -1008 822 -1007
rect 835 -1008 836 -1007
rect 891 -1008 892 -1007
rect 926 -1008 927 -1007
rect 1045 -1008 1046 -1007
rect 1080 -1008 1081 -1007
rect 1129 -1008 1130 -1007
rect 128 -1010 129 -1009
rect 737 -1010 738 -1009
rect 747 -1010 748 -1009
rect 1227 -1010 1228 -1009
rect 37 -1012 38 -1011
rect 128 -1012 129 -1011
rect 142 -1012 143 -1011
rect 289 -1012 290 -1011
rect 303 -1012 304 -1011
rect 415 -1012 416 -1011
rect 506 -1012 507 -1011
rect 562 -1012 563 -1011
rect 632 -1012 633 -1011
rect 1332 -1012 1333 -1011
rect 86 -1014 87 -1013
rect 303 -1014 304 -1013
rect 306 -1014 307 -1013
rect 310 -1014 311 -1013
rect 317 -1014 318 -1013
rect 481 -1014 482 -1013
rect 513 -1014 514 -1013
rect 646 -1014 647 -1013
rect 656 -1014 657 -1013
rect 800 -1014 801 -1013
rect 814 -1014 815 -1013
rect 849 -1014 850 -1013
rect 996 -1014 997 -1013
rect 1108 -1014 1109 -1013
rect 86 -1016 87 -1015
rect 544 -1016 545 -1015
rect 597 -1016 598 -1015
rect 646 -1016 647 -1015
rect 751 -1016 752 -1015
rect 779 -1016 780 -1015
rect 807 -1016 808 -1015
rect 814 -1016 815 -1015
rect 989 -1016 990 -1015
rect 996 -1016 997 -1015
rect 1031 -1016 1032 -1015
rect 1129 -1016 1130 -1015
rect 40 -1018 41 -1017
rect 597 -1018 598 -1017
rect 635 -1018 636 -1017
rect 1346 -1018 1347 -1017
rect 310 -1020 311 -1019
rect 338 -1020 339 -1019
rect 345 -1020 346 -1019
rect 702 -1020 703 -1019
rect 730 -1020 731 -1019
rect 751 -1020 752 -1019
rect 758 -1020 759 -1019
rect 1003 -1020 1004 -1019
rect 345 -1022 346 -1021
rect 373 -1022 374 -1021
rect 376 -1022 377 -1021
rect 1178 -1022 1179 -1021
rect 352 -1024 353 -1023
rect 530 -1024 531 -1023
rect 569 -1024 570 -1023
rect 758 -1024 759 -1023
rect 765 -1024 766 -1023
rect 1143 -1024 1144 -1023
rect 9 -1026 10 -1025
rect 530 -1026 531 -1025
rect 569 -1026 570 -1025
rect 604 -1026 605 -1025
rect 639 -1026 640 -1025
rect 681 -1026 682 -1025
rect 793 -1026 794 -1025
rect 989 -1026 990 -1025
rect 1024 -1026 1025 -1025
rect 1178 -1026 1179 -1025
rect 261 -1028 262 -1027
rect 352 -1028 353 -1027
rect 359 -1028 360 -1027
rect 667 -1028 668 -1027
rect 677 -1028 678 -1027
rect 765 -1028 766 -1027
rect 793 -1028 794 -1027
rect 824 -1028 825 -1027
rect 898 -1028 899 -1027
rect 1024 -1028 1025 -1027
rect 68 -1030 69 -1029
rect 898 -1030 899 -1029
rect 905 -1030 906 -1029
rect 1031 -1030 1032 -1029
rect 107 -1032 108 -1031
rect 359 -1032 360 -1031
rect 366 -1032 367 -1031
rect 1010 -1032 1011 -1031
rect 107 -1034 108 -1033
rect 625 -1034 626 -1033
rect 842 -1034 843 -1033
rect 905 -1034 906 -1033
rect 100 -1036 101 -1035
rect 842 -1036 843 -1035
rect 100 -1038 101 -1037
rect 1038 -1038 1039 -1037
rect 296 -1040 297 -1039
rect 639 -1040 640 -1039
rect 947 -1040 948 -1039
rect 1038 -1040 1039 -1039
rect 135 -1042 136 -1041
rect 296 -1042 297 -1041
rect 366 -1042 367 -1041
rect 1199 -1042 1200 -1041
rect 65 -1044 66 -1043
rect 135 -1044 136 -1043
rect 369 -1044 370 -1043
rect 1283 -1044 1284 -1043
rect 65 -1046 66 -1045
rect 495 -1046 496 -1045
rect 520 -1046 521 -1045
rect 1066 -1046 1067 -1045
rect 373 -1048 374 -1047
rect 394 -1048 395 -1047
rect 401 -1048 402 -1047
rect 457 -1048 458 -1047
rect 464 -1048 465 -1047
rect 730 -1048 731 -1047
rect 828 -1048 829 -1047
rect 947 -1048 948 -1047
rect 191 -1050 192 -1049
rect 394 -1050 395 -1049
rect 429 -1050 430 -1049
rect 457 -1050 458 -1049
rect 481 -1050 482 -1049
rect 1199 -1050 1200 -1049
rect 163 -1052 164 -1051
rect 191 -1052 192 -1051
rect 261 -1052 262 -1051
rect 464 -1052 465 -1051
rect 492 -1052 493 -1051
rect 520 -1052 521 -1051
rect 527 -1052 528 -1051
rect 1164 -1052 1165 -1051
rect 163 -1054 164 -1053
rect 926 -1054 927 -1053
rect 184 -1056 185 -1055
rect 429 -1056 430 -1055
rect 492 -1056 493 -1055
rect 835 -1056 836 -1055
rect 184 -1058 185 -1057
rect 247 -1058 248 -1057
rect 380 -1058 381 -1057
rect 541 -1058 542 -1057
rect 583 -1058 584 -1057
rect 807 -1058 808 -1057
rect 233 -1060 234 -1059
rect 247 -1060 248 -1059
rect 380 -1060 381 -1059
rect 516 -1060 517 -1059
rect 527 -1060 528 -1059
rect 709 -1060 710 -1059
rect 54 -1062 55 -1061
rect 233 -1062 234 -1061
rect 534 -1062 535 -1061
rect 625 -1062 626 -1061
rect 674 -1062 675 -1061
rect 828 -1062 829 -1061
rect 443 -1064 444 -1063
rect 674 -1064 675 -1063
rect 93 -1066 94 -1065
rect 443 -1066 444 -1065
rect 583 -1066 584 -1065
rect 635 -1066 636 -1065
rect 93 -1068 94 -1067
rect 142 -1068 143 -1067
rect 590 -1068 591 -1067
rect 604 -1068 605 -1067
rect 226 -1070 227 -1069
rect 590 -1070 591 -1069
rect 226 -1072 227 -1071
rect 275 -1072 276 -1071
rect 58 -1074 59 -1073
rect 275 -1074 276 -1073
rect 58 -1076 59 -1075
rect 72 -1076 73 -1075
rect 72 -1078 73 -1077
rect 205 -1078 206 -1077
rect 2 -1089 3 -1088
rect 982 -1089 983 -1088
rect 1241 -1089 1242 -1088
rect 1367 -1089 1368 -1088
rect 1444 -1089 1445 -1088
rect 1451 -1089 1452 -1088
rect 9 -1091 10 -1090
rect 338 -1091 339 -1090
rect 404 -1091 405 -1090
rect 667 -1091 668 -1090
rect 674 -1091 675 -1090
rect 1269 -1091 1270 -1090
rect 1318 -1091 1319 -1090
rect 1353 -1091 1354 -1090
rect 9 -1093 10 -1092
rect 33 -1093 34 -1092
rect 37 -1093 38 -1092
rect 121 -1093 122 -1092
rect 149 -1093 150 -1092
rect 226 -1093 227 -1092
rect 247 -1093 248 -1092
rect 264 -1093 265 -1092
rect 439 -1093 440 -1092
rect 520 -1093 521 -1092
rect 527 -1093 528 -1092
rect 1143 -1093 1144 -1092
rect 1213 -1093 1214 -1092
rect 1241 -1093 1242 -1092
rect 1325 -1093 1326 -1092
rect 1360 -1093 1361 -1092
rect 30 -1095 31 -1094
rect 562 -1095 563 -1094
rect 569 -1095 570 -1094
rect 1318 -1095 1319 -1094
rect 1339 -1095 1340 -1094
rect 1374 -1095 1375 -1094
rect 54 -1097 55 -1096
rect 842 -1097 843 -1096
rect 845 -1097 846 -1096
rect 982 -1097 983 -1096
rect 1220 -1097 1221 -1096
rect 1269 -1097 1270 -1096
rect 1311 -1097 1312 -1096
rect 1339 -1097 1340 -1096
rect 58 -1099 59 -1098
rect 100 -1099 101 -1098
rect 121 -1099 122 -1098
rect 289 -1099 290 -1098
rect 408 -1099 409 -1098
rect 562 -1099 563 -1098
rect 572 -1099 573 -1098
rect 772 -1099 773 -1098
rect 786 -1099 787 -1098
rect 1311 -1099 1312 -1098
rect 58 -1101 59 -1100
rect 177 -1101 178 -1100
rect 212 -1101 213 -1100
rect 523 -1101 524 -1100
rect 530 -1101 531 -1100
rect 618 -1101 619 -1100
rect 628 -1101 629 -1100
rect 1136 -1101 1137 -1100
rect 1192 -1101 1193 -1100
rect 1220 -1101 1221 -1100
rect 75 -1103 76 -1102
rect 1101 -1103 1102 -1102
rect 75 -1105 76 -1104
rect 660 -1105 661 -1104
rect 667 -1105 668 -1104
rect 730 -1105 731 -1104
rect 733 -1105 734 -1104
rect 1136 -1105 1137 -1104
rect 79 -1107 80 -1106
rect 544 -1107 545 -1106
rect 558 -1107 559 -1106
rect 765 -1107 766 -1106
rect 863 -1107 864 -1106
rect 1325 -1107 1326 -1106
rect 79 -1109 80 -1108
rect 443 -1109 444 -1108
rect 471 -1109 472 -1108
rect 635 -1109 636 -1108
rect 653 -1109 654 -1108
rect 674 -1109 675 -1108
rect 684 -1109 685 -1108
rect 1206 -1109 1207 -1108
rect 93 -1111 94 -1110
rect 516 -1111 517 -1110
rect 541 -1111 542 -1110
rect 569 -1111 570 -1110
rect 576 -1111 577 -1110
rect 723 -1111 724 -1110
rect 726 -1111 727 -1110
rect 1150 -1111 1151 -1110
rect 1178 -1111 1179 -1110
rect 1206 -1111 1207 -1110
rect 93 -1113 94 -1112
rect 170 -1113 171 -1112
rect 177 -1113 178 -1112
rect 296 -1113 297 -1112
rect 310 -1113 311 -1112
rect 443 -1113 444 -1112
rect 450 -1113 451 -1112
rect 653 -1113 654 -1112
rect 660 -1113 661 -1112
rect 761 -1113 762 -1112
rect 765 -1113 766 -1112
rect 1234 -1113 1235 -1112
rect 72 -1115 73 -1114
rect 170 -1115 171 -1114
rect 205 -1115 206 -1114
rect 471 -1115 472 -1114
rect 478 -1115 479 -1114
rect 485 -1115 486 -1114
rect 492 -1115 493 -1114
rect 989 -1115 990 -1114
rect 1087 -1115 1088 -1114
rect 1101 -1115 1102 -1114
rect 1150 -1115 1151 -1114
rect 1157 -1115 1158 -1114
rect 44 -1117 45 -1116
rect 478 -1117 479 -1116
rect 499 -1117 500 -1116
rect 877 -1117 878 -1116
rect 929 -1117 930 -1116
rect 1304 -1117 1305 -1116
rect 44 -1119 45 -1118
rect 380 -1119 381 -1118
rect 408 -1119 409 -1118
rect 422 -1119 423 -1118
rect 457 -1119 458 -1118
rect 485 -1119 486 -1118
rect 499 -1119 500 -1118
rect 611 -1119 612 -1118
rect 632 -1119 633 -1118
rect 1248 -1119 1249 -1118
rect 1290 -1119 1291 -1118
rect 1304 -1119 1305 -1118
rect 23 -1121 24 -1120
rect 380 -1121 381 -1120
rect 394 -1121 395 -1120
rect 422 -1121 423 -1120
rect 457 -1121 458 -1120
rect 506 -1121 507 -1120
rect 541 -1121 542 -1120
rect 1297 -1121 1298 -1120
rect 23 -1123 24 -1122
rect 366 -1123 367 -1122
rect 464 -1123 465 -1122
rect 611 -1123 612 -1122
rect 695 -1123 696 -1122
rect 754 -1123 755 -1122
rect 828 -1123 829 -1122
rect 877 -1123 878 -1122
rect 954 -1123 955 -1122
rect 1143 -1123 1144 -1122
rect 1227 -1123 1228 -1122
rect 1248 -1123 1249 -1122
rect 1283 -1123 1284 -1122
rect 1297 -1123 1298 -1122
rect 72 -1125 73 -1124
rect 758 -1125 759 -1124
rect 821 -1125 822 -1124
rect 828 -1125 829 -1124
rect 849 -1125 850 -1124
rect 989 -1125 990 -1124
rect 1045 -1125 1046 -1124
rect 1087 -1125 1088 -1124
rect 1171 -1125 1172 -1124
rect 1283 -1125 1284 -1124
rect 96 -1127 97 -1126
rect 639 -1127 640 -1126
rect 681 -1127 682 -1126
rect 695 -1127 696 -1126
rect 712 -1127 713 -1126
rect 1192 -1127 1193 -1126
rect 1199 -1127 1200 -1126
rect 1227 -1127 1228 -1126
rect 100 -1129 101 -1128
rect 849 -1129 850 -1128
rect 866 -1129 867 -1128
rect 1185 -1129 1186 -1128
rect 117 -1131 118 -1130
rect 1185 -1131 1186 -1130
rect 128 -1133 129 -1132
rect 394 -1133 395 -1132
rect 464 -1133 465 -1132
rect 1276 -1133 1277 -1132
rect 128 -1135 129 -1134
rect 632 -1135 633 -1134
rect 716 -1135 717 -1134
rect 723 -1135 724 -1134
rect 730 -1135 731 -1134
rect 1115 -1135 1116 -1134
rect 1262 -1135 1263 -1134
rect 1276 -1135 1277 -1134
rect 149 -1137 150 -1136
rect 646 -1137 647 -1136
rect 702 -1137 703 -1136
rect 716 -1137 717 -1136
rect 744 -1137 745 -1136
rect 835 -1137 836 -1136
rect 870 -1137 871 -1136
rect 1178 -1137 1179 -1136
rect 163 -1139 164 -1138
rect 205 -1139 206 -1138
rect 212 -1139 213 -1138
rect 677 -1139 678 -1138
rect 688 -1139 689 -1138
rect 702 -1139 703 -1138
rect 744 -1139 745 -1138
rect 1122 -1139 1123 -1138
rect 163 -1141 164 -1140
rect 495 -1141 496 -1140
rect 502 -1141 503 -1140
rect 1066 -1141 1067 -1140
rect 1073 -1141 1074 -1140
rect 1115 -1141 1116 -1140
rect 226 -1143 227 -1142
rect 275 -1143 276 -1142
rect 282 -1143 283 -1142
rect 527 -1143 528 -1142
rect 548 -1143 549 -1142
rect 576 -1143 577 -1142
rect 600 -1143 601 -1142
rect 1255 -1143 1256 -1142
rect 152 -1145 153 -1144
rect 275 -1145 276 -1144
rect 289 -1145 290 -1144
rect 467 -1145 468 -1144
rect 495 -1145 496 -1144
rect 870 -1145 871 -1144
rect 905 -1145 906 -1144
rect 954 -1145 955 -1144
rect 968 -1145 969 -1144
rect 1157 -1145 1158 -1144
rect 1255 -1145 1256 -1144
rect 1332 -1145 1333 -1144
rect 184 -1147 185 -1146
rect 282 -1147 283 -1146
rect 296 -1147 297 -1146
rect 352 -1147 353 -1146
rect 373 -1147 374 -1146
rect 639 -1147 640 -1146
rect 649 -1147 650 -1146
rect 688 -1147 689 -1146
rect 747 -1147 748 -1146
rect 940 -1147 941 -1146
rect 1010 -1147 1011 -1146
rect 1045 -1147 1046 -1146
rect 1066 -1147 1067 -1146
rect 1129 -1147 1130 -1146
rect 103 -1149 104 -1148
rect 373 -1149 374 -1148
rect 506 -1149 507 -1148
rect 796 -1149 797 -1148
rect 800 -1149 801 -1148
rect 821 -1149 822 -1148
rect 856 -1149 857 -1148
rect 905 -1149 906 -1148
rect 933 -1149 934 -1148
rect 1073 -1149 1074 -1148
rect 1080 -1149 1081 -1148
rect 1262 -1149 1263 -1148
rect 5 -1151 6 -1150
rect 856 -1151 857 -1150
rect 891 -1151 892 -1150
rect 940 -1151 941 -1150
rect 961 -1151 962 -1150
rect 1010 -1151 1011 -1150
rect 1017 -1151 1018 -1150
rect 1171 -1151 1172 -1150
rect 5 -1153 6 -1152
rect 1290 -1153 1291 -1152
rect 103 -1155 104 -1154
rect 215 -1155 216 -1154
rect 233 -1155 234 -1154
rect 450 -1155 451 -1154
rect 534 -1155 535 -1154
rect 968 -1155 969 -1154
rect 1017 -1155 1018 -1154
rect 1094 -1155 1095 -1154
rect 1108 -1155 1109 -1154
rect 1332 -1155 1333 -1154
rect 135 -1157 136 -1156
rect 233 -1157 234 -1156
rect 240 -1157 241 -1156
rect 247 -1157 248 -1156
rect 254 -1157 255 -1156
rect 376 -1157 377 -1156
rect 534 -1157 535 -1156
rect 646 -1157 647 -1156
rect 709 -1157 710 -1156
rect 891 -1157 892 -1156
rect 912 -1157 913 -1156
rect 961 -1157 962 -1156
rect 1031 -1157 1032 -1156
rect 1199 -1157 1200 -1156
rect 40 -1159 41 -1158
rect 135 -1159 136 -1158
rect 156 -1159 157 -1158
rect 184 -1159 185 -1158
rect 240 -1159 241 -1158
rect 583 -1159 584 -1158
rect 604 -1159 605 -1158
rect 618 -1159 619 -1158
rect 747 -1159 748 -1158
rect 1080 -1159 1081 -1158
rect 156 -1161 157 -1160
rect 436 -1161 437 -1160
rect 481 -1161 482 -1160
rect 583 -1161 584 -1160
rect 607 -1161 608 -1160
rect 1164 -1161 1165 -1160
rect 261 -1163 262 -1162
rect 786 -1163 787 -1162
rect 814 -1163 815 -1162
rect 933 -1163 934 -1162
rect 1052 -1163 1053 -1162
rect 1094 -1163 1095 -1162
rect 191 -1165 192 -1164
rect 261 -1165 262 -1164
rect 303 -1165 304 -1164
rect 835 -1165 836 -1164
rect 884 -1165 885 -1164
rect 1108 -1165 1109 -1164
rect 142 -1167 143 -1166
rect 191 -1167 192 -1166
rect 219 -1167 220 -1166
rect 303 -1167 304 -1166
rect 310 -1167 311 -1166
rect 597 -1167 598 -1166
rect 751 -1167 752 -1166
rect 800 -1167 801 -1166
rect 807 -1167 808 -1166
rect 884 -1167 885 -1166
rect 919 -1167 920 -1166
rect 1031 -1167 1032 -1166
rect 1059 -1167 1060 -1166
rect 1129 -1167 1130 -1166
rect 107 -1169 108 -1168
rect 142 -1169 143 -1168
rect 219 -1169 220 -1168
rect 555 -1169 556 -1168
rect 558 -1169 559 -1168
rect 1122 -1169 1123 -1168
rect 107 -1171 108 -1170
rect 198 -1171 199 -1170
rect 317 -1171 318 -1170
rect 366 -1171 367 -1170
rect 401 -1171 402 -1170
rect 436 -1171 437 -1170
rect 513 -1171 514 -1170
rect 1052 -1171 1053 -1170
rect 180 -1173 181 -1172
rect 513 -1173 514 -1172
rect 530 -1173 531 -1172
rect 1164 -1173 1165 -1172
rect 198 -1175 199 -1174
rect 268 -1175 269 -1174
rect 317 -1175 318 -1174
rect 324 -1175 325 -1174
rect 341 -1175 342 -1174
rect 352 -1175 353 -1174
rect 359 -1175 360 -1174
rect 807 -1175 808 -1174
rect 1024 -1175 1025 -1174
rect 1059 -1175 1060 -1174
rect 254 -1177 255 -1176
rect 401 -1177 402 -1176
rect 555 -1177 556 -1176
rect 1213 -1177 1214 -1176
rect 268 -1179 269 -1178
rect 429 -1179 430 -1178
rect 565 -1179 566 -1178
rect 772 -1179 773 -1178
rect 779 -1179 780 -1178
rect 912 -1179 913 -1178
rect 975 -1179 976 -1178
rect 1024 -1179 1025 -1178
rect 324 -1181 325 -1180
rect 345 -1181 346 -1180
rect 359 -1181 360 -1180
rect 681 -1181 682 -1180
rect 751 -1181 752 -1180
rect 926 -1181 927 -1180
rect 975 -1181 976 -1180
rect 1038 -1181 1039 -1180
rect 331 -1183 332 -1182
rect 779 -1183 780 -1182
rect 793 -1183 794 -1182
rect 814 -1183 815 -1182
rect 1003 -1183 1004 -1182
rect 1038 -1183 1039 -1182
rect 331 -1185 332 -1184
rect 415 -1185 416 -1184
rect 429 -1185 430 -1184
rect 635 -1185 636 -1184
rect 758 -1185 759 -1184
rect 1346 -1185 1347 -1184
rect 51 -1187 52 -1186
rect 1346 -1187 1347 -1186
rect 345 -1189 346 -1188
rect 737 -1189 738 -1188
rect 793 -1189 794 -1188
rect 863 -1189 864 -1188
rect 996 -1189 997 -1188
rect 1003 -1189 1004 -1188
rect 65 -1191 66 -1190
rect 737 -1191 738 -1190
rect 947 -1191 948 -1190
rect 996 -1191 997 -1190
rect 65 -1193 66 -1192
rect 86 -1193 87 -1192
rect 387 -1193 388 -1192
rect 415 -1193 416 -1192
rect 597 -1193 598 -1192
rect 1234 -1193 1235 -1192
rect 86 -1195 87 -1194
rect 114 -1195 115 -1194
rect 387 -1195 388 -1194
rect 492 -1195 493 -1194
rect 625 -1195 626 -1194
rect 919 -1195 920 -1194
rect 51 -1197 52 -1196
rect 625 -1197 626 -1196
rect 898 -1197 899 -1196
rect 947 -1197 948 -1196
rect 114 -1199 115 -1198
rect 590 -1199 591 -1198
rect 551 -1201 552 -1200
rect 898 -1201 899 -1200
rect 590 -1203 591 -1202
rect 709 -1203 710 -1202
rect 2 -1214 3 -1213
rect 303 -1214 304 -1213
rect 366 -1214 367 -1213
rect 558 -1214 559 -1213
rect 607 -1214 608 -1213
rect 968 -1214 969 -1213
rect 1017 -1214 1018 -1213
rect 1020 -1214 1021 -1213
rect 1269 -1214 1270 -1213
rect 1272 -1214 1273 -1213
rect 1360 -1214 1361 -1213
rect 1381 -1214 1382 -1213
rect 1451 -1214 1452 -1213
rect 1458 -1214 1459 -1213
rect 5 -1216 6 -1215
rect 779 -1216 780 -1215
rect 793 -1216 794 -1215
rect 849 -1216 850 -1215
rect 870 -1216 871 -1215
rect 968 -1216 969 -1215
rect 1017 -1216 1018 -1215
rect 1115 -1216 1116 -1215
rect 1269 -1216 1270 -1215
rect 1283 -1216 1284 -1215
rect 30 -1218 31 -1217
rect 551 -1218 552 -1217
rect 614 -1218 615 -1217
rect 618 -1218 619 -1217
rect 628 -1218 629 -1217
rect 695 -1218 696 -1217
rect 698 -1218 699 -1217
rect 1073 -1218 1074 -1217
rect 1283 -1218 1284 -1217
rect 1318 -1218 1319 -1217
rect 30 -1220 31 -1219
rect 562 -1220 563 -1219
rect 632 -1220 633 -1219
rect 1143 -1220 1144 -1219
rect 1272 -1220 1273 -1219
rect 1318 -1220 1319 -1219
rect 37 -1222 38 -1221
rect 212 -1222 213 -1221
rect 289 -1222 290 -1221
rect 562 -1222 563 -1221
rect 646 -1222 647 -1221
rect 1374 -1222 1375 -1221
rect 37 -1224 38 -1223
rect 58 -1224 59 -1223
rect 72 -1224 73 -1223
rect 121 -1224 122 -1223
rect 124 -1224 125 -1223
rect 352 -1224 353 -1223
rect 366 -1224 367 -1223
rect 635 -1224 636 -1223
rect 653 -1224 654 -1223
rect 1388 -1224 1389 -1223
rect 44 -1226 45 -1225
rect 649 -1226 650 -1225
rect 653 -1226 654 -1225
rect 716 -1226 717 -1225
rect 719 -1226 720 -1225
rect 1143 -1226 1144 -1225
rect 44 -1228 45 -1227
rect 93 -1228 94 -1227
rect 100 -1228 101 -1227
rect 117 -1228 118 -1227
rect 121 -1228 122 -1227
rect 555 -1228 556 -1227
rect 600 -1228 601 -1227
rect 646 -1228 647 -1227
rect 684 -1228 685 -1227
rect 1297 -1228 1298 -1227
rect 51 -1230 52 -1229
rect 93 -1230 94 -1229
rect 138 -1230 139 -1229
rect 569 -1230 570 -1229
rect 709 -1230 710 -1229
rect 737 -1230 738 -1229
rect 751 -1230 752 -1229
rect 1374 -1230 1375 -1229
rect 51 -1232 52 -1231
rect 418 -1232 419 -1231
rect 432 -1232 433 -1231
rect 534 -1232 535 -1231
rect 544 -1232 545 -1231
rect 1360 -1232 1361 -1231
rect 58 -1234 59 -1233
rect 478 -1234 479 -1233
rect 492 -1234 493 -1233
rect 884 -1234 885 -1233
rect 915 -1234 916 -1233
rect 1080 -1234 1081 -1233
rect 1150 -1234 1151 -1233
rect 1297 -1234 1298 -1233
rect 75 -1236 76 -1235
rect 422 -1236 423 -1235
rect 436 -1236 437 -1235
rect 464 -1236 465 -1235
rect 520 -1236 521 -1235
rect 709 -1236 710 -1235
rect 712 -1236 713 -1235
rect 1094 -1236 1095 -1235
rect 1150 -1236 1151 -1235
rect 1157 -1236 1158 -1235
rect 89 -1238 90 -1237
rect 226 -1238 227 -1237
rect 289 -1238 290 -1237
rect 373 -1238 374 -1237
rect 394 -1238 395 -1237
rect 530 -1238 531 -1237
rect 534 -1238 535 -1237
rect 705 -1238 706 -1237
rect 754 -1238 755 -1237
rect 1339 -1238 1340 -1237
rect 149 -1240 150 -1239
rect 597 -1240 598 -1239
rect 604 -1240 605 -1239
rect 884 -1240 885 -1239
rect 1010 -1240 1011 -1239
rect 1073 -1240 1074 -1239
rect 1080 -1240 1081 -1239
rect 1108 -1240 1109 -1239
rect 1157 -1240 1158 -1239
rect 1171 -1240 1172 -1239
rect 149 -1242 150 -1241
rect 345 -1242 346 -1241
rect 352 -1242 353 -1241
rect 387 -1242 388 -1241
rect 436 -1242 437 -1241
rect 541 -1242 542 -1241
rect 548 -1242 549 -1241
rect 996 -1242 997 -1241
rect 1010 -1242 1011 -1241
rect 1038 -1242 1039 -1241
rect 1094 -1242 1095 -1241
rect 1178 -1242 1179 -1241
rect 173 -1244 174 -1243
rect 1199 -1244 1200 -1243
rect 177 -1246 178 -1245
rect 254 -1246 255 -1245
rect 282 -1246 283 -1245
rect 387 -1246 388 -1245
rect 446 -1246 447 -1245
rect 1199 -1246 1200 -1245
rect 191 -1248 192 -1247
rect 303 -1248 304 -1247
rect 310 -1248 311 -1247
rect 618 -1248 619 -1247
rect 660 -1248 661 -1247
rect 751 -1248 752 -1247
rect 765 -1248 766 -1247
rect 1024 -1248 1025 -1247
rect 1038 -1248 1039 -1247
rect 1045 -1248 1046 -1247
rect 1129 -1248 1130 -1247
rect 1171 -1248 1172 -1247
rect 1178 -1248 1179 -1247
rect 1192 -1248 1193 -1247
rect 170 -1250 171 -1249
rect 191 -1250 192 -1249
rect 198 -1250 199 -1249
rect 681 -1250 682 -1249
rect 695 -1250 696 -1249
rect 737 -1250 738 -1249
rect 758 -1250 759 -1249
rect 1045 -1250 1046 -1249
rect 1164 -1250 1165 -1249
rect 1339 -1250 1340 -1249
rect 198 -1252 199 -1251
rect 296 -1252 297 -1251
rect 310 -1252 311 -1251
rect 495 -1252 496 -1251
rect 520 -1252 521 -1251
rect 572 -1252 573 -1251
rect 604 -1252 605 -1251
rect 611 -1252 612 -1251
rect 660 -1252 661 -1251
rect 702 -1252 703 -1251
rect 758 -1252 759 -1251
rect 786 -1252 787 -1251
rect 796 -1252 797 -1251
rect 1206 -1252 1207 -1251
rect 205 -1254 206 -1253
rect 394 -1254 395 -1253
rect 450 -1254 451 -1253
rect 492 -1254 493 -1253
rect 527 -1254 528 -1253
rect 1234 -1254 1235 -1253
rect 135 -1256 136 -1255
rect 205 -1256 206 -1255
rect 212 -1256 213 -1255
rect 317 -1256 318 -1255
rect 331 -1256 332 -1255
rect 422 -1256 423 -1255
rect 464 -1256 465 -1255
rect 471 -1256 472 -1255
rect 527 -1256 528 -1255
rect 544 -1256 545 -1255
rect 548 -1256 549 -1255
rect 733 -1256 734 -1255
rect 765 -1256 766 -1255
rect 807 -1256 808 -1255
rect 842 -1256 843 -1255
rect 1262 -1256 1263 -1255
rect 135 -1258 136 -1257
rect 1220 -1258 1221 -1257
rect 1234 -1258 1235 -1257
rect 1248 -1258 1249 -1257
rect 219 -1260 220 -1259
rect 597 -1260 598 -1259
rect 621 -1260 622 -1259
rect 1248 -1260 1249 -1259
rect 156 -1262 157 -1261
rect 219 -1262 220 -1261
rect 226 -1262 227 -1261
rect 467 -1262 468 -1261
rect 555 -1262 556 -1261
rect 576 -1262 577 -1261
rect 681 -1262 682 -1261
rect 1367 -1262 1368 -1261
rect 103 -1264 104 -1263
rect 156 -1264 157 -1263
rect 233 -1264 234 -1263
rect 282 -1264 283 -1263
rect 296 -1264 297 -1263
rect 408 -1264 409 -1263
rect 457 -1264 458 -1263
rect 471 -1264 472 -1263
rect 569 -1264 570 -1263
rect 1332 -1264 1333 -1263
rect 1353 -1264 1354 -1263
rect 1367 -1264 1368 -1263
rect 16 -1266 17 -1265
rect 457 -1266 458 -1265
rect 576 -1266 577 -1265
rect 590 -1266 591 -1265
rect 779 -1266 780 -1265
rect 800 -1266 801 -1265
rect 807 -1266 808 -1265
rect 821 -1266 822 -1265
rect 828 -1266 829 -1265
rect 842 -1266 843 -1265
rect 845 -1266 846 -1265
rect 954 -1266 955 -1265
rect 989 -1266 990 -1265
rect 996 -1266 997 -1265
rect 1003 -1266 1004 -1265
rect 1129 -1266 1130 -1265
rect 1164 -1266 1165 -1265
rect 1185 -1266 1186 -1265
rect 1332 -1266 1333 -1265
rect 1346 -1266 1347 -1265
rect 16 -1268 17 -1267
rect 639 -1268 640 -1267
rect 786 -1268 787 -1267
rect 835 -1268 836 -1267
rect 849 -1268 850 -1267
rect 891 -1268 892 -1267
rect 961 -1268 962 -1267
rect 989 -1268 990 -1267
rect 1003 -1268 1004 -1267
rect 1031 -1268 1032 -1267
rect 1066 -1268 1067 -1267
rect 1206 -1268 1207 -1267
rect 1255 -1268 1256 -1267
rect 1346 -1268 1347 -1267
rect 61 -1270 62 -1269
rect 1353 -1270 1354 -1269
rect 170 -1272 171 -1271
rect 1066 -1272 1067 -1271
rect 1087 -1272 1088 -1271
rect 1220 -1272 1221 -1271
rect 1255 -1272 1256 -1271
rect 1276 -1272 1277 -1271
rect 233 -1274 234 -1273
rect 506 -1274 507 -1273
rect 625 -1274 626 -1273
rect 835 -1274 836 -1273
rect 866 -1274 867 -1273
rect 1262 -1274 1263 -1273
rect 1276 -1274 1277 -1273
rect 1290 -1274 1291 -1273
rect 240 -1276 241 -1275
rect 450 -1276 451 -1275
rect 485 -1276 486 -1275
rect 506 -1276 507 -1275
rect 583 -1276 584 -1275
rect 625 -1276 626 -1275
rect 639 -1276 640 -1275
rect 674 -1276 675 -1275
rect 800 -1276 801 -1275
rect 898 -1276 899 -1275
rect 933 -1276 934 -1275
rect 961 -1276 962 -1275
rect 975 -1276 976 -1275
rect 1031 -1276 1032 -1275
rect 1087 -1276 1088 -1275
rect 1101 -1276 1102 -1275
rect 1122 -1276 1123 -1275
rect 1185 -1276 1186 -1275
rect 1290 -1276 1291 -1275
rect 1325 -1276 1326 -1275
rect 68 -1278 69 -1277
rect 1122 -1278 1123 -1277
rect 1311 -1278 1312 -1277
rect 1325 -1278 1326 -1277
rect 114 -1280 115 -1279
rect 1101 -1280 1102 -1279
rect 65 -1282 66 -1281
rect 114 -1282 115 -1281
rect 240 -1282 241 -1281
rect 632 -1282 633 -1281
rect 744 -1282 745 -1281
rect 933 -1282 934 -1281
rect 1024 -1282 1025 -1281
rect 1052 -1282 1053 -1281
rect 247 -1284 248 -1283
rect 317 -1284 318 -1283
rect 324 -1284 325 -1283
rect 485 -1284 486 -1283
rect 499 -1284 500 -1283
rect 674 -1284 675 -1283
rect 730 -1284 731 -1283
rect 1052 -1284 1053 -1283
rect 79 -1286 80 -1285
rect 499 -1286 500 -1285
rect 583 -1286 584 -1285
rect 768 -1286 769 -1285
rect 821 -1286 822 -1285
rect 856 -1286 857 -1285
rect 870 -1286 871 -1285
rect 947 -1286 948 -1285
rect 79 -1288 80 -1287
rect 254 -1288 255 -1287
rect 331 -1288 332 -1287
rect 429 -1288 430 -1287
rect 443 -1288 444 -1287
rect 590 -1288 591 -1287
rect 730 -1288 731 -1287
rect 1059 -1288 1060 -1287
rect 107 -1290 108 -1289
rect 443 -1290 444 -1289
rect 513 -1290 514 -1289
rect 947 -1290 948 -1289
rect 1059 -1290 1060 -1289
rect 1227 -1290 1228 -1289
rect 86 -1292 87 -1291
rect 107 -1292 108 -1291
rect 184 -1292 185 -1291
rect 324 -1292 325 -1291
rect 338 -1292 339 -1291
rect 478 -1292 479 -1291
rect 513 -1292 514 -1291
rect 688 -1292 689 -1291
rect 744 -1292 745 -1291
rect 817 -1292 818 -1291
rect 828 -1292 829 -1291
rect 926 -1292 927 -1291
rect 1213 -1292 1214 -1291
rect 1227 -1292 1228 -1291
rect 86 -1294 87 -1293
rect 1108 -1294 1109 -1293
rect 1213 -1294 1214 -1293
rect 1241 -1294 1242 -1293
rect 184 -1296 185 -1295
rect 733 -1296 734 -1295
rect 747 -1296 748 -1295
rect 975 -1296 976 -1295
rect 247 -1298 248 -1297
rect 611 -1298 612 -1297
rect 688 -1298 689 -1297
rect 723 -1298 724 -1297
rect 856 -1298 857 -1297
rect 863 -1298 864 -1297
rect 891 -1298 892 -1297
rect 905 -1298 906 -1297
rect 338 -1300 339 -1299
rect 401 -1300 402 -1299
rect 523 -1300 524 -1299
rect 1241 -1300 1242 -1299
rect 9 -1302 10 -1301
rect 401 -1302 402 -1301
rect 702 -1302 703 -1301
rect 926 -1302 927 -1301
rect 9 -1304 10 -1303
rect 772 -1304 773 -1303
rect 863 -1304 864 -1303
rect 1311 -1304 1312 -1303
rect 345 -1306 346 -1305
rect 415 -1306 416 -1305
rect 772 -1306 773 -1305
rect 814 -1306 815 -1305
rect 898 -1306 899 -1305
rect 954 -1306 955 -1305
rect 268 -1308 269 -1307
rect 415 -1308 416 -1307
rect 814 -1308 815 -1307
rect 1136 -1308 1137 -1307
rect 268 -1310 269 -1309
rect 359 -1310 360 -1309
rect 369 -1310 370 -1309
rect 1192 -1310 1193 -1309
rect 359 -1312 360 -1311
rect 541 -1312 542 -1311
rect 905 -1312 906 -1311
rect 919 -1312 920 -1311
rect 376 -1314 377 -1313
rect 723 -1314 724 -1313
rect 912 -1314 913 -1313
rect 919 -1314 920 -1313
rect 380 -1316 381 -1315
rect 408 -1316 409 -1315
rect 761 -1316 762 -1315
rect 912 -1316 913 -1315
rect 23 -1318 24 -1317
rect 380 -1318 381 -1317
rect 404 -1318 405 -1317
rect 1136 -1318 1137 -1317
rect 23 -1320 24 -1319
rect 128 -1320 129 -1319
rect 128 -1322 129 -1321
rect 275 -1322 276 -1321
rect 275 -1324 276 -1323
rect 390 -1324 391 -1323
rect 33 -1335 34 -1334
rect 107 -1335 108 -1334
rect 121 -1335 122 -1334
rect 1353 -1335 1354 -1334
rect 1423 -1335 1424 -1334
rect 1451 -1335 1452 -1334
rect 1458 -1335 1459 -1334
rect 1465 -1335 1466 -1334
rect 44 -1337 45 -1336
rect 373 -1337 374 -1336
rect 387 -1337 388 -1336
rect 1066 -1337 1067 -1336
rect 1122 -1337 1123 -1336
rect 1402 -1337 1403 -1336
rect 44 -1339 45 -1338
rect 751 -1339 752 -1338
rect 814 -1339 815 -1338
rect 1227 -1339 1228 -1338
rect 1255 -1339 1256 -1338
rect 1353 -1339 1354 -1338
rect 1360 -1339 1361 -1338
rect 1458 -1339 1459 -1338
rect 65 -1341 66 -1340
rect 555 -1341 556 -1340
rect 583 -1341 584 -1340
rect 618 -1341 619 -1340
rect 635 -1341 636 -1340
rect 877 -1341 878 -1340
rect 887 -1341 888 -1340
rect 1374 -1341 1375 -1340
rect 65 -1343 66 -1342
rect 124 -1343 125 -1342
rect 135 -1343 136 -1342
rect 1430 -1343 1431 -1342
rect 61 -1345 62 -1344
rect 135 -1345 136 -1344
rect 163 -1345 164 -1344
rect 782 -1345 783 -1344
rect 793 -1345 794 -1344
rect 877 -1345 878 -1344
rect 898 -1345 899 -1344
rect 1073 -1345 1074 -1344
rect 1129 -1345 1130 -1344
rect 1409 -1345 1410 -1344
rect 68 -1347 69 -1346
rect 446 -1347 447 -1346
rect 464 -1347 465 -1346
rect 569 -1347 570 -1346
rect 614 -1347 615 -1346
rect 1080 -1347 1081 -1346
rect 1150 -1347 1151 -1346
rect 1227 -1347 1228 -1346
rect 1262 -1347 1263 -1346
rect 1360 -1347 1361 -1346
rect 30 -1349 31 -1348
rect 569 -1349 570 -1348
rect 646 -1349 647 -1348
rect 817 -1349 818 -1348
rect 821 -1349 822 -1348
rect 898 -1349 899 -1348
rect 912 -1349 913 -1348
rect 1367 -1349 1368 -1348
rect 79 -1351 80 -1350
rect 324 -1351 325 -1350
rect 380 -1351 381 -1350
rect 446 -1351 447 -1350
rect 509 -1351 510 -1350
rect 1304 -1351 1305 -1350
rect 1332 -1351 1333 -1350
rect 1437 -1351 1438 -1350
rect 82 -1353 83 -1352
rect 1220 -1353 1221 -1352
rect 1234 -1353 1235 -1352
rect 1332 -1353 1333 -1352
rect 1339 -1353 1340 -1352
rect 1374 -1353 1375 -1352
rect 82 -1355 83 -1354
rect 747 -1355 748 -1354
rect 821 -1355 822 -1354
rect 1248 -1355 1249 -1354
rect 1269 -1355 1270 -1354
rect 1367 -1355 1368 -1354
rect 86 -1357 87 -1356
rect 100 -1357 101 -1356
rect 107 -1357 108 -1356
rect 366 -1357 367 -1356
rect 380 -1357 381 -1356
rect 684 -1357 685 -1356
rect 695 -1357 696 -1356
rect 723 -1357 724 -1356
rect 852 -1357 853 -1356
rect 1052 -1357 1053 -1356
rect 1094 -1357 1095 -1356
rect 1248 -1357 1249 -1356
rect 1297 -1357 1298 -1356
rect 1416 -1357 1417 -1356
rect 86 -1359 87 -1358
rect 219 -1359 220 -1358
rect 254 -1359 255 -1358
rect 366 -1359 367 -1358
rect 376 -1359 377 -1358
rect 1052 -1359 1053 -1358
rect 1059 -1359 1060 -1358
rect 1297 -1359 1298 -1358
rect 1318 -1359 1319 -1358
rect 1339 -1359 1340 -1358
rect 1346 -1359 1347 -1358
rect 1444 -1359 1445 -1358
rect 100 -1361 101 -1360
rect 296 -1361 297 -1360
rect 317 -1361 318 -1360
rect 373 -1361 374 -1360
rect 415 -1361 416 -1360
rect 1311 -1361 1312 -1360
rect 23 -1363 24 -1362
rect 296 -1363 297 -1362
rect 324 -1363 325 -1362
rect 331 -1363 332 -1362
rect 418 -1363 419 -1362
rect 856 -1363 857 -1362
rect 866 -1363 867 -1362
rect 968 -1363 969 -1362
rect 982 -1363 983 -1362
rect 1066 -1363 1067 -1362
rect 1157 -1363 1158 -1362
rect 1220 -1363 1221 -1362
rect 1241 -1363 1242 -1362
rect 1346 -1363 1347 -1362
rect 23 -1365 24 -1364
rect 247 -1365 248 -1364
rect 429 -1365 430 -1364
rect 859 -1365 860 -1364
rect 968 -1365 969 -1364
rect 975 -1365 976 -1364
rect 996 -1365 997 -1364
rect 1073 -1365 1074 -1364
rect 1164 -1365 1165 -1364
rect 1234 -1365 1235 -1364
rect 37 -1367 38 -1366
rect 317 -1367 318 -1366
rect 429 -1367 430 -1366
rect 572 -1367 573 -1366
rect 583 -1367 584 -1366
rect 646 -1367 647 -1366
rect 649 -1367 650 -1366
rect 1038 -1367 1039 -1366
rect 1045 -1367 1046 -1366
rect 1048 -1367 1049 -1366
rect 1164 -1367 1165 -1366
rect 1171 -1367 1172 -1366
rect 1178 -1367 1179 -1366
rect 1262 -1367 1263 -1366
rect 37 -1369 38 -1368
rect 534 -1369 535 -1368
rect 541 -1369 542 -1368
rect 947 -1369 948 -1368
rect 954 -1369 955 -1368
rect 1038 -1369 1039 -1368
rect 1045 -1369 1046 -1368
rect 1388 -1369 1389 -1368
rect 93 -1371 94 -1370
rect 331 -1371 332 -1370
rect 436 -1371 437 -1370
rect 695 -1371 696 -1370
rect 698 -1371 699 -1370
rect 954 -1371 955 -1370
rect 1017 -1371 1018 -1370
rect 1129 -1371 1130 -1370
rect 1192 -1371 1193 -1370
rect 1255 -1371 1256 -1370
rect 1276 -1371 1277 -1370
rect 1388 -1371 1389 -1370
rect 93 -1373 94 -1372
rect 460 -1373 461 -1372
rect 534 -1373 535 -1372
rect 555 -1373 556 -1372
rect 632 -1373 633 -1372
rect 1311 -1373 1312 -1372
rect 121 -1375 122 -1374
rect 149 -1375 150 -1374
rect 152 -1375 153 -1374
rect 415 -1375 416 -1374
rect 436 -1375 437 -1374
rect 457 -1375 458 -1374
rect 541 -1375 542 -1374
rect 786 -1375 787 -1374
rect 793 -1375 794 -1374
rect 982 -1375 983 -1374
rect 1024 -1375 1025 -1374
rect 1094 -1375 1095 -1374
rect 1101 -1375 1102 -1374
rect 1171 -1375 1172 -1374
rect 1192 -1375 1193 -1374
rect 1283 -1375 1284 -1374
rect 128 -1377 129 -1376
rect 254 -1377 255 -1376
rect 443 -1377 444 -1376
rect 1157 -1377 1158 -1376
rect 1199 -1377 1200 -1376
rect 1283 -1377 1284 -1376
rect 128 -1379 129 -1378
rect 310 -1379 311 -1378
rect 457 -1379 458 -1378
rect 1318 -1379 1319 -1378
rect 131 -1381 132 -1380
rect 1269 -1381 1270 -1380
rect 149 -1383 150 -1382
rect 590 -1383 591 -1382
rect 632 -1383 633 -1382
rect 856 -1383 857 -1382
rect 870 -1383 871 -1382
rect 1024 -1383 1025 -1382
rect 1031 -1383 1032 -1382
rect 1122 -1383 1123 -1382
rect 1199 -1383 1200 -1382
rect 1290 -1383 1291 -1382
rect 163 -1385 164 -1384
rect 411 -1385 412 -1384
rect 527 -1385 528 -1384
rect 870 -1385 871 -1384
rect 884 -1385 885 -1384
rect 947 -1385 948 -1384
rect 1010 -1385 1011 -1384
rect 1101 -1385 1102 -1384
rect 1206 -1385 1207 -1384
rect 1276 -1385 1277 -1384
rect 170 -1387 171 -1386
rect 912 -1387 913 -1386
rect 933 -1387 934 -1386
rect 996 -1387 997 -1386
rect 1143 -1387 1144 -1386
rect 1206 -1387 1207 -1386
rect 170 -1389 171 -1388
rect 681 -1389 682 -1388
rect 702 -1389 703 -1388
rect 989 -1389 990 -1388
rect 1048 -1389 1049 -1388
rect 1143 -1389 1144 -1388
rect 198 -1391 199 -1390
rect 397 -1391 398 -1390
rect 513 -1391 514 -1390
rect 681 -1391 682 -1390
rect 705 -1391 706 -1390
rect 961 -1391 962 -1390
rect 184 -1393 185 -1392
rect 198 -1393 199 -1392
rect 212 -1393 213 -1392
rect 369 -1393 370 -1392
rect 394 -1393 395 -1392
rect 527 -1393 528 -1392
rect 544 -1393 545 -1392
rect 660 -1393 661 -1392
rect 667 -1393 668 -1392
rect 751 -1393 752 -1392
rect 758 -1393 759 -1392
rect 786 -1393 787 -1392
rect 814 -1393 815 -1392
rect 1290 -1393 1291 -1392
rect 184 -1395 185 -1394
rect 240 -1395 241 -1394
rect 247 -1395 248 -1394
rect 565 -1395 566 -1394
rect 590 -1395 591 -1394
rect 653 -1395 654 -1394
rect 667 -1395 668 -1394
rect 800 -1395 801 -1394
rect 828 -1395 829 -1394
rect 1010 -1395 1011 -1394
rect 191 -1397 192 -1396
rect 212 -1397 213 -1396
rect 219 -1397 220 -1396
rect 320 -1397 321 -1396
rect 401 -1397 402 -1396
rect 513 -1397 514 -1396
rect 551 -1397 552 -1396
rect 1080 -1397 1081 -1396
rect 2 -1399 3 -1398
rect 191 -1399 192 -1398
rect 240 -1399 241 -1398
rect 485 -1399 486 -1398
rect 492 -1399 493 -1398
rect 653 -1399 654 -1398
rect 716 -1399 717 -1398
rect 779 -1399 780 -1398
rect 831 -1399 832 -1398
rect 1178 -1399 1179 -1398
rect 2 -1401 3 -1400
rect 51 -1401 52 -1400
rect 275 -1401 276 -1400
rect 800 -1401 801 -1400
rect 842 -1401 843 -1400
rect 933 -1401 934 -1400
rect 940 -1401 941 -1400
rect 1017 -1401 1018 -1400
rect 51 -1403 52 -1402
rect 261 -1403 262 -1402
rect 275 -1403 276 -1402
rect 548 -1403 549 -1402
rect 625 -1403 626 -1402
rect 702 -1403 703 -1402
rect 716 -1403 717 -1402
rect 744 -1403 745 -1402
rect 758 -1403 759 -1402
rect 772 -1403 773 -1402
rect 779 -1403 780 -1402
rect 1150 -1403 1151 -1402
rect 79 -1405 80 -1404
rect 261 -1405 262 -1404
rect 303 -1405 304 -1404
rect 394 -1405 395 -1404
rect 450 -1405 451 -1404
rect 485 -1405 486 -1404
rect 492 -1405 493 -1404
rect 520 -1405 521 -1404
rect 548 -1405 549 -1404
rect 1325 -1405 1326 -1404
rect 89 -1407 90 -1406
rect 940 -1407 941 -1406
rect 1213 -1407 1214 -1406
rect 1325 -1407 1326 -1406
rect 138 -1409 139 -1408
rect 842 -1409 843 -1408
rect 866 -1409 867 -1408
rect 1031 -1409 1032 -1408
rect 1185 -1409 1186 -1408
rect 1213 -1409 1214 -1408
rect 282 -1411 283 -1410
rect 450 -1411 451 -1410
rect 464 -1411 465 -1410
rect 744 -1411 745 -1410
rect 891 -1411 892 -1410
rect 961 -1411 962 -1410
rect 1115 -1411 1116 -1410
rect 1185 -1411 1186 -1410
rect 282 -1413 283 -1412
rect 289 -1413 290 -1412
rect 303 -1413 304 -1412
rect 352 -1413 353 -1412
rect 520 -1413 521 -1412
rect 1395 -1413 1396 -1412
rect 289 -1415 290 -1414
rect 765 -1415 766 -1414
rect 796 -1415 797 -1414
rect 1115 -1415 1116 -1414
rect 310 -1417 311 -1416
rect 726 -1417 727 -1416
rect 730 -1417 731 -1416
rect 1059 -1417 1060 -1416
rect 352 -1419 353 -1418
rect 359 -1419 360 -1418
rect 562 -1419 563 -1418
rect 765 -1419 766 -1418
rect 905 -1419 906 -1418
rect 975 -1419 976 -1418
rect 338 -1421 339 -1420
rect 562 -1421 563 -1420
rect 597 -1421 598 -1420
rect 625 -1421 626 -1420
rect 639 -1421 640 -1420
rect 660 -1421 661 -1420
rect 688 -1421 689 -1420
rect 730 -1421 731 -1420
rect 737 -1421 738 -1420
rect 772 -1421 773 -1420
rect 905 -1421 906 -1420
rect 1108 -1421 1109 -1420
rect 166 -1423 167 -1422
rect 597 -1423 598 -1422
rect 604 -1423 605 -1422
rect 688 -1423 689 -1422
rect 709 -1423 710 -1422
rect 737 -1423 738 -1422
rect 926 -1423 927 -1422
rect 989 -1423 990 -1422
rect 1087 -1423 1088 -1422
rect 1108 -1423 1109 -1422
rect 268 -1425 269 -1424
rect 338 -1425 339 -1424
rect 359 -1425 360 -1424
rect 499 -1425 500 -1424
rect 576 -1425 577 -1424
rect 604 -1425 605 -1424
rect 642 -1425 643 -1424
rect 891 -1425 892 -1424
rect 915 -1425 916 -1424
rect 926 -1425 927 -1424
rect 1003 -1425 1004 -1424
rect 1087 -1425 1088 -1424
rect 58 -1427 59 -1426
rect 1003 -1427 1004 -1426
rect 58 -1429 59 -1428
rect 72 -1429 73 -1428
rect 114 -1429 115 -1428
rect 268 -1429 269 -1428
rect 387 -1429 388 -1428
rect 639 -1429 640 -1428
rect 674 -1429 675 -1428
rect 709 -1429 710 -1428
rect 719 -1429 720 -1428
rect 1381 -1429 1382 -1428
rect 72 -1431 73 -1430
rect 226 -1431 227 -1430
rect 499 -1431 500 -1430
rect 506 -1431 507 -1430
rect 611 -1431 612 -1430
rect 674 -1431 675 -1430
rect 723 -1431 724 -1430
rect 1304 -1431 1305 -1430
rect 16 -1433 17 -1432
rect 611 -1433 612 -1432
rect 919 -1433 920 -1432
rect 1381 -1433 1382 -1432
rect 16 -1435 17 -1434
rect 408 -1435 409 -1434
rect 506 -1435 507 -1434
rect 1241 -1435 1242 -1434
rect 114 -1437 115 -1436
rect 345 -1437 346 -1436
rect 408 -1437 409 -1436
rect 807 -1437 808 -1436
rect 835 -1437 836 -1436
rect 919 -1437 920 -1436
rect 173 -1439 174 -1438
rect 576 -1439 577 -1438
rect 807 -1439 808 -1438
rect 849 -1439 850 -1438
rect 226 -1441 227 -1440
rect 233 -1441 234 -1440
rect 345 -1441 346 -1440
rect 422 -1441 423 -1440
rect 828 -1441 829 -1440
rect 835 -1441 836 -1440
rect 156 -1443 157 -1442
rect 233 -1443 234 -1442
rect 401 -1443 402 -1442
rect 849 -1443 850 -1442
rect 156 -1445 157 -1444
rect 177 -1445 178 -1444
rect 422 -1445 423 -1444
rect 471 -1445 472 -1444
rect 142 -1447 143 -1446
rect 177 -1447 178 -1446
rect 390 -1447 391 -1446
rect 471 -1447 472 -1446
rect 142 -1449 143 -1448
rect 824 -1449 825 -1448
rect 9 -1460 10 -1459
rect 33 -1460 34 -1459
rect 44 -1460 45 -1459
rect 457 -1460 458 -1459
rect 460 -1460 461 -1459
rect 940 -1460 941 -1459
rect 1454 -1460 1455 -1459
rect 1465 -1460 1466 -1459
rect 12 -1462 13 -1461
rect 268 -1462 269 -1461
rect 282 -1462 283 -1461
rect 520 -1462 521 -1461
rect 523 -1462 524 -1461
rect 709 -1462 710 -1461
rect 723 -1462 724 -1461
rect 835 -1462 836 -1461
rect 852 -1462 853 -1461
rect 1276 -1462 1277 -1461
rect 19 -1464 20 -1463
rect 1402 -1464 1403 -1463
rect 44 -1466 45 -1465
rect 485 -1466 486 -1465
rect 520 -1466 521 -1465
rect 688 -1466 689 -1465
rect 702 -1466 703 -1465
rect 782 -1466 783 -1465
rect 793 -1466 794 -1465
rect 1269 -1466 1270 -1465
rect 51 -1468 52 -1467
rect 509 -1468 510 -1467
rect 534 -1468 535 -1467
rect 590 -1468 591 -1467
rect 621 -1468 622 -1467
rect 1297 -1468 1298 -1467
rect 51 -1470 52 -1469
rect 730 -1470 731 -1469
rect 744 -1470 745 -1469
rect 1227 -1470 1228 -1469
rect 1269 -1470 1270 -1469
rect 1367 -1470 1368 -1469
rect 65 -1472 66 -1471
rect 537 -1472 538 -1471
rect 558 -1472 559 -1471
rect 1010 -1472 1011 -1471
rect 1297 -1472 1298 -1471
rect 1395 -1472 1396 -1471
rect 65 -1474 66 -1473
rect 870 -1474 871 -1473
rect 884 -1474 885 -1473
rect 1038 -1474 1039 -1473
rect 93 -1476 94 -1475
rect 488 -1476 489 -1475
rect 534 -1476 535 -1475
rect 667 -1476 668 -1475
rect 688 -1476 689 -1475
rect 695 -1476 696 -1475
rect 705 -1476 706 -1475
rect 1052 -1476 1053 -1475
rect 37 -1478 38 -1477
rect 93 -1478 94 -1477
rect 100 -1478 101 -1477
rect 548 -1478 549 -1477
rect 562 -1478 563 -1477
rect 1234 -1478 1235 -1477
rect 37 -1480 38 -1479
rect 898 -1480 899 -1479
rect 940 -1480 941 -1479
rect 996 -1480 997 -1479
rect 1010 -1480 1011 -1479
rect 1073 -1480 1074 -1479
rect 1234 -1480 1235 -1479
rect 1318 -1480 1319 -1479
rect 103 -1482 104 -1481
rect 450 -1482 451 -1481
rect 548 -1482 549 -1481
rect 604 -1482 605 -1481
rect 639 -1482 640 -1481
rect 1381 -1482 1382 -1481
rect 107 -1484 108 -1483
rect 117 -1484 118 -1483
rect 121 -1484 122 -1483
rect 152 -1484 153 -1483
rect 180 -1484 181 -1483
rect 730 -1484 731 -1483
rect 779 -1484 780 -1483
rect 1332 -1484 1333 -1483
rect 100 -1486 101 -1485
rect 107 -1486 108 -1485
rect 121 -1486 122 -1485
rect 415 -1486 416 -1485
rect 443 -1486 444 -1485
rect 765 -1486 766 -1485
rect 793 -1486 794 -1485
rect 842 -1486 843 -1485
rect 859 -1486 860 -1485
rect 1325 -1486 1326 -1485
rect 1332 -1486 1333 -1485
rect 1430 -1486 1431 -1485
rect 128 -1488 129 -1487
rect 1171 -1488 1172 -1487
rect 1318 -1488 1319 -1487
rect 1416 -1488 1417 -1487
rect 128 -1490 129 -1489
rect 422 -1490 423 -1489
rect 446 -1490 447 -1489
rect 1227 -1490 1228 -1489
rect 1325 -1490 1326 -1489
rect 1423 -1490 1424 -1489
rect 131 -1492 132 -1491
rect 432 -1492 433 -1491
rect 450 -1492 451 -1491
rect 653 -1492 654 -1491
rect 663 -1492 664 -1491
rect 1451 -1492 1452 -1491
rect 138 -1494 139 -1493
rect 800 -1494 801 -1493
rect 814 -1494 815 -1493
rect 1157 -1494 1158 -1493
rect 1171 -1494 1172 -1493
rect 1255 -1494 1256 -1493
rect 149 -1496 150 -1495
rect 849 -1496 850 -1495
rect 863 -1496 864 -1495
rect 1409 -1496 1410 -1495
rect 149 -1498 150 -1497
rect 170 -1498 171 -1497
rect 240 -1498 241 -1497
rect 537 -1498 538 -1497
rect 562 -1498 563 -1497
rect 618 -1498 619 -1497
rect 639 -1498 640 -1497
rect 660 -1498 661 -1497
rect 667 -1498 668 -1497
rect 737 -1498 738 -1497
rect 758 -1498 759 -1497
rect 779 -1498 780 -1497
rect 796 -1498 797 -1497
rect 1045 -1498 1046 -1497
rect 1052 -1498 1053 -1497
rect 1101 -1498 1102 -1497
rect 1157 -1498 1158 -1497
rect 1213 -1498 1214 -1497
rect 72 -1500 73 -1499
rect 170 -1500 171 -1499
rect 191 -1500 192 -1499
rect 240 -1500 241 -1499
rect 261 -1500 262 -1499
rect 604 -1500 605 -1499
rect 653 -1500 654 -1499
rect 681 -1500 682 -1499
rect 702 -1500 703 -1499
rect 1213 -1500 1214 -1499
rect 58 -1502 59 -1501
rect 72 -1502 73 -1501
rect 86 -1502 87 -1501
rect 191 -1502 192 -1501
rect 254 -1502 255 -1501
rect 261 -1502 262 -1501
rect 268 -1502 269 -1501
rect 408 -1502 409 -1501
rect 415 -1502 416 -1501
rect 611 -1502 612 -1501
rect 709 -1502 710 -1501
rect 747 -1502 748 -1501
rect 765 -1502 766 -1501
rect 786 -1502 787 -1501
rect 800 -1502 801 -1501
rect 1346 -1502 1347 -1501
rect 23 -1504 24 -1503
rect 786 -1504 787 -1503
rect 814 -1504 815 -1503
rect 877 -1504 878 -1503
rect 898 -1504 899 -1503
rect 1094 -1504 1095 -1503
rect 1192 -1504 1193 -1503
rect 1255 -1504 1256 -1503
rect 1346 -1504 1347 -1503
rect 1444 -1504 1445 -1503
rect 23 -1506 24 -1505
rect 54 -1506 55 -1505
rect 58 -1506 59 -1505
rect 310 -1506 311 -1505
rect 331 -1506 332 -1505
rect 695 -1506 696 -1505
rect 716 -1506 717 -1505
rect 744 -1506 745 -1505
rect 817 -1506 818 -1505
rect 1087 -1506 1088 -1505
rect 1094 -1506 1095 -1505
rect 1311 -1506 1312 -1505
rect 16 -1508 17 -1507
rect 310 -1508 311 -1507
rect 338 -1508 339 -1507
rect 422 -1508 423 -1507
rect 478 -1508 479 -1507
rect 618 -1508 619 -1507
rect 716 -1508 717 -1507
rect 751 -1508 752 -1507
rect 821 -1508 822 -1507
rect 894 -1508 895 -1507
rect 982 -1508 983 -1507
rect 1276 -1508 1277 -1507
rect 16 -1510 17 -1509
rect 681 -1510 682 -1509
rect 723 -1510 724 -1509
rect 772 -1510 773 -1509
rect 824 -1510 825 -1509
rect 1374 -1510 1375 -1509
rect 219 -1512 220 -1511
rect 331 -1512 332 -1511
rect 338 -1512 339 -1511
rect 499 -1512 500 -1511
rect 565 -1512 566 -1511
rect 751 -1512 752 -1511
rect 828 -1512 829 -1511
rect 1185 -1512 1186 -1511
rect 1192 -1512 1193 -1511
rect 1290 -1512 1291 -1511
rect 2 -1514 3 -1513
rect 219 -1514 220 -1513
rect 247 -1514 248 -1513
rect 254 -1514 255 -1513
rect 282 -1514 283 -1513
rect 345 -1514 346 -1513
rect 380 -1514 381 -1513
rect 443 -1514 444 -1513
rect 478 -1514 479 -1513
rect 492 -1514 493 -1513
rect 572 -1514 573 -1513
rect 866 -1514 867 -1513
rect 870 -1514 871 -1513
rect 1017 -1514 1018 -1513
rect 1038 -1514 1039 -1513
rect 1080 -1514 1081 -1513
rect 1185 -1514 1186 -1513
rect 1283 -1514 1284 -1513
rect 2 -1516 3 -1515
rect 275 -1516 276 -1515
rect 289 -1516 290 -1515
rect 772 -1516 773 -1515
rect 831 -1516 832 -1515
rect 1122 -1516 1123 -1515
rect 1199 -1516 1200 -1515
rect 1311 -1516 1312 -1515
rect 9 -1518 10 -1517
rect 275 -1518 276 -1517
rect 289 -1518 290 -1517
rect 457 -1518 458 -1517
rect 485 -1518 486 -1517
rect 758 -1518 759 -1517
rect 831 -1518 832 -1517
rect 1360 -1518 1361 -1517
rect 114 -1520 115 -1519
rect 499 -1520 500 -1519
rect 583 -1520 584 -1519
rect 642 -1520 643 -1519
rect 835 -1520 836 -1519
rect 891 -1520 892 -1519
rect 905 -1520 906 -1519
rect 1122 -1520 1123 -1519
rect 1129 -1520 1130 -1519
rect 1199 -1520 1200 -1519
rect 1283 -1520 1284 -1519
rect 1388 -1520 1389 -1519
rect 40 -1522 41 -1521
rect 583 -1522 584 -1521
rect 590 -1522 591 -1521
rect 674 -1522 675 -1521
rect 842 -1522 843 -1521
rect 912 -1522 913 -1521
rect 954 -1522 955 -1521
rect 982 -1522 983 -1521
rect 996 -1522 997 -1521
rect 1150 -1522 1151 -1521
rect 89 -1524 90 -1523
rect 912 -1524 913 -1523
rect 1059 -1524 1060 -1523
rect 1101 -1524 1102 -1523
rect 1129 -1524 1130 -1523
rect 1178 -1524 1179 -1523
rect 30 -1526 31 -1525
rect 1178 -1526 1179 -1525
rect 30 -1528 31 -1527
rect 359 -1528 360 -1527
rect 380 -1528 381 -1527
rect 597 -1528 598 -1527
rect 611 -1528 612 -1527
rect 646 -1528 647 -1527
rect 649 -1528 650 -1527
rect 674 -1528 675 -1527
rect 807 -1528 808 -1527
rect 954 -1528 955 -1527
rect 1073 -1528 1074 -1527
rect 1304 -1528 1305 -1527
rect 114 -1530 115 -1529
rect 737 -1530 738 -1529
rect 849 -1530 850 -1529
rect 919 -1530 920 -1529
rect 1080 -1530 1081 -1529
rect 1220 -1530 1221 -1529
rect 1304 -1530 1305 -1529
rect 1339 -1530 1340 -1529
rect 142 -1532 143 -1531
rect 1017 -1532 1018 -1531
rect 1115 -1532 1116 -1531
rect 1220 -1532 1221 -1531
rect 1339 -1532 1340 -1531
rect 1437 -1532 1438 -1531
rect 142 -1534 143 -1533
rect 233 -1534 234 -1533
rect 317 -1534 318 -1533
rect 1059 -1534 1060 -1533
rect 1108 -1534 1109 -1533
rect 1115 -1534 1116 -1533
rect 1150 -1534 1151 -1533
rect 1241 -1534 1242 -1533
rect 198 -1536 199 -1535
rect 247 -1536 248 -1535
rect 324 -1536 325 -1535
rect 905 -1536 906 -1535
rect 919 -1536 920 -1535
rect 961 -1536 962 -1535
rect 82 -1538 83 -1537
rect 324 -1538 325 -1537
rect 345 -1538 346 -1537
rect 366 -1538 367 -1537
rect 397 -1538 398 -1537
rect 1136 -1538 1137 -1537
rect 198 -1540 199 -1539
rect 212 -1540 213 -1539
rect 233 -1540 234 -1539
rect 303 -1540 304 -1539
rect 352 -1540 353 -1539
rect 359 -1540 360 -1539
rect 366 -1540 367 -1539
rect 576 -1540 577 -1539
rect 625 -1540 626 -1539
rect 646 -1540 647 -1539
rect 859 -1540 860 -1539
rect 1136 -1540 1137 -1539
rect 177 -1542 178 -1541
rect 212 -1542 213 -1541
rect 296 -1542 297 -1541
rect 303 -1542 304 -1541
rect 352 -1542 353 -1541
rect 373 -1542 374 -1541
rect 404 -1542 405 -1541
rect 632 -1542 633 -1541
rect 863 -1542 864 -1541
rect 933 -1542 934 -1541
rect 961 -1542 962 -1541
rect 1024 -1542 1025 -1541
rect 135 -1544 136 -1543
rect 296 -1544 297 -1543
rect 373 -1544 374 -1543
rect 387 -1544 388 -1543
rect 408 -1544 409 -1543
rect 492 -1544 493 -1543
rect 513 -1544 514 -1543
rect 576 -1544 577 -1543
rect 625 -1544 626 -1543
rect 926 -1544 927 -1543
rect 933 -1544 934 -1543
rect 989 -1544 990 -1543
rect 1024 -1544 1025 -1543
rect 1206 -1544 1207 -1543
rect 79 -1546 80 -1545
rect 513 -1546 514 -1545
rect 541 -1546 542 -1545
rect 807 -1546 808 -1545
rect 877 -1546 878 -1545
rect 947 -1546 948 -1545
rect 968 -1546 969 -1545
rect 989 -1546 990 -1545
rect 1143 -1546 1144 -1545
rect 1206 -1546 1207 -1545
rect 79 -1548 80 -1547
rect 86 -1548 87 -1547
rect 135 -1548 136 -1547
rect 1241 -1548 1242 -1547
rect 205 -1550 206 -1549
rect 317 -1550 318 -1549
rect 387 -1550 388 -1549
rect 464 -1550 465 -1549
rect 541 -1550 542 -1549
rect 569 -1550 570 -1549
rect 891 -1550 892 -1549
rect 1262 -1550 1263 -1549
rect 205 -1552 206 -1551
rect 551 -1552 552 -1551
rect 555 -1552 556 -1551
rect 597 -1552 598 -1551
rect 926 -1552 927 -1551
rect 975 -1552 976 -1551
rect 1143 -1552 1144 -1551
rect 1164 -1552 1165 -1551
rect 1262 -1552 1263 -1551
rect 1353 -1552 1354 -1551
rect 394 -1554 395 -1553
rect 464 -1554 465 -1553
rect 555 -1554 556 -1553
rect 1045 -1554 1046 -1553
rect 1353 -1554 1354 -1553
rect 1458 -1554 1459 -1553
rect 394 -1556 395 -1555
rect 436 -1556 437 -1555
rect 569 -1556 570 -1555
rect 1290 -1556 1291 -1555
rect 401 -1558 402 -1557
rect 436 -1558 437 -1557
rect 856 -1558 857 -1557
rect 975 -1558 976 -1557
rect 163 -1560 164 -1559
rect 401 -1560 402 -1559
rect 429 -1560 430 -1559
rect 632 -1560 633 -1559
rect 856 -1560 857 -1559
rect 1108 -1560 1109 -1559
rect 163 -1562 164 -1561
rect 1003 -1562 1004 -1561
rect 429 -1564 430 -1563
rect 1087 -1564 1088 -1563
rect 887 -1566 888 -1565
rect 1164 -1566 1165 -1565
rect 947 -1568 948 -1567
rect 1048 -1568 1049 -1567
rect 968 -1570 969 -1569
rect 1031 -1570 1032 -1569
rect 145 -1572 146 -1571
rect 1031 -1572 1032 -1571
rect 1003 -1574 1004 -1573
rect 1066 -1574 1067 -1573
rect 1066 -1576 1067 -1575
rect 1248 -1576 1249 -1575
rect 506 -1578 507 -1577
rect 1248 -1578 1249 -1577
rect 471 -1580 472 -1579
rect 506 -1580 507 -1579
rect 184 -1582 185 -1581
rect 471 -1582 472 -1581
rect 156 -1584 157 -1583
rect 184 -1584 185 -1583
rect 156 -1586 157 -1585
rect 803 -1586 804 -1585
rect 2 -1597 3 -1596
rect 558 -1597 559 -1596
rect 569 -1597 570 -1596
rect 849 -1597 850 -1596
rect 856 -1597 857 -1596
rect 1066 -1597 1067 -1596
rect 1094 -1597 1095 -1596
rect 1097 -1597 1098 -1596
rect 1255 -1597 1256 -1596
rect 1258 -1597 1259 -1596
rect 2 -1599 3 -1598
rect 401 -1599 402 -1598
rect 415 -1599 416 -1598
rect 569 -1599 570 -1598
rect 572 -1599 573 -1598
rect 576 -1599 577 -1598
rect 632 -1599 633 -1598
rect 663 -1599 664 -1598
rect 705 -1599 706 -1598
rect 954 -1599 955 -1598
rect 1045 -1599 1046 -1598
rect 1346 -1599 1347 -1598
rect 9 -1601 10 -1600
rect 940 -1601 941 -1600
rect 954 -1601 955 -1600
rect 1129 -1601 1130 -1600
rect 1255 -1601 1256 -1600
rect 1283 -1601 1284 -1600
rect 12 -1603 13 -1602
rect 163 -1603 164 -1602
rect 177 -1603 178 -1602
rect 212 -1603 213 -1602
rect 320 -1603 321 -1602
rect 905 -1603 906 -1602
rect 940 -1603 941 -1602
rect 1318 -1603 1319 -1602
rect 51 -1605 52 -1604
rect 583 -1605 584 -1604
rect 632 -1605 633 -1604
rect 716 -1605 717 -1604
rect 754 -1605 755 -1604
rect 1136 -1605 1137 -1604
rect 1304 -1605 1305 -1604
rect 1318 -1605 1319 -1604
rect 58 -1607 59 -1606
rect 415 -1607 416 -1606
rect 485 -1607 486 -1606
rect 639 -1607 640 -1606
rect 660 -1607 661 -1606
rect 688 -1607 689 -1606
rect 716 -1607 717 -1606
rect 737 -1607 738 -1606
rect 775 -1607 776 -1606
rect 863 -1607 864 -1606
rect 884 -1607 885 -1606
rect 905 -1607 906 -1606
rect 975 -1607 976 -1606
rect 1136 -1607 1137 -1606
rect 1304 -1607 1305 -1606
rect 1332 -1607 1333 -1606
rect 58 -1609 59 -1608
rect 513 -1609 514 -1608
rect 534 -1609 535 -1608
rect 982 -1609 983 -1608
rect 1045 -1609 1046 -1608
rect 1108 -1609 1109 -1608
rect 1129 -1609 1130 -1608
rect 1171 -1609 1172 -1608
rect 65 -1611 66 -1610
rect 551 -1611 552 -1610
rect 639 -1611 640 -1610
rect 674 -1611 675 -1610
rect 688 -1611 689 -1610
rect 765 -1611 766 -1610
rect 800 -1611 801 -1610
rect 1199 -1611 1200 -1610
rect 65 -1613 66 -1612
rect 702 -1613 703 -1612
rect 765 -1613 766 -1612
rect 779 -1613 780 -1612
rect 803 -1613 804 -1612
rect 1108 -1613 1109 -1612
rect 1199 -1613 1200 -1612
rect 1234 -1613 1235 -1612
rect 79 -1615 80 -1614
rect 800 -1615 801 -1614
rect 849 -1615 850 -1614
rect 870 -1615 871 -1614
rect 884 -1615 885 -1614
rect 898 -1615 899 -1614
rect 975 -1615 976 -1614
rect 1052 -1615 1053 -1614
rect 1094 -1615 1095 -1614
rect 1150 -1615 1151 -1614
rect 1234 -1615 1235 -1614
rect 1325 -1615 1326 -1614
rect 86 -1617 87 -1616
rect 488 -1617 489 -1616
rect 495 -1617 496 -1616
rect 548 -1617 549 -1616
rect 625 -1617 626 -1616
rect 674 -1617 675 -1616
rect 779 -1617 780 -1616
rect 814 -1617 815 -1616
rect 856 -1617 857 -1616
rect 1328 -1617 1329 -1616
rect 86 -1619 87 -1618
rect 107 -1619 108 -1618
rect 110 -1619 111 -1618
rect 576 -1619 577 -1618
rect 621 -1619 622 -1618
rect 625 -1619 626 -1618
rect 660 -1619 661 -1618
rect 1003 -1619 1004 -1618
rect 1052 -1619 1053 -1618
rect 1122 -1619 1123 -1618
rect 1220 -1619 1221 -1618
rect 1325 -1619 1326 -1618
rect 40 -1621 41 -1620
rect 1003 -1621 1004 -1620
rect 1220 -1621 1221 -1620
rect 1276 -1621 1277 -1620
rect 89 -1623 90 -1622
rect 709 -1623 710 -1622
rect 814 -1623 815 -1622
rect 842 -1623 843 -1622
rect 859 -1623 860 -1622
rect 1059 -1623 1060 -1622
rect 1258 -1623 1259 -1622
rect 1283 -1623 1284 -1622
rect 100 -1625 101 -1624
rect 1185 -1625 1186 -1624
rect 1276 -1625 1277 -1624
rect 1353 -1625 1354 -1624
rect 23 -1627 24 -1626
rect 100 -1627 101 -1626
rect 107 -1627 108 -1626
rect 583 -1627 584 -1626
rect 709 -1627 710 -1626
rect 744 -1627 745 -1626
rect 842 -1627 843 -1626
rect 877 -1627 878 -1626
rect 891 -1627 892 -1626
rect 1262 -1627 1263 -1626
rect 117 -1629 118 -1628
rect 184 -1629 185 -1628
rect 194 -1629 195 -1628
rect 380 -1629 381 -1628
rect 499 -1629 500 -1628
rect 534 -1629 535 -1628
rect 537 -1629 538 -1628
rect 702 -1629 703 -1628
rect 737 -1629 738 -1628
rect 744 -1629 745 -1628
rect 863 -1629 864 -1628
rect 919 -1629 920 -1628
rect 947 -1629 948 -1628
rect 1185 -1629 1186 -1628
rect 1262 -1629 1263 -1628
rect 1290 -1629 1291 -1628
rect 138 -1631 139 -1630
rect 471 -1631 472 -1630
rect 485 -1631 486 -1630
rect 499 -1631 500 -1630
rect 506 -1631 507 -1630
rect 523 -1631 524 -1630
rect 730 -1631 731 -1630
rect 947 -1631 948 -1630
rect 982 -1631 983 -1630
rect 1038 -1631 1039 -1630
rect 1290 -1631 1291 -1630
rect 1311 -1631 1312 -1630
rect 142 -1633 143 -1632
rect 1101 -1633 1102 -1632
rect 1311 -1633 1312 -1632
rect 1339 -1633 1340 -1632
rect 47 -1635 48 -1634
rect 142 -1635 143 -1634
rect 145 -1635 146 -1634
rect 254 -1635 255 -1634
rect 338 -1635 339 -1634
rect 457 -1635 458 -1634
rect 471 -1635 472 -1634
rect 611 -1635 612 -1634
rect 730 -1635 731 -1634
rect 747 -1635 748 -1634
rect 870 -1635 871 -1634
rect 968 -1635 969 -1634
rect 996 -1635 997 -1634
rect 1038 -1635 1039 -1634
rect 1080 -1635 1081 -1634
rect 1101 -1635 1102 -1634
rect 93 -1637 94 -1636
rect 338 -1637 339 -1636
rect 352 -1637 353 -1636
rect 457 -1637 458 -1636
rect 506 -1637 507 -1636
rect 961 -1637 962 -1636
rect 968 -1637 969 -1636
rect 989 -1637 990 -1636
rect 996 -1637 997 -1636
rect 1164 -1637 1165 -1636
rect 93 -1639 94 -1638
rect 1206 -1639 1207 -1638
rect 103 -1641 104 -1640
rect 989 -1641 990 -1640
rect 1164 -1641 1165 -1640
rect 1213 -1641 1214 -1640
rect 135 -1643 136 -1642
rect 1213 -1643 1214 -1642
rect 135 -1645 136 -1644
rect 198 -1645 199 -1644
rect 212 -1645 213 -1644
rect 247 -1645 248 -1644
rect 254 -1645 255 -1644
rect 429 -1645 430 -1644
rect 443 -1645 444 -1644
rect 611 -1645 612 -1644
rect 877 -1645 878 -1644
rect 933 -1645 934 -1644
rect 961 -1645 962 -1644
rect 1031 -1645 1032 -1644
rect 1206 -1645 1207 -1644
rect 1227 -1645 1228 -1644
rect 121 -1647 122 -1646
rect 443 -1647 444 -1646
rect 460 -1647 461 -1646
rect 933 -1647 934 -1646
rect 1031 -1647 1032 -1646
rect 1087 -1647 1088 -1646
rect 1157 -1647 1158 -1646
rect 1227 -1647 1228 -1646
rect 114 -1649 115 -1648
rect 1087 -1649 1088 -1648
rect 96 -1651 97 -1650
rect 114 -1651 115 -1650
rect 121 -1651 122 -1650
rect 240 -1651 241 -1650
rect 247 -1651 248 -1650
rect 275 -1651 276 -1650
rect 352 -1651 353 -1650
rect 492 -1651 493 -1650
rect 513 -1651 514 -1650
rect 758 -1651 759 -1650
rect 894 -1651 895 -1650
rect 1178 -1651 1179 -1650
rect 152 -1653 153 -1652
rect 282 -1653 283 -1652
rect 366 -1653 367 -1652
rect 432 -1653 433 -1652
rect 492 -1653 493 -1652
rect 527 -1653 528 -1652
rect 758 -1653 759 -1652
rect 772 -1653 773 -1652
rect 1066 -1653 1067 -1652
rect 1178 -1653 1179 -1652
rect 159 -1655 160 -1654
rect 1059 -1655 1060 -1654
rect 1073 -1655 1074 -1654
rect 1157 -1655 1158 -1654
rect 163 -1657 164 -1656
rect 831 -1657 832 -1656
rect 1024 -1657 1025 -1656
rect 1073 -1657 1074 -1656
rect 177 -1659 178 -1658
rect 751 -1659 752 -1658
rect 772 -1659 773 -1658
rect 1115 -1659 1116 -1658
rect 180 -1661 181 -1660
rect 359 -1661 360 -1660
rect 366 -1661 367 -1660
rect 562 -1661 563 -1660
rect 751 -1661 752 -1660
rect 919 -1661 920 -1660
rect 1024 -1661 1025 -1660
rect 1241 -1661 1242 -1660
rect 44 -1663 45 -1662
rect 359 -1663 360 -1662
rect 373 -1663 374 -1662
rect 429 -1663 430 -1662
rect 523 -1663 524 -1662
rect 1171 -1663 1172 -1662
rect 1241 -1663 1242 -1662
rect 1269 -1663 1270 -1662
rect 44 -1665 45 -1664
rect 54 -1665 55 -1664
rect 184 -1665 185 -1664
rect 205 -1665 206 -1664
rect 240 -1665 241 -1664
rect 296 -1665 297 -1664
rect 376 -1665 377 -1664
rect 1017 -1665 1018 -1664
rect 1115 -1665 1116 -1664
rect 1143 -1665 1144 -1664
rect 54 -1667 55 -1666
rect 79 -1667 80 -1666
rect 198 -1667 199 -1666
rect 331 -1667 332 -1666
rect 380 -1667 381 -1666
rect 422 -1667 423 -1666
rect 450 -1667 451 -1666
rect 1017 -1667 1018 -1666
rect 1143 -1667 1144 -1666
rect 1192 -1667 1193 -1666
rect 51 -1669 52 -1668
rect 1192 -1669 1193 -1668
rect 205 -1671 206 -1670
rect 404 -1671 405 -1670
rect 422 -1671 423 -1670
rect 436 -1671 437 -1670
rect 450 -1671 451 -1670
rect 695 -1671 696 -1670
rect 828 -1671 829 -1670
rect 1269 -1671 1270 -1670
rect 226 -1673 227 -1672
rect 296 -1673 297 -1672
rect 324 -1673 325 -1672
rect 828 -1673 829 -1672
rect 226 -1675 227 -1674
rect 310 -1675 311 -1674
rect 324 -1675 325 -1674
rect 387 -1675 388 -1674
rect 394 -1675 395 -1674
rect 436 -1675 437 -1674
rect 527 -1675 528 -1674
rect 541 -1675 542 -1674
rect 562 -1675 563 -1674
rect 670 -1675 671 -1674
rect 695 -1675 696 -1674
rect 901 -1675 902 -1674
rect 128 -1677 129 -1676
rect 387 -1677 388 -1676
rect 394 -1677 395 -1676
rect 597 -1677 598 -1676
rect 72 -1679 73 -1678
rect 128 -1679 129 -1678
rect 275 -1679 276 -1678
rect 289 -1679 290 -1678
rect 303 -1679 304 -1678
rect 310 -1679 311 -1678
rect 331 -1679 332 -1678
rect 520 -1679 521 -1678
rect 541 -1679 542 -1678
rect 786 -1679 787 -1678
rect 72 -1681 73 -1680
rect 261 -1681 262 -1680
rect 282 -1681 283 -1680
rect 618 -1681 619 -1680
rect 786 -1681 787 -1680
rect 821 -1681 822 -1680
rect 156 -1683 157 -1682
rect 261 -1683 262 -1682
rect 404 -1683 405 -1682
rect 460 -1683 461 -1682
rect 555 -1683 556 -1682
rect 618 -1683 619 -1682
rect 821 -1683 822 -1682
rect 898 -1683 899 -1682
rect 30 -1685 31 -1684
rect 555 -1685 556 -1684
rect 590 -1685 591 -1684
rect 597 -1685 598 -1684
rect 16 -1687 17 -1686
rect 30 -1687 31 -1686
rect 170 -1687 171 -1686
rect 303 -1687 304 -1686
rect 408 -1687 409 -1686
rect 590 -1687 591 -1686
rect 170 -1689 171 -1688
rect 268 -1689 269 -1688
rect 408 -1689 409 -1688
rect 604 -1689 605 -1688
rect 149 -1691 150 -1690
rect 268 -1691 269 -1690
rect 604 -1691 605 -1690
rect 646 -1691 647 -1690
rect 149 -1693 150 -1692
rect 912 -1693 913 -1692
rect 219 -1695 220 -1694
rect 289 -1695 290 -1694
rect 520 -1695 521 -1694
rect 912 -1695 913 -1694
rect 191 -1697 192 -1696
rect 219 -1697 220 -1696
rect 646 -1697 647 -1696
rect 681 -1697 682 -1696
rect 191 -1699 192 -1698
rect 653 -1699 654 -1698
rect 681 -1699 682 -1698
rect 723 -1699 724 -1698
rect 653 -1701 654 -1700
rect 667 -1701 668 -1700
rect 723 -1701 724 -1700
rect 793 -1701 794 -1700
rect 667 -1703 668 -1702
rect 1297 -1703 1298 -1702
rect 793 -1705 794 -1704
rect 807 -1705 808 -1704
rect 1248 -1705 1249 -1704
rect 1297 -1705 1298 -1704
rect 37 -1707 38 -1706
rect 1248 -1707 1249 -1706
rect 37 -1709 38 -1708
rect 317 -1709 318 -1708
rect 807 -1709 808 -1708
rect 835 -1709 836 -1708
rect 317 -1711 318 -1710
rect 1080 -1711 1081 -1710
rect 835 -1713 836 -1712
rect 926 -1713 927 -1712
rect 926 -1715 927 -1714
rect 1010 -1715 1011 -1714
rect 373 -1717 374 -1716
rect 1010 -1717 1011 -1716
rect 9 -1728 10 -1727
rect 110 -1728 111 -1727
rect 117 -1728 118 -1727
rect 646 -1728 647 -1727
rect 667 -1728 668 -1727
rect 933 -1728 934 -1727
rect 940 -1728 941 -1727
rect 968 -1728 969 -1727
rect 1069 -1728 1070 -1727
rect 1241 -1728 1242 -1727
rect 1318 -1728 1319 -1727
rect 1328 -1728 1329 -1727
rect 16 -1730 17 -1729
rect 30 -1730 31 -1729
rect 33 -1730 34 -1729
rect 68 -1730 69 -1729
rect 72 -1730 73 -1729
rect 373 -1730 374 -1729
rect 390 -1730 391 -1729
rect 856 -1730 857 -1729
rect 898 -1730 899 -1729
rect 1101 -1730 1102 -1729
rect 1122 -1730 1123 -1729
rect 1276 -1730 1277 -1729
rect 16 -1732 17 -1731
rect 149 -1732 150 -1731
rect 152 -1732 153 -1731
rect 1101 -1732 1102 -1731
rect 1122 -1732 1123 -1731
rect 1171 -1732 1172 -1731
rect 1227 -1732 1228 -1731
rect 1286 -1732 1287 -1731
rect 9 -1734 10 -1733
rect 152 -1734 153 -1733
rect 205 -1734 206 -1733
rect 355 -1734 356 -1733
rect 359 -1734 360 -1733
rect 646 -1734 647 -1733
rect 667 -1734 668 -1733
rect 702 -1734 703 -1733
rect 712 -1734 713 -1733
rect 765 -1734 766 -1733
rect 814 -1734 815 -1733
rect 891 -1734 892 -1733
rect 898 -1734 899 -1733
rect 975 -1734 976 -1733
rect 1171 -1734 1172 -1733
rect 1213 -1734 1214 -1733
rect 1241 -1734 1242 -1733
rect 1290 -1734 1291 -1733
rect 19 -1736 20 -1735
rect 793 -1736 794 -1735
rect 835 -1736 836 -1735
rect 856 -1736 857 -1735
rect 901 -1736 902 -1735
rect 1276 -1736 1277 -1735
rect 23 -1738 24 -1737
rect 611 -1738 612 -1737
rect 702 -1738 703 -1737
rect 723 -1738 724 -1737
rect 744 -1738 745 -1737
rect 849 -1738 850 -1737
rect 933 -1738 934 -1737
rect 947 -1738 948 -1737
rect 968 -1738 969 -1737
rect 1045 -1738 1046 -1737
rect 1213 -1738 1214 -1737
rect 1255 -1738 1256 -1737
rect 26 -1740 27 -1739
rect 100 -1740 101 -1739
rect 107 -1740 108 -1739
rect 1017 -1740 1018 -1739
rect 1255 -1740 1256 -1739
rect 1304 -1740 1305 -1739
rect 26 -1742 27 -1741
rect 982 -1742 983 -1741
rect 1010 -1742 1011 -1741
rect 1045 -1742 1046 -1741
rect 30 -1744 31 -1743
rect 268 -1744 269 -1743
rect 324 -1744 325 -1743
rect 376 -1744 377 -1743
rect 404 -1744 405 -1743
rect 534 -1744 535 -1743
rect 548 -1744 549 -1743
rect 793 -1744 794 -1743
rect 835 -1744 836 -1743
rect 870 -1744 871 -1743
rect 940 -1744 941 -1743
rect 996 -1744 997 -1743
rect 1017 -1744 1018 -1743
rect 1073 -1744 1074 -1743
rect 37 -1746 38 -1745
rect 159 -1746 160 -1745
rect 205 -1746 206 -1745
rect 310 -1746 311 -1745
rect 359 -1746 360 -1745
rect 387 -1746 388 -1745
rect 457 -1746 458 -1745
rect 1297 -1746 1298 -1745
rect 44 -1748 45 -1747
rect 240 -1748 241 -1747
rect 268 -1748 269 -1747
rect 415 -1748 416 -1747
rect 457 -1748 458 -1747
rect 551 -1748 552 -1747
rect 555 -1748 556 -1747
rect 632 -1748 633 -1747
rect 719 -1748 720 -1747
rect 884 -1748 885 -1747
rect 975 -1748 976 -1747
rect 1031 -1748 1032 -1747
rect 1073 -1748 1074 -1747
rect 1115 -1748 1116 -1747
rect 44 -1750 45 -1749
rect 1059 -1750 1060 -1749
rect 1115 -1750 1116 -1749
rect 1164 -1750 1165 -1749
rect 47 -1752 48 -1751
rect 996 -1752 997 -1751
rect 1031 -1752 1032 -1751
rect 1094 -1752 1095 -1751
rect 1164 -1752 1165 -1751
rect 1192 -1752 1193 -1751
rect 54 -1754 55 -1753
rect 1248 -1754 1249 -1753
rect 72 -1756 73 -1755
rect 93 -1756 94 -1755
rect 100 -1756 101 -1755
rect 467 -1756 468 -1755
rect 485 -1756 486 -1755
rect 1227 -1756 1228 -1755
rect 1234 -1756 1235 -1755
rect 1248 -1756 1249 -1755
rect 51 -1758 52 -1757
rect 93 -1758 94 -1757
rect 107 -1758 108 -1757
rect 289 -1758 290 -1757
rect 369 -1758 370 -1757
rect 744 -1758 745 -1757
rect 747 -1758 748 -1757
rect 821 -1758 822 -1757
rect 849 -1758 850 -1757
rect 912 -1758 913 -1757
rect 1059 -1758 1060 -1757
rect 1108 -1758 1109 -1757
rect 1192 -1758 1193 -1757
rect 1220 -1758 1221 -1757
rect 1234 -1758 1235 -1757
rect 1283 -1758 1284 -1757
rect 51 -1760 52 -1759
rect 842 -1760 843 -1759
rect 912 -1760 913 -1759
rect 989 -1760 990 -1759
rect 1108 -1760 1109 -1759
rect 1150 -1760 1151 -1759
rect 1220 -1760 1221 -1759
rect 1269 -1760 1270 -1759
rect 58 -1762 59 -1761
rect 842 -1762 843 -1761
rect 989 -1762 990 -1761
rect 1052 -1762 1053 -1761
rect 1269 -1762 1270 -1761
rect 1311 -1762 1312 -1761
rect 58 -1764 59 -1763
rect 184 -1764 185 -1763
rect 226 -1764 227 -1763
rect 523 -1764 524 -1763
rect 534 -1764 535 -1763
rect 807 -1764 808 -1763
rect 821 -1764 822 -1763
rect 926 -1764 927 -1763
rect 1052 -1764 1053 -1763
rect 1087 -1764 1088 -1763
rect 2 -1766 3 -1765
rect 226 -1766 227 -1765
rect 233 -1766 234 -1765
rect 240 -1766 241 -1765
rect 275 -1766 276 -1765
rect 324 -1766 325 -1765
rect 373 -1766 374 -1765
rect 614 -1766 615 -1765
rect 625 -1766 626 -1765
rect 807 -1766 808 -1765
rect 926 -1766 927 -1765
rect 1003 -1766 1004 -1765
rect 1087 -1766 1088 -1765
rect 1143 -1766 1144 -1765
rect 2 -1768 3 -1767
rect 54 -1768 55 -1767
rect 79 -1768 80 -1767
rect 586 -1768 587 -1767
rect 604 -1768 605 -1767
rect 947 -1768 948 -1767
rect 1143 -1768 1144 -1767
rect 1185 -1768 1186 -1767
rect 79 -1770 80 -1769
rect 86 -1770 87 -1769
rect 121 -1770 122 -1769
rect 317 -1770 318 -1769
rect 401 -1770 402 -1769
rect 1185 -1770 1186 -1769
rect 86 -1772 87 -1771
rect 299 -1772 300 -1771
rect 317 -1772 318 -1771
rect 331 -1772 332 -1771
rect 401 -1772 402 -1771
rect 422 -1772 423 -1771
rect 488 -1772 489 -1771
rect 894 -1772 895 -1771
rect 114 -1774 115 -1773
rect 121 -1774 122 -1773
rect 128 -1774 129 -1773
rect 289 -1774 290 -1773
rect 331 -1774 332 -1773
rect 345 -1774 346 -1773
rect 415 -1774 416 -1773
rect 436 -1774 437 -1773
rect 506 -1774 507 -1773
rect 642 -1774 643 -1773
rect 660 -1774 661 -1773
rect 884 -1774 885 -1773
rect 128 -1776 129 -1775
rect 261 -1776 262 -1775
rect 345 -1776 346 -1775
rect 380 -1776 381 -1775
rect 436 -1776 437 -1775
rect 471 -1776 472 -1775
rect 506 -1776 507 -1775
rect 541 -1776 542 -1775
rect 555 -1776 556 -1775
rect 772 -1776 773 -1775
rect 138 -1778 139 -1777
rect 303 -1778 304 -1777
rect 464 -1778 465 -1777
rect 471 -1778 472 -1777
rect 513 -1778 514 -1777
rect 548 -1778 549 -1777
rect 576 -1778 577 -1777
rect 1094 -1778 1095 -1777
rect 142 -1780 143 -1779
rect 1283 -1780 1284 -1779
rect 142 -1782 143 -1781
rect 481 -1782 482 -1781
rect 513 -1782 514 -1781
rect 527 -1782 528 -1781
rect 541 -1782 542 -1781
rect 562 -1782 563 -1781
rect 576 -1782 577 -1781
rect 597 -1782 598 -1781
rect 611 -1782 612 -1781
rect 688 -1782 689 -1781
rect 723 -1782 724 -1781
rect 775 -1782 776 -1781
rect 149 -1784 150 -1783
rect 590 -1784 591 -1783
rect 597 -1784 598 -1783
rect 639 -1784 640 -1783
rect 660 -1784 661 -1783
rect 681 -1784 682 -1783
rect 730 -1784 731 -1783
rect 1010 -1784 1011 -1783
rect 156 -1786 157 -1785
rect 590 -1786 591 -1785
rect 625 -1786 626 -1785
rect 863 -1786 864 -1785
rect 156 -1788 157 -1787
rect 170 -1788 171 -1787
rect 177 -1788 178 -1787
rect 681 -1788 682 -1787
rect 730 -1788 731 -1787
rect 919 -1788 920 -1787
rect 96 -1790 97 -1789
rect 919 -1790 920 -1789
rect 163 -1792 164 -1791
rect 380 -1792 381 -1791
rect 408 -1792 409 -1791
rect 527 -1792 528 -1791
rect 562 -1792 563 -1791
rect 618 -1792 619 -1791
rect 628 -1792 629 -1791
rect 1003 -1792 1004 -1791
rect 170 -1794 171 -1793
rect 282 -1794 283 -1793
rect 394 -1794 395 -1793
rect 408 -1794 409 -1793
rect 464 -1794 465 -1793
rect 982 -1794 983 -1793
rect 177 -1796 178 -1795
rect 296 -1796 297 -1795
rect 394 -1796 395 -1795
rect 460 -1796 461 -1795
rect 520 -1796 521 -1795
rect 1206 -1796 1207 -1795
rect 184 -1798 185 -1797
rect 219 -1798 220 -1797
rect 233 -1798 234 -1797
rect 450 -1798 451 -1797
rect 520 -1798 521 -1797
rect 943 -1798 944 -1797
rect 65 -1800 66 -1799
rect 219 -1800 220 -1799
rect 247 -1800 248 -1799
rect 275 -1800 276 -1799
rect 282 -1800 283 -1799
rect 499 -1800 500 -1799
rect 569 -1800 570 -1799
rect 688 -1800 689 -1799
rect 733 -1800 734 -1799
rect 772 -1800 773 -1799
rect 863 -1800 864 -1799
rect 954 -1800 955 -1799
rect 40 -1802 41 -1801
rect 65 -1802 66 -1801
rect 191 -1802 192 -1801
rect 1206 -1802 1207 -1801
rect 114 -1804 115 -1803
rect 191 -1804 192 -1803
rect 198 -1804 199 -1803
rect 303 -1804 304 -1803
rect 338 -1804 339 -1803
rect 450 -1804 451 -1803
rect 569 -1804 570 -1803
rect 695 -1804 696 -1803
rect 737 -1804 738 -1803
rect 870 -1804 871 -1803
rect 135 -1806 136 -1805
rect 198 -1806 199 -1805
rect 247 -1806 248 -1805
rect 254 -1806 255 -1805
rect 261 -1806 262 -1805
rect 492 -1806 493 -1805
rect 583 -1806 584 -1805
rect 954 -1806 955 -1805
rect 135 -1808 136 -1807
rect 163 -1808 164 -1807
rect 254 -1808 255 -1807
rect 387 -1808 388 -1807
rect 443 -1808 444 -1807
rect 499 -1808 500 -1807
rect 583 -1808 584 -1807
rect 758 -1808 759 -1807
rect 761 -1808 762 -1807
rect 877 -1808 878 -1807
rect 296 -1810 297 -1809
rect 716 -1810 717 -1809
rect 751 -1810 752 -1809
rect 1157 -1810 1158 -1809
rect 310 -1812 311 -1811
rect 758 -1812 759 -1811
rect 765 -1812 766 -1811
rect 800 -1812 801 -1811
rect 877 -1812 878 -1811
rect 905 -1812 906 -1811
rect 1024 -1812 1025 -1811
rect 1157 -1812 1158 -1811
rect 338 -1814 339 -1813
rect 352 -1814 353 -1813
rect 366 -1814 367 -1813
rect 492 -1814 493 -1813
rect 618 -1814 619 -1813
rect 653 -1814 654 -1813
rect 674 -1814 675 -1813
rect 800 -1814 801 -1813
rect 905 -1814 906 -1813
rect 961 -1814 962 -1813
rect 1024 -1814 1025 -1813
rect 1080 -1814 1081 -1813
rect 320 -1816 321 -1815
rect 674 -1816 675 -1815
rect 695 -1816 696 -1815
rect 709 -1816 710 -1815
rect 716 -1816 717 -1815
rect 1150 -1816 1151 -1815
rect 352 -1818 353 -1817
rect 754 -1818 755 -1817
rect 961 -1818 962 -1817
rect 1038 -1818 1039 -1817
rect 1080 -1818 1081 -1817
rect 1136 -1818 1137 -1817
rect 366 -1820 367 -1819
rect 429 -1820 430 -1819
rect 443 -1820 444 -1819
rect 604 -1820 605 -1819
rect 607 -1820 608 -1819
rect 1136 -1820 1137 -1819
rect 23 -1822 24 -1821
rect 429 -1822 430 -1821
rect 485 -1822 486 -1821
rect 754 -1822 755 -1821
rect 1038 -1822 1039 -1821
rect 1066 -1822 1067 -1821
rect 422 -1824 423 -1823
rect 709 -1824 710 -1823
rect 737 -1824 738 -1823
rect 751 -1824 752 -1823
rect 1066 -1824 1067 -1823
rect 1129 -1824 1130 -1823
rect 632 -1826 633 -1825
rect 779 -1826 780 -1825
rect 1129 -1826 1130 -1825
rect 1178 -1826 1179 -1825
rect 639 -1828 640 -1827
rect 1125 -1828 1126 -1827
rect 1178 -1828 1179 -1827
rect 1199 -1828 1200 -1827
rect 653 -1830 654 -1829
rect 814 -1830 815 -1829
rect 1199 -1830 1200 -1829
rect 1262 -1830 1263 -1829
rect 558 -1832 559 -1831
rect 1262 -1832 1263 -1831
rect 779 -1834 780 -1833
rect 786 -1834 787 -1833
rect 194 -1836 195 -1835
rect 786 -1836 787 -1835
rect 2 -1847 3 -1846
rect 523 -1847 524 -1846
rect 604 -1847 605 -1846
rect 646 -1847 647 -1846
rect 653 -1847 654 -1846
rect 695 -1847 696 -1846
rect 712 -1847 713 -1846
rect 877 -1847 878 -1846
rect 16 -1849 17 -1848
rect 387 -1849 388 -1848
rect 432 -1849 433 -1848
rect 1010 -1849 1011 -1848
rect 9 -1851 10 -1850
rect 16 -1851 17 -1850
rect 23 -1851 24 -1850
rect 30 -1851 31 -1850
rect 37 -1851 38 -1850
rect 1178 -1851 1179 -1850
rect 9 -1853 10 -1852
rect 79 -1853 80 -1852
rect 89 -1853 90 -1852
rect 247 -1853 248 -1852
rect 254 -1853 255 -1852
rect 366 -1853 367 -1852
rect 387 -1853 388 -1852
rect 555 -1853 556 -1852
rect 558 -1853 559 -1852
rect 653 -1853 654 -1852
rect 656 -1853 657 -1852
rect 891 -1853 892 -1852
rect 1178 -1853 1179 -1852
rect 1269 -1853 1270 -1852
rect 23 -1855 24 -1854
rect 93 -1855 94 -1854
rect 103 -1855 104 -1854
rect 1094 -1855 1095 -1854
rect 30 -1857 31 -1856
rect 520 -1857 521 -1856
rect 555 -1857 556 -1856
rect 1052 -1857 1053 -1856
rect 1094 -1857 1095 -1856
rect 1241 -1857 1242 -1856
rect 37 -1859 38 -1858
rect 338 -1859 339 -1858
rect 366 -1859 367 -1858
rect 436 -1859 437 -1858
rect 464 -1859 465 -1858
rect 506 -1859 507 -1858
rect 513 -1859 514 -1858
rect 541 -1859 542 -1858
rect 607 -1859 608 -1858
rect 856 -1859 857 -1858
rect 877 -1859 878 -1858
rect 996 -1859 997 -1858
rect 1052 -1859 1053 -1858
rect 1157 -1859 1158 -1858
rect 40 -1861 41 -1860
rect 289 -1861 290 -1860
rect 296 -1861 297 -1860
rect 467 -1861 468 -1860
rect 478 -1861 479 -1860
rect 632 -1861 633 -1860
rect 639 -1861 640 -1860
rect 765 -1861 766 -1860
rect 856 -1861 857 -1860
rect 1059 -1861 1060 -1860
rect 1157 -1861 1158 -1860
rect 1234 -1861 1235 -1860
rect 44 -1863 45 -1862
rect 1003 -1863 1004 -1862
rect 1115 -1863 1116 -1862
rect 1234 -1863 1235 -1862
rect 44 -1865 45 -1864
rect 96 -1865 97 -1864
rect 114 -1865 115 -1864
rect 233 -1865 234 -1864
rect 254 -1865 255 -1864
rect 324 -1865 325 -1864
rect 408 -1865 409 -1864
rect 464 -1865 465 -1864
rect 471 -1865 472 -1864
rect 478 -1865 479 -1864
rect 492 -1865 493 -1864
rect 705 -1865 706 -1864
rect 719 -1865 720 -1864
rect 947 -1865 948 -1864
rect 996 -1865 997 -1864
rect 1080 -1865 1081 -1864
rect 1115 -1865 1116 -1864
rect 1199 -1865 1200 -1864
rect 47 -1867 48 -1866
rect 919 -1867 920 -1866
rect 933 -1867 934 -1866
rect 1059 -1867 1060 -1866
rect 1080 -1867 1081 -1866
rect 1192 -1867 1193 -1866
rect 79 -1869 80 -1868
rect 415 -1869 416 -1868
rect 429 -1869 430 -1868
rect 639 -1869 640 -1868
rect 646 -1869 647 -1868
rect 926 -1869 927 -1868
rect 933 -1869 934 -1868
rect 1031 -1869 1032 -1868
rect 1143 -1869 1144 -1868
rect 1199 -1869 1200 -1868
rect 93 -1871 94 -1870
rect 100 -1871 101 -1870
rect 114 -1871 115 -1870
rect 562 -1871 563 -1870
rect 597 -1871 598 -1870
rect 607 -1871 608 -1870
rect 614 -1871 615 -1870
rect 842 -1871 843 -1870
rect 891 -1871 892 -1870
rect 922 -1871 923 -1870
rect 926 -1871 927 -1870
rect 1185 -1871 1186 -1870
rect 100 -1873 101 -1872
rect 527 -1873 528 -1872
rect 534 -1873 535 -1872
rect 562 -1873 563 -1872
rect 597 -1873 598 -1872
rect 618 -1873 619 -1872
rect 628 -1873 629 -1872
rect 1031 -1873 1032 -1872
rect 1038 -1873 1039 -1872
rect 1185 -1873 1186 -1872
rect 135 -1875 136 -1874
rect 807 -1875 808 -1874
rect 842 -1875 843 -1874
rect 968 -1875 969 -1874
rect 1164 -1875 1165 -1874
rect 1192 -1875 1193 -1874
rect 135 -1877 136 -1876
rect 1143 -1877 1144 -1876
rect 149 -1879 150 -1878
rect 233 -1879 234 -1878
rect 264 -1879 265 -1878
rect 282 -1879 283 -1878
rect 289 -1879 290 -1878
rect 310 -1879 311 -1878
rect 324 -1879 325 -1878
rect 394 -1879 395 -1878
rect 408 -1879 409 -1878
rect 674 -1879 675 -1878
rect 677 -1879 678 -1878
rect 688 -1879 689 -1878
rect 695 -1879 696 -1878
rect 786 -1879 787 -1878
rect 919 -1879 920 -1878
rect 1010 -1879 1011 -1878
rect 1073 -1879 1074 -1878
rect 1164 -1879 1165 -1878
rect 86 -1881 87 -1880
rect 282 -1881 283 -1880
rect 299 -1881 300 -1880
rect 572 -1881 573 -1880
rect 688 -1881 689 -1880
rect 772 -1881 773 -1880
rect 786 -1881 787 -1880
rect 898 -1881 899 -1880
rect 947 -1881 948 -1880
rect 1101 -1881 1102 -1880
rect 86 -1883 87 -1882
rect 1227 -1883 1228 -1882
rect 149 -1885 150 -1884
rect 198 -1885 199 -1884
rect 226 -1885 227 -1884
rect 625 -1885 626 -1884
rect 730 -1885 731 -1884
rect 828 -1885 829 -1884
rect 863 -1885 864 -1884
rect 1101 -1885 1102 -1884
rect 152 -1887 153 -1886
rect 268 -1887 269 -1886
rect 275 -1887 276 -1886
rect 415 -1887 416 -1886
rect 436 -1887 437 -1886
rect 450 -1887 451 -1886
rect 457 -1887 458 -1886
rect 625 -1887 626 -1886
rect 709 -1887 710 -1886
rect 828 -1887 829 -1886
rect 863 -1887 864 -1886
rect 961 -1887 962 -1886
rect 968 -1887 969 -1886
rect 1108 -1887 1109 -1886
rect 163 -1889 164 -1888
rect 296 -1889 297 -1888
rect 303 -1889 304 -1888
rect 310 -1889 311 -1888
rect 352 -1889 353 -1888
rect 961 -1889 962 -1888
rect 1073 -1889 1074 -1888
rect 1255 -1889 1256 -1888
rect 163 -1891 164 -1890
rect 355 -1891 356 -1890
rect 422 -1891 423 -1890
rect 450 -1891 451 -1890
rect 471 -1891 472 -1890
rect 838 -1891 839 -1890
rect 898 -1891 899 -1890
rect 1087 -1891 1088 -1890
rect 177 -1893 178 -1892
rect 268 -1893 269 -1892
rect 275 -1893 276 -1892
rect 1223 -1893 1224 -1892
rect 177 -1895 178 -1894
rect 212 -1895 213 -1894
rect 285 -1895 286 -1894
rect 1108 -1895 1109 -1894
rect 184 -1897 185 -1896
rect 226 -1897 227 -1896
rect 303 -1897 304 -1896
rect 520 -1897 521 -1896
rect 527 -1897 528 -1896
rect 576 -1897 577 -1896
rect 709 -1897 710 -1896
rect 744 -1897 745 -1896
rect 751 -1897 752 -1896
rect 975 -1897 976 -1896
rect 1066 -1897 1067 -1896
rect 1087 -1897 1088 -1896
rect 128 -1899 129 -1898
rect 184 -1899 185 -1898
rect 198 -1899 199 -1898
rect 205 -1899 206 -1898
rect 212 -1899 213 -1898
rect 219 -1899 220 -1898
rect 345 -1899 346 -1898
rect 352 -1899 353 -1898
rect 380 -1899 381 -1898
rect 422 -1899 423 -1898
rect 443 -1899 444 -1898
rect 618 -1899 619 -1898
rect 737 -1899 738 -1898
rect 807 -1899 808 -1898
rect 912 -1899 913 -1898
rect 1227 -1899 1228 -1898
rect 128 -1901 129 -1900
rect 142 -1901 143 -1900
rect 205 -1901 206 -1900
rect 240 -1901 241 -1900
rect 345 -1901 346 -1900
rect 401 -1901 402 -1900
rect 495 -1901 496 -1900
rect 793 -1901 794 -1900
rect 912 -1901 913 -1900
rect 1045 -1901 1046 -1900
rect 1066 -1901 1067 -1900
rect 1171 -1901 1172 -1900
rect 51 -1903 52 -1902
rect 401 -1903 402 -1902
rect 506 -1903 507 -1902
rect 723 -1903 724 -1902
rect 737 -1903 738 -1902
rect 849 -1903 850 -1902
rect 975 -1903 976 -1902
rect 1136 -1903 1137 -1902
rect 1171 -1903 1172 -1902
rect 1262 -1903 1263 -1902
rect 51 -1905 52 -1904
rect 457 -1905 458 -1904
rect 516 -1905 517 -1904
rect 1003 -1905 1004 -1904
rect 1045 -1905 1046 -1904
rect 1150 -1905 1151 -1904
rect 58 -1907 59 -1906
rect 142 -1907 143 -1906
rect 219 -1907 220 -1906
rect 317 -1907 318 -1906
rect 359 -1907 360 -1906
rect 443 -1907 444 -1906
rect 534 -1907 535 -1906
rect 590 -1907 591 -1906
rect 744 -1907 745 -1906
rect 835 -1907 836 -1906
rect 849 -1907 850 -1906
rect 1024 -1907 1025 -1906
rect 1150 -1907 1151 -1906
rect 1248 -1907 1249 -1906
rect 58 -1909 59 -1908
rect 499 -1909 500 -1908
rect 541 -1909 542 -1908
rect 667 -1909 668 -1908
rect 751 -1909 752 -1908
rect 761 -1909 762 -1908
rect 765 -1909 766 -1908
rect 884 -1909 885 -1908
rect 1024 -1909 1025 -1908
rect 1129 -1909 1130 -1908
rect 65 -1911 66 -1910
rect 793 -1911 794 -1910
rect 835 -1911 836 -1910
rect 1213 -1911 1214 -1910
rect 138 -1913 139 -1912
rect 723 -1913 724 -1912
rect 754 -1913 755 -1912
rect 940 -1913 941 -1912
rect 1213 -1913 1214 -1912
rect 1276 -1913 1277 -1912
rect 138 -1915 139 -1914
rect 156 -1915 157 -1914
rect 191 -1915 192 -1914
rect 499 -1915 500 -1914
rect 548 -1915 549 -1914
rect 632 -1915 633 -1914
rect 667 -1915 668 -1914
rect 702 -1915 703 -1914
rect 758 -1915 759 -1914
rect 779 -1915 780 -1914
rect 156 -1917 157 -1916
rect 481 -1917 482 -1916
rect 548 -1917 549 -1916
rect 642 -1917 643 -1916
rect 702 -1917 703 -1916
rect 1038 -1917 1039 -1916
rect 191 -1919 192 -1918
rect 369 -1919 370 -1918
rect 380 -1919 381 -1918
rect 604 -1919 605 -1918
rect 761 -1919 762 -1918
rect 884 -1919 885 -1918
rect 72 -1921 73 -1920
rect 369 -1921 370 -1920
rect 429 -1921 430 -1920
rect 1136 -1921 1137 -1920
rect 68 -1923 69 -1922
rect 72 -1923 73 -1922
rect 240 -1923 241 -1922
rect 261 -1923 262 -1922
rect 317 -1923 318 -1922
rect 338 -1923 339 -1922
rect 359 -1923 360 -1922
rect 583 -1923 584 -1922
rect 590 -1923 591 -1922
rect 660 -1923 661 -1922
rect 772 -1923 773 -1922
rect 989 -1923 990 -1922
rect 54 -1925 55 -1924
rect 68 -1925 69 -1924
rect 107 -1925 108 -1924
rect 261 -1925 262 -1924
rect 320 -1925 321 -1924
rect 660 -1925 661 -1924
rect 779 -1925 780 -1924
rect 821 -1925 822 -1924
rect 107 -1927 108 -1926
rect 121 -1927 122 -1926
rect 247 -1927 248 -1926
rect 758 -1927 759 -1926
rect 821 -1927 822 -1926
rect 954 -1927 955 -1926
rect 121 -1929 122 -1928
rect 170 -1929 171 -1928
rect 460 -1929 461 -1928
rect 1129 -1929 1130 -1928
rect 170 -1931 171 -1930
rect 394 -1931 395 -1930
rect 492 -1931 493 -1930
rect 989 -1931 990 -1930
rect 569 -1933 570 -1932
rect 583 -1933 584 -1932
rect 954 -1933 955 -1932
rect 1220 -1933 1221 -1932
rect 569 -1935 570 -1934
rect 940 -1935 941 -1934
rect 576 -1937 577 -1936
rect 814 -1937 815 -1936
rect 814 -1939 815 -1938
rect 870 -1939 871 -1938
rect 870 -1941 871 -1940
rect 982 -1941 983 -1940
rect 611 -1943 612 -1942
rect 982 -1943 983 -1942
rect 611 -1945 612 -1944
rect 681 -1945 682 -1944
rect 681 -1947 682 -1946
rect 716 -1947 717 -1946
rect 716 -1949 717 -1948
rect 800 -1949 801 -1948
rect 800 -1951 801 -1950
rect 905 -1951 906 -1950
rect 905 -1953 906 -1952
rect 1017 -1953 1018 -1952
rect 1017 -1955 1018 -1954
rect 1122 -1955 1123 -1954
rect 1122 -1957 1123 -1956
rect 1206 -1957 1207 -1956
rect 586 -1959 587 -1958
rect 1206 -1959 1207 -1958
rect 2 -1970 3 -1969
rect 646 -1970 647 -1969
rect 674 -1970 675 -1969
rect 954 -1970 955 -1969
rect 964 -1970 965 -1969
rect 1094 -1970 1095 -1969
rect 1164 -1970 1165 -1969
rect 1220 -1970 1221 -1969
rect 9 -1972 10 -1971
rect 135 -1972 136 -1971
rect 142 -1972 143 -1971
rect 285 -1972 286 -1971
rect 310 -1972 311 -1971
rect 317 -1972 318 -1971
rect 320 -1972 321 -1971
rect 331 -1972 332 -1971
rect 373 -1972 374 -1971
rect 376 -1972 377 -1971
rect 401 -1972 402 -1971
rect 674 -1972 675 -1971
rect 702 -1972 703 -1971
rect 1101 -1972 1102 -1971
rect 9 -1974 10 -1973
rect 166 -1974 167 -1973
rect 184 -1974 185 -1973
rect 492 -1974 493 -1973
rect 499 -1974 500 -1973
rect 621 -1974 622 -1973
rect 702 -1974 703 -1973
rect 737 -1974 738 -1973
rect 758 -1974 759 -1973
rect 1087 -1974 1088 -1973
rect 1094 -1974 1095 -1973
rect 1136 -1974 1137 -1973
rect 16 -1976 17 -1975
rect 261 -1976 262 -1975
rect 282 -1976 283 -1975
rect 457 -1976 458 -1975
rect 464 -1976 465 -1975
rect 492 -1976 493 -1975
rect 499 -1976 500 -1975
rect 1213 -1976 1214 -1975
rect 37 -1978 38 -1977
rect 173 -1978 174 -1977
rect 184 -1978 185 -1977
rect 324 -1978 325 -1977
rect 331 -1978 332 -1977
rect 394 -1978 395 -1977
rect 408 -1978 409 -1977
rect 411 -1978 412 -1977
rect 464 -1978 465 -1977
rect 541 -1978 542 -1977
rect 569 -1978 570 -1977
rect 716 -1978 717 -1977
rect 737 -1978 738 -1977
rect 891 -1978 892 -1977
rect 919 -1978 920 -1977
rect 996 -1978 997 -1977
rect 1027 -1978 1028 -1977
rect 1192 -1978 1193 -1977
rect 37 -1980 38 -1979
rect 163 -1980 164 -1979
rect 191 -1980 192 -1979
rect 369 -1980 370 -1979
rect 373 -1980 374 -1979
rect 380 -1980 381 -1979
rect 394 -1980 395 -1979
rect 688 -1980 689 -1979
rect 716 -1980 717 -1979
rect 800 -1980 801 -1979
rect 891 -1980 892 -1979
rect 933 -1980 934 -1979
rect 954 -1980 955 -1979
rect 961 -1980 962 -1979
rect 968 -1980 969 -1979
rect 971 -1980 972 -1979
rect 996 -1980 997 -1979
rect 1122 -1980 1123 -1979
rect 16 -1982 17 -1981
rect 163 -1982 164 -1981
rect 198 -1982 199 -1981
rect 429 -1982 430 -1981
rect 481 -1982 482 -1981
rect 1010 -1982 1011 -1981
rect 1073 -1982 1074 -1981
rect 1122 -1982 1123 -1981
rect 51 -1984 52 -1983
rect 240 -1984 241 -1983
rect 243 -1984 244 -1983
rect 688 -1984 689 -1983
rect 758 -1984 759 -1983
rect 786 -1984 787 -1983
rect 800 -1984 801 -1983
rect 842 -1984 843 -1983
rect 919 -1984 920 -1983
rect 940 -1984 941 -1983
rect 968 -1984 969 -1983
rect 975 -1984 976 -1983
rect 1010 -1984 1011 -1983
rect 1143 -1984 1144 -1983
rect 54 -1986 55 -1985
rect 744 -1986 745 -1985
rect 761 -1986 762 -1985
rect 989 -1986 990 -1985
rect 1059 -1986 1060 -1985
rect 1143 -1986 1144 -1985
rect 58 -1988 59 -1987
rect 457 -1988 458 -1987
rect 488 -1988 489 -1987
rect 772 -1988 773 -1987
rect 786 -1988 787 -1987
rect 870 -1988 871 -1987
rect 940 -1988 941 -1987
rect 947 -1988 948 -1987
rect 982 -1988 983 -1987
rect 1059 -1988 1060 -1987
rect 1073 -1988 1074 -1987
rect 1108 -1988 1109 -1987
rect 58 -1990 59 -1989
rect 366 -1990 367 -1989
rect 408 -1990 409 -1989
rect 415 -1990 416 -1989
rect 429 -1990 430 -1989
rect 478 -1990 479 -1989
rect 502 -1990 503 -1989
rect 646 -1990 647 -1989
rect 677 -1990 678 -1989
rect 961 -1990 962 -1989
rect 982 -1990 983 -1989
rect 1045 -1990 1046 -1989
rect 1087 -1990 1088 -1989
rect 1227 -1990 1228 -1989
rect 65 -1992 66 -1991
rect 96 -1992 97 -1991
rect 100 -1992 101 -1991
rect 289 -1992 290 -1991
rect 310 -1992 311 -1991
rect 597 -1992 598 -1991
rect 604 -1992 605 -1991
rect 1199 -1992 1200 -1991
rect 23 -1994 24 -1993
rect 96 -1994 97 -1993
rect 110 -1994 111 -1993
rect 485 -1994 486 -1993
rect 513 -1994 514 -1993
rect 558 -1994 559 -1993
rect 569 -1994 570 -1993
rect 611 -1994 612 -1993
rect 744 -1994 745 -1993
rect 835 -1994 836 -1993
rect 842 -1994 843 -1993
rect 1017 -1994 1018 -1993
rect 1101 -1994 1102 -1993
rect 1171 -1994 1172 -1993
rect 23 -1996 24 -1995
rect 506 -1996 507 -1995
rect 520 -1996 521 -1995
rect 898 -1996 899 -1995
rect 947 -1996 948 -1995
rect 1003 -1996 1004 -1995
rect 1017 -1996 1018 -1995
rect 1066 -1996 1067 -1995
rect 1108 -1996 1109 -1995
rect 1178 -1996 1179 -1995
rect 44 -1998 45 -1997
rect 65 -1998 66 -1997
rect 68 -1998 69 -1997
rect 730 -1998 731 -1997
rect 772 -1998 773 -1997
rect 838 -1998 839 -1997
rect 849 -1998 850 -1997
rect 870 -1998 871 -1997
rect 898 -1998 899 -1997
rect 1038 -1998 1039 -1997
rect 1066 -1998 1067 -1997
rect 1080 -1998 1081 -1997
rect 72 -2000 73 -1999
rect 663 -2000 664 -1999
rect 835 -2000 836 -1999
rect 877 -2000 878 -1999
rect 971 -2000 972 -1999
rect 975 -2000 976 -1999
rect 989 -2000 990 -1999
rect 1024 -2000 1025 -1999
rect 1031 -2000 1032 -1999
rect 1038 -2000 1039 -1999
rect 1080 -2000 1081 -1999
rect 1115 -2000 1116 -1999
rect 72 -2002 73 -2001
rect 107 -2002 108 -2001
rect 114 -2002 115 -2001
rect 366 -2002 367 -2001
rect 478 -2002 479 -2001
rect 730 -2002 731 -2001
rect 877 -2002 878 -2001
rect 884 -2002 885 -2001
rect 1003 -2002 1004 -2001
rect 1052 -2002 1053 -2001
rect 1115 -2002 1116 -2001
rect 1206 -2002 1207 -2001
rect 86 -2004 87 -2003
rect 135 -2004 136 -2003
rect 142 -2004 143 -2003
rect 268 -2004 269 -2003
rect 282 -2004 283 -2003
rect 450 -2004 451 -2003
rect 506 -2004 507 -2003
rect 698 -2004 699 -2003
rect 926 -2004 927 -2003
rect 1052 -2004 1053 -2003
rect 86 -2006 87 -2005
rect 562 -2006 563 -2005
rect 576 -2006 577 -2005
rect 884 -2006 885 -2005
rect 1031 -2006 1032 -2005
rect 1150 -2006 1151 -2005
rect 44 -2008 45 -2007
rect 576 -2008 577 -2007
rect 579 -2008 580 -2007
rect 814 -2008 815 -2007
rect 856 -2008 857 -2007
rect 926 -2008 927 -2007
rect 1136 -2008 1137 -2007
rect 1150 -2008 1151 -2007
rect 51 -2010 52 -2009
rect 814 -2010 815 -2009
rect 856 -2010 857 -2009
rect 905 -2010 906 -2009
rect 89 -2012 90 -2011
rect 107 -2012 108 -2011
rect 117 -2012 118 -2011
rect 212 -2012 213 -2011
rect 226 -2012 227 -2011
rect 278 -2012 279 -2011
rect 317 -2012 318 -2011
rect 345 -2012 346 -2011
rect 450 -2012 451 -2011
rect 471 -2012 472 -2011
rect 534 -2012 535 -2011
rect 933 -2012 934 -2011
rect 93 -2014 94 -2013
rect 709 -2014 710 -2013
rect 905 -2014 906 -2013
rect 912 -2014 913 -2013
rect 93 -2016 94 -2015
rect 303 -2016 304 -2015
rect 338 -2016 339 -2015
rect 604 -2016 605 -2015
rect 611 -2016 612 -2015
rect 625 -2016 626 -2015
rect 709 -2016 710 -2015
rect 765 -2016 766 -2015
rect 30 -2018 31 -2017
rect 303 -2018 304 -2017
rect 471 -2018 472 -2017
rect 548 -2018 549 -2017
rect 562 -2018 563 -2017
rect 681 -2018 682 -2017
rect 751 -2018 752 -2017
rect 912 -2018 913 -2017
rect 30 -2020 31 -2019
rect 359 -2020 360 -2019
rect 534 -2020 535 -2019
rect 590 -2020 591 -2019
rect 597 -2020 598 -2019
rect 632 -2020 633 -2019
rect 681 -2020 682 -2019
rect 695 -2020 696 -2019
rect 751 -2020 752 -2019
rect 779 -2020 780 -2019
rect 114 -2022 115 -2021
rect 338 -2022 339 -2021
rect 432 -2022 433 -2021
rect 590 -2022 591 -2021
rect 625 -2022 626 -2021
rect 660 -2022 661 -2021
rect 765 -2022 766 -2021
rect 821 -2022 822 -2021
rect 121 -2024 122 -2023
rect 520 -2024 521 -2023
rect 541 -2024 542 -2023
rect 583 -2024 584 -2023
rect 632 -2024 633 -2023
rect 639 -2024 640 -2023
rect 660 -2024 661 -2023
rect 667 -2024 668 -2023
rect 821 -2024 822 -2023
rect 863 -2024 864 -2023
rect 103 -2026 104 -2025
rect 667 -2026 668 -2025
rect 863 -2026 864 -2025
rect 1185 -2026 1186 -2025
rect 121 -2028 122 -2027
rect 653 -2028 654 -2027
rect 1185 -2028 1186 -2027
rect 1234 -2028 1235 -2027
rect 128 -2030 129 -2029
rect 572 -2030 573 -2029
rect 583 -2030 584 -2029
rect 779 -2030 780 -2029
rect 152 -2032 153 -2031
rect 849 -2032 850 -2031
rect 170 -2034 171 -2033
rect 345 -2034 346 -2033
rect 548 -2034 549 -2033
rect 618 -2034 619 -2033
rect 639 -2034 640 -2033
rect 1024 -2034 1025 -2033
rect 149 -2036 150 -2035
rect 170 -2036 171 -2035
rect 177 -2036 178 -2035
rect 212 -2036 213 -2035
rect 226 -2036 227 -2035
rect 275 -2036 276 -2035
rect 618 -2036 619 -2035
rect 1045 -2036 1046 -2035
rect 128 -2038 129 -2037
rect 149 -2038 150 -2037
rect 177 -2038 178 -2037
rect 695 -2038 696 -2037
rect 191 -2040 192 -2039
rect 240 -2040 241 -2039
rect 247 -2040 248 -2039
rect 513 -2040 514 -2039
rect 653 -2040 654 -2039
rect 807 -2040 808 -2039
rect 198 -2042 199 -2041
rect 387 -2042 388 -2041
rect 807 -2042 808 -2041
rect 828 -2042 829 -2041
rect 205 -2044 206 -2043
rect 261 -2044 262 -2043
rect 268 -2044 269 -2043
rect 352 -2044 353 -2043
rect 828 -2044 829 -2043
rect 1129 -2044 1130 -2043
rect 156 -2046 157 -2045
rect 205 -2046 206 -2045
rect 233 -2046 234 -2045
rect 359 -2046 360 -2045
rect 723 -2046 724 -2045
rect 1129 -2046 1130 -2045
rect 79 -2048 80 -2047
rect 156 -2048 157 -2047
rect 233 -2048 234 -2047
rect 523 -2048 524 -2047
rect 723 -2048 724 -2047
rect 793 -2048 794 -2047
rect 79 -2050 80 -2049
rect 334 -2050 335 -2049
rect 352 -2050 353 -2049
rect 422 -2050 423 -2049
rect 555 -2050 556 -2049
rect 793 -2050 794 -2049
rect 247 -2052 248 -2051
rect 460 -2052 461 -2051
rect 555 -2052 556 -2051
rect 1223 -2052 1224 -2051
rect 254 -2054 255 -2053
rect 289 -2054 290 -2053
rect 296 -2054 297 -2053
rect 387 -2054 388 -2053
rect 422 -2054 423 -2053
rect 527 -2054 528 -2053
rect 138 -2056 139 -2055
rect 296 -2056 297 -2055
rect 436 -2056 437 -2055
rect 527 -2056 528 -2055
rect 219 -2058 220 -2057
rect 254 -2058 255 -2057
rect 275 -2058 276 -2057
rect 401 -2058 402 -2057
rect 436 -2058 437 -2057
rect 443 -2058 444 -2057
rect 89 -2060 90 -2059
rect 443 -2060 444 -2059
rect 219 -2062 220 -2061
rect 607 -2062 608 -2061
rect 2 -2073 3 -2072
rect 93 -2073 94 -2072
rect 103 -2073 104 -2072
rect 744 -2073 745 -2072
rect 789 -2073 790 -2072
rect 1122 -2073 1123 -2072
rect 1136 -2073 1137 -2072
rect 1185 -2073 1186 -2072
rect 30 -2075 31 -2074
rect 243 -2075 244 -2074
rect 247 -2075 248 -2074
rect 278 -2075 279 -2074
rect 394 -2075 395 -2074
rect 618 -2075 619 -2074
rect 621 -2075 622 -2074
rect 800 -2075 801 -2074
rect 817 -2075 818 -2074
rect 975 -2075 976 -2074
rect 1122 -2075 1123 -2074
rect 1150 -2075 1151 -2074
rect 30 -2077 31 -2076
rect 86 -2077 87 -2076
rect 93 -2077 94 -2076
rect 163 -2077 164 -2076
rect 166 -2077 167 -2076
rect 996 -2077 997 -2076
rect 1139 -2077 1140 -2076
rect 1157 -2077 1158 -2076
rect 37 -2079 38 -2078
rect 324 -2079 325 -2078
rect 394 -2079 395 -2078
rect 471 -2079 472 -2078
rect 481 -2079 482 -2078
rect 527 -2079 528 -2078
rect 562 -2079 563 -2078
rect 565 -2079 566 -2078
rect 576 -2079 577 -2078
rect 877 -2079 878 -2078
rect 975 -2079 976 -2078
rect 1038 -2079 1039 -2078
rect 65 -2081 66 -2080
rect 152 -2081 153 -2080
rect 156 -2081 157 -2080
rect 499 -2081 500 -2080
rect 509 -2081 510 -2080
rect 639 -2081 640 -2080
rect 653 -2081 654 -2080
rect 1024 -2081 1025 -2080
rect 65 -2083 66 -2082
rect 296 -2083 297 -2082
rect 387 -2083 388 -2082
rect 481 -2083 482 -2082
rect 492 -2083 493 -2082
rect 530 -2083 531 -2082
rect 562 -2083 563 -2082
rect 590 -2083 591 -2082
rect 600 -2083 601 -2082
rect 632 -2083 633 -2082
rect 639 -2083 640 -2082
rect 884 -2083 885 -2082
rect 86 -2085 87 -2084
rect 135 -2085 136 -2084
rect 138 -2085 139 -2084
rect 793 -2085 794 -2084
rect 863 -2085 864 -2084
rect 1087 -2085 1088 -2084
rect 37 -2087 38 -2086
rect 135 -2087 136 -2086
rect 142 -2087 143 -2086
rect 488 -2087 489 -2086
rect 565 -2087 566 -2086
rect 590 -2087 591 -2086
rect 614 -2087 615 -2086
rect 996 -2087 997 -2086
rect 100 -2089 101 -2088
rect 247 -2089 248 -2088
rect 254 -2089 255 -2088
rect 299 -2089 300 -2088
rect 387 -2089 388 -2088
rect 450 -2089 451 -2088
rect 457 -2089 458 -2088
rect 499 -2089 500 -2088
rect 576 -2089 577 -2088
rect 625 -2089 626 -2088
rect 632 -2089 633 -2088
rect 667 -2089 668 -2088
rect 695 -2089 696 -2088
rect 758 -2089 759 -2088
rect 793 -2089 794 -2088
rect 1129 -2089 1130 -2088
rect 100 -2091 101 -2090
rect 163 -2091 164 -2090
rect 170 -2091 171 -2090
rect 240 -2091 241 -2090
rect 254 -2091 255 -2090
rect 289 -2091 290 -2090
rect 401 -2091 402 -2090
rect 492 -2091 493 -2090
rect 579 -2091 580 -2090
rect 611 -2091 612 -2090
rect 618 -2091 619 -2090
rect 674 -2091 675 -2090
rect 695 -2091 696 -2090
rect 947 -2091 948 -2090
rect 107 -2093 108 -2092
rect 114 -2093 115 -2092
rect 117 -2093 118 -2092
rect 282 -2093 283 -2092
rect 289 -2093 290 -2092
rect 303 -2093 304 -2092
rect 401 -2093 402 -2092
rect 464 -2093 465 -2092
rect 467 -2093 468 -2092
rect 1038 -2093 1039 -2092
rect 58 -2095 59 -2094
rect 107 -2095 108 -2094
rect 114 -2095 115 -2094
rect 380 -2095 381 -2094
rect 429 -2095 430 -2094
rect 450 -2095 451 -2094
rect 457 -2095 458 -2094
rect 646 -2095 647 -2094
rect 656 -2095 657 -2094
rect 709 -2095 710 -2094
rect 716 -2095 717 -2094
rect 800 -2095 801 -2094
rect 863 -2095 864 -2094
rect 926 -2095 927 -2094
rect 947 -2095 948 -2094
rect 1101 -2095 1102 -2094
rect 23 -2097 24 -2096
rect 58 -2097 59 -2096
rect 142 -2097 143 -2096
rect 233 -2097 234 -2096
rect 240 -2097 241 -2096
rect 334 -2097 335 -2096
rect 373 -2097 374 -2096
rect 380 -2097 381 -2096
rect 408 -2097 409 -2096
rect 646 -2097 647 -2096
rect 660 -2097 661 -2096
rect 842 -2097 843 -2096
rect 877 -2097 878 -2096
rect 954 -2097 955 -2096
rect 23 -2099 24 -2098
rect 89 -2099 90 -2098
rect 96 -2099 97 -2098
rect 373 -2099 374 -2098
rect 429 -2099 430 -2098
rect 436 -2099 437 -2098
rect 443 -2099 444 -2098
rect 611 -2099 612 -2098
rect 625 -2099 626 -2098
rect 688 -2099 689 -2098
rect 709 -2099 710 -2098
rect 807 -2099 808 -2098
rect 842 -2099 843 -2098
rect 891 -2099 892 -2098
rect 926 -2099 927 -2098
rect 982 -2099 983 -2098
rect 149 -2101 150 -2100
rect 485 -2101 486 -2100
rect 583 -2101 584 -2100
rect 912 -2101 913 -2100
rect 933 -2101 934 -2100
rect 954 -2101 955 -2100
rect 982 -2101 983 -2100
rect 1066 -2101 1067 -2100
rect 44 -2103 45 -2102
rect 149 -2103 150 -2102
rect 156 -2103 157 -2102
rect 219 -2103 220 -2102
rect 233 -2103 234 -2102
rect 317 -2103 318 -2102
rect 345 -2103 346 -2102
rect 408 -2103 409 -2102
rect 443 -2103 444 -2102
rect 691 -2103 692 -2102
rect 716 -2103 717 -2102
rect 772 -2103 773 -2102
rect 807 -2103 808 -2102
rect 821 -2103 822 -2102
rect 884 -2103 885 -2102
rect 961 -2103 962 -2102
rect 1066 -2103 1067 -2102
rect 1080 -2103 1081 -2102
rect 44 -2105 45 -2104
rect 698 -2105 699 -2104
rect 737 -2105 738 -2104
rect 758 -2105 759 -2104
rect 772 -2105 773 -2104
rect 786 -2105 787 -2104
rect 821 -2105 822 -2104
rect 905 -2105 906 -2104
rect 933 -2105 934 -2104
rect 1017 -2105 1018 -2104
rect 51 -2107 52 -2106
rect 219 -2107 220 -2106
rect 261 -2107 262 -2106
rect 320 -2107 321 -2106
rect 338 -2107 339 -2106
rect 961 -2107 962 -2106
rect 1017 -2107 1018 -2106
rect 1115 -2107 1116 -2106
rect 16 -2109 17 -2108
rect 51 -2109 52 -2108
rect 173 -2109 174 -2108
rect 681 -2109 682 -2108
rect 737 -2109 738 -2108
rect 765 -2109 766 -2108
rect 891 -2109 892 -2108
rect 968 -2109 969 -2108
rect 110 -2111 111 -2110
rect 765 -2111 766 -2110
rect 898 -2111 899 -2110
rect 912 -2111 913 -2110
rect 968 -2111 969 -2110
rect 1031 -2111 1032 -2110
rect 184 -2113 185 -2112
rect 282 -2113 283 -2112
rect 303 -2113 304 -2112
rect 516 -2113 517 -2112
rect 583 -2113 584 -2112
rect 597 -2113 598 -2112
rect 660 -2113 661 -2112
rect 663 -2113 664 -2112
rect 667 -2113 668 -2112
rect 702 -2113 703 -2112
rect 744 -2113 745 -2112
rect 751 -2113 752 -2112
rect 814 -2113 815 -2112
rect 898 -2113 899 -2112
rect 905 -2113 906 -2112
rect 1059 -2113 1060 -2112
rect 184 -2115 185 -2114
rect 534 -2115 535 -2114
rect 674 -2115 675 -2114
rect 723 -2115 724 -2114
rect 751 -2115 752 -2114
rect 779 -2115 780 -2114
rect 814 -2115 815 -2114
rect 856 -2115 857 -2114
rect 866 -2115 867 -2114
rect 1059 -2115 1060 -2114
rect 205 -2117 206 -2116
rect 324 -2117 325 -2116
rect 338 -2117 339 -2116
rect 502 -2117 503 -2116
rect 681 -2117 682 -2116
rect 849 -2117 850 -2116
rect 856 -2117 857 -2116
rect 1003 -2117 1004 -2116
rect 1031 -2117 1032 -2116
rect 1104 -2117 1105 -2116
rect 205 -2119 206 -2118
rect 226 -2119 227 -2118
rect 261 -2119 262 -2118
rect 527 -2119 528 -2118
rect 702 -2119 703 -2118
rect 870 -2119 871 -2118
rect 1003 -2119 1004 -2118
rect 1143 -2119 1144 -2118
rect 79 -2121 80 -2120
rect 226 -2121 227 -2120
rect 268 -2121 269 -2120
rect 331 -2121 332 -2120
rect 345 -2121 346 -2120
rect 422 -2121 423 -2120
rect 471 -2121 472 -2120
rect 548 -2121 549 -2120
rect 723 -2121 724 -2120
rect 835 -2121 836 -2120
rect 849 -2121 850 -2120
rect 1052 -2121 1053 -2120
rect 79 -2123 80 -2122
rect 478 -2123 479 -2122
rect 548 -2123 549 -2122
rect 642 -2123 643 -2122
rect 730 -2123 731 -2122
rect 779 -2123 780 -2122
rect 835 -2123 836 -2122
rect 1045 -2123 1046 -2122
rect 1052 -2123 1053 -2122
rect 1101 -2123 1102 -2122
rect 128 -2125 129 -2124
rect 331 -2125 332 -2124
rect 352 -2125 353 -2124
rect 436 -2125 437 -2124
rect 478 -2125 479 -2124
rect 989 -2125 990 -2124
rect 128 -2127 129 -2126
rect 177 -2127 178 -2126
rect 212 -2127 213 -2126
rect 327 -2127 328 -2126
rect 352 -2127 353 -2126
rect 513 -2127 514 -2126
rect 597 -2127 598 -2126
rect 1045 -2127 1046 -2126
rect 9 -2129 10 -2128
rect 513 -2129 514 -2128
rect 730 -2129 731 -2128
rect 828 -2129 829 -2128
rect 870 -2129 871 -2128
rect 940 -2129 941 -2128
rect 989 -2129 990 -2128
rect 1073 -2129 1074 -2128
rect 177 -2131 178 -2130
rect 191 -2131 192 -2130
rect 212 -2131 213 -2130
rect 359 -2131 360 -2130
rect 366 -2131 367 -2130
rect 422 -2131 423 -2130
rect 485 -2131 486 -2130
rect 940 -2131 941 -2130
rect 121 -2133 122 -2132
rect 191 -2133 192 -2132
rect 268 -2133 269 -2132
rect 506 -2133 507 -2132
rect 828 -2133 829 -2132
rect 919 -2133 920 -2132
rect 117 -2135 118 -2134
rect 121 -2135 122 -2134
rect 275 -2135 276 -2134
rect 555 -2135 556 -2134
rect 919 -2135 920 -2134
rect 1094 -2135 1095 -2134
rect 310 -2137 311 -2136
rect 534 -2137 535 -2136
rect 555 -2137 556 -2136
rect 569 -2137 570 -2136
rect 198 -2139 199 -2138
rect 310 -2139 311 -2138
rect 359 -2139 360 -2138
rect 415 -2139 416 -2138
rect 464 -2139 465 -2138
rect 569 -2139 570 -2138
rect 198 -2141 199 -2140
rect 317 -2141 318 -2140
rect 366 -2141 367 -2140
rect 520 -2141 521 -2140
rect 415 -2143 416 -2142
rect 604 -2143 605 -2142
rect 520 -2145 521 -2144
rect 541 -2145 542 -2144
rect 604 -2145 605 -2144
rect 688 -2145 689 -2144
rect 541 -2147 542 -2146
rect 786 -2147 787 -2146
rect 23 -2158 24 -2157
rect 117 -2158 118 -2157
rect 124 -2158 125 -2157
rect 303 -2158 304 -2157
rect 317 -2158 318 -2157
rect 324 -2158 325 -2157
rect 331 -2158 332 -2157
rect 971 -2158 972 -2157
rect 975 -2158 976 -2157
rect 996 -2158 997 -2157
rect 1101 -2158 1102 -2157
rect 1108 -2158 1109 -2157
rect 37 -2160 38 -2159
rect 100 -2160 101 -2159
rect 103 -2160 104 -2159
rect 156 -2160 157 -2159
rect 198 -2160 199 -2159
rect 303 -2160 304 -2159
rect 324 -2160 325 -2159
rect 380 -2160 381 -2159
rect 387 -2160 388 -2159
rect 488 -2160 489 -2159
rect 509 -2160 510 -2159
rect 849 -2160 850 -2159
rect 933 -2160 934 -2159
rect 968 -2160 969 -2159
rect 982 -2160 983 -2159
rect 996 -2160 997 -2159
rect 1104 -2160 1105 -2159
rect 1122 -2160 1123 -2159
rect 37 -2162 38 -2161
rect 86 -2162 87 -2161
rect 93 -2162 94 -2161
rect 261 -2162 262 -2161
rect 275 -2162 276 -2161
rect 464 -2162 465 -2161
rect 485 -2162 486 -2161
rect 583 -2162 584 -2161
rect 597 -2162 598 -2161
rect 702 -2162 703 -2161
rect 786 -2162 787 -2161
rect 898 -2162 899 -2161
rect 933 -2162 934 -2161
rect 1038 -2162 1039 -2161
rect 30 -2164 31 -2163
rect 93 -2164 94 -2163
rect 100 -2164 101 -2163
rect 142 -2164 143 -2163
rect 198 -2164 199 -2163
rect 247 -2164 248 -2163
rect 254 -2164 255 -2163
rect 467 -2164 468 -2163
rect 513 -2164 514 -2163
rect 695 -2164 696 -2163
rect 702 -2164 703 -2163
rect 737 -2164 738 -2163
rect 786 -2164 787 -2163
rect 884 -2164 885 -2163
rect 943 -2164 944 -2163
rect 1059 -2164 1060 -2163
rect 30 -2166 31 -2165
rect 527 -2166 528 -2165
rect 597 -2166 598 -2165
rect 632 -2166 633 -2165
rect 639 -2166 640 -2165
rect 674 -2166 675 -2165
rect 688 -2166 689 -2165
rect 919 -2166 920 -2165
rect 982 -2166 983 -2165
rect 1003 -2166 1004 -2165
rect 51 -2168 52 -2167
rect 156 -2168 157 -2167
rect 233 -2168 234 -2167
rect 478 -2168 479 -2167
rect 513 -2168 514 -2167
rect 541 -2168 542 -2167
rect 611 -2168 612 -2167
rect 954 -2168 955 -2167
rect 1003 -2168 1004 -2167
rect 1052 -2168 1053 -2167
rect 44 -2170 45 -2169
rect 51 -2170 52 -2169
rect 65 -2170 66 -2169
rect 261 -2170 262 -2169
rect 289 -2170 290 -2169
rect 488 -2170 489 -2169
rect 541 -2170 542 -2169
rect 569 -2170 570 -2169
rect 611 -2170 612 -2169
rect 698 -2170 699 -2169
rect 842 -2170 843 -2169
rect 975 -2170 976 -2169
rect 58 -2172 59 -2171
rect 65 -2172 66 -2171
rect 72 -2172 73 -2171
rect 135 -2172 136 -2171
rect 138 -2172 139 -2171
rect 583 -2172 584 -2171
rect 614 -2172 615 -2171
rect 898 -2172 899 -2171
rect 919 -2172 920 -2171
rect 1031 -2172 1032 -2171
rect 58 -2174 59 -2173
rect 397 -2174 398 -2173
rect 408 -2174 409 -2173
rect 481 -2174 482 -2173
rect 632 -2174 633 -2173
rect 709 -2174 710 -2173
rect 842 -2174 843 -2173
rect 961 -2174 962 -2173
rect 72 -2176 73 -2175
rect 184 -2176 185 -2175
rect 240 -2176 241 -2175
rect 247 -2176 248 -2175
rect 254 -2176 255 -2175
rect 268 -2176 269 -2175
rect 289 -2176 290 -2175
rect 394 -2176 395 -2175
rect 401 -2176 402 -2175
rect 408 -2176 409 -2175
rect 429 -2176 430 -2175
rect 506 -2176 507 -2175
rect 646 -2176 647 -2175
rect 884 -2176 885 -2175
rect 96 -2178 97 -2177
rect 184 -2178 185 -2177
rect 205 -2178 206 -2177
rect 240 -2178 241 -2177
rect 268 -2178 269 -2177
rect 789 -2178 790 -2177
rect 96 -2180 97 -2179
rect 656 -2180 657 -2179
rect 674 -2180 675 -2179
rect 681 -2180 682 -2179
rect 688 -2180 689 -2179
rect 765 -2180 766 -2179
rect 114 -2182 115 -2181
rect 275 -2182 276 -2181
rect 296 -2182 297 -2181
rect 331 -2182 332 -2181
rect 355 -2182 356 -2181
rect 604 -2182 605 -2181
rect 646 -2182 647 -2181
rect 667 -2182 668 -2181
rect 681 -2182 682 -2181
rect 758 -2182 759 -2181
rect 114 -2184 115 -2183
rect 121 -2184 122 -2183
rect 131 -2184 132 -2183
rect 359 -2184 360 -2183
rect 366 -2184 367 -2183
rect 394 -2184 395 -2183
rect 401 -2184 402 -2183
rect 450 -2184 451 -2183
rect 464 -2184 465 -2183
rect 499 -2184 500 -2183
rect 506 -2184 507 -2183
rect 555 -2184 556 -2183
rect 604 -2184 605 -2183
rect 747 -2184 748 -2183
rect 751 -2184 752 -2183
rect 961 -2184 962 -2183
rect 121 -2186 122 -2185
rect 443 -2186 444 -2185
rect 457 -2186 458 -2185
rect 555 -2186 556 -2185
rect 656 -2186 657 -2185
rect 856 -2186 857 -2185
rect 135 -2188 136 -2187
rect 219 -2188 220 -2187
rect 282 -2188 283 -2187
rect 296 -2188 297 -2187
rect 310 -2188 311 -2187
rect 366 -2188 367 -2187
rect 373 -2188 374 -2187
rect 429 -2188 430 -2187
rect 443 -2188 444 -2187
rect 492 -2188 493 -2187
rect 499 -2188 500 -2187
rect 530 -2188 531 -2187
rect 691 -2188 692 -2187
rect 800 -2188 801 -2187
rect 856 -2188 857 -2187
rect 905 -2188 906 -2187
rect 79 -2190 80 -2189
rect 282 -2190 283 -2189
rect 310 -2190 311 -2189
rect 352 -2190 353 -2189
rect 359 -2190 360 -2189
rect 548 -2190 549 -2189
rect 695 -2190 696 -2189
rect 1045 -2190 1046 -2189
rect 79 -2192 80 -2191
rect 128 -2192 129 -2191
rect 142 -2192 143 -2191
rect 149 -2192 150 -2191
rect 163 -2192 164 -2191
rect 569 -2192 570 -2191
rect 709 -2192 710 -2191
rect 779 -2192 780 -2191
rect 800 -2192 801 -2191
rect 807 -2192 808 -2191
rect 905 -2192 906 -2191
rect 1024 -2192 1025 -2191
rect 44 -2194 45 -2193
rect 128 -2194 129 -2193
rect 163 -2194 164 -2193
rect 653 -2194 654 -2193
rect 751 -2194 752 -2193
rect 870 -2194 871 -2193
rect 86 -2196 87 -2195
rect 149 -2196 150 -2195
rect 170 -2196 171 -2195
rect 233 -2196 234 -2195
rect 320 -2196 321 -2195
rect 849 -2196 850 -2195
rect 870 -2196 871 -2195
rect 1017 -2196 1018 -2195
rect 170 -2198 171 -2197
rect 177 -2198 178 -2197
rect 180 -2198 181 -2197
rect 492 -2198 493 -2197
rect 548 -2198 549 -2197
rect 590 -2198 591 -2197
rect 653 -2198 654 -2197
rect 772 -2198 773 -2197
rect 779 -2198 780 -2197
rect 821 -2198 822 -2197
rect 954 -2198 955 -2197
rect 1017 -2198 1018 -2197
rect 177 -2200 178 -2199
rect 212 -2200 213 -2199
rect 219 -2200 220 -2199
rect 345 -2200 346 -2199
rect 373 -2200 374 -2199
rect 471 -2200 472 -2199
rect 590 -2200 591 -2199
rect 625 -2200 626 -2199
rect 758 -2200 759 -2199
rect 877 -2200 878 -2199
rect 107 -2202 108 -2201
rect 345 -2202 346 -2201
rect 380 -2202 381 -2201
rect 576 -2202 577 -2201
rect 618 -2202 619 -2201
rect 625 -2202 626 -2201
rect 772 -2202 773 -2201
rect 828 -2202 829 -2201
rect 877 -2202 878 -2201
rect 947 -2202 948 -2201
rect 107 -2204 108 -2203
rect 299 -2204 300 -2203
rect 387 -2204 388 -2203
rect 436 -2204 437 -2203
rect 450 -2204 451 -2203
rect 576 -2204 577 -2203
rect 618 -2204 619 -2203
rect 793 -2204 794 -2203
rect 807 -2204 808 -2203
rect 814 -2204 815 -2203
rect 821 -2204 822 -2203
rect 891 -2204 892 -2203
rect 191 -2206 192 -2205
rect 667 -2206 668 -2205
rect 670 -2206 671 -2205
rect 891 -2206 892 -2205
rect 191 -2208 192 -2207
rect 562 -2208 563 -2207
rect 793 -2208 794 -2207
rect 835 -2208 836 -2207
rect 205 -2210 206 -2209
rect 660 -2210 661 -2209
rect 814 -2210 815 -2209
rect 912 -2210 913 -2209
rect 212 -2212 213 -2211
rect 453 -2212 454 -2211
rect 471 -2212 472 -2211
rect 520 -2212 521 -2211
rect 660 -2212 661 -2211
rect 716 -2212 717 -2211
rect 828 -2212 829 -2211
rect 940 -2212 941 -2211
rect 338 -2214 339 -2213
rect 716 -2214 717 -2213
rect 765 -2214 766 -2213
rect 940 -2214 941 -2213
rect 338 -2216 339 -2215
rect 740 -2216 741 -2215
rect 835 -2216 836 -2215
rect 926 -2216 927 -2215
rect 422 -2218 423 -2217
rect 457 -2218 458 -2217
rect 485 -2218 486 -2217
rect 947 -2218 948 -2217
rect 415 -2220 416 -2219
rect 422 -2220 423 -2219
rect 436 -2220 437 -2219
rect 723 -2220 724 -2219
rect 912 -2220 913 -2219
rect 989 -2220 990 -2219
rect 415 -2222 416 -2221
rect 527 -2222 528 -2221
rect 723 -2222 724 -2221
rect 863 -2222 864 -2221
rect 926 -2222 927 -2221
rect 1010 -2222 1011 -2221
rect 516 -2224 517 -2223
rect 562 -2224 563 -2223
rect 730 -2224 731 -2223
rect 863 -2224 864 -2223
rect 520 -2226 521 -2225
rect 534 -2226 535 -2225
rect 730 -2226 731 -2225
rect 744 -2226 745 -2225
rect 534 -2228 535 -2227
rect 600 -2228 601 -2227
rect 30 -2239 31 -2238
rect 128 -2239 129 -2238
rect 131 -2239 132 -2238
rect 338 -2239 339 -2238
rect 345 -2239 346 -2238
rect 348 -2239 349 -2238
rect 359 -2239 360 -2238
rect 656 -2239 657 -2238
rect 667 -2239 668 -2238
rect 835 -2239 836 -2238
rect 940 -2239 941 -2238
rect 961 -2239 962 -2238
rect 989 -2239 990 -2238
rect 1003 -2239 1004 -2238
rect 1017 -2239 1018 -2238
rect 1038 -2239 1039 -2238
rect 1059 -2239 1060 -2238
rect 1066 -2239 1067 -2238
rect 44 -2241 45 -2240
rect 47 -2241 48 -2240
rect 51 -2241 52 -2240
rect 89 -2241 90 -2240
rect 93 -2241 94 -2240
rect 450 -2241 451 -2240
rect 481 -2241 482 -2240
rect 632 -2241 633 -2240
rect 667 -2241 668 -2240
rect 688 -2241 689 -2240
rect 695 -2241 696 -2240
rect 751 -2241 752 -2240
rect 800 -2241 801 -2240
rect 803 -2241 804 -2240
rect 807 -2241 808 -2240
rect 810 -2241 811 -2240
rect 835 -2241 836 -2240
rect 870 -2241 871 -2240
rect 943 -2241 944 -2240
rect 982 -2241 983 -2240
rect 37 -2243 38 -2242
rect 89 -2243 90 -2242
rect 135 -2243 136 -2242
rect 338 -2243 339 -2242
rect 359 -2243 360 -2242
rect 373 -2243 374 -2242
rect 429 -2243 430 -2242
rect 478 -2243 479 -2242
rect 527 -2243 528 -2242
rect 660 -2243 661 -2242
rect 674 -2243 675 -2242
rect 677 -2243 678 -2242
rect 681 -2243 682 -2242
rect 684 -2243 685 -2242
rect 688 -2243 689 -2242
rect 765 -2243 766 -2242
rect 800 -2243 801 -2242
rect 926 -2243 927 -2242
rect 957 -2243 958 -2242
rect 975 -2243 976 -2242
rect 44 -2245 45 -2244
rect 58 -2245 59 -2244
rect 65 -2245 66 -2244
rect 128 -2245 129 -2244
rect 135 -2245 136 -2244
rect 156 -2245 157 -2244
rect 177 -2245 178 -2244
rect 240 -2245 241 -2244
rect 261 -2245 262 -2244
rect 355 -2245 356 -2244
rect 429 -2245 430 -2244
rect 506 -2245 507 -2244
rect 527 -2245 528 -2244
rect 548 -2245 549 -2244
rect 583 -2245 584 -2244
rect 586 -2245 587 -2244
rect 632 -2245 633 -2244
rect 646 -2245 647 -2244
rect 674 -2245 675 -2244
rect 758 -2245 759 -2244
rect 765 -2245 766 -2244
rect 814 -2245 815 -2244
rect 870 -2245 871 -2244
rect 954 -2245 955 -2244
rect 51 -2247 52 -2246
rect 114 -2247 115 -2246
rect 138 -2247 139 -2246
rect 565 -2247 566 -2246
rect 583 -2247 584 -2246
rect 597 -2247 598 -2246
rect 621 -2247 622 -2246
rect 646 -2247 647 -2246
rect 681 -2247 682 -2246
rect 716 -2247 717 -2246
rect 723 -2247 724 -2246
rect 758 -2247 759 -2246
rect 807 -2247 808 -2246
rect 842 -2247 843 -2246
rect 65 -2249 66 -2248
rect 100 -2249 101 -2248
rect 114 -2249 115 -2248
rect 142 -2249 143 -2248
rect 170 -2249 171 -2248
rect 177 -2249 178 -2248
rect 180 -2249 181 -2248
rect 240 -2249 241 -2248
rect 247 -2249 248 -2248
rect 261 -2249 262 -2248
rect 303 -2249 304 -2248
rect 352 -2249 353 -2248
rect 436 -2249 437 -2248
rect 453 -2249 454 -2248
rect 478 -2249 479 -2248
rect 572 -2249 573 -2248
rect 639 -2249 640 -2248
rect 660 -2249 661 -2248
rect 698 -2249 699 -2248
rect 912 -2249 913 -2248
rect 72 -2251 73 -2250
rect 530 -2251 531 -2250
rect 534 -2251 535 -2250
rect 548 -2251 549 -2250
rect 611 -2251 612 -2250
rect 639 -2251 640 -2250
rect 702 -2251 703 -2250
rect 716 -2251 717 -2250
rect 730 -2251 731 -2250
rect 744 -2251 745 -2250
rect 747 -2251 748 -2250
rect 884 -2251 885 -2250
rect 72 -2253 73 -2252
rect 163 -2253 164 -2252
rect 184 -2253 185 -2252
rect 394 -2253 395 -2252
rect 408 -2253 409 -2252
rect 436 -2253 437 -2252
rect 446 -2253 447 -2252
rect 457 -2253 458 -2252
rect 499 -2253 500 -2252
rect 506 -2253 507 -2252
rect 604 -2253 605 -2252
rect 611 -2253 612 -2252
rect 656 -2253 657 -2252
rect 884 -2253 885 -2252
rect 79 -2255 80 -2254
rect 212 -2255 213 -2254
rect 226 -2255 227 -2254
rect 653 -2255 654 -2254
rect 709 -2255 710 -2254
rect 723 -2255 724 -2254
rect 730 -2255 731 -2254
rect 772 -2255 773 -2254
rect 814 -2255 815 -2254
rect 863 -2255 864 -2254
rect 96 -2257 97 -2256
rect 226 -2257 227 -2256
rect 247 -2257 248 -2256
rect 387 -2257 388 -2256
rect 408 -2257 409 -2256
rect 541 -2257 542 -2256
rect 576 -2257 577 -2256
rect 604 -2257 605 -2256
rect 737 -2257 738 -2256
rect 751 -2257 752 -2256
rect 772 -2257 773 -2256
rect 779 -2257 780 -2256
rect 842 -2257 843 -2256
rect 891 -2257 892 -2256
rect 100 -2259 101 -2258
rect 289 -2259 290 -2258
rect 303 -2259 304 -2258
rect 376 -2259 377 -2258
rect 387 -2259 388 -2258
rect 537 -2259 538 -2258
rect 737 -2259 738 -2258
rect 786 -2259 787 -2258
rect 810 -2259 811 -2258
rect 891 -2259 892 -2258
rect 107 -2261 108 -2260
rect 142 -2261 143 -2260
rect 156 -2261 157 -2260
rect 446 -2261 447 -2260
rect 471 -2261 472 -2260
rect 499 -2261 500 -2260
rect 740 -2261 741 -2260
rect 856 -2261 857 -2260
rect 863 -2261 864 -2260
rect 947 -2261 948 -2260
rect 107 -2263 108 -2262
rect 191 -2263 192 -2262
rect 198 -2263 199 -2262
rect 292 -2263 293 -2262
rect 310 -2263 311 -2262
rect 352 -2263 353 -2262
rect 366 -2263 367 -2262
rect 394 -2263 395 -2262
rect 492 -2263 493 -2262
rect 541 -2263 542 -2262
rect 744 -2263 745 -2262
rect 793 -2263 794 -2262
rect 856 -2263 857 -2262
rect 919 -2263 920 -2262
rect 124 -2265 125 -2264
rect 170 -2265 171 -2264
rect 198 -2265 199 -2264
rect 268 -2265 269 -2264
rect 275 -2265 276 -2264
rect 453 -2265 454 -2264
rect 779 -2265 780 -2264
rect 821 -2265 822 -2264
rect 149 -2267 150 -2266
rect 191 -2267 192 -2266
rect 212 -2267 213 -2266
rect 233 -2267 234 -2266
rect 254 -2267 255 -2266
rect 534 -2267 535 -2266
rect 653 -2267 654 -2266
rect 821 -2267 822 -2266
rect 149 -2269 150 -2268
rect 187 -2269 188 -2268
rect 219 -2269 220 -2268
rect 576 -2269 577 -2268
rect 786 -2269 787 -2268
rect 828 -2269 829 -2268
rect 163 -2271 164 -2270
rect 397 -2271 398 -2270
rect 793 -2271 794 -2270
rect 905 -2271 906 -2270
rect 184 -2273 185 -2272
rect 254 -2273 255 -2272
rect 268 -2273 269 -2272
rect 485 -2273 486 -2272
rect 828 -2273 829 -2272
rect 849 -2273 850 -2272
rect 219 -2275 220 -2274
rect 373 -2275 374 -2274
rect 443 -2275 444 -2274
rect 485 -2275 486 -2274
rect 849 -2275 850 -2274
rect 898 -2275 899 -2274
rect 93 -2277 94 -2276
rect 443 -2277 444 -2276
rect 877 -2277 878 -2276
rect 898 -2277 899 -2276
rect 233 -2279 234 -2278
rect 296 -2279 297 -2278
rect 310 -2279 311 -2278
rect 380 -2279 381 -2278
rect 877 -2279 878 -2278
rect 933 -2279 934 -2278
rect 275 -2281 276 -2280
rect 282 -2281 283 -2280
rect 296 -2281 297 -2280
rect 492 -2281 493 -2280
rect 282 -2283 283 -2282
rect 317 -2283 318 -2282
rect 324 -2283 325 -2282
rect 380 -2283 381 -2282
rect 317 -2285 318 -2284
rect 579 -2285 580 -2284
rect 324 -2287 325 -2286
rect 401 -2287 402 -2286
rect 345 -2289 346 -2288
rect 457 -2289 458 -2288
rect 366 -2291 367 -2290
rect 415 -2291 416 -2290
rect 121 -2293 122 -2292
rect 415 -2293 416 -2292
rect 121 -2295 122 -2294
rect 513 -2295 514 -2294
rect 401 -2297 402 -2296
rect 555 -2297 556 -2296
rect 422 -2299 423 -2298
rect 513 -2299 514 -2298
rect 555 -2299 556 -2298
rect 569 -2299 570 -2298
rect 422 -2301 423 -2300
rect 625 -2301 626 -2300
rect 464 -2303 465 -2302
rect 569 -2303 570 -2302
rect 590 -2303 591 -2302
rect 625 -2303 626 -2302
rect 464 -2305 465 -2304
rect 670 -2305 671 -2304
rect 590 -2307 591 -2306
rect 618 -2307 619 -2306
rect 562 -2309 563 -2308
rect 618 -2309 619 -2308
rect 471 -2311 472 -2310
rect 562 -2311 563 -2310
rect 51 -2322 52 -2321
rect 184 -2322 185 -2321
rect 187 -2322 188 -2321
rect 376 -2322 377 -2321
rect 383 -2322 384 -2321
rect 471 -2322 472 -2321
rect 492 -2322 493 -2321
rect 793 -2322 794 -2321
rect 884 -2322 885 -2321
rect 940 -2322 941 -2321
rect 968 -2322 969 -2321
rect 978 -2322 979 -2321
rect 982 -2322 983 -2321
rect 989 -2322 990 -2321
rect 996 -2322 997 -2321
rect 1003 -2322 1004 -2321
rect 1038 -2322 1039 -2321
rect 1059 -2322 1060 -2321
rect 65 -2324 66 -2323
rect 86 -2324 87 -2323
rect 89 -2324 90 -2323
rect 751 -2324 752 -2323
rect 772 -2324 773 -2323
rect 800 -2324 801 -2323
rect 898 -2324 899 -2323
rect 905 -2324 906 -2323
rect 989 -2324 990 -2323
rect 1006 -2324 1007 -2323
rect 44 -2326 45 -2325
rect 86 -2326 87 -2325
rect 135 -2326 136 -2325
rect 282 -2326 283 -2325
rect 306 -2326 307 -2325
rect 471 -2326 472 -2325
rect 492 -2326 493 -2325
rect 621 -2326 622 -2325
rect 632 -2326 633 -2325
rect 656 -2326 657 -2325
rect 698 -2326 699 -2325
rect 870 -2326 871 -2325
rect 891 -2326 892 -2325
rect 898 -2326 899 -2325
rect 138 -2328 139 -2327
rect 296 -2328 297 -2327
rect 310 -2328 311 -2327
rect 450 -2328 451 -2327
rect 457 -2328 458 -2327
rect 803 -2328 804 -2327
rect 152 -2330 153 -2329
rect 261 -2330 262 -2329
rect 275 -2330 276 -2329
rect 495 -2330 496 -2329
rect 558 -2330 559 -2329
rect 828 -2330 829 -2329
rect 114 -2332 115 -2331
rect 261 -2332 262 -2331
rect 292 -2332 293 -2331
rect 296 -2332 297 -2331
rect 338 -2332 339 -2331
rect 348 -2332 349 -2331
rect 352 -2332 353 -2331
rect 443 -2332 444 -2331
rect 446 -2332 447 -2331
rect 709 -2332 710 -2331
rect 716 -2332 717 -2331
rect 719 -2332 720 -2331
rect 751 -2332 752 -2331
rect 835 -2332 836 -2331
rect 114 -2334 115 -2333
rect 184 -2334 185 -2333
rect 205 -2334 206 -2333
rect 275 -2334 276 -2333
rect 338 -2334 339 -2333
rect 366 -2334 367 -2333
rect 387 -2334 388 -2333
rect 530 -2334 531 -2333
rect 548 -2334 549 -2333
rect 709 -2334 710 -2333
rect 716 -2334 717 -2333
rect 814 -2334 815 -2333
rect 93 -2336 94 -2335
rect 205 -2336 206 -2335
rect 233 -2336 234 -2335
rect 282 -2336 283 -2335
rect 359 -2336 360 -2335
rect 373 -2336 374 -2335
rect 387 -2336 388 -2335
rect 422 -2336 423 -2335
rect 429 -2336 430 -2335
rect 534 -2336 535 -2335
rect 562 -2336 563 -2335
rect 702 -2336 703 -2335
rect 772 -2336 773 -2335
rect 863 -2336 864 -2335
rect 93 -2338 94 -2337
rect 149 -2338 150 -2337
rect 163 -2338 164 -2337
rect 352 -2338 353 -2337
rect 359 -2338 360 -2337
rect 485 -2338 486 -2337
rect 534 -2338 535 -2337
rect 625 -2338 626 -2337
rect 632 -2338 633 -2337
rect 667 -2338 668 -2337
rect 702 -2338 703 -2337
rect 821 -2338 822 -2337
rect 121 -2340 122 -2339
rect 366 -2340 367 -2339
rect 401 -2340 402 -2339
rect 443 -2340 444 -2339
rect 453 -2340 454 -2339
rect 548 -2340 549 -2339
rect 555 -2340 556 -2339
rect 562 -2340 563 -2339
rect 569 -2340 570 -2339
rect 590 -2340 591 -2339
rect 604 -2340 605 -2339
rect 607 -2340 608 -2339
rect 614 -2340 615 -2339
rect 758 -2340 759 -2339
rect 779 -2340 780 -2339
rect 814 -2340 815 -2339
rect 121 -2342 122 -2341
rect 212 -2342 213 -2341
rect 226 -2342 227 -2341
rect 401 -2342 402 -2341
rect 415 -2342 416 -2341
rect 565 -2342 566 -2341
rect 569 -2342 570 -2341
rect 611 -2342 612 -2341
rect 618 -2342 619 -2341
rect 877 -2342 878 -2341
rect 149 -2344 150 -2343
rect 310 -2344 311 -2343
rect 324 -2344 325 -2343
rect 422 -2344 423 -2343
rect 429 -2344 430 -2343
rect 464 -2344 465 -2343
rect 485 -2344 486 -2343
rect 513 -2344 514 -2343
rect 555 -2344 556 -2343
rect 618 -2344 619 -2343
rect 667 -2344 668 -2343
rect 849 -2344 850 -2343
rect 72 -2346 73 -2345
rect 513 -2346 514 -2345
rect 572 -2346 573 -2345
rect 695 -2346 696 -2345
rect 730 -2346 731 -2345
rect 779 -2346 780 -2345
rect 793 -2346 794 -2345
rect 856 -2346 857 -2345
rect 72 -2348 73 -2347
rect 317 -2348 318 -2347
rect 457 -2348 458 -2347
rect 506 -2348 507 -2347
rect 576 -2348 577 -2347
rect 660 -2348 661 -2347
rect 730 -2348 731 -2347
rect 737 -2348 738 -2347
rect 758 -2348 759 -2347
rect 765 -2348 766 -2347
rect 107 -2350 108 -2349
rect 324 -2350 325 -2349
rect 464 -2350 465 -2349
rect 527 -2350 528 -2349
rect 576 -2350 577 -2349
rect 583 -2350 584 -2349
rect 590 -2350 591 -2349
rect 597 -2350 598 -2349
rect 604 -2350 605 -2349
rect 646 -2350 647 -2349
rect 660 -2350 661 -2349
rect 674 -2350 675 -2349
rect 765 -2350 766 -2349
rect 842 -2350 843 -2349
rect 107 -2352 108 -2351
rect 380 -2352 381 -2351
rect 478 -2352 479 -2351
rect 506 -2352 507 -2351
rect 583 -2352 584 -2351
rect 688 -2352 689 -2351
rect 719 -2352 720 -2351
rect 737 -2352 738 -2351
rect 156 -2354 157 -2353
rect 212 -2354 213 -2353
rect 226 -2354 227 -2353
rect 233 -2354 234 -2353
rect 236 -2354 237 -2353
rect 695 -2354 696 -2353
rect 128 -2356 129 -2355
rect 156 -2356 157 -2355
rect 247 -2356 248 -2355
rect 425 -2356 426 -2355
rect 478 -2356 479 -2355
rect 541 -2356 542 -2355
rect 597 -2356 598 -2355
rect 639 -2356 640 -2355
rect 674 -2356 675 -2355
rect 786 -2356 787 -2355
rect 128 -2358 129 -2357
rect 219 -2358 220 -2357
rect 254 -2358 255 -2357
rect 373 -2358 374 -2357
rect 499 -2358 500 -2357
rect 611 -2358 612 -2357
rect 639 -2358 640 -2357
rect 681 -2358 682 -2357
rect 191 -2360 192 -2359
rect 247 -2360 248 -2359
rect 254 -2360 255 -2359
rect 450 -2360 451 -2359
rect 527 -2360 528 -2359
rect 688 -2360 689 -2359
rect 170 -2362 171 -2361
rect 191 -2362 192 -2361
rect 219 -2362 220 -2361
rect 268 -2362 269 -2361
rect 271 -2362 272 -2361
rect 415 -2362 416 -2361
rect 681 -2362 682 -2361
rect 744 -2362 745 -2361
rect 142 -2364 143 -2363
rect 170 -2364 171 -2363
rect 289 -2364 290 -2363
rect 541 -2364 542 -2363
rect 723 -2364 724 -2363
rect 744 -2364 745 -2363
rect 100 -2366 101 -2365
rect 289 -2366 290 -2365
rect 303 -2366 304 -2365
rect 625 -2366 626 -2365
rect 79 -2368 80 -2367
rect 303 -2368 304 -2367
rect 317 -2368 318 -2367
rect 345 -2368 346 -2367
rect 408 -2368 409 -2367
rect 499 -2368 500 -2367
rect 58 -2370 59 -2369
rect 79 -2370 80 -2369
rect 100 -2370 101 -2369
rect 163 -2370 164 -2369
rect 331 -2370 332 -2369
rect 345 -2370 346 -2369
rect 408 -2370 409 -2369
rect 653 -2370 654 -2369
rect 142 -2372 143 -2371
rect 516 -2372 517 -2371
rect 653 -2372 654 -2371
rect 807 -2372 808 -2371
rect 198 -2374 199 -2373
rect 331 -2374 332 -2373
rect 177 -2376 178 -2375
rect 198 -2376 199 -2375
rect 72 -2387 73 -2386
rect 163 -2387 164 -2386
rect 166 -2387 167 -2386
rect 198 -2387 199 -2386
rect 303 -2387 304 -2386
rect 345 -2387 346 -2386
rect 355 -2387 356 -2386
rect 541 -2387 542 -2386
rect 646 -2387 647 -2386
rect 684 -2387 685 -2386
rect 723 -2387 724 -2386
rect 730 -2387 731 -2386
rect 800 -2387 801 -2386
rect 807 -2387 808 -2386
rect 814 -2387 815 -2386
rect 828 -2387 829 -2386
rect 891 -2387 892 -2386
rect 905 -2387 906 -2386
rect 940 -2387 941 -2386
rect 1006 -2387 1007 -2386
rect 79 -2389 80 -2388
rect 187 -2389 188 -2388
rect 191 -2389 192 -2388
rect 236 -2389 237 -2388
rect 303 -2389 304 -2388
rect 401 -2389 402 -2388
rect 418 -2389 419 -2388
rect 698 -2389 699 -2388
rect 730 -2389 731 -2388
rect 744 -2389 745 -2388
rect 779 -2389 780 -2388
rect 800 -2389 801 -2388
rect 975 -2389 976 -2388
rect 989 -2389 990 -2388
rect 86 -2391 87 -2390
rect 149 -2391 150 -2390
rect 156 -2391 157 -2390
rect 173 -2391 174 -2390
rect 177 -2391 178 -2390
rect 247 -2391 248 -2390
rect 282 -2391 283 -2390
rect 401 -2391 402 -2390
rect 422 -2391 423 -2390
rect 614 -2391 615 -2390
rect 688 -2391 689 -2390
rect 744 -2391 745 -2390
rect 978 -2391 979 -2390
rect 982 -2391 983 -2390
rect 93 -2393 94 -2392
rect 184 -2393 185 -2392
rect 219 -2393 220 -2392
rect 422 -2393 423 -2392
rect 429 -2393 430 -2392
rect 488 -2393 489 -2392
rect 499 -2393 500 -2392
rect 527 -2393 528 -2392
rect 530 -2393 531 -2392
rect 625 -2393 626 -2392
rect 691 -2393 692 -2392
rect 905 -2393 906 -2392
rect 121 -2395 122 -2394
rect 268 -2395 269 -2394
rect 310 -2395 311 -2394
rect 383 -2395 384 -2394
rect 394 -2395 395 -2394
rect 509 -2395 510 -2394
rect 516 -2395 517 -2394
rect 702 -2395 703 -2394
rect 135 -2397 136 -2396
rect 450 -2397 451 -2396
rect 453 -2397 454 -2396
rect 653 -2397 654 -2396
rect 142 -2399 143 -2398
rect 198 -2399 199 -2398
rect 205 -2399 206 -2398
rect 219 -2399 220 -2398
rect 247 -2399 248 -2398
rect 261 -2399 262 -2398
rect 268 -2399 269 -2398
rect 306 -2399 307 -2398
rect 310 -2399 311 -2398
rect 408 -2399 409 -2398
rect 443 -2399 444 -2398
rect 558 -2399 559 -2398
rect 576 -2399 577 -2398
rect 625 -2399 626 -2398
rect 653 -2399 654 -2398
rect 674 -2399 675 -2398
rect 261 -2401 262 -2400
rect 324 -2401 325 -2400
rect 345 -2401 346 -2400
rect 383 -2401 384 -2400
rect 436 -2401 437 -2400
rect 443 -2401 444 -2400
rect 450 -2401 451 -2400
rect 464 -2401 465 -2400
rect 499 -2401 500 -2400
rect 506 -2401 507 -2400
rect 516 -2401 517 -2400
rect 583 -2401 584 -2400
rect 674 -2401 675 -2400
rect 716 -2401 717 -2400
rect 254 -2403 255 -2402
rect 324 -2403 325 -2402
rect 352 -2403 353 -2402
rect 541 -2403 542 -2402
rect 548 -2403 549 -2402
rect 646 -2403 647 -2402
rect 716 -2403 717 -2402
rect 751 -2403 752 -2402
rect 128 -2405 129 -2404
rect 254 -2405 255 -2404
rect 296 -2405 297 -2404
rect 394 -2405 395 -2404
rect 415 -2405 416 -2404
rect 464 -2405 465 -2404
rect 492 -2405 493 -2404
rect 506 -2405 507 -2404
rect 513 -2405 514 -2404
rect 583 -2405 584 -2404
rect 709 -2405 710 -2404
rect 751 -2405 752 -2404
rect 212 -2407 213 -2406
rect 296 -2407 297 -2406
rect 359 -2407 360 -2406
rect 408 -2407 409 -2406
rect 436 -2407 437 -2406
rect 457 -2407 458 -2406
rect 460 -2407 461 -2406
rect 485 -2407 486 -2406
rect 492 -2407 493 -2406
rect 534 -2407 535 -2406
rect 548 -2407 549 -2406
rect 555 -2407 556 -2406
rect 576 -2407 577 -2406
rect 597 -2407 598 -2406
rect 289 -2409 290 -2408
rect 359 -2409 360 -2408
rect 366 -2409 367 -2408
rect 611 -2409 612 -2408
rect 100 -2411 101 -2410
rect 289 -2411 290 -2410
rect 369 -2411 370 -2410
rect 387 -2411 388 -2410
rect 478 -2411 479 -2410
rect 534 -2411 535 -2410
rect 555 -2411 556 -2410
rect 688 -2411 689 -2410
rect 114 -2413 115 -2412
rect 387 -2413 388 -2412
rect 523 -2413 524 -2412
rect 569 -2413 570 -2412
rect 597 -2413 598 -2412
rect 604 -2413 605 -2412
rect 611 -2413 612 -2412
rect 632 -2413 633 -2412
rect 331 -2415 332 -2414
rect 478 -2415 479 -2414
rect 604 -2415 605 -2414
rect 667 -2415 668 -2414
rect 233 -2417 234 -2416
rect 331 -2417 332 -2416
rect 373 -2417 374 -2416
rect 513 -2417 514 -2416
rect 632 -2417 633 -2416
rect 660 -2417 661 -2416
rect 667 -2417 668 -2416
rect 681 -2417 682 -2416
rect 226 -2419 227 -2418
rect 233 -2419 234 -2418
rect 338 -2419 339 -2418
rect 373 -2419 374 -2418
rect 471 -2419 472 -2418
rect 569 -2419 570 -2418
rect 618 -2419 619 -2418
rect 660 -2419 661 -2418
rect 681 -2419 682 -2418
rect 765 -2419 766 -2418
rect 107 -2421 108 -2420
rect 226 -2421 227 -2420
rect 317 -2421 318 -2420
rect 338 -2421 339 -2420
rect 471 -2421 472 -2420
rect 562 -2421 563 -2420
rect 618 -2421 619 -2420
rect 639 -2421 640 -2420
rect 758 -2421 759 -2420
rect 765 -2421 766 -2420
rect 275 -2423 276 -2422
rect 317 -2423 318 -2422
rect 562 -2423 563 -2422
rect 590 -2423 591 -2422
rect 737 -2423 738 -2422
rect 758 -2423 759 -2422
rect 275 -2425 276 -2424
rect 380 -2425 381 -2424
rect 520 -2425 521 -2424
rect 590 -2425 591 -2424
rect 737 -2425 738 -2424
rect 772 -2425 773 -2424
rect 282 -2427 283 -2426
rect 380 -2427 381 -2426
rect 429 -2427 430 -2426
rect 520 -2427 521 -2426
rect 772 -2427 773 -2426
rect 793 -2427 794 -2426
rect 226 -2438 227 -2437
rect 352 -2438 353 -2437
rect 380 -2438 381 -2437
rect 471 -2438 472 -2437
rect 509 -2438 510 -2437
rect 576 -2438 577 -2437
rect 607 -2438 608 -2437
rect 618 -2438 619 -2437
rect 639 -2438 640 -2437
rect 691 -2438 692 -2437
rect 702 -2438 703 -2437
rect 716 -2438 717 -2437
rect 744 -2438 745 -2437
rect 758 -2438 759 -2437
rect 807 -2438 808 -2437
rect 817 -2438 818 -2437
rect 898 -2438 899 -2437
rect 905 -2438 906 -2437
rect 219 -2440 220 -2439
rect 226 -2440 227 -2439
rect 233 -2440 234 -2439
rect 243 -2440 244 -2439
rect 261 -2440 262 -2439
rect 366 -2440 367 -2439
rect 387 -2440 388 -2439
rect 513 -2440 514 -2439
rect 569 -2440 570 -2439
rect 611 -2440 612 -2439
rect 614 -2440 615 -2439
rect 908 -2440 909 -2439
rect 233 -2442 234 -2441
rect 247 -2442 248 -2441
rect 275 -2442 276 -2441
rect 369 -2442 370 -2441
rect 387 -2442 388 -2441
rect 429 -2442 430 -2441
rect 432 -2442 433 -2441
rect 562 -2442 563 -2441
rect 572 -2442 573 -2441
rect 597 -2442 598 -2441
rect 611 -2442 612 -2441
rect 653 -2442 654 -2441
rect 660 -2442 661 -2441
rect 663 -2442 664 -2441
rect 688 -2442 689 -2441
rect 737 -2442 738 -2441
rect 747 -2442 748 -2441
rect 765 -2442 766 -2441
rect 800 -2442 801 -2441
rect 807 -2442 808 -2441
rect 891 -2442 892 -2441
rect 898 -2442 899 -2441
rect 236 -2444 237 -2443
rect 327 -2444 328 -2443
rect 331 -2444 332 -2443
rect 457 -2444 458 -2443
rect 460 -2444 461 -2443
rect 838 -2444 839 -2443
rect 282 -2446 283 -2445
rect 418 -2446 419 -2445
rect 450 -2446 451 -2445
rect 506 -2446 507 -2445
rect 509 -2446 510 -2445
rect 583 -2446 584 -2445
rect 590 -2446 591 -2445
rect 618 -2446 619 -2445
rect 625 -2446 626 -2445
rect 653 -2446 654 -2445
rect 660 -2446 661 -2445
rect 674 -2446 675 -2445
rect 730 -2446 731 -2445
rect 744 -2446 745 -2445
rect 751 -2446 752 -2445
rect 754 -2446 755 -2445
rect 296 -2448 297 -2447
rect 331 -2448 332 -2447
rect 338 -2448 339 -2447
rect 366 -2448 367 -2447
rect 401 -2448 402 -2447
rect 453 -2448 454 -2447
rect 457 -2448 458 -2447
rect 523 -2448 524 -2447
rect 576 -2448 577 -2447
rect 604 -2448 605 -2447
rect 625 -2448 626 -2447
rect 649 -2448 650 -2447
rect 663 -2448 664 -2447
rect 674 -2448 675 -2447
rect 751 -2448 752 -2447
rect 772 -2448 773 -2447
rect 254 -2450 255 -2449
rect 296 -2450 297 -2449
rect 310 -2450 311 -2449
rect 352 -2450 353 -2449
rect 373 -2450 374 -2449
rect 401 -2450 402 -2449
rect 453 -2450 454 -2449
rect 499 -2450 500 -2449
rect 597 -2450 598 -2449
rect 632 -2450 633 -2449
rect 646 -2450 647 -2449
rect 688 -2450 689 -2449
rect 198 -2452 199 -2451
rect 254 -2452 255 -2451
rect 268 -2452 269 -2451
rect 310 -2452 311 -2451
rect 317 -2452 318 -2451
rect 450 -2452 451 -2451
rect 464 -2452 465 -2451
rect 471 -2452 472 -2451
rect 499 -2452 500 -2451
rect 534 -2452 535 -2451
rect 541 -2452 542 -2451
rect 632 -2452 633 -2451
rect 646 -2452 647 -2451
rect 667 -2452 668 -2451
rect 341 -2454 342 -2453
rect 548 -2454 549 -2453
rect 345 -2456 346 -2455
rect 373 -2456 374 -2455
rect 443 -2456 444 -2455
rect 464 -2456 465 -2455
rect 478 -2456 479 -2455
rect 548 -2456 549 -2455
rect 303 -2458 304 -2457
rect 345 -2458 346 -2457
rect 348 -2458 349 -2457
rect 555 -2458 556 -2457
rect 394 -2460 395 -2459
rect 443 -2460 444 -2459
rect 478 -2460 479 -2459
rect 485 -2460 486 -2459
rect 527 -2460 528 -2459
rect 541 -2460 542 -2459
rect 359 -2462 360 -2461
rect 394 -2462 395 -2461
rect 422 -2462 423 -2461
rect 485 -2462 486 -2461
rect 492 -2462 493 -2461
rect 527 -2462 528 -2461
rect 289 -2464 290 -2463
rect 359 -2464 360 -2463
rect 415 -2464 416 -2463
rect 492 -2464 493 -2463
rect 422 -2466 423 -2465
rect 436 -2466 437 -2465
rect 436 -2468 437 -2467
rect 516 -2468 517 -2467
rect 247 -2479 248 -2478
rect 254 -2479 255 -2478
rect 296 -2479 297 -2478
rect 341 -2479 342 -2478
rect 359 -2479 360 -2478
rect 380 -2479 381 -2478
rect 390 -2479 391 -2478
rect 457 -2479 458 -2478
rect 492 -2479 493 -2478
rect 509 -2479 510 -2478
rect 513 -2479 514 -2478
rect 611 -2479 612 -2478
rect 649 -2479 650 -2478
rect 653 -2479 654 -2478
rect 674 -2479 675 -2478
rect 691 -2479 692 -2478
rect 726 -2479 727 -2478
rect 901 -2479 902 -2478
rect 310 -2481 311 -2480
rect 348 -2481 349 -2480
rect 359 -2481 360 -2480
rect 387 -2481 388 -2480
rect 394 -2481 395 -2480
rect 429 -2481 430 -2480
rect 432 -2481 433 -2480
rect 499 -2481 500 -2480
rect 527 -2481 528 -2480
rect 534 -2481 535 -2480
rect 541 -2481 542 -2480
rect 555 -2481 556 -2480
rect 604 -2481 605 -2480
rect 639 -2481 640 -2480
rect 653 -2481 654 -2480
rect 660 -2481 661 -2480
rect 688 -2481 689 -2480
rect 695 -2481 696 -2480
rect 744 -2481 745 -2480
rect 751 -2481 752 -2480
rect 807 -2481 808 -2480
rect 817 -2481 818 -2480
rect 828 -2481 829 -2480
rect 835 -2481 836 -2480
rect 898 -2481 899 -2480
rect 905 -2481 906 -2480
rect 331 -2483 332 -2482
rect 369 -2483 370 -2482
rect 373 -2483 374 -2482
rect 394 -2483 395 -2482
rect 401 -2483 402 -2482
rect 408 -2483 409 -2482
rect 443 -2483 444 -2482
rect 471 -2483 472 -2482
rect 548 -2483 549 -2482
rect 614 -2483 615 -2482
rect 632 -2483 633 -2482
rect 660 -2483 661 -2482
rect 688 -2483 689 -2482
rect 702 -2483 703 -2482
rect 352 -2485 353 -2484
rect 373 -2485 374 -2484
rect 404 -2485 405 -2484
rect 422 -2485 423 -2484
rect 446 -2485 447 -2484
rect 464 -2485 465 -2484
rect 485 -2485 486 -2484
rect 548 -2485 549 -2484
rect 551 -2485 552 -2484
rect 576 -2485 577 -2484
rect 597 -2485 598 -2484
rect 604 -2485 605 -2484
rect 614 -2485 615 -2484
rect 625 -2485 626 -2484
rect 695 -2485 696 -2484
rect 702 -2485 703 -2484
rect 366 -2487 367 -2486
rect 387 -2487 388 -2486
rect 453 -2487 454 -2486
rect 478 -2487 479 -2486
rect 618 -2487 619 -2486
rect 632 -2487 633 -2486
rect 366 -2489 367 -2488
rect 436 -2489 437 -2488
rect 226 -2500 227 -2499
rect 233 -2500 234 -2499
rect 236 -2500 237 -2499
rect 240 -2500 241 -2499
rect 359 -2500 360 -2499
rect 366 -2500 367 -2499
rect 373 -2500 374 -2499
rect 394 -2500 395 -2499
rect 397 -2500 398 -2499
rect 408 -2500 409 -2499
rect 534 -2500 535 -2499
rect 548 -2500 549 -2499
rect 558 -2500 559 -2499
rect 901 -2500 902 -2499
rect 380 -2502 381 -2501
rect 401 -2502 402 -2501
rect 604 -2502 605 -2501
rect 611 -2502 612 -2501
rect 632 -2502 633 -2501
rect 653 -2502 654 -2501
rect 660 -2502 661 -2501
rect 691 -2502 692 -2501
rect 702 -2502 703 -2501
rect 726 -2502 727 -2501
rect 898 -2502 899 -2501
rect 905 -2502 906 -2501
<< metal2 >>
rect 152 -5 153 1
rect 205 -5 206 1
rect 338 -5 339 1
rect 352 -5 353 1
rect 366 -5 367 1
rect 411 -5 412 1
rect 432 -5 433 1
rect 513 -5 514 1
rect 341 -5 342 -1
rect 359 -5 360 -1
rect 394 -5 395 -1
rect 471 -5 472 -1
rect 492 -5 493 -1
rect 576 -5 577 -1
rect 345 -5 346 -3
rect 376 -5 377 -3
rect 408 -5 409 -3
rect 450 -5 451 -3
rect 464 -5 465 -3
rect 481 -5 482 -3
rect 128 -36 129 -14
rect 149 -15 150 -13
rect 198 -36 199 -14
rect 289 -36 290 -14
rect 292 -36 293 -14
rect 310 -36 311 -14
rect 320 -36 321 -14
rect 457 -36 458 -14
rect 464 -15 465 -13
rect 485 -36 486 -14
rect 502 -36 503 -14
rect 548 -36 549 -14
rect 576 -15 577 -13
rect 625 -36 626 -14
rect 208 -17 209 -13
rect 219 -36 220 -16
rect 243 -36 244 -16
rect 254 -36 255 -16
rect 282 -36 283 -16
rect 341 -17 342 -13
rect 352 -17 353 -13
rect 380 -36 381 -16
rect 415 -36 416 -16
rect 492 -17 493 -13
rect 513 -17 514 -13
rect 541 -36 542 -16
rect 593 -36 594 -16
rect 618 -36 619 -16
rect 296 -36 297 -18
rect 446 -36 447 -18
rect 450 -19 451 -13
rect 471 -36 472 -18
rect 474 -19 475 -13
rect 527 -36 528 -18
rect 303 -36 304 -20
rect 432 -21 433 -13
rect 450 -36 451 -20
rect 478 -21 479 -13
rect 324 -36 325 -22
rect 345 -23 346 -13
rect 352 -36 353 -22
rect 432 -36 433 -22
rect 436 -23 437 -13
rect 478 -36 479 -22
rect 327 -36 328 -24
rect 408 -36 409 -24
rect 429 -25 430 -13
rect 513 -36 514 -24
rect 331 -36 332 -26
rect 366 -27 367 -13
rect 376 -36 377 -26
rect 387 -36 388 -26
rect 401 -27 402 -13
rect 436 -36 437 -26
rect 464 -36 465 -26
rect 534 -36 535 -26
rect 338 -36 339 -28
rect 394 -29 395 -13
rect 401 -36 402 -28
rect 439 -29 440 -13
rect 345 -36 346 -30
rect 404 -31 405 -13
rect 359 -33 360 -13
rect 359 -36 360 -32
rect 359 -33 360 -13
rect 359 -36 360 -32
rect 366 -36 367 -32
rect 373 -33 374 -13
rect 394 -36 395 -32
rect 422 -36 423 -32
rect 373 -36 374 -34
rect 506 -36 507 -34
rect 114 -89 115 -45
rect 128 -46 129 -44
rect 142 -89 143 -45
rect 198 -46 199 -44
rect 205 -89 206 -45
rect 219 -46 220 -44
rect 233 -89 234 -45
rect 243 -46 244 -44
rect 247 -89 248 -45
rect 390 -89 391 -45
rect 415 -46 416 -44
rect 429 -89 430 -45
rect 432 -46 433 -44
rect 569 -89 570 -45
rect 593 -46 594 -44
rect 681 -89 682 -45
rect 170 -89 171 -47
rect 240 -48 241 -44
rect 254 -48 255 -44
rect 275 -89 276 -47
rect 317 -89 318 -47
rect 387 -48 388 -44
rect 443 -48 444 -44
rect 555 -89 556 -47
rect 593 -89 594 -47
rect 597 -89 598 -47
rect 618 -48 619 -44
rect 646 -89 647 -47
rect 653 -89 654 -47
rect 691 -89 692 -47
rect 191 -89 192 -49
rect 296 -50 297 -44
rect 331 -50 332 -44
rect 415 -89 416 -49
rect 443 -89 444 -49
rect 492 -50 493 -44
rect 495 -50 496 -44
rect 618 -89 619 -49
rect 625 -50 626 -44
rect 660 -89 661 -49
rect 674 -89 675 -49
rect 688 -89 689 -49
rect 198 -89 199 -51
rect 334 -89 335 -51
rect 338 -52 339 -44
rect 373 -52 374 -44
rect 394 -52 395 -44
rect 492 -89 493 -51
rect 502 -52 503 -44
rect 583 -89 584 -51
rect 212 -89 213 -53
rect 303 -54 304 -44
rect 338 -89 339 -53
rect 380 -54 381 -44
rect 478 -54 479 -44
rect 639 -89 640 -53
rect 219 -89 220 -55
rect 310 -56 311 -44
rect 359 -56 360 -44
rect 359 -89 360 -55
rect 359 -56 360 -44
rect 359 -89 360 -55
rect 369 -89 370 -55
rect 520 -89 521 -55
rect 527 -56 528 -44
rect 530 -74 531 -55
rect 534 -56 535 -44
rect 667 -89 668 -55
rect 240 -89 241 -57
rect 324 -58 325 -44
rect 380 -89 381 -57
rect 576 -89 577 -57
rect 254 -89 255 -59
rect 450 -60 451 -44
rect 478 -89 479 -59
rect 625 -89 626 -59
rect 177 -89 178 -61
rect 450 -89 451 -61
rect 485 -62 486 -44
rect 562 -89 563 -61
rect 261 -89 262 -63
rect 366 -64 367 -44
rect 408 -64 409 -44
rect 485 -89 486 -63
rect 499 -64 500 -44
rect 534 -89 535 -63
rect 541 -64 542 -44
rect 541 -89 542 -63
rect 541 -64 542 -44
rect 541 -89 542 -63
rect 548 -64 549 -44
rect 632 -89 633 -63
rect 226 -89 227 -65
rect 366 -89 367 -65
rect 387 -89 388 -65
rect 548 -89 549 -65
rect 268 -89 269 -67
rect 320 -68 321 -44
rect 408 -89 409 -67
rect 457 -68 458 -44
rect 506 -68 507 -44
rect 604 -89 605 -67
rect 282 -70 283 -44
rect 310 -89 311 -69
rect 436 -70 437 -44
rect 457 -89 458 -69
rect 474 -89 475 -69
rect 506 -89 507 -69
rect 513 -70 514 -44
rect 611 -89 612 -69
rect 282 -89 283 -71
rect 345 -72 346 -44
rect 422 -72 423 -44
rect 436 -89 437 -71
rect 446 -72 447 -44
rect 499 -89 500 -71
rect 527 -89 528 -71
rect 590 -72 591 -44
rect 163 -89 164 -73
rect 345 -89 346 -73
rect 422 -89 423 -73
rect 471 -74 472 -44
rect 590 -89 591 -73
rect 289 -76 290 -44
rect 324 -89 325 -75
rect 464 -76 465 -44
rect 513 -89 514 -75
rect 289 -89 290 -77
rect 401 -78 402 -44
rect 296 -89 297 -79
rect 397 -80 398 -44
rect 184 -89 185 -81
rect 397 -89 398 -81
rect 303 -89 304 -83
rect 352 -84 353 -44
rect 373 -89 374 -83
rect 401 -89 402 -83
rect 348 -89 349 -85
rect 464 -89 465 -85
rect 352 -89 353 -87
rect 481 -89 482 -87
rect 51 -156 52 -98
rect 411 -156 412 -98
rect 464 -99 465 -97
rect 723 -156 724 -98
rect 58 -156 59 -100
rect 453 -101 454 -97
rect 471 -101 472 -97
rect 814 -156 815 -100
rect 65 -156 66 -102
rect 142 -103 143 -97
rect 145 -156 146 -102
rect 184 -103 185 -97
rect 198 -103 199 -97
rect 208 -145 209 -102
rect 275 -103 276 -97
rect 376 -103 377 -97
rect 394 -103 395 -97
rect 772 -156 773 -102
rect 72 -156 73 -104
rect 82 -156 83 -104
rect 86 -156 87 -104
rect 117 -105 118 -97
rect 121 -156 122 -104
rect 194 -156 195 -104
rect 198 -156 199 -104
rect 268 -105 269 -97
rect 275 -156 276 -104
rect 474 -105 475 -97
rect 485 -105 486 -97
rect 807 -156 808 -104
rect 93 -156 94 -106
rect 296 -107 297 -97
rect 331 -107 332 -97
rect 383 -107 384 -97
rect 485 -156 486 -106
rect 611 -107 612 -97
rect 632 -107 633 -97
rect 779 -156 780 -106
rect 107 -156 108 -108
rect 247 -109 248 -97
rect 268 -156 269 -108
rect 338 -109 339 -97
rect 345 -109 346 -97
rect 429 -109 430 -97
rect 492 -109 493 -97
rect 695 -156 696 -108
rect 114 -111 115 -97
rect 135 -156 136 -110
rect 156 -156 157 -110
rect 289 -111 290 -97
rect 359 -111 360 -97
rect 394 -156 395 -110
rect 418 -156 419 -110
rect 611 -156 612 -110
rect 639 -111 640 -97
rect 786 -156 787 -110
rect 114 -156 115 -112
rect 278 -113 279 -97
rect 324 -113 325 -97
rect 359 -156 360 -112
rect 366 -156 367 -112
rect 387 -113 388 -97
rect 450 -113 451 -97
rect 639 -156 640 -112
rect 653 -113 654 -97
rect 737 -156 738 -112
rect 128 -156 129 -114
rect 254 -115 255 -97
rect 261 -115 262 -97
rect 289 -156 290 -114
rect 310 -115 311 -97
rect 324 -156 325 -114
rect 369 -115 370 -97
rect 429 -156 430 -114
rect 495 -156 496 -114
rect 709 -156 710 -114
rect 152 -156 153 -116
rect 261 -156 262 -116
rect 303 -117 304 -97
rect 310 -156 311 -116
rect 387 -156 388 -116
rect 401 -117 402 -97
rect 520 -117 521 -97
rect 653 -156 654 -116
rect 660 -117 661 -97
rect 716 -156 717 -116
rect 170 -119 171 -97
rect 296 -156 297 -118
rect 303 -156 304 -118
rect 464 -156 465 -118
rect 478 -156 479 -118
rect 660 -156 661 -118
rect 667 -119 668 -97
rect 751 -156 752 -118
rect 170 -156 171 -120
rect 226 -121 227 -97
rect 247 -156 248 -120
rect 380 -121 381 -97
rect 534 -121 535 -97
rect 765 -156 766 -120
rect 100 -156 101 -122
rect 226 -156 227 -122
rect 254 -156 255 -122
rect 471 -156 472 -122
rect 534 -156 535 -122
rect 579 -156 580 -122
rect 583 -123 584 -97
rect 632 -156 633 -122
rect 646 -123 647 -97
rect 667 -156 668 -122
rect 674 -123 675 -97
rect 730 -156 731 -122
rect 184 -156 185 -124
rect 187 -156 188 -124
rect 201 -156 202 -124
rect 331 -156 332 -124
rect 380 -156 381 -124
rect 474 -156 475 -124
rect 499 -125 500 -97
rect 646 -156 647 -124
rect 681 -125 682 -97
rect 821 -156 822 -124
rect 219 -127 220 -97
rect 338 -156 339 -126
rect 436 -127 437 -97
rect 499 -156 500 -126
rect 513 -127 514 -97
rect 681 -156 682 -126
rect 688 -127 689 -97
rect 793 -156 794 -126
rect 191 -129 192 -97
rect 436 -156 437 -128
rect 467 -156 468 -128
rect 583 -156 584 -128
rect 590 -156 591 -128
rect 618 -129 619 -97
rect 625 -129 626 -97
rect 688 -156 689 -128
rect 219 -156 220 -130
rect 240 -131 241 -97
rect 317 -131 318 -97
rect 401 -156 402 -130
rect 453 -156 454 -130
rect 618 -156 619 -130
rect 205 -133 206 -97
rect 240 -156 241 -132
rect 282 -133 283 -97
rect 317 -156 318 -132
rect 481 -133 482 -97
rect 513 -156 514 -132
rect 527 -133 528 -97
rect 674 -156 675 -132
rect 177 -135 178 -97
rect 282 -156 283 -134
rect 506 -135 507 -97
rect 527 -156 528 -134
rect 548 -135 549 -97
rect 744 -156 745 -134
rect 177 -156 178 -136
rect 212 -137 213 -97
rect 373 -137 374 -97
rect 548 -156 549 -136
rect 562 -137 563 -97
rect 800 -156 801 -136
rect 163 -139 164 -97
rect 212 -156 213 -138
rect 334 -139 335 -97
rect 562 -156 563 -138
rect 569 -139 570 -97
rect 758 -156 759 -138
rect 163 -156 164 -140
rect 352 -141 353 -97
rect 373 -156 374 -140
rect 597 -141 598 -97
rect 205 -156 206 -142
rect 233 -143 234 -97
rect 352 -156 353 -142
rect 625 -156 626 -142
rect 233 -156 234 -144
rect 415 -145 416 -97
rect 506 -156 507 -144
rect 541 -145 542 -97
rect 569 -156 570 -144
rect 576 -145 577 -97
rect 702 -156 703 -144
rect 345 -156 346 -146
rect 415 -156 416 -146
rect 422 -147 423 -97
rect 541 -156 542 -146
rect 555 -147 556 -97
rect 597 -156 598 -146
rect 422 -156 423 -148
rect 457 -149 458 -97
rect 520 -156 521 -148
rect 576 -156 577 -148
rect 443 -151 444 -97
rect 555 -156 556 -150
rect 408 -153 409 -97
rect 443 -156 444 -152
rect 457 -156 458 -152
rect 604 -153 605 -97
rect 593 -155 594 -97
rect 604 -156 605 -154
rect 44 -237 45 -165
rect 184 -166 185 -164
rect 191 -166 192 -164
rect 212 -166 213 -164
rect 240 -166 241 -164
rect 240 -237 241 -165
rect 240 -166 241 -164
rect 240 -237 241 -165
rect 268 -166 269 -164
rect 352 -166 353 -164
rect 362 -237 363 -165
rect 765 -166 766 -164
rect 793 -166 794 -164
rect 849 -237 850 -165
rect 65 -168 66 -164
rect 166 -237 167 -167
rect 184 -237 185 -167
rect 310 -168 311 -164
rect 348 -237 349 -167
rect 695 -168 696 -164
rect 751 -168 752 -164
rect 793 -237 794 -167
rect 800 -168 801 -164
rect 863 -237 864 -167
rect 65 -237 66 -169
rect 72 -170 73 -164
rect 79 -237 80 -169
rect 86 -170 87 -164
rect 100 -170 101 -164
rect 257 -237 258 -169
rect 310 -237 311 -169
rect 324 -170 325 -164
rect 352 -237 353 -169
rect 453 -170 454 -164
rect 464 -170 465 -164
rect 807 -170 808 -164
rect 814 -170 815 -164
rect 835 -237 836 -169
rect 72 -237 73 -171
rect 359 -172 360 -164
rect 408 -172 409 -164
rect 786 -172 787 -164
rect 821 -172 822 -164
rect 842 -237 843 -171
rect 86 -237 87 -173
rect 194 -174 195 -164
rect 198 -237 199 -173
rect 233 -174 234 -164
rect 324 -237 325 -173
rect 422 -174 423 -164
rect 471 -237 472 -173
rect 807 -237 808 -173
rect 103 -176 104 -164
rect 355 -237 356 -175
rect 411 -176 412 -164
rect 723 -176 724 -164
rect 730 -176 731 -164
rect 786 -237 787 -175
rect 117 -237 118 -177
rect 765 -237 766 -177
rect 772 -178 773 -164
rect 814 -237 815 -177
rect 121 -180 122 -164
rect 201 -180 202 -164
rect 212 -237 213 -179
rect 275 -180 276 -164
rect 285 -237 286 -179
rect 422 -237 423 -179
rect 492 -180 493 -164
rect 548 -180 549 -164
rect 576 -180 577 -164
rect 828 -237 829 -179
rect 121 -237 122 -181
rect 124 -237 125 -181
rect 128 -182 129 -164
rect 464 -237 465 -181
rect 495 -182 496 -164
rect 744 -182 745 -164
rect 779 -182 780 -164
rect 821 -237 822 -181
rect 128 -237 129 -183
rect 226 -184 227 -164
rect 275 -237 276 -183
rect 317 -184 318 -164
rect 415 -184 416 -164
rect 758 -184 759 -164
rect 138 -237 139 -185
rect 425 -237 426 -185
rect 460 -237 461 -185
rect 758 -237 759 -185
rect 145 -188 146 -164
rect 366 -188 367 -164
rect 415 -237 416 -187
rect 478 -188 479 -164
rect 495 -237 496 -187
rect 737 -188 738 -164
rect 163 -190 164 -164
rect 408 -237 409 -189
rect 443 -190 444 -164
rect 478 -237 479 -189
rect 499 -190 500 -164
rect 576 -237 577 -189
rect 632 -190 633 -164
rect 800 -237 801 -189
rect 58 -192 59 -164
rect 163 -237 164 -191
rect 177 -192 178 -164
rect 233 -237 234 -191
rect 296 -192 297 -164
rect 317 -237 318 -191
rect 359 -237 360 -191
rect 737 -237 738 -191
rect 51 -194 52 -164
rect 58 -237 59 -193
rect 177 -237 178 -193
rect 247 -194 248 -164
rect 282 -194 283 -164
rect 296 -237 297 -193
rect 366 -237 367 -193
rect 401 -194 402 -164
rect 443 -237 444 -193
rect 481 -194 482 -164
rect 520 -194 521 -164
rect 523 -212 524 -193
rect 548 -237 549 -193
rect 562 -194 563 -164
rect 660 -194 661 -164
rect 723 -237 724 -193
rect 730 -237 731 -193
rect 859 -237 860 -193
rect 51 -237 52 -195
rect 387 -196 388 -164
rect 450 -196 451 -164
rect 632 -237 633 -195
rect 667 -196 668 -164
rect 695 -237 696 -195
rect 709 -196 710 -164
rect 751 -237 752 -195
rect 191 -237 192 -197
rect 219 -198 220 -164
rect 247 -237 248 -197
rect 380 -198 381 -164
rect 429 -198 430 -164
rect 450 -237 451 -197
rect 457 -198 458 -164
rect 499 -237 500 -197
rect 520 -237 521 -197
rect 534 -198 535 -164
rect 618 -198 619 -164
rect 660 -237 661 -197
rect 681 -198 682 -164
rect 779 -237 780 -197
rect 205 -200 206 -164
rect 219 -237 220 -199
rect 226 -237 227 -199
rect 457 -237 458 -199
rect 474 -200 475 -164
rect 667 -237 668 -199
rect 688 -200 689 -164
rect 744 -237 745 -199
rect 205 -237 206 -201
rect 254 -202 255 -164
rect 303 -202 304 -164
rect 380 -237 381 -201
rect 394 -202 395 -164
rect 429 -237 430 -201
rect 439 -237 440 -201
rect 618 -237 619 -201
rect 646 -202 647 -164
rect 688 -237 689 -201
rect 702 -202 703 -164
rect 709 -237 710 -201
rect 716 -202 717 -164
rect 772 -237 773 -201
rect 156 -204 157 -164
rect 394 -237 395 -203
rect 474 -237 475 -203
rect 541 -204 542 -164
rect 653 -204 654 -164
rect 681 -237 682 -203
rect 114 -206 115 -164
rect 156 -237 157 -205
rect 254 -237 255 -205
rect 268 -237 269 -205
rect 289 -206 290 -164
rect 303 -237 304 -205
rect 331 -206 332 -164
rect 401 -237 402 -205
rect 404 -237 405 -205
rect 541 -237 542 -205
rect 639 -206 640 -164
rect 653 -237 654 -205
rect 674 -206 675 -164
rect 702 -237 703 -205
rect 289 -237 290 -207
rect 646 -237 647 -207
rect 331 -237 332 -209
rect 436 -210 437 -164
rect 492 -237 493 -209
rect 716 -237 717 -209
rect 338 -212 339 -164
rect 436 -237 437 -211
rect 534 -237 535 -211
rect 569 -212 570 -164
rect 639 -237 640 -211
rect 261 -214 262 -164
rect 338 -237 339 -213
rect 373 -214 374 -164
rect 387 -237 388 -213
rect 527 -214 528 -164
rect 562 -237 563 -213
rect 611 -214 612 -164
rect 674 -237 675 -213
rect 261 -237 262 -215
rect 345 -216 346 -164
rect 506 -216 507 -164
rect 527 -237 528 -215
rect 555 -216 556 -164
rect 569 -237 570 -215
rect 583 -216 584 -164
rect 611 -237 612 -215
rect 107 -218 108 -164
rect 583 -237 584 -217
rect 107 -237 108 -219
rect 282 -237 283 -219
rect 345 -237 346 -219
rect 625 -220 626 -164
rect 142 -222 143 -164
rect 506 -237 507 -221
rect 597 -222 598 -164
rect 625 -237 626 -221
rect 142 -237 143 -223
rect 376 -237 377 -223
rect 597 -237 598 -223
rect 604 -224 605 -164
rect 149 -226 150 -164
rect 555 -237 556 -225
rect 590 -226 591 -164
rect 604 -237 605 -225
rect 149 -237 150 -227
rect 170 -228 171 -164
rect 513 -228 514 -164
rect 590 -237 591 -227
rect 135 -230 136 -164
rect 170 -237 171 -229
rect 485 -230 486 -164
rect 513 -237 514 -229
rect 93 -232 94 -164
rect 485 -237 486 -231
rect 93 -237 94 -233
rect 152 -234 153 -164
rect 135 -237 136 -235
rect 292 -237 293 -235
rect 2 -326 3 -246
rect 68 -326 69 -246
rect 72 -247 73 -245
rect 348 -247 349 -245
rect 352 -247 353 -245
rect 779 -247 780 -245
rect 807 -247 808 -245
rect 905 -326 906 -246
rect 9 -326 10 -248
rect 285 -249 286 -245
rect 289 -249 290 -245
rect 310 -249 311 -245
rect 352 -326 353 -248
rect 534 -249 535 -245
rect 569 -249 570 -245
rect 940 -326 941 -248
rect 16 -326 17 -250
rect 359 -251 360 -245
rect 383 -326 384 -250
rect 674 -251 675 -245
rect 681 -251 682 -245
rect 891 -326 892 -250
rect 23 -326 24 -252
rect 58 -253 59 -245
rect 72 -326 73 -252
rect 268 -253 269 -245
rect 289 -326 290 -252
rect 450 -253 451 -245
rect 471 -326 472 -252
rect 856 -326 857 -252
rect 30 -326 31 -254
rect 453 -326 454 -254
rect 492 -255 493 -245
rect 611 -255 612 -245
rect 730 -255 731 -245
rect 884 -326 885 -254
rect 37 -326 38 -256
rect 65 -257 66 -245
rect 86 -257 87 -245
rect 292 -257 293 -245
rect 303 -257 304 -245
rect 310 -326 311 -256
rect 359 -326 360 -256
rect 495 -257 496 -245
rect 513 -257 514 -245
rect 513 -326 514 -256
rect 513 -257 514 -245
rect 513 -326 514 -256
rect 520 -257 521 -245
rect 523 -295 524 -256
rect 548 -257 549 -245
rect 611 -326 612 -256
rect 667 -257 668 -245
rect 730 -326 731 -256
rect 744 -257 745 -245
rect 779 -326 780 -256
rect 814 -257 815 -245
rect 954 -326 955 -256
rect 51 -259 52 -245
rect 254 -259 255 -245
rect 268 -326 269 -258
rect 338 -259 339 -245
rect 401 -259 402 -245
rect 590 -259 591 -245
rect 597 -259 598 -245
rect 681 -326 682 -258
rect 758 -259 759 -245
rect 870 -326 871 -258
rect 51 -326 52 -260
rect 394 -261 395 -245
rect 418 -326 419 -260
rect 807 -326 808 -260
rect 821 -261 822 -245
rect 919 -326 920 -260
rect 58 -326 59 -262
rect 499 -263 500 -245
rect 506 -263 507 -245
rect 744 -326 745 -262
rect 758 -326 759 -262
rect 800 -263 801 -245
rect 828 -263 829 -245
rect 926 -326 927 -262
rect 65 -326 66 -264
rect 912 -326 913 -264
rect 79 -267 80 -245
rect 86 -326 87 -266
rect 93 -267 94 -245
rect 282 -267 283 -245
rect 303 -326 304 -266
rect 306 -326 307 -266
rect 376 -267 377 -245
rect 499 -326 500 -266
rect 520 -326 521 -266
rect 555 -267 556 -245
rect 674 -326 675 -266
rect 751 -267 752 -245
rect 800 -326 801 -266
rect 835 -267 836 -245
rect 933 -326 934 -266
rect 79 -326 80 -268
rect 443 -269 444 -245
rect 464 -269 465 -245
rect 506 -326 507 -268
rect 541 -269 542 -245
rect 555 -326 556 -268
rect 569 -326 570 -268
rect 597 -326 598 -268
rect 653 -269 654 -245
rect 667 -326 668 -268
rect 723 -269 724 -245
rect 751 -326 752 -268
rect 765 -269 766 -245
rect 828 -326 829 -268
rect 842 -269 843 -245
rect 947 -326 948 -268
rect 93 -326 94 -270
rect 100 -271 101 -245
rect 103 -271 104 -245
rect 590 -326 591 -270
rect 632 -271 633 -245
rect 653 -326 654 -270
rect 709 -271 710 -245
rect 723 -326 724 -270
rect 793 -271 794 -245
rect 814 -326 815 -270
rect 849 -271 850 -245
rect 877 -326 878 -270
rect 100 -326 101 -272
rect 415 -273 416 -245
rect 425 -273 426 -245
rect 863 -273 864 -245
rect 121 -275 122 -245
rect 163 -275 164 -245
rect 170 -275 171 -245
rect 282 -326 283 -274
rect 338 -326 339 -274
rect 376 -326 377 -274
rect 387 -275 388 -245
rect 443 -326 444 -274
rect 450 -326 451 -274
rect 842 -326 843 -274
rect 121 -326 122 -276
rect 366 -277 367 -245
rect 394 -326 395 -276
rect 688 -277 689 -245
rect 702 -277 703 -245
rect 863 -326 864 -276
rect 142 -279 143 -245
rect 257 -279 258 -245
rect 366 -326 367 -278
rect 548 -326 549 -278
rect 576 -279 577 -245
rect 579 -279 580 -245
rect 583 -279 584 -245
rect 632 -326 633 -278
rect 646 -279 647 -245
rect 702 -326 703 -278
rect 772 -279 773 -245
rect 849 -326 850 -278
rect 142 -326 143 -280
rect 467 -326 468 -280
rect 474 -281 475 -245
rect 541 -326 542 -280
rect 576 -326 577 -280
rect 604 -281 605 -245
rect 625 -281 626 -245
rect 646 -326 647 -280
rect 660 -281 661 -245
rect 709 -326 710 -280
rect 716 -281 717 -245
rect 772 -326 773 -280
rect 786 -281 787 -245
rect 793 -326 794 -280
rect 149 -283 150 -245
rect 149 -326 150 -282
rect 149 -283 150 -245
rect 149 -326 150 -282
rect 156 -283 157 -245
rect 387 -326 388 -282
rect 397 -326 398 -282
rect 821 -326 822 -282
rect 156 -326 157 -284
rect 275 -285 276 -245
rect 425 -326 426 -284
rect 534 -326 535 -284
rect 551 -326 552 -284
rect 716 -326 717 -284
rect 737 -285 738 -245
rect 786 -326 787 -284
rect 163 -326 164 -286
rect 261 -287 262 -245
rect 275 -326 276 -286
rect 345 -287 346 -245
rect 436 -287 437 -245
rect 835 -326 836 -286
rect 44 -289 45 -245
rect 436 -326 437 -288
rect 439 -326 440 -288
rect 765 -326 766 -288
rect 170 -326 171 -290
rect 331 -291 332 -245
rect 457 -291 458 -245
rect 583 -326 584 -290
rect 639 -291 640 -245
rect 660 -326 661 -290
rect 688 -326 689 -290
rect 898 -326 899 -290
rect 128 -293 129 -245
rect 331 -326 332 -292
rect 457 -326 458 -292
rect 639 -326 640 -292
rect 695 -293 696 -245
rect 737 -326 738 -292
rect 177 -295 178 -245
rect 177 -326 178 -294
rect 177 -295 178 -245
rect 177 -326 178 -294
rect 184 -295 185 -245
rect 362 -295 363 -245
rect 478 -295 479 -245
rect 492 -326 493 -294
rect 579 -326 580 -294
rect 604 -326 605 -294
rect 618 -295 619 -245
rect 695 -326 696 -294
rect 166 -297 167 -245
rect 618 -326 619 -296
rect 184 -326 185 -298
rect 191 -299 192 -245
rect 205 -299 206 -245
rect 404 -326 405 -298
rect 478 -326 479 -298
rect 485 -299 486 -245
rect 488 -326 489 -298
rect 625 -326 626 -298
rect 107 -301 108 -245
rect 191 -326 192 -300
rect 205 -326 206 -300
rect 219 -301 220 -245
rect 240 -301 241 -245
rect 240 -326 241 -300
rect 240 -301 241 -245
rect 240 -326 241 -300
rect 254 -326 255 -300
rect 474 -326 475 -300
rect 485 -326 486 -300
rect 562 -301 563 -245
rect 107 -326 108 -302
rect 124 -303 125 -245
rect 219 -326 220 -302
rect 233 -303 234 -245
rect 261 -326 262 -302
rect 422 -303 423 -245
rect 446 -326 447 -302
rect 562 -326 563 -302
rect 198 -305 199 -245
rect 233 -326 234 -304
rect 247 -305 248 -245
rect 422 -326 423 -304
rect 114 -307 115 -245
rect 247 -326 248 -306
rect 317 -307 318 -245
rect 345 -326 346 -306
rect 114 -326 115 -308
rect 429 -309 430 -245
rect 198 -326 199 -310
rect 296 -311 297 -245
rect 380 -311 381 -245
rect 429 -326 430 -310
rect 44 -326 45 -312
rect 380 -326 381 -312
rect 135 -315 136 -245
rect 296 -326 297 -314
rect 135 -326 136 -316
rect 212 -317 213 -245
rect 226 -317 227 -245
rect 317 -326 318 -316
rect 212 -326 213 -318
rect 324 -319 325 -245
rect 226 -326 227 -320
rect 408 -321 409 -245
rect 117 -323 118 -245
rect 408 -326 409 -322
rect 324 -326 325 -324
rect 355 -325 356 -245
rect 16 -336 17 -334
rect 415 -336 416 -334
rect 436 -336 437 -334
rect 681 -336 682 -334
rect 905 -336 906 -334
rect 961 -413 962 -335
rect 16 -413 17 -337
rect 107 -338 108 -334
rect 124 -413 125 -337
rect 282 -338 283 -334
rect 289 -338 290 -334
rect 397 -338 398 -334
rect 401 -338 402 -334
rect 695 -338 696 -334
rect 758 -338 759 -334
rect 905 -413 906 -337
rect 912 -338 913 -334
rect 1024 -413 1025 -337
rect 44 -340 45 -334
rect 75 -413 76 -339
rect 79 -340 80 -334
rect 415 -413 416 -339
rect 439 -340 440 -334
rect 572 -340 573 -334
rect 618 -340 619 -334
rect 1003 -413 1004 -339
rect 37 -342 38 -334
rect 79 -413 80 -341
rect 96 -413 97 -341
rect 681 -413 682 -341
rect 730 -342 731 -334
rect 758 -413 759 -341
rect 779 -342 780 -334
rect 912 -413 913 -341
rect 919 -342 920 -334
rect 982 -413 983 -341
rect 2 -344 3 -334
rect 37 -413 38 -343
rect 44 -413 45 -343
rect 93 -344 94 -334
rect 100 -344 101 -334
rect 282 -413 283 -343
rect 296 -344 297 -334
rect 303 -413 304 -343
rect 310 -344 311 -334
rect 460 -344 461 -334
rect 467 -344 468 -334
rect 884 -344 885 -334
rect 926 -344 927 -334
rect 989 -413 990 -343
rect 2 -413 3 -345
rect 345 -346 346 -334
rect 355 -413 356 -345
rect 436 -413 437 -345
rect 443 -346 444 -334
rect 996 -413 997 -345
rect 51 -348 52 -334
rect 460 -413 461 -347
rect 467 -413 468 -347
rect 898 -348 899 -334
rect 933 -348 934 -334
rect 975 -413 976 -347
rect 51 -413 52 -349
rect 488 -350 489 -334
rect 548 -350 549 -334
rect 968 -413 969 -349
rect 65 -413 66 -351
rect 163 -352 164 -334
rect 191 -413 192 -351
rect 310 -413 311 -351
rect 331 -352 332 -334
rect 401 -413 402 -351
rect 411 -413 412 -351
rect 940 -352 941 -334
rect 947 -352 948 -334
rect 947 -413 948 -351
rect 947 -352 948 -334
rect 947 -413 948 -351
rect 93 -413 94 -353
rect 198 -354 199 -334
rect 205 -354 206 -334
rect 205 -413 206 -353
rect 205 -354 206 -334
rect 205 -413 206 -353
rect 212 -354 213 -334
rect 453 -354 454 -334
rect 457 -354 458 -334
rect 954 -354 955 -334
rect 100 -413 101 -355
rect 142 -356 143 -334
rect 149 -356 150 -334
rect 163 -413 164 -355
rect 198 -413 199 -355
rect 233 -356 234 -334
rect 243 -413 244 -355
rect 289 -413 290 -355
rect 296 -413 297 -355
rect 530 -413 531 -355
rect 583 -356 584 -334
rect 618 -413 619 -355
rect 621 -413 622 -355
rect 779 -413 780 -355
rect 793 -356 794 -334
rect 933 -413 934 -355
rect 107 -413 108 -357
rect 131 -358 132 -334
rect 142 -413 143 -357
rect 219 -358 220 -334
rect 226 -358 227 -334
rect 418 -358 419 -334
rect 422 -358 423 -334
rect 884 -413 885 -357
rect 72 -360 73 -334
rect 226 -413 227 -359
rect 233 -413 234 -359
rect 376 -360 377 -334
rect 380 -413 381 -359
rect 551 -360 552 -334
rect 667 -360 668 -334
rect 695 -413 696 -359
rect 751 -360 752 -334
rect 793 -413 794 -359
rect 800 -360 801 -334
rect 919 -413 920 -359
rect 114 -362 115 -334
rect 397 -413 398 -361
rect 446 -362 447 -334
rect 632 -362 633 -334
rect 744 -362 745 -334
rect 800 -413 801 -361
rect 842 -362 843 -334
rect 898 -413 899 -361
rect 86 -364 87 -334
rect 114 -413 115 -363
rect 177 -364 178 -334
rect 219 -413 220 -363
rect 254 -364 255 -334
rect 383 -364 384 -334
rect 387 -364 388 -334
rect 422 -413 423 -363
rect 457 -413 458 -363
rect 576 -364 577 -334
rect 597 -364 598 -334
rect 667 -413 668 -363
rect 702 -364 703 -334
rect 744 -413 745 -363
rect 786 -364 787 -334
rect 842 -413 843 -363
rect 849 -364 850 -334
rect 926 -413 927 -363
rect 177 -413 178 -365
rect 184 -366 185 -334
rect 194 -413 195 -365
rect 702 -413 703 -365
rect 737 -366 738 -334
rect 786 -413 787 -365
rect 814 -366 815 -334
rect 849 -413 850 -365
rect 856 -366 857 -334
rect 940 -413 941 -365
rect 128 -368 129 -334
rect 184 -413 185 -367
rect 254 -413 255 -367
rect 275 -368 276 -334
rect 338 -368 339 -334
rect 443 -413 444 -367
rect 464 -368 465 -334
rect 856 -413 857 -367
rect 877 -368 878 -334
rect 954 -413 955 -367
rect 128 -413 129 -369
rect 135 -370 136 -334
rect 156 -370 157 -334
rect 338 -413 339 -369
rect 352 -370 353 -334
rect 597 -413 598 -369
rect 632 -413 633 -369
rect 639 -370 640 -334
rect 660 -370 661 -334
rect 737 -413 738 -369
rect 835 -370 836 -334
rect 877 -413 878 -369
rect 86 -413 87 -371
rect 135 -413 136 -371
rect 156 -413 157 -371
rect 317 -372 318 -334
rect 359 -372 360 -334
rect 474 -372 475 -334
rect 485 -372 486 -334
rect 730 -413 731 -371
rect 772 -372 773 -334
rect 835 -413 836 -371
rect 170 -374 171 -334
rect 352 -413 353 -373
rect 373 -374 374 -334
rect 870 -374 871 -334
rect 82 -413 83 -375
rect 170 -413 171 -375
rect 212 -413 213 -375
rect 359 -413 360 -375
rect 387 -413 388 -375
rect 429 -376 430 -334
rect 464 -413 465 -375
rect 485 -413 486 -375
rect 516 -413 517 -375
rect 639 -413 640 -375
rect 646 -376 647 -334
rect 660 -413 661 -375
rect 709 -376 710 -334
rect 870 -413 871 -375
rect 261 -378 262 -334
rect 345 -413 346 -377
rect 425 -378 426 -334
rect 576 -413 577 -377
rect 653 -378 654 -334
rect 709 -413 710 -377
rect 723 -378 724 -334
rect 814 -413 815 -377
rect 247 -380 248 -334
rect 261 -413 262 -379
rect 268 -380 269 -334
rect 373 -413 374 -379
rect 429 -413 430 -379
rect 450 -413 451 -379
rect 471 -380 472 -334
rect 863 -380 864 -334
rect 72 -413 73 -381
rect 471 -413 472 -381
rect 541 -382 542 -334
rect 583 -413 584 -381
rect 625 -382 626 -334
rect 653 -413 654 -381
rect 674 -382 675 -334
rect 723 -413 724 -381
rect 821 -382 822 -334
rect 863 -413 864 -381
rect 121 -384 122 -334
rect 268 -413 269 -383
rect 275 -413 276 -383
rect 394 -384 395 -334
rect 506 -384 507 -334
rect 541 -413 542 -383
rect 551 -413 552 -383
rect 772 -413 773 -383
rect 23 -386 24 -334
rect 121 -413 122 -385
rect 240 -386 241 -334
rect 247 -413 248 -385
rect 306 -386 307 -334
rect 646 -413 647 -385
rect 765 -386 766 -334
rect 821 -413 822 -385
rect 23 -413 24 -387
rect 30 -388 31 -334
rect 58 -388 59 -334
rect 506 -413 507 -387
rect 520 -388 521 -334
rect 625 -413 626 -387
rect 716 -388 717 -334
rect 765 -413 766 -387
rect 30 -413 31 -389
rect 68 -390 69 -334
rect 149 -413 150 -389
rect 240 -413 241 -389
rect 317 -413 318 -389
rect 366 -390 367 -334
rect 394 -413 395 -389
rect 807 -390 808 -334
rect 58 -413 59 -391
rect 324 -392 325 -334
rect 362 -413 363 -391
rect 674 -413 675 -391
rect 688 -392 689 -334
rect 716 -413 717 -391
rect 68 -413 69 -393
rect 331 -413 332 -393
rect 366 -413 367 -393
rect 432 -413 433 -393
rect 513 -394 514 -334
rect 520 -413 521 -393
rect 562 -394 563 -334
rect 688 -413 689 -393
rect 324 -413 325 -395
rect 555 -396 556 -334
rect 569 -396 570 -334
rect 751 -413 752 -395
rect 499 -398 500 -334
rect 562 -413 563 -397
rect 569 -413 570 -397
rect 611 -398 612 -334
rect 478 -400 479 -334
rect 499 -413 500 -399
rect 513 -413 514 -399
rect 891 -400 892 -334
rect 478 -413 479 -401
rect 492 -402 493 -334
rect 527 -402 528 -334
rect 555 -413 556 -401
rect 590 -402 591 -334
rect 611 -413 612 -401
rect 828 -402 829 -334
rect 891 -413 892 -401
rect 9 -404 10 -334
rect 527 -413 528 -403
rect 534 -404 535 -334
rect 590 -413 591 -403
rect 604 -404 605 -334
rect 807 -413 808 -403
rect 9 -413 10 -405
rect 89 -413 90 -405
rect 159 -413 160 -405
rect 828 -413 829 -405
rect 404 -408 405 -334
rect 604 -413 605 -407
rect 408 -410 409 -334
rect 534 -413 535 -409
rect 408 -413 409 -411
rect 492 -413 493 -411
rect 9 -423 10 -421
rect 131 -508 132 -422
rect 142 -423 143 -421
rect 243 -423 244 -421
rect 275 -423 276 -421
rect 352 -508 353 -422
rect 362 -423 363 -421
rect 625 -423 626 -421
rect 695 -423 696 -421
rect 695 -508 696 -422
rect 695 -423 696 -421
rect 695 -508 696 -422
rect 814 -423 815 -421
rect 1073 -508 1074 -422
rect 9 -508 10 -424
rect 639 -425 640 -421
rect 849 -425 850 -421
rect 1045 -508 1046 -424
rect 16 -427 17 -421
rect 93 -427 94 -421
rect 114 -427 115 -421
rect 114 -508 115 -426
rect 114 -427 115 -421
rect 114 -508 115 -426
rect 156 -427 157 -421
rect 282 -427 283 -421
rect 324 -427 325 -421
rect 411 -427 412 -421
rect 415 -427 416 -421
rect 814 -508 815 -426
rect 912 -427 913 -421
rect 1031 -508 1032 -426
rect 16 -508 17 -428
rect 653 -429 654 -421
rect 765 -429 766 -421
rect 849 -508 850 -428
rect 926 -429 927 -421
rect 1052 -508 1053 -428
rect 23 -431 24 -421
rect 152 -508 153 -430
rect 191 -431 192 -421
rect 422 -431 423 -421
rect 429 -431 430 -421
rect 807 -431 808 -421
rect 828 -431 829 -421
rect 926 -508 927 -430
rect 933 -431 934 -421
rect 1010 -508 1011 -430
rect 1024 -431 1025 -421
rect 1087 -508 1088 -430
rect 23 -508 24 -432
rect 390 -508 391 -432
rect 394 -433 395 -421
rect 807 -508 808 -432
rect 828 -508 829 -432
rect 891 -433 892 -421
rect 940 -433 941 -421
rect 1038 -508 1039 -432
rect 30 -435 31 -421
rect 184 -435 185 -421
rect 198 -435 199 -421
rect 198 -508 199 -434
rect 198 -435 199 -421
rect 198 -508 199 -434
rect 226 -435 227 -421
rect 327 -508 328 -434
rect 373 -435 374 -421
rect 481 -508 482 -434
rect 513 -508 514 -434
rect 534 -435 535 -421
rect 548 -435 549 -421
rect 919 -435 920 -421
rect 940 -508 941 -434
rect 1003 -435 1004 -421
rect 30 -508 31 -436
rect 58 -437 59 -421
rect 65 -437 66 -421
rect 359 -437 360 -421
rect 397 -437 398 -421
rect 667 -437 668 -421
rect 670 -508 671 -436
rect 1003 -508 1004 -436
rect 37 -439 38 -421
rect 72 -439 73 -421
rect 86 -508 87 -438
rect 100 -439 101 -421
rect 163 -439 164 -421
rect 191 -508 192 -438
rect 219 -439 220 -421
rect 226 -508 227 -438
rect 275 -508 276 -438
rect 397 -508 398 -438
rect 401 -439 402 -421
rect 415 -508 416 -438
rect 432 -439 433 -421
rect 716 -439 717 -421
rect 730 -439 731 -421
rect 1024 -508 1025 -438
rect 37 -508 38 -440
rect 93 -508 94 -440
rect 100 -508 101 -440
rect 107 -441 108 -421
rect 184 -508 185 -440
rect 317 -441 318 -421
rect 324 -508 325 -440
rect 422 -508 423 -440
rect 450 -441 451 -421
rect 453 -505 454 -440
rect 467 -441 468 -421
rect 478 -441 479 -421
rect 523 -508 524 -440
rect 1101 -508 1102 -440
rect 44 -443 45 -421
rect 79 -443 80 -421
rect 187 -443 188 -421
rect 219 -508 220 -442
rect 296 -443 297 -421
rect 429 -508 430 -442
rect 450 -508 451 -442
rect 723 -443 724 -421
rect 730 -508 731 -442
rect 751 -443 752 -421
rect 786 -443 787 -421
rect 891 -508 892 -442
rect 954 -443 955 -421
rect 1059 -508 1060 -442
rect 44 -508 45 -444
rect 250 -508 251 -444
rect 310 -445 311 -421
rect 317 -508 318 -444
rect 331 -445 332 -421
rect 373 -508 374 -444
rect 401 -508 402 -444
rect 411 -508 412 -444
rect 478 -508 479 -444
rect 905 -445 906 -421
rect 961 -445 962 -421
rect 1094 -508 1095 -444
rect 51 -447 52 -421
rect 240 -447 241 -421
rect 247 -447 248 -421
rect 296 -508 297 -446
rect 331 -508 332 -446
rect 366 -447 367 -421
rect 460 -447 461 -421
rect 961 -508 962 -446
rect 968 -447 969 -421
rect 1108 -508 1109 -446
rect 51 -508 52 -448
rect 485 -449 486 -421
rect 530 -449 531 -421
rect 870 -449 871 -421
rect 975 -449 976 -421
rect 1080 -508 1081 -448
rect 58 -508 59 -450
rect 551 -451 552 -421
rect 555 -451 556 -421
rect 555 -508 556 -450
rect 555 -451 556 -421
rect 555 -508 556 -450
rect 562 -451 563 -421
rect 639 -508 640 -450
rect 649 -508 650 -450
rect 765 -508 766 -450
rect 772 -451 773 -421
rect 870 -508 871 -450
rect 884 -451 885 -421
rect 975 -508 976 -450
rect 982 -451 983 -421
rect 1115 -508 1116 -450
rect 65 -508 66 -452
rect 387 -453 388 -421
rect 408 -453 409 -421
rect 562 -508 563 -452
rect 576 -453 577 -421
rect 625 -508 626 -452
rect 674 -453 675 -421
rect 905 -508 906 -452
rect 989 -453 990 -421
rect 1122 -508 1123 -452
rect 68 -455 69 -421
rect 716 -508 717 -454
rect 737 -455 738 -421
rect 989 -508 990 -454
rect 996 -455 997 -421
rect 1066 -508 1067 -454
rect 72 -508 73 -456
rect 667 -508 668 -456
rect 709 -457 710 -421
rect 786 -508 787 -456
rect 800 -457 801 -421
rect 912 -508 913 -456
rect 75 -459 76 -421
rect 107 -508 108 -458
rect 121 -459 122 -421
rect 884 -508 885 -458
rect 79 -508 80 -460
rect 170 -461 171 -421
rect 205 -461 206 -421
rect 247 -508 248 -460
rect 261 -461 262 -421
rect 366 -508 367 -460
rect 387 -508 388 -460
rect 1017 -508 1018 -460
rect 82 -463 83 -421
rect 772 -508 773 -462
rect 779 -463 780 -421
rect 954 -508 955 -462
rect 121 -508 122 -464
rect 177 -465 178 -421
rect 233 -465 234 -421
rect 408 -508 409 -464
rect 485 -508 486 -464
rect 576 -508 577 -464
rect 597 -465 598 -421
rect 653 -508 654 -464
rect 702 -465 703 -421
rect 709 -508 710 -464
rect 744 -465 745 -421
rect 800 -508 801 -464
rect 821 -465 822 -421
rect 919 -508 920 -464
rect 128 -467 129 -421
rect 170 -508 171 -466
rect 177 -508 178 -466
rect 380 -467 381 -421
rect 520 -467 521 -421
rect 597 -508 598 -466
rect 604 -467 605 -421
rect 674 -508 675 -466
rect 681 -467 682 -421
rect 744 -508 745 -466
rect 835 -467 836 -421
rect 933 -508 934 -466
rect 96 -469 97 -421
rect 128 -508 129 -468
rect 135 -469 136 -421
rect 310 -508 311 -468
rect 338 -469 339 -421
rect 359 -508 360 -468
rect 464 -469 465 -421
rect 835 -508 836 -468
rect 856 -469 857 -421
rect 982 -508 983 -468
rect 96 -508 97 -470
rect 163 -508 164 -470
rect 212 -471 213 -421
rect 380 -508 381 -470
rect 464 -508 465 -470
rect 527 -471 528 -421
rect 534 -508 535 -470
rect 579 -508 580 -470
rect 607 -508 608 -470
rect 702 -508 703 -470
rect 793 -471 794 -421
rect 856 -508 857 -470
rect 863 -471 864 -421
rect 968 -508 969 -470
rect 156 -508 157 -472
rect 338 -508 339 -472
rect 471 -473 472 -421
rect 527 -508 528 -472
rect 548 -508 549 -472
rect 751 -508 752 -472
rect 758 -473 759 -421
rect 863 -508 864 -472
rect 877 -473 878 -421
rect 996 -508 997 -472
rect 149 -475 150 -421
rect 471 -508 472 -474
rect 509 -508 510 -474
rect 793 -508 794 -474
rect 212 -508 213 -476
rect 303 -477 304 -421
rect 516 -477 517 -421
rect 877 -508 878 -476
rect 2 -479 3 -421
rect 303 -508 304 -478
rect 520 -508 521 -478
rect 688 -479 689 -421
rect 2 -508 3 -480
rect 138 -508 139 -480
rect 233 -508 234 -480
rect 254 -481 255 -421
rect 261 -508 262 -480
rect 268 -481 269 -421
rect 572 -508 573 -480
rect 758 -508 759 -480
rect 124 -483 125 -421
rect 268 -508 269 -482
rect 604 -508 605 -482
rect 688 -508 689 -482
rect 240 -508 241 -484
rect 289 -485 290 -421
rect 611 -485 612 -421
rect 779 -508 780 -484
rect 254 -508 255 -486
rect 443 -487 444 -421
rect 618 -487 619 -421
rect 723 -508 724 -486
rect 205 -508 206 -488
rect 443 -508 444 -488
rect 569 -489 570 -421
rect 618 -508 619 -488
rect 621 -489 622 -421
rect 947 -489 948 -421
rect 289 -508 290 -490
rect 499 -491 500 -421
rect 569 -508 570 -490
rect 898 -491 899 -421
rect 345 -493 346 -421
rect 611 -508 612 -492
rect 632 -493 633 -421
rect 737 -508 738 -492
rect 842 -493 843 -421
rect 947 -508 948 -492
rect 159 -495 160 -421
rect 345 -508 346 -494
rect 436 -495 437 -421
rect 499 -508 500 -494
rect 583 -495 584 -421
rect 842 -508 843 -494
rect 394 -508 395 -496
rect 436 -508 437 -496
rect 446 -508 447 -496
rect 632 -508 633 -496
rect 646 -497 647 -421
rect 821 -508 822 -496
rect 457 -499 458 -421
rect 898 -508 899 -498
rect 457 -508 458 -500
rect 541 -501 542 -421
rect 583 -508 584 -500
rect 590 -501 591 -421
rect 660 -501 661 -421
rect 681 -508 682 -500
rect 492 -503 493 -421
rect 541 -508 542 -502
rect 565 -508 566 -502
rect 660 -508 661 -502
rect 492 -508 493 -504
rect 506 -505 507 -421
rect 590 -508 591 -504
rect 282 -508 283 -506
rect 506 -508 507 -506
rect 2 -518 3 -516
rect 142 -607 143 -517
rect 149 -607 150 -517
rect 383 -607 384 -517
rect 390 -607 391 -517
rect 408 -607 409 -517
rect 411 -518 412 -516
rect 821 -518 822 -516
rect 1087 -518 1088 -516
rect 1087 -607 1088 -517
rect 1087 -518 1088 -516
rect 1087 -607 1088 -517
rect 2 -607 3 -519
rect 404 -607 405 -519
rect 425 -607 426 -519
rect 478 -520 479 -516
rect 509 -520 510 -516
rect 1115 -520 1116 -516
rect 9 -522 10 -516
rect 138 -522 139 -516
rect 159 -522 160 -516
rect 450 -522 451 -516
rect 544 -607 545 -521
rect 1108 -522 1109 -516
rect 9 -607 10 -523
rect 786 -524 787 -516
rect 821 -607 822 -523
rect 849 -524 850 -516
rect 16 -526 17 -516
rect 93 -526 94 -516
rect 107 -526 108 -516
rect 128 -526 129 -516
rect 177 -526 178 -516
rect 478 -607 479 -525
rect 572 -526 573 -516
rect 989 -526 990 -516
rect 58 -528 59 -516
rect 562 -528 563 -516
rect 576 -528 577 -516
rect 842 -528 843 -516
rect 989 -607 990 -527
rect 1017 -528 1018 -516
rect 72 -530 73 -516
rect 156 -530 157 -516
rect 177 -607 178 -529
rect 187 -607 188 -529
rect 212 -530 213 -516
rect 562 -607 563 -529
rect 579 -530 580 -516
rect 1122 -530 1123 -516
rect 75 -607 76 -531
rect 380 -532 381 -516
rect 429 -532 430 -516
rect 621 -607 622 -531
rect 628 -607 629 -531
rect 1073 -532 1074 -516
rect 79 -534 80 -516
rect 387 -534 388 -516
rect 415 -534 416 -516
rect 429 -607 430 -533
rect 443 -607 444 -533
rect 464 -534 465 -516
rect 555 -534 556 -516
rect 576 -607 577 -533
rect 646 -534 647 -516
rect 1031 -534 1032 -516
rect 58 -607 59 -535
rect 79 -607 80 -535
rect 86 -536 87 -516
rect 93 -607 94 -535
rect 128 -607 129 -535
rect 303 -536 304 -516
rect 317 -536 318 -516
rect 450 -607 451 -535
rect 464 -607 465 -535
rect 779 -536 780 -516
rect 786 -607 787 -535
rect 947 -536 948 -516
rect 1017 -607 1018 -535
rect 1038 -536 1039 -516
rect 86 -607 87 -537
rect 131 -538 132 -516
rect 145 -538 146 -516
rect 212 -607 213 -537
rect 240 -538 241 -516
rect 324 -607 325 -537
rect 331 -538 332 -516
rect 331 -607 332 -537
rect 331 -538 332 -516
rect 331 -607 332 -537
rect 387 -607 388 -537
rect 590 -538 591 -516
rect 667 -538 668 -516
rect 1094 -538 1095 -516
rect 51 -540 52 -516
rect 590 -607 591 -539
rect 674 -540 675 -516
rect 849 -607 850 -539
rect 947 -607 948 -539
rect 996 -540 997 -516
rect 1031 -607 1032 -539
rect 1045 -540 1046 -516
rect 51 -607 52 -541
rect 597 -542 598 -516
rect 674 -607 675 -541
rect 730 -542 731 -516
rect 754 -542 755 -516
rect 1101 -542 1102 -516
rect 121 -544 122 -516
rect 303 -607 304 -543
rect 446 -544 447 -516
rect 814 -544 815 -516
rect 828 -544 829 -516
rect 1073 -607 1074 -543
rect 72 -607 73 -545
rect 121 -607 122 -545
rect 135 -546 136 -516
rect 240 -607 241 -545
rect 247 -546 248 -516
rect 296 -546 297 -516
rect 481 -546 482 -516
rect 667 -607 668 -545
rect 695 -546 696 -516
rect 698 -552 699 -545
rect 730 -607 731 -545
rect 772 -546 773 -516
rect 807 -546 808 -516
rect 1045 -607 1046 -545
rect 135 -607 136 -547
rect 205 -548 206 -516
rect 247 -607 248 -547
rect 415 -607 416 -547
rect 520 -548 521 -516
rect 646 -607 647 -547
rect 695 -607 696 -547
rect 702 -548 703 -516
rect 772 -607 773 -547
rect 884 -548 885 -516
rect 996 -607 997 -547
rect 1024 -548 1025 -516
rect 1038 -607 1039 -547
rect 1059 -548 1060 -516
rect 145 -607 146 -549
rect 226 -550 227 -516
rect 250 -550 251 -516
rect 317 -607 318 -549
rect 471 -550 472 -516
rect 520 -607 521 -549
rect 551 -607 552 -549
rect 884 -607 885 -549
rect 1059 -607 1060 -549
rect 1066 -550 1067 -516
rect 37 -552 38 -516
rect 226 -607 227 -551
rect 261 -552 262 -516
rect 506 -552 507 -516
rect 555 -607 556 -551
rect 569 -552 570 -516
rect 597 -607 598 -551
rect 639 -552 640 -516
rect 702 -607 703 -551
rect 723 -552 724 -516
rect 1024 -607 1025 -551
rect 44 -554 45 -516
rect 569 -607 570 -553
rect 632 -554 633 -516
rect 807 -607 808 -553
rect 814 -607 815 -553
rect 891 -554 892 -516
rect 940 -554 941 -516
rect 1066 -607 1067 -553
rect 44 -607 45 -555
rect 422 -556 423 -516
rect 436 -556 437 -516
rect 471 -607 472 -555
rect 492 -556 493 -516
rect 506 -607 507 -555
rect 583 -556 584 -516
rect 632 -607 633 -555
rect 639 -607 640 -555
rect 653 -556 654 -516
rect 723 -607 724 -555
rect 800 -556 801 -516
rect 828 -607 829 -555
rect 856 -556 857 -516
rect 940 -607 941 -555
rect 968 -556 969 -516
rect 156 -607 157 -557
rect 191 -558 192 -516
rect 205 -607 206 -557
rect 275 -558 276 -516
rect 289 -558 290 -516
rect 380 -607 381 -557
rect 422 -607 423 -557
rect 779 -607 780 -557
rect 800 -607 801 -557
rect 863 -558 864 -516
rect 114 -560 115 -516
rect 289 -607 290 -559
rect 296 -607 297 -559
rect 401 -560 402 -516
rect 492 -607 493 -559
rect 499 -560 500 -516
rect 583 -607 584 -559
rect 607 -560 608 -516
rect 653 -607 654 -559
rect 660 -560 661 -516
rect 835 -560 836 -516
rect 968 -607 969 -559
rect 100 -562 101 -516
rect 114 -607 115 -561
rect 152 -562 153 -516
rect 275 -607 276 -561
rect 338 -562 339 -516
rect 436 -607 437 -561
rect 499 -607 500 -561
rect 527 -562 528 -516
rect 604 -562 605 -516
rect 891 -607 892 -561
rect 30 -564 31 -516
rect 338 -607 339 -563
rect 401 -607 402 -563
rect 611 -564 612 -516
rect 660 -607 661 -563
rect 688 -564 689 -516
rect 835 -607 836 -563
rect 870 -564 871 -516
rect 30 -607 31 -565
rect 485 -566 486 -516
rect 513 -566 514 -516
rect 527 -607 528 -565
rect 604 -607 605 -565
rect 625 -566 626 -516
rect 842 -607 843 -565
rect 877 -566 878 -516
rect 16 -607 17 -567
rect 625 -607 626 -567
rect 856 -607 857 -567
rect 954 -568 955 -516
rect 100 -607 101 -569
rect 219 -570 220 -516
rect 261 -607 262 -569
rect 278 -607 279 -569
rect 352 -570 353 -516
rect 485 -607 486 -569
rect 513 -607 514 -569
rect 541 -570 542 -516
rect 863 -607 864 -569
rect 898 -570 899 -516
rect 954 -607 955 -569
rect 1003 -570 1004 -516
rect 37 -607 38 -571
rect 219 -607 220 -571
rect 254 -572 255 -516
rect 352 -607 353 -571
rect 394 -572 395 -516
rect 688 -607 689 -571
rect 870 -607 871 -571
rect 905 -572 906 -516
rect 975 -572 976 -516
rect 1003 -607 1004 -571
rect 191 -607 192 -573
rect 233 -574 234 -516
rect 254 -607 255 -573
rect 282 -574 283 -516
rect 394 -607 395 -573
rect 534 -574 535 -516
rect 541 -607 542 -573
rect 716 -574 717 -516
rect 877 -607 878 -573
rect 912 -574 913 -516
rect 975 -607 976 -573
rect 1010 -574 1011 -516
rect 233 -607 234 -575
rect 670 -576 671 -516
rect 716 -607 717 -575
rect 737 -576 738 -516
rect 898 -607 899 -575
rect 919 -576 920 -516
rect 1010 -607 1011 -575
rect 1080 -576 1081 -516
rect 107 -607 108 -577
rect 1080 -607 1081 -577
rect 268 -580 269 -516
rect 268 -607 269 -579
rect 268 -580 269 -516
rect 268 -607 269 -579
rect 282 -607 283 -579
rect 366 -580 367 -516
rect 457 -580 458 -516
rect 534 -607 535 -579
rect 565 -580 566 -516
rect 912 -607 913 -579
rect 919 -607 920 -579
rect 926 -580 927 -516
rect 65 -582 66 -516
rect 366 -607 367 -581
rect 457 -607 458 -581
rect 982 -582 983 -516
rect 65 -607 66 -583
rect 310 -584 311 -516
rect 523 -584 524 -516
rect 611 -607 612 -583
rect 709 -584 710 -516
rect 737 -607 738 -583
rect 751 -584 752 -516
rect 982 -607 983 -583
rect 170 -586 171 -516
rect 310 -607 311 -585
rect 373 -586 374 -516
rect 523 -607 524 -585
rect 565 -607 566 -585
rect 905 -607 906 -585
rect 170 -607 171 -587
rect 198 -588 199 -516
rect 345 -588 346 -516
rect 373 -607 374 -587
rect 681 -588 682 -516
rect 709 -607 710 -587
rect 751 -607 752 -587
rect 765 -588 766 -516
rect 198 -607 199 -589
rect 460 -607 461 -589
rect 618 -590 619 -516
rect 765 -607 766 -589
rect 345 -607 346 -591
rect 359 -592 360 -516
rect 453 -607 454 -591
rect 681 -607 682 -591
rect 758 -592 759 -516
rect 926 -607 927 -591
rect 184 -594 185 -516
rect 359 -607 360 -593
rect 618 -607 619 -593
rect 1052 -594 1053 -516
rect 23 -596 24 -516
rect 184 -607 185 -595
rect 744 -596 745 -516
rect 758 -607 759 -595
rect 933 -596 934 -516
rect 1052 -607 1053 -595
rect 23 -607 24 -597
rect 163 -598 164 -516
rect 744 -607 745 -597
rect 793 -598 794 -516
rect 933 -607 934 -597
rect 961 -598 962 -516
rect 163 -607 164 -599
rect 548 -600 549 -516
rect 334 -607 335 -601
rect 793 -607 794 -601
rect 467 -607 468 -603
rect 961 -607 962 -603
rect 548 -607 549 -605
rect 649 -606 650 -516
rect 23 -617 24 -615
rect 380 -617 381 -615
rect 415 -716 416 -616
rect 436 -617 437 -615
rect 453 -617 454 -615
rect 765 -617 766 -615
rect 905 -617 906 -615
rect 1213 -716 1214 -616
rect 1216 -716 1217 -616
rect 1360 -716 1361 -616
rect 30 -619 31 -615
rect 30 -716 31 -618
rect 30 -619 31 -615
rect 30 -716 31 -618
rect 40 -619 41 -615
rect 586 -619 587 -615
rect 618 -619 619 -615
rect 674 -619 675 -615
rect 716 -619 717 -615
rect 765 -716 766 -618
rect 814 -619 815 -615
rect 905 -716 906 -618
rect 961 -619 962 -615
rect 1157 -716 1158 -618
rect 2 -621 3 -615
rect 674 -716 675 -620
rect 702 -621 703 -615
rect 716 -716 717 -620
rect 723 -621 724 -615
rect 814 -716 815 -620
rect 961 -716 962 -620
rect 982 -621 983 -615
rect 989 -621 990 -615
rect 1101 -716 1102 -620
rect 2 -716 3 -622
rect 940 -623 941 -615
rect 975 -623 976 -615
rect 1094 -716 1095 -622
rect 44 -625 45 -615
rect 618 -716 619 -624
rect 621 -625 622 -615
rect 982 -716 983 -624
rect 996 -625 997 -615
rect 1108 -716 1109 -624
rect 44 -716 45 -626
rect 338 -627 339 -615
rect 352 -627 353 -615
rect 352 -716 353 -626
rect 352 -627 353 -615
rect 352 -716 353 -626
rect 380 -716 381 -626
rect 611 -627 612 -615
rect 635 -716 636 -626
rect 1052 -627 1053 -615
rect 1059 -627 1060 -615
rect 1192 -716 1193 -626
rect 47 -716 48 -628
rect 205 -629 206 -615
rect 229 -716 230 -628
rect 303 -629 304 -615
rect 324 -629 325 -615
rect 338 -716 339 -628
rect 387 -629 388 -615
rect 723 -716 724 -628
rect 726 -716 727 -628
rect 856 -629 857 -615
rect 884 -629 885 -615
rect 975 -716 976 -628
rect 1010 -629 1011 -615
rect 1185 -716 1186 -628
rect 51 -631 52 -615
rect 432 -716 433 -630
rect 460 -631 461 -615
rect 625 -631 626 -615
rect 649 -716 650 -630
rect 1171 -716 1172 -630
rect 58 -633 59 -615
rect 786 -633 787 -615
rect 821 -633 822 -615
rect 856 -716 857 -632
rect 870 -633 871 -615
rect 884 -716 885 -632
rect 891 -633 892 -615
rect 989 -716 990 -632
rect 1031 -633 1032 -615
rect 1129 -716 1130 -632
rect 51 -716 52 -634
rect 58 -716 59 -634
rect 65 -635 66 -615
rect 548 -635 549 -615
rect 551 -635 552 -615
rect 849 -635 850 -615
rect 898 -635 899 -615
rect 1010 -716 1011 -634
rect 1038 -635 1039 -615
rect 1122 -716 1123 -634
rect 65 -716 66 -636
rect 107 -637 108 -615
rect 121 -637 122 -615
rect 324 -716 325 -636
rect 331 -637 332 -615
rect 345 -637 346 -615
rect 404 -637 405 -615
rect 1052 -716 1053 -636
rect 1066 -637 1067 -615
rect 1199 -716 1200 -636
rect 16 -639 17 -615
rect 107 -716 108 -638
rect 121 -716 122 -638
rect 656 -716 657 -638
rect 667 -639 668 -615
rect 702 -716 703 -638
rect 730 -639 731 -615
rect 996 -716 997 -638
rect 1045 -639 1046 -615
rect 1080 -716 1081 -638
rect 1083 -639 1084 -615
rect 1087 -639 1088 -615
rect 16 -716 17 -640
rect 187 -641 188 -615
rect 226 -641 227 -615
rect 387 -716 388 -640
rect 418 -641 419 -615
rect 425 -641 426 -615
rect 464 -641 465 -615
rect 1164 -716 1165 -640
rect 75 -643 76 -615
rect 1003 -643 1004 -615
rect 86 -645 87 -615
rect 205 -716 206 -644
rect 247 -645 248 -615
rect 345 -716 346 -644
rect 422 -645 423 -615
rect 443 -645 444 -615
rect 464 -716 465 -644
rect 513 -645 514 -615
rect 523 -645 524 -615
rect 1024 -645 1025 -615
rect 37 -716 38 -646
rect 86 -716 87 -646
rect 89 -716 90 -646
rect 1178 -716 1179 -646
rect 100 -649 101 -615
rect 467 -649 468 -615
rect 492 -649 493 -615
rect 513 -716 514 -648
rect 541 -649 542 -615
rect 786 -716 787 -648
rect 800 -649 801 -615
rect 870 -716 871 -648
rect 912 -649 913 -615
rect 1003 -716 1004 -648
rect 100 -716 101 -650
rect 390 -651 391 -615
rect 408 -651 409 -615
rect 422 -716 423 -650
rect 478 -651 479 -615
rect 541 -716 542 -650
rect 544 -651 545 -615
rect 751 -651 752 -615
rect 779 -651 780 -615
rect 940 -716 941 -650
rect 947 -651 948 -615
rect 1066 -716 1067 -650
rect 128 -653 129 -615
rect 275 -653 276 -615
rect 289 -653 290 -615
rect 408 -716 409 -652
rect 492 -716 493 -652
rect 660 -653 661 -615
rect 709 -653 710 -615
rect 751 -716 752 -652
rect 807 -653 808 -615
rect 849 -716 850 -652
rect 912 -716 913 -652
rect 926 -653 927 -615
rect 947 -716 948 -652
rect 1017 -653 1018 -615
rect 93 -655 94 -615
rect 128 -716 129 -654
rect 142 -655 143 -615
rect 1143 -716 1144 -654
rect 61 -657 62 -615
rect 142 -716 143 -656
rect 240 -657 241 -615
rect 443 -716 444 -656
rect 502 -716 503 -656
rect 1038 -716 1039 -656
rect 9 -659 10 -615
rect 61 -716 62 -658
rect 93 -716 94 -658
rect 198 -659 199 -615
rect 247 -716 248 -658
rect 282 -659 283 -615
rect 289 -716 290 -658
rect 366 -659 367 -615
rect 394 -659 395 -615
rect 478 -716 479 -658
rect 520 -659 521 -615
rect 800 -716 801 -658
rect 810 -716 811 -658
rect 1087 -716 1088 -658
rect 9 -716 10 -660
rect 369 -716 370 -660
rect 418 -716 419 -660
rect 520 -716 521 -660
rect 548 -716 549 -660
rect 569 -661 570 -615
rect 590 -661 591 -615
rect 611 -716 612 -660
rect 632 -661 633 -615
rect 660 -716 661 -660
rect 709 -716 710 -660
rect 744 -661 745 -615
rect 821 -716 822 -660
rect 919 -661 920 -615
rect 933 -661 934 -615
rect 1017 -716 1018 -660
rect 23 -716 24 -662
rect 366 -716 367 -662
rect 534 -663 535 -615
rect 569 -716 570 -662
rect 576 -663 577 -615
rect 590 -716 591 -662
rect 597 -663 598 -615
rect 625 -716 626 -662
rect 632 -716 633 -662
rect 1115 -716 1116 -662
rect 110 -716 111 -664
rect 394 -716 395 -664
rect 534 -716 535 -664
rect 555 -665 556 -615
rect 558 -716 559 -664
rect 1031 -716 1032 -664
rect 145 -667 146 -615
rect 240 -716 241 -666
rect 261 -667 262 -615
rect 282 -716 283 -666
rect 296 -667 297 -615
rect 436 -716 437 -666
rect 555 -716 556 -666
rect 576 -716 577 -666
rect 597 -716 598 -666
rect 730 -716 731 -666
rect 733 -716 734 -666
rect 1045 -716 1046 -666
rect 198 -716 199 -668
rect 236 -716 237 -668
rect 254 -669 255 -615
rect 261 -716 262 -668
rect 275 -716 276 -668
rect 404 -716 405 -668
rect 562 -669 563 -615
rect 1073 -669 1074 -615
rect 278 -671 279 -615
rect 296 -716 297 -670
rect 303 -716 304 -670
rect 310 -671 311 -615
rect 317 -671 318 -615
rect 331 -716 332 -670
rect 334 -671 335 -615
rect 891 -716 892 -670
rect 954 -671 955 -615
rect 1059 -716 1060 -670
rect 163 -673 164 -615
rect 317 -716 318 -672
rect 457 -673 458 -615
rect 1073 -716 1074 -672
rect 163 -716 164 -674
rect 212 -675 213 -615
rect 268 -675 269 -615
rect 457 -716 458 -674
rect 562 -716 563 -674
rect 758 -675 759 -615
rect 772 -675 773 -615
rect 919 -716 920 -674
rect 968 -675 969 -615
rect 1024 -716 1025 -674
rect 191 -677 192 -615
rect 212 -716 213 -676
rect 219 -677 220 -615
rect 268 -716 269 -676
rect 310 -716 311 -676
rect 485 -677 486 -615
rect 565 -677 566 -615
rect 1136 -716 1137 -676
rect 177 -679 178 -615
rect 191 -716 192 -678
rect 383 -679 384 -615
rect 968 -716 969 -678
rect 177 -716 178 -680
rect 499 -681 500 -615
rect 565 -716 566 -680
rect 1150 -716 1151 -680
rect 149 -683 150 -615
rect 499 -716 500 -682
rect 583 -683 584 -615
rect 772 -716 773 -682
rect 842 -683 843 -615
rect 898 -716 899 -682
rect 149 -716 150 -684
rect 156 -685 157 -615
rect 184 -685 185 -615
rect 219 -716 220 -684
rect 485 -716 486 -684
rect 527 -685 528 -615
rect 583 -716 584 -684
rect 1206 -716 1207 -684
rect 156 -716 157 -686
rect 429 -687 430 -615
rect 506 -687 507 -615
rect 527 -716 528 -686
rect 586 -716 587 -686
rect 758 -716 759 -686
rect 863 -687 864 -615
rect 926 -716 927 -686
rect 72 -689 73 -615
rect 506 -716 507 -688
rect 628 -689 629 -615
rect 842 -716 843 -688
rect 877 -689 878 -615
rect 954 -716 955 -688
rect 72 -716 73 -690
rect 79 -691 80 -615
rect 170 -691 171 -615
rect 184 -716 185 -690
rect 429 -716 430 -690
rect 667 -716 668 -690
rect 695 -691 696 -615
rect 744 -716 745 -690
rect 828 -691 829 -615
rect 863 -716 864 -690
rect 68 -693 69 -615
rect 79 -716 80 -692
rect 114 -693 115 -615
rect 170 -716 171 -692
rect 646 -693 647 -615
rect 933 -716 934 -692
rect 114 -716 115 -694
rect 373 -695 374 -615
rect 681 -695 682 -615
rect 695 -716 696 -694
rect 737 -695 738 -615
rect 779 -716 780 -694
rect 835 -695 836 -615
rect 877 -716 878 -694
rect 373 -716 374 -696
rect 471 -697 472 -615
rect 688 -697 689 -615
rect 828 -716 829 -696
rect 233 -699 234 -615
rect 471 -716 472 -698
rect 653 -699 654 -615
rect 688 -716 689 -698
rect 793 -699 794 -615
rect 835 -716 836 -698
rect 233 -716 234 -700
rect 359 -701 360 -615
rect 383 -716 384 -700
rect 737 -716 738 -700
rect 226 -716 227 -702
rect 359 -716 360 -702
rect 446 -716 447 -702
rect 681 -716 682 -702
rect 254 -716 255 -704
rect 653 -716 654 -704
rect 639 -707 640 -615
rect 793 -716 794 -706
rect 135 -709 136 -615
rect 639 -716 640 -708
rect 135 -716 136 -710
rect 604 -711 605 -615
rect 450 -713 451 -615
rect 604 -716 605 -712
rect 450 -716 451 -714
rect 646 -716 647 -714
rect 2 -726 3 -724
rect 107 -726 108 -724
rect 131 -833 132 -725
rect 310 -726 311 -724
rect 338 -726 339 -724
rect 446 -726 447 -724
rect 464 -726 465 -724
rect 555 -833 556 -725
rect 569 -726 570 -724
rect 572 -833 573 -725
rect 586 -726 587 -724
rect 933 -726 934 -724
rect 1136 -726 1137 -724
rect 1220 -833 1221 -725
rect 1360 -726 1361 -724
rect 1416 -833 1417 -725
rect 2 -833 3 -727
rect 79 -728 80 -724
rect 89 -728 90 -724
rect 194 -728 195 -724
rect 198 -728 199 -724
rect 201 -794 202 -727
rect 254 -728 255 -724
rect 733 -728 734 -724
rect 737 -728 738 -724
rect 737 -833 738 -727
rect 737 -728 738 -724
rect 737 -833 738 -727
rect 828 -728 829 -724
rect 1262 -833 1263 -727
rect 9 -730 10 -724
rect 723 -730 724 -724
rect 726 -730 727 -724
rect 1087 -730 1088 -724
rect 1143 -730 1144 -724
rect 1227 -833 1228 -729
rect 9 -833 10 -731
rect 51 -732 52 -724
rect 79 -833 80 -731
rect 240 -732 241 -724
rect 254 -833 255 -731
rect 373 -732 374 -724
rect 390 -732 391 -724
rect 1206 -732 1207 -724
rect 16 -734 17 -724
rect 61 -734 62 -724
rect 89 -833 90 -733
rect 695 -734 696 -724
rect 705 -833 706 -733
rect 1199 -734 1200 -724
rect 16 -833 17 -735
rect 369 -736 370 -724
rect 401 -833 402 -735
rect 989 -736 990 -724
rect 1017 -736 1018 -724
rect 1087 -833 1088 -735
rect 1164 -736 1165 -724
rect 1241 -833 1242 -735
rect 30 -738 31 -724
rect 110 -738 111 -724
rect 156 -738 157 -724
rect 240 -833 241 -737
rect 338 -833 339 -737
rect 408 -738 409 -724
rect 422 -738 423 -724
rect 464 -833 465 -737
rect 485 -738 486 -724
rect 565 -738 566 -724
rect 611 -738 612 -724
rect 632 -738 633 -724
rect 635 -738 636 -724
rect 1150 -738 1151 -724
rect 1178 -738 1179 -724
rect 1248 -833 1249 -737
rect 37 -740 38 -724
rect 380 -740 381 -724
rect 390 -833 391 -739
rect 422 -833 423 -739
rect 436 -740 437 -724
rect 485 -833 486 -739
rect 495 -833 496 -739
rect 534 -740 535 -724
rect 576 -740 577 -724
rect 611 -833 612 -739
rect 646 -833 647 -739
rect 744 -740 745 -724
rect 828 -833 829 -739
rect 1206 -833 1207 -739
rect 37 -833 38 -741
rect 93 -742 94 -724
rect 100 -742 101 -724
rect 558 -742 559 -724
rect 576 -833 577 -741
rect 625 -742 626 -724
rect 649 -742 650 -724
rect 821 -742 822 -724
rect 905 -742 906 -724
rect 933 -833 934 -741
rect 975 -742 976 -724
rect 989 -833 990 -741
rect 1017 -833 1018 -741
rect 1045 -742 1046 -724
rect 1080 -742 1081 -724
rect 1199 -833 1200 -741
rect 51 -833 52 -743
rect 1213 -744 1214 -724
rect 65 -746 66 -724
rect 93 -833 94 -745
rect 100 -833 101 -745
rect 128 -746 129 -724
rect 142 -746 143 -724
rect 156 -833 157 -745
rect 163 -746 164 -724
rect 366 -746 367 -724
rect 380 -833 381 -745
rect 415 -746 416 -724
rect 443 -746 444 -724
rect 1234 -833 1235 -745
rect 65 -833 66 -747
rect 233 -748 234 -724
rect 289 -748 290 -724
rect 443 -833 444 -747
rect 457 -748 458 -724
rect 632 -833 633 -747
rect 649 -833 650 -747
rect 1171 -748 1172 -724
rect 1185 -748 1186 -724
rect 1255 -833 1256 -747
rect 86 -833 87 -749
rect 1080 -833 1081 -749
rect 1094 -750 1095 -724
rect 1150 -833 1151 -749
rect 1157 -750 1158 -724
rect 1185 -833 1186 -749
rect 107 -833 108 -751
rect 149 -752 150 -724
rect 170 -752 171 -724
rect 173 -794 174 -751
rect 177 -752 178 -724
rect 534 -833 535 -751
rect 590 -752 591 -724
rect 975 -833 976 -751
rect 1101 -752 1102 -724
rect 1178 -833 1179 -751
rect 142 -833 143 -753
rect 387 -754 388 -724
rect 408 -833 409 -753
rect 478 -754 479 -724
rect 502 -754 503 -724
rect 996 -754 997 -724
rect 1108 -754 1109 -724
rect 1171 -833 1172 -753
rect 149 -833 150 -755
rect 513 -756 514 -724
rect 516 -833 517 -755
rect 695 -833 696 -755
rect 709 -756 710 -724
rect 744 -833 745 -755
rect 856 -756 857 -724
rect 905 -833 906 -755
rect 912 -756 913 -724
rect 1045 -833 1046 -755
rect 1115 -756 1116 -724
rect 1164 -833 1165 -755
rect 170 -833 171 -757
rect 205 -758 206 -724
rect 212 -758 213 -724
rect 233 -833 234 -757
rect 299 -833 300 -757
rect 821 -833 822 -757
rect 856 -833 857 -757
rect 968 -758 969 -724
rect 1059 -758 1060 -724
rect 1115 -833 1116 -757
rect 1122 -758 1123 -724
rect 1213 -833 1214 -757
rect 44 -760 45 -724
rect 968 -833 969 -759
rect 44 -833 45 -761
rect 383 -762 384 -724
rect 415 -833 416 -761
rect 681 -762 682 -724
rect 709 -833 710 -761
rect 716 -762 717 -724
rect 723 -833 724 -761
rect 751 -762 752 -724
rect 765 -762 766 -724
rect 912 -833 913 -761
rect 961 -762 962 -724
rect 1094 -833 1095 -761
rect 33 -833 34 -763
rect 751 -833 752 -763
rect 765 -833 766 -763
rect 1052 -764 1053 -724
rect 114 -766 115 -724
rect 681 -833 682 -765
rect 702 -766 703 -724
rect 716 -833 717 -765
rect 730 -766 731 -724
rect 1010 -766 1011 -724
rect 114 -833 115 -767
rect 499 -768 500 -724
rect 506 -768 507 -724
rect 625 -833 626 -767
rect 639 -768 640 -724
rect 1157 -833 1158 -767
rect 128 -833 129 -769
rect 1059 -833 1060 -769
rect 135 -772 136 -724
rect 639 -833 640 -771
rect 653 -772 654 -724
rect 1143 -833 1144 -771
rect 75 -833 76 -773
rect 135 -833 136 -773
rect 191 -774 192 -724
rect 212 -833 213 -773
rect 352 -774 353 -724
rect 404 -774 405 -724
rect 457 -833 458 -773
rect 506 -833 507 -773
rect 513 -833 514 -773
rect 1192 -774 1193 -724
rect 121 -776 122 -724
rect 191 -833 192 -775
rect 198 -833 199 -775
rect 219 -776 220 -724
rect 359 -776 360 -724
rect 373 -833 374 -775
rect 478 -833 479 -775
rect 597 -776 598 -724
rect 656 -776 657 -724
rect 1129 -776 1130 -724
rect 121 -833 122 -777
rect 761 -833 762 -777
rect 870 -778 871 -724
rect 996 -833 997 -777
rect 1024 -778 1025 -724
rect 1129 -833 1130 -777
rect 177 -833 178 -779
rect 352 -833 353 -779
rect 359 -833 360 -779
rect 397 -833 398 -779
rect 432 -780 433 -724
rect 1024 -833 1025 -779
rect 205 -833 206 -781
rect 345 -782 346 -724
rect 366 -833 367 -781
rect 450 -782 451 -724
rect 492 -782 493 -724
rect 1108 -833 1109 -781
rect 184 -784 185 -724
rect 345 -833 346 -783
rect 492 -833 493 -783
rect 793 -784 794 -724
rect 870 -833 871 -783
rect 940 -784 941 -724
rect 947 -784 948 -724
rect 1192 -833 1193 -783
rect 184 -833 185 -785
rect 303 -786 304 -724
rect 520 -786 521 -724
rect 565 -833 566 -785
rect 569 -833 570 -785
rect 1101 -833 1102 -785
rect 23 -788 24 -724
rect 520 -833 521 -787
rect 523 -833 524 -787
rect 919 -788 920 -724
rect 926 -788 927 -724
rect 940 -833 941 -787
rect 954 -788 955 -724
rect 1010 -833 1011 -787
rect 219 -833 220 -789
rect 261 -790 262 -724
rect 275 -790 276 -724
rect 450 -833 451 -789
rect 527 -790 528 -724
rect 954 -833 955 -789
rect 961 -833 962 -789
rect 1003 -790 1004 -724
rect 261 -833 262 -791
rect 282 -792 283 -724
rect 527 -833 528 -791
rect 786 -792 787 -724
rect 877 -792 878 -724
rect 926 -833 927 -791
rect 282 -833 283 -793
rect 583 -794 584 -724
rect 947 -833 948 -793
rect 268 -796 269 -724
rect 275 -833 276 -795
rect 499 -833 500 -795
rect 583 -833 584 -795
rect 586 -833 587 -795
rect 1122 -833 1123 -795
rect 268 -833 269 -797
rect 394 -798 395 -724
rect 590 -833 591 -797
rect 618 -798 619 -724
rect 653 -833 654 -797
rect 793 -833 794 -797
rect 849 -798 850 -724
rect 877 -833 878 -797
rect 898 -798 899 -724
rect 1003 -833 1004 -797
rect 163 -833 164 -799
rect 618 -833 619 -799
rect 656 -833 657 -799
rect 1052 -833 1053 -799
rect 387 -833 388 -801
rect 394 -833 395 -801
rect 429 -802 430 -724
rect 898 -833 899 -801
rect 919 -833 920 -801
rect 982 -802 983 -724
rect 429 -833 430 -803
rect 1136 -833 1137 -803
rect 597 -833 598 -805
rect 674 -806 675 -724
rect 688 -806 689 -724
rect 786 -833 787 -805
rect 814 -806 815 -724
rect 849 -833 850 -805
rect 884 -806 885 -724
rect 982 -833 983 -805
rect 58 -808 59 -724
rect 688 -833 689 -807
rect 702 -833 703 -807
rect 891 -808 892 -724
rect 58 -833 59 -809
rect 72 -810 73 -724
rect 404 -833 405 -809
rect 674 -833 675 -809
rect 779 -810 780 -724
rect 891 -833 892 -809
rect 72 -833 73 -811
rect 289 -833 290 -811
rect 471 -812 472 -724
rect 779 -833 780 -811
rect 800 -812 801 -724
rect 814 -833 815 -811
rect 863 -812 864 -724
rect 884 -833 885 -811
rect 317 -814 318 -724
rect 471 -833 472 -813
rect 604 -814 605 -724
rect 800 -833 801 -813
rect 842 -814 843 -724
rect 863 -833 864 -813
rect 226 -816 227 -724
rect 317 -833 318 -815
rect 548 -816 549 -724
rect 604 -833 605 -815
rect 667 -816 668 -724
rect 730 -833 731 -815
rect 835 -816 836 -724
rect 842 -833 843 -815
rect 226 -833 227 -817
rect 247 -818 248 -724
rect 541 -818 542 -724
rect 548 -833 549 -817
rect 660 -818 661 -724
rect 667 -833 668 -817
rect 807 -818 808 -724
rect 835 -833 836 -817
rect 247 -833 248 -819
rect 324 -820 325 -724
rect 509 -833 510 -819
rect 541 -833 542 -819
rect 562 -820 563 -724
rect 660 -833 661 -819
rect 758 -820 759 -724
rect 807 -833 808 -819
rect 324 -833 325 -821
rect 331 -822 332 -724
rect 562 -833 563 -821
rect 621 -833 622 -821
rect 758 -833 759 -821
rect 1066 -822 1067 -724
rect 296 -824 297 -724
rect 331 -833 332 -823
rect 1031 -824 1032 -724
rect 1066 -833 1067 -823
rect 296 -833 297 -825
rect 1073 -826 1074 -724
rect 432 -833 433 -827
rect 1031 -833 1032 -827
rect 1038 -828 1039 -724
rect 1073 -833 1074 -827
rect 772 -830 773 -724
rect 1038 -833 1039 -829
rect 310 -833 311 -831
rect 772 -833 773 -831
rect 16 -843 17 -841
rect 635 -950 636 -842
rect 649 -843 650 -841
rect 779 -843 780 -841
rect 824 -950 825 -842
rect 1248 -843 1249 -841
rect 1416 -843 1417 -841
rect 1437 -950 1438 -842
rect 16 -950 17 -844
rect 58 -845 59 -841
rect 68 -950 69 -844
rect 338 -845 339 -841
rect 390 -845 391 -841
rect 898 -845 899 -841
rect 961 -845 962 -841
rect 964 -869 965 -844
rect 26 -847 27 -841
rect 44 -847 45 -841
rect 58 -950 59 -846
rect 163 -847 164 -841
rect 170 -847 171 -841
rect 432 -847 433 -841
rect 439 -847 440 -841
rect 1136 -847 1137 -841
rect 30 -849 31 -841
rect 93 -849 94 -841
rect 124 -950 125 -848
rect 1143 -849 1144 -841
rect 30 -950 31 -850
rect 415 -851 416 -841
rect 425 -950 426 -850
rect 786 -851 787 -841
rect 828 -851 829 -841
rect 1220 -851 1221 -841
rect 33 -853 34 -841
rect 947 -853 948 -841
rect 961 -950 962 -852
rect 989 -853 990 -841
rect 1143 -950 1144 -852
rect 1199 -853 1200 -841
rect 37 -855 38 -841
rect 520 -855 521 -841
rect 537 -950 538 -854
rect 576 -855 577 -841
rect 586 -855 587 -841
rect 1010 -855 1011 -841
rect 1129 -855 1130 -841
rect 1199 -950 1200 -854
rect 37 -950 38 -856
rect 51 -857 52 -841
rect 72 -857 73 -841
rect 184 -857 185 -841
rect 198 -857 199 -841
rect 401 -857 402 -841
rect 443 -857 444 -841
rect 516 -857 517 -841
rect 544 -950 545 -856
rect 625 -857 626 -841
rect 653 -857 654 -841
rect 891 -857 892 -841
rect 898 -950 899 -856
rect 940 -857 941 -841
rect 947 -950 948 -856
rect 968 -857 969 -841
rect 1010 -950 1011 -856
rect 1052 -857 1053 -841
rect 44 -950 45 -858
rect 737 -859 738 -841
rect 758 -859 759 -841
rect 1227 -859 1228 -841
rect 51 -950 52 -860
rect 201 -950 202 -860
rect 205 -861 206 -841
rect 583 -861 584 -841
rect 618 -861 619 -841
rect 1003 -861 1004 -841
rect 1052 -950 1053 -860
rect 1202 -950 1203 -860
rect 65 -863 66 -841
rect 72 -950 73 -862
rect 79 -863 80 -841
rect 583 -950 584 -862
rect 611 -863 612 -841
rect 618 -950 619 -862
rect 625 -950 626 -862
rect 1171 -863 1172 -841
rect 65 -950 66 -864
rect 100 -865 101 -841
rect 121 -865 122 -841
rect 415 -950 416 -864
rect 443 -950 444 -864
rect 695 -865 696 -841
rect 702 -865 703 -841
rect 1038 -865 1039 -841
rect 1164 -865 1165 -841
rect 1171 -950 1172 -864
rect 79 -950 80 -866
rect 478 -867 479 -841
rect 485 -867 486 -841
rect 520 -950 521 -866
rect 565 -867 566 -841
rect 1087 -867 1088 -841
rect 86 -869 87 -841
rect 828 -950 829 -868
rect 856 -869 857 -841
rect 940 -950 941 -868
rect 989 -950 990 -868
rect 1003 -950 1004 -868
rect 1045 -869 1046 -841
rect 1059 -869 1060 -841
rect 1164 -950 1165 -868
rect 9 -871 10 -841
rect 86 -950 87 -870
rect 89 -871 90 -841
rect 303 -871 304 -841
rect 380 -871 381 -841
rect 401 -950 402 -870
rect 471 -871 472 -841
rect 485 -950 486 -870
rect 506 -871 507 -841
rect 954 -871 955 -841
rect 968 -950 969 -870
rect 1073 -871 1074 -841
rect 1087 -950 1088 -870
rect 1122 -871 1123 -841
rect 2 -873 3 -841
rect 303 -950 304 -872
rect 331 -873 332 -841
rect 380 -950 381 -872
rect 397 -873 398 -841
rect 1157 -873 1158 -841
rect 23 -875 24 -841
rect 856 -950 857 -874
rect 982 -875 983 -841
rect 1122 -950 1123 -874
rect 23 -950 24 -876
rect 495 -877 496 -841
rect 509 -877 510 -841
rect 660 -877 661 -841
rect 674 -877 675 -841
rect 1059 -950 1060 -876
rect 93 -950 94 -878
rect 215 -950 216 -878
rect 233 -879 234 -841
rect 233 -950 234 -878
rect 233 -879 234 -841
rect 233 -950 234 -878
rect 240 -879 241 -841
rect 394 -879 395 -841
rect 408 -879 409 -841
rect 506 -950 507 -878
rect 569 -879 570 -841
rect 1178 -879 1179 -841
rect 100 -950 101 -880
rect 499 -881 500 -841
rect 572 -881 573 -841
rect 758 -950 759 -880
rect 761 -881 762 -841
rect 954 -950 955 -880
rect 1017 -881 1018 -841
rect 1045 -950 1046 -880
rect 121 -950 122 -882
rect 674 -950 675 -882
rect 688 -883 689 -841
rect 1129 -950 1130 -882
rect 131 -885 132 -841
rect 1178 -950 1179 -884
rect 152 -950 153 -886
rect 982 -950 983 -886
rect 1017 -950 1018 -886
rect 1066 -887 1067 -841
rect 156 -889 157 -841
rect 331 -950 332 -888
rect 369 -950 370 -888
rect 394 -950 395 -888
rect 422 -889 423 -841
rect 471 -950 472 -888
rect 478 -950 479 -888
rect 912 -889 913 -841
rect 1031 -889 1032 -841
rect 1038 -950 1039 -888
rect 2 -950 3 -890
rect 422 -950 423 -890
rect 499 -950 500 -890
rect 975 -891 976 -841
rect 1031 -950 1032 -890
rect 1080 -891 1081 -841
rect 156 -950 157 -892
rect 712 -950 713 -892
rect 723 -893 724 -841
rect 737 -950 738 -892
rect 765 -893 766 -841
rect 1066 -950 1067 -892
rect 1080 -950 1081 -892
rect 1115 -893 1116 -841
rect 89 -950 90 -894
rect 1115 -950 1116 -894
rect 131 -950 132 -896
rect 723 -950 724 -896
rect 730 -897 731 -841
rect 779 -950 780 -896
rect 786 -950 787 -896
rect 863 -897 864 -841
rect 919 -897 920 -841
rect 975 -950 976 -896
rect 163 -950 164 -898
rect 191 -899 192 -841
rect 198 -950 199 -898
rect 240 -950 241 -898
rect 254 -899 255 -841
rect 387 -899 388 -841
rect 611 -950 612 -898
rect 1192 -899 1193 -841
rect 114 -901 115 -841
rect 191 -950 192 -900
rect 205 -950 206 -900
rect 289 -901 290 -841
rect 296 -901 297 -841
rect 345 -901 346 -841
rect 632 -901 633 -841
rect 660 -950 661 -900
rect 695 -950 696 -900
rect 716 -901 717 -841
rect 765 -950 766 -900
rect 800 -901 801 -841
rect 807 -901 808 -841
rect 891 -950 892 -900
rect 919 -950 920 -900
rect 926 -901 927 -841
rect 1094 -901 1095 -841
rect 1192 -950 1193 -900
rect 107 -903 108 -841
rect 114 -950 115 -902
rect 170 -950 171 -902
rect 404 -903 405 -841
rect 569 -950 570 -902
rect 632 -950 633 -902
rect 646 -903 647 -841
rect 1073 -950 1074 -902
rect 1094 -950 1095 -902
rect 1150 -903 1151 -841
rect 107 -950 108 -904
rect 359 -905 360 -841
rect 590 -905 591 -841
rect 646 -950 647 -904
rect 653 -950 654 -904
rect 996 -905 997 -841
rect 1150 -950 1151 -904
rect 1206 -905 1207 -841
rect 177 -950 178 -906
rect 275 -907 276 -841
rect 282 -907 283 -841
rect 320 -950 321 -906
rect 345 -950 346 -906
rect 562 -907 563 -841
rect 614 -950 615 -906
rect 926 -950 927 -906
rect 996 -950 997 -906
rect 1024 -907 1025 -841
rect 1185 -907 1186 -841
rect 1206 -950 1207 -906
rect 180 -909 181 -841
rect 681 -909 682 -841
rect 702 -950 703 -908
rect 842 -909 843 -841
rect 863 -950 864 -908
rect 933 -909 934 -841
rect 1024 -950 1025 -908
rect 1101 -909 1102 -841
rect 1185 -950 1186 -908
rect 1234 -909 1235 -841
rect 184 -950 185 -910
rect 691 -950 692 -910
rect 709 -911 710 -841
rect 730 -950 731 -910
rect 751 -911 752 -841
rect 800 -950 801 -910
rect 807 -950 808 -910
rect 814 -911 815 -841
rect 870 -911 871 -841
rect 933 -950 934 -910
rect 212 -913 213 -841
rect 359 -950 360 -912
rect 513 -913 514 -841
rect 814 -950 815 -912
rect 870 -950 871 -912
rect 1262 -913 1263 -841
rect 212 -950 213 -914
rect 429 -915 430 -841
rect 555 -915 556 -841
rect 590 -950 591 -914
rect 656 -915 657 -841
rect 905 -915 906 -841
rect 219 -917 220 -841
rect 296 -950 297 -916
rect 299 -917 300 -841
rect 387 -950 388 -916
rect 450 -917 451 -841
rect 555 -950 556 -916
rect 562 -950 563 -916
rect 747 -950 748 -916
rect 772 -917 773 -841
rect 1241 -917 1242 -841
rect 219 -950 220 -918
rect 502 -950 503 -918
rect 527 -919 528 -841
rect 772 -950 773 -918
rect 775 -919 776 -841
rect 842 -950 843 -918
rect 247 -921 248 -841
rect 254 -950 255 -920
rect 261 -921 262 -841
rect 275 -950 276 -920
rect 282 -950 283 -920
rect 436 -921 437 -841
rect 450 -950 451 -920
rect 1136 -950 1137 -920
rect 247 -950 248 -922
rect 831 -923 832 -841
rect 261 -950 262 -924
rect 366 -925 367 -841
rect 373 -925 374 -841
rect 513 -950 514 -924
rect 576 -950 577 -924
rect 656 -950 657 -924
rect 667 -925 668 -841
rect 681 -950 682 -924
rect 709 -950 710 -924
rect 1255 -925 1256 -841
rect 226 -927 227 -841
rect 366 -950 367 -926
rect 436 -950 437 -926
rect 541 -927 542 -841
rect 597 -927 598 -841
rect 905 -950 906 -926
rect 135 -929 136 -841
rect 226 -950 227 -928
rect 268 -929 269 -841
rect 338 -950 339 -928
rect 352 -929 353 -841
rect 429 -950 430 -928
rect 541 -950 542 -928
rect 849 -929 850 -841
rect 135 -950 136 -930
rect 492 -931 493 -841
rect 548 -931 549 -841
rect 597 -950 598 -930
rect 639 -931 640 -841
rect 667 -950 668 -930
rect 716 -950 717 -930
rect 1108 -931 1109 -841
rect 142 -933 143 -841
rect 352 -950 353 -932
rect 457 -933 458 -841
rect 548 -950 549 -932
rect 604 -933 605 -841
rect 639 -950 640 -932
rect 688 -950 689 -932
rect 1108 -950 1109 -932
rect 142 -950 143 -934
rect 705 -935 706 -841
rect 719 -950 720 -934
rect 1101 -950 1102 -934
rect 149 -937 150 -841
rect 492 -950 493 -936
rect 534 -937 535 -841
rect 604 -950 605 -936
rect 744 -937 745 -841
rect 751 -950 752 -936
rect 793 -937 794 -841
rect 912 -950 913 -936
rect 268 -950 269 -938
rect 481 -950 482 -938
rect 534 -950 535 -938
rect 1157 -950 1158 -938
rect 289 -950 290 -940
rect 324 -941 325 -841
rect 457 -950 458 -940
rect 464 -941 465 -841
rect 793 -950 794 -940
rect 835 -941 836 -841
rect 849 -950 850 -940
rect 877 -941 878 -841
rect 310 -943 311 -841
rect 373 -950 374 -942
rect 464 -950 465 -942
rect 523 -943 524 -841
rect 821 -943 822 -841
rect 835 -950 836 -942
rect 877 -950 878 -942
rect 884 -943 885 -841
rect 75 -945 76 -841
rect 310 -950 311 -944
rect 317 -945 318 -841
rect 408 -950 409 -944
rect 821 -950 822 -944
rect 1213 -945 1214 -841
rect 9 -950 10 -946
rect 317 -950 318 -946
rect 324 -950 325 -946
rect 628 -950 629 -946
rect 128 -950 129 -948
rect 884 -950 885 -948
rect 2 -960 3 -958
rect 149 -960 150 -958
rect 152 -960 153 -958
rect 439 -1079 440 -959
rect 485 -960 486 -958
rect 485 -1079 486 -959
rect 485 -960 486 -958
rect 485 -1079 486 -959
rect 502 -960 503 -958
rect 681 -960 682 -958
rect 688 -960 689 -958
rect 919 -960 920 -958
rect 929 -1079 930 -959
rect 1325 -1079 1326 -959
rect 1437 -960 1438 -958
rect 1444 -1079 1445 -959
rect 5 -1079 6 -961
rect 408 -962 409 -958
rect 541 -962 542 -958
rect 1262 -1079 1263 -961
rect 9 -964 10 -958
rect 422 -964 423 -958
rect 548 -964 549 -958
rect 712 -964 713 -958
rect 719 -964 720 -958
rect 1290 -1079 1291 -963
rect 16 -966 17 -958
rect 89 -966 90 -958
rect 103 -1079 104 -965
rect 716 -1079 717 -965
rect 744 -966 745 -958
rect 1122 -966 1123 -958
rect 1136 -966 1137 -958
rect 1269 -1079 1270 -965
rect 16 -1079 17 -967
rect 534 -968 535 -958
rect 558 -1079 559 -967
rect 786 -968 787 -958
rect 863 -968 864 -958
rect 1136 -1079 1137 -967
rect 1143 -968 1144 -958
rect 1304 -1079 1305 -967
rect 30 -970 31 -958
rect 537 -970 538 -958
rect 565 -1079 566 -969
rect 1059 -970 1060 -958
rect 1073 -970 1074 -958
rect 1220 -1079 1221 -969
rect 2 -1079 3 -971
rect 30 -1079 31 -971
rect 33 -1079 34 -971
rect 772 -972 773 -958
rect 866 -1079 867 -971
rect 968 -972 969 -958
rect 1087 -972 1088 -958
rect 1213 -1079 1214 -971
rect 44 -974 45 -958
rect 317 -974 318 -958
rect 320 -974 321 -958
rect 422 -1079 423 -973
rect 502 -1079 503 -973
rect 786 -1079 787 -973
rect 877 -974 878 -958
rect 1122 -1079 1123 -973
rect 1157 -974 1158 -958
rect 1311 -1079 1312 -973
rect 44 -1079 45 -975
rect 170 -976 171 -958
rect 198 -976 199 -958
rect 198 -1079 199 -975
rect 198 -976 199 -958
rect 198 -1079 199 -975
rect 201 -976 202 -958
rect 387 -976 388 -958
rect 611 -976 612 -958
rect 1276 -1079 1277 -975
rect 37 -978 38 -958
rect 170 -1079 171 -977
rect 212 -978 213 -958
rect 726 -1079 727 -977
rect 744 -1079 745 -977
rect 863 -1079 864 -977
rect 870 -978 871 -958
rect 877 -1079 878 -977
rect 912 -978 913 -958
rect 919 -1079 920 -977
rect 954 -978 955 -958
rect 1073 -1079 1074 -977
rect 1094 -978 1095 -958
rect 1248 -1079 1249 -977
rect 75 -1079 76 -979
rect 660 -980 661 -958
rect 667 -980 668 -958
rect 772 -1079 773 -979
rect 849 -980 850 -958
rect 954 -1079 955 -979
rect 961 -980 962 -958
rect 1255 -1079 1256 -979
rect 51 -982 52 -958
rect 660 -1079 661 -981
rect 695 -982 696 -958
rect 1297 -1079 1298 -981
rect 51 -1079 52 -983
rect 884 -984 885 -958
rect 968 -1079 969 -983
rect 1010 -984 1011 -958
rect 1052 -984 1053 -958
rect 1094 -1079 1095 -983
rect 1101 -984 1102 -958
rect 1234 -1079 1235 -983
rect 79 -986 80 -958
rect 450 -986 451 -958
rect 572 -1079 573 -985
rect 870 -1079 871 -985
rect 884 -1079 885 -985
rect 940 -986 941 -958
rect 975 -986 976 -958
rect 1087 -1079 1088 -985
rect 1115 -986 1116 -958
rect 1241 -1079 1242 -985
rect 23 -988 24 -958
rect 450 -1079 451 -987
rect 576 -988 577 -958
rect 912 -1079 913 -987
rect 933 -988 934 -958
rect 1052 -1079 1053 -987
rect 1150 -988 1151 -958
rect 1157 -1079 1158 -987
rect 1164 -988 1165 -958
rect 1318 -1079 1319 -987
rect 23 -1079 24 -989
rect 268 -990 269 -958
rect 282 -990 283 -958
rect 425 -990 426 -958
rect 436 -990 437 -958
rect 695 -1079 696 -989
rect 702 -990 703 -958
rect 933 -1079 934 -989
rect 1003 -990 1004 -958
rect 1115 -1079 1116 -989
rect 1171 -990 1172 -958
rect 1171 -1079 1172 -989
rect 1171 -990 1172 -958
rect 1171 -1079 1172 -989
rect 1185 -990 1186 -958
rect 1339 -1079 1340 -989
rect 79 -1079 80 -991
rect 219 -992 220 -958
rect 254 -992 255 -958
rect 614 -992 615 -958
rect 618 -992 619 -958
rect 688 -1079 689 -991
rect 709 -992 710 -958
rect 1059 -1079 1060 -991
rect 1192 -992 1193 -958
rect 1206 -992 1207 -958
rect 114 -994 115 -958
rect 131 -994 132 -958
rect 149 -1079 150 -993
rect 408 -1079 409 -993
rect 436 -1079 437 -993
rect 576 -1079 577 -993
rect 611 -1079 612 -993
rect 821 -994 822 -958
rect 856 -994 857 -958
rect 1101 -1079 1102 -993
rect 96 -1079 97 -995
rect 114 -1079 115 -995
rect 121 -996 122 -958
rect 121 -1079 122 -995
rect 121 -996 122 -958
rect 121 -1079 122 -995
rect 124 -996 125 -958
rect 653 -996 654 -958
rect 723 -996 724 -958
rect 940 -1079 941 -995
rect 1017 -996 1018 -958
rect 1150 -1079 1151 -995
rect 156 -998 157 -958
rect 156 -1079 157 -997
rect 156 -998 157 -958
rect 156 -1079 157 -997
rect 177 -998 178 -958
rect 254 -1079 255 -997
rect 264 -1079 265 -997
rect 478 -998 479 -958
rect 499 -998 500 -958
rect 856 -1079 857 -997
rect 891 -998 892 -958
rect 975 -1079 976 -997
rect 982 -998 983 -958
rect 1017 -1079 1018 -997
rect 1045 -998 1046 -958
rect 1185 -1079 1186 -997
rect 177 -1079 178 -999
rect 240 -1000 241 -958
rect 268 -1079 269 -999
rect 453 -1000 454 -958
rect 471 -1000 472 -958
rect 982 -1079 983 -999
rect 1066 -1000 1067 -958
rect 1192 -1079 1193 -999
rect 205 -1002 206 -958
rect 212 -1079 213 -1001
rect 219 -1079 220 -1001
rect 1195 -1002 1196 -958
rect 240 -1079 241 -1003
rect 324 -1004 325 -958
rect 331 -1004 332 -958
rect 331 -1079 332 -1003
rect 331 -1004 332 -958
rect 331 -1079 332 -1003
rect 338 -1004 339 -958
rect 387 -1079 388 -1003
rect 471 -1079 472 -1003
rect 506 -1004 507 -958
rect 513 -1004 514 -958
rect 653 -1079 654 -1003
rect 723 -1079 724 -1003
rect 961 -1079 962 -1003
rect 1080 -1004 1081 -958
rect 1206 -1079 1207 -1003
rect 282 -1079 283 -1005
rect 415 -1006 416 -958
rect 478 -1079 479 -1005
rect 1108 -1006 1109 -958
rect 289 -1008 290 -958
rect 324 -1079 325 -1007
rect 341 -1079 342 -1007
rect 401 -1008 402 -958
rect 499 -1079 500 -1007
rect 548 -1079 549 -1007
rect 555 -1008 556 -958
rect 618 -1079 619 -1007
rect 628 -1079 629 -1007
rect 737 -1008 738 -958
rect 747 -1008 748 -958
rect 779 -1008 780 -958
rect 800 -1008 801 -958
rect 821 -1079 822 -1007
rect 835 -1008 836 -958
rect 891 -1079 892 -1007
rect 926 -1008 927 -958
rect 1045 -1079 1046 -1007
rect 1080 -1079 1081 -1007
rect 1129 -1008 1130 -958
rect 128 -1010 129 -958
rect 737 -1079 738 -1009
rect 747 -1079 748 -1009
rect 1227 -1079 1228 -1009
rect 37 -1079 38 -1011
rect 128 -1079 129 -1011
rect 142 -1012 143 -958
rect 289 -1079 290 -1011
rect 303 -1012 304 -958
rect 415 -1079 416 -1011
rect 506 -1079 507 -1011
rect 562 -1012 563 -958
rect 632 -1012 633 -958
rect 1332 -1079 1333 -1011
rect 86 -1014 87 -958
rect 303 -1079 304 -1013
rect 306 -1079 307 -1013
rect 310 -1014 311 -958
rect 317 -1079 318 -1013
rect 481 -1014 482 -958
rect 513 -1079 514 -1013
rect 646 -1014 647 -958
rect 656 -1014 657 -958
rect 800 -1079 801 -1013
rect 814 -1014 815 -958
rect 849 -1079 850 -1013
rect 996 -1014 997 -958
rect 1108 -1079 1109 -1013
rect 86 -1079 87 -1015
rect 544 -1016 545 -958
rect 597 -1016 598 -958
rect 646 -1079 647 -1015
rect 751 -1016 752 -958
rect 779 -1079 780 -1015
rect 807 -1016 808 -958
rect 814 -1079 815 -1015
rect 989 -1016 990 -958
rect 996 -1079 997 -1015
rect 1031 -1016 1032 -958
rect 1129 -1079 1130 -1015
rect 40 -1079 41 -1017
rect 597 -1079 598 -1017
rect 635 -1018 636 -958
rect 1346 -1079 1347 -1017
rect 310 -1079 311 -1019
rect 338 -1079 339 -1019
rect 345 -1020 346 -958
rect 702 -1079 703 -1019
rect 730 -1020 731 -958
rect 751 -1079 752 -1019
rect 758 -1020 759 -958
rect 1003 -1079 1004 -1019
rect 345 -1079 346 -1021
rect 373 -1022 374 -958
rect 376 -1079 377 -1021
rect 1178 -1022 1179 -958
rect 352 -1024 353 -958
rect 530 -1024 531 -958
rect 569 -1024 570 -958
rect 758 -1079 759 -1023
rect 765 -1024 766 -958
rect 1143 -1079 1144 -1023
rect 9 -1079 10 -1025
rect 530 -1079 531 -1025
rect 569 -1079 570 -1025
rect 604 -1026 605 -958
rect 639 -1026 640 -958
rect 681 -1079 682 -1025
rect 793 -1026 794 -958
rect 989 -1079 990 -1025
rect 1024 -1026 1025 -958
rect 1178 -1079 1179 -1025
rect 261 -1028 262 -958
rect 352 -1079 353 -1027
rect 359 -1028 360 -958
rect 667 -1079 668 -1027
rect 677 -1079 678 -1027
rect 765 -1079 766 -1027
rect 793 -1079 794 -1027
rect 824 -1028 825 -958
rect 898 -1028 899 -958
rect 1024 -1079 1025 -1027
rect 68 -1030 69 -958
rect 898 -1079 899 -1029
rect 905 -1030 906 -958
rect 1031 -1079 1032 -1029
rect 107 -1032 108 -958
rect 359 -1079 360 -1031
rect 366 -1032 367 -958
rect 1010 -1079 1011 -1031
rect 107 -1079 108 -1033
rect 625 -1034 626 -958
rect 842 -1034 843 -958
rect 905 -1079 906 -1033
rect 100 -1036 101 -958
rect 842 -1079 843 -1035
rect 100 -1079 101 -1037
rect 1038 -1038 1039 -958
rect 296 -1040 297 -958
rect 639 -1079 640 -1039
rect 947 -1040 948 -958
rect 1038 -1079 1039 -1039
rect 135 -1042 136 -958
rect 296 -1079 297 -1041
rect 366 -1079 367 -1041
rect 1199 -1042 1200 -958
rect 65 -1044 66 -958
rect 135 -1079 136 -1043
rect 369 -1044 370 -958
rect 1283 -1079 1284 -1043
rect 65 -1079 66 -1045
rect 495 -1079 496 -1045
rect 520 -1046 521 -958
rect 1066 -1079 1067 -1045
rect 373 -1079 374 -1047
rect 394 -1048 395 -958
rect 401 -1079 402 -1047
rect 457 -1048 458 -958
rect 464 -1048 465 -958
rect 730 -1079 731 -1047
rect 828 -1048 829 -958
rect 947 -1079 948 -1047
rect 191 -1050 192 -958
rect 394 -1079 395 -1049
rect 429 -1050 430 -958
rect 457 -1079 458 -1049
rect 481 -1079 482 -1049
rect 1199 -1079 1200 -1049
rect 163 -1052 164 -958
rect 191 -1079 192 -1051
rect 261 -1079 262 -1051
rect 464 -1079 465 -1051
rect 492 -1052 493 -958
rect 520 -1079 521 -1051
rect 527 -1052 528 -958
rect 1164 -1079 1165 -1051
rect 163 -1079 164 -1053
rect 926 -1079 927 -1053
rect 184 -1056 185 -958
rect 429 -1079 430 -1055
rect 492 -1079 493 -1055
rect 835 -1079 836 -1055
rect 184 -1079 185 -1057
rect 247 -1058 248 -958
rect 380 -1058 381 -958
rect 541 -1079 542 -1057
rect 583 -1058 584 -958
rect 807 -1079 808 -1057
rect 233 -1060 234 -958
rect 247 -1079 248 -1059
rect 380 -1079 381 -1059
rect 516 -1079 517 -1059
rect 527 -1079 528 -1059
rect 709 -1079 710 -1059
rect 54 -1079 55 -1061
rect 233 -1079 234 -1061
rect 534 -1079 535 -1061
rect 625 -1079 626 -1061
rect 674 -1062 675 -958
rect 828 -1079 829 -1061
rect 443 -1064 444 -958
rect 674 -1079 675 -1063
rect 93 -1066 94 -958
rect 443 -1079 444 -1065
rect 583 -1079 584 -1065
rect 635 -1079 636 -1065
rect 93 -1079 94 -1067
rect 142 -1079 143 -1067
rect 590 -1068 591 -958
rect 604 -1079 605 -1067
rect 226 -1070 227 -958
rect 590 -1079 591 -1069
rect 226 -1079 227 -1071
rect 275 -1072 276 -958
rect 58 -1074 59 -958
rect 275 -1079 276 -1073
rect 58 -1079 59 -1075
rect 72 -1076 73 -958
rect 72 -1079 73 -1077
rect 205 -1079 206 -1077
rect 2 -1204 3 -1088
rect 982 -1089 983 -1087
rect 1241 -1089 1242 -1087
rect 1367 -1204 1368 -1088
rect 1444 -1089 1445 -1087
rect 1451 -1204 1452 -1088
rect 9 -1091 10 -1087
rect 338 -1204 339 -1090
rect 404 -1204 405 -1090
rect 667 -1091 668 -1087
rect 674 -1091 675 -1087
rect 1269 -1091 1270 -1087
rect 1318 -1091 1319 -1087
rect 1353 -1204 1354 -1090
rect 9 -1204 10 -1092
rect 33 -1093 34 -1087
rect 37 -1204 38 -1092
rect 121 -1093 122 -1087
rect 149 -1093 150 -1087
rect 226 -1093 227 -1087
rect 247 -1093 248 -1087
rect 264 -1093 265 -1087
rect 439 -1093 440 -1087
rect 520 -1093 521 -1087
rect 527 -1093 528 -1087
rect 1143 -1093 1144 -1087
rect 1213 -1093 1214 -1087
rect 1241 -1204 1242 -1092
rect 1325 -1093 1326 -1087
rect 1360 -1204 1361 -1092
rect 16 -1095 17 -1087
rect 16 -1204 17 -1094
rect 16 -1095 17 -1087
rect 16 -1204 17 -1094
rect 30 -1204 31 -1094
rect 562 -1095 563 -1087
rect 569 -1095 570 -1087
rect 1318 -1204 1319 -1094
rect 1339 -1095 1340 -1087
rect 1374 -1204 1375 -1094
rect 54 -1097 55 -1087
rect 842 -1097 843 -1087
rect 845 -1204 846 -1096
rect 982 -1204 983 -1096
rect 1220 -1097 1221 -1087
rect 1269 -1204 1270 -1096
rect 1311 -1097 1312 -1087
rect 1339 -1204 1340 -1096
rect 58 -1099 59 -1087
rect 100 -1099 101 -1087
rect 121 -1204 122 -1098
rect 289 -1099 290 -1087
rect 408 -1099 409 -1087
rect 562 -1204 563 -1098
rect 572 -1099 573 -1087
rect 772 -1099 773 -1087
rect 786 -1099 787 -1087
rect 1311 -1204 1312 -1098
rect 58 -1204 59 -1100
rect 177 -1101 178 -1087
rect 212 -1101 213 -1087
rect 523 -1204 524 -1100
rect 530 -1101 531 -1087
rect 618 -1101 619 -1087
rect 628 -1204 629 -1100
rect 1136 -1101 1137 -1087
rect 1192 -1101 1193 -1087
rect 1220 -1204 1221 -1100
rect 75 -1103 76 -1087
rect 1101 -1103 1102 -1087
rect 75 -1204 76 -1104
rect 660 -1105 661 -1087
rect 667 -1204 668 -1104
rect 730 -1105 731 -1087
rect 733 -1204 734 -1104
rect 1136 -1204 1137 -1104
rect 79 -1107 80 -1087
rect 544 -1204 545 -1106
rect 558 -1107 559 -1087
rect 765 -1107 766 -1087
rect 863 -1107 864 -1087
rect 1325 -1204 1326 -1106
rect 79 -1204 80 -1108
rect 443 -1109 444 -1087
rect 471 -1109 472 -1087
rect 635 -1109 636 -1087
rect 653 -1109 654 -1087
rect 674 -1204 675 -1108
rect 684 -1204 685 -1108
rect 1206 -1109 1207 -1087
rect 93 -1111 94 -1087
rect 516 -1111 517 -1087
rect 541 -1111 542 -1087
rect 569 -1204 570 -1110
rect 576 -1111 577 -1087
rect 723 -1111 724 -1087
rect 726 -1111 727 -1087
rect 1150 -1111 1151 -1087
rect 1178 -1111 1179 -1087
rect 1206 -1204 1207 -1110
rect 93 -1204 94 -1112
rect 170 -1113 171 -1087
rect 177 -1204 178 -1112
rect 296 -1113 297 -1087
rect 310 -1113 311 -1087
rect 443 -1204 444 -1112
rect 450 -1113 451 -1087
rect 653 -1204 654 -1112
rect 660 -1204 661 -1112
rect 761 -1204 762 -1112
rect 765 -1204 766 -1112
rect 1234 -1113 1235 -1087
rect 72 -1115 73 -1087
rect 170 -1204 171 -1114
rect 205 -1115 206 -1087
rect 471 -1204 472 -1114
rect 478 -1115 479 -1087
rect 485 -1115 486 -1087
rect 492 -1115 493 -1087
rect 989 -1115 990 -1087
rect 1087 -1115 1088 -1087
rect 1101 -1204 1102 -1114
rect 1150 -1204 1151 -1114
rect 1157 -1115 1158 -1087
rect 44 -1117 45 -1087
rect 478 -1204 479 -1116
rect 499 -1117 500 -1087
rect 877 -1117 878 -1087
rect 929 -1117 930 -1087
rect 1304 -1117 1305 -1087
rect 44 -1204 45 -1118
rect 380 -1119 381 -1087
rect 408 -1204 409 -1118
rect 422 -1119 423 -1087
rect 457 -1119 458 -1087
rect 485 -1204 486 -1118
rect 499 -1204 500 -1118
rect 611 -1119 612 -1087
rect 632 -1119 633 -1087
rect 1248 -1119 1249 -1087
rect 1290 -1119 1291 -1087
rect 1304 -1204 1305 -1118
rect 23 -1121 24 -1087
rect 380 -1204 381 -1120
rect 394 -1121 395 -1087
rect 422 -1204 423 -1120
rect 457 -1204 458 -1120
rect 506 -1121 507 -1087
rect 541 -1204 542 -1120
rect 1297 -1121 1298 -1087
rect 23 -1204 24 -1122
rect 366 -1123 367 -1087
rect 464 -1123 465 -1087
rect 611 -1204 612 -1122
rect 695 -1123 696 -1087
rect 754 -1204 755 -1122
rect 828 -1123 829 -1087
rect 877 -1204 878 -1122
rect 954 -1123 955 -1087
rect 1143 -1204 1144 -1122
rect 1227 -1123 1228 -1087
rect 1248 -1204 1249 -1122
rect 1283 -1123 1284 -1087
rect 1297 -1204 1298 -1122
rect 72 -1204 73 -1124
rect 758 -1125 759 -1087
rect 821 -1125 822 -1087
rect 828 -1204 829 -1124
rect 849 -1125 850 -1087
rect 989 -1204 990 -1124
rect 1045 -1125 1046 -1087
rect 1087 -1204 1088 -1124
rect 1171 -1125 1172 -1087
rect 1283 -1204 1284 -1124
rect 96 -1127 97 -1087
rect 639 -1127 640 -1087
rect 681 -1127 682 -1087
rect 695 -1204 696 -1126
rect 712 -1204 713 -1126
rect 1192 -1204 1193 -1126
rect 1199 -1127 1200 -1087
rect 1227 -1204 1228 -1126
rect 100 -1204 101 -1128
rect 849 -1204 850 -1128
rect 866 -1129 867 -1087
rect 1185 -1129 1186 -1087
rect 117 -1204 118 -1130
rect 1185 -1204 1186 -1130
rect 128 -1133 129 -1087
rect 394 -1204 395 -1132
rect 464 -1204 465 -1132
rect 1276 -1133 1277 -1087
rect 128 -1204 129 -1134
rect 632 -1204 633 -1134
rect 716 -1135 717 -1087
rect 723 -1204 724 -1134
rect 730 -1204 731 -1134
rect 1115 -1135 1116 -1087
rect 1262 -1135 1263 -1087
rect 1276 -1204 1277 -1134
rect 149 -1204 150 -1136
rect 646 -1137 647 -1087
rect 702 -1137 703 -1087
rect 716 -1204 717 -1136
rect 744 -1137 745 -1087
rect 835 -1137 836 -1087
rect 870 -1137 871 -1087
rect 1178 -1204 1179 -1136
rect 163 -1139 164 -1087
rect 205 -1204 206 -1138
rect 212 -1204 213 -1138
rect 677 -1139 678 -1087
rect 688 -1139 689 -1087
rect 702 -1204 703 -1138
rect 744 -1204 745 -1138
rect 1122 -1139 1123 -1087
rect 163 -1204 164 -1140
rect 495 -1141 496 -1087
rect 502 -1141 503 -1087
rect 1066 -1141 1067 -1087
rect 1073 -1141 1074 -1087
rect 1115 -1204 1116 -1140
rect 226 -1204 227 -1142
rect 275 -1143 276 -1087
rect 282 -1143 283 -1087
rect 527 -1204 528 -1142
rect 548 -1143 549 -1087
rect 576 -1204 577 -1142
rect 600 -1204 601 -1142
rect 1255 -1143 1256 -1087
rect 152 -1145 153 -1087
rect 275 -1204 276 -1144
rect 289 -1204 290 -1144
rect 467 -1204 468 -1144
rect 495 -1204 496 -1144
rect 870 -1204 871 -1144
rect 905 -1145 906 -1087
rect 954 -1204 955 -1144
rect 968 -1145 969 -1087
rect 1157 -1204 1158 -1144
rect 1255 -1204 1256 -1144
rect 1332 -1145 1333 -1087
rect 184 -1147 185 -1087
rect 282 -1204 283 -1146
rect 296 -1204 297 -1146
rect 352 -1147 353 -1087
rect 373 -1147 374 -1087
rect 639 -1204 640 -1146
rect 649 -1204 650 -1146
rect 688 -1204 689 -1146
rect 747 -1147 748 -1087
rect 940 -1147 941 -1087
rect 1010 -1147 1011 -1087
rect 1045 -1204 1046 -1146
rect 1066 -1204 1067 -1146
rect 1129 -1147 1130 -1087
rect 103 -1149 104 -1087
rect 373 -1204 374 -1148
rect 506 -1204 507 -1148
rect 796 -1204 797 -1148
rect 800 -1149 801 -1087
rect 821 -1204 822 -1148
rect 856 -1149 857 -1087
rect 905 -1204 906 -1148
rect 933 -1149 934 -1087
rect 1073 -1204 1074 -1148
rect 1080 -1149 1081 -1087
rect 1262 -1204 1263 -1148
rect 5 -1151 6 -1087
rect 856 -1204 857 -1150
rect 891 -1151 892 -1087
rect 940 -1204 941 -1150
rect 961 -1151 962 -1087
rect 1010 -1204 1011 -1150
rect 1017 -1151 1018 -1087
rect 1171 -1204 1172 -1150
rect 5 -1204 6 -1152
rect 1290 -1204 1291 -1152
rect 103 -1204 104 -1154
rect 215 -1204 216 -1154
rect 233 -1155 234 -1087
rect 450 -1204 451 -1154
rect 534 -1155 535 -1087
rect 968 -1204 969 -1154
rect 1017 -1204 1018 -1154
rect 1094 -1155 1095 -1087
rect 1108 -1155 1109 -1087
rect 1332 -1204 1333 -1154
rect 135 -1157 136 -1087
rect 233 -1204 234 -1156
rect 240 -1157 241 -1087
rect 247 -1204 248 -1156
rect 254 -1157 255 -1087
rect 376 -1157 377 -1087
rect 534 -1204 535 -1156
rect 646 -1204 647 -1156
rect 709 -1157 710 -1087
rect 891 -1204 892 -1156
rect 912 -1157 913 -1087
rect 961 -1204 962 -1156
rect 1031 -1157 1032 -1087
rect 1199 -1204 1200 -1156
rect 40 -1159 41 -1087
rect 135 -1204 136 -1158
rect 156 -1159 157 -1087
rect 184 -1204 185 -1158
rect 240 -1204 241 -1158
rect 583 -1159 584 -1087
rect 604 -1159 605 -1087
rect 618 -1204 619 -1158
rect 747 -1204 748 -1158
rect 1080 -1204 1081 -1158
rect 156 -1204 157 -1160
rect 436 -1161 437 -1087
rect 481 -1161 482 -1087
rect 583 -1204 584 -1160
rect 607 -1204 608 -1160
rect 1164 -1161 1165 -1087
rect 261 -1163 262 -1087
rect 786 -1204 787 -1162
rect 814 -1163 815 -1087
rect 933 -1204 934 -1162
rect 1052 -1163 1053 -1087
rect 1094 -1204 1095 -1162
rect 191 -1165 192 -1087
rect 261 -1204 262 -1164
rect 303 -1165 304 -1087
rect 835 -1204 836 -1164
rect 884 -1165 885 -1087
rect 1108 -1204 1109 -1164
rect 142 -1167 143 -1087
rect 191 -1204 192 -1166
rect 219 -1167 220 -1087
rect 303 -1204 304 -1166
rect 310 -1204 311 -1166
rect 597 -1167 598 -1087
rect 751 -1167 752 -1087
rect 800 -1204 801 -1166
rect 807 -1167 808 -1087
rect 884 -1204 885 -1166
rect 919 -1167 920 -1087
rect 1031 -1204 1032 -1166
rect 1059 -1167 1060 -1087
rect 1129 -1204 1130 -1166
rect 107 -1169 108 -1087
rect 142 -1204 143 -1168
rect 219 -1204 220 -1168
rect 555 -1169 556 -1087
rect 558 -1204 559 -1168
rect 1122 -1204 1123 -1168
rect 107 -1204 108 -1170
rect 198 -1171 199 -1087
rect 317 -1171 318 -1087
rect 366 -1204 367 -1170
rect 401 -1171 402 -1087
rect 436 -1204 437 -1170
rect 513 -1171 514 -1087
rect 1052 -1204 1053 -1170
rect 180 -1204 181 -1172
rect 513 -1204 514 -1172
rect 530 -1204 531 -1172
rect 1164 -1204 1165 -1172
rect 198 -1204 199 -1174
rect 268 -1175 269 -1087
rect 317 -1204 318 -1174
rect 324 -1175 325 -1087
rect 341 -1175 342 -1087
rect 352 -1204 353 -1174
rect 359 -1175 360 -1087
rect 807 -1204 808 -1174
rect 1024 -1175 1025 -1087
rect 1059 -1204 1060 -1174
rect 254 -1204 255 -1176
rect 401 -1204 402 -1176
rect 555 -1204 556 -1176
rect 1213 -1204 1214 -1176
rect 268 -1204 269 -1178
rect 429 -1179 430 -1087
rect 565 -1179 566 -1087
rect 772 -1204 773 -1178
rect 779 -1179 780 -1087
rect 912 -1204 913 -1178
rect 975 -1179 976 -1087
rect 1024 -1204 1025 -1178
rect 324 -1204 325 -1180
rect 345 -1181 346 -1087
rect 359 -1204 360 -1180
rect 681 -1204 682 -1180
rect 751 -1204 752 -1180
rect 926 -1204 927 -1180
rect 975 -1204 976 -1180
rect 1038 -1181 1039 -1087
rect 331 -1183 332 -1087
rect 779 -1204 780 -1182
rect 793 -1183 794 -1087
rect 814 -1204 815 -1182
rect 1003 -1183 1004 -1087
rect 1038 -1204 1039 -1182
rect 331 -1204 332 -1184
rect 415 -1185 416 -1087
rect 429 -1204 430 -1184
rect 635 -1204 636 -1184
rect 758 -1204 759 -1184
rect 1346 -1185 1347 -1087
rect 51 -1187 52 -1087
rect 1346 -1204 1347 -1186
rect 345 -1204 346 -1188
rect 737 -1189 738 -1087
rect 793 -1204 794 -1188
rect 863 -1204 864 -1188
rect 996 -1189 997 -1087
rect 1003 -1204 1004 -1188
rect 65 -1191 66 -1087
rect 737 -1204 738 -1190
rect 947 -1191 948 -1087
rect 996 -1204 997 -1190
rect 65 -1204 66 -1192
rect 86 -1193 87 -1087
rect 387 -1193 388 -1087
rect 415 -1204 416 -1192
rect 597 -1204 598 -1192
rect 1234 -1204 1235 -1192
rect 86 -1204 87 -1194
rect 114 -1195 115 -1087
rect 387 -1204 388 -1194
rect 492 -1204 493 -1194
rect 625 -1195 626 -1087
rect 919 -1204 920 -1194
rect 51 -1204 52 -1196
rect 625 -1204 626 -1196
rect 898 -1197 899 -1087
rect 947 -1204 948 -1196
rect 114 -1204 115 -1198
rect 590 -1199 591 -1087
rect 551 -1204 552 -1200
rect 898 -1204 899 -1200
rect 590 -1204 591 -1202
rect 709 -1204 710 -1202
rect 2 -1325 3 -1213
rect 303 -1214 304 -1212
rect 366 -1214 367 -1212
rect 558 -1214 559 -1212
rect 607 -1214 608 -1212
rect 968 -1214 969 -1212
rect 982 -1214 983 -1212
rect 982 -1325 983 -1213
rect 982 -1214 983 -1212
rect 982 -1325 983 -1213
rect 1017 -1214 1018 -1212
rect 1020 -1220 1021 -1213
rect 1269 -1214 1270 -1212
rect 1272 -1214 1273 -1212
rect 1304 -1214 1305 -1212
rect 1304 -1325 1305 -1213
rect 1304 -1214 1305 -1212
rect 1304 -1325 1305 -1213
rect 1360 -1214 1361 -1212
rect 1381 -1325 1382 -1213
rect 1451 -1214 1452 -1212
rect 1458 -1325 1459 -1213
rect 5 -1216 6 -1212
rect 779 -1216 780 -1212
rect 793 -1325 794 -1215
rect 849 -1216 850 -1212
rect 870 -1216 871 -1212
rect 968 -1325 969 -1215
rect 1017 -1325 1018 -1215
rect 1269 -1325 1270 -1215
rect 1283 -1216 1284 -1212
rect 30 -1218 31 -1212
rect 551 -1218 552 -1212
rect 614 -1325 615 -1217
rect 618 -1218 619 -1212
rect 628 -1218 629 -1212
rect 695 -1218 696 -1212
rect 698 -1325 699 -1217
rect 1073 -1218 1074 -1212
rect 1283 -1325 1284 -1217
rect 1318 -1218 1319 -1212
rect 30 -1325 31 -1219
rect 562 -1220 563 -1212
rect 632 -1220 633 -1212
rect 1143 -1220 1144 -1212
rect 1272 -1325 1273 -1219
rect 1318 -1325 1319 -1219
rect 37 -1222 38 -1212
rect 212 -1222 213 -1212
rect 261 -1222 262 -1212
rect 261 -1325 262 -1221
rect 261 -1222 262 -1212
rect 261 -1325 262 -1221
rect 289 -1222 290 -1212
rect 562 -1325 563 -1221
rect 646 -1222 647 -1212
rect 1374 -1222 1375 -1212
rect 37 -1325 38 -1223
rect 58 -1224 59 -1212
rect 72 -1325 73 -1223
rect 121 -1224 122 -1212
rect 124 -1325 125 -1223
rect 352 -1224 353 -1212
rect 366 -1325 367 -1223
rect 635 -1325 636 -1223
rect 653 -1224 654 -1212
rect 1388 -1325 1389 -1223
rect 44 -1226 45 -1212
rect 649 -1226 650 -1212
rect 653 -1325 654 -1225
rect 716 -1226 717 -1212
rect 719 -1325 720 -1225
rect 1143 -1325 1144 -1225
rect 44 -1325 45 -1227
rect 93 -1228 94 -1212
rect 100 -1325 101 -1227
rect 117 -1228 118 -1212
rect 121 -1325 122 -1227
rect 555 -1228 556 -1212
rect 600 -1228 601 -1212
rect 646 -1325 647 -1227
rect 667 -1228 668 -1212
rect 667 -1325 668 -1227
rect 667 -1228 668 -1212
rect 667 -1325 668 -1227
rect 684 -1325 685 -1227
rect 1297 -1228 1298 -1212
rect 51 -1230 52 -1212
rect 93 -1325 94 -1229
rect 138 -1325 139 -1229
rect 569 -1230 570 -1212
rect 709 -1230 710 -1212
rect 737 -1230 738 -1212
rect 751 -1230 752 -1212
rect 1374 -1325 1375 -1229
rect 51 -1325 52 -1231
rect 418 -1325 419 -1231
rect 432 -1325 433 -1231
rect 534 -1232 535 -1212
rect 544 -1232 545 -1212
rect 1360 -1325 1361 -1231
rect 58 -1325 59 -1233
rect 478 -1234 479 -1212
rect 492 -1234 493 -1212
rect 884 -1234 885 -1212
rect 915 -1325 916 -1233
rect 1080 -1234 1081 -1212
rect 1150 -1234 1151 -1212
rect 1297 -1325 1298 -1233
rect 75 -1236 76 -1212
rect 422 -1236 423 -1212
rect 436 -1236 437 -1212
rect 464 -1236 465 -1212
rect 520 -1236 521 -1212
rect 709 -1325 710 -1235
rect 712 -1236 713 -1212
rect 1094 -1236 1095 -1212
rect 1150 -1325 1151 -1235
rect 1157 -1236 1158 -1212
rect 89 -1325 90 -1237
rect 226 -1238 227 -1212
rect 289 -1325 290 -1237
rect 373 -1238 374 -1212
rect 394 -1238 395 -1212
rect 530 -1238 531 -1212
rect 534 -1325 535 -1237
rect 705 -1325 706 -1237
rect 754 -1238 755 -1212
rect 1339 -1238 1340 -1212
rect 142 -1240 143 -1212
rect 142 -1325 143 -1239
rect 142 -1240 143 -1212
rect 142 -1325 143 -1239
rect 149 -1240 150 -1212
rect 597 -1240 598 -1212
rect 604 -1240 605 -1212
rect 884 -1325 885 -1239
rect 940 -1240 941 -1212
rect 940 -1325 941 -1239
rect 940 -1240 941 -1212
rect 940 -1325 941 -1239
rect 1010 -1240 1011 -1212
rect 1073 -1325 1074 -1239
rect 1080 -1325 1081 -1239
rect 1108 -1240 1109 -1212
rect 1157 -1325 1158 -1239
rect 1171 -1240 1172 -1212
rect 149 -1325 150 -1241
rect 345 -1242 346 -1212
rect 352 -1325 353 -1241
rect 387 -1242 388 -1212
rect 436 -1325 437 -1241
rect 541 -1242 542 -1212
rect 548 -1242 549 -1212
rect 996 -1242 997 -1212
rect 1010 -1325 1011 -1241
rect 1038 -1242 1039 -1212
rect 1094 -1325 1095 -1241
rect 1178 -1242 1179 -1212
rect 163 -1244 164 -1212
rect 163 -1325 164 -1243
rect 163 -1244 164 -1212
rect 163 -1325 164 -1243
rect 173 -1325 174 -1243
rect 1199 -1244 1200 -1212
rect 177 -1325 178 -1245
rect 254 -1246 255 -1212
rect 282 -1246 283 -1212
rect 387 -1325 388 -1245
rect 446 -1325 447 -1245
rect 1199 -1325 1200 -1245
rect 191 -1248 192 -1212
rect 303 -1325 304 -1247
rect 310 -1248 311 -1212
rect 618 -1325 619 -1247
rect 660 -1248 661 -1212
rect 751 -1325 752 -1247
rect 765 -1248 766 -1212
rect 1024 -1248 1025 -1212
rect 1038 -1325 1039 -1247
rect 1045 -1248 1046 -1212
rect 1129 -1248 1130 -1212
rect 1171 -1325 1172 -1247
rect 1178 -1325 1179 -1247
rect 1192 -1248 1193 -1212
rect 170 -1250 171 -1212
rect 191 -1325 192 -1249
rect 198 -1250 199 -1212
rect 681 -1250 682 -1212
rect 695 -1325 696 -1249
rect 737 -1325 738 -1249
rect 758 -1250 759 -1212
rect 1045 -1325 1046 -1249
rect 1164 -1250 1165 -1212
rect 1339 -1325 1340 -1249
rect 198 -1325 199 -1251
rect 296 -1252 297 -1212
rect 310 -1325 311 -1251
rect 495 -1252 496 -1212
rect 520 -1325 521 -1251
rect 572 -1325 573 -1251
rect 604 -1325 605 -1251
rect 611 -1252 612 -1212
rect 660 -1325 661 -1251
rect 702 -1252 703 -1212
rect 758 -1325 759 -1251
rect 786 -1252 787 -1212
rect 796 -1252 797 -1212
rect 1206 -1252 1207 -1212
rect 205 -1254 206 -1212
rect 394 -1325 395 -1253
rect 450 -1254 451 -1212
rect 492 -1325 493 -1253
rect 527 -1254 528 -1212
rect 1234 -1254 1235 -1212
rect 135 -1256 136 -1212
rect 205 -1325 206 -1255
rect 212 -1325 213 -1255
rect 317 -1256 318 -1212
rect 331 -1256 332 -1212
rect 422 -1325 423 -1255
rect 464 -1325 465 -1255
rect 471 -1256 472 -1212
rect 527 -1325 528 -1255
rect 544 -1325 545 -1255
rect 548 -1325 549 -1255
rect 733 -1256 734 -1212
rect 765 -1325 766 -1255
rect 807 -1256 808 -1212
rect 842 -1256 843 -1212
rect 1262 -1256 1263 -1212
rect 135 -1325 136 -1257
rect 1220 -1258 1221 -1212
rect 1234 -1325 1235 -1257
rect 1248 -1258 1249 -1212
rect 219 -1260 220 -1212
rect 597 -1325 598 -1259
rect 621 -1325 622 -1259
rect 1248 -1325 1249 -1259
rect 156 -1262 157 -1212
rect 219 -1325 220 -1261
rect 226 -1325 227 -1261
rect 467 -1262 468 -1212
rect 555 -1325 556 -1261
rect 576 -1262 577 -1212
rect 681 -1325 682 -1261
rect 1367 -1262 1368 -1212
rect 103 -1264 104 -1212
rect 156 -1325 157 -1263
rect 233 -1264 234 -1212
rect 282 -1325 283 -1263
rect 296 -1325 297 -1263
rect 408 -1264 409 -1212
rect 457 -1264 458 -1212
rect 471 -1325 472 -1263
rect 569 -1325 570 -1263
rect 1332 -1264 1333 -1212
rect 1353 -1264 1354 -1212
rect 1367 -1325 1368 -1263
rect 16 -1266 17 -1212
rect 457 -1325 458 -1265
rect 576 -1325 577 -1265
rect 590 -1266 591 -1212
rect 779 -1325 780 -1265
rect 800 -1266 801 -1212
rect 807 -1325 808 -1265
rect 821 -1266 822 -1212
rect 828 -1266 829 -1212
rect 842 -1325 843 -1265
rect 845 -1266 846 -1212
rect 954 -1266 955 -1212
rect 989 -1266 990 -1212
rect 996 -1325 997 -1265
rect 1003 -1266 1004 -1212
rect 1129 -1325 1130 -1265
rect 1164 -1325 1165 -1265
rect 1185 -1266 1186 -1212
rect 1332 -1325 1333 -1265
rect 1346 -1266 1347 -1212
rect 16 -1325 17 -1267
rect 639 -1268 640 -1212
rect 786 -1325 787 -1267
rect 835 -1268 836 -1212
rect 849 -1325 850 -1267
rect 891 -1268 892 -1212
rect 961 -1268 962 -1212
rect 989 -1325 990 -1267
rect 1003 -1325 1004 -1267
rect 1031 -1268 1032 -1212
rect 1066 -1268 1067 -1212
rect 1206 -1325 1207 -1267
rect 1255 -1268 1256 -1212
rect 1346 -1325 1347 -1267
rect 61 -1325 62 -1269
rect 1353 -1325 1354 -1269
rect 170 -1325 171 -1271
rect 1066 -1325 1067 -1271
rect 1087 -1272 1088 -1212
rect 1220 -1325 1221 -1271
rect 1255 -1325 1256 -1271
rect 1276 -1272 1277 -1212
rect 233 -1325 234 -1273
rect 506 -1274 507 -1212
rect 625 -1274 626 -1212
rect 835 -1325 836 -1273
rect 866 -1325 867 -1273
rect 1262 -1325 1263 -1273
rect 1276 -1325 1277 -1273
rect 1290 -1274 1291 -1212
rect 240 -1276 241 -1212
rect 450 -1325 451 -1275
rect 485 -1276 486 -1212
rect 506 -1325 507 -1275
rect 583 -1276 584 -1212
rect 625 -1325 626 -1275
rect 639 -1325 640 -1275
rect 674 -1276 675 -1212
rect 800 -1325 801 -1275
rect 898 -1276 899 -1212
rect 933 -1276 934 -1212
rect 961 -1325 962 -1275
rect 975 -1276 976 -1212
rect 1031 -1325 1032 -1275
rect 1087 -1325 1088 -1275
rect 1101 -1276 1102 -1212
rect 1122 -1276 1123 -1212
rect 1185 -1325 1186 -1275
rect 1290 -1325 1291 -1275
rect 1325 -1276 1326 -1212
rect 68 -1325 69 -1277
rect 1122 -1325 1123 -1277
rect 1311 -1278 1312 -1212
rect 1325 -1325 1326 -1277
rect 114 -1280 115 -1212
rect 1101 -1325 1102 -1279
rect 65 -1282 66 -1212
rect 114 -1325 115 -1281
rect 240 -1325 241 -1281
rect 632 -1325 633 -1281
rect 744 -1282 745 -1212
rect 933 -1325 934 -1281
rect 1024 -1325 1025 -1281
rect 1052 -1282 1053 -1212
rect 247 -1284 248 -1212
rect 317 -1325 318 -1283
rect 324 -1284 325 -1212
rect 485 -1325 486 -1283
rect 499 -1284 500 -1212
rect 674 -1325 675 -1283
rect 730 -1284 731 -1212
rect 1052 -1325 1053 -1283
rect 79 -1286 80 -1212
rect 499 -1325 500 -1285
rect 583 -1325 584 -1285
rect 768 -1286 769 -1212
rect 821 -1325 822 -1285
rect 856 -1286 857 -1212
rect 870 -1325 871 -1285
rect 947 -1286 948 -1212
rect 79 -1325 80 -1287
rect 254 -1325 255 -1287
rect 331 -1325 332 -1287
rect 429 -1288 430 -1212
rect 443 -1288 444 -1212
rect 590 -1325 591 -1287
rect 730 -1325 731 -1287
rect 1059 -1288 1060 -1212
rect 107 -1290 108 -1212
rect 443 -1325 444 -1289
rect 513 -1290 514 -1212
rect 947 -1325 948 -1289
rect 1059 -1325 1060 -1289
rect 1227 -1290 1228 -1212
rect 86 -1292 87 -1212
rect 107 -1325 108 -1291
rect 184 -1292 185 -1212
rect 324 -1325 325 -1291
rect 338 -1292 339 -1212
rect 478 -1325 479 -1291
rect 513 -1325 514 -1291
rect 688 -1292 689 -1212
rect 744 -1325 745 -1291
rect 817 -1325 818 -1291
rect 828 -1325 829 -1291
rect 926 -1292 927 -1212
rect 1213 -1292 1214 -1212
rect 1227 -1325 1228 -1291
rect 86 -1325 87 -1293
rect 1108 -1325 1109 -1293
rect 1213 -1325 1214 -1293
rect 1241 -1294 1242 -1212
rect 184 -1325 185 -1295
rect 733 -1325 734 -1295
rect 747 -1296 748 -1212
rect 975 -1325 976 -1295
rect 247 -1325 248 -1297
rect 611 -1325 612 -1297
rect 688 -1325 689 -1297
rect 723 -1298 724 -1212
rect 856 -1325 857 -1297
rect 863 -1298 864 -1212
rect 877 -1298 878 -1212
rect 877 -1325 878 -1297
rect 877 -1298 878 -1212
rect 877 -1325 878 -1297
rect 891 -1325 892 -1297
rect 905 -1298 906 -1212
rect 338 -1325 339 -1299
rect 401 -1300 402 -1212
rect 523 -1300 524 -1212
rect 1241 -1325 1242 -1299
rect 9 -1302 10 -1212
rect 401 -1325 402 -1301
rect 702 -1325 703 -1301
rect 926 -1325 927 -1301
rect 9 -1325 10 -1303
rect 772 -1304 773 -1212
rect 863 -1325 864 -1303
rect 1311 -1325 1312 -1303
rect 345 -1325 346 -1305
rect 415 -1306 416 -1212
rect 772 -1325 773 -1305
rect 814 -1306 815 -1212
rect 898 -1325 899 -1305
rect 954 -1325 955 -1305
rect 268 -1308 269 -1212
rect 415 -1325 416 -1307
rect 814 -1325 815 -1307
rect 1136 -1308 1137 -1212
rect 268 -1325 269 -1309
rect 359 -1310 360 -1212
rect 369 -1325 370 -1309
rect 1192 -1325 1193 -1309
rect 359 -1325 360 -1311
rect 541 -1325 542 -1311
rect 905 -1325 906 -1311
rect 919 -1312 920 -1212
rect 376 -1325 377 -1313
rect 723 -1325 724 -1313
rect 912 -1314 913 -1212
rect 919 -1325 920 -1313
rect 380 -1316 381 -1212
rect 408 -1325 409 -1315
rect 761 -1316 762 -1212
rect 912 -1325 913 -1315
rect 23 -1318 24 -1212
rect 380 -1325 381 -1317
rect 404 -1318 405 -1212
rect 1136 -1325 1137 -1317
rect 23 -1325 24 -1319
rect 128 -1320 129 -1212
rect 128 -1325 129 -1321
rect 275 -1322 276 -1212
rect 275 -1325 276 -1323
rect 390 -1325 391 -1323
rect 9 -1335 10 -1333
rect 9 -1450 10 -1334
rect 9 -1335 10 -1333
rect 9 -1450 10 -1334
rect 33 -1450 34 -1334
rect 107 -1335 108 -1333
rect 121 -1335 122 -1333
rect 1353 -1335 1354 -1333
rect 1423 -1450 1424 -1334
rect 1451 -1450 1452 -1334
rect 1458 -1335 1459 -1333
rect 1465 -1450 1466 -1334
rect 44 -1337 45 -1333
rect 373 -1337 374 -1333
rect 387 -1337 388 -1333
rect 1066 -1337 1067 -1333
rect 1122 -1337 1123 -1333
rect 1402 -1450 1403 -1336
rect 44 -1450 45 -1338
rect 751 -1339 752 -1333
rect 814 -1339 815 -1333
rect 1227 -1339 1228 -1333
rect 1255 -1339 1256 -1333
rect 1353 -1450 1354 -1338
rect 1360 -1339 1361 -1333
rect 1458 -1450 1459 -1338
rect 65 -1341 66 -1333
rect 555 -1341 556 -1333
rect 583 -1341 584 -1333
rect 618 -1450 619 -1340
rect 635 -1341 636 -1333
rect 877 -1341 878 -1333
rect 887 -1450 888 -1340
rect 1374 -1341 1375 -1333
rect 65 -1450 66 -1342
rect 124 -1343 125 -1333
rect 135 -1343 136 -1333
rect 1430 -1450 1431 -1342
rect 61 -1345 62 -1333
rect 135 -1450 136 -1344
rect 163 -1345 164 -1333
rect 782 -1450 783 -1344
rect 793 -1345 794 -1333
rect 877 -1450 878 -1344
rect 898 -1345 899 -1333
rect 1073 -1345 1074 -1333
rect 1129 -1345 1130 -1333
rect 1409 -1450 1410 -1344
rect 68 -1347 69 -1333
rect 446 -1347 447 -1333
rect 464 -1347 465 -1333
rect 569 -1347 570 -1333
rect 614 -1347 615 -1333
rect 1080 -1347 1081 -1333
rect 1136 -1347 1137 -1333
rect 1136 -1450 1137 -1346
rect 1136 -1347 1137 -1333
rect 1136 -1450 1137 -1346
rect 1150 -1347 1151 -1333
rect 1227 -1450 1228 -1346
rect 1262 -1347 1263 -1333
rect 1360 -1450 1361 -1346
rect 30 -1349 31 -1333
rect 569 -1450 570 -1348
rect 646 -1349 647 -1333
rect 817 -1450 818 -1348
rect 821 -1349 822 -1333
rect 898 -1450 899 -1348
rect 912 -1349 913 -1333
rect 1367 -1349 1368 -1333
rect 79 -1351 80 -1333
rect 324 -1351 325 -1333
rect 380 -1351 381 -1333
rect 446 -1450 447 -1350
rect 478 -1351 479 -1333
rect 478 -1450 479 -1350
rect 478 -1351 479 -1333
rect 478 -1450 479 -1350
rect 509 -1450 510 -1350
rect 1304 -1351 1305 -1333
rect 1332 -1351 1333 -1333
rect 1437 -1450 1438 -1350
rect 82 -1353 83 -1333
rect 1220 -1353 1221 -1333
rect 1234 -1353 1235 -1333
rect 1332 -1450 1333 -1352
rect 1339 -1353 1340 -1333
rect 1374 -1450 1375 -1352
rect 82 -1450 83 -1354
rect 747 -1450 748 -1354
rect 821 -1450 822 -1354
rect 1248 -1355 1249 -1333
rect 1269 -1355 1270 -1333
rect 1367 -1450 1368 -1354
rect 86 -1357 87 -1333
rect 100 -1357 101 -1333
rect 107 -1450 108 -1356
rect 366 -1357 367 -1333
rect 380 -1450 381 -1356
rect 684 -1357 685 -1333
rect 695 -1357 696 -1333
rect 723 -1357 724 -1333
rect 852 -1450 853 -1356
rect 1052 -1357 1053 -1333
rect 1094 -1357 1095 -1333
rect 1248 -1450 1249 -1356
rect 1297 -1357 1298 -1333
rect 1416 -1450 1417 -1356
rect 86 -1450 87 -1358
rect 219 -1359 220 -1333
rect 254 -1359 255 -1333
rect 366 -1450 367 -1358
rect 376 -1359 377 -1333
rect 1052 -1450 1053 -1358
rect 1059 -1359 1060 -1333
rect 1297 -1450 1298 -1358
rect 1318 -1359 1319 -1333
rect 1339 -1450 1340 -1358
rect 1346 -1359 1347 -1333
rect 1444 -1450 1445 -1358
rect 100 -1450 101 -1360
rect 296 -1361 297 -1333
rect 317 -1361 318 -1333
rect 373 -1450 374 -1360
rect 415 -1361 416 -1333
rect 1311 -1361 1312 -1333
rect 23 -1363 24 -1333
rect 296 -1450 297 -1362
rect 324 -1450 325 -1362
rect 331 -1363 332 -1333
rect 418 -1363 419 -1333
rect 856 -1363 857 -1333
rect 866 -1363 867 -1333
rect 968 -1363 969 -1333
rect 982 -1363 983 -1333
rect 1066 -1450 1067 -1362
rect 1157 -1363 1158 -1333
rect 1220 -1450 1221 -1362
rect 1241 -1363 1242 -1333
rect 1346 -1450 1347 -1362
rect 23 -1450 24 -1364
rect 247 -1365 248 -1333
rect 429 -1365 430 -1333
rect 859 -1450 860 -1364
rect 968 -1450 969 -1364
rect 975 -1365 976 -1333
rect 996 -1365 997 -1333
rect 1073 -1450 1074 -1364
rect 1164 -1365 1165 -1333
rect 1234 -1450 1235 -1364
rect 37 -1367 38 -1333
rect 317 -1450 318 -1366
rect 429 -1450 430 -1366
rect 572 -1367 573 -1333
rect 583 -1450 584 -1366
rect 646 -1450 647 -1366
rect 649 -1450 650 -1366
rect 1038 -1367 1039 -1333
rect 1045 -1367 1046 -1333
rect 1048 -1389 1049 -1366
rect 1164 -1450 1165 -1366
rect 1171 -1367 1172 -1333
rect 1178 -1367 1179 -1333
rect 1262 -1450 1263 -1366
rect 37 -1450 38 -1368
rect 534 -1369 535 -1333
rect 541 -1369 542 -1333
rect 947 -1369 948 -1333
rect 954 -1369 955 -1333
rect 1038 -1450 1039 -1368
rect 1045 -1450 1046 -1368
rect 1388 -1369 1389 -1333
rect 93 -1371 94 -1333
rect 331 -1450 332 -1370
rect 436 -1371 437 -1333
rect 695 -1450 696 -1370
rect 698 -1371 699 -1333
rect 954 -1450 955 -1370
rect 1017 -1371 1018 -1333
rect 1129 -1450 1130 -1370
rect 1192 -1371 1193 -1333
rect 1255 -1450 1256 -1370
rect 1276 -1371 1277 -1333
rect 1388 -1450 1389 -1370
rect 93 -1450 94 -1372
rect 460 -1450 461 -1372
rect 534 -1450 535 -1372
rect 555 -1450 556 -1372
rect 632 -1373 633 -1333
rect 1311 -1450 1312 -1372
rect 121 -1450 122 -1374
rect 149 -1375 150 -1333
rect 152 -1450 153 -1374
rect 415 -1450 416 -1374
rect 436 -1450 437 -1374
rect 457 -1375 458 -1333
rect 541 -1450 542 -1374
rect 786 -1375 787 -1333
rect 793 -1450 794 -1374
rect 982 -1450 983 -1374
rect 1024 -1375 1025 -1333
rect 1094 -1450 1095 -1374
rect 1101 -1375 1102 -1333
rect 1171 -1450 1172 -1374
rect 1192 -1450 1193 -1374
rect 1283 -1375 1284 -1333
rect 128 -1377 129 -1333
rect 254 -1450 255 -1376
rect 443 -1377 444 -1333
rect 1157 -1450 1158 -1376
rect 1199 -1377 1200 -1333
rect 1283 -1450 1284 -1376
rect 128 -1450 129 -1378
rect 310 -1379 311 -1333
rect 457 -1450 458 -1378
rect 1318 -1450 1319 -1378
rect 131 -1450 132 -1380
rect 1269 -1450 1270 -1380
rect 149 -1450 150 -1382
rect 590 -1383 591 -1333
rect 632 -1450 633 -1382
rect 856 -1450 857 -1382
rect 870 -1383 871 -1333
rect 1024 -1450 1025 -1382
rect 1031 -1383 1032 -1333
rect 1122 -1450 1123 -1382
rect 1199 -1450 1200 -1382
rect 1290 -1383 1291 -1333
rect 163 -1450 164 -1384
rect 411 -1450 412 -1384
rect 527 -1385 528 -1333
rect 870 -1450 871 -1384
rect 884 -1385 885 -1333
rect 947 -1450 948 -1384
rect 1010 -1385 1011 -1333
rect 1101 -1450 1102 -1384
rect 1206 -1385 1207 -1333
rect 1276 -1450 1277 -1384
rect 170 -1387 171 -1333
rect 912 -1450 913 -1386
rect 933 -1387 934 -1333
rect 996 -1450 997 -1386
rect 1143 -1387 1144 -1333
rect 1206 -1450 1207 -1386
rect 170 -1450 171 -1388
rect 681 -1389 682 -1333
rect 702 -1389 703 -1333
rect 989 -1389 990 -1333
rect 1143 -1450 1144 -1388
rect 198 -1391 199 -1333
rect 397 -1450 398 -1390
rect 513 -1391 514 -1333
rect 681 -1450 682 -1390
rect 705 -1391 706 -1333
rect 961 -1391 962 -1333
rect 184 -1393 185 -1333
rect 198 -1450 199 -1392
rect 205 -1393 206 -1333
rect 205 -1450 206 -1392
rect 205 -1393 206 -1333
rect 205 -1450 206 -1392
rect 212 -1393 213 -1333
rect 369 -1393 370 -1333
rect 394 -1393 395 -1333
rect 527 -1450 528 -1392
rect 544 -1393 545 -1333
rect 660 -1393 661 -1333
rect 667 -1393 668 -1333
rect 751 -1450 752 -1392
rect 758 -1393 759 -1333
rect 786 -1450 787 -1392
rect 814 -1450 815 -1392
rect 1290 -1450 1291 -1392
rect 184 -1450 185 -1394
rect 240 -1395 241 -1333
rect 247 -1450 248 -1394
rect 565 -1450 566 -1394
rect 590 -1450 591 -1394
rect 653 -1395 654 -1333
rect 667 -1450 668 -1394
rect 800 -1395 801 -1333
rect 828 -1395 829 -1333
rect 1010 -1450 1011 -1394
rect 191 -1397 192 -1333
rect 212 -1450 213 -1396
rect 219 -1450 220 -1396
rect 320 -1450 321 -1396
rect 401 -1397 402 -1333
rect 513 -1450 514 -1396
rect 551 -1450 552 -1396
rect 1080 -1450 1081 -1396
rect 2 -1399 3 -1333
rect 191 -1450 192 -1398
rect 240 -1450 241 -1398
rect 485 -1399 486 -1333
rect 492 -1399 493 -1333
rect 653 -1450 654 -1398
rect 716 -1399 717 -1333
rect 779 -1399 780 -1333
rect 831 -1450 832 -1398
rect 1178 -1450 1179 -1398
rect 2 -1450 3 -1400
rect 51 -1401 52 -1333
rect 275 -1401 276 -1333
rect 800 -1450 801 -1400
rect 842 -1401 843 -1333
rect 933 -1450 934 -1400
rect 940 -1401 941 -1333
rect 1017 -1450 1018 -1400
rect 51 -1450 52 -1402
rect 261 -1403 262 -1333
rect 275 -1450 276 -1402
rect 548 -1403 549 -1333
rect 625 -1403 626 -1333
rect 702 -1450 703 -1402
rect 716 -1450 717 -1402
rect 744 -1403 745 -1333
rect 758 -1450 759 -1402
rect 772 -1403 773 -1333
rect 779 -1450 780 -1402
rect 1150 -1450 1151 -1402
rect 79 -1450 80 -1404
rect 261 -1450 262 -1404
rect 303 -1405 304 -1333
rect 394 -1450 395 -1404
rect 450 -1405 451 -1333
rect 485 -1450 486 -1404
rect 492 -1450 493 -1404
rect 520 -1405 521 -1333
rect 548 -1450 549 -1404
rect 1325 -1405 1326 -1333
rect 89 -1407 90 -1333
rect 940 -1450 941 -1406
rect 1213 -1407 1214 -1333
rect 1325 -1450 1326 -1406
rect 138 -1409 139 -1333
rect 842 -1450 843 -1408
rect 866 -1450 867 -1408
rect 1031 -1450 1032 -1408
rect 1185 -1409 1186 -1333
rect 1213 -1450 1214 -1408
rect 282 -1411 283 -1333
rect 450 -1450 451 -1410
rect 464 -1450 465 -1410
rect 744 -1450 745 -1410
rect 891 -1411 892 -1333
rect 961 -1450 962 -1410
rect 1115 -1411 1116 -1333
rect 1185 -1450 1186 -1410
rect 282 -1450 283 -1412
rect 289 -1413 290 -1333
rect 303 -1450 304 -1412
rect 352 -1413 353 -1333
rect 520 -1450 521 -1412
rect 1395 -1450 1396 -1412
rect 289 -1450 290 -1414
rect 765 -1415 766 -1333
rect 796 -1450 797 -1414
rect 1115 -1450 1116 -1414
rect 310 -1450 311 -1416
rect 726 -1450 727 -1416
rect 730 -1417 731 -1333
rect 1059 -1450 1060 -1416
rect 352 -1450 353 -1418
rect 359 -1419 360 -1333
rect 562 -1419 563 -1333
rect 765 -1450 766 -1418
rect 905 -1419 906 -1333
rect 975 -1450 976 -1418
rect 338 -1421 339 -1333
rect 562 -1450 563 -1420
rect 597 -1421 598 -1333
rect 625 -1450 626 -1420
rect 639 -1421 640 -1333
rect 660 -1450 661 -1420
rect 688 -1421 689 -1333
rect 730 -1450 731 -1420
rect 737 -1421 738 -1333
rect 772 -1450 773 -1420
rect 905 -1450 906 -1420
rect 1108 -1421 1109 -1333
rect 166 -1423 167 -1333
rect 597 -1450 598 -1422
rect 604 -1423 605 -1333
rect 688 -1450 689 -1422
rect 709 -1423 710 -1333
rect 737 -1450 738 -1422
rect 926 -1423 927 -1333
rect 989 -1450 990 -1422
rect 1087 -1423 1088 -1333
rect 1108 -1450 1109 -1422
rect 268 -1425 269 -1333
rect 338 -1450 339 -1424
rect 359 -1450 360 -1424
rect 499 -1425 500 -1333
rect 576 -1425 577 -1333
rect 604 -1450 605 -1424
rect 642 -1450 643 -1424
rect 891 -1450 892 -1424
rect 915 -1425 916 -1333
rect 926 -1450 927 -1424
rect 1003 -1425 1004 -1333
rect 1087 -1450 1088 -1424
rect 58 -1427 59 -1333
rect 1003 -1450 1004 -1426
rect 58 -1450 59 -1428
rect 72 -1429 73 -1333
rect 114 -1429 115 -1333
rect 268 -1450 269 -1428
rect 387 -1450 388 -1428
rect 639 -1450 640 -1428
rect 674 -1429 675 -1333
rect 709 -1450 710 -1428
rect 719 -1429 720 -1333
rect 1381 -1429 1382 -1333
rect 72 -1450 73 -1430
rect 226 -1431 227 -1333
rect 499 -1450 500 -1430
rect 506 -1431 507 -1333
rect 611 -1431 612 -1333
rect 674 -1450 675 -1430
rect 723 -1450 724 -1430
rect 1304 -1450 1305 -1430
rect 16 -1433 17 -1333
rect 611 -1450 612 -1432
rect 919 -1433 920 -1333
rect 1381 -1450 1382 -1432
rect 16 -1450 17 -1434
rect 408 -1435 409 -1333
rect 506 -1450 507 -1434
rect 1241 -1450 1242 -1434
rect 114 -1450 115 -1436
rect 345 -1437 346 -1333
rect 408 -1450 409 -1436
rect 807 -1437 808 -1333
rect 835 -1437 836 -1333
rect 919 -1450 920 -1436
rect 173 -1439 174 -1333
rect 576 -1450 577 -1438
rect 807 -1450 808 -1438
rect 849 -1439 850 -1333
rect 226 -1450 227 -1440
rect 233 -1441 234 -1333
rect 345 -1450 346 -1440
rect 422 -1441 423 -1333
rect 828 -1450 829 -1440
rect 835 -1450 836 -1440
rect 156 -1443 157 -1333
rect 233 -1450 234 -1442
rect 401 -1450 402 -1442
rect 849 -1450 850 -1442
rect 156 -1450 157 -1444
rect 177 -1445 178 -1333
rect 422 -1450 423 -1444
rect 471 -1445 472 -1333
rect 142 -1447 143 -1333
rect 177 -1450 178 -1446
rect 390 -1447 391 -1333
rect 471 -1450 472 -1446
rect 142 -1450 143 -1448
rect 824 -1450 825 -1448
rect 9 -1460 10 -1458
rect 33 -1460 34 -1458
rect 44 -1460 45 -1458
rect 457 -1460 458 -1458
rect 460 -1587 461 -1459
rect 940 -1460 941 -1458
rect 1454 -1460 1455 -1458
rect 1465 -1460 1466 -1458
rect 12 -1587 13 -1461
rect 268 -1462 269 -1458
rect 282 -1462 283 -1458
rect 520 -1462 521 -1458
rect 523 -1587 524 -1461
rect 709 -1462 710 -1458
rect 723 -1462 724 -1458
rect 835 -1462 836 -1458
rect 852 -1462 853 -1458
rect 1276 -1462 1277 -1458
rect 19 -1587 20 -1463
rect 1402 -1464 1403 -1458
rect 44 -1587 45 -1465
rect 485 -1466 486 -1458
rect 520 -1587 521 -1465
rect 688 -1466 689 -1458
rect 702 -1466 703 -1458
rect 782 -1466 783 -1458
rect 793 -1466 794 -1458
rect 1269 -1466 1270 -1458
rect 51 -1468 52 -1458
rect 509 -1468 510 -1458
rect 527 -1468 528 -1458
rect 527 -1587 528 -1467
rect 527 -1468 528 -1458
rect 527 -1587 528 -1467
rect 534 -1468 535 -1458
rect 590 -1468 591 -1458
rect 621 -1587 622 -1467
rect 1297 -1468 1298 -1458
rect 51 -1587 52 -1469
rect 730 -1470 731 -1458
rect 744 -1470 745 -1458
rect 1227 -1470 1228 -1458
rect 1269 -1587 1270 -1469
rect 1367 -1470 1368 -1458
rect 65 -1472 66 -1458
rect 537 -1472 538 -1458
rect 558 -1587 559 -1471
rect 1010 -1472 1011 -1458
rect 1297 -1587 1298 -1471
rect 1395 -1472 1396 -1458
rect 65 -1587 66 -1473
rect 870 -1474 871 -1458
rect 884 -1587 885 -1473
rect 1038 -1474 1039 -1458
rect 93 -1476 94 -1458
rect 488 -1587 489 -1475
rect 534 -1587 535 -1475
rect 667 -1476 668 -1458
rect 688 -1587 689 -1475
rect 695 -1476 696 -1458
rect 705 -1587 706 -1475
rect 1052 -1476 1053 -1458
rect 37 -1478 38 -1458
rect 93 -1587 94 -1477
rect 100 -1478 101 -1458
rect 548 -1478 549 -1458
rect 562 -1478 563 -1458
rect 1234 -1478 1235 -1458
rect 37 -1587 38 -1479
rect 898 -1480 899 -1458
rect 940 -1587 941 -1479
rect 996 -1480 997 -1458
rect 1010 -1587 1011 -1479
rect 1073 -1480 1074 -1458
rect 1234 -1587 1235 -1479
rect 1318 -1480 1319 -1458
rect 103 -1587 104 -1481
rect 450 -1482 451 -1458
rect 548 -1587 549 -1481
rect 604 -1482 605 -1458
rect 639 -1482 640 -1458
rect 1381 -1482 1382 -1458
rect 107 -1484 108 -1458
rect 117 -1587 118 -1483
rect 121 -1484 122 -1458
rect 152 -1484 153 -1458
rect 180 -1587 181 -1483
rect 730 -1587 731 -1483
rect 779 -1484 780 -1458
rect 1332 -1484 1333 -1458
rect 100 -1587 101 -1485
rect 107 -1587 108 -1485
rect 121 -1587 122 -1485
rect 415 -1486 416 -1458
rect 443 -1486 444 -1458
rect 765 -1486 766 -1458
rect 793 -1587 794 -1485
rect 842 -1486 843 -1458
rect 859 -1486 860 -1458
rect 1325 -1486 1326 -1458
rect 1332 -1587 1333 -1485
rect 1430 -1486 1431 -1458
rect 128 -1488 129 -1458
rect 1171 -1488 1172 -1458
rect 1318 -1587 1319 -1487
rect 1416 -1488 1417 -1458
rect 128 -1587 129 -1489
rect 422 -1490 423 -1458
rect 446 -1490 447 -1458
rect 1227 -1587 1228 -1489
rect 1325 -1587 1326 -1489
rect 1423 -1490 1424 -1458
rect 131 -1492 132 -1458
rect 432 -1587 433 -1491
rect 450 -1587 451 -1491
rect 653 -1492 654 -1458
rect 663 -1587 664 -1491
rect 1451 -1492 1452 -1458
rect 138 -1587 139 -1493
rect 800 -1494 801 -1458
rect 814 -1494 815 -1458
rect 1157 -1494 1158 -1458
rect 1171 -1587 1172 -1493
rect 1255 -1494 1256 -1458
rect 149 -1496 150 -1458
rect 849 -1496 850 -1458
rect 863 -1496 864 -1458
rect 1409 -1496 1410 -1458
rect 149 -1587 150 -1497
rect 170 -1498 171 -1458
rect 226 -1498 227 -1458
rect 226 -1587 227 -1497
rect 226 -1498 227 -1458
rect 226 -1587 227 -1497
rect 240 -1498 241 -1458
rect 537 -1587 538 -1497
rect 562 -1587 563 -1497
rect 618 -1498 619 -1458
rect 639 -1587 640 -1497
rect 660 -1498 661 -1458
rect 667 -1587 668 -1497
rect 737 -1498 738 -1458
rect 758 -1498 759 -1458
rect 779 -1587 780 -1497
rect 796 -1498 797 -1458
rect 1045 -1498 1046 -1458
rect 1052 -1587 1053 -1497
rect 1101 -1498 1102 -1458
rect 1157 -1587 1158 -1497
rect 1213 -1498 1214 -1458
rect 72 -1500 73 -1458
rect 170 -1587 171 -1499
rect 191 -1500 192 -1458
rect 240 -1587 241 -1499
rect 261 -1500 262 -1458
rect 604 -1587 605 -1499
rect 653 -1587 654 -1499
rect 681 -1500 682 -1458
rect 702 -1587 703 -1499
rect 1213 -1587 1214 -1499
rect 58 -1502 59 -1458
rect 72 -1587 73 -1501
rect 86 -1502 87 -1458
rect 191 -1587 192 -1501
rect 254 -1502 255 -1458
rect 261 -1587 262 -1501
rect 268 -1587 269 -1501
rect 408 -1502 409 -1458
rect 415 -1587 416 -1501
rect 611 -1502 612 -1458
rect 709 -1587 710 -1501
rect 747 -1502 748 -1458
rect 765 -1587 766 -1501
rect 786 -1502 787 -1458
rect 800 -1587 801 -1501
rect 1346 -1502 1347 -1458
rect 23 -1504 24 -1458
rect 786 -1587 787 -1503
rect 814 -1587 815 -1503
rect 877 -1504 878 -1458
rect 898 -1587 899 -1503
rect 1094 -1504 1095 -1458
rect 1192 -1504 1193 -1458
rect 1255 -1587 1256 -1503
rect 1346 -1587 1347 -1503
rect 1444 -1504 1445 -1458
rect 23 -1587 24 -1505
rect 54 -1587 55 -1505
rect 58 -1587 59 -1505
rect 310 -1506 311 -1458
rect 331 -1506 332 -1458
rect 695 -1587 696 -1505
rect 716 -1506 717 -1458
rect 744 -1587 745 -1505
rect 817 -1506 818 -1458
rect 1087 -1506 1088 -1458
rect 1094 -1587 1095 -1505
rect 1311 -1506 1312 -1458
rect 16 -1508 17 -1458
rect 310 -1587 311 -1507
rect 338 -1508 339 -1458
rect 422 -1587 423 -1507
rect 478 -1508 479 -1458
rect 618 -1587 619 -1507
rect 716 -1587 717 -1507
rect 751 -1508 752 -1458
rect 821 -1587 822 -1507
rect 894 -1587 895 -1507
rect 982 -1508 983 -1458
rect 1276 -1587 1277 -1507
rect 16 -1587 17 -1509
rect 681 -1587 682 -1509
rect 723 -1587 724 -1509
rect 772 -1510 773 -1458
rect 824 -1510 825 -1458
rect 1374 -1510 1375 -1458
rect 219 -1512 220 -1458
rect 331 -1587 332 -1511
rect 338 -1587 339 -1511
rect 499 -1512 500 -1458
rect 565 -1512 566 -1458
rect 751 -1587 752 -1511
rect 828 -1587 829 -1511
rect 1185 -1512 1186 -1458
rect 1192 -1587 1193 -1511
rect 1290 -1512 1291 -1458
rect 2 -1514 3 -1458
rect 219 -1587 220 -1513
rect 247 -1514 248 -1458
rect 254 -1587 255 -1513
rect 282 -1587 283 -1513
rect 345 -1514 346 -1458
rect 380 -1514 381 -1458
rect 443 -1587 444 -1513
rect 478 -1587 479 -1513
rect 492 -1514 493 -1458
rect 572 -1587 573 -1513
rect 866 -1514 867 -1458
rect 870 -1587 871 -1513
rect 1017 -1514 1018 -1458
rect 1038 -1587 1039 -1513
rect 1080 -1514 1081 -1458
rect 1185 -1587 1186 -1513
rect 1283 -1514 1284 -1458
rect 2 -1587 3 -1515
rect 275 -1516 276 -1458
rect 289 -1516 290 -1458
rect 772 -1587 773 -1515
rect 831 -1516 832 -1458
rect 1122 -1516 1123 -1458
rect 1199 -1516 1200 -1458
rect 1311 -1587 1312 -1515
rect 9 -1587 10 -1517
rect 275 -1587 276 -1517
rect 289 -1587 290 -1517
rect 457 -1587 458 -1517
rect 485 -1587 486 -1517
rect 758 -1587 759 -1517
rect 831 -1587 832 -1517
rect 1360 -1518 1361 -1458
rect 114 -1520 115 -1458
rect 499 -1587 500 -1519
rect 583 -1520 584 -1458
rect 642 -1520 643 -1458
rect 835 -1587 836 -1519
rect 891 -1520 892 -1458
rect 905 -1520 906 -1458
rect 1122 -1587 1123 -1519
rect 1129 -1520 1130 -1458
rect 1199 -1587 1200 -1519
rect 1283 -1587 1284 -1519
rect 1388 -1520 1389 -1458
rect 40 -1587 41 -1521
rect 583 -1587 584 -1521
rect 590 -1587 591 -1521
rect 674 -1522 675 -1458
rect 842 -1587 843 -1521
rect 912 -1522 913 -1458
rect 954 -1522 955 -1458
rect 982 -1587 983 -1521
rect 996 -1587 997 -1521
rect 1150 -1522 1151 -1458
rect 89 -1587 90 -1523
rect 912 -1587 913 -1523
rect 1059 -1524 1060 -1458
rect 1101 -1587 1102 -1523
rect 1129 -1587 1130 -1523
rect 1178 -1524 1179 -1458
rect 30 -1526 31 -1458
rect 1178 -1587 1179 -1525
rect 30 -1587 31 -1527
rect 359 -1528 360 -1458
rect 380 -1587 381 -1527
rect 597 -1528 598 -1458
rect 611 -1587 612 -1527
rect 646 -1528 647 -1458
rect 649 -1528 650 -1458
rect 674 -1587 675 -1527
rect 807 -1528 808 -1458
rect 954 -1587 955 -1527
rect 1073 -1587 1074 -1527
rect 1304 -1528 1305 -1458
rect 114 -1587 115 -1529
rect 737 -1587 738 -1529
rect 849 -1587 850 -1529
rect 919 -1530 920 -1458
rect 1080 -1587 1081 -1529
rect 1220 -1530 1221 -1458
rect 1304 -1587 1305 -1529
rect 1339 -1530 1340 -1458
rect 142 -1532 143 -1458
rect 1017 -1587 1018 -1531
rect 1115 -1532 1116 -1458
rect 1220 -1587 1221 -1531
rect 1339 -1587 1340 -1531
rect 1437 -1532 1438 -1458
rect 142 -1587 143 -1533
rect 233 -1534 234 -1458
rect 317 -1534 318 -1458
rect 1059 -1587 1060 -1533
rect 1108 -1534 1109 -1458
rect 1115 -1587 1116 -1533
rect 1150 -1587 1151 -1533
rect 1241 -1534 1242 -1458
rect 198 -1536 199 -1458
rect 247 -1587 248 -1535
rect 324 -1536 325 -1458
rect 905 -1587 906 -1535
rect 919 -1587 920 -1535
rect 961 -1536 962 -1458
rect 82 -1538 83 -1458
rect 324 -1587 325 -1537
rect 345 -1587 346 -1537
rect 366 -1538 367 -1458
rect 397 -1538 398 -1458
rect 1136 -1538 1137 -1458
rect 198 -1587 199 -1539
rect 212 -1540 213 -1458
rect 233 -1587 234 -1539
rect 303 -1540 304 -1458
rect 352 -1540 353 -1458
rect 359 -1587 360 -1539
rect 366 -1587 367 -1539
rect 576 -1540 577 -1458
rect 625 -1540 626 -1458
rect 646 -1587 647 -1539
rect 859 -1587 860 -1539
rect 1136 -1587 1137 -1539
rect 177 -1542 178 -1458
rect 212 -1587 213 -1541
rect 296 -1542 297 -1458
rect 303 -1587 304 -1541
rect 352 -1587 353 -1541
rect 373 -1542 374 -1458
rect 404 -1587 405 -1541
rect 632 -1542 633 -1458
rect 863 -1587 864 -1541
rect 933 -1542 934 -1458
rect 961 -1587 962 -1541
rect 1024 -1542 1025 -1458
rect 135 -1544 136 -1458
rect 296 -1587 297 -1543
rect 373 -1587 374 -1543
rect 387 -1544 388 -1458
rect 408 -1587 409 -1543
rect 492 -1587 493 -1543
rect 513 -1544 514 -1458
rect 576 -1587 577 -1543
rect 625 -1587 626 -1543
rect 926 -1544 927 -1458
rect 933 -1587 934 -1543
rect 989 -1544 990 -1458
rect 1024 -1587 1025 -1543
rect 1206 -1544 1207 -1458
rect 79 -1546 80 -1458
rect 513 -1587 514 -1545
rect 541 -1546 542 -1458
rect 807 -1587 808 -1545
rect 877 -1587 878 -1545
rect 947 -1546 948 -1458
rect 968 -1546 969 -1458
rect 989 -1587 990 -1545
rect 1143 -1546 1144 -1458
rect 1206 -1587 1207 -1545
rect 79 -1587 80 -1547
rect 86 -1587 87 -1547
rect 135 -1587 136 -1547
rect 1241 -1587 1242 -1547
rect 205 -1550 206 -1458
rect 317 -1587 318 -1549
rect 387 -1587 388 -1549
rect 464 -1550 465 -1458
rect 541 -1587 542 -1549
rect 569 -1550 570 -1458
rect 891 -1587 892 -1549
rect 1262 -1550 1263 -1458
rect 205 -1587 206 -1551
rect 551 -1552 552 -1458
rect 555 -1552 556 -1458
rect 597 -1587 598 -1551
rect 926 -1587 927 -1551
rect 975 -1552 976 -1458
rect 1143 -1587 1144 -1551
rect 1164 -1552 1165 -1458
rect 1262 -1587 1263 -1551
rect 1353 -1552 1354 -1458
rect 394 -1554 395 -1458
rect 464 -1587 465 -1553
rect 555 -1587 556 -1553
rect 1045 -1587 1046 -1553
rect 1353 -1587 1354 -1553
rect 1458 -1554 1459 -1458
rect 394 -1587 395 -1555
rect 436 -1556 437 -1458
rect 569 -1587 570 -1555
rect 1290 -1587 1291 -1555
rect 401 -1558 402 -1458
rect 436 -1587 437 -1557
rect 856 -1558 857 -1458
rect 975 -1587 976 -1557
rect 163 -1560 164 -1458
rect 401 -1587 402 -1559
rect 429 -1560 430 -1458
rect 632 -1587 633 -1559
rect 856 -1587 857 -1559
rect 1108 -1587 1109 -1559
rect 163 -1587 164 -1561
rect 1003 -1562 1004 -1458
rect 429 -1587 430 -1563
rect 1087 -1587 1088 -1563
rect 887 -1566 888 -1458
rect 1164 -1587 1165 -1565
rect 947 -1587 948 -1567
rect 1048 -1587 1049 -1567
rect 968 -1587 969 -1569
rect 1031 -1570 1032 -1458
rect 145 -1587 146 -1571
rect 1031 -1587 1032 -1571
rect 1003 -1587 1004 -1573
rect 1066 -1574 1067 -1458
rect 1066 -1587 1067 -1575
rect 1248 -1576 1249 -1458
rect 506 -1578 507 -1458
rect 1248 -1587 1249 -1577
rect 471 -1580 472 -1458
rect 506 -1587 507 -1579
rect 184 -1582 185 -1458
rect 471 -1587 472 -1581
rect 156 -1584 157 -1458
rect 184 -1587 185 -1583
rect 156 -1587 157 -1585
rect 803 -1587 804 -1585
rect 2 -1597 3 -1595
rect 558 -1597 559 -1595
rect 569 -1597 570 -1595
rect 849 -1597 850 -1595
rect 856 -1597 857 -1595
rect 1066 -1597 1067 -1595
rect 1094 -1597 1095 -1595
rect 1097 -1623 1098 -1596
rect 1255 -1597 1256 -1595
rect 1258 -1597 1259 -1595
rect 2 -1718 3 -1598
rect 401 -1718 402 -1598
rect 415 -1599 416 -1595
rect 569 -1718 570 -1598
rect 572 -1599 573 -1595
rect 576 -1599 577 -1595
rect 632 -1599 633 -1595
rect 663 -1599 664 -1595
rect 705 -1599 706 -1595
rect 954 -1599 955 -1595
rect 1045 -1599 1046 -1595
rect 1346 -1599 1347 -1595
rect 9 -1718 10 -1600
rect 940 -1601 941 -1595
rect 954 -1718 955 -1600
rect 1129 -1601 1130 -1595
rect 1255 -1718 1256 -1600
rect 1283 -1601 1284 -1595
rect 12 -1603 13 -1595
rect 163 -1603 164 -1595
rect 177 -1603 178 -1595
rect 212 -1603 213 -1595
rect 233 -1603 234 -1595
rect 233 -1718 234 -1602
rect 233 -1603 234 -1595
rect 233 -1718 234 -1602
rect 320 -1718 321 -1602
rect 905 -1603 906 -1595
rect 940 -1718 941 -1602
rect 1318 -1603 1319 -1595
rect 51 -1605 52 -1595
rect 583 -1605 584 -1595
rect 632 -1718 633 -1604
rect 716 -1605 717 -1595
rect 754 -1718 755 -1604
rect 1136 -1605 1137 -1595
rect 1304 -1605 1305 -1595
rect 1318 -1718 1319 -1604
rect 58 -1607 59 -1595
rect 415 -1718 416 -1606
rect 464 -1607 465 -1595
rect 464 -1718 465 -1606
rect 464 -1607 465 -1595
rect 464 -1718 465 -1606
rect 478 -1607 479 -1595
rect 478 -1718 479 -1606
rect 478 -1607 479 -1595
rect 478 -1718 479 -1606
rect 485 -1607 486 -1595
rect 639 -1607 640 -1595
rect 660 -1607 661 -1595
rect 688 -1607 689 -1595
rect 716 -1718 717 -1606
rect 737 -1607 738 -1595
rect 775 -1718 776 -1606
rect 863 -1607 864 -1595
rect 884 -1607 885 -1595
rect 905 -1718 906 -1606
rect 975 -1607 976 -1595
rect 1136 -1718 1137 -1606
rect 1304 -1718 1305 -1606
rect 1332 -1607 1333 -1595
rect 58 -1718 59 -1608
rect 513 -1609 514 -1595
rect 534 -1609 535 -1595
rect 982 -1609 983 -1595
rect 1045 -1718 1046 -1608
rect 1108 -1609 1109 -1595
rect 1129 -1718 1130 -1608
rect 1171 -1609 1172 -1595
rect 65 -1611 66 -1595
rect 551 -1718 552 -1610
rect 639 -1718 640 -1610
rect 674 -1611 675 -1595
rect 688 -1718 689 -1610
rect 765 -1611 766 -1595
rect 800 -1611 801 -1595
rect 1199 -1611 1200 -1595
rect 65 -1718 66 -1612
rect 702 -1613 703 -1595
rect 765 -1718 766 -1612
rect 779 -1613 780 -1595
rect 803 -1613 804 -1595
rect 1108 -1718 1109 -1612
rect 1199 -1718 1200 -1612
rect 1234 -1613 1235 -1595
rect 79 -1615 80 -1595
rect 800 -1718 801 -1614
rect 849 -1718 850 -1614
rect 870 -1615 871 -1595
rect 884 -1718 885 -1614
rect 898 -1615 899 -1595
rect 975 -1718 976 -1614
rect 1052 -1615 1053 -1595
rect 1094 -1718 1095 -1614
rect 1234 -1718 1235 -1614
rect 1325 -1615 1326 -1595
rect 86 -1617 87 -1595
rect 488 -1718 489 -1616
rect 495 -1617 496 -1595
rect 548 -1617 549 -1595
rect 625 -1617 626 -1595
rect 674 -1718 675 -1616
rect 779 -1718 780 -1616
rect 814 -1617 815 -1595
rect 856 -1718 857 -1616
rect 1328 -1718 1329 -1616
rect 86 -1718 87 -1618
rect 107 -1619 108 -1595
rect 110 -1718 111 -1618
rect 576 -1718 577 -1618
rect 621 -1619 622 -1595
rect 625 -1718 626 -1618
rect 660 -1718 661 -1618
rect 1003 -1619 1004 -1595
rect 1052 -1718 1053 -1618
rect 1122 -1619 1123 -1595
rect 1220 -1619 1221 -1595
rect 1325 -1718 1326 -1618
rect 40 -1621 41 -1595
rect 1003 -1718 1004 -1620
rect 1220 -1718 1221 -1620
rect 1276 -1621 1277 -1595
rect 89 -1623 90 -1595
rect 709 -1623 710 -1595
rect 814 -1718 815 -1622
rect 842 -1623 843 -1595
rect 859 -1623 860 -1595
rect 1059 -1623 1060 -1595
rect 1258 -1718 1259 -1622
rect 1283 -1718 1284 -1622
rect 100 -1625 101 -1595
rect 1185 -1625 1186 -1595
rect 1276 -1718 1277 -1624
rect 1353 -1625 1354 -1595
rect 23 -1627 24 -1595
rect 100 -1718 101 -1626
rect 107 -1718 108 -1626
rect 583 -1718 584 -1626
rect 709 -1718 710 -1626
rect 744 -1627 745 -1595
rect 842 -1718 843 -1626
rect 877 -1627 878 -1595
rect 891 -1718 892 -1626
rect 1262 -1627 1263 -1595
rect 117 -1629 118 -1595
rect 184 -1629 185 -1595
rect 194 -1718 195 -1628
rect 380 -1629 381 -1595
rect 499 -1629 500 -1595
rect 534 -1718 535 -1628
rect 537 -1629 538 -1595
rect 702 -1718 703 -1628
rect 737 -1718 738 -1628
rect 744 -1718 745 -1628
rect 863 -1718 864 -1628
rect 919 -1629 920 -1595
rect 947 -1629 948 -1595
rect 1185 -1718 1186 -1628
rect 1262 -1718 1263 -1628
rect 1290 -1629 1291 -1595
rect 138 -1631 139 -1595
rect 471 -1631 472 -1595
rect 485 -1718 486 -1630
rect 499 -1718 500 -1630
rect 506 -1631 507 -1595
rect 523 -1631 524 -1595
rect 730 -1631 731 -1595
rect 947 -1718 948 -1630
rect 982 -1718 983 -1630
rect 1038 -1631 1039 -1595
rect 1290 -1718 1291 -1630
rect 1311 -1631 1312 -1595
rect 142 -1633 143 -1595
rect 1101 -1633 1102 -1595
rect 1311 -1718 1312 -1632
rect 1339 -1633 1340 -1595
rect 47 -1718 48 -1634
rect 142 -1718 143 -1634
rect 145 -1635 146 -1595
rect 254 -1635 255 -1595
rect 338 -1635 339 -1595
rect 457 -1635 458 -1595
rect 471 -1718 472 -1634
rect 611 -1635 612 -1595
rect 730 -1718 731 -1634
rect 747 -1718 748 -1634
rect 870 -1718 871 -1634
rect 968 -1635 969 -1595
rect 996 -1635 997 -1595
rect 1038 -1718 1039 -1634
rect 1080 -1635 1081 -1595
rect 1101 -1718 1102 -1634
rect 93 -1637 94 -1595
rect 338 -1718 339 -1636
rect 345 -1637 346 -1595
rect 345 -1718 346 -1636
rect 345 -1637 346 -1595
rect 345 -1718 346 -1636
rect 352 -1637 353 -1595
rect 457 -1718 458 -1636
rect 506 -1718 507 -1636
rect 961 -1637 962 -1595
rect 968 -1718 969 -1636
rect 989 -1637 990 -1595
rect 996 -1718 997 -1636
rect 1164 -1637 1165 -1595
rect 93 -1718 94 -1638
rect 1206 -1639 1207 -1595
rect 103 -1641 104 -1595
rect 989 -1718 990 -1640
rect 1164 -1718 1165 -1640
rect 1213 -1641 1214 -1595
rect 135 -1643 136 -1595
rect 1213 -1718 1214 -1642
rect 135 -1718 136 -1644
rect 198 -1645 199 -1595
rect 212 -1718 213 -1644
rect 247 -1645 248 -1595
rect 254 -1718 255 -1644
rect 429 -1645 430 -1595
rect 443 -1645 444 -1595
rect 611 -1718 612 -1644
rect 877 -1718 878 -1644
rect 933 -1645 934 -1595
rect 961 -1718 962 -1644
rect 1031 -1645 1032 -1595
rect 1206 -1718 1207 -1644
rect 1227 -1645 1228 -1595
rect 121 -1647 122 -1595
rect 443 -1718 444 -1646
rect 460 -1647 461 -1595
rect 933 -1718 934 -1646
rect 1031 -1718 1032 -1646
rect 1087 -1647 1088 -1595
rect 1157 -1647 1158 -1595
rect 1227 -1718 1228 -1646
rect 114 -1649 115 -1595
rect 1087 -1718 1088 -1648
rect 96 -1718 97 -1650
rect 114 -1718 115 -1650
rect 121 -1718 122 -1650
rect 240 -1651 241 -1595
rect 247 -1718 248 -1650
rect 275 -1651 276 -1595
rect 352 -1718 353 -1650
rect 492 -1651 493 -1595
rect 513 -1718 514 -1650
rect 758 -1651 759 -1595
rect 894 -1718 895 -1650
rect 1178 -1651 1179 -1595
rect 152 -1718 153 -1652
rect 282 -1653 283 -1595
rect 366 -1653 367 -1595
rect 432 -1653 433 -1595
rect 492 -1718 493 -1652
rect 527 -1653 528 -1595
rect 758 -1718 759 -1652
rect 772 -1653 773 -1595
rect 1066 -1718 1067 -1652
rect 1178 -1718 1179 -1652
rect 159 -1718 160 -1654
rect 1059 -1718 1060 -1654
rect 1073 -1655 1074 -1595
rect 1157 -1718 1158 -1654
rect 163 -1718 164 -1656
rect 831 -1657 832 -1595
rect 1024 -1657 1025 -1595
rect 1073 -1718 1074 -1656
rect 177 -1718 178 -1658
rect 751 -1659 752 -1595
rect 772 -1718 773 -1658
rect 1115 -1659 1116 -1595
rect 180 -1661 181 -1595
rect 359 -1661 360 -1595
rect 366 -1718 367 -1660
rect 562 -1661 563 -1595
rect 751 -1718 752 -1660
rect 919 -1718 920 -1660
rect 1024 -1718 1025 -1660
rect 1241 -1661 1242 -1595
rect 44 -1663 45 -1595
rect 359 -1718 360 -1662
rect 373 -1663 374 -1595
rect 429 -1718 430 -1662
rect 523 -1718 524 -1662
rect 1171 -1718 1172 -1662
rect 1241 -1718 1242 -1662
rect 1269 -1663 1270 -1595
rect 44 -1718 45 -1664
rect 54 -1665 55 -1595
rect 184 -1718 185 -1664
rect 205 -1665 206 -1595
rect 240 -1718 241 -1664
rect 296 -1665 297 -1595
rect 376 -1718 377 -1664
rect 1017 -1665 1018 -1595
rect 1115 -1718 1116 -1664
rect 1143 -1665 1144 -1595
rect 54 -1718 55 -1666
rect 79 -1718 80 -1666
rect 198 -1718 199 -1666
rect 331 -1667 332 -1595
rect 380 -1718 381 -1666
rect 422 -1667 423 -1595
rect 450 -1667 451 -1595
rect 1017 -1718 1018 -1666
rect 1143 -1718 1144 -1666
rect 1192 -1667 1193 -1595
rect 51 -1718 52 -1668
rect 1192 -1718 1193 -1668
rect 205 -1718 206 -1670
rect 404 -1671 405 -1595
rect 422 -1718 423 -1670
rect 436 -1671 437 -1595
rect 450 -1718 451 -1670
rect 695 -1671 696 -1595
rect 828 -1671 829 -1595
rect 1269 -1718 1270 -1670
rect 226 -1673 227 -1595
rect 296 -1718 297 -1672
rect 324 -1673 325 -1595
rect 828 -1718 829 -1672
rect 226 -1718 227 -1674
rect 310 -1675 311 -1595
rect 324 -1718 325 -1674
rect 387 -1675 388 -1595
rect 394 -1675 395 -1595
rect 436 -1718 437 -1674
rect 527 -1718 528 -1674
rect 541 -1675 542 -1595
rect 562 -1718 563 -1674
rect 670 -1718 671 -1674
rect 695 -1718 696 -1674
rect 901 -1718 902 -1674
rect 128 -1677 129 -1595
rect 387 -1718 388 -1676
rect 394 -1718 395 -1676
rect 597 -1677 598 -1595
rect 72 -1679 73 -1595
rect 128 -1718 129 -1678
rect 275 -1718 276 -1678
rect 289 -1679 290 -1595
rect 303 -1679 304 -1595
rect 310 -1718 311 -1678
rect 331 -1718 332 -1678
rect 520 -1679 521 -1595
rect 541 -1718 542 -1678
rect 786 -1679 787 -1595
rect 72 -1718 73 -1680
rect 261 -1681 262 -1595
rect 282 -1718 283 -1680
rect 618 -1681 619 -1595
rect 786 -1718 787 -1680
rect 821 -1681 822 -1595
rect 156 -1683 157 -1595
rect 261 -1718 262 -1682
rect 404 -1718 405 -1682
rect 460 -1718 461 -1682
rect 555 -1683 556 -1595
rect 618 -1718 619 -1682
rect 821 -1718 822 -1682
rect 898 -1718 899 -1682
rect 30 -1685 31 -1595
rect 555 -1718 556 -1684
rect 590 -1685 591 -1595
rect 597 -1718 598 -1684
rect 16 -1687 17 -1595
rect 30 -1718 31 -1686
rect 170 -1687 171 -1595
rect 303 -1718 304 -1686
rect 408 -1687 409 -1595
rect 590 -1718 591 -1686
rect 170 -1718 171 -1688
rect 268 -1689 269 -1595
rect 408 -1718 409 -1688
rect 604 -1689 605 -1595
rect 149 -1691 150 -1595
rect 268 -1718 269 -1690
rect 604 -1718 605 -1690
rect 646 -1691 647 -1595
rect 149 -1718 150 -1692
rect 912 -1693 913 -1595
rect 219 -1695 220 -1595
rect 289 -1718 290 -1694
rect 520 -1718 521 -1694
rect 912 -1718 913 -1694
rect 191 -1697 192 -1595
rect 219 -1718 220 -1696
rect 646 -1718 647 -1696
rect 681 -1697 682 -1595
rect 191 -1718 192 -1698
rect 653 -1699 654 -1595
rect 681 -1718 682 -1698
rect 723 -1699 724 -1595
rect 653 -1718 654 -1700
rect 667 -1701 668 -1595
rect 723 -1718 724 -1700
rect 793 -1701 794 -1595
rect 667 -1718 668 -1702
rect 1297 -1703 1298 -1595
rect 793 -1718 794 -1704
rect 807 -1705 808 -1595
rect 1248 -1705 1249 -1595
rect 1297 -1718 1298 -1704
rect 37 -1707 38 -1595
rect 1248 -1718 1249 -1706
rect 37 -1718 38 -1708
rect 317 -1709 318 -1595
rect 807 -1718 808 -1708
rect 835 -1709 836 -1595
rect 317 -1718 318 -1710
rect 1080 -1718 1081 -1710
rect 835 -1718 836 -1712
rect 926 -1713 927 -1595
rect 926 -1718 927 -1714
rect 1010 -1715 1011 -1595
rect 373 -1718 374 -1716
rect 1010 -1718 1011 -1716
rect 9 -1728 10 -1726
rect 110 -1728 111 -1726
rect 117 -1837 118 -1727
rect 646 -1728 647 -1726
rect 667 -1728 668 -1726
rect 933 -1728 934 -1726
rect 940 -1728 941 -1726
rect 968 -1728 969 -1726
rect 1069 -1728 1070 -1726
rect 1241 -1728 1242 -1726
rect 1318 -1728 1319 -1726
rect 1328 -1728 1329 -1726
rect 16 -1730 17 -1726
rect 30 -1730 31 -1726
rect 33 -1730 34 -1726
rect 68 -1837 69 -1729
rect 72 -1730 73 -1726
rect 373 -1730 374 -1726
rect 390 -1837 391 -1729
rect 856 -1730 857 -1726
rect 898 -1730 899 -1726
rect 1101 -1730 1102 -1726
rect 1122 -1730 1123 -1726
rect 1276 -1730 1277 -1726
rect 16 -1837 17 -1731
rect 149 -1732 150 -1726
rect 152 -1732 153 -1726
rect 1101 -1837 1102 -1731
rect 1122 -1837 1123 -1731
rect 1171 -1732 1172 -1726
rect 1227 -1732 1228 -1726
rect 1286 -1837 1287 -1731
rect 9 -1837 10 -1733
rect 152 -1837 153 -1733
rect 205 -1734 206 -1726
rect 355 -1837 356 -1733
rect 359 -1734 360 -1726
rect 646 -1837 647 -1733
rect 667 -1837 668 -1733
rect 702 -1734 703 -1726
rect 712 -1837 713 -1733
rect 765 -1734 766 -1726
rect 814 -1734 815 -1726
rect 891 -1837 892 -1733
rect 898 -1837 899 -1733
rect 975 -1734 976 -1726
rect 1171 -1837 1172 -1733
rect 1213 -1734 1214 -1726
rect 1241 -1837 1242 -1733
rect 1290 -1734 1291 -1726
rect 19 -1736 20 -1726
rect 793 -1736 794 -1726
rect 828 -1736 829 -1726
rect 828 -1837 829 -1735
rect 828 -1736 829 -1726
rect 828 -1837 829 -1735
rect 835 -1736 836 -1726
rect 856 -1837 857 -1735
rect 901 -1736 902 -1726
rect 1276 -1837 1277 -1735
rect 23 -1738 24 -1726
rect 611 -1738 612 -1726
rect 702 -1837 703 -1737
rect 723 -1738 724 -1726
rect 744 -1738 745 -1726
rect 849 -1738 850 -1726
rect 933 -1837 934 -1737
rect 947 -1738 948 -1726
rect 968 -1837 969 -1737
rect 1045 -1738 1046 -1726
rect 1213 -1837 1214 -1737
rect 1255 -1738 1256 -1726
rect 26 -1740 27 -1726
rect 100 -1740 101 -1726
rect 107 -1740 108 -1726
rect 1017 -1740 1018 -1726
rect 1255 -1837 1256 -1739
rect 1304 -1740 1305 -1726
rect 26 -1837 27 -1741
rect 982 -1742 983 -1726
rect 1010 -1742 1011 -1726
rect 1045 -1837 1046 -1741
rect 30 -1837 31 -1743
rect 268 -1744 269 -1726
rect 324 -1744 325 -1726
rect 376 -1744 377 -1726
rect 404 -1744 405 -1726
rect 534 -1744 535 -1726
rect 548 -1744 549 -1726
rect 793 -1837 794 -1743
rect 835 -1837 836 -1743
rect 870 -1744 871 -1726
rect 940 -1837 941 -1743
rect 996 -1744 997 -1726
rect 1017 -1837 1018 -1743
rect 1073 -1744 1074 -1726
rect 37 -1746 38 -1726
rect 159 -1746 160 -1726
rect 205 -1837 206 -1745
rect 310 -1746 311 -1726
rect 359 -1837 360 -1745
rect 387 -1746 388 -1726
rect 457 -1746 458 -1726
rect 1297 -1746 1298 -1726
rect 44 -1748 45 -1726
rect 240 -1748 241 -1726
rect 268 -1837 269 -1747
rect 415 -1748 416 -1726
rect 457 -1837 458 -1747
rect 551 -1748 552 -1726
rect 555 -1748 556 -1726
rect 632 -1748 633 -1726
rect 719 -1837 720 -1747
rect 884 -1748 885 -1726
rect 975 -1837 976 -1747
rect 1031 -1748 1032 -1726
rect 1073 -1837 1074 -1747
rect 1115 -1748 1116 -1726
rect 44 -1837 45 -1749
rect 1059 -1750 1060 -1726
rect 1115 -1837 1116 -1749
rect 1164 -1750 1165 -1726
rect 47 -1837 48 -1751
rect 996 -1837 997 -1751
rect 1031 -1837 1032 -1751
rect 1094 -1752 1095 -1726
rect 1164 -1837 1165 -1751
rect 1192 -1752 1193 -1726
rect 54 -1754 55 -1726
rect 1248 -1754 1249 -1726
rect 72 -1837 73 -1755
rect 93 -1756 94 -1726
rect 100 -1837 101 -1755
rect 467 -1837 468 -1755
rect 478 -1756 479 -1726
rect 478 -1837 479 -1755
rect 478 -1756 479 -1726
rect 478 -1837 479 -1755
rect 485 -1756 486 -1726
rect 1227 -1837 1228 -1755
rect 1234 -1756 1235 -1726
rect 1248 -1837 1249 -1755
rect 51 -1758 52 -1726
rect 93 -1837 94 -1757
rect 107 -1837 108 -1757
rect 289 -1758 290 -1726
rect 369 -1837 370 -1757
rect 744 -1837 745 -1757
rect 747 -1758 748 -1726
rect 821 -1758 822 -1726
rect 849 -1837 850 -1757
rect 912 -1758 913 -1726
rect 1059 -1837 1060 -1757
rect 1108 -1758 1109 -1726
rect 1192 -1837 1193 -1757
rect 1220 -1758 1221 -1726
rect 1234 -1837 1235 -1757
rect 1283 -1758 1284 -1726
rect 51 -1837 52 -1759
rect 842 -1760 843 -1726
rect 912 -1837 913 -1759
rect 989 -1760 990 -1726
rect 1108 -1837 1109 -1759
rect 1150 -1760 1151 -1726
rect 1220 -1837 1221 -1759
rect 1269 -1760 1270 -1726
rect 58 -1762 59 -1726
rect 842 -1837 843 -1761
rect 989 -1837 990 -1761
rect 1052 -1762 1053 -1726
rect 1269 -1837 1270 -1761
rect 1311 -1762 1312 -1726
rect 58 -1837 59 -1763
rect 184 -1764 185 -1726
rect 212 -1764 213 -1726
rect 212 -1837 213 -1763
rect 212 -1764 213 -1726
rect 212 -1837 213 -1763
rect 226 -1764 227 -1726
rect 523 -1764 524 -1726
rect 534 -1837 535 -1763
rect 807 -1764 808 -1726
rect 821 -1837 822 -1763
rect 926 -1764 927 -1726
rect 1052 -1837 1053 -1763
rect 1087 -1764 1088 -1726
rect 2 -1766 3 -1726
rect 226 -1837 227 -1765
rect 233 -1766 234 -1726
rect 240 -1837 241 -1765
rect 275 -1766 276 -1726
rect 324 -1837 325 -1765
rect 373 -1837 374 -1765
rect 614 -1837 615 -1765
rect 625 -1766 626 -1726
rect 807 -1837 808 -1765
rect 926 -1837 927 -1765
rect 1003 -1766 1004 -1726
rect 1087 -1837 1088 -1765
rect 1143 -1766 1144 -1726
rect 2 -1837 3 -1767
rect 54 -1837 55 -1767
rect 79 -1768 80 -1726
rect 586 -1837 587 -1767
rect 604 -1768 605 -1726
rect 947 -1837 948 -1767
rect 1143 -1837 1144 -1767
rect 1185 -1768 1186 -1726
rect 79 -1837 80 -1769
rect 86 -1770 87 -1726
rect 121 -1770 122 -1726
rect 317 -1770 318 -1726
rect 401 -1770 402 -1726
rect 1185 -1837 1186 -1769
rect 86 -1837 87 -1771
rect 299 -1837 300 -1771
rect 317 -1837 318 -1771
rect 331 -1772 332 -1726
rect 401 -1837 402 -1771
rect 422 -1772 423 -1726
rect 488 -1772 489 -1726
rect 894 -1772 895 -1726
rect 114 -1774 115 -1726
rect 121 -1837 122 -1773
rect 128 -1774 129 -1726
rect 289 -1837 290 -1773
rect 331 -1837 332 -1773
rect 345 -1774 346 -1726
rect 415 -1837 416 -1773
rect 436 -1774 437 -1726
rect 506 -1774 507 -1726
rect 642 -1837 643 -1773
rect 660 -1774 661 -1726
rect 884 -1837 885 -1773
rect 128 -1837 129 -1775
rect 261 -1776 262 -1726
rect 345 -1837 346 -1775
rect 380 -1776 381 -1726
rect 436 -1837 437 -1775
rect 471 -1776 472 -1726
rect 506 -1837 507 -1775
rect 541 -1776 542 -1726
rect 555 -1837 556 -1775
rect 772 -1776 773 -1726
rect 138 -1837 139 -1777
rect 303 -1778 304 -1726
rect 464 -1778 465 -1726
rect 471 -1837 472 -1777
rect 513 -1778 514 -1726
rect 548 -1837 549 -1777
rect 576 -1778 577 -1726
rect 1094 -1837 1095 -1777
rect 142 -1780 143 -1726
rect 1283 -1837 1284 -1779
rect 142 -1837 143 -1781
rect 481 -1837 482 -1781
rect 513 -1837 514 -1781
rect 527 -1782 528 -1726
rect 541 -1837 542 -1781
rect 562 -1782 563 -1726
rect 576 -1837 577 -1781
rect 597 -1782 598 -1726
rect 611 -1837 612 -1781
rect 688 -1782 689 -1726
rect 723 -1837 724 -1781
rect 775 -1782 776 -1726
rect 149 -1837 150 -1783
rect 590 -1784 591 -1726
rect 597 -1837 598 -1783
rect 639 -1784 640 -1726
rect 660 -1837 661 -1783
rect 681 -1784 682 -1726
rect 730 -1784 731 -1726
rect 1010 -1837 1011 -1783
rect 156 -1786 157 -1726
rect 590 -1837 591 -1785
rect 625 -1837 626 -1785
rect 863 -1786 864 -1726
rect 156 -1837 157 -1787
rect 170 -1788 171 -1726
rect 177 -1788 178 -1726
rect 681 -1837 682 -1787
rect 730 -1837 731 -1787
rect 919 -1788 920 -1726
rect 96 -1790 97 -1726
rect 919 -1837 920 -1789
rect 163 -1792 164 -1726
rect 380 -1837 381 -1791
rect 408 -1792 409 -1726
rect 527 -1837 528 -1791
rect 562 -1837 563 -1791
rect 618 -1792 619 -1726
rect 628 -1837 629 -1791
rect 1003 -1837 1004 -1791
rect 170 -1837 171 -1793
rect 282 -1794 283 -1726
rect 394 -1794 395 -1726
rect 408 -1837 409 -1793
rect 464 -1837 465 -1793
rect 982 -1837 983 -1793
rect 177 -1837 178 -1795
rect 296 -1796 297 -1726
rect 394 -1837 395 -1795
rect 460 -1796 461 -1726
rect 520 -1796 521 -1726
rect 1206 -1796 1207 -1726
rect 184 -1837 185 -1797
rect 219 -1798 220 -1726
rect 233 -1837 234 -1797
rect 450 -1798 451 -1726
rect 520 -1837 521 -1797
rect 943 -1798 944 -1726
rect 65 -1800 66 -1726
rect 219 -1837 220 -1799
rect 247 -1800 248 -1726
rect 275 -1837 276 -1799
rect 282 -1837 283 -1799
rect 499 -1800 500 -1726
rect 569 -1800 570 -1726
rect 688 -1837 689 -1799
rect 733 -1837 734 -1799
rect 772 -1837 773 -1799
rect 863 -1837 864 -1799
rect 954 -1800 955 -1726
rect 40 -1837 41 -1801
rect 65 -1837 66 -1801
rect 191 -1802 192 -1726
rect 1206 -1837 1207 -1801
rect 114 -1837 115 -1803
rect 191 -1837 192 -1803
rect 198 -1804 199 -1726
rect 303 -1837 304 -1803
rect 338 -1804 339 -1726
rect 450 -1837 451 -1803
rect 569 -1837 570 -1803
rect 695 -1804 696 -1726
rect 737 -1804 738 -1726
rect 870 -1837 871 -1803
rect 135 -1806 136 -1726
rect 198 -1837 199 -1805
rect 247 -1837 248 -1805
rect 254 -1806 255 -1726
rect 261 -1837 262 -1805
rect 492 -1806 493 -1726
rect 583 -1806 584 -1726
rect 954 -1837 955 -1805
rect 135 -1837 136 -1807
rect 163 -1837 164 -1807
rect 254 -1837 255 -1807
rect 387 -1837 388 -1807
rect 443 -1808 444 -1726
rect 499 -1837 500 -1807
rect 583 -1837 584 -1807
rect 758 -1808 759 -1726
rect 761 -1837 762 -1807
rect 877 -1808 878 -1726
rect 296 -1837 297 -1809
rect 716 -1810 717 -1726
rect 751 -1810 752 -1726
rect 1157 -1810 1158 -1726
rect 310 -1837 311 -1811
rect 758 -1837 759 -1811
rect 765 -1837 766 -1811
rect 800 -1812 801 -1726
rect 877 -1837 878 -1811
rect 905 -1812 906 -1726
rect 1024 -1812 1025 -1726
rect 1157 -1837 1158 -1811
rect 338 -1837 339 -1813
rect 352 -1814 353 -1726
rect 366 -1814 367 -1726
rect 492 -1837 493 -1813
rect 618 -1837 619 -1813
rect 653 -1814 654 -1726
rect 674 -1814 675 -1726
rect 800 -1837 801 -1813
rect 905 -1837 906 -1813
rect 961 -1814 962 -1726
rect 1024 -1837 1025 -1813
rect 1080 -1814 1081 -1726
rect 320 -1816 321 -1726
rect 674 -1837 675 -1815
rect 695 -1837 696 -1815
rect 709 -1816 710 -1726
rect 716 -1837 717 -1815
rect 1150 -1837 1151 -1815
rect 352 -1837 353 -1817
rect 754 -1818 755 -1726
rect 961 -1837 962 -1817
rect 1038 -1818 1039 -1726
rect 1080 -1837 1081 -1817
rect 1136 -1818 1137 -1726
rect 366 -1837 367 -1819
rect 429 -1820 430 -1726
rect 443 -1837 444 -1819
rect 604 -1837 605 -1819
rect 607 -1837 608 -1819
rect 1136 -1837 1137 -1819
rect 23 -1837 24 -1821
rect 429 -1837 430 -1821
rect 485 -1837 486 -1821
rect 754 -1837 755 -1821
rect 1038 -1837 1039 -1821
rect 1066 -1822 1067 -1726
rect 422 -1837 423 -1823
rect 709 -1837 710 -1823
rect 737 -1837 738 -1823
rect 751 -1837 752 -1823
rect 1066 -1837 1067 -1823
rect 1129 -1824 1130 -1726
rect 632 -1837 633 -1825
rect 779 -1826 780 -1726
rect 1129 -1837 1130 -1825
rect 1178 -1826 1179 -1726
rect 639 -1837 640 -1827
rect 1125 -1828 1126 -1726
rect 1178 -1837 1179 -1827
rect 1199 -1828 1200 -1726
rect 653 -1837 654 -1829
rect 814 -1837 815 -1829
rect 1199 -1837 1200 -1829
rect 1262 -1830 1263 -1726
rect 558 -1832 559 -1726
rect 1262 -1837 1263 -1831
rect 779 -1837 780 -1833
rect 786 -1834 787 -1726
rect 194 -1836 195 -1726
rect 786 -1837 787 -1835
rect 2 -1847 3 -1845
rect 523 -1960 524 -1846
rect 604 -1847 605 -1845
rect 646 -1847 647 -1845
rect 653 -1847 654 -1845
rect 695 -1847 696 -1845
rect 712 -1847 713 -1845
rect 877 -1847 878 -1845
rect 16 -1849 17 -1845
rect 387 -1849 388 -1845
rect 432 -1960 433 -1848
rect 1010 -1849 1011 -1845
rect 9 -1851 10 -1845
rect 16 -1960 17 -1850
rect 23 -1851 24 -1845
rect 30 -1851 31 -1845
rect 37 -1851 38 -1845
rect 1178 -1851 1179 -1845
rect 9 -1960 10 -1852
rect 79 -1853 80 -1845
rect 89 -1960 90 -1852
rect 247 -1853 248 -1845
rect 254 -1853 255 -1845
rect 366 -1853 367 -1845
rect 373 -1853 374 -1845
rect 373 -1960 374 -1852
rect 373 -1853 374 -1845
rect 373 -1960 374 -1852
rect 387 -1960 388 -1852
rect 555 -1853 556 -1845
rect 558 -1960 559 -1852
rect 653 -1960 654 -1852
rect 656 -1853 657 -1845
rect 891 -1853 892 -1845
rect 1178 -1960 1179 -1852
rect 1269 -1853 1270 -1845
rect 23 -1960 24 -1854
rect 93 -1855 94 -1845
rect 103 -1960 104 -1854
rect 1094 -1855 1095 -1845
rect 30 -1960 31 -1856
rect 520 -1857 521 -1845
rect 555 -1960 556 -1856
rect 1052 -1857 1053 -1845
rect 1094 -1960 1095 -1856
rect 1241 -1857 1242 -1845
rect 37 -1960 38 -1858
rect 338 -1859 339 -1845
rect 366 -1960 367 -1858
rect 436 -1859 437 -1845
rect 464 -1859 465 -1845
rect 506 -1859 507 -1845
rect 513 -1960 514 -1858
rect 541 -1859 542 -1845
rect 607 -1859 608 -1845
rect 856 -1859 857 -1845
rect 877 -1960 878 -1858
rect 996 -1859 997 -1845
rect 1052 -1960 1053 -1858
rect 1157 -1859 1158 -1845
rect 40 -1861 41 -1845
rect 289 -1861 290 -1845
rect 296 -1861 297 -1845
rect 467 -1861 468 -1845
rect 478 -1861 479 -1845
rect 632 -1861 633 -1845
rect 639 -1861 640 -1845
rect 765 -1861 766 -1845
rect 856 -1960 857 -1860
rect 1059 -1861 1060 -1845
rect 1157 -1960 1158 -1860
rect 1234 -1861 1235 -1845
rect 44 -1863 45 -1845
rect 1003 -1863 1004 -1845
rect 1115 -1863 1116 -1845
rect 1234 -1960 1235 -1862
rect 44 -1960 45 -1864
rect 96 -1960 97 -1864
rect 114 -1865 115 -1845
rect 233 -1865 234 -1845
rect 254 -1960 255 -1864
rect 324 -1865 325 -1845
rect 331 -1865 332 -1845
rect 331 -1960 332 -1864
rect 331 -1865 332 -1845
rect 331 -1960 332 -1864
rect 408 -1865 409 -1845
rect 464 -1960 465 -1864
rect 471 -1865 472 -1845
rect 478 -1960 479 -1864
rect 485 -1865 486 -1845
rect 485 -1960 486 -1864
rect 485 -1865 486 -1845
rect 485 -1960 486 -1864
rect 492 -1865 493 -1845
rect 705 -1960 706 -1864
rect 719 -1865 720 -1845
rect 947 -1865 948 -1845
rect 996 -1960 997 -1864
rect 1080 -1865 1081 -1845
rect 1115 -1960 1116 -1864
rect 1199 -1865 1200 -1845
rect 47 -1867 48 -1845
rect 919 -1867 920 -1845
rect 933 -1867 934 -1845
rect 1059 -1960 1060 -1866
rect 1080 -1960 1081 -1866
rect 1192 -1867 1193 -1845
rect 79 -1960 80 -1868
rect 415 -1869 416 -1845
rect 429 -1869 430 -1845
rect 639 -1960 640 -1868
rect 646 -1960 647 -1868
rect 926 -1869 927 -1845
rect 933 -1960 934 -1868
rect 1031 -1869 1032 -1845
rect 1143 -1869 1144 -1845
rect 1199 -1960 1200 -1868
rect 93 -1960 94 -1870
rect 100 -1871 101 -1845
rect 114 -1960 115 -1870
rect 562 -1871 563 -1845
rect 597 -1871 598 -1845
rect 607 -1960 608 -1870
rect 614 -1871 615 -1845
rect 842 -1871 843 -1845
rect 891 -1960 892 -1870
rect 922 -1960 923 -1870
rect 926 -1960 927 -1870
rect 1185 -1871 1186 -1845
rect 100 -1960 101 -1872
rect 527 -1873 528 -1845
rect 534 -1873 535 -1845
rect 562 -1960 563 -1872
rect 597 -1960 598 -1872
rect 618 -1873 619 -1845
rect 628 -1873 629 -1845
rect 1031 -1960 1032 -1872
rect 1038 -1873 1039 -1845
rect 1185 -1960 1186 -1872
rect 135 -1875 136 -1845
rect 807 -1875 808 -1845
rect 842 -1960 843 -1874
rect 968 -1875 969 -1845
rect 1164 -1875 1165 -1845
rect 1192 -1960 1193 -1874
rect 135 -1960 136 -1876
rect 1143 -1960 1144 -1876
rect 149 -1879 150 -1845
rect 233 -1960 234 -1878
rect 264 -1960 265 -1878
rect 282 -1879 283 -1845
rect 289 -1960 290 -1878
rect 310 -1879 311 -1845
rect 324 -1960 325 -1878
rect 394 -1879 395 -1845
rect 408 -1960 409 -1878
rect 674 -1879 675 -1845
rect 677 -1960 678 -1878
rect 688 -1879 689 -1845
rect 695 -1960 696 -1878
rect 786 -1879 787 -1845
rect 919 -1960 920 -1878
rect 1010 -1960 1011 -1878
rect 1073 -1879 1074 -1845
rect 1164 -1960 1165 -1878
rect 86 -1881 87 -1845
rect 282 -1960 283 -1880
rect 299 -1881 300 -1845
rect 572 -1960 573 -1880
rect 688 -1960 689 -1880
rect 772 -1881 773 -1845
rect 786 -1960 787 -1880
rect 898 -1881 899 -1845
rect 947 -1960 948 -1880
rect 1101 -1881 1102 -1845
rect 86 -1960 87 -1882
rect 1227 -1883 1228 -1845
rect 149 -1960 150 -1884
rect 198 -1885 199 -1845
rect 226 -1885 227 -1845
rect 625 -1885 626 -1845
rect 730 -1960 731 -1884
rect 828 -1885 829 -1845
rect 863 -1885 864 -1845
rect 1101 -1960 1102 -1884
rect 152 -1887 153 -1845
rect 268 -1887 269 -1845
rect 275 -1887 276 -1845
rect 415 -1960 416 -1886
rect 436 -1960 437 -1886
rect 450 -1887 451 -1845
rect 457 -1887 458 -1845
rect 625 -1960 626 -1886
rect 709 -1887 710 -1845
rect 828 -1960 829 -1886
rect 863 -1960 864 -1886
rect 961 -1887 962 -1845
rect 968 -1960 969 -1886
rect 1108 -1887 1109 -1845
rect 163 -1889 164 -1845
rect 296 -1960 297 -1888
rect 303 -1889 304 -1845
rect 310 -1960 311 -1888
rect 352 -1889 353 -1845
rect 961 -1960 962 -1888
rect 1073 -1960 1074 -1888
rect 1255 -1889 1256 -1845
rect 163 -1960 164 -1890
rect 355 -1891 356 -1845
rect 422 -1891 423 -1845
rect 450 -1960 451 -1890
rect 471 -1960 472 -1890
rect 838 -1960 839 -1890
rect 898 -1960 899 -1890
rect 1087 -1891 1088 -1845
rect 177 -1893 178 -1845
rect 268 -1960 269 -1892
rect 275 -1960 276 -1892
rect 1223 -1960 1224 -1892
rect 177 -1960 178 -1894
rect 212 -1895 213 -1845
rect 285 -1960 286 -1894
rect 1108 -1960 1109 -1894
rect 184 -1897 185 -1845
rect 226 -1960 227 -1896
rect 303 -1960 304 -1896
rect 520 -1960 521 -1896
rect 527 -1960 528 -1896
rect 576 -1897 577 -1845
rect 709 -1960 710 -1896
rect 744 -1897 745 -1845
rect 751 -1897 752 -1845
rect 975 -1897 976 -1845
rect 1066 -1897 1067 -1845
rect 1087 -1960 1088 -1896
rect 128 -1899 129 -1845
rect 184 -1960 185 -1898
rect 198 -1960 199 -1898
rect 205 -1899 206 -1845
rect 212 -1960 213 -1898
rect 219 -1899 220 -1845
rect 345 -1899 346 -1845
rect 352 -1960 353 -1898
rect 380 -1899 381 -1845
rect 422 -1960 423 -1898
rect 443 -1899 444 -1845
rect 618 -1960 619 -1898
rect 737 -1899 738 -1845
rect 807 -1960 808 -1898
rect 912 -1899 913 -1845
rect 1227 -1960 1228 -1898
rect 128 -1960 129 -1900
rect 142 -1901 143 -1845
rect 205 -1960 206 -1900
rect 240 -1901 241 -1845
rect 345 -1960 346 -1900
rect 401 -1901 402 -1845
rect 495 -1960 496 -1900
rect 793 -1901 794 -1845
rect 912 -1960 913 -1900
rect 1045 -1901 1046 -1845
rect 1066 -1960 1067 -1900
rect 1171 -1901 1172 -1845
rect 51 -1903 52 -1845
rect 401 -1960 402 -1902
rect 506 -1960 507 -1902
rect 723 -1903 724 -1845
rect 737 -1960 738 -1902
rect 849 -1903 850 -1845
rect 975 -1960 976 -1902
rect 1136 -1903 1137 -1845
rect 1171 -1960 1172 -1902
rect 1262 -1903 1263 -1845
rect 51 -1960 52 -1904
rect 457 -1960 458 -1904
rect 516 -1905 517 -1845
rect 1003 -1960 1004 -1904
rect 1045 -1960 1046 -1904
rect 1150 -1905 1151 -1845
rect 58 -1907 59 -1845
rect 142 -1960 143 -1906
rect 219 -1960 220 -1906
rect 317 -1907 318 -1845
rect 359 -1907 360 -1845
rect 443 -1960 444 -1906
rect 534 -1960 535 -1906
rect 590 -1907 591 -1845
rect 744 -1960 745 -1906
rect 835 -1907 836 -1845
rect 849 -1960 850 -1906
rect 1024 -1907 1025 -1845
rect 1150 -1960 1151 -1906
rect 1248 -1907 1249 -1845
rect 58 -1960 59 -1908
rect 499 -1909 500 -1845
rect 541 -1960 542 -1908
rect 667 -1909 668 -1845
rect 751 -1960 752 -1908
rect 761 -1909 762 -1845
rect 765 -1960 766 -1908
rect 884 -1909 885 -1845
rect 1024 -1960 1025 -1908
rect 1129 -1909 1130 -1845
rect 65 -1960 66 -1910
rect 793 -1960 794 -1910
rect 835 -1960 836 -1910
rect 1213 -1911 1214 -1845
rect 138 -1913 139 -1845
rect 723 -1960 724 -1912
rect 754 -1913 755 -1845
rect 940 -1913 941 -1845
rect 1213 -1960 1214 -1912
rect 1276 -1913 1277 -1845
rect 138 -1960 139 -1914
rect 156 -1915 157 -1845
rect 191 -1915 192 -1845
rect 499 -1960 500 -1914
rect 548 -1915 549 -1845
rect 632 -1960 633 -1914
rect 667 -1960 668 -1914
rect 702 -1915 703 -1845
rect 758 -1915 759 -1845
rect 779 -1915 780 -1845
rect 156 -1960 157 -1916
rect 481 -1917 482 -1845
rect 548 -1960 549 -1916
rect 642 -1917 643 -1845
rect 702 -1960 703 -1916
rect 1038 -1960 1039 -1916
rect 191 -1960 192 -1918
rect 369 -1919 370 -1845
rect 380 -1960 381 -1918
rect 604 -1960 605 -1918
rect 761 -1960 762 -1918
rect 884 -1960 885 -1918
rect 72 -1921 73 -1845
rect 369 -1960 370 -1920
rect 429 -1960 430 -1920
rect 1136 -1960 1137 -1920
rect 68 -1923 69 -1845
rect 72 -1960 73 -1922
rect 240 -1960 241 -1922
rect 261 -1923 262 -1845
rect 317 -1960 318 -1922
rect 338 -1960 339 -1922
rect 359 -1960 360 -1922
rect 583 -1923 584 -1845
rect 590 -1960 591 -1922
rect 660 -1923 661 -1845
rect 772 -1960 773 -1922
rect 989 -1923 990 -1845
rect 54 -1925 55 -1845
rect 68 -1960 69 -1924
rect 107 -1925 108 -1845
rect 261 -1960 262 -1924
rect 320 -1960 321 -1924
rect 660 -1960 661 -1924
rect 779 -1960 780 -1924
rect 821 -1925 822 -1845
rect 107 -1960 108 -1926
rect 121 -1927 122 -1845
rect 247 -1960 248 -1926
rect 758 -1960 759 -1926
rect 821 -1960 822 -1926
rect 954 -1927 955 -1845
rect 121 -1960 122 -1928
rect 170 -1929 171 -1845
rect 460 -1960 461 -1928
rect 1129 -1960 1130 -1928
rect 170 -1960 171 -1930
rect 394 -1960 395 -1930
rect 492 -1960 493 -1930
rect 989 -1960 990 -1930
rect 569 -1933 570 -1845
rect 583 -1960 584 -1932
rect 954 -1960 955 -1932
rect 1220 -1933 1221 -1845
rect 569 -1960 570 -1934
rect 940 -1960 941 -1934
rect 576 -1960 577 -1936
rect 814 -1937 815 -1845
rect 814 -1960 815 -1938
rect 870 -1939 871 -1845
rect 870 -1960 871 -1940
rect 982 -1941 983 -1845
rect 611 -1943 612 -1845
rect 982 -1960 983 -1942
rect 611 -1960 612 -1944
rect 681 -1945 682 -1845
rect 681 -1960 682 -1946
rect 716 -1947 717 -1845
rect 716 -1960 717 -1948
rect 800 -1949 801 -1845
rect 800 -1960 801 -1950
rect 905 -1951 906 -1845
rect 905 -1960 906 -1952
rect 1017 -1953 1018 -1845
rect 1017 -1960 1018 -1954
rect 1122 -1955 1123 -1845
rect 1122 -1960 1123 -1956
rect 1206 -1957 1207 -1845
rect 586 -1959 587 -1845
rect 1206 -1960 1207 -1958
rect 2 -2063 3 -1969
rect 646 -1970 647 -1968
rect 674 -1970 675 -1968
rect 954 -1970 955 -1968
rect 964 -1970 965 -1968
rect 1094 -1970 1095 -1968
rect 1157 -1970 1158 -1968
rect 1157 -2063 1158 -1969
rect 1157 -1970 1158 -1968
rect 1157 -2063 1158 -1969
rect 1164 -1970 1165 -1968
rect 1220 -1970 1221 -1968
rect 9 -1972 10 -1968
rect 135 -1972 136 -1968
rect 142 -1972 143 -1968
rect 285 -1972 286 -1968
rect 310 -1972 311 -1968
rect 317 -1972 318 -1968
rect 320 -1972 321 -1968
rect 331 -1972 332 -1968
rect 373 -1972 374 -1968
rect 376 -2000 377 -1971
rect 401 -1972 402 -1968
rect 674 -2063 675 -1971
rect 702 -1972 703 -1968
rect 1101 -1972 1102 -1968
rect 9 -2063 10 -1973
rect 166 -2063 167 -1973
rect 184 -1974 185 -1968
rect 492 -1974 493 -1968
rect 499 -1974 500 -1968
rect 621 -2063 622 -1973
rect 702 -2063 703 -1973
rect 737 -1974 738 -1968
rect 758 -1974 759 -1968
rect 1087 -1974 1088 -1968
rect 1094 -2063 1095 -1973
rect 1136 -1974 1137 -1968
rect 16 -1976 17 -1968
rect 261 -1976 262 -1968
rect 282 -1976 283 -1968
rect 457 -1976 458 -1968
rect 464 -1976 465 -1968
rect 492 -2063 493 -1975
rect 499 -2063 500 -1975
rect 1213 -1976 1214 -1968
rect 37 -1978 38 -1968
rect 173 -1978 174 -1968
rect 184 -2063 185 -1977
rect 324 -1978 325 -1968
rect 331 -2063 332 -1977
rect 394 -1978 395 -1968
rect 408 -1978 409 -1968
rect 411 -2000 412 -1977
rect 464 -2063 465 -1977
rect 541 -1978 542 -1968
rect 569 -1978 570 -1968
rect 716 -1978 717 -1968
rect 737 -2063 738 -1977
rect 891 -1978 892 -1968
rect 919 -1978 920 -1968
rect 996 -1978 997 -1968
rect 1027 -2063 1028 -1977
rect 1192 -1978 1193 -1968
rect 37 -2063 38 -1979
rect 163 -1980 164 -1968
rect 191 -1980 192 -1968
rect 369 -1980 370 -1968
rect 373 -2063 374 -1979
rect 394 -2063 395 -1979
rect 688 -1980 689 -1968
rect 716 -2063 717 -1979
rect 800 -1980 801 -1968
rect 891 -2063 892 -1979
rect 933 -1980 934 -1968
rect 954 -2063 955 -1979
rect 961 -1980 962 -1968
rect 968 -1980 969 -1968
rect 971 -1980 972 -1968
rect 996 -2063 997 -1979
rect 1122 -1980 1123 -1968
rect 16 -2063 17 -1981
rect 163 -2063 164 -1981
rect 198 -1982 199 -1968
rect 429 -1982 430 -1968
rect 481 -2063 482 -1981
rect 1010 -1982 1011 -1968
rect 1073 -1982 1074 -1968
rect 1122 -2063 1123 -1981
rect 51 -1984 52 -1968
rect 240 -1984 241 -1968
rect 243 -2063 244 -1983
rect 688 -2063 689 -1983
rect 758 -2063 759 -1983
rect 786 -1984 787 -1968
rect 800 -2063 801 -1983
rect 842 -1984 843 -1968
rect 919 -2063 920 -1983
rect 940 -1984 941 -1968
rect 968 -2063 969 -1983
rect 975 -1984 976 -1968
rect 1010 -2063 1011 -1983
rect 1143 -1984 1144 -1968
rect 54 -1986 55 -1968
rect 744 -1986 745 -1968
rect 761 -1986 762 -1968
rect 989 -1986 990 -1968
rect 1059 -1986 1060 -1968
rect 1143 -2063 1144 -1985
rect 58 -1988 59 -1968
rect 457 -2063 458 -1987
rect 488 -2063 489 -1987
rect 772 -1988 773 -1968
rect 786 -2063 787 -1987
rect 870 -1988 871 -1968
rect 940 -2063 941 -1987
rect 947 -1988 948 -1968
rect 982 -1988 983 -1968
rect 1059 -2063 1060 -1987
rect 1073 -2063 1074 -1987
rect 1108 -1988 1109 -1968
rect 58 -2063 59 -1989
rect 366 -1990 367 -1968
rect 408 -2063 409 -1989
rect 415 -1990 416 -1968
rect 429 -2063 430 -1989
rect 478 -1990 479 -1968
rect 502 -2063 503 -1989
rect 646 -2063 647 -1989
rect 677 -1990 678 -1968
rect 961 -2063 962 -1989
rect 982 -2063 983 -1989
rect 1045 -1990 1046 -1968
rect 1087 -2063 1088 -1989
rect 1227 -1990 1228 -1968
rect 65 -1992 66 -1968
rect 96 -1992 97 -1968
rect 100 -2063 101 -1991
rect 289 -1992 290 -1968
rect 310 -2063 311 -1991
rect 597 -1992 598 -1968
rect 604 -1992 605 -1968
rect 1199 -1992 1200 -1968
rect 23 -1994 24 -1968
rect 96 -2063 97 -1993
rect 110 -2063 111 -1993
rect 485 -1994 486 -1968
rect 513 -1994 514 -1968
rect 558 -1994 559 -1968
rect 569 -2063 570 -1993
rect 611 -1994 612 -1968
rect 744 -2063 745 -1993
rect 835 -1994 836 -1968
rect 842 -2063 843 -1993
rect 1017 -1994 1018 -1968
rect 1101 -2063 1102 -1993
rect 1171 -1994 1172 -1968
rect 23 -2063 24 -1995
rect 506 -1996 507 -1968
rect 520 -1996 521 -1968
rect 898 -1996 899 -1968
rect 947 -2063 948 -1995
rect 1003 -1996 1004 -1968
rect 1017 -2063 1018 -1995
rect 1066 -1996 1067 -1968
rect 1108 -2063 1109 -1995
rect 1178 -1996 1179 -1968
rect 44 -1998 45 -1968
rect 65 -2063 66 -1997
rect 68 -1998 69 -1968
rect 730 -1998 731 -1968
rect 772 -2063 773 -1997
rect 838 -1998 839 -1968
rect 849 -1998 850 -1968
rect 870 -2063 871 -1997
rect 898 -2063 899 -1997
rect 1038 -1998 1039 -1968
rect 1066 -2063 1067 -1997
rect 1080 -1998 1081 -1968
rect 72 -2000 73 -1968
rect 663 -2063 664 -1999
rect 835 -2063 836 -1999
rect 877 -2000 878 -1968
rect 971 -2063 972 -1999
rect 975 -2063 976 -1999
rect 989 -2063 990 -1999
rect 1024 -2000 1025 -1968
rect 1031 -2000 1032 -1968
rect 1038 -2063 1039 -1999
rect 1080 -2063 1081 -1999
rect 1115 -2000 1116 -1968
rect 72 -2063 73 -2001
rect 107 -2002 108 -1968
rect 114 -2002 115 -1968
rect 366 -2063 367 -2001
rect 478 -2063 479 -2001
rect 730 -2063 731 -2001
rect 877 -2063 878 -2001
rect 884 -2002 885 -1968
rect 1003 -2063 1004 -2001
rect 1052 -2002 1053 -1968
rect 1115 -2063 1116 -2001
rect 1206 -2002 1207 -1968
rect 86 -2004 87 -1968
rect 135 -2063 136 -2003
rect 142 -2063 143 -2003
rect 268 -2004 269 -1968
rect 282 -2063 283 -2003
rect 450 -2004 451 -1968
rect 506 -2063 507 -2003
rect 698 -2063 699 -2003
rect 926 -2004 927 -1968
rect 1052 -2063 1053 -2003
rect 86 -2063 87 -2005
rect 562 -2006 563 -1968
rect 576 -2006 577 -1968
rect 884 -2063 885 -2005
rect 1031 -2063 1032 -2005
rect 1150 -2006 1151 -1968
rect 44 -2063 45 -2007
rect 576 -2063 577 -2007
rect 579 -2063 580 -2007
rect 814 -2008 815 -1968
rect 856 -2008 857 -1968
rect 926 -2063 927 -2007
rect 1136 -2063 1137 -2007
rect 1150 -2063 1151 -2007
rect 51 -2063 52 -2009
rect 814 -2063 815 -2009
rect 856 -2063 857 -2009
rect 905 -2010 906 -1968
rect 89 -2012 90 -1968
rect 107 -2063 108 -2011
rect 117 -2063 118 -2011
rect 212 -2012 213 -1968
rect 226 -2012 227 -1968
rect 278 -2063 279 -2011
rect 317 -2063 318 -2011
rect 345 -2012 346 -1968
rect 450 -2063 451 -2011
rect 471 -2012 472 -1968
rect 534 -2012 535 -1968
rect 933 -2063 934 -2011
rect 93 -2014 94 -1968
rect 709 -2014 710 -1968
rect 905 -2063 906 -2013
rect 912 -2014 913 -1968
rect 93 -2063 94 -2015
rect 303 -2016 304 -1968
rect 338 -2016 339 -1968
rect 604 -2063 605 -2015
rect 611 -2063 612 -2015
rect 625 -2016 626 -1968
rect 709 -2063 710 -2015
rect 765 -2016 766 -1968
rect 30 -2018 31 -1968
rect 303 -2063 304 -2017
rect 471 -2063 472 -2017
rect 548 -2018 549 -1968
rect 562 -2063 563 -2017
rect 681 -2018 682 -1968
rect 751 -2018 752 -1968
rect 912 -2063 913 -2017
rect 30 -2063 31 -2019
rect 359 -2020 360 -1968
rect 534 -2063 535 -2019
rect 590 -2020 591 -1968
rect 597 -2063 598 -2019
rect 632 -2020 633 -1968
rect 681 -2063 682 -2019
rect 695 -2020 696 -1968
rect 751 -2063 752 -2019
rect 779 -2020 780 -1968
rect 114 -2063 115 -2021
rect 338 -2063 339 -2021
rect 432 -2022 433 -1968
rect 590 -2063 591 -2021
rect 625 -2063 626 -2021
rect 660 -2022 661 -1968
rect 765 -2063 766 -2021
rect 821 -2022 822 -1968
rect 121 -2024 122 -1968
rect 520 -2063 521 -2023
rect 541 -2063 542 -2023
rect 583 -2024 584 -1968
rect 632 -2063 633 -2023
rect 639 -2024 640 -1968
rect 660 -2063 661 -2023
rect 667 -2024 668 -1968
rect 821 -2063 822 -2023
rect 863 -2024 864 -1968
rect 103 -2026 104 -1968
rect 667 -2063 668 -2025
rect 863 -2063 864 -2025
rect 1185 -2026 1186 -1968
rect 121 -2063 122 -2027
rect 653 -2028 654 -1968
rect 1185 -2063 1186 -2027
rect 1234 -2028 1235 -1968
rect 128 -2030 129 -1968
rect 572 -2030 573 -1968
rect 583 -2063 584 -2029
rect 779 -2063 780 -2029
rect 152 -2063 153 -2031
rect 849 -2063 850 -2031
rect 170 -2034 171 -1968
rect 345 -2063 346 -2033
rect 548 -2063 549 -2033
rect 618 -2034 619 -1968
rect 639 -2063 640 -2033
rect 1024 -2063 1025 -2033
rect 149 -2036 150 -1968
rect 170 -2063 171 -2035
rect 177 -2036 178 -1968
rect 212 -2063 213 -2035
rect 226 -2063 227 -2035
rect 275 -2036 276 -1968
rect 618 -2063 619 -2035
rect 1045 -2063 1046 -2035
rect 128 -2063 129 -2037
rect 149 -2063 150 -2037
rect 177 -2063 178 -2037
rect 695 -2063 696 -2037
rect 191 -2063 192 -2039
rect 240 -2063 241 -2039
rect 247 -2040 248 -1968
rect 513 -2063 514 -2039
rect 653 -2063 654 -2039
rect 807 -2040 808 -1968
rect 198 -2063 199 -2041
rect 387 -2042 388 -1968
rect 807 -2063 808 -2041
rect 828 -2042 829 -1968
rect 205 -2044 206 -1968
rect 261 -2063 262 -2043
rect 268 -2063 269 -2043
rect 352 -2044 353 -1968
rect 828 -2063 829 -2043
rect 1129 -2044 1130 -1968
rect 156 -2046 157 -1968
rect 205 -2063 206 -2045
rect 233 -2046 234 -1968
rect 359 -2063 360 -2045
rect 723 -2046 724 -1968
rect 1129 -2063 1130 -2045
rect 79 -2048 80 -1968
rect 156 -2063 157 -2047
rect 233 -2063 234 -2047
rect 523 -2048 524 -1968
rect 723 -2063 724 -2047
rect 793 -2048 794 -1968
rect 79 -2063 80 -2049
rect 334 -2063 335 -2049
rect 352 -2063 353 -2049
rect 422 -2050 423 -1968
rect 555 -2050 556 -1968
rect 793 -2063 794 -2049
rect 247 -2063 248 -2051
rect 460 -2052 461 -1968
rect 555 -2063 556 -2051
rect 1223 -2052 1224 -1968
rect 254 -2054 255 -1968
rect 289 -2063 290 -2053
rect 296 -2054 297 -1968
rect 387 -2063 388 -2053
rect 422 -2063 423 -2053
rect 527 -2054 528 -1968
rect 138 -2056 139 -1968
rect 296 -2063 297 -2055
rect 436 -2056 437 -1968
rect 527 -2063 528 -2055
rect 219 -2058 220 -1968
rect 254 -2063 255 -2057
rect 275 -2063 276 -2057
rect 401 -2063 402 -2057
rect 436 -2063 437 -2057
rect 443 -2058 444 -1968
rect 89 -2063 90 -2059
rect 443 -2063 444 -2059
rect 219 -2063 220 -2061
rect 607 -2062 608 -1968
rect 2 -2073 3 -2071
rect 93 -2073 94 -2071
rect 103 -2148 104 -2072
rect 744 -2073 745 -2071
rect 789 -2148 790 -2072
rect 1122 -2073 1123 -2071
rect 1136 -2073 1137 -2071
rect 1185 -2073 1186 -2071
rect 30 -2075 31 -2071
rect 243 -2075 244 -2071
rect 247 -2075 248 -2071
rect 278 -2075 279 -2071
rect 394 -2075 395 -2071
rect 618 -2075 619 -2071
rect 621 -2075 622 -2071
rect 800 -2075 801 -2071
rect 817 -2075 818 -2071
rect 975 -2075 976 -2071
rect 1010 -2075 1011 -2071
rect 1010 -2148 1011 -2074
rect 1010 -2075 1011 -2071
rect 1010 -2148 1011 -2074
rect 1108 -2075 1109 -2071
rect 1108 -2148 1109 -2074
rect 1108 -2075 1109 -2071
rect 1108 -2148 1109 -2074
rect 1122 -2148 1123 -2074
rect 1150 -2075 1151 -2071
rect 30 -2148 31 -2076
rect 86 -2077 87 -2071
rect 93 -2148 94 -2076
rect 163 -2077 164 -2071
rect 166 -2077 167 -2071
rect 996 -2077 997 -2071
rect 1139 -2077 1140 -2071
rect 1157 -2077 1158 -2071
rect 37 -2079 38 -2071
rect 324 -2079 325 -2071
rect 394 -2148 395 -2078
rect 471 -2079 472 -2071
rect 481 -2079 482 -2071
rect 527 -2079 528 -2071
rect 562 -2079 563 -2071
rect 565 -2087 566 -2078
rect 576 -2079 577 -2071
rect 877 -2079 878 -2071
rect 975 -2148 976 -2078
rect 1038 -2079 1039 -2071
rect 65 -2081 66 -2071
rect 152 -2081 153 -2071
rect 156 -2081 157 -2071
rect 499 -2081 500 -2071
rect 509 -2148 510 -2080
rect 639 -2081 640 -2071
rect 653 -2148 654 -2080
rect 1024 -2148 1025 -2080
rect 65 -2148 66 -2082
rect 296 -2083 297 -2071
rect 387 -2083 388 -2071
rect 481 -2148 482 -2082
rect 492 -2083 493 -2071
rect 530 -2148 531 -2082
rect 562 -2148 563 -2082
rect 590 -2083 591 -2071
rect 600 -2148 601 -2082
rect 632 -2083 633 -2071
rect 639 -2148 640 -2082
rect 884 -2083 885 -2071
rect 72 -2085 73 -2071
rect 72 -2148 73 -2084
rect 72 -2085 73 -2071
rect 72 -2148 73 -2084
rect 86 -2148 87 -2084
rect 135 -2085 136 -2071
rect 138 -2148 139 -2084
rect 793 -2085 794 -2071
rect 863 -2085 864 -2071
rect 1087 -2085 1088 -2071
rect 37 -2148 38 -2086
rect 135 -2148 136 -2086
rect 142 -2087 143 -2071
rect 488 -2087 489 -2071
rect 590 -2148 591 -2086
rect 614 -2148 615 -2086
rect 996 -2148 997 -2086
rect 100 -2089 101 -2071
rect 247 -2148 248 -2088
rect 254 -2089 255 -2071
rect 299 -2148 300 -2088
rect 387 -2148 388 -2088
rect 450 -2089 451 -2071
rect 457 -2089 458 -2071
rect 499 -2148 500 -2088
rect 576 -2148 577 -2088
rect 625 -2089 626 -2071
rect 632 -2148 633 -2088
rect 667 -2089 668 -2071
rect 695 -2089 696 -2071
rect 758 -2089 759 -2071
rect 793 -2148 794 -2088
rect 1129 -2089 1130 -2071
rect 100 -2148 101 -2090
rect 163 -2148 164 -2090
rect 170 -2091 171 -2071
rect 240 -2091 241 -2071
rect 254 -2148 255 -2090
rect 289 -2091 290 -2071
rect 401 -2091 402 -2071
rect 492 -2148 493 -2090
rect 579 -2091 580 -2071
rect 611 -2091 612 -2071
rect 618 -2148 619 -2090
rect 674 -2091 675 -2071
rect 695 -2148 696 -2090
rect 947 -2091 948 -2071
rect 107 -2093 108 -2071
rect 114 -2093 115 -2071
rect 117 -2093 118 -2071
rect 282 -2093 283 -2071
rect 289 -2148 290 -2092
rect 303 -2093 304 -2071
rect 401 -2148 402 -2092
rect 464 -2093 465 -2071
rect 467 -2148 468 -2092
rect 1038 -2148 1039 -2092
rect 58 -2095 59 -2071
rect 107 -2148 108 -2094
rect 114 -2148 115 -2094
rect 380 -2095 381 -2071
rect 429 -2095 430 -2071
rect 450 -2148 451 -2094
rect 457 -2148 458 -2094
rect 646 -2095 647 -2071
rect 656 -2148 657 -2094
rect 709 -2095 710 -2071
rect 716 -2095 717 -2071
rect 800 -2148 801 -2094
rect 863 -2148 864 -2094
rect 926 -2095 927 -2071
rect 947 -2148 948 -2094
rect 1101 -2095 1102 -2071
rect 23 -2097 24 -2071
rect 58 -2148 59 -2096
rect 142 -2148 143 -2096
rect 233 -2097 234 -2071
rect 240 -2148 241 -2096
rect 334 -2097 335 -2071
rect 373 -2097 374 -2071
rect 380 -2148 381 -2096
rect 408 -2097 409 -2071
rect 646 -2148 647 -2096
rect 660 -2097 661 -2071
rect 842 -2097 843 -2071
rect 877 -2148 878 -2096
rect 954 -2097 955 -2071
rect 23 -2148 24 -2098
rect 89 -2099 90 -2071
rect 96 -2148 97 -2098
rect 373 -2148 374 -2098
rect 429 -2148 430 -2098
rect 436 -2099 437 -2071
rect 443 -2099 444 -2071
rect 611 -2148 612 -2098
rect 625 -2148 626 -2098
rect 688 -2099 689 -2071
rect 709 -2148 710 -2098
rect 807 -2099 808 -2071
rect 842 -2148 843 -2098
rect 891 -2099 892 -2071
rect 926 -2148 927 -2098
rect 982 -2099 983 -2071
rect 149 -2101 150 -2071
rect 485 -2101 486 -2071
rect 583 -2101 584 -2071
rect 912 -2101 913 -2071
rect 933 -2101 934 -2071
rect 954 -2148 955 -2100
rect 982 -2148 983 -2100
rect 1066 -2101 1067 -2071
rect 44 -2103 45 -2071
rect 149 -2148 150 -2102
rect 156 -2148 157 -2102
rect 219 -2103 220 -2071
rect 233 -2148 234 -2102
rect 317 -2103 318 -2071
rect 345 -2103 346 -2071
rect 408 -2148 409 -2102
rect 443 -2148 444 -2102
rect 691 -2148 692 -2102
rect 716 -2148 717 -2102
rect 772 -2103 773 -2071
rect 807 -2148 808 -2102
rect 821 -2103 822 -2071
rect 884 -2148 885 -2102
rect 961 -2103 962 -2071
rect 1066 -2148 1067 -2102
rect 1080 -2103 1081 -2071
rect 44 -2148 45 -2104
rect 698 -2105 699 -2071
rect 737 -2105 738 -2071
rect 758 -2148 759 -2104
rect 772 -2148 773 -2104
rect 786 -2105 787 -2071
rect 821 -2148 822 -2104
rect 905 -2105 906 -2071
rect 933 -2148 934 -2104
rect 1017 -2105 1018 -2071
rect 51 -2107 52 -2071
rect 219 -2148 220 -2106
rect 261 -2107 262 -2071
rect 320 -2148 321 -2106
rect 338 -2107 339 -2071
rect 961 -2148 962 -2106
rect 1017 -2148 1018 -2106
rect 1115 -2107 1116 -2071
rect 16 -2109 17 -2071
rect 51 -2148 52 -2108
rect 173 -2148 174 -2108
rect 681 -2109 682 -2071
rect 737 -2148 738 -2108
rect 765 -2109 766 -2071
rect 891 -2148 892 -2108
rect 968 -2109 969 -2071
rect 110 -2111 111 -2071
rect 765 -2148 766 -2110
rect 898 -2111 899 -2071
rect 912 -2148 913 -2110
rect 968 -2148 969 -2110
rect 1031 -2111 1032 -2071
rect 184 -2113 185 -2071
rect 282 -2148 283 -2112
rect 303 -2148 304 -2112
rect 516 -2148 517 -2112
rect 583 -2148 584 -2112
rect 597 -2113 598 -2071
rect 660 -2148 661 -2112
rect 663 -2113 664 -2071
rect 667 -2148 668 -2112
rect 702 -2113 703 -2071
rect 744 -2148 745 -2112
rect 751 -2113 752 -2071
rect 814 -2113 815 -2071
rect 898 -2148 899 -2112
rect 905 -2148 906 -2112
rect 1059 -2113 1060 -2071
rect 184 -2148 185 -2114
rect 534 -2115 535 -2071
rect 674 -2148 675 -2114
rect 723 -2115 724 -2071
rect 751 -2148 752 -2114
rect 779 -2115 780 -2071
rect 814 -2148 815 -2114
rect 856 -2115 857 -2071
rect 866 -2115 867 -2071
rect 1059 -2148 1060 -2114
rect 205 -2117 206 -2071
rect 324 -2148 325 -2116
rect 338 -2148 339 -2116
rect 502 -2117 503 -2071
rect 681 -2148 682 -2116
rect 849 -2117 850 -2071
rect 856 -2148 857 -2116
rect 1003 -2117 1004 -2071
rect 1031 -2148 1032 -2116
rect 1104 -2148 1105 -2116
rect 205 -2148 206 -2118
rect 226 -2119 227 -2071
rect 261 -2148 262 -2118
rect 527 -2148 528 -2118
rect 702 -2148 703 -2118
rect 870 -2119 871 -2071
rect 1003 -2148 1004 -2118
rect 1143 -2119 1144 -2071
rect 79 -2121 80 -2071
rect 226 -2148 227 -2120
rect 268 -2121 269 -2071
rect 331 -2121 332 -2071
rect 345 -2148 346 -2120
rect 422 -2121 423 -2071
rect 471 -2148 472 -2120
rect 548 -2121 549 -2071
rect 723 -2148 724 -2120
rect 835 -2121 836 -2071
rect 849 -2148 850 -2120
rect 1052 -2121 1053 -2071
rect 79 -2148 80 -2122
rect 478 -2123 479 -2071
rect 548 -2148 549 -2122
rect 642 -2148 643 -2122
rect 730 -2123 731 -2071
rect 779 -2148 780 -2122
rect 835 -2148 836 -2122
rect 1045 -2123 1046 -2071
rect 1052 -2148 1053 -2122
rect 1101 -2148 1102 -2122
rect 128 -2125 129 -2071
rect 331 -2148 332 -2124
rect 352 -2125 353 -2071
rect 436 -2148 437 -2124
rect 478 -2148 479 -2124
rect 989 -2125 990 -2071
rect 128 -2148 129 -2126
rect 177 -2127 178 -2071
rect 212 -2127 213 -2071
rect 327 -2127 328 -2071
rect 352 -2148 353 -2126
rect 513 -2127 514 -2071
rect 597 -2148 598 -2126
rect 1045 -2148 1046 -2126
rect 9 -2129 10 -2071
rect 513 -2148 514 -2128
rect 730 -2148 731 -2128
rect 828 -2129 829 -2071
rect 870 -2148 871 -2128
rect 940 -2129 941 -2071
rect 989 -2148 990 -2128
rect 1073 -2129 1074 -2071
rect 177 -2148 178 -2130
rect 191 -2131 192 -2071
rect 212 -2148 213 -2130
rect 359 -2131 360 -2071
rect 366 -2131 367 -2071
rect 422 -2148 423 -2130
rect 485 -2148 486 -2130
rect 940 -2148 941 -2130
rect 121 -2133 122 -2071
rect 191 -2148 192 -2132
rect 268 -2148 269 -2132
rect 506 -2133 507 -2071
rect 828 -2148 829 -2132
rect 919 -2133 920 -2071
rect 117 -2148 118 -2134
rect 121 -2148 122 -2134
rect 275 -2148 276 -2134
rect 555 -2135 556 -2071
rect 919 -2148 920 -2134
rect 1094 -2135 1095 -2071
rect 310 -2137 311 -2071
rect 534 -2148 535 -2136
rect 555 -2148 556 -2136
rect 569 -2137 570 -2071
rect 198 -2139 199 -2071
rect 310 -2148 311 -2138
rect 359 -2148 360 -2138
rect 415 -2139 416 -2071
rect 464 -2148 465 -2138
rect 569 -2148 570 -2138
rect 198 -2148 199 -2140
rect 317 -2148 318 -2140
rect 366 -2148 367 -2140
rect 520 -2141 521 -2071
rect 415 -2148 416 -2142
rect 604 -2143 605 -2071
rect 520 -2148 521 -2144
rect 541 -2145 542 -2071
rect 604 -2148 605 -2144
rect 688 -2148 689 -2144
rect 541 -2148 542 -2146
rect 786 -2148 787 -2146
rect 23 -2158 24 -2156
rect 117 -2158 118 -2156
rect 124 -2229 125 -2157
rect 303 -2158 304 -2156
rect 317 -2229 318 -2157
rect 324 -2158 325 -2156
rect 331 -2158 332 -2156
rect 971 -2158 972 -2156
rect 975 -2158 976 -2156
rect 996 -2158 997 -2156
rect 1066 -2158 1067 -2156
rect 1066 -2229 1067 -2157
rect 1066 -2158 1067 -2156
rect 1066 -2229 1067 -2157
rect 1101 -2158 1102 -2156
rect 1108 -2158 1109 -2156
rect 37 -2160 38 -2156
rect 100 -2160 101 -2156
rect 103 -2160 104 -2156
rect 156 -2160 157 -2156
rect 198 -2160 199 -2156
rect 303 -2229 304 -2159
rect 324 -2229 325 -2159
rect 380 -2160 381 -2156
rect 387 -2160 388 -2156
rect 488 -2160 489 -2156
rect 509 -2160 510 -2156
rect 849 -2160 850 -2156
rect 933 -2160 934 -2156
rect 968 -2229 969 -2159
rect 982 -2160 983 -2156
rect 996 -2229 997 -2159
rect 1104 -2160 1105 -2156
rect 1122 -2160 1123 -2156
rect 37 -2229 38 -2161
rect 86 -2162 87 -2156
rect 93 -2162 94 -2156
rect 261 -2162 262 -2156
rect 275 -2162 276 -2156
rect 464 -2162 465 -2156
rect 485 -2162 486 -2156
rect 583 -2162 584 -2156
rect 597 -2162 598 -2156
rect 702 -2162 703 -2156
rect 786 -2162 787 -2156
rect 898 -2162 899 -2156
rect 933 -2229 934 -2161
rect 1038 -2162 1039 -2156
rect 30 -2164 31 -2156
rect 93 -2229 94 -2163
rect 100 -2229 101 -2163
rect 142 -2164 143 -2156
rect 198 -2229 199 -2163
rect 247 -2164 248 -2156
rect 254 -2164 255 -2156
rect 467 -2164 468 -2156
rect 513 -2164 514 -2156
rect 695 -2164 696 -2156
rect 702 -2229 703 -2163
rect 737 -2164 738 -2156
rect 786 -2229 787 -2163
rect 884 -2164 885 -2156
rect 943 -2229 944 -2163
rect 1059 -2164 1060 -2156
rect 30 -2229 31 -2165
rect 527 -2166 528 -2156
rect 597 -2229 598 -2165
rect 632 -2166 633 -2156
rect 639 -2229 640 -2165
rect 674 -2166 675 -2156
rect 688 -2166 689 -2156
rect 919 -2166 920 -2156
rect 982 -2229 983 -2165
rect 1003 -2166 1004 -2156
rect 51 -2168 52 -2156
rect 156 -2229 157 -2167
rect 226 -2168 227 -2156
rect 226 -2229 227 -2167
rect 226 -2168 227 -2156
rect 226 -2229 227 -2167
rect 233 -2168 234 -2156
rect 478 -2168 479 -2156
rect 513 -2229 514 -2167
rect 541 -2168 542 -2156
rect 611 -2168 612 -2156
rect 954 -2168 955 -2156
rect 1003 -2229 1004 -2167
rect 1052 -2168 1053 -2156
rect 44 -2170 45 -2156
rect 51 -2229 52 -2169
rect 65 -2170 66 -2156
rect 261 -2229 262 -2169
rect 289 -2170 290 -2156
rect 488 -2229 489 -2169
rect 541 -2229 542 -2169
rect 569 -2170 570 -2156
rect 611 -2229 612 -2169
rect 698 -2229 699 -2169
rect 842 -2170 843 -2156
rect 975 -2229 976 -2169
rect 58 -2172 59 -2156
rect 65 -2229 66 -2171
rect 72 -2172 73 -2156
rect 135 -2172 136 -2156
rect 138 -2172 139 -2156
rect 583 -2229 584 -2171
rect 614 -2172 615 -2156
rect 898 -2229 899 -2171
rect 919 -2229 920 -2171
rect 1031 -2172 1032 -2156
rect 58 -2229 59 -2173
rect 397 -2229 398 -2173
rect 408 -2174 409 -2156
rect 481 -2229 482 -2173
rect 632 -2229 633 -2173
rect 709 -2174 710 -2156
rect 842 -2229 843 -2173
rect 961 -2174 962 -2156
rect 72 -2229 73 -2175
rect 184 -2176 185 -2156
rect 240 -2176 241 -2156
rect 247 -2229 248 -2175
rect 254 -2229 255 -2175
rect 268 -2176 269 -2156
rect 289 -2229 290 -2175
rect 394 -2176 395 -2156
rect 401 -2176 402 -2156
rect 408 -2229 409 -2175
rect 429 -2176 430 -2156
rect 506 -2176 507 -2156
rect 646 -2176 647 -2156
rect 884 -2229 885 -2175
rect 96 -2178 97 -2156
rect 184 -2229 185 -2177
rect 205 -2178 206 -2156
rect 240 -2229 241 -2177
rect 268 -2229 269 -2177
rect 789 -2178 790 -2156
rect 96 -2229 97 -2179
rect 656 -2180 657 -2156
rect 674 -2229 675 -2179
rect 681 -2180 682 -2156
rect 688 -2229 689 -2179
rect 765 -2180 766 -2156
rect 114 -2182 115 -2156
rect 275 -2229 276 -2181
rect 296 -2182 297 -2156
rect 331 -2229 332 -2181
rect 355 -2229 356 -2181
rect 604 -2182 605 -2156
rect 646 -2229 647 -2181
rect 667 -2182 668 -2156
rect 681 -2229 682 -2181
rect 758 -2182 759 -2156
rect 114 -2229 115 -2183
rect 121 -2184 122 -2156
rect 131 -2229 132 -2183
rect 359 -2184 360 -2156
rect 366 -2184 367 -2156
rect 394 -2229 395 -2183
rect 401 -2229 402 -2183
rect 450 -2184 451 -2156
rect 464 -2229 465 -2183
rect 499 -2184 500 -2156
rect 506 -2229 507 -2183
rect 555 -2184 556 -2156
rect 604 -2229 605 -2183
rect 747 -2229 748 -2183
rect 751 -2184 752 -2156
rect 961 -2229 962 -2183
rect 121 -2229 122 -2185
rect 443 -2186 444 -2156
rect 457 -2186 458 -2156
rect 555 -2229 556 -2185
rect 656 -2229 657 -2185
rect 856 -2186 857 -2156
rect 135 -2229 136 -2187
rect 219 -2188 220 -2156
rect 282 -2188 283 -2156
rect 296 -2229 297 -2187
rect 310 -2188 311 -2156
rect 366 -2229 367 -2187
rect 373 -2188 374 -2156
rect 429 -2229 430 -2187
rect 443 -2229 444 -2187
rect 492 -2188 493 -2156
rect 499 -2229 500 -2187
rect 530 -2229 531 -2187
rect 691 -2188 692 -2156
rect 800 -2188 801 -2156
rect 856 -2229 857 -2187
rect 905 -2188 906 -2156
rect 79 -2190 80 -2156
rect 282 -2229 283 -2189
rect 310 -2229 311 -2189
rect 352 -2190 353 -2156
rect 359 -2229 360 -2189
rect 548 -2190 549 -2156
rect 695 -2229 696 -2189
rect 1045 -2190 1046 -2156
rect 79 -2229 80 -2191
rect 128 -2192 129 -2156
rect 142 -2229 143 -2191
rect 149 -2192 150 -2156
rect 163 -2192 164 -2156
rect 569 -2229 570 -2191
rect 709 -2229 710 -2191
rect 779 -2192 780 -2156
rect 800 -2229 801 -2191
rect 807 -2192 808 -2156
rect 905 -2229 906 -2191
rect 1024 -2192 1025 -2156
rect 44 -2229 45 -2193
rect 128 -2229 129 -2193
rect 163 -2229 164 -2193
rect 653 -2194 654 -2156
rect 751 -2229 752 -2193
rect 870 -2194 871 -2156
rect 86 -2229 87 -2195
rect 149 -2229 150 -2195
rect 170 -2196 171 -2156
rect 233 -2229 234 -2195
rect 320 -2196 321 -2156
rect 849 -2229 850 -2195
rect 870 -2229 871 -2195
rect 1017 -2196 1018 -2156
rect 170 -2229 171 -2197
rect 177 -2198 178 -2156
rect 180 -2229 181 -2197
rect 492 -2229 493 -2197
rect 548 -2229 549 -2197
rect 590 -2198 591 -2156
rect 653 -2229 654 -2197
rect 772 -2198 773 -2156
rect 779 -2229 780 -2197
rect 821 -2198 822 -2156
rect 954 -2229 955 -2197
rect 1017 -2229 1018 -2197
rect 177 -2229 178 -2199
rect 212 -2200 213 -2156
rect 219 -2229 220 -2199
rect 345 -2200 346 -2156
rect 373 -2229 374 -2199
rect 471 -2200 472 -2156
rect 590 -2229 591 -2199
rect 625 -2200 626 -2156
rect 758 -2229 759 -2199
rect 877 -2200 878 -2156
rect 107 -2202 108 -2156
rect 345 -2229 346 -2201
rect 380 -2229 381 -2201
rect 576 -2202 577 -2156
rect 618 -2202 619 -2156
rect 625 -2229 626 -2201
rect 772 -2229 773 -2201
rect 828 -2202 829 -2156
rect 877 -2229 878 -2201
rect 947 -2202 948 -2156
rect 107 -2229 108 -2203
rect 299 -2204 300 -2156
rect 387 -2229 388 -2203
rect 436 -2204 437 -2156
rect 450 -2229 451 -2203
rect 576 -2229 577 -2203
rect 618 -2229 619 -2203
rect 793 -2204 794 -2156
rect 807 -2229 808 -2203
rect 814 -2204 815 -2156
rect 821 -2229 822 -2203
rect 891 -2204 892 -2156
rect 191 -2206 192 -2156
rect 667 -2229 668 -2205
rect 670 -2229 671 -2205
rect 891 -2229 892 -2205
rect 191 -2229 192 -2207
rect 562 -2208 563 -2156
rect 793 -2229 794 -2207
rect 835 -2208 836 -2156
rect 205 -2229 206 -2209
rect 660 -2210 661 -2156
rect 814 -2229 815 -2209
rect 912 -2210 913 -2156
rect 212 -2229 213 -2211
rect 453 -2229 454 -2211
rect 471 -2229 472 -2211
rect 520 -2212 521 -2156
rect 660 -2229 661 -2211
rect 716 -2212 717 -2156
rect 828 -2229 829 -2211
rect 940 -2212 941 -2156
rect 338 -2214 339 -2156
rect 716 -2229 717 -2213
rect 765 -2229 766 -2213
rect 940 -2229 941 -2213
rect 338 -2229 339 -2215
rect 740 -2229 741 -2215
rect 835 -2229 836 -2215
rect 926 -2216 927 -2156
rect 422 -2218 423 -2156
rect 457 -2229 458 -2217
rect 485 -2229 486 -2217
rect 947 -2229 948 -2217
rect 415 -2220 416 -2156
rect 422 -2229 423 -2219
rect 436 -2229 437 -2219
rect 723 -2220 724 -2156
rect 912 -2229 913 -2219
rect 989 -2220 990 -2156
rect 415 -2229 416 -2221
rect 527 -2229 528 -2221
rect 723 -2229 724 -2221
rect 863 -2222 864 -2156
rect 926 -2229 927 -2221
rect 1010 -2222 1011 -2156
rect 516 -2224 517 -2156
rect 562 -2229 563 -2223
rect 730 -2224 731 -2156
rect 863 -2229 864 -2223
rect 520 -2229 521 -2225
rect 534 -2226 535 -2156
rect 730 -2229 731 -2225
rect 744 -2226 745 -2156
rect 534 -2229 535 -2227
rect 600 -2228 601 -2156
rect 30 -2239 31 -2237
rect 128 -2239 129 -2237
rect 131 -2239 132 -2237
rect 338 -2239 339 -2237
rect 345 -2239 346 -2237
rect 348 -2312 349 -2238
rect 359 -2239 360 -2237
rect 656 -2239 657 -2237
rect 667 -2239 668 -2237
rect 835 -2239 836 -2237
rect 940 -2239 941 -2237
rect 961 -2239 962 -2237
rect 968 -2239 969 -2237
rect 968 -2312 969 -2238
rect 968 -2239 969 -2237
rect 968 -2312 969 -2238
rect 989 -2312 990 -2238
rect 1003 -2239 1004 -2237
rect 1017 -2239 1018 -2237
rect 1038 -2312 1039 -2238
rect 1059 -2312 1060 -2238
rect 1066 -2239 1067 -2237
rect 44 -2241 45 -2237
rect 47 -2259 48 -2240
rect 51 -2241 52 -2237
rect 89 -2241 90 -2237
rect 93 -2241 94 -2237
rect 450 -2241 451 -2237
rect 481 -2241 482 -2237
rect 632 -2241 633 -2237
rect 667 -2312 668 -2240
rect 688 -2241 689 -2237
rect 695 -2312 696 -2240
rect 751 -2241 752 -2237
rect 800 -2241 801 -2237
rect 803 -2312 804 -2240
rect 807 -2241 808 -2237
rect 810 -2241 811 -2237
rect 835 -2312 836 -2240
rect 870 -2241 871 -2237
rect 943 -2241 944 -2237
rect 982 -2241 983 -2237
rect 996 -2241 997 -2237
rect 996 -2312 997 -2240
rect 996 -2241 997 -2237
rect 996 -2312 997 -2240
rect 37 -2243 38 -2237
rect 89 -2312 90 -2242
rect 135 -2243 136 -2237
rect 338 -2312 339 -2242
rect 359 -2312 360 -2242
rect 373 -2243 374 -2237
rect 429 -2243 430 -2237
rect 478 -2243 479 -2237
rect 520 -2243 521 -2237
rect 520 -2312 521 -2242
rect 520 -2243 521 -2237
rect 520 -2312 521 -2242
rect 527 -2243 528 -2237
rect 660 -2243 661 -2237
rect 674 -2243 675 -2237
rect 677 -2259 678 -2242
rect 681 -2243 682 -2237
rect 684 -2243 685 -2237
rect 688 -2312 689 -2242
rect 765 -2243 766 -2237
rect 800 -2312 801 -2242
rect 926 -2243 927 -2237
rect 957 -2243 958 -2237
rect 975 -2243 976 -2237
rect 44 -2312 45 -2244
rect 65 -2245 66 -2237
rect 128 -2312 129 -2244
rect 135 -2312 136 -2244
rect 156 -2245 157 -2237
rect 177 -2245 178 -2237
rect 240 -2245 241 -2237
rect 261 -2245 262 -2237
rect 355 -2245 356 -2237
rect 429 -2312 430 -2244
rect 506 -2245 507 -2237
rect 527 -2312 528 -2244
rect 548 -2245 549 -2237
rect 583 -2245 584 -2237
rect 586 -2259 587 -2244
rect 632 -2312 633 -2244
rect 646 -2245 647 -2237
rect 674 -2312 675 -2244
rect 758 -2245 759 -2237
rect 765 -2312 766 -2244
rect 814 -2245 815 -2237
rect 870 -2312 871 -2244
rect 954 -2245 955 -2237
rect 51 -2312 52 -2246
rect 114 -2247 115 -2237
rect 138 -2312 139 -2246
rect 565 -2312 566 -2246
rect 583 -2312 584 -2246
rect 621 -2312 622 -2246
rect 646 -2312 647 -2246
rect 681 -2312 682 -2246
rect 716 -2247 717 -2237
rect 723 -2247 724 -2237
rect 758 -2312 759 -2246
rect 807 -2312 808 -2246
rect 842 -2247 843 -2237
rect 65 -2312 66 -2248
rect 100 -2249 101 -2237
rect 114 -2312 115 -2248
rect 142 -2249 143 -2237
rect 170 -2249 171 -2237
rect 177 -2312 178 -2248
rect 180 -2249 181 -2237
rect 240 -2312 241 -2248
rect 247 -2249 248 -2237
rect 261 -2312 262 -2248
rect 303 -2249 304 -2237
rect 352 -2249 353 -2237
rect 436 -2249 437 -2237
rect 453 -2249 454 -2237
rect 478 -2312 479 -2248
rect 572 -2312 573 -2248
rect 639 -2249 640 -2237
rect 660 -2312 661 -2248
rect 698 -2249 699 -2237
rect 912 -2249 913 -2237
rect 72 -2251 73 -2237
rect 530 -2251 531 -2237
rect 534 -2251 535 -2237
rect 548 -2312 549 -2250
rect 611 -2251 612 -2237
rect 639 -2312 640 -2250
rect 702 -2251 703 -2237
rect 716 -2312 717 -2250
rect 730 -2251 731 -2237
rect 744 -2251 745 -2237
rect 747 -2251 748 -2237
rect 884 -2251 885 -2237
rect 72 -2312 73 -2252
rect 163 -2253 164 -2237
rect 184 -2253 185 -2237
rect 394 -2253 395 -2237
rect 408 -2253 409 -2237
rect 436 -2312 437 -2252
rect 446 -2253 447 -2237
rect 457 -2253 458 -2237
rect 499 -2253 500 -2237
rect 506 -2312 507 -2252
rect 604 -2253 605 -2237
rect 611 -2312 612 -2252
rect 656 -2312 657 -2252
rect 884 -2312 885 -2252
rect 79 -2312 80 -2254
rect 212 -2255 213 -2237
rect 226 -2255 227 -2237
rect 653 -2255 654 -2237
rect 709 -2255 710 -2237
rect 723 -2312 724 -2254
rect 730 -2312 731 -2254
rect 772 -2255 773 -2237
rect 814 -2312 815 -2254
rect 863 -2255 864 -2237
rect 96 -2257 97 -2237
rect 226 -2312 227 -2256
rect 247 -2312 248 -2256
rect 387 -2257 388 -2237
rect 408 -2312 409 -2256
rect 541 -2257 542 -2237
rect 576 -2257 577 -2237
rect 604 -2312 605 -2256
rect 737 -2257 738 -2237
rect 751 -2312 752 -2256
rect 772 -2312 773 -2256
rect 779 -2257 780 -2237
rect 842 -2312 843 -2256
rect 891 -2257 892 -2237
rect 100 -2312 101 -2258
rect 289 -2259 290 -2237
rect 303 -2312 304 -2258
rect 376 -2312 377 -2258
rect 387 -2312 388 -2258
rect 537 -2312 538 -2258
rect 737 -2312 738 -2258
rect 786 -2259 787 -2237
rect 810 -2312 811 -2258
rect 891 -2312 892 -2258
rect 107 -2261 108 -2237
rect 142 -2312 143 -2260
rect 156 -2312 157 -2260
rect 446 -2312 447 -2260
rect 471 -2261 472 -2237
rect 499 -2312 500 -2260
rect 740 -2261 741 -2237
rect 856 -2261 857 -2237
rect 863 -2312 864 -2260
rect 947 -2261 948 -2237
rect 107 -2312 108 -2262
rect 191 -2263 192 -2237
rect 198 -2263 199 -2237
rect 292 -2312 293 -2262
rect 310 -2263 311 -2237
rect 352 -2312 353 -2262
rect 366 -2263 367 -2237
rect 394 -2312 395 -2262
rect 492 -2263 493 -2237
rect 541 -2312 542 -2262
rect 744 -2312 745 -2262
rect 793 -2263 794 -2237
rect 856 -2312 857 -2262
rect 919 -2263 920 -2237
rect 124 -2265 125 -2237
rect 170 -2312 171 -2264
rect 198 -2312 199 -2264
rect 268 -2265 269 -2237
rect 275 -2265 276 -2237
rect 453 -2312 454 -2264
rect 779 -2312 780 -2264
rect 821 -2265 822 -2237
rect 149 -2267 150 -2237
rect 191 -2312 192 -2266
rect 205 -2267 206 -2237
rect 205 -2312 206 -2266
rect 205 -2267 206 -2237
rect 205 -2312 206 -2266
rect 212 -2312 213 -2266
rect 233 -2267 234 -2237
rect 254 -2267 255 -2237
rect 534 -2312 535 -2266
rect 653 -2312 654 -2266
rect 821 -2312 822 -2266
rect 149 -2312 150 -2268
rect 187 -2312 188 -2268
rect 219 -2269 220 -2237
rect 576 -2312 577 -2268
rect 786 -2312 787 -2268
rect 828 -2269 829 -2237
rect 163 -2312 164 -2270
rect 397 -2271 398 -2237
rect 793 -2312 794 -2270
rect 905 -2271 906 -2237
rect 184 -2312 185 -2272
rect 254 -2312 255 -2272
rect 268 -2312 269 -2272
rect 485 -2273 486 -2237
rect 828 -2312 829 -2272
rect 849 -2273 850 -2237
rect 219 -2312 220 -2274
rect 373 -2312 374 -2274
rect 443 -2275 444 -2237
rect 485 -2312 486 -2274
rect 849 -2312 850 -2274
rect 898 -2275 899 -2237
rect 93 -2312 94 -2276
rect 443 -2312 444 -2276
rect 877 -2277 878 -2237
rect 898 -2312 899 -2276
rect 233 -2312 234 -2278
rect 296 -2279 297 -2237
rect 310 -2312 311 -2278
rect 380 -2279 381 -2237
rect 877 -2312 878 -2278
rect 933 -2279 934 -2237
rect 275 -2312 276 -2280
rect 282 -2281 283 -2237
rect 296 -2312 297 -2280
rect 492 -2312 493 -2280
rect 282 -2312 283 -2282
rect 317 -2283 318 -2237
rect 324 -2283 325 -2237
rect 380 -2312 381 -2282
rect 317 -2312 318 -2284
rect 579 -2312 580 -2284
rect 324 -2312 325 -2286
rect 401 -2287 402 -2237
rect 331 -2289 332 -2237
rect 331 -2312 332 -2288
rect 331 -2289 332 -2237
rect 331 -2312 332 -2288
rect 345 -2312 346 -2288
rect 457 -2312 458 -2288
rect 366 -2312 367 -2290
rect 415 -2291 416 -2237
rect 121 -2293 122 -2237
rect 415 -2312 416 -2292
rect 121 -2312 122 -2294
rect 513 -2295 514 -2237
rect 401 -2312 402 -2296
rect 555 -2297 556 -2237
rect 422 -2299 423 -2237
rect 513 -2312 514 -2298
rect 555 -2312 556 -2298
rect 569 -2299 570 -2237
rect 422 -2312 423 -2300
rect 625 -2301 626 -2237
rect 464 -2303 465 -2237
rect 569 -2312 570 -2302
rect 590 -2303 591 -2237
rect 625 -2312 626 -2302
rect 464 -2312 465 -2304
rect 670 -2305 671 -2237
rect 590 -2312 591 -2306
rect 618 -2307 619 -2237
rect 562 -2309 563 -2237
rect 618 -2312 619 -2308
rect 471 -2312 472 -2310
rect 562 -2312 563 -2310
rect 51 -2322 52 -2320
rect 184 -2322 185 -2320
rect 187 -2377 188 -2321
rect 376 -2322 377 -2320
rect 383 -2377 384 -2321
rect 471 -2322 472 -2320
rect 492 -2322 493 -2320
rect 793 -2322 794 -2320
rect 884 -2322 885 -2320
rect 940 -2377 941 -2321
rect 968 -2322 969 -2320
rect 978 -2377 979 -2321
rect 982 -2377 983 -2321
rect 989 -2322 990 -2320
rect 996 -2322 997 -2320
rect 1003 -2377 1004 -2321
rect 1038 -2322 1039 -2320
rect 1059 -2322 1060 -2320
rect 65 -2324 66 -2320
rect 86 -2324 87 -2320
rect 89 -2324 90 -2320
rect 751 -2324 752 -2320
rect 772 -2324 773 -2320
rect 800 -2377 801 -2323
rect 898 -2324 899 -2320
rect 905 -2377 906 -2323
rect 989 -2377 990 -2323
rect 1006 -2377 1007 -2323
rect 44 -2326 45 -2320
rect 86 -2377 87 -2325
rect 135 -2377 136 -2325
rect 282 -2326 283 -2320
rect 306 -2377 307 -2325
rect 471 -2377 472 -2325
rect 492 -2377 493 -2325
rect 621 -2326 622 -2320
rect 632 -2326 633 -2320
rect 656 -2326 657 -2320
rect 698 -2377 699 -2325
rect 870 -2326 871 -2320
rect 891 -2326 892 -2320
rect 898 -2377 899 -2325
rect 138 -2328 139 -2320
rect 296 -2328 297 -2320
rect 310 -2328 311 -2320
rect 450 -2328 451 -2320
rect 457 -2328 458 -2320
rect 803 -2328 804 -2320
rect 152 -2377 153 -2329
rect 261 -2330 262 -2320
rect 275 -2330 276 -2320
rect 495 -2330 496 -2320
rect 520 -2330 521 -2320
rect 520 -2377 521 -2329
rect 520 -2330 521 -2320
rect 520 -2377 521 -2329
rect 558 -2377 559 -2329
rect 828 -2330 829 -2320
rect 114 -2332 115 -2320
rect 261 -2377 262 -2331
rect 292 -2332 293 -2320
rect 296 -2377 297 -2331
rect 338 -2332 339 -2320
rect 348 -2332 349 -2320
rect 352 -2332 353 -2320
rect 443 -2332 444 -2320
rect 446 -2332 447 -2320
rect 709 -2332 710 -2320
rect 716 -2332 717 -2320
rect 719 -2332 720 -2320
rect 751 -2377 752 -2331
rect 835 -2332 836 -2320
rect 114 -2377 115 -2333
rect 184 -2377 185 -2333
rect 205 -2334 206 -2320
rect 275 -2377 276 -2333
rect 338 -2377 339 -2333
rect 366 -2334 367 -2320
rect 387 -2334 388 -2320
rect 530 -2377 531 -2333
rect 548 -2334 549 -2320
rect 709 -2377 710 -2333
rect 716 -2377 717 -2333
rect 814 -2334 815 -2320
rect 93 -2336 94 -2320
rect 205 -2377 206 -2335
rect 233 -2336 234 -2320
rect 282 -2377 283 -2335
rect 359 -2336 360 -2320
rect 373 -2336 374 -2320
rect 387 -2377 388 -2335
rect 422 -2336 423 -2320
rect 429 -2336 430 -2320
rect 534 -2336 535 -2320
rect 562 -2336 563 -2320
rect 702 -2336 703 -2320
rect 772 -2377 773 -2335
rect 863 -2336 864 -2320
rect 93 -2377 94 -2337
rect 149 -2338 150 -2320
rect 163 -2338 164 -2320
rect 352 -2377 353 -2337
rect 359 -2377 360 -2337
rect 485 -2338 486 -2320
rect 534 -2377 535 -2337
rect 625 -2338 626 -2320
rect 632 -2377 633 -2337
rect 667 -2338 668 -2320
rect 702 -2377 703 -2337
rect 821 -2338 822 -2320
rect 121 -2340 122 -2320
rect 366 -2377 367 -2339
rect 394 -2340 395 -2320
rect 394 -2377 395 -2339
rect 394 -2340 395 -2320
rect 394 -2377 395 -2339
rect 401 -2340 402 -2320
rect 443 -2377 444 -2339
rect 453 -2340 454 -2320
rect 548 -2377 549 -2339
rect 555 -2340 556 -2320
rect 562 -2377 563 -2339
rect 569 -2340 570 -2320
rect 590 -2340 591 -2320
rect 604 -2340 605 -2320
rect 607 -2352 608 -2339
rect 614 -2377 615 -2339
rect 758 -2340 759 -2320
rect 779 -2340 780 -2320
rect 814 -2377 815 -2339
rect 121 -2377 122 -2341
rect 212 -2342 213 -2320
rect 226 -2342 227 -2320
rect 401 -2377 402 -2341
rect 415 -2342 416 -2320
rect 565 -2342 566 -2320
rect 569 -2377 570 -2341
rect 611 -2342 612 -2320
rect 618 -2342 619 -2320
rect 877 -2342 878 -2320
rect 149 -2377 150 -2343
rect 310 -2377 311 -2343
rect 324 -2344 325 -2320
rect 422 -2377 423 -2343
rect 429 -2377 430 -2343
rect 464 -2344 465 -2320
rect 485 -2377 486 -2343
rect 513 -2344 514 -2320
rect 555 -2377 556 -2343
rect 618 -2377 619 -2343
rect 667 -2377 668 -2343
rect 849 -2344 850 -2320
rect 72 -2346 73 -2320
rect 513 -2377 514 -2345
rect 572 -2346 573 -2320
rect 695 -2346 696 -2320
rect 730 -2346 731 -2320
rect 779 -2377 780 -2345
rect 793 -2377 794 -2345
rect 856 -2346 857 -2320
rect 72 -2377 73 -2347
rect 317 -2348 318 -2320
rect 436 -2348 437 -2320
rect 436 -2377 437 -2347
rect 436 -2348 437 -2320
rect 436 -2377 437 -2347
rect 457 -2377 458 -2347
rect 506 -2348 507 -2320
rect 576 -2348 577 -2320
rect 660 -2348 661 -2320
rect 730 -2377 731 -2347
rect 737 -2348 738 -2320
rect 758 -2377 759 -2347
rect 765 -2348 766 -2320
rect 107 -2350 108 -2320
rect 324 -2377 325 -2349
rect 464 -2377 465 -2349
rect 527 -2350 528 -2320
rect 576 -2377 577 -2349
rect 583 -2350 584 -2320
rect 590 -2377 591 -2349
rect 597 -2350 598 -2320
rect 604 -2377 605 -2349
rect 660 -2377 661 -2349
rect 674 -2350 675 -2320
rect 765 -2377 766 -2349
rect 842 -2350 843 -2320
rect 107 -2377 108 -2351
rect 380 -2352 381 -2320
rect 478 -2352 479 -2320
rect 506 -2377 507 -2351
rect 583 -2377 584 -2351
rect 688 -2352 689 -2320
rect 719 -2377 720 -2351
rect 737 -2377 738 -2351
rect 156 -2354 157 -2320
rect 212 -2377 213 -2353
rect 226 -2377 227 -2353
rect 233 -2377 234 -2353
rect 236 -2377 237 -2353
rect 695 -2377 696 -2353
rect 128 -2356 129 -2320
rect 156 -2377 157 -2355
rect 240 -2356 241 -2320
rect 240 -2377 241 -2355
rect 240 -2356 241 -2320
rect 240 -2377 241 -2355
rect 247 -2356 248 -2320
rect 425 -2356 426 -2320
rect 478 -2377 479 -2355
rect 541 -2356 542 -2320
rect 597 -2377 598 -2355
rect 639 -2356 640 -2320
rect 674 -2377 675 -2355
rect 786 -2356 787 -2320
rect 128 -2377 129 -2357
rect 219 -2358 220 -2320
rect 254 -2358 255 -2320
rect 373 -2377 374 -2357
rect 499 -2358 500 -2320
rect 611 -2377 612 -2357
rect 639 -2377 640 -2357
rect 681 -2358 682 -2320
rect 191 -2360 192 -2320
rect 247 -2377 248 -2359
rect 254 -2377 255 -2359
rect 450 -2377 451 -2359
rect 527 -2377 528 -2359
rect 688 -2377 689 -2359
rect 170 -2362 171 -2320
rect 191 -2377 192 -2361
rect 219 -2377 220 -2361
rect 268 -2362 269 -2320
rect 271 -2377 272 -2361
rect 415 -2377 416 -2361
rect 681 -2377 682 -2361
rect 744 -2362 745 -2320
rect 142 -2364 143 -2320
rect 170 -2377 171 -2363
rect 289 -2364 290 -2320
rect 541 -2377 542 -2363
rect 723 -2364 724 -2320
rect 744 -2377 745 -2363
rect 100 -2366 101 -2320
rect 289 -2377 290 -2365
rect 303 -2366 304 -2320
rect 625 -2377 626 -2365
rect 79 -2368 80 -2320
rect 303 -2377 304 -2367
rect 317 -2377 318 -2367
rect 345 -2368 346 -2320
rect 408 -2368 409 -2320
rect 499 -2377 500 -2367
rect 58 -2370 59 -2320
rect 79 -2377 80 -2369
rect 100 -2377 101 -2369
rect 163 -2377 164 -2369
rect 331 -2370 332 -2320
rect 345 -2377 346 -2369
rect 408 -2377 409 -2369
rect 653 -2370 654 -2320
rect 142 -2377 143 -2371
rect 516 -2377 517 -2371
rect 653 -2377 654 -2371
rect 807 -2372 808 -2320
rect 198 -2374 199 -2320
rect 331 -2377 332 -2373
rect 177 -2376 178 -2320
rect 198 -2377 199 -2375
rect 72 -2387 73 -2385
rect 163 -2387 164 -2385
rect 166 -2387 167 -2385
rect 198 -2387 199 -2385
rect 240 -2387 241 -2385
rect 240 -2428 241 -2386
rect 240 -2387 241 -2385
rect 240 -2428 241 -2386
rect 303 -2387 304 -2385
rect 345 -2387 346 -2385
rect 355 -2428 356 -2386
rect 541 -2387 542 -2385
rect 646 -2387 647 -2385
rect 684 -2428 685 -2386
rect 723 -2428 724 -2386
rect 730 -2387 731 -2385
rect 800 -2387 801 -2385
rect 807 -2428 808 -2386
rect 814 -2387 815 -2385
rect 828 -2428 829 -2386
rect 891 -2428 892 -2386
rect 905 -2387 906 -2385
rect 940 -2387 941 -2385
rect 1006 -2387 1007 -2385
rect 79 -2389 80 -2385
rect 187 -2389 188 -2385
rect 191 -2389 192 -2385
rect 236 -2389 237 -2385
rect 303 -2428 304 -2388
rect 401 -2389 402 -2385
rect 418 -2428 419 -2388
rect 698 -2389 699 -2385
rect 730 -2428 731 -2388
rect 744 -2389 745 -2385
rect 779 -2389 780 -2385
rect 800 -2428 801 -2388
rect 898 -2389 899 -2385
rect 898 -2428 899 -2388
rect 898 -2389 899 -2385
rect 898 -2428 899 -2388
rect 975 -2389 976 -2385
rect 989 -2389 990 -2385
rect 86 -2391 87 -2385
rect 149 -2391 150 -2385
rect 156 -2391 157 -2385
rect 173 -2391 174 -2385
rect 177 -2391 178 -2385
rect 247 -2391 248 -2385
rect 282 -2391 283 -2385
rect 401 -2428 402 -2390
rect 422 -2391 423 -2385
rect 614 -2391 615 -2385
rect 688 -2391 689 -2385
rect 744 -2428 745 -2390
rect 978 -2391 979 -2385
rect 982 -2391 983 -2385
rect 93 -2393 94 -2385
rect 184 -2393 185 -2385
rect 219 -2393 220 -2385
rect 422 -2428 423 -2392
rect 429 -2393 430 -2385
rect 488 -2428 489 -2392
rect 499 -2393 500 -2385
rect 527 -2428 528 -2392
rect 530 -2393 531 -2385
rect 625 -2393 626 -2385
rect 691 -2428 692 -2392
rect 905 -2428 906 -2392
rect 121 -2395 122 -2385
rect 268 -2395 269 -2385
rect 310 -2395 311 -2385
rect 383 -2395 384 -2385
rect 394 -2395 395 -2385
rect 509 -2428 510 -2394
rect 516 -2395 517 -2385
rect 702 -2395 703 -2385
rect 135 -2397 136 -2385
rect 450 -2397 451 -2385
rect 453 -2397 454 -2385
rect 653 -2397 654 -2385
rect 142 -2399 143 -2385
rect 198 -2428 199 -2398
rect 205 -2399 206 -2385
rect 219 -2428 220 -2398
rect 247 -2428 248 -2398
rect 261 -2399 262 -2385
rect 268 -2428 269 -2398
rect 306 -2399 307 -2385
rect 310 -2428 311 -2398
rect 408 -2399 409 -2385
rect 443 -2399 444 -2385
rect 558 -2399 559 -2385
rect 576 -2399 577 -2385
rect 625 -2428 626 -2398
rect 653 -2428 654 -2398
rect 674 -2399 675 -2385
rect 261 -2428 262 -2400
rect 324 -2401 325 -2385
rect 345 -2428 346 -2400
rect 383 -2428 384 -2400
rect 436 -2401 437 -2385
rect 443 -2428 444 -2400
rect 450 -2428 451 -2400
rect 464 -2401 465 -2385
rect 499 -2428 500 -2400
rect 506 -2401 507 -2385
rect 516 -2428 517 -2400
rect 583 -2401 584 -2385
rect 674 -2428 675 -2400
rect 716 -2401 717 -2385
rect 254 -2403 255 -2385
rect 324 -2428 325 -2402
rect 352 -2403 353 -2385
rect 541 -2428 542 -2402
rect 548 -2403 549 -2385
rect 646 -2428 647 -2402
rect 716 -2428 717 -2402
rect 751 -2403 752 -2385
rect 128 -2405 129 -2385
rect 254 -2428 255 -2404
rect 296 -2405 297 -2385
rect 394 -2428 395 -2404
rect 415 -2405 416 -2385
rect 464 -2428 465 -2404
rect 492 -2405 493 -2385
rect 506 -2428 507 -2404
rect 513 -2405 514 -2385
rect 583 -2428 584 -2404
rect 709 -2405 710 -2385
rect 751 -2428 752 -2404
rect 212 -2407 213 -2385
rect 296 -2428 297 -2406
rect 359 -2407 360 -2385
rect 408 -2428 409 -2406
rect 436 -2428 437 -2406
rect 457 -2407 458 -2385
rect 460 -2428 461 -2406
rect 485 -2407 486 -2385
rect 492 -2428 493 -2406
rect 534 -2407 535 -2385
rect 548 -2428 549 -2406
rect 555 -2407 556 -2385
rect 576 -2428 577 -2406
rect 597 -2407 598 -2385
rect 289 -2409 290 -2385
rect 359 -2428 360 -2408
rect 366 -2409 367 -2385
rect 611 -2409 612 -2385
rect 100 -2411 101 -2385
rect 289 -2428 290 -2410
rect 369 -2428 370 -2410
rect 387 -2411 388 -2385
rect 478 -2411 479 -2385
rect 534 -2428 535 -2410
rect 555 -2428 556 -2410
rect 688 -2428 689 -2410
rect 114 -2413 115 -2385
rect 387 -2428 388 -2412
rect 523 -2428 524 -2412
rect 569 -2413 570 -2385
rect 597 -2428 598 -2412
rect 604 -2413 605 -2385
rect 611 -2428 612 -2412
rect 632 -2413 633 -2385
rect 331 -2415 332 -2385
rect 478 -2428 479 -2414
rect 604 -2428 605 -2414
rect 667 -2415 668 -2385
rect 233 -2417 234 -2385
rect 331 -2428 332 -2416
rect 373 -2417 374 -2385
rect 513 -2428 514 -2416
rect 632 -2428 633 -2416
rect 660 -2417 661 -2385
rect 667 -2428 668 -2416
rect 681 -2417 682 -2385
rect 226 -2419 227 -2385
rect 233 -2428 234 -2418
rect 338 -2419 339 -2385
rect 373 -2428 374 -2418
rect 471 -2419 472 -2385
rect 569 -2428 570 -2418
rect 618 -2419 619 -2385
rect 660 -2428 661 -2418
rect 681 -2428 682 -2418
rect 765 -2419 766 -2385
rect 107 -2421 108 -2385
rect 226 -2428 227 -2420
rect 317 -2421 318 -2385
rect 338 -2428 339 -2420
rect 471 -2428 472 -2420
rect 562 -2421 563 -2385
rect 618 -2428 619 -2420
rect 639 -2421 640 -2385
rect 758 -2421 759 -2385
rect 765 -2428 766 -2420
rect 275 -2423 276 -2385
rect 317 -2428 318 -2422
rect 562 -2428 563 -2422
rect 590 -2423 591 -2385
rect 737 -2423 738 -2385
rect 758 -2428 759 -2422
rect 275 -2428 276 -2424
rect 380 -2425 381 -2385
rect 520 -2425 521 -2385
rect 590 -2428 591 -2424
rect 737 -2428 738 -2424
rect 772 -2425 773 -2385
rect 282 -2428 283 -2426
rect 380 -2428 381 -2426
rect 429 -2428 430 -2426
rect 520 -2428 521 -2426
rect 772 -2428 773 -2426
rect 793 -2427 794 -2385
rect 226 -2438 227 -2436
rect 352 -2438 353 -2436
rect 380 -2438 381 -2436
rect 471 -2438 472 -2436
rect 509 -2438 510 -2436
rect 576 -2438 577 -2436
rect 607 -2469 608 -2437
rect 618 -2438 619 -2436
rect 639 -2469 640 -2437
rect 691 -2438 692 -2436
rect 702 -2469 703 -2437
rect 716 -2438 717 -2436
rect 723 -2438 724 -2436
rect 723 -2469 724 -2437
rect 723 -2438 724 -2436
rect 723 -2469 724 -2437
rect 744 -2438 745 -2436
rect 758 -2438 759 -2436
rect 807 -2438 808 -2436
rect 817 -2469 818 -2437
rect 828 -2438 829 -2436
rect 828 -2469 829 -2437
rect 828 -2438 829 -2436
rect 828 -2469 829 -2437
rect 898 -2438 899 -2436
rect 905 -2438 906 -2436
rect 219 -2440 220 -2436
rect 226 -2469 227 -2439
rect 233 -2440 234 -2436
rect 243 -2448 244 -2439
rect 261 -2440 262 -2436
rect 366 -2440 367 -2436
rect 387 -2440 388 -2436
rect 513 -2469 514 -2439
rect 569 -2440 570 -2436
rect 611 -2440 612 -2436
rect 614 -2469 615 -2439
rect 908 -2440 909 -2436
rect 233 -2469 234 -2441
rect 275 -2442 276 -2436
rect 369 -2442 370 -2436
rect 387 -2469 388 -2441
rect 429 -2442 430 -2436
rect 432 -2469 433 -2441
rect 562 -2442 563 -2436
rect 572 -2442 573 -2436
rect 597 -2442 598 -2436
rect 611 -2469 612 -2441
rect 653 -2442 654 -2436
rect 660 -2442 661 -2436
rect 663 -2442 664 -2436
rect 688 -2442 689 -2436
rect 737 -2442 738 -2436
rect 747 -2442 748 -2436
rect 765 -2442 766 -2436
rect 800 -2442 801 -2436
rect 807 -2469 808 -2441
rect 891 -2442 892 -2436
rect 898 -2469 899 -2441
rect 236 -2469 237 -2443
rect 327 -2444 328 -2436
rect 331 -2444 332 -2436
rect 457 -2444 458 -2436
rect 460 -2444 461 -2436
rect 838 -2469 839 -2443
rect 240 -2446 241 -2436
rect 240 -2469 241 -2445
rect 240 -2446 241 -2436
rect 240 -2469 241 -2445
rect 282 -2446 283 -2436
rect 418 -2446 419 -2436
rect 450 -2446 451 -2436
rect 506 -2446 507 -2436
rect 509 -2469 510 -2445
rect 583 -2446 584 -2436
rect 590 -2446 591 -2436
rect 618 -2469 619 -2445
rect 625 -2446 626 -2436
rect 653 -2469 654 -2445
rect 660 -2469 661 -2445
rect 674 -2446 675 -2436
rect 730 -2446 731 -2436
rect 744 -2469 745 -2445
rect 751 -2446 752 -2436
rect 754 -2469 755 -2445
rect 296 -2448 297 -2436
rect 331 -2469 332 -2447
rect 338 -2448 339 -2436
rect 366 -2469 367 -2447
rect 401 -2448 402 -2436
rect 453 -2448 454 -2436
rect 457 -2469 458 -2447
rect 523 -2448 524 -2436
rect 576 -2469 577 -2447
rect 604 -2448 605 -2436
rect 625 -2469 626 -2447
rect 649 -2469 650 -2447
rect 663 -2469 664 -2447
rect 674 -2469 675 -2447
rect 751 -2469 752 -2447
rect 772 -2448 773 -2436
rect 254 -2450 255 -2436
rect 296 -2469 297 -2449
rect 310 -2450 311 -2436
rect 352 -2469 353 -2449
rect 373 -2450 374 -2436
rect 401 -2469 402 -2449
rect 408 -2450 409 -2436
rect 408 -2469 409 -2449
rect 408 -2450 409 -2436
rect 408 -2469 409 -2449
rect 453 -2469 454 -2449
rect 499 -2450 500 -2436
rect 597 -2469 598 -2449
rect 632 -2450 633 -2436
rect 646 -2450 647 -2436
rect 688 -2469 689 -2449
rect 198 -2452 199 -2436
rect 254 -2469 255 -2451
rect 268 -2452 269 -2436
rect 310 -2469 311 -2451
rect 317 -2452 318 -2436
rect 450 -2469 451 -2451
rect 464 -2452 465 -2436
rect 471 -2469 472 -2451
rect 499 -2469 500 -2451
rect 534 -2452 535 -2436
rect 541 -2452 542 -2436
rect 632 -2469 633 -2451
rect 646 -2469 647 -2451
rect 667 -2452 668 -2436
rect 341 -2469 342 -2453
rect 548 -2454 549 -2436
rect 345 -2456 346 -2436
rect 373 -2469 374 -2455
rect 443 -2456 444 -2436
rect 464 -2469 465 -2455
rect 478 -2456 479 -2436
rect 548 -2469 549 -2455
rect 303 -2458 304 -2436
rect 345 -2469 346 -2457
rect 348 -2469 349 -2457
rect 555 -2458 556 -2436
rect 394 -2460 395 -2436
rect 443 -2469 444 -2459
rect 478 -2469 479 -2459
rect 485 -2460 486 -2436
rect 527 -2460 528 -2436
rect 541 -2469 542 -2459
rect 359 -2462 360 -2436
rect 394 -2469 395 -2461
rect 422 -2462 423 -2436
rect 485 -2469 486 -2461
rect 492 -2462 493 -2436
rect 527 -2469 528 -2461
rect 289 -2464 290 -2436
rect 359 -2469 360 -2463
rect 415 -2464 416 -2436
rect 492 -2469 493 -2463
rect 422 -2469 423 -2465
rect 436 -2466 437 -2436
rect 436 -2469 437 -2467
rect 516 -2468 517 -2436
rect 226 -2479 227 -2477
rect 226 -2490 227 -2478
rect 226 -2479 227 -2477
rect 226 -2490 227 -2478
rect 240 -2479 241 -2477
rect 240 -2490 241 -2478
rect 240 -2479 241 -2477
rect 240 -2490 241 -2478
rect 247 -2479 248 -2477
rect 254 -2479 255 -2477
rect 296 -2479 297 -2477
rect 341 -2479 342 -2477
rect 359 -2479 360 -2477
rect 380 -2490 381 -2478
rect 390 -2490 391 -2478
rect 457 -2479 458 -2477
rect 492 -2479 493 -2477
rect 509 -2479 510 -2477
rect 513 -2479 514 -2477
rect 611 -2490 612 -2478
rect 649 -2479 650 -2477
rect 653 -2479 654 -2477
rect 674 -2479 675 -2477
rect 691 -2490 692 -2478
rect 723 -2479 724 -2477
rect 723 -2490 724 -2478
rect 723 -2479 724 -2477
rect 723 -2490 724 -2478
rect 726 -2490 727 -2478
rect 901 -2490 902 -2478
rect 310 -2481 311 -2477
rect 348 -2481 349 -2477
rect 359 -2490 360 -2480
rect 387 -2481 388 -2477
rect 394 -2481 395 -2477
rect 429 -2481 430 -2477
rect 432 -2481 433 -2477
rect 499 -2481 500 -2477
rect 527 -2481 528 -2477
rect 534 -2490 535 -2480
rect 541 -2481 542 -2477
rect 555 -2490 556 -2480
rect 604 -2481 605 -2477
rect 639 -2481 640 -2477
rect 653 -2490 654 -2480
rect 660 -2481 661 -2477
rect 688 -2481 689 -2477
rect 695 -2485 696 -2480
rect 744 -2481 745 -2477
rect 751 -2481 752 -2477
rect 807 -2481 808 -2477
rect 817 -2481 818 -2477
rect 828 -2481 829 -2477
rect 835 -2481 836 -2477
rect 898 -2481 899 -2477
rect 905 -2490 906 -2480
rect 331 -2483 332 -2477
rect 369 -2490 370 -2482
rect 373 -2483 374 -2477
rect 394 -2490 395 -2482
rect 401 -2490 402 -2482
rect 408 -2483 409 -2477
rect 443 -2483 444 -2477
rect 471 -2483 472 -2477
rect 548 -2483 549 -2477
rect 614 -2483 615 -2477
rect 632 -2483 633 -2477
rect 660 -2490 661 -2482
rect 688 -2490 689 -2482
rect 702 -2483 703 -2477
rect 352 -2485 353 -2477
rect 373 -2490 374 -2484
rect 404 -2490 405 -2484
rect 422 -2485 423 -2477
rect 446 -2485 447 -2477
rect 464 -2485 465 -2477
rect 485 -2485 486 -2477
rect 548 -2490 549 -2484
rect 551 -2490 552 -2484
rect 576 -2485 577 -2477
rect 597 -2485 598 -2477
rect 604 -2490 605 -2484
rect 614 -2490 615 -2484
rect 625 -2485 626 -2477
rect 702 -2490 703 -2484
rect 366 -2487 367 -2477
rect 387 -2490 388 -2486
rect 453 -2487 454 -2477
rect 478 -2487 479 -2477
rect 618 -2487 619 -2477
rect 632 -2490 633 -2486
rect 366 -2490 367 -2488
rect 436 -2489 437 -2477
rect 226 -2500 227 -2498
rect 233 -2500 234 -2498
rect 236 -2500 237 -2498
rect 240 -2500 241 -2498
rect 359 -2500 360 -2498
rect 366 -2500 367 -2498
rect 373 -2500 374 -2498
rect 394 -2500 395 -2498
rect 397 -2500 398 -2498
rect 408 -2500 409 -2498
rect 534 -2500 535 -2498
rect 548 -2500 549 -2498
rect 558 -2500 559 -2498
rect 901 -2500 902 -2498
rect 380 -2502 381 -2498
rect 401 -2502 402 -2498
rect 604 -2502 605 -2498
rect 611 -2502 612 -2498
rect 632 -2502 633 -2498
rect 653 -2502 654 -2498
rect 660 -2502 661 -2498
rect 691 -2502 692 -2498
rect 702 -2502 703 -2498
rect 726 -2502 727 -2498
rect 898 -2502 899 -2498
rect 905 -2502 906 -2498
<< labels >>
rlabel pdiffusion 150 -10 150 -10 0 cellNo=295
rlabel pdiffusion 206 -10 206 -10 0 cellNo=151
rlabel pdiffusion 339 -10 339 -10 0 cellNo=65
rlabel pdiffusion 346 -10 346 -10 0 feedthrough
rlabel pdiffusion 353 -10 353 -10 0 feedthrough
rlabel pdiffusion 360 -10 360 -10 0 feedthrough
rlabel pdiffusion 367 -10 367 -10 0 feedthrough
rlabel pdiffusion 374 -10 374 -10 0 cellNo=500
rlabel pdiffusion 395 -10 395 -10 0 feedthrough
rlabel pdiffusion 402 -10 402 -10 0 cellNo=82
rlabel pdiffusion 409 -10 409 -10 0 cellNo=237
rlabel pdiffusion 430 -10 430 -10 0 cellNo=267
rlabel pdiffusion 437 -10 437 -10 0 cellNo=363
rlabel pdiffusion 451 -10 451 -10 0 feedthrough
rlabel pdiffusion 465 -10 465 -10 0 feedthrough
rlabel pdiffusion 472 -10 472 -10 0 cellNo=527
rlabel pdiffusion 479 -10 479 -10 0 cellNo=169
rlabel pdiffusion 493 -10 493 -10 0 cellNo=153
rlabel pdiffusion 514 -10 514 -10 0 feedthrough
rlabel pdiffusion 577 -10 577 -10 0 feedthrough
rlabel pdiffusion 129 -41 129 -41 0 feedthrough
rlabel pdiffusion 199 -41 199 -41 0 feedthrough
rlabel pdiffusion 220 -41 220 -41 0 feedthrough
rlabel pdiffusion 241 -41 241 -41 0 cellNo=468
rlabel pdiffusion 255 -41 255 -41 0 feedthrough
rlabel pdiffusion 283 -41 283 -41 0 feedthrough
rlabel pdiffusion 290 -41 290 -41 0 cellNo=271
rlabel pdiffusion 297 -41 297 -41 0 feedthrough
rlabel pdiffusion 304 -41 304 -41 0 feedthrough
rlabel pdiffusion 311 -41 311 -41 0 feedthrough
rlabel pdiffusion 318 -41 318 -41 0 cellNo=465
rlabel pdiffusion 325 -41 325 -41 0 cellNo=216
rlabel pdiffusion 332 -41 332 -41 0 feedthrough
rlabel pdiffusion 339 -41 339 -41 0 feedthrough
rlabel pdiffusion 346 -41 346 -41 0 feedthrough
rlabel pdiffusion 353 -41 353 -41 0 feedthrough
rlabel pdiffusion 360 -41 360 -41 0 feedthrough
rlabel pdiffusion 367 -41 367 -41 0 feedthrough
rlabel pdiffusion 374 -41 374 -41 0 cellNo=272
rlabel pdiffusion 381 -41 381 -41 0 feedthrough
rlabel pdiffusion 388 -41 388 -41 0 feedthrough
rlabel pdiffusion 395 -41 395 -41 0 cellNo=565
rlabel pdiffusion 402 -41 402 -41 0 feedthrough
rlabel pdiffusion 409 -41 409 -41 0 feedthrough
rlabel pdiffusion 416 -41 416 -41 0 feedthrough
rlabel pdiffusion 423 -41 423 -41 0 feedthrough
rlabel pdiffusion 430 -41 430 -41 0 cellNo=442
rlabel pdiffusion 437 -41 437 -41 0 feedthrough
rlabel pdiffusion 444 -41 444 -41 0 cellNo=457
rlabel pdiffusion 451 -41 451 -41 0 feedthrough
rlabel pdiffusion 458 -41 458 -41 0 feedthrough
rlabel pdiffusion 465 -41 465 -41 0 feedthrough
rlabel pdiffusion 472 -41 472 -41 0 feedthrough
rlabel pdiffusion 479 -41 479 -41 0 feedthrough
rlabel pdiffusion 486 -41 486 -41 0 feedthrough
rlabel pdiffusion 493 -41 493 -41 0 cellNo=262
rlabel pdiffusion 500 -41 500 -41 0 cellNo=492
rlabel pdiffusion 507 -41 507 -41 0 feedthrough
rlabel pdiffusion 514 -41 514 -41 0 feedthrough
rlabel pdiffusion 528 -41 528 -41 0 feedthrough
rlabel pdiffusion 535 -41 535 -41 0 cellNo=242
rlabel pdiffusion 542 -41 542 -41 0 feedthrough
rlabel pdiffusion 549 -41 549 -41 0 feedthrough
rlabel pdiffusion 591 -41 591 -41 0 cellNo=208
rlabel pdiffusion 619 -41 619 -41 0 feedthrough
rlabel pdiffusion 626 -41 626 -41 0 feedthrough
rlabel pdiffusion 115 -94 115 -94 0 cellNo=469
rlabel pdiffusion 143 -94 143 -94 0 feedthrough
rlabel pdiffusion 164 -94 164 -94 0 feedthrough
rlabel pdiffusion 171 -94 171 -94 0 feedthrough
rlabel pdiffusion 178 -94 178 -94 0 feedthrough
rlabel pdiffusion 185 -94 185 -94 0 feedthrough
rlabel pdiffusion 192 -94 192 -94 0 feedthrough
rlabel pdiffusion 199 -94 199 -94 0 feedthrough
rlabel pdiffusion 206 -94 206 -94 0 feedthrough
rlabel pdiffusion 213 -94 213 -94 0 feedthrough
rlabel pdiffusion 220 -94 220 -94 0 feedthrough
rlabel pdiffusion 227 -94 227 -94 0 feedthrough
rlabel pdiffusion 234 -94 234 -94 0 feedthrough
rlabel pdiffusion 241 -94 241 -94 0 feedthrough
rlabel pdiffusion 248 -94 248 -94 0 feedthrough
rlabel pdiffusion 255 -94 255 -94 0 feedthrough
rlabel pdiffusion 262 -94 262 -94 0 feedthrough
rlabel pdiffusion 269 -94 269 -94 0 feedthrough
rlabel pdiffusion 276 -94 276 -94 0 cellNo=510
rlabel pdiffusion 283 -94 283 -94 0 feedthrough
rlabel pdiffusion 290 -94 290 -94 0 feedthrough
rlabel pdiffusion 297 -94 297 -94 0 feedthrough
rlabel pdiffusion 304 -94 304 -94 0 feedthrough
rlabel pdiffusion 311 -94 311 -94 0 feedthrough
rlabel pdiffusion 318 -94 318 -94 0 feedthrough
rlabel pdiffusion 325 -94 325 -94 0 feedthrough
rlabel pdiffusion 332 -94 332 -94 0 cellNo=258
rlabel pdiffusion 339 -94 339 -94 0 feedthrough
rlabel pdiffusion 346 -94 346 -94 0 cellNo=241
rlabel pdiffusion 353 -94 353 -94 0 feedthrough
rlabel pdiffusion 360 -94 360 -94 0 feedthrough
rlabel pdiffusion 367 -94 367 -94 0 cellNo=319
rlabel pdiffusion 374 -94 374 -94 0 cellNo=357
rlabel pdiffusion 381 -94 381 -94 0 cellNo=563
rlabel pdiffusion 388 -94 388 -94 0 cellNo=270
rlabel pdiffusion 395 -94 395 -94 0 cellNo=335
rlabel pdiffusion 402 -94 402 -94 0 feedthrough
rlabel pdiffusion 409 -94 409 -94 0 feedthrough
rlabel pdiffusion 416 -94 416 -94 0 feedthrough
rlabel pdiffusion 423 -94 423 -94 0 feedthrough
rlabel pdiffusion 430 -94 430 -94 0 feedthrough
rlabel pdiffusion 437 -94 437 -94 0 feedthrough
rlabel pdiffusion 444 -94 444 -94 0 feedthrough
rlabel pdiffusion 451 -94 451 -94 0 cellNo=539
rlabel pdiffusion 458 -94 458 -94 0 feedthrough
rlabel pdiffusion 465 -94 465 -94 0 feedthrough
rlabel pdiffusion 472 -94 472 -94 0 cellNo=392
rlabel pdiffusion 479 -94 479 -94 0 cellNo=536
rlabel pdiffusion 486 -94 486 -94 0 feedthrough
rlabel pdiffusion 493 -94 493 -94 0 feedthrough
rlabel pdiffusion 500 -94 500 -94 0 feedthrough
rlabel pdiffusion 507 -94 507 -94 0 feedthrough
rlabel pdiffusion 514 -94 514 -94 0 feedthrough
rlabel pdiffusion 521 -94 521 -94 0 feedthrough
rlabel pdiffusion 528 -94 528 -94 0 feedthrough
rlabel pdiffusion 535 -94 535 -94 0 feedthrough
rlabel pdiffusion 542 -94 542 -94 0 feedthrough
rlabel pdiffusion 549 -94 549 -94 0 feedthrough
rlabel pdiffusion 556 -94 556 -94 0 feedthrough
rlabel pdiffusion 563 -94 563 -94 0 feedthrough
rlabel pdiffusion 570 -94 570 -94 0 feedthrough
rlabel pdiffusion 577 -94 577 -94 0 feedthrough
rlabel pdiffusion 584 -94 584 -94 0 feedthrough
rlabel pdiffusion 591 -94 591 -94 0 cellNo=545
rlabel pdiffusion 598 -94 598 -94 0 feedthrough
rlabel pdiffusion 605 -94 605 -94 0 feedthrough
rlabel pdiffusion 612 -94 612 -94 0 feedthrough
rlabel pdiffusion 619 -94 619 -94 0 feedthrough
rlabel pdiffusion 626 -94 626 -94 0 feedthrough
rlabel pdiffusion 633 -94 633 -94 0 feedthrough
rlabel pdiffusion 640 -94 640 -94 0 feedthrough
rlabel pdiffusion 647 -94 647 -94 0 feedthrough
rlabel pdiffusion 654 -94 654 -94 0 feedthrough
rlabel pdiffusion 661 -94 661 -94 0 feedthrough
rlabel pdiffusion 668 -94 668 -94 0 feedthrough
rlabel pdiffusion 675 -94 675 -94 0 feedthrough
rlabel pdiffusion 682 -94 682 -94 0 feedthrough
rlabel pdiffusion 689 -94 689 -94 0 cellNo=164
rlabel pdiffusion 52 -161 52 -161 0 feedthrough
rlabel pdiffusion 59 -161 59 -161 0 feedthrough
rlabel pdiffusion 66 -161 66 -161 0 feedthrough
rlabel pdiffusion 73 -161 73 -161 0 feedthrough
rlabel pdiffusion 80 -161 80 -161 0 cellNo=25
rlabel pdiffusion 87 -161 87 -161 0 feedthrough
rlabel pdiffusion 94 -161 94 -161 0 feedthrough
rlabel pdiffusion 101 -161 101 -161 0 cellNo=449
rlabel pdiffusion 108 -161 108 -161 0 feedthrough
rlabel pdiffusion 115 -161 115 -161 0 feedthrough
rlabel pdiffusion 122 -161 122 -161 0 feedthrough
rlabel pdiffusion 129 -161 129 -161 0 feedthrough
rlabel pdiffusion 136 -161 136 -161 0 feedthrough
rlabel pdiffusion 143 -161 143 -161 0 cellNo=578
rlabel pdiffusion 150 -161 150 -161 0 cellNo=291
rlabel pdiffusion 157 -161 157 -161 0 feedthrough
rlabel pdiffusion 164 -161 164 -161 0 feedthrough
rlabel pdiffusion 171 -161 171 -161 0 feedthrough
rlabel pdiffusion 178 -161 178 -161 0 feedthrough
rlabel pdiffusion 185 -161 185 -161 0 cellNo=353
rlabel pdiffusion 192 -161 192 -161 0 cellNo=87
rlabel pdiffusion 199 -161 199 -161 0 cellNo=192
rlabel pdiffusion 206 -161 206 -161 0 feedthrough
rlabel pdiffusion 213 -161 213 -161 0 feedthrough
rlabel pdiffusion 220 -161 220 -161 0 feedthrough
rlabel pdiffusion 227 -161 227 -161 0 feedthrough
rlabel pdiffusion 234 -161 234 -161 0 feedthrough
rlabel pdiffusion 241 -161 241 -161 0 feedthrough
rlabel pdiffusion 248 -161 248 -161 0 feedthrough
rlabel pdiffusion 255 -161 255 -161 0 feedthrough
rlabel pdiffusion 262 -161 262 -161 0 feedthrough
rlabel pdiffusion 269 -161 269 -161 0 feedthrough
rlabel pdiffusion 276 -161 276 -161 0 feedthrough
rlabel pdiffusion 283 -161 283 -161 0 feedthrough
rlabel pdiffusion 290 -161 290 -161 0 feedthrough
rlabel pdiffusion 297 -161 297 -161 0 feedthrough
rlabel pdiffusion 304 -161 304 -161 0 feedthrough
rlabel pdiffusion 311 -161 311 -161 0 feedthrough
rlabel pdiffusion 318 -161 318 -161 0 feedthrough
rlabel pdiffusion 325 -161 325 -161 0 feedthrough
rlabel pdiffusion 332 -161 332 -161 0 feedthrough
rlabel pdiffusion 339 -161 339 -161 0 feedthrough
rlabel pdiffusion 346 -161 346 -161 0 feedthrough
rlabel pdiffusion 353 -161 353 -161 0 cellNo=175
rlabel pdiffusion 360 -161 360 -161 0 feedthrough
rlabel pdiffusion 367 -161 367 -161 0 feedthrough
rlabel pdiffusion 374 -161 374 -161 0 feedthrough
rlabel pdiffusion 381 -161 381 -161 0 feedthrough
rlabel pdiffusion 388 -161 388 -161 0 feedthrough
rlabel pdiffusion 395 -161 395 -161 0 feedthrough
rlabel pdiffusion 402 -161 402 -161 0 feedthrough
rlabel pdiffusion 409 -161 409 -161 0 cellNo=276
rlabel pdiffusion 416 -161 416 -161 0 cellNo=478
rlabel pdiffusion 423 -161 423 -161 0 feedthrough
rlabel pdiffusion 430 -161 430 -161 0 feedthrough
rlabel pdiffusion 437 -161 437 -161 0 feedthrough
rlabel pdiffusion 444 -161 444 -161 0 feedthrough
rlabel pdiffusion 451 -161 451 -161 0 cellNo=215
rlabel pdiffusion 458 -161 458 -161 0 feedthrough
rlabel pdiffusion 465 -161 465 -161 0 cellNo=34
rlabel pdiffusion 472 -161 472 -161 0 cellNo=591
rlabel pdiffusion 479 -161 479 -161 0 cellNo=548
rlabel pdiffusion 486 -161 486 -161 0 feedthrough
rlabel pdiffusion 493 -161 493 -161 0 cellNo=141
rlabel pdiffusion 500 -161 500 -161 0 feedthrough
rlabel pdiffusion 507 -161 507 -161 0 feedthrough
rlabel pdiffusion 514 -161 514 -161 0 feedthrough
rlabel pdiffusion 521 -161 521 -161 0 feedthrough
rlabel pdiffusion 528 -161 528 -161 0 feedthrough
rlabel pdiffusion 535 -161 535 -161 0 feedthrough
rlabel pdiffusion 542 -161 542 -161 0 feedthrough
rlabel pdiffusion 549 -161 549 -161 0 feedthrough
rlabel pdiffusion 556 -161 556 -161 0 feedthrough
rlabel pdiffusion 563 -161 563 -161 0 feedthrough
rlabel pdiffusion 570 -161 570 -161 0 feedthrough
rlabel pdiffusion 577 -161 577 -161 0 cellNo=185
rlabel pdiffusion 584 -161 584 -161 0 feedthrough
rlabel pdiffusion 591 -161 591 -161 0 feedthrough
rlabel pdiffusion 598 -161 598 -161 0 feedthrough
rlabel pdiffusion 605 -161 605 -161 0 feedthrough
rlabel pdiffusion 612 -161 612 -161 0 feedthrough
rlabel pdiffusion 619 -161 619 -161 0 feedthrough
rlabel pdiffusion 626 -161 626 -161 0 feedthrough
rlabel pdiffusion 633 -161 633 -161 0 feedthrough
rlabel pdiffusion 640 -161 640 -161 0 feedthrough
rlabel pdiffusion 647 -161 647 -161 0 feedthrough
rlabel pdiffusion 654 -161 654 -161 0 feedthrough
rlabel pdiffusion 661 -161 661 -161 0 feedthrough
rlabel pdiffusion 668 -161 668 -161 0 feedthrough
rlabel pdiffusion 675 -161 675 -161 0 feedthrough
rlabel pdiffusion 682 -161 682 -161 0 feedthrough
rlabel pdiffusion 689 -161 689 -161 0 feedthrough
rlabel pdiffusion 696 -161 696 -161 0 feedthrough
rlabel pdiffusion 703 -161 703 -161 0 feedthrough
rlabel pdiffusion 710 -161 710 -161 0 feedthrough
rlabel pdiffusion 717 -161 717 -161 0 feedthrough
rlabel pdiffusion 724 -161 724 -161 0 feedthrough
rlabel pdiffusion 731 -161 731 -161 0 feedthrough
rlabel pdiffusion 738 -161 738 -161 0 feedthrough
rlabel pdiffusion 745 -161 745 -161 0 feedthrough
rlabel pdiffusion 752 -161 752 -161 0 feedthrough
rlabel pdiffusion 759 -161 759 -161 0 feedthrough
rlabel pdiffusion 766 -161 766 -161 0 feedthrough
rlabel pdiffusion 773 -161 773 -161 0 feedthrough
rlabel pdiffusion 780 -161 780 -161 0 feedthrough
rlabel pdiffusion 787 -161 787 -161 0 feedthrough
rlabel pdiffusion 794 -161 794 -161 0 feedthrough
rlabel pdiffusion 801 -161 801 -161 0 feedthrough
rlabel pdiffusion 808 -161 808 -161 0 feedthrough
rlabel pdiffusion 815 -161 815 -161 0 feedthrough
rlabel pdiffusion 822 -161 822 -161 0 feedthrough
rlabel pdiffusion 45 -242 45 -242 0 feedthrough
rlabel pdiffusion 52 -242 52 -242 0 feedthrough
rlabel pdiffusion 59 -242 59 -242 0 feedthrough
rlabel pdiffusion 66 -242 66 -242 0 feedthrough
rlabel pdiffusion 73 -242 73 -242 0 feedthrough
rlabel pdiffusion 80 -242 80 -242 0 feedthrough
rlabel pdiffusion 87 -242 87 -242 0 feedthrough
rlabel pdiffusion 94 -242 94 -242 0 feedthrough
rlabel pdiffusion 101 -242 101 -242 0 cellNo=201
rlabel pdiffusion 108 -242 108 -242 0 feedthrough
rlabel pdiffusion 115 -242 115 -242 0 cellNo=54
rlabel pdiffusion 122 -242 122 -242 0 cellNo=26
rlabel pdiffusion 129 -242 129 -242 0 feedthrough
rlabel pdiffusion 136 -242 136 -242 0 cellNo=214
rlabel pdiffusion 143 -242 143 -242 0 feedthrough
rlabel pdiffusion 150 -242 150 -242 0 feedthrough
rlabel pdiffusion 157 -242 157 -242 0 feedthrough
rlabel pdiffusion 164 -242 164 -242 0 cellNo=179
rlabel pdiffusion 171 -242 171 -242 0 feedthrough
rlabel pdiffusion 178 -242 178 -242 0 feedthrough
rlabel pdiffusion 185 -242 185 -242 0 feedthrough
rlabel pdiffusion 192 -242 192 -242 0 feedthrough
rlabel pdiffusion 199 -242 199 -242 0 feedthrough
rlabel pdiffusion 206 -242 206 -242 0 feedthrough
rlabel pdiffusion 213 -242 213 -242 0 feedthrough
rlabel pdiffusion 220 -242 220 -242 0 feedthrough
rlabel pdiffusion 227 -242 227 -242 0 feedthrough
rlabel pdiffusion 234 -242 234 -242 0 feedthrough
rlabel pdiffusion 241 -242 241 -242 0 feedthrough
rlabel pdiffusion 248 -242 248 -242 0 feedthrough
rlabel pdiffusion 255 -242 255 -242 0 cellNo=401
rlabel pdiffusion 262 -242 262 -242 0 feedthrough
rlabel pdiffusion 269 -242 269 -242 0 feedthrough
rlabel pdiffusion 276 -242 276 -242 0 feedthrough
rlabel pdiffusion 283 -242 283 -242 0 cellNo=487
rlabel pdiffusion 290 -242 290 -242 0 cellNo=414
rlabel pdiffusion 297 -242 297 -242 0 feedthrough
rlabel pdiffusion 304 -242 304 -242 0 feedthrough
rlabel pdiffusion 311 -242 311 -242 0 feedthrough
rlabel pdiffusion 318 -242 318 -242 0 feedthrough
rlabel pdiffusion 325 -242 325 -242 0 feedthrough
rlabel pdiffusion 332 -242 332 -242 0 feedthrough
rlabel pdiffusion 339 -242 339 -242 0 feedthrough
rlabel pdiffusion 346 -242 346 -242 0 cellNo=315
rlabel pdiffusion 353 -242 353 -242 0 cellNo=191
rlabel pdiffusion 360 -242 360 -242 0 cellNo=119
rlabel pdiffusion 367 -242 367 -242 0 feedthrough
rlabel pdiffusion 374 -242 374 -242 0 cellNo=341
rlabel pdiffusion 381 -242 381 -242 0 feedthrough
rlabel pdiffusion 388 -242 388 -242 0 feedthrough
rlabel pdiffusion 395 -242 395 -242 0 feedthrough
rlabel pdiffusion 402 -242 402 -242 0 cellNo=394
rlabel pdiffusion 409 -242 409 -242 0 feedthrough
rlabel pdiffusion 416 -242 416 -242 0 feedthrough
rlabel pdiffusion 423 -242 423 -242 0 cellNo=395
rlabel pdiffusion 430 -242 430 -242 0 feedthrough
rlabel pdiffusion 437 -242 437 -242 0 cellNo=297
rlabel pdiffusion 444 -242 444 -242 0 feedthrough
rlabel pdiffusion 451 -242 451 -242 0 feedthrough
rlabel pdiffusion 458 -242 458 -242 0 cellNo=186
rlabel pdiffusion 465 -242 465 -242 0 feedthrough
rlabel pdiffusion 472 -242 472 -242 0 cellNo=110
rlabel pdiffusion 479 -242 479 -242 0 feedthrough
rlabel pdiffusion 486 -242 486 -242 0 feedthrough
rlabel pdiffusion 493 -242 493 -242 0 cellNo=562
rlabel pdiffusion 500 -242 500 -242 0 feedthrough
rlabel pdiffusion 507 -242 507 -242 0 feedthrough
rlabel pdiffusion 514 -242 514 -242 0 feedthrough
rlabel pdiffusion 521 -242 521 -242 0 feedthrough
rlabel pdiffusion 528 -242 528 -242 0 feedthrough
rlabel pdiffusion 535 -242 535 -242 0 feedthrough
rlabel pdiffusion 542 -242 542 -242 0 feedthrough
rlabel pdiffusion 549 -242 549 -242 0 feedthrough
rlabel pdiffusion 556 -242 556 -242 0 feedthrough
rlabel pdiffusion 563 -242 563 -242 0 feedthrough
rlabel pdiffusion 570 -242 570 -242 0 feedthrough
rlabel pdiffusion 577 -242 577 -242 0 feedthrough
rlabel pdiffusion 584 -242 584 -242 0 feedthrough
rlabel pdiffusion 591 -242 591 -242 0 feedthrough
rlabel pdiffusion 598 -242 598 -242 0 feedthrough
rlabel pdiffusion 605 -242 605 -242 0 feedthrough
rlabel pdiffusion 612 -242 612 -242 0 feedthrough
rlabel pdiffusion 619 -242 619 -242 0 feedthrough
rlabel pdiffusion 626 -242 626 -242 0 feedthrough
rlabel pdiffusion 633 -242 633 -242 0 feedthrough
rlabel pdiffusion 640 -242 640 -242 0 feedthrough
rlabel pdiffusion 647 -242 647 -242 0 feedthrough
rlabel pdiffusion 654 -242 654 -242 0 feedthrough
rlabel pdiffusion 661 -242 661 -242 0 feedthrough
rlabel pdiffusion 668 -242 668 -242 0 feedthrough
rlabel pdiffusion 675 -242 675 -242 0 feedthrough
rlabel pdiffusion 682 -242 682 -242 0 feedthrough
rlabel pdiffusion 689 -242 689 -242 0 feedthrough
rlabel pdiffusion 696 -242 696 -242 0 feedthrough
rlabel pdiffusion 703 -242 703 -242 0 feedthrough
rlabel pdiffusion 710 -242 710 -242 0 feedthrough
rlabel pdiffusion 717 -242 717 -242 0 feedthrough
rlabel pdiffusion 724 -242 724 -242 0 feedthrough
rlabel pdiffusion 731 -242 731 -242 0 feedthrough
rlabel pdiffusion 738 -242 738 -242 0 feedthrough
rlabel pdiffusion 745 -242 745 -242 0 feedthrough
rlabel pdiffusion 752 -242 752 -242 0 feedthrough
rlabel pdiffusion 759 -242 759 -242 0 feedthrough
rlabel pdiffusion 766 -242 766 -242 0 feedthrough
rlabel pdiffusion 773 -242 773 -242 0 feedthrough
rlabel pdiffusion 780 -242 780 -242 0 feedthrough
rlabel pdiffusion 787 -242 787 -242 0 feedthrough
rlabel pdiffusion 794 -242 794 -242 0 feedthrough
rlabel pdiffusion 801 -242 801 -242 0 feedthrough
rlabel pdiffusion 808 -242 808 -242 0 feedthrough
rlabel pdiffusion 815 -242 815 -242 0 feedthrough
rlabel pdiffusion 822 -242 822 -242 0 feedthrough
rlabel pdiffusion 829 -242 829 -242 0 feedthrough
rlabel pdiffusion 836 -242 836 -242 0 feedthrough
rlabel pdiffusion 843 -242 843 -242 0 feedthrough
rlabel pdiffusion 850 -242 850 -242 0 feedthrough
rlabel pdiffusion 857 -242 857 -242 0 cellNo=447
rlabel pdiffusion 864 -242 864 -242 0 feedthrough
rlabel pdiffusion 3 -331 3 -331 0 feedthrough
rlabel pdiffusion 10 -331 10 -331 0 feedthrough
rlabel pdiffusion 17 -331 17 -331 0 feedthrough
rlabel pdiffusion 24 -331 24 -331 0 feedthrough
rlabel pdiffusion 31 -331 31 -331 0 feedthrough
rlabel pdiffusion 38 -331 38 -331 0 feedthrough
rlabel pdiffusion 45 -331 45 -331 0 feedthrough
rlabel pdiffusion 52 -331 52 -331 0 feedthrough
rlabel pdiffusion 59 -331 59 -331 0 feedthrough
rlabel pdiffusion 66 -331 66 -331 0 cellNo=421
rlabel pdiffusion 73 -331 73 -331 0 feedthrough
rlabel pdiffusion 80 -331 80 -331 0 feedthrough
rlabel pdiffusion 87 -331 87 -331 0 feedthrough
rlabel pdiffusion 94 -331 94 -331 0 feedthrough
rlabel pdiffusion 101 -331 101 -331 0 feedthrough
rlabel pdiffusion 108 -331 108 -331 0 feedthrough
rlabel pdiffusion 115 -331 115 -331 0 feedthrough
rlabel pdiffusion 122 -331 122 -331 0 feedthrough
rlabel pdiffusion 129 -331 129 -331 0 cellNo=107
rlabel pdiffusion 136 -331 136 -331 0 feedthrough
rlabel pdiffusion 143 -331 143 -331 0 feedthrough
rlabel pdiffusion 150 -331 150 -331 0 feedthrough
rlabel pdiffusion 157 -331 157 -331 0 feedthrough
rlabel pdiffusion 164 -331 164 -331 0 feedthrough
rlabel pdiffusion 171 -331 171 -331 0 feedthrough
rlabel pdiffusion 178 -331 178 -331 0 feedthrough
rlabel pdiffusion 185 -331 185 -331 0 feedthrough
rlabel pdiffusion 192 -331 192 -331 0 cellNo=425
rlabel pdiffusion 199 -331 199 -331 0 feedthrough
rlabel pdiffusion 206 -331 206 -331 0 feedthrough
rlabel pdiffusion 213 -331 213 -331 0 feedthrough
rlabel pdiffusion 220 -331 220 -331 0 feedthrough
rlabel pdiffusion 227 -331 227 -331 0 feedthrough
rlabel pdiffusion 234 -331 234 -331 0 feedthrough
rlabel pdiffusion 241 -331 241 -331 0 feedthrough
rlabel pdiffusion 248 -331 248 -331 0 feedthrough
rlabel pdiffusion 255 -331 255 -331 0 feedthrough
rlabel pdiffusion 262 -331 262 -331 0 feedthrough
rlabel pdiffusion 269 -331 269 -331 0 feedthrough
rlabel pdiffusion 276 -331 276 -331 0 feedthrough
rlabel pdiffusion 283 -331 283 -331 0 feedthrough
rlabel pdiffusion 290 -331 290 -331 0 feedthrough
rlabel pdiffusion 297 -331 297 -331 0 feedthrough
rlabel pdiffusion 304 -331 304 -331 0 cellNo=182
rlabel pdiffusion 311 -331 311 -331 0 feedthrough
rlabel pdiffusion 318 -331 318 -331 0 feedthrough
rlabel pdiffusion 325 -331 325 -331 0 feedthrough
rlabel pdiffusion 332 -331 332 -331 0 feedthrough
rlabel pdiffusion 339 -331 339 -331 0 feedthrough
rlabel pdiffusion 346 -331 346 -331 0 feedthrough
rlabel pdiffusion 353 -331 353 -331 0 feedthrough
rlabel pdiffusion 360 -331 360 -331 0 feedthrough
rlabel pdiffusion 367 -331 367 -331 0 feedthrough
rlabel pdiffusion 374 -331 374 -331 0 cellNo=170
rlabel pdiffusion 381 -331 381 -331 0 cellNo=306
rlabel pdiffusion 388 -331 388 -331 0 feedthrough
rlabel pdiffusion 395 -331 395 -331 0 cellNo=423
rlabel pdiffusion 402 -331 402 -331 0 cellNo=249
rlabel pdiffusion 409 -331 409 -331 0 feedthrough
rlabel pdiffusion 416 -331 416 -331 0 cellNo=320
rlabel pdiffusion 423 -331 423 -331 0 cellNo=504
rlabel pdiffusion 430 -331 430 -331 0 feedthrough
rlabel pdiffusion 437 -331 437 -331 0 cellNo=313
rlabel pdiffusion 444 -331 444 -331 0 cellNo=260
rlabel pdiffusion 451 -331 451 -331 0 cellNo=156
rlabel pdiffusion 458 -331 458 -331 0 cellNo=8
rlabel pdiffusion 465 -331 465 -331 0 cellNo=489
rlabel pdiffusion 472 -331 472 -331 0 cellNo=168
rlabel pdiffusion 479 -331 479 -331 0 feedthrough
rlabel pdiffusion 486 -331 486 -331 0 cellNo=358
rlabel pdiffusion 493 -331 493 -331 0 feedthrough
rlabel pdiffusion 500 -331 500 -331 0 feedthrough
rlabel pdiffusion 507 -331 507 -331 0 feedthrough
rlabel pdiffusion 514 -331 514 -331 0 feedthrough
rlabel pdiffusion 521 -331 521 -331 0 feedthrough
rlabel pdiffusion 528 -331 528 -331 0 feedthrough
rlabel pdiffusion 535 -331 535 -331 0 feedthrough
rlabel pdiffusion 542 -331 542 -331 0 feedthrough
rlabel pdiffusion 549 -331 549 -331 0 cellNo=480
rlabel pdiffusion 556 -331 556 -331 0 feedthrough
rlabel pdiffusion 563 -331 563 -331 0 feedthrough
rlabel pdiffusion 570 -331 570 -331 0 cellNo=45
rlabel pdiffusion 577 -331 577 -331 0 feedthrough
rlabel pdiffusion 584 -331 584 -331 0 feedthrough
rlabel pdiffusion 591 -331 591 -331 0 feedthrough
rlabel pdiffusion 598 -331 598 -331 0 feedthrough
rlabel pdiffusion 605 -331 605 -331 0 feedthrough
rlabel pdiffusion 612 -331 612 -331 0 feedthrough
rlabel pdiffusion 619 -331 619 -331 0 feedthrough
rlabel pdiffusion 626 -331 626 -331 0 feedthrough
rlabel pdiffusion 633 -331 633 -331 0 feedthrough
rlabel pdiffusion 640 -331 640 -331 0 feedthrough
rlabel pdiffusion 647 -331 647 -331 0 feedthrough
rlabel pdiffusion 654 -331 654 -331 0 feedthrough
rlabel pdiffusion 661 -331 661 -331 0 feedthrough
rlabel pdiffusion 668 -331 668 -331 0 feedthrough
rlabel pdiffusion 675 -331 675 -331 0 feedthrough
rlabel pdiffusion 682 -331 682 -331 0 feedthrough
rlabel pdiffusion 689 -331 689 -331 0 cellNo=109
rlabel pdiffusion 696 -331 696 -331 0 feedthrough
rlabel pdiffusion 703 -331 703 -331 0 feedthrough
rlabel pdiffusion 710 -331 710 -331 0 feedthrough
rlabel pdiffusion 717 -331 717 -331 0 feedthrough
rlabel pdiffusion 724 -331 724 -331 0 feedthrough
rlabel pdiffusion 731 -331 731 -331 0 feedthrough
rlabel pdiffusion 738 -331 738 -331 0 feedthrough
rlabel pdiffusion 745 -331 745 -331 0 feedthrough
rlabel pdiffusion 752 -331 752 -331 0 feedthrough
rlabel pdiffusion 759 -331 759 -331 0 feedthrough
rlabel pdiffusion 766 -331 766 -331 0 feedthrough
rlabel pdiffusion 773 -331 773 -331 0 feedthrough
rlabel pdiffusion 780 -331 780 -331 0 feedthrough
rlabel pdiffusion 787 -331 787 -331 0 feedthrough
rlabel pdiffusion 794 -331 794 -331 0 feedthrough
rlabel pdiffusion 801 -331 801 -331 0 feedthrough
rlabel pdiffusion 808 -331 808 -331 0 feedthrough
rlabel pdiffusion 815 -331 815 -331 0 feedthrough
rlabel pdiffusion 822 -331 822 -331 0 feedthrough
rlabel pdiffusion 829 -331 829 -331 0 feedthrough
rlabel pdiffusion 836 -331 836 -331 0 feedthrough
rlabel pdiffusion 843 -331 843 -331 0 feedthrough
rlabel pdiffusion 850 -331 850 -331 0 feedthrough
rlabel pdiffusion 857 -331 857 -331 0 feedthrough
rlabel pdiffusion 864 -331 864 -331 0 feedthrough
rlabel pdiffusion 871 -331 871 -331 0 feedthrough
rlabel pdiffusion 878 -331 878 -331 0 feedthrough
rlabel pdiffusion 885 -331 885 -331 0 feedthrough
rlabel pdiffusion 892 -331 892 -331 0 feedthrough
rlabel pdiffusion 899 -331 899 -331 0 feedthrough
rlabel pdiffusion 906 -331 906 -331 0 feedthrough
rlabel pdiffusion 913 -331 913 -331 0 feedthrough
rlabel pdiffusion 920 -331 920 -331 0 feedthrough
rlabel pdiffusion 927 -331 927 -331 0 feedthrough
rlabel pdiffusion 934 -331 934 -331 0 feedthrough
rlabel pdiffusion 941 -331 941 -331 0 feedthrough
rlabel pdiffusion 948 -331 948 -331 0 feedthrough
rlabel pdiffusion 955 -331 955 -331 0 feedthrough
rlabel pdiffusion 3 -418 3 -418 0 feedthrough
rlabel pdiffusion 10 -418 10 -418 0 feedthrough
rlabel pdiffusion 17 -418 17 -418 0 feedthrough
rlabel pdiffusion 24 -418 24 -418 0 feedthrough
rlabel pdiffusion 31 -418 31 -418 0 feedthrough
rlabel pdiffusion 38 -418 38 -418 0 feedthrough
rlabel pdiffusion 45 -418 45 -418 0 feedthrough
rlabel pdiffusion 52 -418 52 -418 0 feedthrough
rlabel pdiffusion 59 -418 59 -418 0 feedthrough
rlabel pdiffusion 66 -418 66 -418 0 cellNo=411
rlabel pdiffusion 73 -418 73 -418 0 cellNo=515
rlabel pdiffusion 80 -418 80 -418 0 cellNo=70
rlabel pdiffusion 87 -418 87 -418 0 cellNo=116
rlabel pdiffusion 94 -418 94 -418 0 cellNo=446
rlabel pdiffusion 101 -418 101 -418 0 feedthrough
rlabel pdiffusion 108 -418 108 -418 0 feedthrough
rlabel pdiffusion 115 -418 115 -418 0 feedthrough
rlabel pdiffusion 122 -418 122 -418 0 cellNo=393
rlabel pdiffusion 129 -418 129 -418 0 feedthrough
rlabel pdiffusion 136 -418 136 -418 0 feedthrough
rlabel pdiffusion 143 -418 143 -418 0 feedthrough
rlabel pdiffusion 150 -418 150 -418 0 feedthrough
rlabel pdiffusion 157 -418 157 -418 0 cellNo=596
rlabel pdiffusion 164 -418 164 -418 0 feedthrough
rlabel pdiffusion 171 -418 171 -418 0 feedthrough
rlabel pdiffusion 178 -418 178 -418 0 feedthrough
rlabel pdiffusion 185 -418 185 -418 0 cellNo=78
rlabel pdiffusion 192 -418 192 -418 0 cellNo=22
rlabel pdiffusion 199 -418 199 -418 0 feedthrough
rlabel pdiffusion 206 -418 206 -418 0 feedthrough
rlabel pdiffusion 213 -418 213 -418 0 feedthrough
rlabel pdiffusion 220 -418 220 -418 0 feedthrough
rlabel pdiffusion 227 -418 227 -418 0 feedthrough
rlabel pdiffusion 234 -418 234 -418 0 feedthrough
rlabel pdiffusion 241 -418 241 -418 0 cellNo=200
rlabel pdiffusion 248 -418 248 -418 0 feedthrough
rlabel pdiffusion 255 -418 255 -418 0 feedthrough
rlabel pdiffusion 262 -418 262 -418 0 feedthrough
rlabel pdiffusion 269 -418 269 -418 0 feedthrough
rlabel pdiffusion 276 -418 276 -418 0 feedthrough
rlabel pdiffusion 283 -418 283 -418 0 feedthrough
rlabel pdiffusion 290 -418 290 -418 0 feedthrough
rlabel pdiffusion 297 -418 297 -418 0 feedthrough
rlabel pdiffusion 304 -418 304 -418 0 feedthrough
rlabel pdiffusion 311 -418 311 -418 0 feedthrough
rlabel pdiffusion 318 -418 318 -418 0 feedthrough
rlabel pdiffusion 325 -418 325 -418 0 feedthrough
rlabel pdiffusion 332 -418 332 -418 0 feedthrough
rlabel pdiffusion 339 -418 339 -418 0 feedthrough
rlabel pdiffusion 346 -418 346 -418 0 feedthrough
rlabel pdiffusion 353 -418 353 -418 0 cellNo=516
rlabel pdiffusion 360 -418 360 -418 0 cellNo=224
rlabel pdiffusion 367 -418 367 -418 0 feedthrough
rlabel pdiffusion 374 -418 374 -418 0 feedthrough
rlabel pdiffusion 381 -418 381 -418 0 feedthrough
rlabel pdiffusion 388 -418 388 -418 0 feedthrough
rlabel pdiffusion 395 -418 395 -418 0 cellNo=448
rlabel pdiffusion 402 -418 402 -418 0 feedthrough
rlabel pdiffusion 409 -418 409 -418 0 cellNo=416
rlabel pdiffusion 416 -418 416 -418 0 feedthrough
rlabel pdiffusion 423 -418 423 -418 0 feedthrough
rlabel pdiffusion 430 -418 430 -418 0 cellNo=184
rlabel pdiffusion 437 -418 437 -418 0 feedthrough
rlabel pdiffusion 444 -418 444 -418 0 feedthrough
rlabel pdiffusion 451 -418 451 -418 0 feedthrough
rlabel pdiffusion 458 -418 458 -418 0 cellNo=415
rlabel pdiffusion 465 -418 465 -418 0 cellNo=354
rlabel pdiffusion 472 -418 472 -418 0 feedthrough
rlabel pdiffusion 479 -418 479 -418 0 feedthrough
rlabel pdiffusion 486 -418 486 -418 0 feedthrough
rlabel pdiffusion 493 -418 493 -418 0 feedthrough
rlabel pdiffusion 500 -418 500 -418 0 feedthrough
rlabel pdiffusion 507 -418 507 -418 0 feedthrough
rlabel pdiffusion 514 -418 514 -418 0 cellNo=4
rlabel pdiffusion 521 -418 521 -418 0 feedthrough
rlabel pdiffusion 528 -418 528 -418 0 cellNo=232
rlabel pdiffusion 535 -418 535 -418 0 feedthrough
rlabel pdiffusion 542 -418 542 -418 0 feedthrough
rlabel pdiffusion 549 -418 549 -418 0 cellNo=400
rlabel pdiffusion 556 -418 556 -418 0 feedthrough
rlabel pdiffusion 563 -418 563 -418 0 feedthrough
rlabel pdiffusion 570 -418 570 -418 0 feedthrough
rlabel pdiffusion 577 -418 577 -418 0 feedthrough
rlabel pdiffusion 584 -418 584 -418 0 feedthrough
rlabel pdiffusion 591 -418 591 -418 0 feedthrough
rlabel pdiffusion 598 -418 598 -418 0 feedthrough
rlabel pdiffusion 605 -418 605 -418 0 feedthrough
rlabel pdiffusion 612 -418 612 -418 0 feedthrough
rlabel pdiffusion 619 -418 619 -418 0 cellNo=138
rlabel pdiffusion 626 -418 626 -418 0 feedthrough
rlabel pdiffusion 633 -418 633 -418 0 feedthrough
rlabel pdiffusion 640 -418 640 -418 0 feedthrough
rlabel pdiffusion 647 -418 647 -418 0 feedthrough
rlabel pdiffusion 654 -418 654 -418 0 feedthrough
rlabel pdiffusion 661 -418 661 -418 0 feedthrough
rlabel pdiffusion 668 -418 668 -418 0 feedthrough
rlabel pdiffusion 675 -418 675 -418 0 feedthrough
rlabel pdiffusion 682 -418 682 -418 0 feedthrough
rlabel pdiffusion 689 -418 689 -418 0 feedthrough
rlabel pdiffusion 696 -418 696 -418 0 feedthrough
rlabel pdiffusion 703 -418 703 -418 0 feedthrough
rlabel pdiffusion 710 -418 710 -418 0 feedthrough
rlabel pdiffusion 717 -418 717 -418 0 feedthrough
rlabel pdiffusion 724 -418 724 -418 0 feedthrough
rlabel pdiffusion 731 -418 731 -418 0 feedthrough
rlabel pdiffusion 738 -418 738 -418 0 feedthrough
rlabel pdiffusion 745 -418 745 -418 0 feedthrough
rlabel pdiffusion 752 -418 752 -418 0 feedthrough
rlabel pdiffusion 759 -418 759 -418 0 feedthrough
rlabel pdiffusion 766 -418 766 -418 0 feedthrough
rlabel pdiffusion 773 -418 773 -418 0 feedthrough
rlabel pdiffusion 780 -418 780 -418 0 feedthrough
rlabel pdiffusion 787 -418 787 -418 0 feedthrough
rlabel pdiffusion 794 -418 794 -418 0 feedthrough
rlabel pdiffusion 801 -418 801 -418 0 feedthrough
rlabel pdiffusion 808 -418 808 -418 0 feedthrough
rlabel pdiffusion 815 -418 815 -418 0 feedthrough
rlabel pdiffusion 822 -418 822 -418 0 feedthrough
rlabel pdiffusion 829 -418 829 -418 0 feedthrough
rlabel pdiffusion 836 -418 836 -418 0 feedthrough
rlabel pdiffusion 843 -418 843 -418 0 feedthrough
rlabel pdiffusion 850 -418 850 -418 0 feedthrough
rlabel pdiffusion 857 -418 857 -418 0 feedthrough
rlabel pdiffusion 864 -418 864 -418 0 feedthrough
rlabel pdiffusion 871 -418 871 -418 0 feedthrough
rlabel pdiffusion 878 -418 878 -418 0 feedthrough
rlabel pdiffusion 885 -418 885 -418 0 feedthrough
rlabel pdiffusion 892 -418 892 -418 0 feedthrough
rlabel pdiffusion 899 -418 899 -418 0 feedthrough
rlabel pdiffusion 906 -418 906 -418 0 feedthrough
rlabel pdiffusion 913 -418 913 -418 0 feedthrough
rlabel pdiffusion 920 -418 920 -418 0 feedthrough
rlabel pdiffusion 927 -418 927 -418 0 feedthrough
rlabel pdiffusion 934 -418 934 -418 0 feedthrough
rlabel pdiffusion 941 -418 941 -418 0 feedthrough
rlabel pdiffusion 948 -418 948 -418 0 feedthrough
rlabel pdiffusion 955 -418 955 -418 0 feedthrough
rlabel pdiffusion 962 -418 962 -418 0 feedthrough
rlabel pdiffusion 969 -418 969 -418 0 feedthrough
rlabel pdiffusion 976 -418 976 -418 0 feedthrough
rlabel pdiffusion 983 -418 983 -418 0 feedthrough
rlabel pdiffusion 990 -418 990 -418 0 feedthrough
rlabel pdiffusion 997 -418 997 -418 0 feedthrough
rlabel pdiffusion 1004 -418 1004 -418 0 feedthrough
rlabel pdiffusion 1025 -418 1025 -418 0 feedthrough
rlabel pdiffusion 3 -513 3 -513 0 feedthrough
rlabel pdiffusion 10 -513 10 -513 0 feedthrough
rlabel pdiffusion 17 -513 17 -513 0 feedthrough
rlabel pdiffusion 24 -513 24 -513 0 feedthrough
rlabel pdiffusion 31 -513 31 -513 0 feedthrough
rlabel pdiffusion 38 -513 38 -513 0 feedthrough
rlabel pdiffusion 45 -513 45 -513 0 feedthrough
rlabel pdiffusion 52 -513 52 -513 0 feedthrough
rlabel pdiffusion 59 -513 59 -513 0 feedthrough
rlabel pdiffusion 66 -513 66 -513 0 feedthrough
rlabel pdiffusion 73 -513 73 -513 0 feedthrough
rlabel pdiffusion 80 -513 80 -513 0 feedthrough
rlabel pdiffusion 87 -513 87 -513 0 feedthrough
rlabel pdiffusion 94 -513 94 -513 0 cellNo=112
rlabel pdiffusion 101 -513 101 -513 0 feedthrough
rlabel pdiffusion 108 -513 108 -513 0 feedthrough
rlabel pdiffusion 115 -513 115 -513 0 feedthrough
rlabel pdiffusion 122 -513 122 -513 0 feedthrough
rlabel pdiffusion 129 -513 129 -513 0 cellNo=51
rlabel pdiffusion 136 -513 136 -513 0 cellNo=66
rlabel pdiffusion 143 -513 143 -513 0 cellNo=343
rlabel pdiffusion 150 -513 150 -513 0 cellNo=19
rlabel pdiffusion 157 -513 157 -513 0 cellNo=332
rlabel pdiffusion 164 -513 164 -513 0 feedthrough
rlabel pdiffusion 171 -513 171 -513 0 feedthrough
rlabel pdiffusion 178 -513 178 -513 0 feedthrough
rlabel pdiffusion 185 -513 185 -513 0 feedthrough
rlabel pdiffusion 192 -513 192 -513 0 feedthrough
rlabel pdiffusion 199 -513 199 -513 0 feedthrough
rlabel pdiffusion 206 -513 206 -513 0 feedthrough
rlabel pdiffusion 213 -513 213 -513 0 feedthrough
rlabel pdiffusion 220 -513 220 -513 0 feedthrough
rlabel pdiffusion 227 -513 227 -513 0 feedthrough
rlabel pdiffusion 234 -513 234 -513 0 feedthrough
rlabel pdiffusion 241 -513 241 -513 0 feedthrough
rlabel pdiffusion 248 -513 248 -513 0 cellNo=240
rlabel pdiffusion 255 -513 255 -513 0 feedthrough
rlabel pdiffusion 262 -513 262 -513 0 feedthrough
rlabel pdiffusion 269 -513 269 -513 0 feedthrough
rlabel pdiffusion 276 -513 276 -513 0 feedthrough
rlabel pdiffusion 283 -513 283 -513 0 feedthrough
rlabel pdiffusion 290 -513 290 -513 0 feedthrough
rlabel pdiffusion 297 -513 297 -513 0 feedthrough
rlabel pdiffusion 304 -513 304 -513 0 feedthrough
rlabel pdiffusion 311 -513 311 -513 0 feedthrough
rlabel pdiffusion 318 -513 318 -513 0 feedthrough
rlabel pdiffusion 325 -513 325 -513 0 cellNo=62
rlabel pdiffusion 332 -513 332 -513 0 feedthrough
rlabel pdiffusion 339 -513 339 -513 0 feedthrough
rlabel pdiffusion 346 -513 346 -513 0 feedthrough
rlabel pdiffusion 353 -513 353 -513 0 feedthrough
rlabel pdiffusion 360 -513 360 -513 0 feedthrough
rlabel pdiffusion 367 -513 367 -513 0 feedthrough
rlabel pdiffusion 374 -513 374 -513 0 feedthrough
rlabel pdiffusion 381 -513 381 -513 0 feedthrough
rlabel pdiffusion 388 -513 388 -513 0 cellNo=310
rlabel pdiffusion 395 -513 395 -513 0 cellNo=554
rlabel pdiffusion 402 -513 402 -513 0 feedthrough
rlabel pdiffusion 409 -513 409 -513 0 cellNo=29
rlabel pdiffusion 416 -513 416 -513 0 feedthrough
rlabel pdiffusion 423 -513 423 -513 0 feedthrough
rlabel pdiffusion 430 -513 430 -513 0 feedthrough
rlabel pdiffusion 437 -513 437 -513 0 feedthrough
rlabel pdiffusion 444 -513 444 -513 0 cellNo=69
rlabel pdiffusion 451 -513 451 -513 0 feedthrough
rlabel pdiffusion 458 -513 458 -513 0 feedthrough
rlabel pdiffusion 465 -513 465 -513 0 feedthrough
rlabel pdiffusion 472 -513 472 -513 0 feedthrough
rlabel pdiffusion 479 -513 479 -513 0 cellNo=413
rlabel pdiffusion 486 -513 486 -513 0 feedthrough
rlabel pdiffusion 493 -513 493 -513 0 feedthrough
rlabel pdiffusion 500 -513 500 -513 0 feedthrough
rlabel pdiffusion 507 -513 507 -513 0 cellNo=350
rlabel pdiffusion 514 -513 514 -513 0 feedthrough
rlabel pdiffusion 521 -513 521 -513 0 cellNo=252
rlabel pdiffusion 528 -513 528 -513 0 feedthrough
rlabel pdiffusion 535 -513 535 -513 0 feedthrough
rlabel pdiffusion 542 -513 542 -513 0 feedthrough
rlabel pdiffusion 549 -513 549 -513 0 feedthrough
rlabel pdiffusion 556 -513 556 -513 0 feedthrough
rlabel pdiffusion 563 -513 563 -513 0 cellNo=331
rlabel pdiffusion 570 -513 570 -513 0 cellNo=535
rlabel pdiffusion 577 -513 577 -513 0 cellNo=132
rlabel pdiffusion 584 -513 584 -513 0 feedthrough
rlabel pdiffusion 591 -513 591 -513 0 feedthrough
rlabel pdiffusion 598 -513 598 -513 0 feedthrough
rlabel pdiffusion 605 -513 605 -513 0 cellNo=369
rlabel pdiffusion 612 -513 612 -513 0 feedthrough
rlabel pdiffusion 619 -513 619 -513 0 feedthrough
rlabel pdiffusion 626 -513 626 -513 0 feedthrough
rlabel pdiffusion 633 -513 633 -513 0 feedthrough
rlabel pdiffusion 640 -513 640 -513 0 feedthrough
rlabel pdiffusion 647 -513 647 -513 0 cellNo=98
rlabel pdiffusion 654 -513 654 -513 0 feedthrough
rlabel pdiffusion 661 -513 661 -513 0 feedthrough
rlabel pdiffusion 668 -513 668 -513 0 cellNo=367
rlabel pdiffusion 675 -513 675 -513 0 feedthrough
rlabel pdiffusion 682 -513 682 -513 0 feedthrough
rlabel pdiffusion 689 -513 689 -513 0 feedthrough
rlabel pdiffusion 696 -513 696 -513 0 feedthrough
rlabel pdiffusion 703 -513 703 -513 0 feedthrough
rlabel pdiffusion 710 -513 710 -513 0 feedthrough
rlabel pdiffusion 717 -513 717 -513 0 feedthrough
rlabel pdiffusion 724 -513 724 -513 0 feedthrough
rlabel pdiffusion 731 -513 731 -513 0 feedthrough
rlabel pdiffusion 738 -513 738 -513 0 feedthrough
rlabel pdiffusion 745 -513 745 -513 0 feedthrough
rlabel pdiffusion 752 -513 752 -513 0 cellNo=235
rlabel pdiffusion 759 -513 759 -513 0 feedthrough
rlabel pdiffusion 766 -513 766 -513 0 feedthrough
rlabel pdiffusion 773 -513 773 -513 0 feedthrough
rlabel pdiffusion 780 -513 780 -513 0 feedthrough
rlabel pdiffusion 787 -513 787 -513 0 feedthrough
rlabel pdiffusion 794 -513 794 -513 0 feedthrough
rlabel pdiffusion 801 -513 801 -513 0 feedthrough
rlabel pdiffusion 808 -513 808 -513 0 feedthrough
rlabel pdiffusion 815 -513 815 -513 0 feedthrough
rlabel pdiffusion 822 -513 822 -513 0 feedthrough
rlabel pdiffusion 829 -513 829 -513 0 feedthrough
rlabel pdiffusion 836 -513 836 -513 0 feedthrough
rlabel pdiffusion 843 -513 843 -513 0 feedthrough
rlabel pdiffusion 850 -513 850 -513 0 feedthrough
rlabel pdiffusion 857 -513 857 -513 0 feedthrough
rlabel pdiffusion 864 -513 864 -513 0 feedthrough
rlabel pdiffusion 871 -513 871 -513 0 feedthrough
rlabel pdiffusion 878 -513 878 -513 0 feedthrough
rlabel pdiffusion 885 -513 885 -513 0 feedthrough
rlabel pdiffusion 892 -513 892 -513 0 feedthrough
rlabel pdiffusion 899 -513 899 -513 0 feedthrough
rlabel pdiffusion 906 -513 906 -513 0 feedthrough
rlabel pdiffusion 913 -513 913 -513 0 feedthrough
rlabel pdiffusion 920 -513 920 -513 0 feedthrough
rlabel pdiffusion 927 -513 927 -513 0 feedthrough
rlabel pdiffusion 934 -513 934 -513 0 feedthrough
rlabel pdiffusion 941 -513 941 -513 0 feedthrough
rlabel pdiffusion 948 -513 948 -513 0 feedthrough
rlabel pdiffusion 955 -513 955 -513 0 feedthrough
rlabel pdiffusion 962 -513 962 -513 0 feedthrough
rlabel pdiffusion 969 -513 969 -513 0 feedthrough
rlabel pdiffusion 976 -513 976 -513 0 feedthrough
rlabel pdiffusion 983 -513 983 -513 0 feedthrough
rlabel pdiffusion 990 -513 990 -513 0 feedthrough
rlabel pdiffusion 997 -513 997 -513 0 feedthrough
rlabel pdiffusion 1004 -513 1004 -513 0 feedthrough
rlabel pdiffusion 1011 -513 1011 -513 0 feedthrough
rlabel pdiffusion 1018 -513 1018 -513 0 feedthrough
rlabel pdiffusion 1025 -513 1025 -513 0 feedthrough
rlabel pdiffusion 1032 -513 1032 -513 0 feedthrough
rlabel pdiffusion 1039 -513 1039 -513 0 feedthrough
rlabel pdiffusion 1046 -513 1046 -513 0 feedthrough
rlabel pdiffusion 1053 -513 1053 -513 0 feedthrough
rlabel pdiffusion 1060 -513 1060 -513 0 feedthrough
rlabel pdiffusion 1067 -513 1067 -513 0 feedthrough
rlabel pdiffusion 1074 -513 1074 -513 0 feedthrough
rlabel pdiffusion 1081 -513 1081 -513 0 feedthrough
rlabel pdiffusion 1088 -513 1088 -513 0 feedthrough
rlabel pdiffusion 1095 -513 1095 -513 0 feedthrough
rlabel pdiffusion 1102 -513 1102 -513 0 feedthrough
rlabel pdiffusion 1109 -513 1109 -513 0 feedthrough
rlabel pdiffusion 1116 -513 1116 -513 0 feedthrough
rlabel pdiffusion 1123 -513 1123 -513 0 feedthrough
rlabel pdiffusion 3 -612 3 -612 0 feedthrough
rlabel pdiffusion 10 -612 10 -612 0 feedthrough
rlabel pdiffusion 17 -612 17 -612 0 feedthrough
rlabel pdiffusion 24 -612 24 -612 0 feedthrough
rlabel pdiffusion 31 -612 31 -612 0 feedthrough
rlabel pdiffusion 38 -612 38 -612 0 cellNo=52
rlabel pdiffusion 45 -612 45 -612 0 feedthrough
rlabel pdiffusion 52 -612 52 -612 0 feedthrough
rlabel pdiffusion 59 -612 59 -612 0 cellNo=32
rlabel pdiffusion 66 -612 66 -612 0 cellNo=344
rlabel pdiffusion 73 -612 73 -612 0 cellNo=177
rlabel pdiffusion 80 -612 80 -612 0 feedthrough
rlabel pdiffusion 87 -612 87 -612 0 feedthrough
rlabel pdiffusion 94 -612 94 -612 0 feedthrough
rlabel pdiffusion 101 -612 101 -612 0 feedthrough
rlabel pdiffusion 108 -612 108 -612 0 feedthrough
rlabel pdiffusion 115 -612 115 -612 0 feedthrough
rlabel pdiffusion 122 -612 122 -612 0 feedthrough
rlabel pdiffusion 129 -612 129 -612 0 feedthrough
rlabel pdiffusion 136 -612 136 -612 0 feedthrough
rlabel pdiffusion 143 -612 143 -612 0 cellNo=125
rlabel pdiffusion 150 -612 150 -612 0 feedthrough
rlabel pdiffusion 157 -612 157 -612 0 feedthrough
rlabel pdiffusion 164 -612 164 -612 0 feedthrough
rlabel pdiffusion 171 -612 171 -612 0 feedthrough
rlabel pdiffusion 178 -612 178 -612 0 feedthrough
rlabel pdiffusion 185 -612 185 -612 0 cellNo=304
rlabel pdiffusion 192 -612 192 -612 0 feedthrough
rlabel pdiffusion 199 -612 199 -612 0 feedthrough
rlabel pdiffusion 206 -612 206 -612 0 feedthrough
rlabel pdiffusion 213 -612 213 -612 0 feedthrough
rlabel pdiffusion 220 -612 220 -612 0 feedthrough
rlabel pdiffusion 227 -612 227 -612 0 feedthrough
rlabel pdiffusion 234 -612 234 -612 0 feedthrough
rlabel pdiffusion 241 -612 241 -612 0 feedthrough
rlabel pdiffusion 248 -612 248 -612 0 feedthrough
rlabel pdiffusion 255 -612 255 -612 0 feedthrough
rlabel pdiffusion 262 -612 262 -612 0 feedthrough
rlabel pdiffusion 269 -612 269 -612 0 feedthrough
rlabel pdiffusion 276 -612 276 -612 0 cellNo=314
rlabel pdiffusion 283 -612 283 -612 0 feedthrough
rlabel pdiffusion 290 -612 290 -612 0 feedthrough
rlabel pdiffusion 297 -612 297 -612 0 feedthrough
rlabel pdiffusion 304 -612 304 -612 0 feedthrough
rlabel pdiffusion 311 -612 311 -612 0 feedthrough
rlabel pdiffusion 318 -612 318 -612 0 feedthrough
rlabel pdiffusion 325 -612 325 -612 0 feedthrough
rlabel pdiffusion 332 -612 332 -612 0 cellNo=518
rlabel pdiffusion 339 -612 339 -612 0 feedthrough
rlabel pdiffusion 346 -612 346 -612 0 feedthrough
rlabel pdiffusion 353 -612 353 -612 0 feedthrough
rlabel pdiffusion 360 -612 360 -612 0 feedthrough
rlabel pdiffusion 367 -612 367 -612 0 feedthrough
rlabel pdiffusion 374 -612 374 -612 0 feedthrough
rlabel pdiffusion 381 -612 381 -612 0 cellNo=274
rlabel pdiffusion 388 -612 388 -612 0 cellNo=127
rlabel pdiffusion 395 -612 395 -612 0 feedthrough
rlabel pdiffusion 402 -612 402 -612 0 cellNo=418
rlabel pdiffusion 409 -612 409 -612 0 feedthrough
rlabel pdiffusion 416 -612 416 -612 0 cellNo=264
rlabel pdiffusion 423 -612 423 -612 0 cellNo=549
rlabel pdiffusion 430 -612 430 -612 0 feedthrough
rlabel pdiffusion 437 -612 437 -612 0 feedthrough
rlabel pdiffusion 444 -612 444 -612 0 feedthrough
rlabel pdiffusion 451 -612 451 -612 0 cellNo=88
rlabel pdiffusion 458 -612 458 -612 0 cellNo=325
rlabel pdiffusion 465 -612 465 -612 0 cellNo=154
rlabel pdiffusion 472 -612 472 -612 0 feedthrough
rlabel pdiffusion 479 -612 479 -612 0 feedthrough
rlabel pdiffusion 486 -612 486 -612 0 feedthrough
rlabel pdiffusion 493 -612 493 -612 0 feedthrough
rlabel pdiffusion 500 -612 500 -612 0 feedthrough
rlabel pdiffusion 507 -612 507 -612 0 feedthrough
rlabel pdiffusion 514 -612 514 -612 0 feedthrough
rlabel pdiffusion 521 -612 521 -612 0 cellNo=173
rlabel pdiffusion 528 -612 528 -612 0 feedthrough
rlabel pdiffusion 535 -612 535 -612 0 feedthrough
rlabel pdiffusion 542 -612 542 -612 0 cellNo=33
rlabel pdiffusion 549 -612 549 -612 0 cellNo=202
rlabel pdiffusion 556 -612 556 -612 0 feedthrough
rlabel pdiffusion 563 -612 563 -612 0 cellNo=595
rlabel pdiffusion 570 -612 570 -612 0 feedthrough
rlabel pdiffusion 577 -612 577 -612 0 feedthrough
rlabel pdiffusion 584 -612 584 -612 0 cellNo=346
rlabel pdiffusion 591 -612 591 -612 0 feedthrough
rlabel pdiffusion 598 -612 598 -612 0 feedthrough
rlabel pdiffusion 605 -612 605 -612 0 feedthrough
rlabel pdiffusion 612 -612 612 -612 0 feedthrough
rlabel pdiffusion 619 -612 619 -612 0 cellNo=540
rlabel pdiffusion 626 -612 626 -612 0 cellNo=178
rlabel pdiffusion 633 -612 633 -612 0 feedthrough
rlabel pdiffusion 640 -612 640 -612 0 feedthrough
rlabel pdiffusion 647 -612 647 -612 0 feedthrough
rlabel pdiffusion 654 -612 654 -612 0 feedthrough
rlabel pdiffusion 661 -612 661 -612 0 feedthrough
rlabel pdiffusion 668 -612 668 -612 0 feedthrough
rlabel pdiffusion 675 -612 675 -612 0 feedthrough
rlabel pdiffusion 682 -612 682 -612 0 feedthrough
rlabel pdiffusion 689 -612 689 -612 0 feedthrough
rlabel pdiffusion 696 -612 696 -612 0 feedthrough
rlabel pdiffusion 703 -612 703 -612 0 feedthrough
rlabel pdiffusion 710 -612 710 -612 0 feedthrough
rlabel pdiffusion 717 -612 717 -612 0 feedthrough
rlabel pdiffusion 724 -612 724 -612 0 feedthrough
rlabel pdiffusion 731 -612 731 -612 0 feedthrough
rlabel pdiffusion 738 -612 738 -612 0 feedthrough
rlabel pdiffusion 745 -612 745 -612 0 feedthrough
rlabel pdiffusion 752 -612 752 -612 0 feedthrough
rlabel pdiffusion 759 -612 759 -612 0 feedthrough
rlabel pdiffusion 766 -612 766 -612 0 feedthrough
rlabel pdiffusion 773 -612 773 -612 0 feedthrough
rlabel pdiffusion 780 -612 780 -612 0 feedthrough
rlabel pdiffusion 787 -612 787 -612 0 feedthrough
rlabel pdiffusion 794 -612 794 -612 0 feedthrough
rlabel pdiffusion 801 -612 801 -612 0 feedthrough
rlabel pdiffusion 808 -612 808 -612 0 feedthrough
rlabel pdiffusion 815 -612 815 -612 0 feedthrough
rlabel pdiffusion 822 -612 822 -612 0 feedthrough
rlabel pdiffusion 829 -612 829 -612 0 feedthrough
rlabel pdiffusion 836 -612 836 -612 0 feedthrough
rlabel pdiffusion 843 -612 843 -612 0 feedthrough
rlabel pdiffusion 850 -612 850 -612 0 feedthrough
rlabel pdiffusion 857 -612 857 -612 0 feedthrough
rlabel pdiffusion 864 -612 864 -612 0 feedthrough
rlabel pdiffusion 871 -612 871 -612 0 feedthrough
rlabel pdiffusion 878 -612 878 -612 0 feedthrough
rlabel pdiffusion 885 -612 885 -612 0 feedthrough
rlabel pdiffusion 892 -612 892 -612 0 feedthrough
rlabel pdiffusion 899 -612 899 -612 0 feedthrough
rlabel pdiffusion 906 -612 906 -612 0 feedthrough
rlabel pdiffusion 913 -612 913 -612 0 feedthrough
rlabel pdiffusion 920 -612 920 -612 0 feedthrough
rlabel pdiffusion 927 -612 927 -612 0 feedthrough
rlabel pdiffusion 934 -612 934 -612 0 feedthrough
rlabel pdiffusion 941 -612 941 -612 0 feedthrough
rlabel pdiffusion 948 -612 948 -612 0 feedthrough
rlabel pdiffusion 955 -612 955 -612 0 feedthrough
rlabel pdiffusion 962 -612 962 -612 0 feedthrough
rlabel pdiffusion 969 -612 969 -612 0 feedthrough
rlabel pdiffusion 976 -612 976 -612 0 feedthrough
rlabel pdiffusion 983 -612 983 -612 0 feedthrough
rlabel pdiffusion 990 -612 990 -612 0 feedthrough
rlabel pdiffusion 997 -612 997 -612 0 feedthrough
rlabel pdiffusion 1004 -612 1004 -612 0 feedthrough
rlabel pdiffusion 1011 -612 1011 -612 0 feedthrough
rlabel pdiffusion 1018 -612 1018 -612 0 feedthrough
rlabel pdiffusion 1025 -612 1025 -612 0 feedthrough
rlabel pdiffusion 1032 -612 1032 -612 0 feedthrough
rlabel pdiffusion 1039 -612 1039 -612 0 feedthrough
rlabel pdiffusion 1046 -612 1046 -612 0 feedthrough
rlabel pdiffusion 1053 -612 1053 -612 0 feedthrough
rlabel pdiffusion 1060 -612 1060 -612 0 feedthrough
rlabel pdiffusion 1067 -612 1067 -612 0 feedthrough
rlabel pdiffusion 1074 -612 1074 -612 0 feedthrough
rlabel pdiffusion 1081 -612 1081 -612 0 cellNo=144
rlabel pdiffusion 1088 -612 1088 -612 0 feedthrough
rlabel pdiffusion 3 -721 3 -721 0 feedthrough
rlabel pdiffusion 10 -721 10 -721 0 feedthrough
rlabel pdiffusion 17 -721 17 -721 0 feedthrough
rlabel pdiffusion 24 -721 24 -721 0 feedthrough
rlabel pdiffusion 31 -721 31 -721 0 feedthrough
rlabel pdiffusion 38 -721 38 -721 0 feedthrough
rlabel pdiffusion 45 -721 45 -721 0 cellNo=124
rlabel pdiffusion 52 -721 52 -721 0 feedthrough
rlabel pdiffusion 59 -721 59 -721 0 cellNo=39
rlabel pdiffusion 66 -721 66 -721 0 feedthrough
rlabel pdiffusion 73 -721 73 -721 0 feedthrough
rlabel pdiffusion 80 -721 80 -721 0 feedthrough
rlabel pdiffusion 87 -721 87 -721 0 cellNo=35
rlabel pdiffusion 94 -721 94 -721 0 feedthrough
rlabel pdiffusion 101 -721 101 -721 0 feedthrough
rlabel pdiffusion 108 -721 108 -721 0 cellNo=183
rlabel pdiffusion 115 -721 115 -721 0 feedthrough
rlabel pdiffusion 122 -721 122 -721 0 feedthrough
rlabel pdiffusion 129 -721 129 -721 0 feedthrough
rlabel pdiffusion 136 -721 136 -721 0 feedthrough
rlabel pdiffusion 143 -721 143 -721 0 feedthrough
rlabel pdiffusion 150 -721 150 -721 0 feedthrough
rlabel pdiffusion 157 -721 157 -721 0 feedthrough
rlabel pdiffusion 164 -721 164 -721 0 feedthrough
rlabel pdiffusion 171 -721 171 -721 0 feedthrough
rlabel pdiffusion 178 -721 178 -721 0 feedthrough
rlabel pdiffusion 185 -721 185 -721 0 feedthrough
rlabel pdiffusion 192 -721 192 -721 0 cellNo=126
rlabel pdiffusion 199 -721 199 -721 0 feedthrough
rlabel pdiffusion 206 -721 206 -721 0 feedthrough
rlabel pdiffusion 213 -721 213 -721 0 feedthrough
rlabel pdiffusion 220 -721 220 -721 0 feedthrough
rlabel pdiffusion 227 -721 227 -721 0 cellNo=505
rlabel pdiffusion 234 -721 234 -721 0 cellNo=137
rlabel pdiffusion 241 -721 241 -721 0 feedthrough
rlabel pdiffusion 248 -721 248 -721 0 feedthrough
rlabel pdiffusion 255 -721 255 -721 0 feedthrough
rlabel pdiffusion 262 -721 262 -721 0 feedthrough
rlabel pdiffusion 269 -721 269 -721 0 feedthrough
rlabel pdiffusion 276 -721 276 -721 0 feedthrough
rlabel pdiffusion 283 -721 283 -721 0 feedthrough
rlabel pdiffusion 290 -721 290 -721 0 feedthrough
rlabel pdiffusion 297 -721 297 -721 0 feedthrough
rlabel pdiffusion 304 -721 304 -721 0 feedthrough
rlabel pdiffusion 311 -721 311 -721 0 feedthrough
rlabel pdiffusion 318 -721 318 -721 0 feedthrough
rlabel pdiffusion 325 -721 325 -721 0 feedthrough
rlabel pdiffusion 332 -721 332 -721 0 feedthrough
rlabel pdiffusion 339 -721 339 -721 0 feedthrough
rlabel pdiffusion 346 -721 346 -721 0 feedthrough
rlabel pdiffusion 353 -721 353 -721 0 feedthrough
rlabel pdiffusion 360 -721 360 -721 0 feedthrough
rlabel pdiffusion 367 -721 367 -721 0 cellNo=94
rlabel pdiffusion 374 -721 374 -721 0 feedthrough
rlabel pdiffusion 381 -721 381 -721 0 cellNo=422
rlabel pdiffusion 388 -721 388 -721 0 cellNo=90
rlabel pdiffusion 395 -721 395 -721 0 feedthrough
rlabel pdiffusion 402 -721 402 -721 0 cellNo=338
rlabel pdiffusion 409 -721 409 -721 0 feedthrough
rlabel pdiffusion 416 -721 416 -721 0 cellNo=122
rlabel pdiffusion 423 -721 423 -721 0 feedthrough
rlabel pdiffusion 430 -721 430 -721 0 cellNo=23
rlabel pdiffusion 437 -721 437 -721 0 feedthrough
rlabel pdiffusion 444 -721 444 -721 0 cellNo=225
rlabel pdiffusion 451 -721 451 -721 0 feedthrough
rlabel pdiffusion 458 -721 458 -721 0 feedthrough
rlabel pdiffusion 465 -721 465 -721 0 feedthrough
rlabel pdiffusion 472 -721 472 -721 0 feedthrough
rlabel pdiffusion 479 -721 479 -721 0 feedthrough
rlabel pdiffusion 486 -721 486 -721 0 feedthrough
rlabel pdiffusion 493 -721 493 -721 0 feedthrough
rlabel pdiffusion 500 -721 500 -721 0 cellNo=426
rlabel pdiffusion 507 -721 507 -721 0 feedthrough
rlabel pdiffusion 514 -721 514 -721 0 feedthrough
rlabel pdiffusion 521 -721 521 -721 0 feedthrough
rlabel pdiffusion 528 -721 528 -721 0 feedthrough
rlabel pdiffusion 535 -721 535 -721 0 feedthrough
rlabel pdiffusion 542 -721 542 -721 0 feedthrough
rlabel pdiffusion 549 -721 549 -721 0 feedthrough
rlabel pdiffusion 556 -721 556 -721 0 cellNo=250
rlabel pdiffusion 563 -721 563 -721 0 cellNo=385
rlabel pdiffusion 570 -721 570 -721 0 feedthrough
rlabel pdiffusion 577 -721 577 -721 0 feedthrough
rlabel pdiffusion 584 -721 584 -721 0 cellNo=160
rlabel pdiffusion 591 -721 591 -721 0 feedthrough
rlabel pdiffusion 598 -721 598 -721 0 feedthrough
rlabel pdiffusion 605 -721 605 -721 0 feedthrough
rlabel pdiffusion 612 -721 612 -721 0 feedthrough
rlabel pdiffusion 619 -721 619 -721 0 feedthrough
rlabel pdiffusion 626 -721 626 -721 0 feedthrough
rlabel pdiffusion 633 -721 633 -721 0 cellNo=218
rlabel pdiffusion 640 -721 640 -721 0 feedthrough
rlabel pdiffusion 647 -721 647 -721 0 cellNo=73
rlabel pdiffusion 654 -721 654 -721 0 cellNo=476
rlabel pdiffusion 661 -721 661 -721 0 feedthrough
rlabel pdiffusion 668 -721 668 -721 0 feedthrough
rlabel pdiffusion 675 -721 675 -721 0 feedthrough
rlabel pdiffusion 682 -721 682 -721 0 feedthrough
rlabel pdiffusion 689 -721 689 -721 0 feedthrough
rlabel pdiffusion 696 -721 696 -721 0 feedthrough
rlabel pdiffusion 703 -721 703 -721 0 feedthrough
rlabel pdiffusion 710 -721 710 -721 0 feedthrough
rlabel pdiffusion 717 -721 717 -721 0 feedthrough
rlabel pdiffusion 724 -721 724 -721 0 cellNo=495
rlabel pdiffusion 731 -721 731 -721 0 cellNo=213
rlabel pdiffusion 738 -721 738 -721 0 feedthrough
rlabel pdiffusion 745 -721 745 -721 0 feedthrough
rlabel pdiffusion 752 -721 752 -721 0 feedthrough
rlabel pdiffusion 759 -721 759 -721 0 feedthrough
rlabel pdiffusion 766 -721 766 -721 0 feedthrough
rlabel pdiffusion 773 -721 773 -721 0 feedthrough
rlabel pdiffusion 780 -721 780 -721 0 feedthrough
rlabel pdiffusion 787 -721 787 -721 0 feedthrough
rlabel pdiffusion 794 -721 794 -721 0 feedthrough
rlabel pdiffusion 801 -721 801 -721 0 feedthrough
rlabel pdiffusion 808 -721 808 -721 0 cellNo=531
rlabel pdiffusion 815 -721 815 -721 0 feedthrough
rlabel pdiffusion 822 -721 822 -721 0 feedthrough
rlabel pdiffusion 829 -721 829 -721 0 feedthrough
rlabel pdiffusion 836 -721 836 -721 0 feedthrough
rlabel pdiffusion 843 -721 843 -721 0 feedthrough
rlabel pdiffusion 850 -721 850 -721 0 feedthrough
rlabel pdiffusion 857 -721 857 -721 0 feedthrough
rlabel pdiffusion 864 -721 864 -721 0 feedthrough
rlabel pdiffusion 871 -721 871 -721 0 feedthrough
rlabel pdiffusion 878 -721 878 -721 0 feedthrough
rlabel pdiffusion 885 -721 885 -721 0 feedthrough
rlabel pdiffusion 892 -721 892 -721 0 feedthrough
rlabel pdiffusion 899 -721 899 -721 0 feedthrough
rlabel pdiffusion 906 -721 906 -721 0 feedthrough
rlabel pdiffusion 913 -721 913 -721 0 feedthrough
rlabel pdiffusion 920 -721 920 -721 0 feedthrough
rlabel pdiffusion 927 -721 927 -721 0 feedthrough
rlabel pdiffusion 934 -721 934 -721 0 feedthrough
rlabel pdiffusion 941 -721 941 -721 0 feedthrough
rlabel pdiffusion 948 -721 948 -721 0 feedthrough
rlabel pdiffusion 955 -721 955 -721 0 feedthrough
rlabel pdiffusion 962 -721 962 -721 0 feedthrough
rlabel pdiffusion 969 -721 969 -721 0 feedthrough
rlabel pdiffusion 976 -721 976 -721 0 feedthrough
rlabel pdiffusion 983 -721 983 -721 0 feedthrough
rlabel pdiffusion 990 -721 990 -721 0 feedthrough
rlabel pdiffusion 997 -721 997 -721 0 feedthrough
rlabel pdiffusion 1004 -721 1004 -721 0 feedthrough
rlabel pdiffusion 1011 -721 1011 -721 0 feedthrough
rlabel pdiffusion 1018 -721 1018 -721 0 feedthrough
rlabel pdiffusion 1025 -721 1025 -721 0 feedthrough
rlabel pdiffusion 1032 -721 1032 -721 0 feedthrough
rlabel pdiffusion 1039 -721 1039 -721 0 feedthrough
rlabel pdiffusion 1046 -721 1046 -721 0 feedthrough
rlabel pdiffusion 1053 -721 1053 -721 0 feedthrough
rlabel pdiffusion 1060 -721 1060 -721 0 feedthrough
rlabel pdiffusion 1067 -721 1067 -721 0 feedthrough
rlabel pdiffusion 1074 -721 1074 -721 0 feedthrough
rlabel pdiffusion 1081 -721 1081 -721 0 feedthrough
rlabel pdiffusion 1088 -721 1088 -721 0 feedthrough
rlabel pdiffusion 1095 -721 1095 -721 0 feedthrough
rlabel pdiffusion 1102 -721 1102 -721 0 feedthrough
rlabel pdiffusion 1109 -721 1109 -721 0 feedthrough
rlabel pdiffusion 1116 -721 1116 -721 0 feedthrough
rlabel pdiffusion 1123 -721 1123 -721 0 feedthrough
rlabel pdiffusion 1130 -721 1130 -721 0 feedthrough
rlabel pdiffusion 1137 -721 1137 -721 0 feedthrough
rlabel pdiffusion 1144 -721 1144 -721 0 feedthrough
rlabel pdiffusion 1151 -721 1151 -721 0 feedthrough
rlabel pdiffusion 1158 -721 1158 -721 0 feedthrough
rlabel pdiffusion 1165 -721 1165 -721 0 feedthrough
rlabel pdiffusion 1172 -721 1172 -721 0 feedthrough
rlabel pdiffusion 1179 -721 1179 -721 0 feedthrough
rlabel pdiffusion 1186 -721 1186 -721 0 feedthrough
rlabel pdiffusion 1193 -721 1193 -721 0 feedthrough
rlabel pdiffusion 1200 -721 1200 -721 0 feedthrough
rlabel pdiffusion 1207 -721 1207 -721 0 feedthrough
rlabel pdiffusion 1214 -721 1214 -721 0 cellNo=63
rlabel pdiffusion 1361 -721 1361 -721 0 feedthrough
rlabel pdiffusion 3 -838 3 -838 0 feedthrough
rlabel pdiffusion 10 -838 10 -838 0 feedthrough
rlabel pdiffusion 17 -838 17 -838 0 feedthrough
rlabel pdiffusion 24 -838 24 -838 0 cellNo=233
rlabel pdiffusion 31 -838 31 -838 0 cellNo=166
rlabel pdiffusion 38 -838 38 -838 0 feedthrough
rlabel pdiffusion 45 -838 45 -838 0 feedthrough
rlabel pdiffusion 52 -838 52 -838 0 feedthrough
rlabel pdiffusion 59 -838 59 -838 0 feedthrough
rlabel pdiffusion 66 -838 66 -838 0 feedthrough
rlabel pdiffusion 73 -838 73 -838 0 cellNo=13
rlabel pdiffusion 80 -838 80 -838 0 feedthrough
rlabel pdiffusion 87 -838 87 -838 0 cellNo=128
rlabel pdiffusion 94 -838 94 -838 0 feedthrough
rlabel pdiffusion 101 -838 101 -838 0 feedthrough
rlabel pdiffusion 108 -838 108 -838 0 feedthrough
rlabel pdiffusion 115 -838 115 -838 0 feedthrough
rlabel pdiffusion 122 -838 122 -838 0 feedthrough
rlabel pdiffusion 129 -838 129 -838 0 cellNo=60
rlabel pdiffusion 136 -838 136 -838 0 feedthrough
rlabel pdiffusion 143 -838 143 -838 0 feedthrough
rlabel pdiffusion 150 -838 150 -838 0 feedthrough
rlabel pdiffusion 157 -838 157 -838 0 feedthrough
rlabel pdiffusion 164 -838 164 -838 0 feedthrough
rlabel pdiffusion 171 -838 171 -838 0 feedthrough
rlabel pdiffusion 178 -838 178 -838 0 cellNo=294
rlabel pdiffusion 185 -838 185 -838 0 feedthrough
rlabel pdiffusion 192 -838 192 -838 0 feedthrough
rlabel pdiffusion 199 -838 199 -838 0 feedthrough
rlabel pdiffusion 206 -838 206 -838 0 feedthrough
rlabel pdiffusion 213 -838 213 -838 0 feedthrough
rlabel pdiffusion 220 -838 220 -838 0 feedthrough
rlabel pdiffusion 227 -838 227 -838 0 feedthrough
rlabel pdiffusion 234 -838 234 -838 0 feedthrough
rlabel pdiffusion 241 -838 241 -838 0 feedthrough
rlabel pdiffusion 248 -838 248 -838 0 feedthrough
rlabel pdiffusion 255 -838 255 -838 0 feedthrough
rlabel pdiffusion 262 -838 262 -838 0 feedthrough
rlabel pdiffusion 269 -838 269 -838 0 feedthrough
rlabel pdiffusion 276 -838 276 -838 0 feedthrough
rlabel pdiffusion 283 -838 283 -838 0 feedthrough
rlabel pdiffusion 290 -838 290 -838 0 feedthrough
rlabel pdiffusion 297 -838 297 -838 0 cellNo=152
rlabel pdiffusion 304 -838 304 -838 0 feedthrough
rlabel pdiffusion 311 -838 311 -838 0 feedthrough
rlabel pdiffusion 318 -838 318 -838 0 feedthrough
rlabel pdiffusion 325 -838 325 -838 0 feedthrough
rlabel pdiffusion 332 -838 332 -838 0 feedthrough
rlabel pdiffusion 339 -838 339 -838 0 feedthrough
rlabel pdiffusion 346 -838 346 -838 0 feedthrough
rlabel pdiffusion 353 -838 353 -838 0 feedthrough
rlabel pdiffusion 360 -838 360 -838 0 feedthrough
rlabel pdiffusion 367 -838 367 -838 0 feedthrough
rlabel pdiffusion 374 -838 374 -838 0 feedthrough
rlabel pdiffusion 381 -838 381 -838 0 feedthrough
rlabel pdiffusion 388 -838 388 -838 0 cellNo=145
rlabel pdiffusion 395 -838 395 -838 0 cellNo=327
rlabel pdiffusion 402 -838 402 -838 0 cellNo=37
rlabel pdiffusion 409 -838 409 -838 0 feedthrough
rlabel pdiffusion 416 -838 416 -838 0 feedthrough
rlabel pdiffusion 423 -838 423 -838 0 feedthrough
rlabel pdiffusion 430 -838 430 -838 0 cellNo=104
rlabel pdiffusion 437 -838 437 -838 0 cellNo=103
rlabel pdiffusion 444 -838 444 -838 0 feedthrough
rlabel pdiffusion 451 -838 451 -838 0 feedthrough
rlabel pdiffusion 458 -838 458 -838 0 feedthrough
rlabel pdiffusion 465 -838 465 -838 0 feedthrough
rlabel pdiffusion 472 -838 472 -838 0 feedthrough
rlabel pdiffusion 479 -838 479 -838 0 feedthrough
rlabel pdiffusion 486 -838 486 -838 0 feedthrough
rlabel pdiffusion 493 -838 493 -838 0 cellNo=445
rlabel pdiffusion 500 -838 500 -838 0 feedthrough
rlabel pdiffusion 507 -838 507 -838 0 cellNo=10
rlabel pdiffusion 514 -838 514 -838 0 cellNo=30
rlabel pdiffusion 521 -838 521 -838 0 cellNo=172
rlabel pdiffusion 528 -838 528 -838 0 feedthrough
rlabel pdiffusion 535 -838 535 -838 0 feedthrough
rlabel pdiffusion 542 -838 542 -838 0 feedthrough
rlabel pdiffusion 549 -838 549 -838 0 feedthrough
rlabel pdiffusion 556 -838 556 -838 0 feedthrough
rlabel pdiffusion 563 -838 563 -838 0 cellNo=481
rlabel pdiffusion 570 -838 570 -838 0 cellNo=261
rlabel pdiffusion 577 -838 577 -838 0 feedthrough
rlabel pdiffusion 584 -838 584 -838 0 cellNo=420
rlabel pdiffusion 591 -838 591 -838 0 feedthrough
rlabel pdiffusion 598 -838 598 -838 0 feedthrough
rlabel pdiffusion 605 -838 605 -838 0 feedthrough
rlabel pdiffusion 612 -838 612 -838 0 feedthrough
rlabel pdiffusion 619 -838 619 -838 0 cellNo=322
rlabel pdiffusion 626 -838 626 -838 0 feedthrough
rlabel pdiffusion 633 -838 633 -838 0 feedthrough
rlabel pdiffusion 640 -838 640 -838 0 feedthrough
rlabel pdiffusion 647 -838 647 -838 0 cellNo=149
rlabel pdiffusion 654 -838 654 -838 0 cellNo=75
rlabel pdiffusion 661 -838 661 -838 0 feedthrough
rlabel pdiffusion 668 -838 668 -838 0 feedthrough
rlabel pdiffusion 675 -838 675 -838 0 feedthrough
rlabel pdiffusion 682 -838 682 -838 0 feedthrough
rlabel pdiffusion 689 -838 689 -838 0 feedthrough
rlabel pdiffusion 696 -838 696 -838 0 feedthrough
rlabel pdiffusion 703 -838 703 -838 0 cellNo=59
rlabel pdiffusion 710 -838 710 -838 0 feedthrough
rlabel pdiffusion 717 -838 717 -838 0 feedthrough
rlabel pdiffusion 724 -838 724 -838 0 feedthrough
rlabel pdiffusion 731 -838 731 -838 0 feedthrough
rlabel pdiffusion 738 -838 738 -838 0 feedthrough
rlabel pdiffusion 745 -838 745 -838 0 feedthrough
rlabel pdiffusion 752 -838 752 -838 0 feedthrough
rlabel pdiffusion 759 -838 759 -838 0 cellNo=77
rlabel pdiffusion 766 -838 766 -838 0 feedthrough
rlabel pdiffusion 773 -838 773 -838 0 cellNo=566
rlabel pdiffusion 780 -838 780 -838 0 feedthrough
rlabel pdiffusion 787 -838 787 -838 0 feedthrough
rlabel pdiffusion 794 -838 794 -838 0 feedthrough
rlabel pdiffusion 801 -838 801 -838 0 feedthrough
rlabel pdiffusion 808 -838 808 -838 0 feedthrough
rlabel pdiffusion 815 -838 815 -838 0 feedthrough
rlabel pdiffusion 822 -838 822 -838 0 feedthrough
rlabel pdiffusion 829 -838 829 -838 0 cellNo=342
rlabel pdiffusion 836 -838 836 -838 0 feedthrough
rlabel pdiffusion 843 -838 843 -838 0 feedthrough
rlabel pdiffusion 850 -838 850 -838 0 feedthrough
rlabel pdiffusion 857 -838 857 -838 0 feedthrough
rlabel pdiffusion 864 -838 864 -838 0 feedthrough
rlabel pdiffusion 871 -838 871 -838 0 feedthrough
rlabel pdiffusion 878 -838 878 -838 0 feedthrough
rlabel pdiffusion 885 -838 885 -838 0 feedthrough
rlabel pdiffusion 892 -838 892 -838 0 feedthrough
rlabel pdiffusion 899 -838 899 -838 0 feedthrough
rlabel pdiffusion 906 -838 906 -838 0 feedthrough
rlabel pdiffusion 913 -838 913 -838 0 feedthrough
rlabel pdiffusion 920 -838 920 -838 0 feedthrough
rlabel pdiffusion 927 -838 927 -838 0 feedthrough
rlabel pdiffusion 934 -838 934 -838 0 feedthrough
rlabel pdiffusion 941 -838 941 -838 0 feedthrough
rlabel pdiffusion 948 -838 948 -838 0 feedthrough
rlabel pdiffusion 955 -838 955 -838 0 feedthrough
rlabel pdiffusion 962 -838 962 -838 0 feedthrough
rlabel pdiffusion 969 -838 969 -838 0 feedthrough
rlabel pdiffusion 976 -838 976 -838 0 feedthrough
rlabel pdiffusion 983 -838 983 -838 0 feedthrough
rlabel pdiffusion 990 -838 990 -838 0 feedthrough
rlabel pdiffusion 997 -838 997 -838 0 feedthrough
rlabel pdiffusion 1004 -838 1004 -838 0 feedthrough
rlabel pdiffusion 1011 -838 1011 -838 0 feedthrough
rlabel pdiffusion 1018 -838 1018 -838 0 feedthrough
rlabel pdiffusion 1025 -838 1025 -838 0 feedthrough
rlabel pdiffusion 1032 -838 1032 -838 0 feedthrough
rlabel pdiffusion 1039 -838 1039 -838 0 feedthrough
rlabel pdiffusion 1046 -838 1046 -838 0 feedthrough
rlabel pdiffusion 1053 -838 1053 -838 0 feedthrough
rlabel pdiffusion 1060 -838 1060 -838 0 feedthrough
rlabel pdiffusion 1067 -838 1067 -838 0 feedthrough
rlabel pdiffusion 1074 -838 1074 -838 0 feedthrough
rlabel pdiffusion 1081 -838 1081 -838 0 feedthrough
rlabel pdiffusion 1088 -838 1088 -838 0 feedthrough
rlabel pdiffusion 1095 -838 1095 -838 0 feedthrough
rlabel pdiffusion 1102 -838 1102 -838 0 feedthrough
rlabel pdiffusion 1109 -838 1109 -838 0 feedthrough
rlabel pdiffusion 1116 -838 1116 -838 0 feedthrough
rlabel pdiffusion 1123 -838 1123 -838 0 feedthrough
rlabel pdiffusion 1130 -838 1130 -838 0 feedthrough
rlabel pdiffusion 1137 -838 1137 -838 0 feedthrough
rlabel pdiffusion 1144 -838 1144 -838 0 feedthrough
rlabel pdiffusion 1151 -838 1151 -838 0 feedthrough
rlabel pdiffusion 1158 -838 1158 -838 0 feedthrough
rlabel pdiffusion 1165 -838 1165 -838 0 feedthrough
rlabel pdiffusion 1172 -838 1172 -838 0 feedthrough
rlabel pdiffusion 1179 -838 1179 -838 0 feedthrough
rlabel pdiffusion 1186 -838 1186 -838 0 feedthrough
rlabel pdiffusion 1193 -838 1193 -838 0 feedthrough
rlabel pdiffusion 1200 -838 1200 -838 0 feedthrough
rlabel pdiffusion 1207 -838 1207 -838 0 feedthrough
rlabel pdiffusion 1214 -838 1214 -838 0 feedthrough
rlabel pdiffusion 1221 -838 1221 -838 0 feedthrough
rlabel pdiffusion 1228 -838 1228 -838 0 feedthrough
rlabel pdiffusion 1235 -838 1235 -838 0 feedthrough
rlabel pdiffusion 1242 -838 1242 -838 0 feedthrough
rlabel pdiffusion 1249 -838 1249 -838 0 feedthrough
rlabel pdiffusion 1256 -838 1256 -838 0 feedthrough
rlabel pdiffusion 1263 -838 1263 -838 0 feedthrough
rlabel pdiffusion 1417 -838 1417 -838 0 feedthrough
rlabel pdiffusion 3 -955 3 -955 0 feedthrough
rlabel pdiffusion 10 -955 10 -955 0 feedthrough
rlabel pdiffusion 17 -955 17 -955 0 feedthrough
rlabel pdiffusion 24 -955 24 -955 0 feedthrough
rlabel pdiffusion 31 -955 31 -955 0 feedthrough
rlabel pdiffusion 38 -955 38 -955 0 feedthrough
rlabel pdiffusion 45 -955 45 -955 0 feedthrough
rlabel pdiffusion 52 -955 52 -955 0 feedthrough
rlabel pdiffusion 59 -955 59 -955 0 feedthrough
rlabel pdiffusion 66 -955 66 -955 0 cellNo=299
rlabel pdiffusion 73 -955 73 -955 0 feedthrough
rlabel pdiffusion 80 -955 80 -955 0 feedthrough
rlabel pdiffusion 87 -955 87 -955 0 cellNo=380
rlabel pdiffusion 94 -955 94 -955 0 feedthrough
rlabel pdiffusion 101 -955 101 -955 0 feedthrough
rlabel pdiffusion 108 -955 108 -955 0 feedthrough
rlabel pdiffusion 115 -955 115 -955 0 feedthrough
rlabel pdiffusion 122 -955 122 -955 0 cellNo=194
rlabel pdiffusion 129 -955 129 -955 0 cellNo=458
rlabel pdiffusion 136 -955 136 -955 0 feedthrough
rlabel pdiffusion 143 -955 143 -955 0 feedthrough
rlabel pdiffusion 150 -955 150 -955 0 cellNo=176
rlabel pdiffusion 157 -955 157 -955 0 feedthrough
rlabel pdiffusion 164 -955 164 -955 0 feedthrough
rlabel pdiffusion 171 -955 171 -955 0 feedthrough
rlabel pdiffusion 178 -955 178 -955 0 feedthrough
rlabel pdiffusion 185 -955 185 -955 0 feedthrough
rlabel pdiffusion 192 -955 192 -955 0 feedthrough
rlabel pdiffusion 199 -955 199 -955 0 cellNo=284
rlabel pdiffusion 206 -955 206 -955 0 feedthrough
rlabel pdiffusion 213 -955 213 -955 0 cellNo=56
rlabel pdiffusion 220 -955 220 -955 0 feedthrough
rlabel pdiffusion 227 -955 227 -955 0 feedthrough
rlabel pdiffusion 234 -955 234 -955 0 feedthrough
rlabel pdiffusion 241 -955 241 -955 0 feedthrough
rlabel pdiffusion 248 -955 248 -955 0 feedthrough
rlabel pdiffusion 255 -955 255 -955 0 feedthrough
rlabel pdiffusion 262 -955 262 -955 0 feedthrough
rlabel pdiffusion 269 -955 269 -955 0 feedthrough
rlabel pdiffusion 276 -955 276 -955 0 feedthrough
rlabel pdiffusion 283 -955 283 -955 0 feedthrough
rlabel pdiffusion 290 -955 290 -955 0 feedthrough
rlabel pdiffusion 297 -955 297 -955 0 feedthrough
rlabel pdiffusion 304 -955 304 -955 0 feedthrough
rlabel pdiffusion 311 -955 311 -955 0 feedthrough
rlabel pdiffusion 318 -955 318 -955 0 cellNo=55
rlabel pdiffusion 325 -955 325 -955 0 feedthrough
rlabel pdiffusion 332 -955 332 -955 0 feedthrough
rlabel pdiffusion 339 -955 339 -955 0 feedthrough
rlabel pdiffusion 346 -955 346 -955 0 feedthrough
rlabel pdiffusion 353 -955 353 -955 0 feedthrough
rlabel pdiffusion 360 -955 360 -955 0 feedthrough
rlabel pdiffusion 367 -955 367 -955 0 cellNo=263
rlabel pdiffusion 374 -955 374 -955 0 feedthrough
rlabel pdiffusion 381 -955 381 -955 0 feedthrough
rlabel pdiffusion 388 -955 388 -955 0 feedthrough
rlabel pdiffusion 395 -955 395 -955 0 feedthrough
rlabel pdiffusion 402 -955 402 -955 0 feedthrough
rlabel pdiffusion 409 -955 409 -955 0 feedthrough
rlabel pdiffusion 416 -955 416 -955 0 feedthrough
rlabel pdiffusion 423 -955 423 -955 0 cellNo=383
rlabel pdiffusion 430 -955 430 -955 0 feedthrough
rlabel pdiffusion 437 -955 437 -955 0 feedthrough
rlabel pdiffusion 444 -955 444 -955 0 feedthrough
rlabel pdiffusion 451 -955 451 -955 0 cellNo=573
rlabel pdiffusion 458 -955 458 -955 0 feedthrough
rlabel pdiffusion 465 -955 465 -955 0 feedthrough
rlabel pdiffusion 472 -955 472 -955 0 feedthrough
rlabel pdiffusion 479 -955 479 -955 0 cellNo=537
rlabel pdiffusion 486 -955 486 -955 0 feedthrough
rlabel pdiffusion 493 -955 493 -955 0 feedthrough
rlabel pdiffusion 500 -955 500 -955 0 cellNo=316
rlabel pdiffusion 507 -955 507 -955 0 feedthrough
rlabel pdiffusion 514 -955 514 -955 0 feedthrough
rlabel pdiffusion 521 -955 521 -955 0 feedthrough
rlabel pdiffusion 528 -955 528 -955 0 cellNo=99
rlabel pdiffusion 535 -955 535 -955 0 cellNo=419
rlabel pdiffusion 542 -955 542 -955 0 cellNo=57
rlabel pdiffusion 549 -955 549 -955 0 feedthrough
rlabel pdiffusion 556 -955 556 -955 0 feedthrough
rlabel pdiffusion 563 -955 563 -955 0 feedthrough
rlabel pdiffusion 570 -955 570 -955 0 feedthrough
rlabel pdiffusion 577 -955 577 -955 0 feedthrough
rlabel pdiffusion 584 -955 584 -955 0 feedthrough
rlabel pdiffusion 591 -955 591 -955 0 feedthrough
rlabel pdiffusion 598 -955 598 -955 0 feedthrough
rlabel pdiffusion 605 -955 605 -955 0 feedthrough
rlabel pdiffusion 612 -955 612 -955 0 cellNo=300
rlabel pdiffusion 619 -955 619 -955 0 feedthrough
rlabel pdiffusion 626 -955 626 -955 0 cellNo=528
rlabel pdiffusion 633 -955 633 -955 0 cellNo=301
rlabel pdiffusion 640 -955 640 -955 0 feedthrough
rlabel pdiffusion 647 -955 647 -955 0 feedthrough
rlabel pdiffusion 654 -955 654 -955 0 cellNo=41
rlabel pdiffusion 661 -955 661 -955 0 feedthrough
rlabel pdiffusion 668 -955 668 -955 0 feedthrough
rlabel pdiffusion 675 -955 675 -955 0 feedthrough
rlabel pdiffusion 682 -955 682 -955 0 feedthrough
rlabel pdiffusion 689 -955 689 -955 0 cellNo=485
rlabel pdiffusion 696 -955 696 -955 0 feedthrough
rlabel pdiffusion 703 -955 703 -955 0 feedthrough
rlabel pdiffusion 710 -955 710 -955 0 cellNo=289
rlabel pdiffusion 717 -955 717 -955 0 cellNo=292
rlabel pdiffusion 724 -955 724 -955 0 feedthrough
rlabel pdiffusion 731 -955 731 -955 0 feedthrough
rlabel pdiffusion 738 -955 738 -955 0 feedthrough
rlabel pdiffusion 745 -955 745 -955 0 cellNo=372
rlabel pdiffusion 752 -955 752 -955 0 feedthrough
rlabel pdiffusion 759 -955 759 -955 0 feedthrough
rlabel pdiffusion 766 -955 766 -955 0 feedthrough
rlabel pdiffusion 773 -955 773 -955 0 feedthrough
rlabel pdiffusion 780 -955 780 -955 0 feedthrough
rlabel pdiffusion 787 -955 787 -955 0 feedthrough
rlabel pdiffusion 794 -955 794 -955 0 feedthrough
rlabel pdiffusion 801 -955 801 -955 0 feedthrough
rlabel pdiffusion 808 -955 808 -955 0 feedthrough
rlabel pdiffusion 815 -955 815 -955 0 feedthrough
rlabel pdiffusion 822 -955 822 -955 0 cellNo=359
rlabel pdiffusion 829 -955 829 -955 0 feedthrough
rlabel pdiffusion 836 -955 836 -955 0 feedthrough
rlabel pdiffusion 843 -955 843 -955 0 feedthrough
rlabel pdiffusion 850 -955 850 -955 0 feedthrough
rlabel pdiffusion 857 -955 857 -955 0 feedthrough
rlabel pdiffusion 864 -955 864 -955 0 feedthrough
rlabel pdiffusion 871 -955 871 -955 0 feedthrough
rlabel pdiffusion 878 -955 878 -955 0 feedthrough
rlabel pdiffusion 885 -955 885 -955 0 feedthrough
rlabel pdiffusion 892 -955 892 -955 0 feedthrough
rlabel pdiffusion 899 -955 899 -955 0 feedthrough
rlabel pdiffusion 906 -955 906 -955 0 feedthrough
rlabel pdiffusion 913 -955 913 -955 0 feedthrough
rlabel pdiffusion 920 -955 920 -955 0 feedthrough
rlabel pdiffusion 927 -955 927 -955 0 feedthrough
rlabel pdiffusion 934 -955 934 -955 0 feedthrough
rlabel pdiffusion 941 -955 941 -955 0 feedthrough
rlabel pdiffusion 948 -955 948 -955 0 feedthrough
rlabel pdiffusion 955 -955 955 -955 0 feedthrough
rlabel pdiffusion 962 -955 962 -955 0 feedthrough
rlabel pdiffusion 969 -955 969 -955 0 feedthrough
rlabel pdiffusion 976 -955 976 -955 0 feedthrough
rlabel pdiffusion 983 -955 983 -955 0 feedthrough
rlabel pdiffusion 990 -955 990 -955 0 feedthrough
rlabel pdiffusion 997 -955 997 -955 0 feedthrough
rlabel pdiffusion 1004 -955 1004 -955 0 feedthrough
rlabel pdiffusion 1011 -955 1011 -955 0 feedthrough
rlabel pdiffusion 1018 -955 1018 -955 0 feedthrough
rlabel pdiffusion 1025 -955 1025 -955 0 feedthrough
rlabel pdiffusion 1032 -955 1032 -955 0 feedthrough
rlabel pdiffusion 1039 -955 1039 -955 0 feedthrough
rlabel pdiffusion 1046 -955 1046 -955 0 feedthrough
rlabel pdiffusion 1053 -955 1053 -955 0 feedthrough
rlabel pdiffusion 1060 -955 1060 -955 0 feedthrough
rlabel pdiffusion 1067 -955 1067 -955 0 feedthrough
rlabel pdiffusion 1074 -955 1074 -955 0 feedthrough
rlabel pdiffusion 1081 -955 1081 -955 0 feedthrough
rlabel pdiffusion 1088 -955 1088 -955 0 feedthrough
rlabel pdiffusion 1095 -955 1095 -955 0 feedthrough
rlabel pdiffusion 1102 -955 1102 -955 0 feedthrough
rlabel pdiffusion 1109 -955 1109 -955 0 feedthrough
rlabel pdiffusion 1116 -955 1116 -955 0 feedthrough
rlabel pdiffusion 1123 -955 1123 -955 0 feedthrough
rlabel pdiffusion 1130 -955 1130 -955 0 feedthrough
rlabel pdiffusion 1137 -955 1137 -955 0 feedthrough
rlabel pdiffusion 1144 -955 1144 -955 0 feedthrough
rlabel pdiffusion 1151 -955 1151 -955 0 feedthrough
rlabel pdiffusion 1158 -955 1158 -955 0 feedthrough
rlabel pdiffusion 1165 -955 1165 -955 0 feedthrough
rlabel pdiffusion 1172 -955 1172 -955 0 feedthrough
rlabel pdiffusion 1179 -955 1179 -955 0 feedthrough
rlabel pdiffusion 1186 -955 1186 -955 0 feedthrough
rlabel pdiffusion 1193 -955 1193 -955 0 cellNo=373
rlabel pdiffusion 1200 -955 1200 -955 0 cellNo=456
rlabel pdiffusion 1207 -955 1207 -955 0 feedthrough
rlabel pdiffusion 1438 -955 1438 -955 0 feedthrough
rlabel pdiffusion 3 -1084 3 -1084 0 cellNo=498
rlabel pdiffusion 10 -1084 10 -1084 0 feedthrough
rlabel pdiffusion 17 -1084 17 -1084 0 feedthrough
rlabel pdiffusion 24 -1084 24 -1084 0 feedthrough
rlabel pdiffusion 31 -1084 31 -1084 0 cellNo=199
rlabel pdiffusion 38 -1084 38 -1084 0 cellNo=18
rlabel pdiffusion 45 -1084 45 -1084 0 feedthrough
rlabel pdiffusion 52 -1084 52 -1084 0 cellNo=408
rlabel pdiffusion 59 -1084 59 -1084 0 feedthrough
rlabel pdiffusion 66 -1084 66 -1084 0 feedthrough
rlabel pdiffusion 73 -1084 73 -1084 0 cellNo=466
rlabel pdiffusion 80 -1084 80 -1084 0 feedthrough
rlabel pdiffusion 87 -1084 87 -1084 0 feedthrough
rlabel pdiffusion 94 -1084 94 -1084 0 cellNo=433
rlabel pdiffusion 101 -1084 101 -1084 0 cellNo=223
rlabel pdiffusion 108 -1084 108 -1084 0 feedthrough
rlabel pdiffusion 115 -1084 115 -1084 0 feedthrough
rlabel pdiffusion 122 -1084 122 -1084 0 feedthrough
rlabel pdiffusion 129 -1084 129 -1084 0 feedthrough
rlabel pdiffusion 136 -1084 136 -1084 0 feedthrough
rlabel pdiffusion 143 -1084 143 -1084 0 feedthrough
rlabel pdiffusion 150 -1084 150 -1084 0 cellNo=483
rlabel pdiffusion 157 -1084 157 -1084 0 feedthrough
rlabel pdiffusion 164 -1084 164 -1084 0 feedthrough
rlabel pdiffusion 171 -1084 171 -1084 0 feedthrough
rlabel pdiffusion 178 -1084 178 -1084 0 feedthrough
rlabel pdiffusion 185 -1084 185 -1084 0 feedthrough
rlabel pdiffusion 192 -1084 192 -1084 0 feedthrough
rlabel pdiffusion 199 -1084 199 -1084 0 feedthrough
rlabel pdiffusion 206 -1084 206 -1084 0 feedthrough
rlabel pdiffusion 213 -1084 213 -1084 0 feedthrough
rlabel pdiffusion 220 -1084 220 -1084 0 feedthrough
rlabel pdiffusion 227 -1084 227 -1084 0 feedthrough
rlabel pdiffusion 234 -1084 234 -1084 0 feedthrough
rlabel pdiffusion 241 -1084 241 -1084 0 feedthrough
rlabel pdiffusion 248 -1084 248 -1084 0 feedthrough
rlabel pdiffusion 255 -1084 255 -1084 0 feedthrough
rlabel pdiffusion 262 -1084 262 -1084 0 cellNo=15
rlabel pdiffusion 269 -1084 269 -1084 0 feedthrough
rlabel pdiffusion 276 -1084 276 -1084 0 feedthrough
rlabel pdiffusion 283 -1084 283 -1084 0 feedthrough
rlabel pdiffusion 290 -1084 290 -1084 0 feedthrough
rlabel pdiffusion 297 -1084 297 -1084 0 feedthrough
rlabel pdiffusion 304 -1084 304 -1084 0 cellNo=462
rlabel pdiffusion 311 -1084 311 -1084 0 feedthrough
rlabel pdiffusion 318 -1084 318 -1084 0 feedthrough
rlabel pdiffusion 325 -1084 325 -1084 0 feedthrough
rlabel pdiffusion 332 -1084 332 -1084 0 feedthrough
rlabel pdiffusion 339 -1084 339 -1084 0 cellNo=309
rlabel pdiffusion 346 -1084 346 -1084 0 feedthrough
rlabel pdiffusion 353 -1084 353 -1084 0 feedthrough
rlabel pdiffusion 360 -1084 360 -1084 0 feedthrough
rlabel pdiffusion 367 -1084 367 -1084 0 feedthrough
rlabel pdiffusion 374 -1084 374 -1084 0 cellNo=1
rlabel pdiffusion 381 -1084 381 -1084 0 feedthrough
rlabel pdiffusion 388 -1084 388 -1084 0 feedthrough
rlabel pdiffusion 395 -1084 395 -1084 0 feedthrough
rlabel pdiffusion 402 -1084 402 -1084 0 feedthrough
rlabel pdiffusion 409 -1084 409 -1084 0 feedthrough
rlabel pdiffusion 416 -1084 416 -1084 0 feedthrough
rlabel pdiffusion 423 -1084 423 -1084 0 feedthrough
rlabel pdiffusion 430 -1084 430 -1084 0 feedthrough
rlabel pdiffusion 437 -1084 437 -1084 0 cellNo=198
rlabel pdiffusion 444 -1084 444 -1084 0 feedthrough
rlabel pdiffusion 451 -1084 451 -1084 0 feedthrough
rlabel pdiffusion 458 -1084 458 -1084 0 feedthrough
rlabel pdiffusion 465 -1084 465 -1084 0 feedthrough
rlabel pdiffusion 472 -1084 472 -1084 0 feedthrough
rlabel pdiffusion 479 -1084 479 -1084 0 cellNo=58
rlabel pdiffusion 486 -1084 486 -1084 0 feedthrough
rlabel pdiffusion 493 -1084 493 -1084 0 cellNo=569
rlabel pdiffusion 500 -1084 500 -1084 0 cellNo=96
rlabel pdiffusion 507 -1084 507 -1084 0 feedthrough
rlabel pdiffusion 514 -1084 514 -1084 0 cellNo=27
rlabel pdiffusion 521 -1084 521 -1084 0 feedthrough
rlabel pdiffusion 528 -1084 528 -1084 0 cellNo=206
rlabel pdiffusion 535 -1084 535 -1084 0 feedthrough
rlabel pdiffusion 542 -1084 542 -1084 0 feedthrough
rlabel pdiffusion 549 -1084 549 -1084 0 feedthrough
rlabel pdiffusion 556 -1084 556 -1084 0 cellNo=379
rlabel pdiffusion 563 -1084 563 -1084 0 cellNo=472
rlabel pdiffusion 570 -1084 570 -1084 0 cellNo=43
rlabel pdiffusion 577 -1084 577 -1084 0 feedthrough
rlabel pdiffusion 584 -1084 584 -1084 0 feedthrough
rlabel pdiffusion 591 -1084 591 -1084 0 feedthrough
rlabel pdiffusion 598 -1084 598 -1084 0 feedthrough
rlabel pdiffusion 605 -1084 605 -1084 0 feedthrough
rlabel pdiffusion 612 -1084 612 -1084 0 feedthrough
rlabel pdiffusion 619 -1084 619 -1084 0 feedthrough
rlabel pdiffusion 626 -1084 626 -1084 0 cellNo=113
rlabel pdiffusion 633 -1084 633 -1084 0 cellNo=234
rlabel pdiffusion 640 -1084 640 -1084 0 feedthrough
rlabel pdiffusion 647 -1084 647 -1084 0 feedthrough
rlabel pdiffusion 654 -1084 654 -1084 0 feedthrough
rlabel pdiffusion 661 -1084 661 -1084 0 feedthrough
rlabel pdiffusion 668 -1084 668 -1084 0 feedthrough
rlabel pdiffusion 675 -1084 675 -1084 0 cellNo=436
rlabel pdiffusion 682 -1084 682 -1084 0 feedthrough
rlabel pdiffusion 689 -1084 689 -1084 0 feedthrough
rlabel pdiffusion 696 -1084 696 -1084 0 feedthrough
rlabel pdiffusion 703 -1084 703 -1084 0 feedthrough
rlabel pdiffusion 710 -1084 710 -1084 0 feedthrough
rlabel pdiffusion 717 -1084 717 -1084 0 feedthrough
rlabel pdiffusion 724 -1084 724 -1084 0 cellNo=92
rlabel pdiffusion 731 -1084 731 -1084 0 feedthrough
rlabel pdiffusion 738 -1084 738 -1084 0 feedthrough
rlabel pdiffusion 745 -1084 745 -1084 0 cellNo=2
rlabel pdiffusion 752 -1084 752 -1084 0 feedthrough
rlabel pdiffusion 759 -1084 759 -1084 0 feedthrough
rlabel pdiffusion 766 -1084 766 -1084 0 feedthrough
rlabel pdiffusion 773 -1084 773 -1084 0 feedthrough
rlabel pdiffusion 780 -1084 780 -1084 0 feedthrough
rlabel pdiffusion 787 -1084 787 -1084 0 feedthrough
rlabel pdiffusion 794 -1084 794 -1084 0 feedthrough
rlabel pdiffusion 801 -1084 801 -1084 0 feedthrough
rlabel pdiffusion 808 -1084 808 -1084 0 feedthrough
rlabel pdiffusion 815 -1084 815 -1084 0 feedthrough
rlabel pdiffusion 822 -1084 822 -1084 0 feedthrough
rlabel pdiffusion 829 -1084 829 -1084 0 feedthrough
rlabel pdiffusion 836 -1084 836 -1084 0 feedthrough
rlabel pdiffusion 843 -1084 843 -1084 0 feedthrough
rlabel pdiffusion 850 -1084 850 -1084 0 feedthrough
rlabel pdiffusion 857 -1084 857 -1084 0 feedthrough
rlabel pdiffusion 864 -1084 864 -1084 0 cellNo=130
rlabel pdiffusion 871 -1084 871 -1084 0 feedthrough
rlabel pdiffusion 878 -1084 878 -1084 0 feedthrough
rlabel pdiffusion 885 -1084 885 -1084 0 feedthrough
rlabel pdiffusion 892 -1084 892 -1084 0 feedthrough
rlabel pdiffusion 899 -1084 899 -1084 0 feedthrough
rlabel pdiffusion 906 -1084 906 -1084 0 feedthrough
rlabel pdiffusion 913 -1084 913 -1084 0 feedthrough
rlabel pdiffusion 920 -1084 920 -1084 0 feedthrough
rlabel pdiffusion 927 -1084 927 -1084 0 cellNo=567
rlabel pdiffusion 934 -1084 934 -1084 0 feedthrough
rlabel pdiffusion 941 -1084 941 -1084 0 feedthrough
rlabel pdiffusion 948 -1084 948 -1084 0 feedthrough
rlabel pdiffusion 955 -1084 955 -1084 0 feedthrough
rlabel pdiffusion 962 -1084 962 -1084 0 feedthrough
rlabel pdiffusion 969 -1084 969 -1084 0 feedthrough
rlabel pdiffusion 976 -1084 976 -1084 0 feedthrough
rlabel pdiffusion 983 -1084 983 -1084 0 feedthrough
rlabel pdiffusion 990 -1084 990 -1084 0 feedthrough
rlabel pdiffusion 997 -1084 997 -1084 0 feedthrough
rlabel pdiffusion 1004 -1084 1004 -1084 0 feedthrough
rlabel pdiffusion 1011 -1084 1011 -1084 0 feedthrough
rlabel pdiffusion 1018 -1084 1018 -1084 0 feedthrough
rlabel pdiffusion 1025 -1084 1025 -1084 0 feedthrough
rlabel pdiffusion 1032 -1084 1032 -1084 0 feedthrough
rlabel pdiffusion 1039 -1084 1039 -1084 0 feedthrough
rlabel pdiffusion 1046 -1084 1046 -1084 0 feedthrough
rlabel pdiffusion 1053 -1084 1053 -1084 0 feedthrough
rlabel pdiffusion 1060 -1084 1060 -1084 0 feedthrough
rlabel pdiffusion 1067 -1084 1067 -1084 0 feedthrough
rlabel pdiffusion 1074 -1084 1074 -1084 0 feedthrough
rlabel pdiffusion 1081 -1084 1081 -1084 0 feedthrough
rlabel pdiffusion 1088 -1084 1088 -1084 0 feedthrough
rlabel pdiffusion 1095 -1084 1095 -1084 0 feedthrough
rlabel pdiffusion 1102 -1084 1102 -1084 0 feedthrough
rlabel pdiffusion 1109 -1084 1109 -1084 0 feedthrough
rlabel pdiffusion 1116 -1084 1116 -1084 0 feedthrough
rlabel pdiffusion 1123 -1084 1123 -1084 0 feedthrough
rlabel pdiffusion 1130 -1084 1130 -1084 0 feedthrough
rlabel pdiffusion 1137 -1084 1137 -1084 0 feedthrough
rlabel pdiffusion 1144 -1084 1144 -1084 0 feedthrough
rlabel pdiffusion 1151 -1084 1151 -1084 0 feedthrough
rlabel pdiffusion 1158 -1084 1158 -1084 0 feedthrough
rlabel pdiffusion 1165 -1084 1165 -1084 0 feedthrough
rlabel pdiffusion 1172 -1084 1172 -1084 0 feedthrough
rlabel pdiffusion 1179 -1084 1179 -1084 0 feedthrough
rlabel pdiffusion 1186 -1084 1186 -1084 0 feedthrough
rlabel pdiffusion 1193 -1084 1193 -1084 0 feedthrough
rlabel pdiffusion 1200 -1084 1200 -1084 0 feedthrough
rlabel pdiffusion 1207 -1084 1207 -1084 0 feedthrough
rlabel pdiffusion 1214 -1084 1214 -1084 0 feedthrough
rlabel pdiffusion 1221 -1084 1221 -1084 0 feedthrough
rlabel pdiffusion 1228 -1084 1228 -1084 0 feedthrough
rlabel pdiffusion 1235 -1084 1235 -1084 0 feedthrough
rlabel pdiffusion 1242 -1084 1242 -1084 0 feedthrough
rlabel pdiffusion 1249 -1084 1249 -1084 0 feedthrough
rlabel pdiffusion 1256 -1084 1256 -1084 0 feedthrough
rlabel pdiffusion 1263 -1084 1263 -1084 0 feedthrough
rlabel pdiffusion 1270 -1084 1270 -1084 0 feedthrough
rlabel pdiffusion 1277 -1084 1277 -1084 0 feedthrough
rlabel pdiffusion 1284 -1084 1284 -1084 0 feedthrough
rlabel pdiffusion 1291 -1084 1291 -1084 0 feedthrough
rlabel pdiffusion 1298 -1084 1298 -1084 0 feedthrough
rlabel pdiffusion 1305 -1084 1305 -1084 0 feedthrough
rlabel pdiffusion 1312 -1084 1312 -1084 0 feedthrough
rlabel pdiffusion 1319 -1084 1319 -1084 0 feedthrough
rlabel pdiffusion 1326 -1084 1326 -1084 0 feedthrough
rlabel pdiffusion 1333 -1084 1333 -1084 0 feedthrough
rlabel pdiffusion 1340 -1084 1340 -1084 0 feedthrough
rlabel pdiffusion 1347 -1084 1347 -1084 0 feedthrough
rlabel pdiffusion 1445 -1084 1445 -1084 0 feedthrough
rlabel pdiffusion 3 -1209 3 -1209 0 cellNo=499
rlabel pdiffusion 10 -1209 10 -1209 0 feedthrough
rlabel pdiffusion 17 -1209 17 -1209 0 feedthrough
rlabel pdiffusion 24 -1209 24 -1209 0 feedthrough
rlabel pdiffusion 31 -1209 31 -1209 0 feedthrough
rlabel pdiffusion 38 -1209 38 -1209 0 feedthrough
rlabel pdiffusion 45 -1209 45 -1209 0 feedthrough
rlabel pdiffusion 52 -1209 52 -1209 0 feedthrough
rlabel pdiffusion 59 -1209 59 -1209 0 feedthrough
rlabel pdiffusion 66 -1209 66 -1209 0 feedthrough
rlabel pdiffusion 73 -1209 73 -1209 0 cellNo=85
rlabel pdiffusion 80 -1209 80 -1209 0 feedthrough
rlabel pdiffusion 87 -1209 87 -1209 0 feedthrough
rlabel pdiffusion 94 -1209 94 -1209 0 feedthrough
rlabel pdiffusion 101 -1209 101 -1209 0 cellNo=490
rlabel pdiffusion 108 -1209 108 -1209 0 feedthrough
rlabel pdiffusion 115 -1209 115 -1209 0 cellNo=265
rlabel pdiffusion 122 -1209 122 -1209 0 feedthrough
rlabel pdiffusion 129 -1209 129 -1209 0 feedthrough
rlabel pdiffusion 136 -1209 136 -1209 0 feedthrough
rlabel pdiffusion 143 -1209 143 -1209 0 feedthrough
rlabel pdiffusion 150 -1209 150 -1209 0 feedthrough
rlabel pdiffusion 157 -1209 157 -1209 0 feedthrough
rlabel pdiffusion 164 -1209 164 -1209 0 feedthrough
rlabel pdiffusion 171 -1209 171 -1209 0 feedthrough
rlabel pdiffusion 178 -1209 178 -1209 0 cellNo=364
rlabel pdiffusion 185 -1209 185 -1209 0 feedthrough
rlabel pdiffusion 192 -1209 192 -1209 0 feedthrough
rlabel pdiffusion 199 -1209 199 -1209 0 feedthrough
rlabel pdiffusion 206 -1209 206 -1209 0 feedthrough
rlabel pdiffusion 213 -1209 213 -1209 0 cellNo=529
rlabel pdiffusion 220 -1209 220 -1209 0 feedthrough
rlabel pdiffusion 227 -1209 227 -1209 0 feedthrough
rlabel pdiffusion 234 -1209 234 -1209 0 feedthrough
rlabel pdiffusion 241 -1209 241 -1209 0 feedthrough
rlabel pdiffusion 248 -1209 248 -1209 0 feedthrough
rlabel pdiffusion 255 -1209 255 -1209 0 feedthrough
rlabel pdiffusion 262 -1209 262 -1209 0 feedthrough
rlabel pdiffusion 269 -1209 269 -1209 0 feedthrough
rlabel pdiffusion 276 -1209 276 -1209 0 feedthrough
rlabel pdiffusion 283 -1209 283 -1209 0 feedthrough
rlabel pdiffusion 290 -1209 290 -1209 0 feedthrough
rlabel pdiffusion 297 -1209 297 -1209 0 feedthrough
rlabel pdiffusion 304 -1209 304 -1209 0 feedthrough
rlabel pdiffusion 311 -1209 311 -1209 0 feedthrough
rlabel pdiffusion 318 -1209 318 -1209 0 feedthrough
rlabel pdiffusion 325 -1209 325 -1209 0 feedthrough
rlabel pdiffusion 332 -1209 332 -1209 0 feedthrough
rlabel pdiffusion 339 -1209 339 -1209 0 feedthrough
rlabel pdiffusion 346 -1209 346 -1209 0 feedthrough
rlabel pdiffusion 353 -1209 353 -1209 0 feedthrough
rlabel pdiffusion 360 -1209 360 -1209 0 feedthrough
rlabel pdiffusion 367 -1209 367 -1209 0 feedthrough
rlabel pdiffusion 374 -1209 374 -1209 0 feedthrough
rlabel pdiffusion 381 -1209 381 -1209 0 feedthrough
rlabel pdiffusion 388 -1209 388 -1209 0 feedthrough
rlabel pdiffusion 395 -1209 395 -1209 0 feedthrough
rlabel pdiffusion 402 -1209 402 -1209 0 cellNo=437
rlabel pdiffusion 409 -1209 409 -1209 0 feedthrough
rlabel pdiffusion 416 -1209 416 -1209 0 feedthrough
rlabel pdiffusion 423 -1209 423 -1209 0 feedthrough
rlabel pdiffusion 430 -1209 430 -1209 0 feedthrough
rlabel pdiffusion 437 -1209 437 -1209 0 feedthrough
rlabel pdiffusion 444 -1209 444 -1209 0 feedthrough
rlabel pdiffusion 451 -1209 451 -1209 0 feedthrough
rlabel pdiffusion 458 -1209 458 -1209 0 feedthrough
rlabel pdiffusion 465 -1209 465 -1209 0 cellNo=17
rlabel pdiffusion 472 -1209 472 -1209 0 feedthrough
rlabel pdiffusion 479 -1209 479 -1209 0 feedthrough
rlabel pdiffusion 486 -1209 486 -1209 0 feedthrough
rlabel pdiffusion 493 -1209 493 -1209 0 cellNo=333
rlabel pdiffusion 500 -1209 500 -1209 0 feedthrough
rlabel pdiffusion 507 -1209 507 -1209 0 feedthrough
rlabel pdiffusion 514 -1209 514 -1209 0 feedthrough
rlabel pdiffusion 521 -1209 521 -1209 0 cellNo=84
rlabel pdiffusion 528 -1209 528 -1209 0 cellNo=283
rlabel pdiffusion 535 -1209 535 -1209 0 feedthrough
rlabel pdiffusion 542 -1209 542 -1209 0 cellNo=226
rlabel pdiffusion 549 -1209 549 -1209 0 cellNo=53
rlabel pdiffusion 556 -1209 556 -1209 0 cellNo=317
rlabel pdiffusion 563 -1209 563 -1209 0 feedthrough
rlabel pdiffusion 570 -1209 570 -1209 0 feedthrough
rlabel pdiffusion 577 -1209 577 -1209 0 feedthrough
rlabel pdiffusion 584 -1209 584 -1209 0 feedthrough
rlabel pdiffusion 591 -1209 591 -1209 0 feedthrough
rlabel pdiffusion 598 -1209 598 -1209 0 cellNo=402
rlabel pdiffusion 605 -1209 605 -1209 0 cellNo=453
rlabel pdiffusion 612 -1209 612 -1209 0 feedthrough
rlabel pdiffusion 619 -1209 619 -1209 0 feedthrough
rlabel pdiffusion 626 -1209 626 -1209 0 cellNo=547
rlabel pdiffusion 633 -1209 633 -1209 0 cellNo=64
rlabel pdiffusion 640 -1209 640 -1209 0 feedthrough
rlabel pdiffusion 647 -1209 647 -1209 0 cellNo=560
rlabel pdiffusion 654 -1209 654 -1209 0 feedthrough
rlabel pdiffusion 661 -1209 661 -1209 0 feedthrough
rlabel pdiffusion 668 -1209 668 -1209 0 feedthrough
rlabel pdiffusion 675 -1209 675 -1209 0 feedthrough
rlabel pdiffusion 682 -1209 682 -1209 0 cellNo=311
rlabel pdiffusion 689 -1209 689 -1209 0 feedthrough
rlabel pdiffusion 696 -1209 696 -1209 0 feedthrough
rlabel pdiffusion 703 -1209 703 -1209 0 feedthrough
rlabel pdiffusion 710 -1209 710 -1209 0 cellNo=471
rlabel pdiffusion 717 -1209 717 -1209 0 feedthrough
rlabel pdiffusion 724 -1209 724 -1209 0 feedthrough
rlabel pdiffusion 731 -1209 731 -1209 0 cellNo=577
rlabel pdiffusion 738 -1209 738 -1209 0 feedthrough
rlabel pdiffusion 745 -1209 745 -1209 0 cellNo=6
rlabel pdiffusion 752 -1209 752 -1209 0 cellNo=220
rlabel pdiffusion 759 -1209 759 -1209 0 cellNo=525
rlabel pdiffusion 766 -1209 766 -1209 0 cellNo=102
rlabel pdiffusion 773 -1209 773 -1209 0 feedthrough
rlabel pdiffusion 780 -1209 780 -1209 0 feedthrough
rlabel pdiffusion 787 -1209 787 -1209 0 feedthrough
rlabel pdiffusion 794 -1209 794 -1209 0 cellNo=28
rlabel pdiffusion 801 -1209 801 -1209 0 feedthrough
rlabel pdiffusion 808 -1209 808 -1209 0 feedthrough
rlabel pdiffusion 815 -1209 815 -1209 0 feedthrough
rlabel pdiffusion 822 -1209 822 -1209 0 feedthrough
rlabel pdiffusion 829 -1209 829 -1209 0 feedthrough
rlabel pdiffusion 836 -1209 836 -1209 0 feedthrough
rlabel pdiffusion 843 -1209 843 -1209 0 cellNo=148
rlabel pdiffusion 850 -1209 850 -1209 0 feedthrough
rlabel pdiffusion 857 -1209 857 -1209 0 feedthrough
rlabel pdiffusion 864 -1209 864 -1209 0 feedthrough
rlabel pdiffusion 871 -1209 871 -1209 0 feedthrough
rlabel pdiffusion 878 -1209 878 -1209 0 feedthrough
rlabel pdiffusion 885 -1209 885 -1209 0 feedthrough
rlabel pdiffusion 892 -1209 892 -1209 0 feedthrough
rlabel pdiffusion 899 -1209 899 -1209 0 feedthrough
rlabel pdiffusion 906 -1209 906 -1209 0 feedthrough
rlabel pdiffusion 913 -1209 913 -1209 0 feedthrough
rlabel pdiffusion 920 -1209 920 -1209 0 feedthrough
rlabel pdiffusion 927 -1209 927 -1209 0 feedthrough
rlabel pdiffusion 934 -1209 934 -1209 0 feedthrough
rlabel pdiffusion 941 -1209 941 -1209 0 feedthrough
rlabel pdiffusion 948 -1209 948 -1209 0 feedthrough
rlabel pdiffusion 955 -1209 955 -1209 0 feedthrough
rlabel pdiffusion 962 -1209 962 -1209 0 feedthrough
rlabel pdiffusion 969 -1209 969 -1209 0 feedthrough
rlabel pdiffusion 976 -1209 976 -1209 0 feedthrough
rlabel pdiffusion 983 -1209 983 -1209 0 feedthrough
rlabel pdiffusion 990 -1209 990 -1209 0 feedthrough
rlabel pdiffusion 997 -1209 997 -1209 0 feedthrough
rlabel pdiffusion 1004 -1209 1004 -1209 0 feedthrough
rlabel pdiffusion 1011 -1209 1011 -1209 0 feedthrough
rlabel pdiffusion 1018 -1209 1018 -1209 0 feedthrough
rlabel pdiffusion 1025 -1209 1025 -1209 0 feedthrough
rlabel pdiffusion 1032 -1209 1032 -1209 0 feedthrough
rlabel pdiffusion 1039 -1209 1039 -1209 0 feedthrough
rlabel pdiffusion 1046 -1209 1046 -1209 0 feedthrough
rlabel pdiffusion 1053 -1209 1053 -1209 0 feedthrough
rlabel pdiffusion 1060 -1209 1060 -1209 0 feedthrough
rlabel pdiffusion 1067 -1209 1067 -1209 0 feedthrough
rlabel pdiffusion 1074 -1209 1074 -1209 0 feedthrough
rlabel pdiffusion 1081 -1209 1081 -1209 0 feedthrough
rlabel pdiffusion 1088 -1209 1088 -1209 0 feedthrough
rlabel pdiffusion 1095 -1209 1095 -1209 0 feedthrough
rlabel pdiffusion 1102 -1209 1102 -1209 0 feedthrough
rlabel pdiffusion 1109 -1209 1109 -1209 0 feedthrough
rlabel pdiffusion 1116 -1209 1116 -1209 0 feedthrough
rlabel pdiffusion 1123 -1209 1123 -1209 0 feedthrough
rlabel pdiffusion 1130 -1209 1130 -1209 0 feedthrough
rlabel pdiffusion 1137 -1209 1137 -1209 0 feedthrough
rlabel pdiffusion 1144 -1209 1144 -1209 0 feedthrough
rlabel pdiffusion 1151 -1209 1151 -1209 0 feedthrough
rlabel pdiffusion 1158 -1209 1158 -1209 0 feedthrough
rlabel pdiffusion 1165 -1209 1165 -1209 0 feedthrough
rlabel pdiffusion 1172 -1209 1172 -1209 0 feedthrough
rlabel pdiffusion 1179 -1209 1179 -1209 0 feedthrough
rlabel pdiffusion 1186 -1209 1186 -1209 0 feedthrough
rlabel pdiffusion 1193 -1209 1193 -1209 0 feedthrough
rlabel pdiffusion 1200 -1209 1200 -1209 0 feedthrough
rlabel pdiffusion 1207 -1209 1207 -1209 0 feedthrough
rlabel pdiffusion 1214 -1209 1214 -1209 0 feedthrough
rlabel pdiffusion 1221 -1209 1221 -1209 0 feedthrough
rlabel pdiffusion 1228 -1209 1228 -1209 0 feedthrough
rlabel pdiffusion 1235 -1209 1235 -1209 0 feedthrough
rlabel pdiffusion 1242 -1209 1242 -1209 0 feedthrough
rlabel pdiffusion 1249 -1209 1249 -1209 0 feedthrough
rlabel pdiffusion 1256 -1209 1256 -1209 0 feedthrough
rlabel pdiffusion 1263 -1209 1263 -1209 0 feedthrough
rlabel pdiffusion 1270 -1209 1270 -1209 0 feedthrough
rlabel pdiffusion 1277 -1209 1277 -1209 0 feedthrough
rlabel pdiffusion 1284 -1209 1284 -1209 0 feedthrough
rlabel pdiffusion 1291 -1209 1291 -1209 0 feedthrough
rlabel pdiffusion 1298 -1209 1298 -1209 0 feedthrough
rlabel pdiffusion 1305 -1209 1305 -1209 0 feedthrough
rlabel pdiffusion 1312 -1209 1312 -1209 0 feedthrough
rlabel pdiffusion 1319 -1209 1319 -1209 0 feedthrough
rlabel pdiffusion 1326 -1209 1326 -1209 0 feedthrough
rlabel pdiffusion 1333 -1209 1333 -1209 0 feedthrough
rlabel pdiffusion 1340 -1209 1340 -1209 0 feedthrough
rlabel pdiffusion 1347 -1209 1347 -1209 0 feedthrough
rlabel pdiffusion 1354 -1209 1354 -1209 0 feedthrough
rlabel pdiffusion 1361 -1209 1361 -1209 0 feedthrough
rlabel pdiffusion 1368 -1209 1368 -1209 0 feedthrough
rlabel pdiffusion 1375 -1209 1375 -1209 0 feedthrough
rlabel pdiffusion 1452 -1209 1452 -1209 0 feedthrough
rlabel pdiffusion 3 -1330 3 -1330 0 feedthrough
rlabel pdiffusion 10 -1330 10 -1330 0 feedthrough
rlabel pdiffusion 17 -1330 17 -1330 0 feedthrough
rlabel pdiffusion 24 -1330 24 -1330 0 feedthrough
rlabel pdiffusion 31 -1330 31 -1330 0 feedthrough
rlabel pdiffusion 38 -1330 38 -1330 0 feedthrough
rlabel pdiffusion 45 -1330 45 -1330 0 feedthrough
rlabel pdiffusion 52 -1330 52 -1330 0 feedthrough
rlabel pdiffusion 59 -1330 59 -1330 0 cellNo=150
rlabel pdiffusion 66 -1330 66 -1330 0 cellNo=507
rlabel pdiffusion 73 -1330 73 -1330 0 feedthrough
rlabel pdiffusion 80 -1330 80 -1330 0 cellNo=146
rlabel pdiffusion 87 -1330 87 -1330 0 cellNo=181
rlabel pdiffusion 94 -1330 94 -1330 0 feedthrough
rlabel pdiffusion 101 -1330 101 -1330 0 feedthrough
rlabel pdiffusion 108 -1330 108 -1330 0 feedthrough
rlabel pdiffusion 115 -1330 115 -1330 0 feedthrough
rlabel pdiffusion 122 -1330 122 -1330 0 cellNo=86
rlabel pdiffusion 129 -1330 129 -1330 0 feedthrough
rlabel pdiffusion 136 -1330 136 -1330 0 cellNo=136
rlabel pdiffusion 143 -1330 143 -1330 0 feedthrough
rlabel pdiffusion 150 -1330 150 -1330 0 feedthrough
rlabel pdiffusion 157 -1330 157 -1330 0 feedthrough
rlabel pdiffusion 164 -1330 164 -1330 0 cellNo=121
rlabel pdiffusion 171 -1330 171 -1330 0 cellNo=543
rlabel pdiffusion 178 -1330 178 -1330 0 feedthrough
rlabel pdiffusion 185 -1330 185 -1330 0 feedthrough
rlabel pdiffusion 192 -1330 192 -1330 0 feedthrough
rlabel pdiffusion 199 -1330 199 -1330 0 feedthrough
rlabel pdiffusion 206 -1330 206 -1330 0 feedthrough
rlabel pdiffusion 213 -1330 213 -1330 0 feedthrough
rlabel pdiffusion 220 -1330 220 -1330 0 feedthrough
rlabel pdiffusion 227 -1330 227 -1330 0 feedthrough
rlabel pdiffusion 234 -1330 234 -1330 0 feedthrough
rlabel pdiffusion 241 -1330 241 -1330 0 feedthrough
rlabel pdiffusion 248 -1330 248 -1330 0 feedthrough
rlabel pdiffusion 255 -1330 255 -1330 0 feedthrough
rlabel pdiffusion 262 -1330 262 -1330 0 feedthrough
rlabel pdiffusion 269 -1330 269 -1330 0 feedthrough
rlabel pdiffusion 276 -1330 276 -1330 0 feedthrough
rlabel pdiffusion 283 -1330 283 -1330 0 feedthrough
rlabel pdiffusion 290 -1330 290 -1330 0 feedthrough
rlabel pdiffusion 297 -1330 297 -1330 0 feedthrough
rlabel pdiffusion 304 -1330 304 -1330 0 feedthrough
rlabel pdiffusion 311 -1330 311 -1330 0 feedthrough
rlabel pdiffusion 318 -1330 318 -1330 0 feedthrough
rlabel pdiffusion 325 -1330 325 -1330 0 feedthrough
rlabel pdiffusion 332 -1330 332 -1330 0 feedthrough
rlabel pdiffusion 339 -1330 339 -1330 0 feedthrough
rlabel pdiffusion 346 -1330 346 -1330 0 feedthrough
rlabel pdiffusion 353 -1330 353 -1330 0 feedthrough
rlabel pdiffusion 360 -1330 360 -1330 0 feedthrough
rlabel pdiffusion 367 -1330 367 -1330 0 cellNo=106
rlabel pdiffusion 374 -1330 374 -1330 0 cellNo=451
rlabel pdiffusion 381 -1330 381 -1330 0 feedthrough
rlabel pdiffusion 388 -1330 388 -1330 0 cellNo=161
rlabel pdiffusion 395 -1330 395 -1330 0 feedthrough
rlabel pdiffusion 402 -1330 402 -1330 0 feedthrough
rlabel pdiffusion 409 -1330 409 -1330 0 feedthrough
rlabel pdiffusion 416 -1330 416 -1330 0 cellNo=134
rlabel pdiffusion 423 -1330 423 -1330 0 feedthrough
rlabel pdiffusion 430 -1330 430 -1330 0 cellNo=143
rlabel pdiffusion 437 -1330 437 -1330 0 feedthrough
rlabel pdiffusion 444 -1330 444 -1330 0 cellNo=388
rlabel pdiffusion 451 -1330 451 -1330 0 feedthrough
rlabel pdiffusion 458 -1330 458 -1330 0 feedthrough
rlabel pdiffusion 465 -1330 465 -1330 0 feedthrough
rlabel pdiffusion 472 -1330 472 -1330 0 feedthrough
rlabel pdiffusion 479 -1330 479 -1330 0 feedthrough
rlabel pdiffusion 486 -1330 486 -1330 0 feedthrough
rlabel pdiffusion 493 -1330 493 -1330 0 feedthrough
rlabel pdiffusion 500 -1330 500 -1330 0 feedthrough
rlabel pdiffusion 507 -1330 507 -1330 0 feedthrough
rlabel pdiffusion 514 -1330 514 -1330 0 feedthrough
rlabel pdiffusion 521 -1330 521 -1330 0 feedthrough
rlabel pdiffusion 528 -1330 528 -1330 0 feedthrough
rlabel pdiffusion 535 -1330 535 -1330 0 feedthrough
rlabel pdiffusion 542 -1330 542 -1330 0 cellNo=582
rlabel pdiffusion 549 -1330 549 -1330 0 feedthrough
rlabel pdiffusion 556 -1330 556 -1330 0 feedthrough
rlabel pdiffusion 563 -1330 563 -1330 0 feedthrough
rlabel pdiffusion 570 -1330 570 -1330 0 cellNo=376
rlabel pdiffusion 577 -1330 577 -1330 0 feedthrough
rlabel pdiffusion 584 -1330 584 -1330 0 feedthrough
rlabel pdiffusion 591 -1330 591 -1330 0 feedthrough
rlabel pdiffusion 598 -1330 598 -1330 0 feedthrough
rlabel pdiffusion 605 -1330 605 -1330 0 feedthrough
rlabel pdiffusion 612 -1330 612 -1330 0 cellNo=71
rlabel pdiffusion 619 -1330 619 -1330 0 cellNo=390
rlabel pdiffusion 626 -1330 626 -1330 0 feedthrough
rlabel pdiffusion 633 -1330 633 -1330 0 cellNo=470
rlabel pdiffusion 640 -1330 640 -1330 0 feedthrough
rlabel pdiffusion 647 -1330 647 -1330 0 feedthrough
rlabel pdiffusion 654 -1330 654 -1330 0 feedthrough
rlabel pdiffusion 661 -1330 661 -1330 0 feedthrough
rlabel pdiffusion 668 -1330 668 -1330 0 feedthrough
rlabel pdiffusion 675 -1330 675 -1330 0 feedthrough
rlabel pdiffusion 682 -1330 682 -1330 0 cellNo=157
rlabel pdiffusion 689 -1330 689 -1330 0 feedthrough
rlabel pdiffusion 696 -1330 696 -1330 0 cellNo=374
rlabel pdiffusion 703 -1330 703 -1330 0 cellNo=83
rlabel pdiffusion 710 -1330 710 -1330 0 feedthrough
rlabel pdiffusion 717 -1330 717 -1330 0 cellNo=118
rlabel pdiffusion 724 -1330 724 -1330 0 feedthrough
rlabel pdiffusion 731 -1330 731 -1330 0 cellNo=9
rlabel pdiffusion 738 -1330 738 -1330 0 feedthrough
rlabel pdiffusion 745 -1330 745 -1330 0 feedthrough
rlabel pdiffusion 752 -1330 752 -1330 0 feedthrough
rlabel pdiffusion 759 -1330 759 -1330 0 feedthrough
rlabel pdiffusion 766 -1330 766 -1330 0 feedthrough
rlabel pdiffusion 773 -1330 773 -1330 0 feedthrough
rlabel pdiffusion 780 -1330 780 -1330 0 feedthrough
rlabel pdiffusion 787 -1330 787 -1330 0 feedthrough
rlabel pdiffusion 794 -1330 794 -1330 0 feedthrough
rlabel pdiffusion 801 -1330 801 -1330 0 feedthrough
rlabel pdiffusion 808 -1330 808 -1330 0 feedthrough
rlabel pdiffusion 815 -1330 815 -1330 0 cellNo=229
rlabel pdiffusion 822 -1330 822 -1330 0 feedthrough
rlabel pdiffusion 829 -1330 829 -1330 0 feedthrough
rlabel pdiffusion 836 -1330 836 -1330 0 feedthrough
rlabel pdiffusion 843 -1330 843 -1330 0 feedthrough
rlabel pdiffusion 850 -1330 850 -1330 0 feedthrough
rlabel pdiffusion 857 -1330 857 -1330 0 feedthrough
rlabel pdiffusion 864 -1330 864 -1330 0 cellNo=377
rlabel pdiffusion 871 -1330 871 -1330 0 feedthrough
rlabel pdiffusion 878 -1330 878 -1330 0 feedthrough
rlabel pdiffusion 885 -1330 885 -1330 0 feedthrough
rlabel pdiffusion 892 -1330 892 -1330 0 feedthrough
rlabel pdiffusion 899 -1330 899 -1330 0 cellNo=49
rlabel pdiffusion 906 -1330 906 -1330 0 feedthrough
rlabel pdiffusion 913 -1330 913 -1330 0 cellNo=108
rlabel pdiffusion 920 -1330 920 -1330 0 feedthrough
rlabel pdiffusion 927 -1330 927 -1330 0 feedthrough
rlabel pdiffusion 934 -1330 934 -1330 0 feedthrough
rlabel pdiffusion 941 -1330 941 -1330 0 feedthrough
rlabel pdiffusion 948 -1330 948 -1330 0 feedthrough
rlabel pdiffusion 955 -1330 955 -1330 0 feedthrough
rlabel pdiffusion 962 -1330 962 -1330 0 feedthrough
rlabel pdiffusion 969 -1330 969 -1330 0 feedthrough
rlabel pdiffusion 976 -1330 976 -1330 0 feedthrough
rlabel pdiffusion 983 -1330 983 -1330 0 feedthrough
rlabel pdiffusion 990 -1330 990 -1330 0 feedthrough
rlabel pdiffusion 997 -1330 997 -1330 0 feedthrough
rlabel pdiffusion 1004 -1330 1004 -1330 0 feedthrough
rlabel pdiffusion 1011 -1330 1011 -1330 0 feedthrough
rlabel pdiffusion 1018 -1330 1018 -1330 0 feedthrough
rlabel pdiffusion 1025 -1330 1025 -1330 0 feedthrough
rlabel pdiffusion 1032 -1330 1032 -1330 0 feedthrough
rlabel pdiffusion 1039 -1330 1039 -1330 0 feedthrough
rlabel pdiffusion 1046 -1330 1046 -1330 0 feedthrough
rlabel pdiffusion 1053 -1330 1053 -1330 0 feedthrough
rlabel pdiffusion 1060 -1330 1060 -1330 0 feedthrough
rlabel pdiffusion 1067 -1330 1067 -1330 0 feedthrough
rlabel pdiffusion 1074 -1330 1074 -1330 0 feedthrough
rlabel pdiffusion 1081 -1330 1081 -1330 0 feedthrough
rlabel pdiffusion 1088 -1330 1088 -1330 0 feedthrough
rlabel pdiffusion 1095 -1330 1095 -1330 0 feedthrough
rlabel pdiffusion 1102 -1330 1102 -1330 0 feedthrough
rlabel pdiffusion 1109 -1330 1109 -1330 0 feedthrough
rlabel pdiffusion 1116 -1330 1116 -1330 0 feedthrough
rlabel pdiffusion 1123 -1330 1123 -1330 0 feedthrough
rlabel pdiffusion 1130 -1330 1130 -1330 0 feedthrough
rlabel pdiffusion 1137 -1330 1137 -1330 0 feedthrough
rlabel pdiffusion 1144 -1330 1144 -1330 0 feedthrough
rlabel pdiffusion 1151 -1330 1151 -1330 0 feedthrough
rlabel pdiffusion 1158 -1330 1158 -1330 0 feedthrough
rlabel pdiffusion 1165 -1330 1165 -1330 0 feedthrough
rlabel pdiffusion 1172 -1330 1172 -1330 0 feedthrough
rlabel pdiffusion 1179 -1330 1179 -1330 0 feedthrough
rlabel pdiffusion 1186 -1330 1186 -1330 0 feedthrough
rlabel pdiffusion 1193 -1330 1193 -1330 0 feedthrough
rlabel pdiffusion 1200 -1330 1200 -1330 0 feedthrough
rlabel pdiffusion 1207 -1330 1207 -1330 0 feedthrough
rlabel pdiffusion 1214 -1330 1214 -1330 0 feedthrough
rlabel pdiffusion 1221 -1330 1221 -1330 0 feedthrough
rlabel pdiffusion 1228 -1330 1228 -1330 0 feedthrough
rlabel pdiffusion 1235 -1330 1235 -1330 0 feedthrough
rlabel pdiffusion 1242 -1330 1242 -1330 0 feedthrough
rlabel pdiffusion 1249 -1330 1249 -1330 0 feedthrough
rlabel pdiffusion 1256 -1330 1256 -1330 0 feedthrough
rlabel pdiffusion 1263 -1330 1263 -1330 0 feedthrough
rlabel pdiffusion 1270 -1330 1270 -1330 0 feedthrough
rlabel pdiffusion 1277 -1330 1277 -1330 0 feedthrough
rlabel pdiffusion 1284 -1330 1284 -1330 0 feedthrough
rlabel pdiffusion 1291 -1330 1291 -1330 0 feedthrough
rlabel pdiffusion 1298 -1330 1298 -1330 0 feedthrough
rlabel pdiffusion 1305 -1330 1305 -1330 0 feedthrough
rlabel pdiffusion 1312 -1330 1312 -1330 0 feedthrough
rlabel pdiffusion 1319 -1330 1319 -1330 0 feedthrough
rlabel pdiffusion 1326 -1330 1326 -1330 0 feedthrough
rlabel pdiffusion 1333 -1330 1333 -1330 0 feedthrough
rlabel pdiffusion 1340 -1330 1340 -1330 0 feedthrough
rlabel pdiffusion 1347 -1330 1347 -1330 0 feedthrough
rlabel pdiffusion 1354 -1330 1354 -1330 0 feedthrough
rlabel pdiffusion 1361 -1330 1361 -1330 0 feedthrough
rlabel pdiffusion 1368 -1330 1368 -1330 0 feedthrough
rlabel pdiffusion 1375 -1330 1375 -1330 0 feedthrough
rlabel pdiffusion 1382 -1330 1382 -1330 0 feedthrough
rlabel pdiffusion 1389 -1330 1389 -1330 0 feedthrough
rlabel pdiffusion 1459 -1330 1459 -1330 0 feedthrough
rlabel pdiffusion 3 -1455 3 -1455 0 feedthrough
rlabel pdiffusion 10 -1455 10 -1455 0 feedthrough
rlabel pdiffusion 17 -1455 17 -1455 0 feedthrough
rlabel pdiffusion 24 -1455 24 -1455 0 feedthrough
rlabel pdiffusion 31 -1455 31 -1455 0 cellNo=512
rlabel pdiffusion 38 -1455 38 -1455 0 feedthrough
rlabel pdiffusion 45 -1455 45 -1455 0 feedthrough
rlabel pdiffusion 52 -1455 52 -1455 0 feedthrough
rlabel pdiffusion 59 -1455 59 -1455 0 feedthrough
rlabel pdiffusion 66 -1455 66 -1455 0 feedthrough
rlabel pdiffusion 73 -1455 73 -1455 0 feedthrough
rlabel pdiffusion 80 -1455 80 -1455 0 cellNo=583
rlabel pdiffusion 87 -1455 87 -1455 0 feedthrough
rlabel pdiffusion 94 -1455 94 -1455 0 feedthrough
rlabel pdiffusion 101 -1455 101 -1455 0 feedthrough
rlabel pdiffusion 108 -1455 108 -1455 0 feedthrough
rlabel pdiffusion 115 -1455 115 -1455 0 feedthrough
rlabel pdiffusion 122 -1455 122 -1455 0 feedthrough
rlabel pdiffusion 129 -1455 129 -1455 0 cellNo=365
rlabel pdiffusion 136 -1455 136 -1455 0 feedthrough
rlabel pdiffusion 143 -1455 143 -1455 0 feedthrough
rlabel pdiffusion 150 -1455 150 -1455 0 cellNo=3
rlabel pdiffusion 157 -1455 157 -1455 0 feedthrough
rlabel pdiffusion 164 -1455 164 -1455 0 feedthrough
rlabel pdiffusion 171 -1455 171 -1455 0 feedthrough
rlabel pdiffusion 178 -1455 178 -1455 0 feedthrough
rlabel pdiffusion 185 -1455 185 -1455 0 feedthrough
rlabel pdiffusion 192 -1455 192 -1455 0 feedthrough
rlabel pdiffusion 199 -1455 199 -1455 0 feedthrough
rlabel pdiffusion 206 -1455 206 -1455 0 feedthrough
rlabel pdiffusion 213 -1455 213 -1455 0 feedthrough
rlabel pdiffusion 220 -1455 220 -1455 0 feedthrough
rlabel pdiffusion 227 -1455 227 -1455 0 feedthrough
rlabel pdiffusion 234 -1455 234 -1455 0 feedthrough
rlabel pdiffusion 241 -1455 241 -1455 0 feedthrough
rlabel pdiffusion 248 -1455 248 -1455 0 feedthrough
rlabel pdiffusion 255 -1455 255 -1455 0 feedthrough
rlabel pdiffusion 262 -1455 262 -1455 0 feedthrough
rlabel pdiffusion 269 -1455 269 -1455 0 feedthrough
rlabel pdiffusion 276 -1455 276 -1455 0 feedthrough
rlabel pdiffusion 283 -1455 283 -1455 0 feedthrough
rlabel pdiffusion 290 -1455 290 -1455 0 feedthrough
rlabel pdiffusion 297 -1455 297 -1455 0 feedthrough
rlabel pdiffusion 304 -1455 304 -1455 0 feedthrough
rlabel pdiffusion 311 -1455 311 -1455 0 feedthrough
rlabel pdiffusion 318 -1455 318 -1455 0 cellNo=514
rlabel pdiffusion 325 -1455 325 -1455 0 feedthrough
rlabel pdiffusion 332 -1455 332 -1455 0 feedthrough
rlabel pdiffusion 339 -1455 339 -1455 0 feedthrough
rlabel pdiffusion 346 -1455 346 -1455 0 feedthrough
rlabel pdiffusion 353 -1455 353 -1455 0 feedthrough
rlabel pdiffusion 360 -1455 360 -1455 0 feedthrough
rlabel pdiffusion 367 -1455 367 -1455 0 feedthrough
rlabel pdiffusion 374 -1455 374 -1455 0 feedthrough
rlabel pdiffusion 381 -1455 381 -1455 0 feedthrough
rlabel pdiffusion 388 -1455 388 -1455 0 feedthrough
rlabel pdiffusion 395 -1455 395 -1455 0 cellNo=171
rlabel pdiffusion 402 -1455 402 -1455 0 feedthrough
rlabel pdiffusion 409 -1455 409 -1455 0 cellNo=79
rlabel pdiffusion 416 -1455 416 -1455 0 feedthrough
rlabel pdiffusion 423 -1455 423 -1455 0 feedthrough
rlabel pdiffusion 430 -1455 430 -1455 0 feedthrough
rlabel pdiffusion 437 -1455 437 -1455 0 feedthrough
rlabel pdiffusion 444 -1455 444 -1455 0 cellNo=600
rlabel pdiffusion 451 -1455 451 -1455 0 feedthrough
rlabel pdiffusion 458 -1455 458 -1455 0 cellNo=31
rlabel pdiffusion 465 -1455 465 -1455 0 feedthrough
rlabel pdiffusion 472 -1455 472 -1455 0 feedthrough
rlabel pdiffusion 479 -1455 479 -1455 0 feedthrough
rlabel pdiffusion 486 -1455 486 -1455 0 feedthrough
rlabel pdiffusion 493 -1455 493 -1455 0 feedthrough
rlabel pdiffusion 500 -1455 500 -1455 0 feedthrough
rlabel pdiffusion 507 -1455 507 -1455 0 cellNo=593
rlabel pdiffusion 514 -1455 514 -1455 0 feedthrough
rlabel pdiffusion 521 -1455 521 -1455 0 cellNo=129
rlabel pdiffusion 528 -1455 528 -1455 0 feedthrough
rlabel pdiffusion 535 -1455 535 -1455 0 cellNo=111
rlabel pdiffusion 542 -1455 542 -1455 0 feedthrough
rlabel pdiffusion 549 -1455 549 -1455 0 cellNo=243
rlabel pdiffusion 556 -1455 556 -1455 0 feedthrough
rlabel pdiffusion 563 -1455 563 -1455 0 cellNo=579
rlabel pdiffusion 570 -1455 570 -1455 0 feedthrough
rlabel pdiffusion 577 -1455 577 -1455 0 feedthrough
rlabel pdiffusion 584 -1455 584 -1455 0 feedthrough
rlabel pdiffusion 591 -1455 591 -1455 0 feedthrough
rlabel pdiffusion 598 -1455 598 -1455 0 feedthrough
rlabel pdiffusion 605 -1455 605 -1455 0 feedthrough
rlabel pdiffusion 612 -1455 612 -1455 0 feedthrough
rlabel pdiffusion 619 -1455 619 -1455 0 feedthrough
rlabel pdiffusion 626 -1455 626 -1455 0 feedthrough
rlabel pdiffusion 633 -1455 633 -1455 0 feedthrough
rlabel pdiffusion 640 -1455 640 -1455 0 cellNo=203
rlabel pdiffusion 647 -1455 647 -1455 0 cellNo=444
rlabel pdiffusion 654 -1455 654 -1455 0 feedthrough
rlabel pdiffusion 661 -1455 661 -1455 0 feedthrough
rlabel pdiffusion 668 -1455 668 -1455 0 feedthrough
rlabel pdiffusion 675 -1455 675 -1455 0 feedthrough
rlabel pdiffusion 682 -1455 682 -1455 0 feedthrough
rlabel pdiffusion 689 -1455 689 -1455 0 feedthrough
rlabel pdiffusion 696 -1455 696 -1455 0 feedthrough
rlabel pdiffusion 703 -1455 703 -1455 0 feedthrough
rlabel pdiffusion 710 -1455 710 -1455 0 feedthrough
rlabel pdiffusion 717 -1455 717 -1455 0 feedthrough
rlabel pdiffusion 724 -1455 724 -1455 0 cellNo=24
rlabel pdiffusion 731 -1455 731 -1455 0 feedthrough
rlabel pdiffusion 738 -1455 738 -1455 0 feedthrough
rlabel pdiffusion 745 -1455 745 -1455 0 cellNo=389
rlabel pdiffusion 752 -1455 752 -1455 0 feedthrough
rlabel pdiffusion 759 -1455 759 -1455 0 feedthrough
rlabel pdiffusion 766 -1455 766 -1455 0 feedthrough
rlabel pdiffusion 773 -1455 773 -1455 0 feedthrough
rlabel pdiffusion 780 -1455 780 -1455 0 cellNo=559
rlabel pdiffusion 787 -1455 787 -1455 0 feedthrough
rlabel pdiffusion 794 -1455 794 -1455 0 cellNo=217
rlabel pdiffusion 801 -1455 801 -1455 0 feedthrough
rlabel pdiffusion 808 -1455 808 -1455 0 feedthrough
rlabel pdiffusion 815 -1455 815 -1455 0 cellNo=526
rlabel pdiffusion 822 -1455 822 -1455 0 cellNo=497
rlabel pdiffusion 829 -1455 829 -1455 0 cellNo=11
rlabel pdiffusion 836 -1455 836 -1455 0 feedthrough
rlabel pdiffusion 843 -1455 843 -1455 0 feedthrough
rlabel pdiffusion 850 -1455 850 -1455 0 cellNo=131
rlabel pdiffusion 857 -1455 857 -1455 0 cellNo=324
rlabel pdiffusion 864 -1455 864 -1455 0 cellNo=293
rlabel pdiffusion 871 -1455 871 -1455 0 feedthrough
rlabel pdiffusion 878 -1455 878 -1455 0 feedthrough
rlabel pdiffusion 885 -1455 885 -1455 0 cellNo=14
rlabel pdiffusion 892 -1455 892 -1455 0 feedthrough
rlabel pdiffusion 899 -1455 899 -1455 0 feedthrough
rlabel pdiffusion 906 -1455 906 -1455 0 feedthrough
rlabel pdiffusion 913 -1455 913 -1455 0 feedthrough
rlabel pdiffusion 920 -1455 920 -1455 0 feedthrough
rlabel pdiffusion 927 -1455 927 -1455 0 feedthrough
rlabel pdiffusion 934 -1455 934 -1455 0 feedthrough
rlabel pdiffusion 941 -1455 941 -1455 0 feedthrough
rlabel pdiffusion 948 -1455 948 -1455 0 feedthrough
rlabel pdiffusion 955 -1455 955 -1455 0 feedthrough
rlabel pdiffusion 962 -1455 962 -1455 0 feedthrough
rlabel pdiffusion 969 -1455 969 -1455 0 feedthrough
rlabel pdiffusion 976 -1455 976 -1455 0 feedthrough
rlabel pdiffusion 983 -1455 983 -1455 0 feedthrough
rlabel pdiffusion 990 -1455 990 -1455 0 feedthrough
rlabel pdiffusion 997 -1455 997 -1455 0 feedthrough
rlabel pdiffusion 1004 -1455 1004 -1455 0 feedthrough
rlabel pdiffusion 1011 -1455 1011 -1455 0 feedthrough
rlabel pdiffusion 1018 -1455 1018 -1455 0 feedthrough
rlabel pdiffusion 1025 -1455 1025 -1455 0 feedthrough
rlabel pdiffusion 1032 -1455 1032 -1455 0 feedthrough
rlabel pdiffusion 1039 -1455 1039 -1455 0 feedthrough
rlabel pdiffusion 1046 -1455 1046 -1455 0 feedthrough
rlabel pdiffusion 1053 -1455 1053 -1455 0 feedthrough
rlabel pdiffusion 1060 -1455 1060 -1455 0 feedthrough
rlabel pdiffusion 1067 -1455 1067 -1455 0 feedthrough
rlabel pdiffusion 1074 -1455 1074 -1455 0 feedthrough
rlabel pdiffusion 1081 -1455 1081 -1455 0 feedthrough
rlabel pdiffusion 1088 -1455 1088 -1455 0 feedthrough
rlabel pdiffusion 1095 -1455 1095 -1455 0 feedthrough
rlabel pdiffusion 1102 -1455 1102 -1455 0 feedthrough
rlabel pdiffusion 1109 -1455 1109 -1455 0 feedthrough
rlabel pdiffusion 1116 -1455 1116 -1455 0 feedthrough
rlabel pdiffusion 1123 -1455 1123 -1455 0 feedthrough
rlabel pdiffusion 1130 -1455 1130 -1455 0 feedthrough
rlabel pdiffusion 1137 -1455 1137 -1455 0 feedthrough
rlabel pdiffusion 1144 -1455 1144 -1455 0 feedthrough
rlabel pdiffusion 1151 -1455 1151 -1455 0 feedthrough
rlabel pdiffusion 1158 -1455 1158 -1455 0 feedthrough
rlabel pdiffusion 1165 -1455 1165 -1455 0 feedthrough
rlabel pdiffusion 1172 -1455 1172 -1455 0 feedthrough
rlabel pdiffusion 1179 -1455 1179 -1455 0 feedthrough
rlabel pdiffusion 1186 -1455 1186 -1455 0 feedthrough
rlabel pdiffusion 1193 -1455 1193 -1455 0 feedthrough
rlabel pdiffusion 1200 -1455 1200 -1455 0 feedthrough
rlabel pdiffusion 1207 -1455 1207 -1455 0 feedthrough
rlabel pdiffusion 1214 -1455 1214 -1455 0 feedthrough
rlabel pdiffusion 1221 -1455 1221 -1455 0 feedthrough
rlabel pdiffusion 1228 -1455 1228 -1455 0 feedthrough
rlabel pdiffusion 1235 -1455 1235 -1455 0 feedthrough
rlabel pdiffusion 1242 -1455 1242 -1455 0 feedthrough
rlabel pdiffusion 1249 -1455 1249 -1455 0 feedthrough
rlabel pdiffusion 1256 -1455 1256 -1455 0 feedthrough
rlabel pdiffusion 1263 -1455 1263 -1455 0 feedthrough
rlabel pdiffusion 1270 -1455 1270 -1455 0 feedthrough
rlabel pdiffusion 1277 -1455 1277 -1455 0 feedthrough
rlabel pdiffusion 1284 -1455 1284 -1455 0 feedthrough
rlabel pdiffusion 1291 -1455 1291 -1455 0 feedthrough
rlabel pdiffusion 1298 -1455 1298 -1455 0 feedthrough
rlabel pdiffusion 1305 -1455 1305 -1455 0 feedthrough
rlabel pdiffusion 1312 -1455 1312 -1455 0 feedthrough
rlabel pdiffusion 1319 -1455 1319 -1455 0 feedthrough
rlabel pdiffusion 1326 -1455 1326 -1455 0 feedthrough
rlabel pdiffusion 1333 -1455 1333 -1455 0 feedthrough
rlabel pdiffusion 1340 -1455 1340 -1455 0 feedthrough
rlabel pdiffusion 1347 -1455 1347 -1455 0 feedthrough
rlabel pdiffusion 1354 -1455 1354 -1455 0 feedthrough
rlabel pdiffusion 1361 -1455 1361 -1455 0 feedthrough
rlabel pdiffusion 1368 -1455 1368 -1455 0 feedthrough
rlabel pdiffusion 1375 -1455 1375 -1455 0 feedthrough
rlabel pdiffusion 1382 -1455 1382 -1455 0 feedthrough
rlabel pdiffusion 1389 -1455 1389 -1455 0 feedthrough
rlabel pdiffusion 1396 -1455 1396 -1455 0 feedthrough
rlabel pdiffusion 1403 -1455 1403 -1455 0 feedthrough
rlabel pdiffusion 1410 -1455 1410 -1455 0 feedthrough
rlabel pdiffusion 1417 -1455 1417 -1455 0 feedthrough
rlabel pdiffusion 1424 -1455 1424 -1455 0 feedthrough
rlabel pdiffusion 1431 -1455 1431 -1455 0 feedthrough
rlabel pdiffusion 1438 -1455 1438 -1455 0 feedthrough
rlabel pdiffusion 1445 -1455 1445 -1455 0 feedthrough
rlabel pdiffusion 1452 -1455 1452 -1455 0 cellNo=286
rlabel pdiffusion 1459 -1455 1459 -1455 0 feedthrough
rlabel pdiffusion 1466 -1455 1466 -1455 0 feedthrough
rlabel pdiffusion 3 -1592 3 -1592 0 feedthrough
rlabel pdiffusion 10 -1592 10 -1592 0 cellNo=564
rlabel pdiffusion 17 -1592 17 -1592 0 cellNo=407
rlabel pdiffusion 24 -1592 24 -1592 0 feedthrough
rlabel pdiffusion 31 -1592 31 -1592 0 feedthrough
rlabel pdiffusion 38 -1592 38 -1592 0 cellNo=352
rlabel pdiffusion 45 -1592 45 -1592 0 feedthrough
rlabel pdiffusion 52 -1592 52 -1592 0 cellNo=193
rlabel pdiffusion 59 -1592 59 -1592 0 feedthrough
rlabel pdiffusion 66 -1592 66 -1592 0 feedthrough
rlabel pdiffusion 73 -1592 73 -1592 0 feedthrough
rlabel pdiffusion 80 -1592 80 -1592 0 feedthrough
rlabel pdiffusion 87 -1592 87 -1592 0 cellNo=279
rlabel pdiffusion 94 -1592 94 -1592 0 feedthrough
rlabel pdiffusion 101 -1592 101 -1592 0 cellNo=105
rlabel pdiffusion 108 -1592 108 -1592 0 feedthrough
rlabel pdiffusion 115 -1592 115 -1592 0 cellNo=273
rlabel pdiffusion 122 -1592 122 -1592 0 feedthrough
rlabel pdiffusion 129 -1592 129 -1592 0 feedthrough
rlabel pdiffusion 136 -1592 136 -1592 0 cellNo=501
rlabel pdiffusion 143 -1592 143 -1592 0 cellNo=139
rlabel pdiffusion 150 -1592 150 -1592 0 feedthrough
rlabel pdiffusion 157 -1592 157 -1592 0 feedthrough
rlabel pdiffusion 164 -1592 164 -1592 0 feedthrough
rlabel pdiffusion 171 -1592 171 -1592 0 feedthrough
rlabel pdiffusion 178 -1592 178 -1592 0 cellNo=67
rlabel pdiffusion 185 -1592 185 -1592 0 feedthrough
rlabel pdiffusion 192 -1592 192 -1592 0 feedthrough
rlabel pdiffusion 199 -1592 199 -1592 0 feedthrough
rlabel pdiffusion 206 -1592 206 -1592 0 feedthrough
rlabel pdiffusion 213 -1592 213 -1592 0 feedthrough
rlabel pdiffusion 220 -1592 220 -1592 0 cellNo=533
rlabel pdiffusion 227 -1592 227 -1592 0 feedthrough
rlabel pdiffusion 234 -1592 234 -1592 0 feedthrough
rlabel pdiffusion 241 -1592 241 -1592 0 feedthrough
rlabel pdiffusion 248 -1592 248 -1592 0 feedthrough
rlabel pdiffusion 255 -1592 255 -1592 0 feedthrough
rlabel pdiffusion 262 -1592 262 -1592 0 feedthrough
rlabel pdiffusion 269 -1592 269 -1592 0 feedthrough
rlabel pdiffusion 276 -1592 276 -1592 0 feedthrough
rlabel pdiffusion 283 -1592 283 -1592 0 feedthrough
rlabel pdiffusion 290 -1592 290 -1592 0 feedthrough
rlabel pdiffusion 297 -1592 297 -1592 0 feedthrough
rlabel pdiffusion 304 -1592 304 -1592 0 feedthrough
rlabel pdiffusion 311 -1592 311 -1592 0 feedthrough
rlabel pdiffusion 318 -1592 318 -1592 0 feedthrough
rlabel pdiffusion 325 -1592 325 -1592 0 feedthrough
rlabel pdiffusion 332 -1592 332 -1592 0 feedthrough
rlabel pdiffusion 339 -1592 339 -1592 0 feedthrough
rlabel pdiffusion 346 -1592 346 -1592 0 feedthrough
rlabel pdiffusion 353 -1592 353 -1592 0 feedthrough
rlabel pdiffusion 360 -1592 360 -1592 0 feedthrough
rlabel pdiffusion 367 -1592 367 -1592 0 feedthrough
rlabel pdiffusion 374 -1592 374 -1592 0 feedthrough
rlabel pdiffusion 381 -1592 381 -1592 0 feedthrough
rlabel pdiffusion 388 -1592 388 -1592 0 feedthrough
rlabel pdiffusion 395 -1592 395 -1592 0 feedthrough
rlabel pdiffusion 402 -1592 402 -1592 0 cellNo=50
rlabel pdiffusion 409 -1592 409 -1592 0 feedthrough
rlabel pdiffusion 416 -1592 416 -1592 0 feedthrough
rlabel pdiffusion 423 -1592 423 -1592 0 feedthrough
rlabel pdiffusion 430 -1592 430 -1592 0 cellNo=74
rlabel pdiffusion 437 -1592 437 -1592 0 feedthrough
rlabel pdiffusion 444 -1592 444 -1592 0 feedthrough
rlabel pdiffusion 451 -1592 451 -1592 0 feedthrough
rlabel pdiffusion 458 -1592 458 -1592 0 cellNo=246
rlabel pdiffusion 465 -1592 465 -1592 0 feedthrough
rlabel pdiffusion 472 -1592 472 -1592 0 feedthrough
rlabel pdiffusion 479 -1592 479 -1592 0 feedthrough
rlabel pdiffusion 486 -1592 486 -1592 0 cellNo=147
rlabel pdiffusion 493 -1592 493 -1592 0 cellNo=384
rlabel pdiffusion 500 -1592 500 -1592 0 feedthrough
rlabel pdiffusion 507 -1592 507 -1592 0 feedthrough
rlabel pdiffusion 514 -1592 514 -1592 0 feedthrough
rlabel pdiffusion 521 -1592 521 -1592 0 cellNo=114
rlabel pdiffusion 528 -1592 528 -1592 0 feedthrough
rlabel pdiffusion 535 -1592 535 -1592 0 cellNo=356
rlabel pdiffusion 542 -1592 542 -1592 0 feedthrough
rlabel pdiffusion 549 -1592 549 -1592 0 feedthrough
rlabel pdiffusion 556 -1592 556 -1592 0 cellNo=406
rlabel pdiffusion 563 -1592 563 -1592 0 feedthrough
rlabel pdiffusion 570 -1592 570 -1592 0 cellNo=123
rlabel pdiffusion 577 -1592 577 -1592 0 feedthrough
rlabel pdiffusion 584 -1592 584 -1592 0 feedthrough
rlabel pdiffusion 591 -1592 591 -1592 0 feedthrough
rlabel pdiffusion 598 -1592 598 -1592 0 feedthrough
rlabel pdiffusion 605 -1592 605 -1592 0 feedthrough
rlabel pdiffusion 612 -1592 612 -1592 0 feedthrough
rlabel pdiffusion 619 -1592 619 -1592 0 cellNo=556
rlabel pdiffusion 626 -1592 626 -1592 0 feedthrough
rlabel pdiffusion 633 -1592 633 -1592 0 feedthrough
rlabel pdiffusion 640 -1592 640 -1592 0 feedthrough
rlabel pdiffusion 647 -1592 647 -1592 0 feedthrough
rlabel pdiffusion 654 -1592 654 -1592 0 feedthrough
rlabel pdiffusion 661 -1592 661 -1592 0 cellNo=210
rlabel pdiffusion 668 -1592 668 -1592 0 feedthrough
rlabel pdiffusion 675 -1592 675 -1592 0 feedthrough
rlabel pdiffusion 682 -1592 682 -1592 0 feedthrough
rlabel pdiffusion 689 -1592 689 -1592 0 feedthrough
rlabel pdiffusion 696 -1592 696 -1592 0 feedthrough
rlabel pdiffusion 703 -1592 703 -1592 0 cellNo=355
rlabel pdiffusion 710 -1592 710 -1592 0 feedthrough
rlabel pdiffusion 717 -1592 717 -1592 0 feedthrough
rlabel pdiffusion 724 -1592 724 -1592 0 feedthrough
rlabel pdiffusion 731 -1592 731 -1592 0 feedthrough
rlabel pdiffusion 738 -1592 738 -1592 0 feedthrough
rlabel pdiffusion 745 -1592 745 -1592 0 feedthrough
rlabel pdiffusion 752 -1592 752 -1592 0 feedthrough
rlabel pdiffusion 759 -1592 759 -1592 0 feedthrough
rlabel pdiffusion 766 -1592 766 -1592 0 feedthrough
rlabel pdiffusion 773 -1592 773 -1592 0 feedthrough
rlabel pdiffusion 780 -1592 780 -1592 0 feedthrough
rlabel pdiffusion 787 -1592 787 -1592 0 feedthrough
rlabel pdiffusion 794 -1592 794 -1592 0 feedthrough
rlabel pdiffusion 801 -1592 801 -1592 0 cellNo=405
rlabel pdiffusion 808 -1592 808 -1592 0 feedthrough
rlabel pdiffusion 815 -1592 815 -1592 0 feedthrough
rlabel pdiffusion 822 -1592 822 -1592 0 feedthrough
rlabel pdiffusion 829 -1592 829 -1592 0 cellNo=397
rlabel pdiffusion 836 -1592 836 -1592 0 feedthrough
rlabel pdiffusion 843 -1592 843 -1592 0 feedthrough
rlabel pdiffusion 850 -1592 850 -1592 0 feedthrough
rlabel pdiffusion 857 -1592 857 -1592 0 cellNo=93
rlabel pdiffusion 864 -1592 864 -1592 0 feedthrough
rlabel pdiffusion 871 -1592 871 -1592 0 feedthrough
rlabel pdiffusion 878 -1592 878 -1592 0 feedthrough
rlabel pdiffusion 885 -1592 885 -1592 0 feedthrough
rlabel pdiffusion 892 -1592 892 -1592 0 cellNo=585
rlabel pdiffusion 899 -1592 899 -1592 0 feedthrough
rlabel pdiffusion 906 -1592 906 -1592 0 feedthrough
rlabel pdiffusion 913 -1592 913 -1592 0 feedthrough
rlabel pdiffusion 920 -1592 920 -1592 0 feedthrough
rlabel pdiffusion 927 -1592 927 -1592 0 feedthrough
rlabel pdiffusion 934 -1592 934 -1592 0 feedthrough
rlabel pdiffusion 941 -1592 941 -1592 0 feedthrough
rlabel pdiffusion 948 -1592 948 -1592 0 feedthrough
rlabel pdiffusion 955 -1592 955 -1592 0 feedthrough
rlabel pdiffusion 962 -1592 962 -1592 0 feedthrough
rlabel pdiffusion 969 -1592 969 -1592 0 feedthrough
rlabel pdiffusion 976 -1592 976 -1592 0 feedthrough
rlabel pdiffusion 983 -1592 983 -1592 0 feedthrough
rlabel pdiffusion 990 -1592 990 -1592 0 feedthrough
rlabel pdiffusion 997 -1592 997 -1592 0 feedthrough
rlabel pdiffusion 1004 -1592 1004 -1592 0 feedthrough
rlabel pdiffusion 1011 -1592 1011 -1592 0 feedthrough
rlabel pdiffusion 1018 -1592 1018 -1592 0 feedthrough
rlabel pdiffusion 1025 -1592 1025 -1592 0 feedthrough
rlabel pdiffusion 1032 -1592 1032 -1592 0 feedthrough
rlabel pdiffusion 1039 -1592 1039 -1592 0 feedthrough
rlabel pdiffusion 1046 -1592 1046 -1592 0 cellNo=195
rlabel pdiffusion 1053 -1592 1053 -1592 0 feedthrough
rlabel pdiffusion 1060 -1592 1060 -1592 0 feedthrough
rlabel pdiffusion 1067 -1592 1067 -1592 0 feedthrough
rlabel pdiffusion 1074 -1592 1074 -1592 0 feedthrough
rlabel pdiffusion 1081 -1592 1081 -1592 0 feedthrough
rlabel pdiffusion 1088 -1592 1088 -1592 0 feedthrough
rlabel pdiffusion 1095 -1592 1095 -1592 0 feedthrough
rlabel pdiffusion 1102 -1592 1102 -1592 0 feedthrough
rlabel pdiffusion 1109 -1592 1109 -1592 0 feedthrough
rlabel pdiffusion 1116 -1592 1116 -1592 0 feedthrough
rlabel pdiffusion 1123 -1592 1123 -1592 0 feedthrough
rlabel pdiffusion 1130 -1592 1130 -1592 0 feedthrough
rlabel pdiffusion 1137 -1592 1137 -1592 0 feedthrough
rlabel pdiffusion 1144 -1592 1144 -1592 0 feedthrough
rlabel pdiffusion 1151 -1592 1151 -1592 0 feedthrough
rlabel pdiffusion 1158 -1592 1158 -1592 0 feedthrough
rlabel pdiffusion 1165 -1592 1165 -1592 0 feedthrough
rlabel pdiffusion 1172 -1592 1172 -1592 0 feedthrough
rlabel pdiffusion 1179 -1592 1179 -1592 0 feedthrough
rlabel pdiffusion 1186 -1592 1186 -1592 0 feedthrough
rlabel pdiffusion 1193 -1592 1193 -1592 0 feedthrough
rlabel pdiffusion 1200 -1592 1200 -1592 0 feedthrough
rlabel pdiffusion 1207 -1592 1207 -1592 0 feedthrough
rlabel pdiffusion 1214 -1592 1214 -1592 0 feedthrough
rlabel pdiffusion 1221 -1592 1221 -1592 0 feedthrough
rlabel pdiffusion 1228 -1592 1228 -1592 0 feedthrough
rlabel pdiffusion 1235 -1592 1235 -1592 0 feedthrough
rlabel pdiffusion 1242 -1592 1242 -1592 0 feedthrough
rlabel pdiffusion 1249 -1592 1249 -1592 0 feedthrough
rlabel pdiffusion 1256 -1592 1256 -1592 0 feedthrough
rlabel pdiffusion 1263 -1592 1263 -1592 0 feedthrough
rlabel pdiffusion 1270 -1592 1270 -1592 0 feedthrough
rlabel pdiffusion 1277 -1592 1277 -1592 0 feedthrough
rlabel pdiffusion 1284 -1592 1284 -1592 0 feedthrough
rlabel pdiffusion 1291 -1592 1291 -1592 0 feedthrough
rlabel pdiffusion 1298 -1592 1298 -1592 0 feedthrough
rlabel pdiffusion 1305 -1592 1305 -1592 0 feedthrough
rlabel pdiffusion 1312 -1592 1312 -1592 0 feedthrough
rlabel pdiffusion 1319 -1592 1319 -1592 0 feedthrough
rlabel pdiffusion 1326 -1592 1326 -1592 0 feedthrough
rlabel pdiffusion 1333 -1592 1333 -1592 0 feedthrough
rlabel pdiffusion 1340 -1592 1340 -1592 0 feedthrough
rlabel pdiffusion 1347 -1592 1347 -1592 0 feedthrough
rlabel pdiffusion 1354 -1592 1354 -1592 0 feedthrough
rlabel pdiffusion 3 -1723 3 -1723 0 feedthrough
rlabel pdiffusion 10 -1723 10 -1723 0 feedthrough
rlabel pdiffusion 17 -1723 17 -1723 0 cellNo=580
rlabel pdiffusion 24 -1723 24 -1723 0 cellNo=496
rlabel pdiffusion 31 -1723 31 -1723 0 cellNo=455
rlabel pdiffusion 38 -1723 38 -1723 0 feedthrough
rlabel pdiffusion 45 -1723 45 -1723 0 cellNo=115
rlabel pdiffusion 52 -1723 52 -1723 0 cellNo=555
rlabel pdiffusion 59 -1723 59 -1723 0 feedthrough
rlabel pdiffusion 66 -1723 66 -1723 0 feedthrough
rlabel pdiffusion 73 -1723 73 -1723 0 feedthrough
rlabel pdiffusion 80 -1723 80 -1723 0 feedthrough
rlabel pdiffusion 87 -1723 87 -1723 0 feedthrough
rlabel pdiffusion 94 -1723 94 -1723 0 cellNo=190
rlabel pdiffusion 101 -1723 101 -1723 0 feedthrough
rlabel pdiffusion 108 -1723 108 -1723 0 cellNo=428
rlabel pdiffusion 115 -1723 115 -1723 0 feedthrough
rlabel pdiffusion 122 -1723 122 -1723 0 feedthrough
rlabel pdiffusion 129 -1723 129 -1723 0 feedthrough
rlabel pdiffusion 136 -1723 136 -1723 0 feedthrough
rlabel pdiffusion 143 -1723 143 -1723 0 feedthrough
rlabel pdiffusion 150 -1723 150 -1723 0 cellNo=452
rlabel pdiffusion 157 -1723 157 -1723 0 cellNo=5
rlabel pdiffusion 164 -1723 164 -1723 0 feedthrough
rlabel pdiffusion 171 -1723 171 -1723 0 feedthrough
rlabel pdiffusion 178 -1723 178 -1723 0 feedthrough
rlabel pdiffusion 185 -1723 185 -1723 0 feedthrough
rlabel pdiffusion 192 -1723 192 -1723 0 cellNo=587
rlabel pdiffusion 199 -1723 199 -1723 0 feedthrough
rlabel pdiffusion 206 -1723 206 -1723 0 feedthrough
rlabel pdiffusion 213 -1723 213 -1723 0 feedthrough
rlabel pdiffusion 220 -1723 220 -1723 0 feedthrough
rlabel pdiffusion 227 -1723 227 -1723 0 feedthrough
rlabel pdiffusion 234 -1723 234 -1723 0 feedthrough
rlabel pdiffusion 241 -1723 241 -1723 0 feedthrough
rlabel pdiffusion 248 -1723 248 -1723 0 feedthrough
rlabel pdiffusion 255 -1723 255 -1723 0 feedthrough
rlabel pdiffusion 262 -1723 262 -1723 0 feedthrough
rlabel pdiffusion 269 -1723 269 -1723 0 feedthrough
rlabel pdiffusion 276 -1723 276 -1723 0 feedthrough
rlabel pdiffusion 283 -1723 283 -1723 0 feedthrough
rlabel pdiffusion 290 -1723 290 -1723 0 feedthrough
rlabel pdiffusion 297 -1723 297 -1723 0 feedthrough
rlabel pdiffusion 304 -1723 304 -1723 0 feedthrough
rlabel pdiffusion 311 -1723 311 -1723 0 feedthrough
rlabel pdiffusion 318 -1723 318 -1723 0 cellNo=187
rlabel pdiffusion 325 -1723 325 -1723 0 feedthrough
rlabel pdiffusion 332 -1723 332 -1723 0 feedthrough
rlabel pdiffusion 339 -1723 339 -1723 0 feedthrough
rlabel pdiffusion 346 -1723 346 -1723 0 feedthrough
rlabel pdiffusion 353 -1723 353 -1723 0 feedthrough
rlabel pdiffusion 360 -1723 360 -1723 0 feedthrough
rlabel pdiffusion 367 -1723 367 -1723 0 feedthrough
rlabel pdiffusion 374 -1723 374 -1723 0 cellNo=238
rlabel pdiffusion 381 -1723 381 -1723 0 feedthrough
rlabel pdiffusion 388 -1723 388 -1723 0 feedthrough
rlabel pdiffusion 395 -1723 395 -1723 0 feedthrough
rlabel pdiffusion 402 -1723 402 -1723 0 cellNo=509
rlabel pdiffusion 409 -1723 409 -1723 0 feedthrough
rlabel pdiffusion 416 -1723 416 -1723 0 feedthrough
rlabel pdiffusion 423 -1723 423 -1723 0 feedthrough
rlabel pdiffusion 430 -1723 430 -1723 0 feedthrough
rlabel pdiffusion 437 -1723 437 -1723 0 feedthrough
rlabel pdiffusion 444 -1723 444 -1723 0 feedthrough
rlabel pdiffusion 451 -1723 451 -1723 0 feedthrough
rlabel pdiffusion 458 -1723 458 -1723 0 cellNo=439
rlabel pdiffusion 465 -1723 465 -1723 0 feedthrough
rlabel pdiffusion 472 -1723 472 -1723 0 feedthrough
rlabel pdiffusion 479 -1723 479 -1723 0 feedthrough
rlabel pdiffusion 486 -1723 486 -1723 0 cellNo=572
rlabel pdiffusion 493 -1723 493 -1723 0 feedthrough
rlabel pdiffusion 500 -1723 500 -1723 0 feedthrough
rlabel pdiffusion 507 -1723 507 -1723 0 feedthrough
rlabel pdiffusion 514 -1723 514 -1723 0 feedthrough
rlabel pdiffusion 521 -1723 521 -1723 0 cellNo=16
rlabel pdiffusion 528 -1723 528 -1723 0 feedthrough
rlabel pdiffusion 535 -1723 535 -1723 0 feedthrough
rlabel pdiffusion 542 -1723 542 -1723 0 feedthrough
rlabel pdiffusion 549 -1723 549 -1723 0 cellNo=576
rlabel pdiffusion 556 -1723 556 -1723 0 cellNo=7
rlabel pdiffusion 563 -1723 563 -1723 0 feedthrough
rlabel pdiffusion 570 -1723 570 -1723 0 feedthrough
rlabel pdiffusion 577 -1723 577 -1723 0 feedthrough
rlabel pdiffusion 584 -1723 584 -1723 0 feedthrough
rlabel pdiffusion 591 -1723 591 -1723 0 feedthrough
rlabel pdiffusion 598 -1723 598 -1723 0 feedthrough
rlabel pdiffusion 605 -1723 605 -1723 0 feedthrough
rlabel pdiffusion 612 -1723 612 -1723 0 feedthrough
rlabel pdiffusion 619 -1723 619 -1723 0 feedthrough
rlabel pdiffusion 626 -1723 626 -1723 0 feedthrough
rlabel pdiffusion 633 -1723 633 -1723 0 feedthrough
rlabel pdiffusion 640 -1723 640 -1723 0 feedthrough
rlabel pdiffusion 647 -1723 647 -1723 0 feedthrough
rlabel pdiffusion 654 -1723 654 -1723 0 feedthrough
rlabel pdiffusion 661 -1723 661 -1723 0 feedthrough
rlabel pdiffusion 668 -1723 668 -1723 0 cellNo=584
rlabel pdiffusion 675 -1723 675 -1723 0 feedthrough
rlabel pdiffusion 682 -1723 682 -1723 0 feedthrough
rlabel pdiffusion 689 -1723 689 -1723 0 feedthrough
rlabel pdiffusion 696 -1723 696 -1723 0 feedthrough
rlabel pdiffusion 703 -1723 703 -1723 0 feedthrough
rlabel pdiffusion 710 -1723 710 -1723 0 feedthrough
rlabel pdiffusion 717 -1723 717 -1723 0 feedthrough
rlabel pdiffusion 724 -1723 724 -1723 0 feedthrough
rlabel pdiffusion 731 -1723 731 -1723 0 feedthrough
rlabel pdiffusion 738 -1723 738 -1723 0 feedthrough
rlabel pdiffusion 745 -1723 745 -1723 0 cellNo=336
rlabel pdiffusion 752 -1723 752 -1723 0 cellNo=76
rlabel pdiffusion 759 -1723 759 -1723 0 feedthrough
rlabel pdiffusion 766 -1723 766 -1723 0 feedthrough
rlabel pdiffusion 773 -1723 773 -1723 0 cellNo=91
rlabel pdiffusion 780 -1723 780 -1723 0 feedthrough
rlabel pdiffusion 787 -1723 787 -1723 0 feedthrough
rlabel pdiffusion 794 -1723 794 -1723 0 feedthrough
rlabel pdiffusion 801 -1723 801 -1723 0 feedthrough
rlabel pdiffusion 808 -1723 808 -1723 0 feedthrough
rlabel pdiffusion 815 -1723 815 -1723 0 feedthrough
rlabel pdiffusion 822 -1723 822 -1723 0 feedthrough
rlabel pdiffusion 829 -1723 829 -1723 0 feedthrough
rlabel pdiffusion 836 -1723 836 -1723 0 feedthrough
rlabel pdiffusion 843 -1723 843 -1723 0 feedthrough
rlabel pdiffusion 850 -1723 850 -1723 0 feedthrough
rlabel pdiffusion 857 -1723 857 -1723 0 feedthrough
rlabel pdiffusion 864 -1723 864 -1723 0 feedthrough
rlabel pdiffusion 871 -1723 871 -1723 0 feedthrough
rlabel pdiffusion 878 -1723 878 -1723 0 feedthrough
rlabel pdiffusion 885 -1723 885 -1723 0 feedthrough
rlabel pdiffusion 892 -1723 892 -1723 0 cellNo=561
rlabel pdiffusion 899 -1723 899 -1723 0 cellNo=254
rlabel pdiffusion 906 -1723 906 -1723 0 feedthrough
rlabel pdiffusion 913 -1723 913 -1723 0 feedthrough
rlabel pdiffusion 920 -1723 920 -1723 0 feedthrough
rlabel pdiffusion 927 -1723 927 -1723 0 feedthrough
rlabel pdiffusion 934 -1723 934 -1723 0 feedthrough
rlabel pdiffusion 941 -1723 941 -1723 0 cellNo=245
rlabel pdiffusion 948 -1723 948 -1723 0 feedthrough
rlabel pdiffusion 955 -1723 955 -1723 0 feedthrough
rlabel pdiffusion 962 -1723 962 -1723 0 feedthrough
rlabel pdiffusion 969 -1723 969 -1723 0 feedthrough
rlabel pdiffusion 976 -1723 976 -1723 0 feedthrough
rlabel pdiffusion 983 -1723 983 -1723 0 feedthrough
rlabel pdiffusion 990 -1723 990 -1723 0 feedthrough
rlabel pdiffusion 997 -1723 997 -1723 0 feedthrough
rlabel pdiffusion 1004 -1723 1004 -1723 0 feedthrough
rlabel pdiffusion 1011 -1723 1011 -1723 0 feedthrough
rlabel pdiffusion 1018 -1723 1018 -1723 0 feedthrough
rlabel pdiffusion 1025 -1723 1025 -1723 0 feedthrough
rlabel pdiffusion 1032 -1723 1032 -1723 0 feedthrough
rlabel pdiffusion 1039 -1723 1039 -1723 0 feedthrough
rlabel pdiffusion 1046 -1723 1046 -1723 0 feedthrough
rlabel pdiffusion 1053 -1723 1053 -1723 0 feedthrough
rlabel pdiffusion 1060 -1723 1060 -1723 0 feedthrough
rlabel pdiffusion 1067 -1723 1067 -1723 0 cellNo=351
rlabel pdiffusion 1074 -1723 1074 -1723 0 feedthrough
rlabel pdiffusion 1081 -1723 1081 -1723 0 feedthrough
rlabel pdiffusion 1088 -1723 1088 -1723 0 feedthrough
rlabel pdiffusion 1095 -1723 1095 -1723 0 feedthrough
rlabel pdiffusion 1102 -1723 1102 -1723 0 feedthrough
rlabel pdiffusion 1109 -1723 1109 -1723 0 feedthrough
rlabel pdiffusion 1116 -1723 1116 -1723 0 feedthrough
rlabel pdiffusion 1123 -1723 1123 -1723 0 cellNo=47
rlabel pdiffusion 1130 -1723 1130 -1723 0 feedthrough
rlabel pdiffusion 1137 -1723 1137 -1723 0 feedthrough
rlabel pdiffusion 1144 -1723 1144 -1723 0 feedthrough
rlabel pdiffusion 1151 -1723 1151 -1723 0 feedthrough
rlabel pdiffusion 1158 -1723 1158 -1723 0 feedthrough
rlabel pdiffusion 1165 -1723 1165 -1723 0 feedthrough
rlabel pdiffusion 1172 -1723 1172 -1723 0 feedthrough
rlabel pdiffusion 1179 -1723 1179 -1723 0 feedthrough
rlabel pdiffusion 1186 -1723 1186 -1723 0 feedthrough
rlabel pdiffusion 1193 -1723 1193 -1723 0 feedthrough
rlabel pdiffusion 1200 -1723 1200 -1723 0 feedthrough
rlabel pdiffusion 1207 -1723 1207 -1723 0 feedthrough
rlabel pdiffusion 1214 -1723 1214 -1723 0 feedthrough
rlabel pdiffusion 1221 -1723 1221 -1723 0 feedthrough
rlabel pdiffusion 1228 -1723 1228 -1723 0 feedthrough
rlabel pdiffusion 1235 -1723 1235 -1723 0 feedthrough
rlabel pdiffusion 1242 -1723 1242 -1723 0 feedthrough
rlabel pdiffusion 1249 -1723 1249 -1723 0 feedthrough
rlabel pdiffusion 1256 -1723 1256 -1723 0 feedthrough
rlabel pdiffusion 1263 -1723 1263 -1723 0 feedthrough
rlabel pdiffusion 1270 -1723 1270 -1723 0 feedthrough
rlabel pdiffusion 1277 -1723 1277 -1723 0 feedthrough
rlabel pdiffusion 1284 -1723 1284 -1723 0 feedthrough
rlabel pdiffusion 1291 -1723 1291 -1723 0 feedthrough
rlabel pdiffusion 1298 -1723 1298 -1723 0 feedthrough
rlabel pdiffusion 1305 -1723 1305 -1723 0 feedthrough
rlabel pdiffusion 1312 -1723 1312 -1723 0 feedthrough
rlabel pdiffusion 1319 -1723 1319 -1723 0 feedthrough
rlabel pdiffusion 1326 -1723 1326 -1723 0 cellNo=221
rlabel pdiffusion 3 -1842 3 -1842 0 feedthrough
rlabel pdiffusion 10 -1842 10 -1842 0 feedthrough
rlabel pdiffusion 17 -1842 17 -1842 0 feedthrough
rlabel pdiffusion 24 -1842 24 -1842 0 cellNo=513
rlabel pdiffusion 31 -1842 31 -1842 0 feedthrough
rlabel pdiffusion 38 -1842 38 -1842 0 cellNo=209
rlabel pdiffusion 45 -1842 45 -1842 0 cellNo=544
rlabel pdiffusion 52 -1842 52 -1842 0 cellNo=323
rlabel pdiffusion 59 -1842 59 -1842 0 feedthrough
rlabel pdiffusion 66 -1842 66 -1842 0 cellNo=81
rlabel pdiffusion 73 -1842 73 -1842 0 feedthrough
rlabel pdiffusion 80 -1842 80 -1842 0 feedthrough
rlabel pdiffusion 87 -1842 87 -1842 0 feedthrough
rlabel pdiffusion 94 -1842 94 -1842 0 feedthrough
rlabel pdiffusion 101 -1842 101 -1842 0 feedthrough
rlabel pdiffusion 108 -1842 108 -1842 0 feedthrough
rlabel pdiffusion 115 -1842 115 -1842 0 cellNo=440
rlabel pdiffusion 122 -1842 122 -1842 0 feedthrough
rlabel pdiffusion 129 -1842 129 -1842 0 feedthrough
rlabel pdiffusion 136 -1842 136 -1842 0 cellNo=266
rlabel pdiffusion 143 -1842 143 -1842 0 feedthrough
rlabel pdiffusion 150 -1842 150 -1842 0 cellNo=188
rlabel pdiffusion 157 -1842 157 -1842 0 feedthrough
rlabel pdiffusion 164 -1842 164 -1842 0 feedthrough
rlabel pdiffusion 171 -1842 171 -1842 0 feedthrough
rlabel pdiffusion 178 -1842 178 -1842 0 feedthrough
rlabel pdiffusion 185 -1842 185 -1842 0 feedthrough
rlabel pdiffusion 192 -1842 192 -1842 0 feedthrough
rlabel pdiffusion 199 -1842 199 -1842 0 feedthrough
rlabel pdiffusion 206 -1842 206 -1842 0 feedthrough
rlabel pdiffusion 213 -1842 213 -1842 0 feedthrough
rlabel pdiffusion 220 -1842 220 -1842 0 feedthrough
rlabel pdiffusion 227 -1842 227 -1842 0 feedthrough
rlabel pdiffusion 234 -1842 234 -1842 0 feedthrough
rlabel pdiffusion 241 -1842 241 -1842 0 feedthrough
rlabel pdiffusion 248 -1842 248 -1842 0 feedthrough
rlabel pdiffusion 255 -1842 255 -1842 0 feedthrough
rlabel pdiffusion 262 -1842 262 -1842 0 feedthrough
rlabel pdiffusion 269 -1842 269 -1842 0 feedthrough
rlabel pdiffusion 276 -1842 276 -1842 0 feedthrough
rlabel pdiffusion 283 -1842 283 -1842 0 feedthrough
rlabel pdiffusion 290 -1842 290 -1842 0 feedthrough
rlabel pdiffusion 297 -1842 297 -1842 0 cellNo=484
rlabel pdiffusion 304 -1842 304 -1842 0 feedthrough
rlabel pdiffusion 311 -1842 311 -1842 0 feedthrough
rlabel pdiffusion 318 -1842 318 -1842 0 feedthrough
rlabel pdiffusion 325 -1842 325 -1842 0 feedthrough
rlabel pdiffusion 332 -1842 332 -1842 0 feedthrough
rlabel pdiffusion 339 -1842 339 -1842 0 feedthrough
rlabel pdiffusion 346 -1842 346 -1842 0 feedthrough
rlabel pdiffusion 353 -1842 353 -1842 0 cellNo=589
rlabel pdiffusion 360 -1842 360 -1842 0 feedthrough
rlabel pdiffusion 367 -1842 367 -1842 0 cellNo=454
rlabel pdiffusion 374 -1842 374 -1842 0 feedthrough
rlabel pdiffusion 381 -1842 381 -1842 0 feedthrough
rlabel pdiffusion 388 -1842 388 -1842 0 cellNo=460
rlabel pdiffusion 395 -1842 395 -1842 0 feedthrough
rlabel pdiffusion 402 -1842 402 -1842 0 feedthrough
rlabel pdiffusion 409 -1842 409 -1842 0 feedthrough
rlabel pdiffusion 416 -1842 416 -1842 0 feedthrough
rlabel pdiffusion 423 -1842 423 -1842 0 feedthrough
rlabel pdiffusion 430 -1842 430 -1842 0 feedthrough
rlabel pdiffusion 437 -1842 437 -1842 0 feedthrough
rlabel pdiffusion 444 -1842 444 -1842 0 feedthrough
rlabel pdiffusion 451 -1842 451 -1842 0 feedthrough
rlabel pdiffusion 458 -1842 458 -1842 0 feedthrough
rlabel pdiffusion 465 -1842 465 -1842 0 cellNo=158
rlabel pdiffusion 472 -1842 472 -1842 0 feedthrough
rlabel pdiffusion 479 -1842 479 -1842 0 cellNo=46
rlabel pdiffusion 486 -1842 486 -1842 0 feedthrough
rlabel pdiffusion 493 -1842 493 -1842 0 feedthrough
rlabel pdiffusion 500 -1842 500 -1842 0 feedthrough
rlabel pdiffusion 507 -1842 507 -1842 0 feedthrough
rlabel pdiffusion 514 -1842 514 -1842 0 cellNo=326
rlabel pdiffusion 521 -1842 521 -1842 0 feedthrough
rlabel pdiffusion 528 -1842 528 -1842 0 feedthrough
rlabel pdiffusion 535 -1842 535 -1842 0 feedthrough
rlabel pdiffusion 542 -1842 542 -1842 0 feedthrough
rlabel pdiffusion 549 -1842 549 -1842 0 feedthrough
rlabel pdiffusion 556 -1842 556 -1842 0 feedthrough
rlabel pdiffusion 563 -1842 563 -1842 0 feedthrough
rlabel pdiffusion 570 -1842 570 -1842 0 feedthrough
rlabel pdiffusion 577 -1842 577 -1842 0 feedthrough
rlabel pdiffusion 584 -1842 584 -1842 0 cellNo=89
rlabel pdiffusion 591 -1842 591 -1842 0 feedthrough
rlabel pdiffusion 598 -1842 598 -1842 0 feedthrough
rlabel pdiffusion 605 -1842 605 -1842 0 cellNo=551
rlabel pdiffusion 612 -1842 612 -1842 0 cellNo=162
rlabel pdiffusion 619 -1842 619 -1842 0 feedthrough
rlabel pdiffusion 626 -1842 626 -1842 0 cellNo=370
rlabel pdiffusion 633 -1842 633 -1842 0 feedthrough
rlabel pdiffusion 640 -1842 640 -1842 0 cellNo=550
rlabel pdiffusion 647 -1842 647 -1842 0 feedthrough
rlabel pdiffusion 654 -1842 654 -1842 0 cellNo=330
rlabel pdiffusion 661 -1842 661 -1842 0 feedthrough
rlabel pdiffusion 668 -1842 668 -1842 0 feedthrough
rlabel pdiffusion 675 -1842 675 -1842 0 feedthrough
rlabel pdiffusion 682 -1842 682 -1842 0 feedthrough
rlabel pdiffusion 689 -1842 689 -1842 0 feedthrough
rlabel pdiffusion 696 -1842 696 -1842 0 feedthrough
rlabel pdiffusion 703 -1842 703 -1842 0 feedthrough
rlabel pdiffusion 710 -1842 710 -1842 0 cellNo=348
rlabel pdiffusion 717 -1842 717 -1842 0 cellNo=443
rlabel pdiffusion 724 -1842 724 -1842 0 feedthrough
rlabel pdiffusion 731 -1842 731 -1842 0 cellNo=42
rlabel pdiffusion 738 -1842 738 -1842 0 feedthrough
rlabel pdiffusion 745 -1842 745 -1842 0 feedthrough
rlabel pdiffusion 752 -1842 752 -1842 0 cellNo=72
rlabel pdiffusion 759 -1842 759 -1842 0 cellNo=180
rlabel pdiffusion 766 -1842 766 -1842 0 feedthrough
rlabel pdiffusion 773 -1842 773 -1842 0 feedthrough
rlabel pdiffusion 780 -1842 780 -1842 0 feedthrough
rlabel pdiffusion 787 -1842 787 -1842 0 feedthrough
rlabel pdiffusion 794 -1842 794 -1842 0 feedthrough
rlabel pdiffusion 801 -1842 801 -1842 0 feedthrough
rlabel pdiffusion 808 -1842 808 -1842 0 feedthrough
rlabel pdiffusion 815 -1842 815 -1842 0 feedthrough
rlabel pdiffusion 822 -1842 822 -1842 0 feedthrough
rlabel pdiffusion 829 -1842 829 -1842 0 feedthrough
rlabel pdiffusion 836 -1842 836 -1842 0 feedthrough
rlabel pdiffusion 843 -1842 843 -1842 0 feedthrough
rlabel pdiffusion 850 -1842 850 -1842 0 feedthrough
rlabel pdiffusion 857 -1842 857 -1842 0 feedthrough
rlabel pdiffusion 864 -1842 864 -1842 0 feedthrough
rlabel pdiffusion 871 -1842 871 -1842 0 feedthrough
rlabel pdiffusion 878 -1842 878 -1842 0 feedthrough
rlabel pdiffusion 885 -1842 885 -1842 0 feedthrough
rlabel pdiffusion 892 -1842 892 -1842 0 feedthrough
rlabel pdiffusion 899 -1842 899 -1842 0 feedthrough
rlabel pdiffusion 906 -1842 906 -1842 0 feedthrough
rlabel pdiffusion 913 -1842 913 -1842 0 feedthrough
rlabel pdiffusion 920 -1842 920 -1842 0 feedthrough
rlabel pdiffusion 927 -1842 927 -1842 0 feedthrough
rlabel pdiffusion 934 -1842 934 -1842 0 feedthrough
rlabel pdiffusion 941 -1842 941 -1842 0 feedthrough
rlabel pdiffusion 948 -1842 948 -1842 0 feedthrough
rlabel pdiffusion 955 -1842 955 -1842 0 feedthrough
rlabel pdiffusion 962 -1842 962 -1842 0 feedthrough
rlabel pdiffusion 969 -1842 969 -1842 0 feedthrough
rlabel pdiffusion 976 -1842 976 -1842 0 feedthrough
rlabel pdiffusion 983 -1842 983 -1842 0 feedthrough
rlabel pdiffusion 990 -1842 990 -1842 0 feedthrough
rlabel pdiffusion 997 -1842 997 -1842 0 feedthrough
rlabel pdiffusion 1004 -1842 1004 -1842 0 feedthrough
rlabel pdiffusion 1011 -1842 1011 -1842 0 feedthrough
rlabel pdiffusion 1018 -1842 1018 -1842 0 feedthrough
rlabel pdiffusion 1025 -1842 1025 -1842 0 feedthrough
rlabel pdiffusion 1032 -1842 1032 -1842 0 feedthrough
rlabel pdiffusion 1039 -1842 1039 -1842 0 feedthrough
rlabel pdiffusion 1046 -1842 1046 -1842 0 feedthrough
rlabel pdiffusion 1053 -1842 1053 -1842 0 feedthrough
rlabel pdiffusion 1060 -1842 1060 -1842 0 feedthrough
rlabel pdiffusion 1067 -1842 1067 -1842 0 feedthrough
rlabel pdiffusion 1074 -1842 1074 -1842 0 feedthrough
rlabel pdiffusion 1081 -1842 1081 -1842 0 feedthrough
rlabel pdiffusion 1088 -1842 1088 -1842 0 feedthrough
rlabel pdiffusion 1095 -1842 1095 -1842 0 feedthrough
rlabel pdiffusion 1102 -1842 1102 -1842 0 feedthrough
rlabel pdiffusion 1109 -1842 1109 -1842 0 feedthrough
rlabel pdiffusion 1116 -1842 1116 -1842 0 feedthrough
rlabel pdiffusion 1123 -1842 1123 -1842 0 feedthrough
rlabel pdiffusion 1130 -1842 1130 -1842 0 feedthrough
rlabel pdiffusion 1137 -1842 1137 -1842 0 feedthrough
rlabel pdiffusion 1144 -1842 1144 -1842 0 feedthrough
rlabel pdiffusion 1151 -1842 1151 -1842 0 feedthrough
rlabel pdiffusion 1158 -1842 1158 -1842 0 feedthrough
rlabel pdiffusion 1165 -1842 1165 -1842 0 feedthrough
rlabel pdiffusion 1172 -1842 1172 -1842 0 feedthrough
rlabel pdiffusion 1179 -1842 1179 -1842 0 feedthrough
rlabel pdiffusion 1186 -1842 1186 -1842 0 feedthrough
rlabel pdiffusion 1193 -1842 1193 -1842 0 feedthrough
rlabel pdiffusion 1200 -1842 1200 -1842 0 feedthrough
rlabel pdiffusion 1207 -1842 1207 -1842 0 feedthrough
rlabel pdiffusion 1214 -1842 1214 -1842 0 feedthrough
rlabel pdiffusion 1221 -1842 1221 -1842 0 feedthrough
rlabel pdiffusion 1228 -1842 1228 -1842 0 feedthrough
rlabel pdiffusion 1235 -1842 1235 -1842 0 feedthrough
rlabel pdiffusion 1242 -1842 1242 -1842 0 feedthrough
rlabel pdiffusion 1249 -1842 1249 -1842 0 feedthrough
rlabel pdiffusion 1256 -1842 1256 -1842 0 feedthrough
rlabel pdiffusion 1263 -1842 1263 -1842 0 feedthrough
rlabel pdiffusion 1270 -1842 1270 -1842 0 feedthrough
rlabel pdiffusion 1277 -1842 1277 -1842 0 feedthrough
rlabel pdiffusion 1284 -1842 1284 -1842 0 cellNo=568
rlabel pdiffusion 10 -1965 10 -1965 0 feedthrough
rlabel pdiffusion 17 -1965 17 -1965 0 feedthrough
rlabel pdiffusion 24 -1965 24 -1965 0 feedthrough
rlabel pdiffusion 31 -1965 31 -1965 0 feedthrough
rlabel pdiffusion 38 -1965 38 -1965 0 feedthrough
rlabel pdiffusion 45 -1965 45 -1965 0 feedthrough
rlabel pdiffusion 52 -1965 52 -1965 0 cellNo=546
rlabel pdiffusion 59 -1965 59 -1965 0 feedthrough
rlabel pdiffusion 66 -1965 66 -1965 0 cellNo=558
rlabel pdiffusion 73 -1965 73 -1965 0 feedthrough
rlabel pdiffusion 80 -1965 80 -1965 0 feedthrough
rlabel pdiffusion 87 -1965 87 -1965 0 cellNo=36
rlabel pdiffusion 94 -1965 94 -1965 0 cellNo=204
rlabel pdiffusion 101 -1965 101 -1965 0 cellNo=189
rlabel pdiffusion 108 -1965 108 -1965 0 feedthrough
rlabel pdiffusion 115 -1965 115 -1965 0 feedthrough
rlabel pdiffusion 122 -1965 122 -1965 0 feedthrough
rlabel pdiffusion 129 -1965 129 -1965 0 feedthrough
rlabel pdiffusion 136 -1965 136 -1965 0 cellNo=523
rlabel pdiffusion 143 -1965 143 -1965 0 feedthrough
rlabel pdiffusion 150 -1965 150 -1965 0 feedthrough
rlabel pdiffusion 157 -1965 157 -1965 0 feedthrough
rlabel pdiffusion 164 -1965 164 -1965 0 feedthrough
rlabel pdiffusion 171 -1965 171 -1965 0 cellNo=211
rlabel pdiffusion 178 -1965 178 -1965 0 feedthrough
rlabel pdiffusion 185 -1965 185 -1965 0 feedthrough
rlabel pdiffusion 192 -1965 192 -1965 0 feedthrough
rlabel pdiffusion 199 -1965 199 -1965 0 feedthrough
rlabel pdiffusion 206 -1965 206 -1965 0 feedthrough
rlabel pdiffusion 213 -1965 213 -1965 0 feedthrough
rlabel pdiffusion 220 -1965 220 -1965 0 feedthrough
rlabel pdiffusion 227 -1965 227 -1965 0 feedthrough
rlabel pdiffusion 234 -1965 234 -1965 0 feedthrough
rlabel pdiffusion 241 -1965 241 -1965 0 feedthrough
rlabel pdiffusion 248 -1965 248 -1965 0 feedthrough
rlabel pdiffusion 255 -1965 255 -1965 0 feedthrough
rlabel pdiffusion 262 -1965 262 -1965 0 cellNo=285
rlabel pdiffusion 269 -1965 269 -1965 0 feedthrough
rlabel pdiffusion 276 -1965 276 -1965 0 feedthrough
rlabel pdiffusion 283 -1965 283 -1965 0 cellNo=594
rlabel pdiffusion 290 -1965 290 -1965 0 feedthrough
rlabel pdiffusion 297 -1965 297 -1965 0 feedthrough
rlabel pdiffusion 304 -1965 304 -1965 0 feedthrough
rlabel pdiffusion 311 -1965 311 -1965 0 feedthrough
rlabel pdiffusion 318 -1965 318 -1965 0 cellNo=387
rlabel pdiffusion 325 -1965 325 -1965 0 feedthrough
rlabel pdiffusion 332 -1965 332 -1965 0 feedthrough
rlabel pdiffusion 339 -1965 339 -1965 0 feedthrough
rlabel pdiffusion 346 -1965 346 -1965 0 feedthrough
rlabel pdiffusion 353 -1965 353 -1965 0 feedthrough
rlabel pdiffusion 360 -1965 360 -1965 0 feedthrough
rlabel pdiffusion 367 -1965 367 -1965 0 cellNo=467
rlabel pdiffusion 374 -1965 374 -1965 0 feedthrough
rlabel pdiffusion 381 -1965 381 -1965 0 feedthrough
rlabel pdiffusion 388 -1965 388 -1965 0 feedthrough
rlabel pdiffusion 395 -1965 395 -1965 0 feedthrough
rlabel pdiffusion 402 -1965 402 -1965 0 feedthrough
rlabel pdiffusion 409 -1965 409 -1965 0 feedthrough
rlabel pdiffusion 416 -1965 416 -1965 0 feedthrough
rlabel pdiffusion 423 -1965 423 -1965 0 feedthrough
rlabel pdiffusion 430 -1965 430 -1965 0 cellNo=337
rlabel pdiffusion 437 -1965 437 -1965 0 feedthrough
rlabel pdiffusion 444 -1965 444 -1965 0 feedthrough
rlabel pdiffusion 451 -1965 451 -1965 0 feedthrough
rlabel pdiffusion 458 -1965 458 -1965 0 cellNo=257
rlabel pdiffusion 465 -1965 465 -1965 0 feedthrough
rlabel pdiffusion 472 -1965 472 -1965 0 feedthrough
rlabel pdiffusion 479 -1965 479 -1965 0 feedthrough
rlabel pdiffusion 486 -1965 486 -1965 0 feedthrough
rlabel pdiffusion 493 -1965 493 -1965 0 cellNo=230
rlabel pdiffusion 500 -1965 500 -1965 0 feedthrough
rlabel pdiffusion 507 -1965 507 -1965 0 feedthrough
rlabel pdiffusion 514 -1965 514 -1965 0 feedthrough
rlabel pdiffusion 521 -1965 521 -1965 0 cellNo=398
rlabel pdiffusion 528 -1965 528 -1965 0 feedthrough
rlabel pdiffusion 535 -1965 535 -1965 0 feedthrough
rlabel pdiffusion 542 -1965 542 -1965 0 feedthrough
rlabel pdiffusion 549 -1965 549 -1965 0 feedthrough
rlabel pdiffusion 556 -1965 556 -1965 0 cellNo=441
rlabel pdiffusion 563 -1965 563 -1965 0 feedthrough
rlabel pdiffusion 570 -1965 570 -1965 0 cellNo=231
rlabel pdiffusion 577 -1965 577 -1965 0 feedthrough
rlabel pdiffusion 584 -1965 584 -1965 0 feedthrough
rlabel pdiffusion 591 -1965 591 -1965 0 feedthrough
rlabel pdiffusion 598 -1965 598 -1965 0 feedthrough
rlabel pdiffusion 605 -1965 605 -1965 0 cellNo=552
rlabel pdiffusion 612 -1965 612 -1965 0 feedthrough
rlabel pdiffusion 619 -1965 619 -1965 0 feedthrough
rlabel pdiffusion 626 -1965 626 -1965 0 feedthrough
rlabel pdiffusion 633 -1965 633 -1965 0 feedthrough
rlabel pdiffusion 640 -1965 640 -1965 0 feedthrough
rlabel pdiffusion 647 -1965 647 -1965 0 feedthrough
rlabel pdiffusion 654 -1965 654 -1965 0 feedthrough
rlabel pdiffusion 661 -1965 661 -1965 0 feedthrough
rlabel pdiffusion 668 -1965 668 -1965 0 feedthrough
rlabel pdiffusion 675 -1965 675 -1965 0 cellNo=399
rlabel pdiffusion 682 -1965 682 -1965 0 feedthrough
rlabel pdiffusion 689 -1965 689 -1965 0 feedthrough
rlabel pdiffusion 696 -1965 696 -1965 0 feedthrough
rlabel pdiffusion 703 -1965 703 -1965 0 cellNo=503
rlabel pdiffusion 710 -1965 710 -1965 0 feedthrough
rlabel pdiffusion 717 -1965 717 -1965 0 feedthrough
rlabel pdiffusion 724 -1965 724 -1965 0 feedthrough
rlabel pdiffusion 731 -1965 731 -1965 0 feedthrough
rlabel pdiffusion 738 -1965 738 -1965 0 feedthrough
rlabel pdiffusion 745 -1965 745 -1965 0 feedthrough
rlabel pdiffusion 752 -1965 752 -1965 0 feedthrough
rlabel pdiffusion 759 -1965 759 -1965 0 cellNo=281
rlabel pdiffusion 766 -1965 766 -1965 0 feedthrough
rlabel pdiffusion 773 -1965 773 -1965 0 feedthrough
rlabel pdiffusion 780 -1965 780 -1965 0 feedthrough
rlabel pdiffusion 787 -1965 787 -1965 0 feedthrough
rlabel pdiffusion 794 -1965 794 -1965 0 feedthrough
rlabel pdiffusion 801 -1965 801 -1965 0 feedthrough
rlabel pdiffusion 808 -1965 808 -1965 0 feedthrough
rlabel pdiffusion 815 -1965 815 -1965 0 feedthrough
rlabel pdiffusion 822 -1965 822 -1965 0 feedthrough
rlabel pdiffusion 829 -1965 829 -1965 0 feedthrough
rlabel pdiffusion 836 -1965 836 -1965 0 cellNo=488
rlabel pdiffusion 843 -1965 843 -1965 0 feedthrough
rlabel pdiffusion 850 -1965 850 -1965 0 feedthrough
rlabel pdiffusion 857 -1965 857 -1965 0 feedthrough
rlabel pdiffusion 864 -1965 864 -1965 0 feedthrough
rlabel pdiffusion 871 -1965 871 -1965 0 feedthrough
rlabel pdiffusion 878 -1965 878 -1965 0 feedthrough
rlabel pdiffusion 885 -1965 885 -1965 0 feedthrough
rlabel pdiffusion 892 -1965 892 -1965 0 feedthrough
rlabel pdiffusion 899 -1965 899 -1965 0 feedthrough
rlabel pdiffusion 906 -1965 906 -1965 0 feedthrough
rlabel pdiffusion 913 -1965 913 -1965 0 feedthrough
rlabel pdiffusion 920 -1965 920 -1965 0 cellNo=524
rlabel pdiffusion 927 -1965 927 -1965 0 feedthrough
rlabel pdiffusion 934 -1965 934 -1965 0 feedthrough
rlabel pdiffusion 941 -1965 941 -1965 0 feedthrough
rlabel pdiffusion 948 -1965 948 -1965 0 feedthrough
rlabel pdiffusion 955 -1965 955 -1965 0 feedthrough
rlabel pdiffusion 962 -1965 962 -1965 0 cellNo=340
rlabel pdiffusion 969 -1965 969 -1965 0 feedthrough
rlabel pdiffusion 976 -1965 976 -1965 0 feedthrough
rlabel pdiffusion 983 -1965 983 -1965 0 feedthrough
rlabel pdiffusion 990 -1965 990 -1965 0 feedthrough
rlabel pdiffusion 997 -1965 997 -1965 0 feedthrough
rlabel pdiffusion 1004 -1965 1004 -1965 0 feedthrough
rlabel pdiffusion 1011 -1965 1011 -1965 0 feedthrough
rlabel pdiffusion 1018 -1965 1018 -1965 0 feedthrough
rlabel pdiffusion 1025 -1965 1025 -1965 0 feedthrough
rlabel pdiffusion 1032 -1965 1032 -1965 0 feedthrough
rlabel pdiffusion 1039 -1965 1039 -1965 0 feedthrough
rlabel pdiffusion 1046 -1965 1046 -1965 0 feedthrough
rlabel pdiffusion 1053 -1965 1053 -1965 0 feedthrough
rlabel pdiffusion 1060 -1965 1060 -1965 0 feedthrough
rlabel pdiffusion 1067 -1965 1067 -1965 0 feedthrough
rlabel pdiffusion 1074 -1965 1074 -1965 0 feedthrough
rlabel pdiffusion 1081 -1965 1081 -1965 0 feedthrough
rlabel pdiffusion 1088 -1965 1088 -1965 0 feedthrough
rlabel pdiffusion 1095 -1965 1095 -1965 0 feedthrough
rlabel pdiffusion 1102 -1965 1102 -1965 0 feedthrough
rlabel pdiffusion 1109 -1965 1109 -1965 0 feedthrough
rlabel pdiffusion 1116 -1965 1116 -1965 0 feedthrough
rlabel pdiffusion 1123 -1965 1123 -1965 0 feedthrough
rlabel pdiffusion 1130 -1965 1130 -1965 0 feedthrough
rlabel pdiffusion 1137 -1965 1137 -1965 0 feedthrough
rlabel pdiffusion 1144 -1965 1144 -1965 0 feedthrough
rlabel pdiffusion 1151 -1965 1151 -1965 0 feedthrough
rlabel pdiffusion 1158 -1965 1158 -1965 0 feedthrough
rlabel pdiffusion 1165 -1965 1165 -1965 0 feedthrough
rlabel pdiffusion 1172 -1965 1172 -1965 0 feedthrough
rlabel pdiffusion 1179 -1965 1179 -1965 0 feedthrough
rlabel pdiffusion 1186 -1965 1186 -1965 0 feedthrough
rlabel pdiffusion 1193 -1965 1193 -1965 0 feedthrough
rlabel pdiffusion 1200 -1965 1200 -1965 0 feedthrough
rlabel pdiffusion 1207 -1965 1207 -1965 0 feedthrough
rlabel pdiffusion 1214 -1965 1214 -1965 0 feedthrough
rlabel pdiffusion 1221 -1965 1221 -1965 0 cellNo=167
rlabel pdiffusion 1228 -1965 1228 -1965 0 feedthrough
rlabel pdiffusion 1235 -1965 1235 -1965 0 feedthrough
rlabel pdiffusion 3 -2068 3 -2068 0 feedthrough
rlabel pdiffusion 10 -2068 10 -2068 0 feedthrough
rlabel pdiffusion 17 -2068 17 -2068 0 feedthrough
rlabel pdiffusion 24 -2068 24 -2068 0 feedthrough
rlabel pdiffusion 31 -2068 31 -2068 0 feedthrough
rlabel pdiffusion 38 -2068 38 -2068 0 feedthrough
rlabel pdiffusion 45 -2068 45 -2068 0 feedthrough
rlabel pdiffusion 52 -2068 52 -2068 0 feedthrough
rlabel pdiffusion 59 -2068 59 -2068 0 feedthrough
rlabel pdiffusion 66 -2068 66 -2068 0 feedthrough
rlabel pdiffusion 73 -2068 73 -2068 0 feedthrough
rlabel pdiffusion 80 -2068 80 -2068 0 feedthrough
rlabel pdiffusion 87 -2068 87 -2068 0 cellNo=197
rlabel pdiffusion 94 -2068 94 -2068 0 cellNo=268
rlabel pdiffusion 101 -2068 101 -2068 0 feedthrough
rlabel pdiffusion 108 -2068 108 -2068 0 cellNo=142
rlabel pdiffusion 115 -2068 115 -2068 0 cellNo=44
rlabel pdiffusion 122 -2068 122 -2068 0 feedthrough
rlabel pdiffusion 129 -2068 129 -2068 0 feedthrough
rlabel pdiffusion 136 -2068 136 -2068 0 feedthrough
rlabel pdiffusion 143 -2068 143 -2068 0 feedthrough
rlabel pdiffusion 150 -2068 150 -2068 0 cellNo=410
rlabel pdiffusion 157 -2068 157 -2068 0 feedthrough
rlabel pdiffusion 164 -2068 164 -2068 0 cellNo=520
rlabel pdiffusion 171 -2068 171 -2068 0 feedthrough
rlabel pdiffusion 178 -2068 178 -2068 0 feedthrough
rlabel pdiffusion 185 -2068 185 -2068 0 feedthrough
rlabel pdiffusion 192 -2068 192 -2068 0 feedthrough
rlabel pdiffusion 199 -2068 199 -2068 0 feedthrough
rlabel pdiffusion 206 -2068 206 -2068 0 feedthrough
rlabel pdiffusion 213 -2068 213 -2068 0 feedthrough
rlabel pdiffusion 220 -2068 220 -2068 0 feedthrough
rlabel pdiffusion 227 -2068 227 -2068 0 feedthrough
rlabel pdiffusion 234 -2068 234 -2068 0 feedthrough
rlabel pdiffusion 241 -2068 241 -2068 0 cellNo=239
rlabel pdiffusion 248 -2068 248 -2068 0 feedthrough
rlabel pdiffusion 255 -2068 255 -2068 0 feedthrough
rlabel pdiffusion 262 -2068 262 -2068 0 feedthrough
rlabel pdiffusion 269 -2068 269 -2068 0 feedthrough
rlabel pdiffusion 276 -2068 276 -2068 0 cellNo=361
rlabel pdiffusion 283 -2068 283 -2068 0 feedthrough
rlabel pdiffusion 290 -2068 290 -2068 0 feedthrough
rlabel pdiffusion 297 -2068 297 -2068 0 feedthrough
rlabel pdiffusion 304 -2068 304 -2068 0 feedthrough
rlabel pdiffusion 311 -2068 311 -2068 0 feedthrough
rlabel pdiffusion 318 -2068 318 -2068 0 feedthrough
rlabel pdiffusion 325 -2068 325 -2068 0 cellNo=302
rlabel pdiffusion 332 -2068 332 -2068 0 cellNo=482
rlabel pdiffusion 339 -2068 339 -2068 0 feedthrough
rlabel pdiffusion 346 -2068 346 -2068 0 feedthrough
rlabel pdiffusion 353 -2068 353 -2068 0 feedthrough
rlabel pdiffusion 360 -2068 360 -2068 0 feedthrough
rlabel pdiffusion 367 -2068 367 -2068 0 feedthrough
rlabel pdiffusion 374 -2068 374 -2068 0 feedthrough
rlabel pdiffusion 381 -2068 381 -2068 0 feedthrough
rlabel pdiffusion 388 -2068 388 -2068 0 feedthrough
rlabel pdiffusion 395 -2068 395 -2068 0 feedthrough
rlabel pdiffusion 402 -2068 402 -2068 0 feedthrough
rlabel pdiffusion 409 -2068 409 -2068 0 cellNo=347
rlabel pdiffusion 416 -2068 416 -2068 0 feedthrough
rlabel pdiffusion 423 -2068 423 -2068 0 feedthrough
rlabel pdiffusion 430 -2068 430 -2068 0 feedthrough
rlabel pdiffusion 437 -2068 437 -2068 0 feedthrough
rlabel pdiffusion 444 -2068 444 -2068 0 feedthrough
rlabel pdiffusion 451 -2068 451 -2068 0 feedthrough
rlabel pdiffusion 458 -2068 458 -2068 0 feedthrough
rlabel pdiffusion 465 -2068 465 -2068 0 feedthrough
rlabel pdiffusion 472 -2068 472 -2068 0 feedthrough
rlabel pdiffusion 479 -2068 479 -2068 0 cellNo=438
rlabel pdiffusion 486 -2068 486 -2068 0 cellNo=222
rlabel pdiffusion 493 -2068 493 -2068 0 feedthrough
rlabel pdiffusion 500 -2068 500 -2068 0 cellNo=219
rlabel pdiffusion 507 -2068 507 -2068 0 feedthrough
rlabel pdiffusion 514 -2068 514 -2068 0 feedthrough
rlabel pdiffusion 521 -2068 521 -2068 0 feedthrough
rlabel pdiffusion 528 -2068 528 -2068 0 feedthrough
rlabel pdiffusion 535 -2068 535 -2068 0 feedthrough
rlabel pdiffusion 542 -2068 542 -2068 0 feedthrough
rlabel pdiffusion 549 -2068 549 -2068 0 feedthrough
rlabel pdiffusion 556 -2068 556 -2068 0 feedthrough
rlabel pdiffusion 563 -2068 563 -2068 0 feedthrough
rlabel pdiffusion 570 -2068 570 -2068 0 feedthrough
rlabel pdiffusion 577 -2068 577 -2068 0 cellNo=21
rlabel pdiffusion 584 -2068 584 -2068 0 cellNo=431
rlabel pdiffusion 591 -2068 591 -2068 0 feedthrough
rlabel pdiffusion 598 -2068 598 -2068 0 feedthrough
rlabel pdiffusion 605 -2068 605 -2068 0 feedthrough
rlabel pdiffusion 612 -2068 612 -2068 0 feedthrough
rlabel pdiffusion 619 -2068 619 -2068 0 cellNo=391
rlabel pdiffusion 626 -2068 626 -2068 0 feedthrough
rlabel pdiffusion 633 -2068 633 -2068 0 feedthrough
rlabel pdiffusion 640 -2068 640 -2068 0 feedthrough
rlabel pdiffusion 647 -2068 647 -2068 0 feedthrough
rlabel pdiffusion 654 -2068 654 -2068 0 cellNo=174
rlabel pdiffusion 661 -2068 661 -2068 0 cellNo=590
rlabel pdiffusion 668 -2068 668 -2068 0 feedthrough
rlabel pdiffusion 675 -2068 675 -2068 0 feedthrough
rlabel pdiffusion 682 -2068 682 -2068 0 feedthrough
rlabel pdiffusion 689 -2068 689 -2068 0 feedthrough
rlabel pdiffusion 696 -2068 696 -2068 0 cellNo=429
rlabel pdiffusion 703 -2068 703 -2068 0 feedthrough
rlabel pdiffusion 710 -2068 710 -2068 0 feedthrough
rlabel pdiffusion 717 -2068 717 -2068 0 feedthrough
rlabel pdiffusion 724 -2068 724 -2068 0 feedthrough
rlabel pdiffusion 731 -2068 731 -2068 0 feedthrough
rlabel pdiffusion 738 -2068 738 -2068 0 feedthrough
rlabel pdiffusion 745 -2068 745 -2068 0 feedthrough
rlabel pdiffusion 752 -2068 752 -2068 0 feedthrough
rlabel pdiffusion 759 -2068 759 -2068 0 feedthrough
rlabel pdiffusion 766 -2068 766 -2068 0 feedthrough
rlabel pdiffusion 773 -2068 773 -2068 0 feedthrough
rlabel pdiffusion 780 -2068 780 -2068 0 feedthrough
rlabel pdiffusion 787 -2068 787 -2068 0 feedthrough
rlabel pdiffusion 794 -2068 794 -2068 0 feedthrough
rlabel pdiffusion 801 -2068 801 -2068 0 feedthrough
rlabel pdiffusion 808 -2068 808 -2068 0 feedthrough
rlabel pdiffusion 815 -2068 815 -2068 0 cellNo=251
rlabel pdiffusion 822 -2068 822 -2068 0 feedthrough
rlabel pdiffusion 829 -2068 829 -2068 0 feedthrough
rlabel pdiffusion 836 -2068 836 -2068 0 feedthrough
rlabel pdiffusion 843 -2068 843 -2068 0 feedthrough
rlabel pdiffusion 850 -2068 850 -2068 0 feedthrough
rlabel pdiffusion 857 -2068 857 -2068 0 feedthrough
rlabel pdiffusion 864 -2068 864 -2068 0 cellNo=517
rlabel pdiffusion 871 -2068 871 -2068 0 feedthrough
rlabel pdiffusion 878 -2068 878 -2068 0 feedthrough
rlabel pdiffusion 885 -2068 885 -2068 0 feedthrough
rlabel pdiffusion 892 -2068 892 -2068 0 feedthrough
rlabel pdiffusion 899 -2068 899 -2068 0 feedthrough
rlabel pdiffusion 906 -2068 906 -2068 0 feedthrough
rlabel pdiffusion 913 -2068 913 -2068 0 feedthrough
rlabel pdiffusion 920 -2068 920 -2068 0 feedthrough
rlabel pdiffusion 927 -2068 927 -2068 0 feedthrough
rlabel pdiffusion 934 -2068 934 -2068 0 feedthrough
rlabel pdiffusion 941 -2068 941 -2068 0 feedthrough
rlabel pdiffusion 948 -2068 948 -2068 0 feedthrough
rlabel pdiffusion 955 -2068 955 -2068 0 feedthrough
rlabel pdiffusion 962 -2068 962 -2068 0 feedthrough
rlabel pdiffusion 969 -2068 969 -2068 0 feedthrough
rlabel pdiffusion 976 -2068 976 -2068 0 feedthrough
rlabel pdiffusion 983 -2068 983 -2068 0 feedthrough
rlabel pdiffusion 990 -2068 990 -2068 0 feedthrough
rlabel pdiffusion 997 -2068 997 -2068 0 feedthrough
rlabel pdiffusion 1004 -2068 1004 -2068 0 feedthrough
rlabel pdiffusion 1011 -2068 1011 -2068 0 feedthrough
rlabel pdiffusion 1018 -2068 1018 -2068 0 feedthrough
rlabel pdiffusion 1025 -2068 1025 -2068 0 cellNo=519
rlabel pdiffusion 1032 -2068 1032 -2068 0 feedthrough
rlabel pdiffusion 1039 -2068 1039 -2068 0 feedthrough
rlabel pdiffusion 1046 -2068 1046 -2068 0 feedthrough
rlabel pdiffusion 1053 -2068 1053 -2068 0 feedthrough
rlabel pdiffusion 1060 -2068 1060 -2068 0 feedthrough
rlabel pdiffusion 1067 -2068 1067 -2068 0 feedthrough
rlabel pdiffusion 1074 -2068 1074 -2068 0 feedthrough
rlabel pdiffusion 1081 -2068 1081 -2068 0 feedthrough
rlabel pdiffusion 1088 -2068 1088 -2068 0 feedthrough
rlabel pdiffusion 1095 -2068 1095 -2068 0 feedthrough
rlabel pdiffusion 1102 -2068 1102 -2068 0 feedthrough
rlabel pdiffusion 1109 -2068 1109 -2068 0 feedthrough
rlabel pdiffusion 1116 -2068 1116 -2068 0 feedthrough
rlabel pdiffusion 1123 -2068 1123 -2068 0 feedthrough
rlabel pdiffusion 1130 -2068 1130 -2068 0 feedthrough
rlabel pdiffusion 1137 -2068 1137 -2068 0 cellNo=288
rlabel pdiffusion 1144 -2068 1144 -2068 0 feedthrough
rlabel pdiffusion 1151 -2068 1151 -2068 0 feedthrough
rlabel pdiffusion 1158 -2068 1158 -2068 0 feedthrough
rlabel pdiffusion 1186 -2068 1186 -2068 0 feedthrough
rlabel pdiffusion 24 -2153 24 -2153 0 feedthrough
rlabel pdiffusion 31 -2153 31 -2153 0 feedthrough
rlabel pdiffusion 38 -2153 38 -2153 0 feedthrough
rlabel pdiffusion 45 -2153 45 -2153 0 feedthrough
rlabel pdiffusion 52 -2153 52 -2153 0 feedthrough
rlabel pdiffusion 59 -2153 59 -2153 0 feedthrough
rlabel pdiffusion 66 -2153 66 -2153 0 feedthrough
rlabel pdiffusion 73 -2153 73 -2153 0 feedthrough
rlabel pdiffusion 80 -2153 80 -2153 0 feedthrough
rlabel pdiffusion 87 -2153 87 -2153 0 feedthrough
rlabel pdiffusion 94 -2153 94 -2153 0 cellNo=228
rlabel pdiffusion 101 -2153 101 -2153 0 cellNo=434
rlabel pdiffusion 108 -2153 108 -2153 0 feedthrough
rlabel pdiffusion 115 -2153 115 -2153 0 cellNo=506
rlabel pdiffusion 122 -2153 122 -2153 0 feedthrough
rlabel pdiffusion 129 -2153 129 -2153 0 feedthrough
rlabel pdiffusion 136 -2153 136 -2153 0 cellNo=459
rlabel pdiffusion 143 -2153 143 -2153 0 feedthrough
rlabel pdiffusion 150 -2153 150 -2153 0 feedthrough
rlabel pdiffusion 157 -2153 157 -2153 0 feedthrough
rlabel pdiffusion 164 -2153 164 -2153 0 feedthrough
rlabel pdiffusion 171 -2153 171 -2153 0 cellNo=196
rlabel pdiffusion 178 -2153 178 -2153 0 feedthrough
rlabel pdiffusion 185 -2153 185 -2153 0 feedthrough
rlabel pdiffusion 192 -2153 192 -2153 0 feedthrough
rlabel pdiffusion 199 -2153 199 -2153 0 feedthrough
rlabel pdiffusion 206 -2153 206 -2153 0 feedthrough
rlabel pdiffusion 213 -2153 213 -2153 0 feedthrough
rlabel pdiffusion 220 -2153 220 -2153 0 feedthrough
rlabel pdiffusion 227 -2153 227 -2153 0 feedthrough
rlabel pdiffusion 234 -2153 234 -2153 0 feedthrough
rlabel pdiffusion 241 -2153 241 -2153 0 feedthrough
rlabel pdiffusion 248 -2153 248 -2153 0 feedthrough
rlabel pdiffusion 255 -2153 255 -2153 0 feedthrough
rlabel pdiffusion 262 -2153 262 -2153 0 feedthrough
rlabel pdiffusion 269 -2153 269 -2153 0 feedthrough
rlabel pdiffusion 276 -2153 276 -2153 0 feedthrough
rlabel pdiffusion 283 -2153 283 -2153 0 feedthrough
rlabel pdiffusion 290 -2153 290 -2153 0 feedthrough
rlabel pdiffusion 297 -2153 297 -2153 0 cellNo=253
rlabel pdiffusion 304 -2153 304 -2153 0 feedthrough
rlabel pdiffusion 311 -2153 311 -2153 0 feedthrough
rlabel pdiffusion 318 -2153 318 -2153 0 cellNo=140
rlabel pdiffusion 325 -2153 325 -2153 0 feedthrough
rlabel pdiffusion 332 -2153 332 -2153 0 feedthrough
rlabel pdiffusion 339 -2153 339 -2153 0 feedthrough
rlabel pdiffusion 346 -2153 346 -2153 0 feedthrough
rlabel pdiffusion 353 -2153 353 -2153 0 feedthrough
rlabel pdiffusion 360 -2153 360 -2153 0 feedthrough
rlabel pdiffusion 367 -2153 367 -2153 0 feedthrough
rlabel pdiffusion 374 -2153 374 -2153 0 feedthrough
rlabel pdiffusion 381 -2153 381 -2153 0 feedthrough
rlabel pdiffusion 388 -2153 388 -2153 0 feedthrough
rlabel pdiffusion 395 -2153 395 -2153 0 feedthrough
rlabel pdiffusion 402 -2153 402 -2153 0 feedthrough
rlabel pdiffusion 409 -2153 409 -2153 0 feedthrough
rlabel pdiffusion 416 -2153 416 -2153 0 feedthrough
rlabel pdiffusion 423 -2153 423 -2153 0 feedthrough
rlabel pdiffusion 430 -2153 430 -2153 0 feedthrough
rlabel pdiffusion 437 -2153 437 -2153 0 feedthrough
rlabel pdiffusion 444 -2153 444 -2153 0 feedthrough
rlabel pdiffusion 451 -2153 451 -2153 0 feedthrough
rlabel pdiffusion 458 -2153 458 -2153 0 feedthrough
rlabel pdiffusion 465 -2153 465 -2153 0 cellNo=277
rlabel pdiffusion 472 -2153 472 -2153 0 feedthrough
rlabel pdiffusion 479 -2153 479 -2153 0 cellNo=474
rlabel pdiffusion 486 -2153 486 -2153 0 cellNo=12
rlabel pdiffusion 493 -2153 493 -2153 0 feedthrough
rlabel pdiffusion 500 -2153 500 -2153 0 feedthrough
rlabel pdiffusion 507 -2153 507 -2153 0 cellNo=321
rlabel pdiffusion 514 -2153 514 -2153 0 cellNo=259
rlabel pdiffusion 521 -2153 521 -2153 0 feedthrough
rlabel pdiffusion 528 -2153 528 -2153 0 cellNo=588
rlabel pdiffusion 535 -2153 535 -2153 0 feedthrough
rlabel pdiffusion 542 -2153 542 -2153 0 feedthrough
rlabel pdiffusion 549 -2153 549 -2153 0 feedthrough
rlabel pdiffusion 556 -2153 556 -2153 0 feedthrough
rlabel pdiffusion 563 -2153 563 -2153 0 feedthrough
rlabel pdiffusion 570 -2153 570 -2153 0 feedthrough
rlabel pdiffusion 577 -2153 577 -2153 0 feedthrough
rlabel pdiffusion 584 -2153 584 -2153 0 feedthrough
rlabel pdiffusion 591 -2153 591 -2153 0 feedthrough
rlabel pdiffusion 598 -2153 598 -2153 0 cellNo=100
rlabel pdiffusion 605 -2153 605 -2153 0 feedthrough
rlabel pdiffusion 612 -2153 612 -2153 0 cellNo=205
rlabel pdiffusion 619 -2153 619 -2153 0 feedthrough
rlabel pdiffusion 626 -2153 626 -2153 0 feedthrough
rlabel pdiffusion 633 -2153 633 -2153 0 feedthrough
rlabel pdiffusion 640 -2153 640 -2153 0 cellNo=534
rlabel pdiffusion 647 -2153 647 -2153 0 feedthrough
rlabel pdiffusion 654 -2153 654 -2153 0 cellNo=307
rlabel pdiffusion 661 -2153 661 -2153 0 feedthrough
rlabel pdiffusion 668 -2153 668 -2153 0 feedthrough
rlabel pdiffusion 675 -2153 675 -2153 0 feedthrough
rlabel pdiffusion 682 -2153 682 -2153 0 feedthrough
rlabel pdiffusion 689 -2153 689 -2153 0 cellNo=522
rlabel pdiffusion 696 -2153 696 -2153 0 feedthrough
rlabel pdiffusion 703 -2153 703 -2153 0 feedthrough
rlabel pdiffusion 710 -2153 710 -2153 0 feedthrough
rlabel pdiffusion 717 -2153 717 -2153 0 feedthrough
rlabel pdiffusion 724 -2153 724 -2153 0 feedthrough
rlabel pdiffusion 731 -2153 731 -2153 0 feedthrough
rlabel pdiffusion 738 -2153 738 -2153 0 feedthrough
rlabel pdiffusion 745 -2153 745 -2153 0 feedthrough
rlabel pdiffusion 752 -2153 752 -2153 0 feedthrough
rlabel pdiffusion 759 -2153 759 -2153 0 feedthrough
rlabel pdiffusion 766 -2153 766 -2153 0 feedthrough
rlabel pdiffusion 773 -2153 773 -2153 0 feedthrough
rlabel pdiffusion 780 -2153 780 -2153 0 feedthrough
rlabel pdiffusion 787 -2153 787 -2153 0 cellNo=290
rlabel pdiffusion 794 -2153 794 -2153 0 feedthrough
rlabel pdiffusion 801 -2153 801 -2153 0 feedthrough
rlabel pdiffusion 808 -2153 808 -2153 0 feedthrough
rlabel pdiffusion 815 -2153 815 -2153 0 feedthrough
rlabel pdiffusion 822 -2153 822 -2153 0 feedthrough
rlabel pdiffusion 829 -2153 829 -2153 0 feedthrough
rlabel pdiffusion 836 -2153 836 -2153 0 feedthrough
rlabel pdiffusion 843 -2153 843 -2153 0 feedthrough
rlabel pdiffusion 850 -2153 850 -2153 0 feedthrough
rlabel pdiffusion 857 -2153 857 -2153 0 feedthrough
rlabel pdiffusion 864 -2153 864 -2153 0 feedthrough
rlabel pdiffusion 871 -2153 871 -2153 0 feedthrough
rlabel pdiffusion 878 -2153 878 -2153 0 feedthrough
rlabel pdiffusion 885 -2153 885 -2153 0 feedthrough
rlabel pdiffusion 892 -2153 892 -2153 0 feedthrough
rlabel pdiffusion 899 -2153 899 -2153 0 feedthrough
rlabel pdiffusion 906 -2153 906 -2153 0 feedthrough
rlabel pdiffusion 913 -2153 913 -2153 0 feedthrough
rlabel pdiffusion 920 -2153 920 -2153 0 feedthrough
rlabel pdiffusion 927 -2153 927 -2153 0 feedthrough
rlabel pdiffusion 934 -2153 934 -2153 0 feedthrough
rlabel pdiffusion 941 -2153 941 -2153 0 feedthrough
rlabel pdiffusion 948 -2153 948 -2153 0 feedthrough
rlabel pdiffusion 955 -2153 955 -2153 0 feedthrough
rlabel pdiffusion 962 -2153 962 -2153 0 feedthrough
rlabel pdiffusion 969 -2153 969 -2153 0 cellNo=282
rlabel pdiffusion 976 -2153 976 -2153 0 feedthrough
rlabel pdiffusion 983 -2153 983 -2153 0 feedthrough
rlabel pdiffusion 990 -2153 990 -2153 0 feedthrough
rlabel pdiffusion 997 -2153 997 -2153 0 cellNo=475
rlabel pdiffusion 1004 -2153 1004 -2153 0 feedthrough
rlabel pdiffusion 1011 -2153 1011 -2153 0 feedthrough
rlabel pdiffusion 1018 -2153 1018 -2153 0 feedthrough
rlabel pdiffusion 1025 -2153 1025 -2153 0 feedthrough
rlabel pdiffusion 1032 -2153 1032 -2153 0 feedthrough
rlabel pdiffusion 1039 -2153 1039 -2153 0 feedthrough
rlabel pdiffusion 1046 -2153 1046 -2153 0 feedthrough
rlabel pdiffusion 1053 -2153 1053 -2153 0 feedthrough
rlabel pdiffusion 1060 -2153 1060 -2153 0 feedthrough
rlabel pdiffusion 1067 -2153 1067 -2153 0 feedthrough
rlabel pdiffusion 1102 -2153 1102 -2153 0 cellNo=396
rlabel pdiffusion 1109 -2153 1109 -2153 0 feedthrough
rlabel pdiffusion 1123 -2153 1123 -2153 0 feedthrough
rlabel pdiffusion 31 -2234 31 -2234 0 feedthrough
rlabel pdiffusion 38 -2234 38 -2234 0 feedthrough
rlabel pdiffusion 45 -2234 45 -2234 0 feedthrough
rlabel pdiffusion 52 -2234 52 -2234 0 feedthrough
rlabel pdiffusion 59 -2234 59 -2234 0 feedthrough
rlabel pdiffusion 66 -2234 66 -2234 0 feedthrough
rlabel pdiffusion 73 -2234 73 -2234 0 feedthrough
rlabel pdiffusion 80 -2234 80 -2234 0 cellNo=486
rlabel pdiffusion 87 -2234 87 -2234 0 cellNo=435
rlabel pdiffusion 94 -2234 94 -2234 0 cellNo=375
rlabel pdiffusion 101 -2234 101 -2234 0 feedthrough
rlabel pdiffusion 108 -2234 108 -2234 0 feedthrough
rlabel pdiffusion 115 -2234 115 -2234 0 feedthrough
rlabel pdiffusion 122 -2234 122 -2234 0 cellNo=553
rlabel pdiffusion 129 -2234 129 -2234 0 cellNo=403
rlabel pdiffusion 136 -2234 136 -2234 0 feedthrough
rlabel pdiffusion 143 -2234 143 -2234 0 feedthrough
rlabel pdiffusion 150 -2234 150 -2234 0 feedthrough
rlabel pdiffusion 157 -2234 157 -2234 0 feedthrough
rlabel pdiffusion 164 -2234 164 -2234 0 feedthrough
rlabel pdiffusion 171 -2234 171 -2234 0 feedthrough
rlabel pdiffusion 178 -2234 178 -2234 0 cellNo=236
rlabel pdiffusion 185 -2234 185 -2234 0 feedthrough
rlabel pdiffusion 192 -2234 192 -2234 0 feedthrough
rlabel pdiffusion 199 -2234 199 -2234 0 feedthrough
rlabel pdiffusion 206 -2234 206 -2234 0 feedthrough
rlabel pdiffusion 213 -2234 213 -2234 0 feedthrough
rlabel pdiffusion 220 -2234 220 -2234 0 feedthrough
rlabel pdiffusion 227 -2234 227 -2234 0 feedthrough
rlabel pdiffusion 234 -2234 234 -2234 0 feedthrough
rlabel pdiffusion 241 -2234 241 -2234 0 feedthrough
rlabel pdiffusion 248 -2234 248 -2234 0 feedthrough
rlabel pdiffusion 255 -2234 255 -2234 0 feedthrough
rlabel pdiffusion 262 -2234 262 -2234 0 feedthrough
rlabel pdiffusion 269 -2234 269 -2234 0 feedthrough
rlabel pdiffusion 276 -2234 276 -2234 0 feedthrough
rlabel pdiffusion 283 -2234 283 -2234 0 feedthrough
rlabel pdiffusion 290 -2234 290 -2234 0 feedthrough
rlabel pdiffusion 297 -2234 297 -2234 0 feedthrough
rlabel pdiffusion 304 -2234 304 -2234 0 feedthrough
rlabel pdiffusion 311 -2234 311 -2234 0 feedthrough
rlabel pdiffusion 318 -2234 318 -2234 0 feedthrough
rlabel pdiffusion 325 -2234 325 -2234 0 feedthrough
rlabel pdiffusion 332 -2234 332 -2234 0 feedthrough
rlabel pdiffusion 339 -2234 339 -2234 0 feedthrough
rlabel pdiffusion 346 -2234 346 -2234 0 feedthrough
rlabel pdiffusion 353 -2234 353 -2234 0 cellNo=386
rlabel pdiffusion 360 -2234 360 -2234 0 feedthrough
rlabel pdiffusion 367 -2234 367 -2234 0 feedthrough
rlabel pdiffusion 374 -2234 374 -2234 0 feedthrough
rlabel pdiffusion 381 -2234 381 -2234 0 feedthrough
rlabel pdiffusion 388 -2234 388 -2234 0 feedthrough
rlabel pdiffusion 395 -2234 395 -2234 0 cellNo=117
rlabel pdiffusion 402 -2234 402 -2234 0 feedthrough
rlabel pdiffusion 409 -2234 409 -2234 0 feedthrough
rlabel pdiffusion 416 -2234 416 -2234 0 feedthrough
rlabel pdiffusion 423 -2234 423 -2234 0 feedthrough
rlabel pdiffusion 430 -2234 430 -2234 0 feedthrough
rlabel pdiffusion 437 -2234 437 -2234 0 feedthrough
rlabel pdiffusion 444 -2234 444 -2234 0 cellNo=287
rlabel pdiffusion 451 -2234 451 -2234 0 cellNo=464
rlabel pdiffusion 458 -2234 458 -2234 0 feedthrough
rlabel pdiffusion 465 -2234 465 -2234 0 feedthrough
rlabel pdiffusion 472 -2234 472 -2234 0 feedthrough
rlabel pdiffusion 479 -2234 479 -2234 0 cellNo=362
rlabel pdiffusion 486 -2234 486 -2234 0 cellNo=412
rlabel pdiffusion 493 -2234 493 -2234 0 feedthrough
rlabel pdiffusion 500 -2234 500 -2234 0 feedthrough
rlabel pdiffusion 507 -2234 507 -2234 0 feedthrough
rlabel pdiffusion 514 -2234 514 -2234 0 feedthrough
rlabel pdiffusion 521 -2234 521 -2234 0 feedthrough
rlabel pdiffusion 528 -2234 528 -2234 0 cellNo=135
rlabel pdiffusion 535 -2234 535 -2234 0 feedthrough
rlabel pdiffusion 542 -2234 542 -2234 0 feedthrough
rlabel pdiffusion 549 -2234 549 -2234 0 feedthrough
rlabel pdiffusion 556 -2234 556 -2234 0 feedthrough
rlabel pdiffusion 563 -2234 563 -2234 0 feedthrough
rlabel pdiffusion 570 -2234 570 -2234 0 feedthrough
rlabel pdiffusion 577 -2234 577 -2234 0 feedthrough
rlabel pdiffusion 584 -2234 584 -2234 0 feedthrough
rlabel pdiffusion 591 -2234 591 -2234 0 feedthrough
rlabel pdiffusion 598 -2234 598 -2234 0 feedthrough
rlabel pdiffusion 605 -2234 605 -2234 0 feedthrough
rlabel pdiffusion 612 -2234 612 -2234 0 feedthrough
rlabel pdiffusion 619 -2234 619 -2234 0 feedthrough
rlabel pdiffusion 626 -2234 626 -2234 0 feedthrough
rlabel pdiffusion 633 -2234 633 -2234 0 feedthrough
rlabel pdiffusion 640 -2234 640 -2234 0 feedthrough
rlabel pdiffusion 647 -2234 647 -2234 0 feedthrough
rlabel pdiffusion 654 -2234 654 -2234 0 cellNo=493
rlabel pdiffusion 661 -2234 661 -2234 0 feedthrough
rlabel pdiffusion 668 -2234 668 -2234 0 cellNo=360
rlabel pdiffusion 675 -2234 675 -2234 0 feedthrough
rlabel pdiffusion 682 -2234 682 -2234 0 feedthrough
rlabel pdiffusion 689 -2234 689 -2234 0 feedthrough
rlabel pdiffusion 696 -2234 696 -2234 0 cellNo=155
rlabel pdiffusion 703 -2234 703 -2234 0 feedthrough
rlabel pdiffusion 710 -2234 710 -2234 0 feedthrough
rlabel pdiffusion 717 -2234 717 -2234 0 feedthrough
rlabel pdiffusion 724 -2234 724 -2234 0 feedthrough
rlabel pdiffusion 731 -2234 731 -2234 0 feedthrough
rlabel pdiffusion 738 -2234 738 -2234 0 cellNo=80
rlabel pdiffusion 745 -2234 745 -2234 0 cellNo=120
rlabel pdiffusion 752 -2234 752 -2234 0 feedthrough
rlabel pdiffusion 759 -2234 759 -2234 0 feedthrough
rlabel pdiffusion 766 -2234 766 -2234 0 feedthrough
rlabel pdiffusion 773 -2234 773 -2234 0 feedthrough
rlabel pdiffusion 780 -2234 780 -2234 0 feedthrough
rlabel pdiffusion 787 -2234 787 -2234 0 feedthrough
rlabel pdiffusion 794 -2234 794 -2234 0 feedthrough
rlabel pdiffusion 801 -2234 801 -2234 0 feedthrough
rlabel pdiffusion 808 -2234 808 -2234 0 feedthrough
rlabel pdiffusion 815 -2234 815 -2234 0 feedthrough
rlabel pdiffusion 822 -2234 822 -2234 0 feedthrough
rlabel pdiffusion 829 -2234 829 -2234 0 feedthrough
rlabel pdiffusion 836 -2234 836 -2234 0 feedthrough
rlabel pdiffusion 843 -2234 843 -2234 0 feedthrough
rlabel pdiffusion 850 -2234 850 -2234 0 feedthrough
rlabel pdiffusion 857 -2234 857 -2234 0 feedthrough
rlabel pdiffusion 864 -2234 864 -2234 0 feedthrough
rlabel pdiffusion 871 -2234 871 -2234 0 feedthrough
rlabel pdiffusion 878 -2234 878 -2234 0 feedthrough
rlabel pdiffusion 885 -2234 885 -2234 0 feedthrough
rlabel pdiffusion 892 -2234 892 -2234 0 feedthrough
rlabel pdiffusion 899 -2234 899 -2234 0 feedthrough
rlabel pdiffusion 906 -2234 906 -2234 0 feedthrough
rlabel pdiffusion 913 -2234 913 -2234 0 feedthrough
rlabel pdiffusion 920 -2234 920 -2234 0 feedthrough
rlabel pdiffusion 927 -2234 927 -2234 0 feedthrough
rlabel pdiffusion 934 -2234 934 -2234 0 feedthrough
rlabel pdiffusion 941 -2234 941 -2234 0 cellNo=598
rlabel pdiffusion 948 -2234 948 -2234 0 feedthrough
rlabel pdiffusion 955 -2234 955 -2234 0 cellNo=212
rlabel pdiffusion 962 -2234 962 -2234 0 feedthrough
rlabel pdiffusion 969 -2234 969 -2234 0 feedthrough
rlabel pdiffusion 976 -2234 976 -2234 0 feedthrough
rlabel pdiffusion 983 -2234 983 -2234 0 feedthrough
rlabel pdiffusion 997 -2234 997 -2234 0 feedthrough
rlabel pdiffusion 1004 -2234 1004 -2234 0 feedthrough
rlabel pdiffusion 1018 -2234 1018 -2234 0 feedthrough
rlabel pdiffusion 1067 -2234 1067 -2234 0 feedthrough
rlabel pdiffusion 45 -2317 45 -2317 0 feedthrough
rlabel pdiffusion 52 -2317 52 -2317 0 feedthrough
rlabel pdiffusion 59 -2317 59 -2317 0 feedthrough
rlabel pdiffusion 66 -2317 66 -2317 0 feedthrough
rlabel pdiffusion 73 -2317 73 -2317 0 feedthrough
rlabel pdiffusion 80 -2317 80 -2317 0 feedthrough
rlabel pdiffusion 87 -2317 87 -2317 0 cellNo=366
rlabel pdiffusion 94 -2317 94 -2317 0 feedthrough
rlabel pdiffusion 101 -2317 101 -2317 0 feedthrough
rlabel pdiffusion 108 -2317 108 -2317 0 feedthrough
rlabel pdiffusion 115 -2317 115 -2317 0 feedthrough
rlabel pdiffusion 122 -2317 122 -2317 0 feedthrough
rlabel pdiffusion 129 -2317 129 -2317 0 feedthrough
rlabel pdiffusion 136 -2317 136 -2317 0 cellNo=303
rlabel pdiffusion 143 -2317 143 -2317 0 feedthrough
rlabel pdiffusion 150 -2317 150 -2317 0 feedthrough
rlabel pdiffusion 157 -2317 157 -2317 0 feedthrough
rlabel pdiffusion 164 -2317 164 -2317 0 feedthrough
rlabel pdiffusion 171 -2317 171 -2317 0 feedthrough
rlabel pdiffusion 178 -2317 178 -2317 0 feedthrough
rlabel pdiffusion 185 -2317 185 -2317 0 cellNo=101
rlabel pdiffusion 192 -2317 192 -2317 0 feedthrough
rlabel pdiffusion 199 -2317 199 -2317 0 feedthrough
rlabel pdiffusion 206 -2317 206 -2317 0 feedthrough
rlabel pdiffusion 213 -2317 213 -2317 0 feedthrough
rlabel pdiffusion 220 -2317 220 -2317 0 feedthrough
rlabel pdiffusion 227 -2317 227 -2317 0 feedthrough
rlabel pdiffusion 234 -2317 234 -2317 0 feedthrough
rlabel pdiffusion 241 -2317 241 -2317 0 feedthrough
rlabel pdiffusion 248 -2317 248 -2317 0 feedthrough
rlabel pdiffusion 255 -2317 255 -2317 0 feedthrough
rlabel pdiffusion 262 -2317 262 -2317 0 feedthrough
rlabel pdiffusion 269 -2317 269 -2317 0 feedthrough
rlabel pdiffusion 276 -2317 276 -2317 0 feedthrough
rlabel pdiffusion 283 -2317 283 -2317 0 feedthrough
rlabel pdiffusion 290 -2317 290 -2317 0 cellNo=38
rlabel pdiffusion 297 -2317 297 -2317 0 feedthrough
rlabel pdiffusion 304 -2317 304 -2317 0 feedthrough
rlabel pdiffusion 311 -2317 311 -2317 0 feedthrough
rlabel pdiffusion 318 -2317 318 -2317 0 feedthrough
rlabel pdiffusion 325 -2317 325 -2317 0 feedthrough
rlabel pdiffusion 332 -2317 332 -2317 0 feedthrough
rlabel pdiffusion 339 -2317 339 -2317 0 feedthrough
rlabel pdiffusion 346 -2317 346 -2317 0 cellNo=570
rlabel pdiffusion 353 -2317 353 -2317 0 feedthrough
rlabel pdiffusion 360 -2317 360 -2317 0 feedthrough
rlabel pdiffusion 367 -2317 367 -2317 0 feedthrough
rlabel pdiffusion 374 -2317 374 -2317 0 cellNo=227
rlabel pdiffusion 381 -2317 381 -2317 0 feedthrough
rlabel pdiffusion 388 -2317 388 -2317 0 feedthrough
rlabel pdiffusion 395 -2317 395 -2317 0 feedthrough
rlabel pdiffusion 402 -2317 402 -2317 0 feedthrough
rlabel pdiffusion 409 -2317 409 -2317 0 feedthrough
rlabel pdiffusion 416 -2317 416 -2317 0 feedthrough
rlabel pdiffusion 423 -2317 423 -2317 0 cellNo=20
rlabel pdiffusion 430 -2317 430 -2317 0 feedthrough
rlabel pdiffusion 437 -2317 437 -2317 0 feedthrough
rlabel pdiffusion 444 -2317 444 -2317 0 cellNo=432
rlabel pdiffusion 451 -2317 451 -2317 0 cellNo=312
rlabel pdiffusion 458 -2317 458 -2317 0 feedthrough
rlabel pdiffusion 465 -2317 465 -2317 0 feedthrough
rlabel pdiffusion 472 -2317 472 -2317 0 feedthrough
rlabel pdiffusion 479 -2317 479 -2317 0 feedthrough
rlabel pdiffusion 486 -2317 486 -2317 0 feedthrough
rlabel pdiffusion 493 -2317 493 -2317 0 cellNo=163
rlabel pdiffusion 500 -2317 500 -2317 0 feedthrough
rlabel pdiffusion 507 -2317 507 -2317 0 feedthrough
rlabel pdiffusion 514 -2317 514 -2317 0 feedthrough
rlabel pdiffusion 521 -2317 521 -2317 0 feedthrough
rlabel pdiffusion 528 -2317 528 -2317 0 feedthrough
rlabel pdiffusion 535 -2317 535 -2317 0 cellNo=450
rlabel pdiffusion 542 -2317 542 -2317 0 feedthrough
rlabel pdiffusion 549 -2317 549 -2317 0 feedthrough
rlabel pdiffusion 556 -2317 556 -2317 0 feedthrough
rlabel pdiffusion 563 -2317 563 -2317 0 cellNo=381
rlabel pdiffusion 570 -2317 570 -2317 0 cellNo=586
rlabel pdiffusion 577 -2317 577 -2317 0 cellNo=328
rlabel pdiffusion 584 -2317 584 -2317 0 feedthrough
rlabel pdiffusion 591 -2317 591 -2317 0 feedthrough
rlabel pdiffusion 598 -2317 598 -2317 0 feedthrough
rlabel pdiffusion 605 -2317 605 -2317 0 feedthrough
rlabel pdiffusion 612 -2317 612 -2317 0 feedthrough
rlabel pdiffusion 619 -2317 619 -2317 0 cellNo=305
rlabel pdiffusion 626 -2317 626 -2317 0 feedthrough
rlabel pdiffusion 633 -2317 633 -2317 0 feedthrough
rlabel pdiffusion 640 -2317 640 -2317 0 feedthrough
rlabel pdiffusion 647 -2317 647 -2317 0 feedthrough
rlabel pdiffusion 654 -2317 654 -2317 0 cellNo=574
rlabel pdiffusion 661 -2317 661 -2317 0 feedthrough
rlabel pdiffusion 668 -2317 668 -2317 0 feedthrough
rlabel pdiffusion 675 -2317 675 -2317 0 feedthrough
rlabel pdiffusion 682 -2317 682 -2317 0 feedthrough
rlabel pdiffusion 689 -2317 689 -2317 0 feedthrough
rlabel pdiffusion 696 -2317 696 -2317 0 feedthrough
rlabel pdiffusion 703 -2317 703 -2317 0 feedthrough
rlabel pdiffusion 710 -2317 710 -2317 0 feedthrough
rlabel pdiffusion 717 -2317 717 -2317 0 feedthrough
rlabel pdiffusion 724 -2317 724 -2317 0 feedthrough
rlabel pdiffusion 731 -2317 731 -2317 0 feedthrough
rlabel pdiffusion 738 -2317 738 -2317 0 feedthrough
rlabel pdiffusion 745 -2317 745 -2317 0 feedthrough
rlabel pdiffusion 752 -2317 752 -2317 0 feedthrough
rlabel pdiffusion 759 -2317 759 -2317 0 feedthrough
rlabel pdiffusion 766 -2317 766 -2317 0 feedthrough
rlabel pdiffusion 773 -2317 773 -2317 0 feedthrough
rlabel pdiffusion 780 -2317 780 -2317 0 feedthrough
rlabel pdiffusion 787 -2317 787 -2317 0 feedthrough
rlabel pdiffusion 794 -2317 794 -2317 0 feedthrough
rlabel pdiffusion 801 -2317 801 -2317 0 cellNo=133
rlabel pdiffusion 808 -2317 808 -2317 0 feedthrough
rlabel pdiffusion 815 -2317 815 -2317 0 feedthrough
rlabel pdiffusion 822 -2317 822 -2317 0 feedthrough
rlabel pdiffusion 829 -2317 829 -2317 0 feedthrough
rlabel pdiffusion 836 -2317 836 -2317 0 feedthrough
rlabel pdiffusion 843 -2317 843 -2317 0 feedthrough
rlabel pdiffusion 850 -2317 850 -2317 0 feedthrough
rlabel pdiffusion 857 -2317 857 -2317 0 feedthrough
rlabel pdiffusion 864 -2317 864 -2317 0 feedthrough
rlabel pdiffusion 871 -2317 871 -2317 0 feedthrough
rlabel pdiffusion 878 -2317 878 -2317 0 feedthrough
rlabel pdiffusion 885 -2317 885 -2317 0 feedthrough
rlabel pdiffusion 892 -2317 892 -2317 0 feedthrough
rlabel pdiffusion 899 -2317 899 -2317 0 feedthrough
rlabel pdiffusion 969 -2317 969 -2317 0 feedthrough
rlabel pdiffusion 990 -2317 990 -2317 0 feedthrough
rlabel pdiffusion 997 -2317 997 -2317 0 feedthrough
rlabel pdiffusion 1039 -2317 1039 -2317 0 feedthrough
rlabel pdiffusion 1060 -2317 1060 -2317 0 cellNo=318
rlabel pdiffusion 73 -2382 73 -2382 0 feedthrough
rlabel pdiffusion 80 -2382 80 -2382 0 feedthrough
rlabel pdiffusion 87 -2382 87 -2382 0 feedthrough
rlabel pdiffusion 94 -2382 94 -2382 0 feedthrough
rlabel pdiffusion 101 -2382 101 -2382 0 feedthrough
rlabel pdiffusion 108 -2382 108 -2382 0 feedthrough
rlabel pdiffusion 115 -2382 115 -2382 0 feedthrough
rlabel pdiffusion 122 -2382 122 -2382 0 feedthrough
rlabel pdiffusion 129 -2382 129 -2382 0 feedthrough
rlabel pdiffusion 136 -2382 136 -2382 0 feedthrough
rlabel pdiffusion 143 -2382 143 -2382 0 feedthrough
rlabel pdiffusion 150 -2382 150 -2382 0 cellNo=461
rlabel pdiffusion 157 -2382 157 -2382 0 feedthrough
rlabel pdiffusion 164 -2382 164 -2382 0 cellNo=345
rlabel pdiffusion 171 -2382 171 -2382 0 cellNo=247
rlabel pdiffusion 178 -2382 178 -2382 0 cellNo=95
rlabel pdiffusion 185 -2382 185 -2382 0 cellNo=404
rlabel pdiffusion 192 -2382 192 -2382 0 feedthrough
rlabel pdiffusion 199 -2382 199 -2382 0 feedthrough
rlabel pdiffusion 206 -2382 206 -2382 0 feedthrough
rlabel pdiffusion 213 -2382 213 -2382 0 feedthrough
rlabel pdiffusion 220 -2382 220 -2382 0 feedthrough
rlabel pdiffusion 227 -2382 227 -2382 0 feedthrough
rlabel pdiffusion 234 -2382 234 -2382 0 cellNo=61
rlabel pdiffusion 241 -2382 241 -2382 0 feedthrough
rlabel pdiffusion 248 -2382 248 -2382 0 feedthrough
rlabel pdiffusion 255 -2382 255 -2382 0 feedthrough
rlabel pdiffusion 262 -2382 262 -2382 0 feedthrough
rlabel pdiffusion 269 -2382 269 -2382 0 cellNo=159
rlabel pdiffusion 276 -2382 276 -2382 0 feedthrough
rlabel pdiffusion 283 -2382 283 -2382 0 feedthrough
rlabel pdiffusion 290 -2382 290 -2382 0 feedthrough
rlabel pdiffusion 297 -2382 297 -2382 0 feedthrough
rlabel pdiffusion 304 -2382 304 -2382 0 cellNo=532
rlabel pdiffusion 311 -2382 311 -2382 0 feedthrough
rlabel pdiffusion 318 -2382 318 -2382 0 feedthrough
rlabel pdiffusion 325 -2382 325 -2382 0 feedthrough
rlabel pdiffusion 332 -2382 332 -2382 0 feedthrough
rlabel pdiffusion 339 -2382 339 -2382 0 feedthrough
rlabel pdiffusion 346 -2382 346 -2382 0 feedthrough
rlabel pdiffusion 353 -2382 353 -2382 0 feedthrough
rlabel pdiffusion 360 -2382 360 -2382 0 feedthrough
rlabel pdiffusion 367 -2382 367 -2382 0 feedthrough
rlabel pdiffusion 374 -2382 374 -2382 0 feedthrough
rlabel pdiffusion 381 -2382 381 -2382 0 cellNo=334
rlabel pdiffusion 388 -2382 388 -2382 0 feedthrough
rlabel pdiffusion 395 -2382 395 -2382 0 feedthrough
rlabel pdiffusion 402 -2382 402 -2382 0 feedthrough
rlabel pdiffusion 409 -2382 409 -2382 0 feedthrough
rlabel pdiffusion 416 -2382 416 -2382 0 feedthrough
rlabel pdiffusion 423 -2382 423 -2382 0 feedthrough
rlabel pdiffusion 430 -2382 430 -2382 0 feedthrough
rlabel pdiffusion 437 -2382 437 -2382 0 feedthrough
rlabel pdiffusion 444 -2382 444 -2382 0 feedthrough
rlabel pdiffusion 451 -2382 451 -2382 0 cellNo=557
rlabel pdiffusion 458 -2382 458 -2382 0 feedthrough
rlabel pdiffusion 465 -2382 465 -2382 0 feedthrough
rlabel pdiffusion 472 -2382 472 -2382 0 feedthrough
rlabel pdiffusion 479 -2382 479 -2382 0 feedthrough
rlabel pdiffusion 486 -2382 486 -2382 0 feedthrough
rlabel pdiffusion 493 -2382 493 -2382 0 feedthrough
rlabel pdiffusion 500 -2382 500 -2382 0 feedthrough
rlabel pdiffusion 507 -2382 507 -2382 0 feedthrough
rlabel pdiffusion 514 -2382 514 -2382 0 cellNo=424
rlabel pdiffusion 521 -2382 521 -2382 0 feedthrough
rlabel pdiffusion 528 -2382 528 -2382 0 cellNo=298
rlabel pdiffusion 535 -2382 535 -2382 0 feedthrough
rlabel pdiffusion 542 -2382 542 -2382 0 feedthrough
rlabel pdiffusion 549 -2382 549 -2382 0 feedthrough
rlabel pdiffusion 556 -2382 556 -2382 0 cellNo=40
rlabel pdiffusion 563 -2382 563 -2382 0 feedthrough
rlabel pdiffusion 570 -2382 570 -2382 0 feedthrough
rlabel pdiffusion 577 -2382 577 -2382 0 feedthrough
rlabel pdiffusion 584 -2382 584 -2382 0 feedthrough
rlabel pdiffusion 591 -2382 591 -2382 0 feedthrough
rlabel pdiffusion 598 -2382 598 -2382 0 feedthrough
rlabel pdiffusion 605 -2382 605 -2382 0 feedthrough
rlabel pdiffusion 612 -2382 612 -2382 0 cellNo=473
rlabel pdiffusion 619 -2382 619 -2382 0 feedthrough
rlabel pdiffusion 626 -2382 626 -2382 0 feedthrough
rlabel pdiffusion 633 -2382 633 -2382 0 feedthrough
rlabel pdiffusion 640 -2382 640 -2382 0 feedthrough
rlabel pdiffusion 647 -2382 647 -2382 0 feedthrough
rlabel pdiffusion 654 -2382 654 -2382 0 feedthrough
rlabel pdiffusion 661 -2382 661 -2382 0 feedthrough
rlabel pdiffusion 668 -2382 668 -2382 0 feedthrough
rlabel pdiffusion 675 -2382 675 -2382 0 feedthrough
rlabel pdiffusion 682 -2382 682 -2382 0 feedthrough
rlabel pdiffusion 689 -2382 689 -2382 0 feedthrough
rlabel pdiffusion 696 -2382 696 -2382 0 cellNo=430
rlabel pdiffusion 703 -2382 703 -2382 0 feedthrough
rlabel pdiffusion 710 -2382 710 -2382 0 feedthrough
rlabel pdiffusion 717 -2382 717 -2382 0 feedthrough
rlabel pdiffusion 731 -2382 731 -2382 0 feedthrough
rlabel pdiffusion 738 -2382 738 -2382 0 feedthrough
rlabel pdiffusion 745 -2382 745 -2382 0 feedthrough
rlabel pdiffusion 752 -2382 752 -2382 0 feedthrough
rlabel pdiffusion 759 -2382 759 -2382 0 feedthrough
rlabel pdiffusion 766 -2382 766 -2382 0 feedthrough
rlabel pdiffusion 773 -2382 773 -2382 0 feedthrough
rlabel pdiffusion 780 -2382 780 -2382 0 feedthrough
rlabel pdiffusion 794 -2382 794 -2382 0 feedthrough
rlabel pdiffusion 801 -2382 801 -2382 0 feedthrough
rlabel pdiffusion 815 -2382 815 -2382 0 feedthrough
rlabel pdiffusion 899 -2382 899 -2382 0 feedthrough
rlabel pdiffusion 906 -2382 906 -2382 0 feedthrough
rlabel pdiffusion 941 -2382 941 -2382 0 feedthrough
rlabel pdiffusion 976 -2382 976 -2382 0 cellNo=269
rlabel pdiffusion 983 -2382 983 -2382 0 feedthrough
rlabel pdiffusion 990 -2382 990 -2382 0 feedthrough
rlabel pdiffusion 1004 -2382 1004 -2382 0 cellNo=409
rlabel pdiffusion 199 -2433 199 -2433 0 feedthrough
rlabel pdiffusion 220 -2433 220 -2433 0 feedthrough
rlabel pdiffusion 227 -2433 227 -2433 0 feedthrough
rlabel pdiffusion 234 -2433 234 -2433 0 feedthrough
rlabel pdiffusion 241 -2433 241 -2433 0 feedthrough
rlabel pdiffusion 248 -2433 248 -2433 0 feedthrough
rlabel pdiffusion 255 -2433 255 -2433 0 feedthrough
rlabel pdiffusion 262 -2433 262 -2433 0 feedthrough
rlabel pdiffusion 269 -2433 269 -2433 0 feedthrough
rlabel pdiffusion 276 -2433 276 -2433 0 feedthrough
rlabel pdiffusion 283 -2433 283 -2433 0 feedthrough
rlabel pdiffusion 290 -2433 290 -2433 0 feedthrough
rlabel pdiffusion 297 -2433 297 -2433 0 feedthrough
rlabel pdiffusion 304 -2433 304 -2433 0 feedthrough
rlabel pdiffusion 311 -2433 311 -2433 0 feedthrough
rlabel pdiffusion 318 -2433 318 -2433 0 feedthrough
rlabel pdiffusion 325 -2433 325 -2433 0 cellNo=339
rlabel pdiffusion 332 -2433 332 -2433 0 feedthrough
rlabel pdiffusion 339 -2433 339 -2433 0 feedthrough
rlabel pdiffusion 346 -2433 346 -2433 0 feedthrough
rlabel pdiffusion 353 -2433 353 -2433 0 cellNo=308
rlabel pdiffusion 360 -2433 360 -2433 0 feedthrough
rlabel pdiffusion 367 -2433 367 -2433 0 cellNo=477
rlabel pdiffusion 374 -2433 374 -2433 0 feedthrough
rlabel pdiffusion 381 -2433 381 -2433 0 cellNo=378
rlabel pdiffusion 388 -2433 388 -2433 0 feedthrough
rlabel pdiffusion 395 -2433 395 -2433 0 feedthrough
rlabel pdiffusion 402 -2433 402 -2433 0 feedthrough
rlabel pdiffusion 409 -2433 409 -2433 0 feedthrough
rlabel pdiffusion 416 -2433 416 -2433 0 cellNo=371
rlabel pdiffusion 423 -2433 423 -2433 0 feedthrough
rlabel pdiffusion 430 -2433 430 -2433 0 feedthrough
rlabel pdiffusion 437 -2433 437 -2433 0 feedthrough
rlabel pdiffusion 444 -2433 444 -2433 0 feedthrough
rlabel pdiffusion 451 -2433 451 -2433 0 cellNo=427
rlabel pdiffusion 458 -2433 458 -2433 0 cellNo=571
rlabel pdiffusion 465 -2433 465 -2433 0 feedthrough
rlabel pdiffusion 472 -2433 472 -2433 0 feedthrough
rlabel pdiffusion 479 -2433 479 -2433 0 feedthrough
rlabel pdiffusion 486 -2433 486 -2433 0 cellNo=280
rlabel pdiffusion 493 -2433 493 -2433 0 feedthrough
rlabel pdiffusion 500 -2433 500 -2433 0 feedthrough
rlabel pdiffusion 507 -2433 507 -2433 0 cellNo=541
rlabel pdiffusion 514 -2433 514 -2433 0 cellNo=382
rlabel pdiffusion 521 -2433 521 -2433 0 cellNo=248
rlabel pdiffusion 528 -2433 528 -2433 0 feedthrough
rlabel pdiffusion 535 -2433 535 -2433 0 feedthrough
rlabel pdiffusion 542 -2433 542 -2433 0 feedthrough
rlabel pdiffusion 549 -2433 549 -2433 0 feedthrough
rlabel pdiffusion 556 -2433 556 -2433 0 feedthrough
rlabel pdiffusion 563 -2433 563 -2433 0 feedthrough
rlabel pdiffusion 570 -2433 570 -2433 0 cellNo=521
rlabel pdiffusion 577 -2433 577 -2433 0 feedthrough
rlabel pdiffusion 584 -2433 584 -2433 0 feedthrough
rlabel pdiffusion 591 -2433 591 -2433 0 feedthrough
rlabel pdiffusion 598 -2433 598 -2433 0 feedthrough
rlabel pdiffusion 605 -2433 605 -2433 0 feedthrough
rlabel pdiffusion 612 -2433 612 -2433 0 feedthrough
rlabel pdiffusion 619 -2433 619 -2433 0 feedthrough
rlabel pdiffusion 626 -2433 626 -2433 0 feedthrough
rlabel pdiffusion 633 -2433 633 -2433 0 feedthrough
rlabel pdiffusion 647 -2433 647 -2433 0 feedthrough
rlabel pdiffusion 654 -2433 654 -2433 0 feedthrough
rlabel pdiffusion 661 -2433 661 -2433 0 feedthrough
rlabel pdiffusion 668 -2433 668 -2433 0 feedthrough
rlabel pdiffusion 675 -2433 675 -2433 0 feedthrough
rlabel pdiffusion 682 -2433 682 -2433 0 cellNo=581
rlabel pdiffusion 689 -2433 689 -2433 0 cellNo=275
rlabel pdiffusion 717 -2433 717 -2433 0 feedthrough
rlabel pdiffusion 724 -2433 724 -2433 0 feedthrough
rlabel pdiffusion 731 -2433 731 -2433 0 feedthrough
rlabel pdiffusion 738 -2433 738 -2433 0 feedthrough
rlabel pdiffusion 745 -2433 745 -2433 0 cellNo=592
rlabel pdiffusion 752 -2433 752 -2433 0 feedthrough
rlabel pdiffusion 759 -2433 759 -2433 0 feedthrough
rlabel pdiffusion 766 -2433 766 -2433 0 feedthrough
rlabel pdiffusion 773 -2433 773 -2433 0 feedthrough
rlabel pdiffusion 801 -2433 801 -2433 0 feedthrough
rlabel pdiffusion 808 -2433 808 -2433 0 feedthrough
rlabel pdiffusion 829 -2433 829 -2433 0 feedthrough
rlabel pdiffusion 892 -2433 892 -2433 0 feedthrough
rlabel pdiffusion 899 -2433 899 -2433 0 feedthrough
rlabel pdiffusion 906 -2433 906 -2433 0 cellNo=575
rlabel pdiffusion 227 -2474 227 -2474 0 feedthrough
rlabel pdiffusion 234 -2474 234 -2474 0 cellNo=48
rlabel pdiffusion 241 -2474 241 -2474 0 feedthrough
rlabel pdiffusion 248 -2474 248 -2474 0 feedthrough
rlabel pdiffusion 255 -2474 255 -2474 0 cellNo=97
rlabel pdiffusion 297 -2474 297 -2474 0 feedthrough
rlabel pdiffusion 311 -2474 311 -2474 0 feedthrough
rlabel pdiffusion 332 -2474 332 -2474 0 feedthrough
rlabel pdiffusion 339 -2474 339 -2474 0 cellNo=165
rlabel pdiffusion 346 -2474 346 -2474 0 cellNo=542
rlabel pdiffusion 353 -2474 353 -2474 0 feedthrough
rlabel pdiffusion 360 -2474 360 -2474 0 feedthrough
rlabel pdiffusion 367 -2474 367 -2474 0 feedthrough
rlabel pdiffusion 374 -2474 374 -2474 0 feedthrough
rlabel pdiffusion 388 -2474 388 -2474 0 feedthrough
rlabel pdiffusion 395 -2474 395 -2474 0 feedthrough
rlabel pdiffusion 402 -2474 402 -2474 0 feedthrough
rlabel pdiffusion 409 -2474 409 -2474 0 feedthrough
rlabel pdiffusion 423 -2474 423 -2474 0 feedthrough
rlabel pdiffusion 430 -2474 430 -2474 0 cellNo=479
rlabel pdiffusion 437 -2474 437 -2474 0 feedthrough
rlabel pdiffusion 444 -2474 444 -2474 0 cellNo=491
rlabel pdiffusion 451 -2474 451 -2474 0 cellNo=463
rlabel pdiffusion 458 -2474 458 -2474 0 feedthrough
rlabel pdiffusion 465 -2474 465 -2474 0 feedthrough
rlabel pdiffusion 472 -2474 472 -2474 0 feedthrough
rlabel pdiffusion 479 -2474 479 -2474 0 feedthrough
rlabel pdiffusion 486 -2474 486 -2474 0 feedthrough
rlabel pdiffusion 493 -2474 493 -2474 0 feedthrough
rlabel pdiffusion 500 -2474 500 -2474 0 feedthrough
rlabel pdiffusion 507 -2474 507 -2474 0 cellNo=68
rlabel pdiffusion 514 -2474 514 -2474 0 feedthrough
rlabel pdiffusion 528 -2474 528 -2474 0 feedthrough
rlabel pdiffusion 542 -2474 542 -2474 0 feedthrough
rlabel pdiffusion 549 -2474 549 -2474 0 feedthrough
rlabel pdiffusion 577 -2474 577 -2474 0 feedthrough
rlabel pdiffusion 598 -2474 598 -2474 0 feedthrough
rlabel pdiffusion 605 -2474 605 -2474 0 cellNo=207
rlabel pdiffusion 612 -2474 612 -2474 0 cellNo=494
rlabel pdiffusion 619 -2474 619 -2474 0 feedthrough
rlabel pdiffusion 626 -2474 626 -2474 0 feedthrough
rlabel pdiffusion 633 -2474 633 -2474 0 feedthrough
rlabel pdiffusion 640 -2474 640 -2474 0 feedthrough
rlabel pdiffusion 647 -2474 647 -2474 0 cellNo=502
rlabel pdiffusion 654 -2474 654 -2474 0 feedthrough
rlabel pdiffusion 661 -2474 661 -2474 0 feedthrough
rlabel pdiffusion 675 -2474 675 -2474 0 feedthrough
rlabel pdiffusion 689 -2474 689 -2474 0 feedthrough
rlabel pdiffusion 703 -2474 703 -2474 0 feedthrough
rlabel pdiffusion 724 -2474 724 -2474 0 feedthrough
rlabel pdiffusion 745 -2474 745 -2474 0 feedthrough
rlabel pdiffusion 752 -2474 752 -2474 0 cellNo=278
rlabel pdiffusion 808 -2474 808 -2474 0 feedthrough
rlabel pdiffusion 815 -2474 815 -2474 0 cellNo=244
rlabel pdiffusion 829 -2474 829 -2474 0 feedthrough
rlabel pdiffusion 836 -2474 836 -2474 0 cellNo=538
rlabel pdiffusion 899 -2474 899 -2474 0 feedthrough
rlabel pdiffusion 227 -2495 227 -2495 0 feedthrough
rlabel pdiffusion 234 -2495 234 -2495 0 cellNo=329
rlabel pdiffusion 241 -2495 241 -2495 0 feedthrough
rlabel pdiffusion 360 -2495 360 -2495 0 feedthrough
rlabel pdiffusion 367 -2495 367 -2495 0 cellNo=255
rlabel pdiffusion 374 -2495 374 -2495 0 feedthrough
rlabel pdiffusion 381 -2495 381 -2495 0 feedthrough
rlabel pdiffusion 388 -2495 388 -2495 0 cellNo=256
rlabel pdiffusion 395 -2495 395 -2495 0 cellNo=349
rlabel pdiffusion 402 -2495 402 -2495 0 cellNo=417
rlabel pdiffusion 409 -2495 409 -2495 0 feedthrough
rlabel pdiffusion 535 -2495 535 -2495 0 feedthrough
rlabel pdiffusion 549 -2495 549 -2495 0 cellNo=597
rlabel pdiffusion 556 -2495 556 -2495 0 cellNo=599
rlabel pdiffusion 605 -2495 605 -2495 0 feedthrough
rlabel pdiffusion 612 -2495 612 -2495 0 cellNo=530
rlabel pdiffusion 633 -2495 633 -2495 0 feedthrough
rlabel pdiffusion 654 -2495 654 -2495 0 cellNo=296
rlabel pdiffusion 661 -2495 661 -2495 0 feedthrough
rlabel pdiffusion 689 -2495 689 -2495 0 cellNo=511
rlabel pdiffusion 703 -2495 703 -2495 0 feedthrough
rlabel pdiffusion 724 -2495 724 -2495 0 cellNo=508
rlabel pdiffusion 899 -2495 899 -2495 0 cellNo=368
rlabel pdiffusion 906 -2495 906 -2495 0 feedthrough
rlabel polysilicon 152 -6 152 -6 0 2
rlabel polysilicon 149 -12 149 -12 0 3
rlabel polysilicon 205 -6 205 -6 0 1
rlabel polysilicon 208 -12 208 -12 0 4
rlabel polysilicon 338 -6 338 -6 0 1
rlabel polysilicon 341 -6 341 -6 0 2
rlabel polysilicon 341 -12 341 -12 0 4
rlabel polysilicon 345 -6 345 -6 0 1
rlabel polysilicon 345 -12 345 -12 0 3
rlabel polysilicon 352 -6 352 -6 0 1
rlabel polysilicon 352 -12 352 -12 0 3
rlabel polysilicon 359 -6 359 -6 0 1
rlabel polysilicon 359 -12 359 -12 0 3
rlabel polysilicon 366 -6 366 -6 0 1
rlabel polysilicon 366 -12 366 -12 0 3
rlabel polysilicon 376 -6 376 -6 0 2
rlabel polysilicon 373 -12 373 -12 0 3
rlabel polysilicon 394 -6 394 -6 0 1
rlabel polysilicon 394 -12 394 -12 0 3
rlabel polysilicon 401 -12 401 -12 0 3
rlabel polysilicon 404 -12 404 -12 0 4
rlabel polysilicon 408 -6 408 -6 0 1
rlabel polysilicon 411 -6 411 -6 0 2
rlabel polysilicon 432 -6 432 -6 0 2
rlabel polysilicon 429 -12 429 -12 0 3
rlabel polysilicon 432 -12 432 -12 0 4
rlabel polysilicon 436 -12 436 -12 0 3
rlabel polysilicon 439 -12 439 -12 0 4
rlabel polysilicon 450 -6 450 -6 0 1
rlabel polysilicon 450 -12 450 -12 0 3
rlabel polysilicon 464 -6 464 -6 0 1
rlabel polysilicon 464 -12 464 -12 0 3
rlabel polysilicon 471 -6 471 -6 0 1
rlabel polysilicon 474 -12 474 -12 0 4
rlabel polysilicon 481 -6 481 -6 0 2
rlabel polysilicon 478 -12 478 -12 0 3
rlabel polysilicon 492 -6 492 -6 0 1
rlabel polysilicon 492 -12 492 -12 0 3
rlabel polysilicon 513 -6 513 -6 0 1
rlabel polysilicon 513 -12 513 -12 0 3
rlabel polysilicon 576 -6 576 -6 0 1
rlabel polysilicon 576 -12 576 -12 0 3
rlabel polysilicon 128 -37 128 -37 0 1
rlabel polysilicon 128 -43 128 -43 0 3
rlabel polysilicon 198 -37 198 -37 0 1
rlabel polysilicon 198 -43 198 -43 0 3
rlabel polysilicon 219 -37 219 -37 0 1
rlabel polysilicon 219 -43 219 -43 0 3
rlabel polysilicon 243 -37 243 -37 0 2
rlabel polysilicon 240 -43 240 -43 0 3
rlabel polysilicon 243 -43 243 -43 0 4
rlabel polysilicon 254 -37 254 -37 0 1
rlabel polysilicon 254 -43 254 -43 0 3
rlabel polysilicon 282 -37 282 -37 0 1
rlabel polysilicon 282 -43 282 -43 0 3
rlabel polysilicon 289 -37 289 -37 0 1
rlabel polysilicon 292 -37 292 -37 0 2
rlabel polysilicon 289 -43 289 -43 0 3
rlabel polysilicon 296 -37 296 -37 0 1
rlabel polysilicon 296 -43 296 -43 0 3
rlabel polysilicon 303 -37 303 -37 0 1
rlabel polysilicon 303 -43 303 -43 0 3
rlabel polysilicon 310 -37 310 -37 0 1
rlabel polysilicon 310 -43 310 -43 0 3
rlabel polysilicon 320 -37 320 -37 0 2
rlabel polysilicon 320 -43 320 -43 0 4
rlabel polysilicon 324 -37 324 -37 0 1
rlabel polysilicon 327 -37 327 -37 0 2
rlabel polysilicon 324 -43 324 -43 0 3
rlabel polysilicon 331 -37 331 -37 0 1
rlabel polysilicon 331 -43 331 -43 0 3
rlabel polysilicon 338 -37 338 -37 0 1
rlabel polysilicon 338 -43 338 -43 0 3
rlabel polysilicon 345 -37 345 -37 0 1
rlabel polysilicon 345 -43 345 -43 0 3
rlabel polysilicon 352 -37 352 -37 0 1
rlabel polysilicon 352 -43 352 -43 0 3
rlabel polysilicon 359 -37 359 -37 0 1
rlabel polysilicon 359 -43 359 -43 0 3
rlabel polysilicon 366 -37 366 -37 0 1
rlabel polysilicon 366 -43 366 -43 0 3
rlabel polysilicon 373 -37 373 -37 0 1
rlabel polysilicon 376 -37 376 -37 0 2
rlabel polysilicon 373 -43 373 -43 0 3
rlabel polysilicon 380 -37 380 -37 0 1
rlabel polysilicon 380 -43 380 -43 0 3
rlabel polysilicon 387 -37 387 -37 0 1
rlabel polysilicon 387 -43 387 -43 0 3
rlabel polysilicon 394 -37 394 -37 0 1
rlabel polysilicon 394 -43 394 -43 0 3
rlabel polysilicon 397 -43 397 -43 0 4
rlabel polysilicon 401 -37 401 -37 0 1
rlabel polysilicon 401 -43 401 -43 0 3
rlabel polysilicon 408 -37 408 -37 0 1
rlabel polysilicon 408 -43 408 -43 0 3
rlabel polysilicon 415 -37 415 -37 0 1
rlabel polysilicon 415 -43 415 -43 0 3
rlabel polysilicon 422 -37 422 -37 0 1
rlabel polysilicon 422 -43 422 -43 0 3
rlabel polysilicon 432 -37 432 -37 0 2
rlabel polysilicon 432 -43 432 -43 0 4
rlabel polysilicon 436 -37 436 -37 0 1
rlabel polysilicon 436 -43 436 -43 0 3
rlabel polysilicon 446 -37 446 -37 0 2
rlabel polysilicon 443 -43 443 -43 0 3
rlabel polysilicon 446 -43 446 -43 0 4
rlabel polysilicon 450 -37 450 -37 0 1
rlabel polysilicon 450 -43 450 -43 0 3
rlabel polysilicon 457 -37 457 -37 0 1
rlabel polysilicon 457 -43 457 -43 0 3
rlabel polysilicon 464 -37 464 -37 0 1
rlabel polysilicon 464 -43 464 -43 0 3
rlabel polysilicon 471 -37 471 -37 0 1
rlabel polysilicon 471 -43 471 -43 0 3
rlabel polysilicon 478 -37 478 -37 0 1
rlabel polysilicon 478 -43 478 -43 0 3
rlabel polysilicon 485 -37 485 -37 0 1
rlabel polysilicon 485 -43 485 -43 0 3
rlabel polysilicon 492 -43 492 -43 0 3
rlabel polysilicon 495 -43 495 -43 0 4
rlabel polysilicon 502 -37 502 -37 0 2
rlabel polysilicon 499 -43 499 -43 0 3
rlabel polysilicon 502 -43 502 -43 0 4
rlabel polysilicon 506 -37 506 -37 0 1
rlabel polysilicon 506 -43 506 -43 0 3
rlabel polysilicon 513 -37 513 -37 0 1
rlabel polysilicon 513 -43 513 -43 0 3
rlabel polysilicon 527 -37 527 -37 0 1
rlabel polysilicon 527 -43 527 -43 0 3
rlabel polysilicon 534 -37 534 -37 0 1
rlabel polysilicon 534 -43 534 -43 0 3
rlabel polysilicon 541 -37 541 -37 0 1
rlabel polysilicon 541 -43 541 -43 0 3
rlabel polysilicon 548 -37 548 -37 0 1
rlabel polysilicon 548 -43 548 -43 0 3
rlabel polysilicon 593 -37 593 -37 0 2
rlabel polysilicon 590 -43 590 -43 0 3
rlabel polysilicon 593 -43 593 -43 0 4
rlabel polysilicon 618 -37 618 -37 0 1
rlabel polysilicon 618 -43 618 -43 0 3
rlabel polysilicon 625 -37 625 -37 0 1
rlabel polysilicon 625 -43 625 -43 0 3
rlabel polysilicon 114 -90 114 -90 0 1
rlabel polysilicon 114 -96 114 -96 0 3
rlabel polysilicon 117 -96 117 -96 0 4
rlabel polysilicon 142 -90 142 -90 0 1
rlabel polysilicon 142 -96 142 -96 0 3
rlabel polysilicon 163 -90 163 -90 0 1
rlabel polysilicon 163 -96 163 -96 0 3
rlabel polysilicon 170 -90 170 -90 0 1
rlabel polysilicon 170 -96 170 -96 0 3
rlabel polysilicon 177 -90 177 -90 0 1
rlabel polysilicon 177 -96 177 -96 0 3
rlabel polysilicon 184 -90 184 -90 0 1
rlabel polysilicon 184 -96 184 -96 0 3
rlabel polysilicon 191 -90 191 -90 0 1
rlabel polysilicon 191 -96 191 -96 0 3
rlabel polysilicon 198 -90 198 -90 0 1
rlabel polysilicon 198 -96 198 -96 0 3
rlabel polysilicon 205 -90 205 -90 0 1
rlabel polysilicon 205 -96 205 -96 0 3
rlabel polysilicon 212 -90 212 -90 0 1
rlabel polysilicon 212 -96 212 -96 0 3
rlabel polysilicon 219 -90 219 -90 0 1
rlabel polysilicon 219 -96 219 -96 0 3
rlabel polysilicon 226 -90 226 -90 0 1
rlabel polysilicon 226 -96 226 -96 0 3
rlabel polysilicon 233 -90 233 -90 0 1
rlabel polysilicon 233 -96 233 -96 0 3
rlabel polysilicon 240 -90 240 -90 0 1
rlabel polysilicon 240 -96 240 -96 0 3
rlabel polysilicon 247 -90 247 -90 0 1
rlabel polysilicon 247 -96 247 -96 0 3
rlabel polysilicon 254 -90 254 -90 0 1
rlabel polysilicon 254 -96 254 -96 0 3
rlabel polysilicon 261 -90 261 -90 0 1
rlabel polysilicon 261 -96 261 -96 0 3
rlabel polysilicon 268 -90 268 -90 0 1
rlabel polysilicon 268 -96 268 -96 0 3
rlabel polysilicon 275 -90 275 -90 0 1
rlabel polysilicon 275 -96 275 -96 0 3
rlabel polysilicon 278 -96 278 -96 0 4
rlabel polysilicon 282 -90 282 -90 0 1
rlabel polysilicon 282 -96 282 -96 0 3
rlabel polysilicon 289 -90 289 -90 0 1
rlabel polysilicon 289 -96 289 -96 0 3
rlabel polysilicon 296 -90 296 -90 0 1
rlabel polysilicon 296 -96 296 -96 0 3
rlabel polysilicon 303 -90 303 -90 0 1
rlabel polysilicon 303 -96 303 -96 0 3
rlabel polysilicon 310 -90 310 -90 0 1
rlabel polysilicon 310 -96 310 -96 0 3
rlabel polysilicon 317 -90 317 -90 0 1
rlabel polysilicon 317 -96 317 -96 0 3
rlabel polysilicon 324 -90 324 -90 0 1
rlabel polysilicon 324 -96 324 -96 0 3
rlabel polysilicon 334 -90 334 -90 0 2
rlabel polysilicon 331 -96 331 -96 0 3
rlabel polysilicon 334 -96 334 -96 0 4
rlabel polysilicon 338 -90 338 -90 0 1
rlabel polysilicon 338 -96 338 -96 0 3
rlabel polysilicon 345 -90 345 -90 0 1
rlabel polysilicon 348 -90 348 -90 0 2
rlabel polysilicon 345 -96 345 -96 0 3
rlabel polysilicon 352 -90 352 -90 0 1
rlabel polysilicon 352 -96 352 -96 0 3
rlabel polysilicon 359 -90 359 -90 0 1
rlabel polysilicon 359 -96 359 -96 0 3
rlabel polysilicon 366 -90 366 -90 0 1
rlabel polysilicon 369 -90 369 -90 0 2
rlabel polysilicon 369 -96 369 -96 0 4
rlabel polysilicon 373 -90 373 -90 0 1
rlabel polysilicon 373 -96 373 -96 0 3
rlabel polysilicon 376 -96 376 -96 0 4
rlabel polysilicon 380 -90 380 -90 0 1
rlabel polysilicon 380 -96 380 -96 0 3
rlabel polysilicon 383 -96 383 -96 0 4
rlabel polysilicon 387 -90 387 -90 0 1
rlabel polysilicon 390 -90 390 -90 0 2
rlabel polysilicon 387 -96 387 -96 0 3
rlabel polysilicon 397 -90 397 -90 0 2
rlabel polysilicon 394 -96 394 -96 0 3
rlabel polysilicon 401 -90 401 -90 0 1
rlabel polysilicon 401 -96 401 -96 0 3
rlabel polysilicon 408 -90 408 -90 0 1
rlabel polysilicon 408 -96 408 -96 0 3
rlabel polysilicon 415 -90 415 -90 0 1
rlabel polysilicon 415 -96 415 -96 0 3
rlabel polysilicon 422 -90 422 -90 0 1
rlabel polysilicon 422 -96 422 -96 0 3
rlabel polysilicon 429 -90 429 -90 0 1
rlabel polysilicon 429 -96 429 -96 0 3
rlabel polysilicon 436 -90 436 -90 0 1
rlabel polysilicon 436 -96 436 -96 0 3
rlabel polysilicon 443 -90 443 -90 0 1
rlabel polysilicon 443 -96 443 -96 0 3
rlabel polysilicon 450 -90 450 -90 0 1
rlabel polysilicon 450 -96 450 -96 0 3
rlabel polysilicon 453 -96 453 -96 0 4
rlabel polysilicon 457 -90 457 -90 0 1
rlabel polysilicon 457 -96 457 -96 0 3
rlabel polysilicon 464 -90 464 -90 0 1
rlabel polysilicon 464 -96 464 -96 0 3
rlabel polysilicon 474 -90 474 -90 0 2
rlabel polysilicon 471 -96 471 -96 0 3
rlabel polysilicon 474 -96 474 -96 0 4
rlabel polysilicon 478 -90 478 -90 0 1
rlabel polysilicon 481 -90 481 -90 0 2
rlabel polysilicon 481 -96 481 -96 0 4
rlabel polysilicon 485 -90 485 -90 0 1
rlabel polysilicon 485 -96 485 -96 0 3
rlabel polysilicon 492 -90 492 -90 0 1
rlabel polysilicon 492 -96 492 -96 0 3
rlabel polysilicon 499 -90 499 -90 0 1
rlabel polysilicon 499 -96 499 -96 0 3
rlabel polysilicon 506 -90 506 -90 0 1
rlabel polysilicon 506 -96 506 -96 0 3
rlabel polysilicon 513 -90 513 -90 0 1
rlabel polysilicon 513 -96 513 -96 0 3
rlabel polysilicon 520 -90 520 -90 0 1
rlabel polysilicon 520 -96 520 -96 0 3
rlabel polysilicon 527 -90 527 -90 0 1
rlabel polysilicon 527 -96 527 -96 0 3
rlabel polysilicon 534 -90 534 -90 0 1
rlabel polysilicon 534 -96 534 -96 0 3
rlabel polysilicon 541 -90 541 -90 0 1
rlabel polysilicon 541 -96 541 -96 0 3
rlabel polysilicon 548 -90 548 -90 0 1
rlabel polysilicon 548 -96 548 -96 0 3
rlabel polysilicon 555 -90 555 -90 0 1
rlabel polysilicon 555 -96 555 -96 0 3
rlabel polysilicon 562 -90 562 -90 0 1
rlabel polysilicon 562 -96 562 -96 0 3
rlabel polysilicon 569 -90 569 -90 0 1
rlabel polysilicon 569 -96 569 -96 0 3
rlabel polysilicon 576 -90 576 -90 0 1
rlabel polysilicon 576 -96 576 -96 0 3
rlabel polysilicon 583 -90 583 -90 0 1
rlabel polysilicon 583 -96 583 -96 0 3
rlabel polysilicon 590 -90 590 -90 0 1
rlabel polysilicon 593 -90 593 -90 0 2
rlabel polysilicon 593 -96 593 -96 0 4
rlabel polysilicon 597 -90 597 -90 0 1
rlabel polysilicon 597 -96 597 -96 0 3
rlabel polysilicon 604 -90 604 -90 0 1
rlabel polysilicon 604 -96 604 -96 0 3
rlabel polysilicon 611 -90 611 -90 0 1
rlabel polysilicon 611 -96 611 -96 0 3
rlabel polysilicon 618 -90 618 -90 0 1
rlabel polysilicon 618 -96 618 -96 0 3
rlabel polysilicon 625 -90 625 -90 0 1
rlabel polysilicon 625 -96 625 -96 0 3
rlabel polysilicon 632 -90 632 -90 0 1
rlabel polysilicon 632 -96 632 -96 0 3
rlabel polysilicon 639 -90 639 -90 0 1
rlabel polysilicon 639 -96 639 -96 0 3
rlabel polysilicon 646 -90 646 -90 0 1
rlabel polysilicon 646 -96 646 -96 0 3
rlabel polysilicon 653 -90 653 -90 0 1
rlabel polysilicon 653 -96 653 -96 0 3
rlabel polysilicon 660 -90 660 -90 0 1
rlabel polysilicon 660 -96 660 -96 0 3
rlabel polysilicon 667 -90 667 -90 0 1
rlabel polysilicon 667 -96 667 -96 0 3
rlabel polysilicon 674 -90 674 -90 0 1
rlabel polysilicon 674 -96 674 -96 0 3
rlabel polysilicon 681 -90 681 -90 0 1
rlabel polysilicon 681 -96 681 -96 0 3
rlabel polysilicon 688 -90 688 -90 0 1
rlabel polysilicon 691 -90 691 -90 0 2
rlabel polysilicon 688 -96 688 -96 0 3
rlabel polysilicon 51 -157 51 -157 0 1
rlabel polysilicon 51 -163 51 -163 0 3
rlabel polysilicon 58 -157 58 -157 0 1
rlabel polysilicon 58 -163 58 -163 0 3
rlabel polysilicon 65 -157 65 -157 0 1
rlabel polysilicon 65 -163 65 -163 0 3
rlabel polysilicon 72 -157 72 -157 0 1
rlabel polysilicon 72 -163 72 -163 0 3
rlabel polysilicon 82 -157 82 -157 0 2
rlabel polysilicon 86 -157 86 -157 0 1
rlabel polysilicon 86 -163 86 -163 0 3
rlabel polysilicon 93 -157 93 -157 0 1
rlabel polysilicon 93 -163 93 -163 0 3
rlabel polysilicon 100 -157 100 -157 0 1
rlabel polysilicon 100 -163 100 -163 0 3
rlabel polysilicon 103 -163 103 -163 0 4
rlabel polysilicon 107 -157 107 -157 0 1
rlabel polysilicon 107 -163 107 -163 0 3
rlabel polysilicon 114 -157 114 -157 0 1
rlabel polysilicon 114 -163 114 -163 0 3
rlabel polysilicon 121 -157 121 -157 0 1
rlabel polysilicon 121 -163 121 -163 0 3
rlabel polysilicon 128 -157 128 -157 0 1
rlabel polysilicon 128 -163 128 -163 0 3
rlabel polysilicon 135 -157 135 -157 0 1
rlabel polysilicon 135 -163 135 -163 0 3
rlabel polysilicon 145 -157 145 -157 0 2
rlabel polysilicon 142 -163 142 -163 0 3
rlabel polysilicon 145 -163 145 -163 0 4
rlabel polysilicon 152 -157 152 -157 0 2
rlabel polysilicon 149 -163 149 -163 0 3
rlabel polysilicon 152 -163 152 -163 0 4
rlabel polysilicon 156 -157 156 -157 0 1
rlabel polysilicon 156 -163 156 -163 0 3
rlabel polysilicon 163 -157 163 -157 0 1
rlabel polysilicon 163 -163 163 -163 0 3
rlabel polysilicon 170 -157 170 -157 0 1
rlabel polysilicon 170 -163 170 -163 0 3
rlabel polysilicon 177 -157 177 -157 0 1
rlabel polysilicon 177 -163 177 -163 0 3
rlabel polysilicon 184 -157 184 -157 0 1
rlabel polysilicon 187 -157 187 -157 0 2
rlabel polysilicon 184 -163 184 -163 0 3
rlabel polysilicon 194 -157 194 -157 0 2
rlabel polysilicon 191 -163 191 -163 0 3
rlabel polysilicon 194 -163 194 -163 0 4
rlabel polysilicon 198 -157 198 -157 0 1
rlabel polysilicon 201 -157 201 -157 0 2
rlabel polysilicon 201 -163 201 -163 0 4
rlabel polysilicon 205 -157 205 -157 0 1
rlabel polysilicon 205 -163 205 -163 0 3
rlabel polysilicon 212 -157 212 -157 0 1
rlabel polysilicon 212 -163 212 -163 0 3
rlabel polysilicon 219 -157 219 -157 0 1
rlabel polysilicon 219 -163 219 -163 0 3
rlabel polysilicon 226 -157 226 -157 0 1
rlabel polysilicon 226 -163 226 -163 0 3
rlabel polysilicon 233 -157 233 -157 0 1
rlabel polysilicon 233 -163 233 -163 0 3
rlabel polysilicon 240 -157 240 -157 0 1
rlabel polysilicon 240 -163 240 -163 0 3
rlabel polysilicon 247 -157 247 -157 0 1
rlabel polysilicon 247 -163 247 -163 0 3
rlabel polysilicon 254 -157 254 -157 0 1
rlabel polysilicon 254 -163 254 -163 0 3
rlabel polysilicon 261 -157 261 -157 0 1
rlabel polysilicon 261 -163 261 -163 0 3
rlabel polysilicon 268 -157 268 -157 0 1
rlabel polysilicon 268 -163 268 -163 0 3
rlabel polysilicon 275 -157 275 -157 0 1
rlabel polysilicon 275 -163 275 -163 0 3
rlabel polysilicon 282 -157 282 -157 0 1
rlabel polysilicon 282 -163 282 -163 0 3
rlabel polysilicon 289 -157 289 -157 0 1
rlabel polysilicon 289 -163 289 -163 0 3
rlabel polysilicon 296 -157 296 -157 0 1
rlabel polysilicon 296 -163 296 -163 0 3
rlabel polysilicon 303 -157 303 -157 0 1
rlabel polysilicon 303 -163 303 -163 0 3
rlabel polysilicon 310 -157 310 -157 0 1
rlabel polysilicon 310 -163 310 -163 0 3
rlabel polysilicon 317 -157 317 -157 0 1
rlabel polysilicon 317 -163 317 -163 0 3
rlabel polysilicon 324 -157 324 -157 0 1
rlabel polysilicon 324 -163 324 -163 0 3
rlabel polysilicon 331 -157 331 -157 0 1
rlabel polysilicon 331 -163 331 -163 0 3
rlabel polysilicon 338 -157 338 -157 0 1
rlabel polysilicon 338 -163 338 -163 0 3
rlabel polysilicon 345 -157 345 -157 0 1
rlabel polysilicon 345 -163 345 -163 0 3
rlabel polysilicon 352 -157 352 -157 0 1
rlabel polysilicon 352 -163 352 -163 0 3
rlabel polysilicon 359 -157 359 -157 0 1
rlabel polysilicon 359 -163 359 -163 0 3
rlabel polysilicon 366 -157 366 -157 0 1
rlabel polysilicon 366 -163 366 -163 0 3
rlabel polysilicon 373 -157 373 -157 0 1
rlabel polysilicon 373 -163 373 -163 0 3
rlabel polysilicon 380 -157 380 -157 0 1
rlabel polysilicon 380 -163 380 -163 0 3
rlabel polysilicon 387 -157 387 -157 0 1
rlabel polysilicon 387 -163 387 -163 0 3
rlabel polysilicon 394 -157 394 -157 0 1
rlabel polysilicon 394 -163 394 -163 0 3
rlabel polysilicon 401 -157 401 -157 0 1
rlabel polysilicon 401 -163 401 -163 0 3
rlabel polysilicon 411 -157 411 -157 0 2
rlabel polysilicon 408 -163 408 -163 0 3
rlabel polysilicon 411 -163 411 -163 0 4
rlabel polysilicon 415 -157 415 -157 0 1
rlabel polysilicon 418 -157 418 -157 0 2
rlabel polysilicon 415 -163 415 -163 0 3
rlabel polysilicon 422 -157 422 -157 0 1
rlabel polysilicon 422 -163 422 -163 0 3
rlabel polysilicon 429 -157 429 -157 0 1
rlabel polysilicon 429 -163 429 -163 0 3
rlabel polysilicon 436 -157 436 -157 0 1
rlabel polysilicon 436 -163 436 -163 0 3
rlabel polysilicon 443 -157 443 -157 0 1
rlabel polysilicon 443 -163 443 -163 0 3
rlabel polysilicon 453 -157 453 -157 0 2
rlabel polysilicon 450 -163 450 -163 0 3
rlabel polysilicon 453 -163 453 -163 0 4
rlabel polysilicon 457 -157 457 -157 0 1
rlabel polysilicon 457 -163 457 -163 0 3
rlabel polysilicon 464 -157 464 -157 0 1
rlabel polysilicon 467 -157 467 -157 0 2
rlabel polysilicon 464 -163 464 -163 0 3
rlabel polysilicon 471 -157 471 -157 0 1
rlabel polysilicon 474 -157 474 -157 0 2
rlabel polysilicon 474 -163 474 -163 0 4
rlabel polysilicon 478 -157 478 -157 0 1
rlabel polysilicon 478 -163 478 -163 0 3
rlabel polysilicon 481 -163 481 -163 0 4
rlabel polysilicon 485 -157 485 -157 0 1
rlabel polysilicon 485 -163 485 -163 0 3
rlabel polysilicon 495 -157 495 -157 0 2
rlabel polysilicon 492 -163 492 -163 0 3
rlabel polysilicon 495 -163 495 -163 0 4
rlabel polysilicon 499 -157 499 -157 0 1
rlabel polysilicon 499 -163 499 -163 0 3
rlabel polysilicon 506 -157 506 -157 0 1
rlabel polysilicon 506 -163 506 -163 0 3
rlabel polysilicon 513 -157 513 -157 0 1
rlabel polysilicon 513 -163 513 -163 0 3
rlabel polysilicon 520 -157 520 -157 0 1
rlabel polysilicon 520 -163 520 -163 0 3
rlabel polysilicon 527 -157 527 -157 0 1
rlabel polysilicon 527 -163 527 -163 0 3
rlabel polysilicon 534 -157 534 -157 0 1
rlabel polysilicon 534 -163 534 -163 0 3
rlabel polysilicon 541 -157 541 -157 0 1
rlabel polysilicon 541 -163 541 -163 0 3
rlabel polysilicon 548 -157 548 -157 0 1
rlabel polysilicon 548 -163 548 -163 0 3
rlabel polysilicon 555 -157 555 -157 0 1
rlabel polysilicon 555 -163 555 -163 0 3
rlabel polysilicon 562 -157 562 -157 0 1
rlabel polysilicon 562 -163 562 -163 0 3
rlabel polysilicon 569 -157 569 -157 0 1
rlabel polysilicon 569 -163 569 -163 0 3
rlabel polysilicon 576 -157 576 -157 0 1
rlabel polysilicon 579 -157 579 -157 0 2
rlabel polysilicon 576 -163 576 -163 0 3
rlabel polysilicon 583 -157 583 -157 0 1
rlabel polysilicon 583 -163 583 -163 0 3
rlabel polysilicon 590 -157 590 -157 0 1
rlabel polysilicon 590 -163 590 -163 0 3
rlabel polysilicon 597 -157 597 -157 0 1
rlabel polysilicon 597 -163 597 -163 0 3
rlabel polysilicon 604 -157 604 -157 0 1
rlabel polysilicon 604 -163 604 -163 0 3
rlabel polysilicon 611 -157 611 -157 0 1
rlabel polysilicon 611 -163 611 -163 0 3
rlabel polysilicon 618 -157 618 -157 0 1
rlabel polysilicon 618 -163 618 -163 0 3
rlabel polysilicon 625 -157 625 -157 0 1
rlabel polysilicon 625 -163 625 -163 0 3
rlabel polysilicon 632 -157 632 -157 0 1
rlabel polysilicon 632 -163 632 -163 0 3
rlabel polysilicon 639 -157 639 -157 0 1
rlabel polysilicon 639 -163 639 -163 0 3
rlabel polysilicon 646 -157 646 -157 0 1
rlabel polysilicon 646 -163 646 -163 0 3
rlabel polysilicon 653 -157 653 -157 0 1
rlabel polysilicon 653 -163 653 -163 0 3
rlabel polysilicon 660 -157 660 -157 0 1
rlabel polysilicon 660 -163 660 -163 0 3
rlabel polysilicon 667 -157 667 -157 0 1
rlabel polysilicon 667 -163 667 -163 0 3
rlabel polysilicon 674 -157 674 -157 0 1
rlabel polysilicon 674 -163 674 -163 0 3
rlabel polysilicon 681 -157 681 -157 0 1
rlabel polysilicon 681 -163 681 -163 0 3
rlabel polysilicon 688 -157 688 -157 0 1
rlabel polysilicon 688 -163 688 -163 0 3
rlabel polysilicon 695 -157 695 -157 0 1
rlabel polysilicon 695 -163 695 -163 0 3
rlabel polysilicon 702 -157 702 -157 0 1
rlabel polysilicon 702 -163 702 -163 0 3
rlabel polysilicon 709 -157 709 -157 0 1
rlabel polysilicon 709 -163 709 -163 0 3
rlabel polysilicon 716 -157 716 -157 0 1
rlabel polysilicon 716 -163 716 -163 0 3
rlabel polysilicon 723 -157 723 -157 0 1
rlabel polysilicon 723 -163 723 -163 0 3
rlabel polysilicon 730 -157 730 -157 0 1
rlabel polysilicon 730 -163 730 -163 0 3
rlabel polysilicon 737 -157 737 -157 0 1
rlabel polysilicon 737 -163 737 -163 0 3
rlabel polysilicon 744 -157 744 -157 0 1
rlabel polysilicon 744 -163 744 -163 0 3
rlabel polysilicon 751 -157 751 -157 0 1
rlabel polysilicon 751 -163 751 -163 0 3
rlabel polysilicon 758 -157 758 -157 0 1
rlabel polysilicon 758 -163 758 -163 0 3
rlabel polysilicon 765 -157 765 -157 0 1
rlabel polysilicon 765 -163 765 -163 0 3
rlabel polysilicon 772 -157 772 -157 0 1
rlabel polysilicon 772 -163 772 -163 0 3
rlabel polysilicon 779 -157 779 -157 0 1
rlabel polysilicon 779 -163 779 -163 0 3
rlabel polysilicon 786 -157 786 -157 0 1
rlabel polysilicon 786 -163 786 -163 0 3
rlabel polysilicon 793 -157 793 -157 0 1
rlabel polysilicon 793 -163 793 -163 0 3
rlabel polysilicon 800 -157 800 -157 0 1
rlabel polysilicon 800 -163 800 -163 0 3
rlabel polysilicon 807 -157 807 -157 0 1
rlabel polysilicon 807 -163 807 -163 0 3
rlabel polysilicon 814 -157 814 -157 0 1
rlabel polysilicon 814 -163 814 -163 0 3
rlabel polysilicon 821 -157 821 -157 0 1
rlabel polysilicon 821 -163 821 -163 0 3
rlabel polysilicon 44 -238 44 -238 0 1
rlabel polysilicon 44 -244 44 -244 0 3
rlabel polysilicon 51 -238 51 -238 0 1
rlabel polysilicon 51 -244 51 -244 0 3
rlabel polysilicon 58 -238 58 -238 0 1
rlabel polysilicon 58 -244 58 -244 0 3
rlabel polysilicon 65 -238 65 -238 0 1
rlabel polysilicon 65 -244 65 -244 0 3
rlabel polysilicon 72 -238 72 -238 0 1
rlabel polysilicon 72 -244 72 -244 0 3
rlabel polysilicon 79 -238 79 -238 0 1
rlabel polysilicon 79 -244 79 -244 0 3
rlabel polysilicon 86 -238 86 -238 0 1
rlabel polysilicon 86 -244 86 -244 0 3
rlabel polysilicon 93 -238 93 -238 0 1
rlabel polysilicon 93 -244 93 -244 0 3
rlabel polysilicon 100 -244 100 -244 0 3
rlabel polysilicon 103 -244 103 -244 0 4
rlabel polysilicon 107 -238 107 -238 0 1
rlabel polysilicon 107 -244 107 -244 0 3
rlabel polysilicon 117 -238 117 -238 0 2
rlabel polysilicon 114 -244 114 -244 0 3
rlabel polysilicon 117 -244 117 -244 0 4
rlabel polysilicon 121 -238 121 -238 0 1
rlabel polysilicon 124 -238 124 -238 0 2
rlabel polysilicon 121 -244 121 -244 0 3
rlabel polysilicon 124 -244 124 -244 0 4
rlabel polysilicon 128 -238 128 -238 0 1
rlabel polysilicon 128 -244 128 -244 0 3
rlabel polysilicon 135 -238 135 -238 0 1
rlabel polysilicon 138 -238 138 -238 0 2
rlabel polysilicon 135 -244 135 -244 0 3
rlabel polysilicon 142 -238 142 -238 0 1
rlabel polysilicon 142 -244 142 -244 0 3
rlabel polysilicon 149 -238 149 -238 0 1
rlabel polysilicon 149 -244 149 -244 0 3
rlabel polysilicon 156 -238 156 -238 0 1
rlabel polysilicon 156 -244 156 -244 0 3
rlabel polysilicon 163 -238 163 -238 0 1
rlabel polysilicon 166 -238 166 -238 0 2
rlabel polysilicon 163 -244 163 -244 0 3
rlabel polysilicon 166 -244 166 -244 0 4
rlabel polysilicon 170 -238 170 -238 0 1
rlabel polysilicon 170 -244 170 -244 0 3
rlabel polysilicon 177 -238 177 -238 0 1
rlabel polysilicon 177 -244 177 -244 0 3
rlabel polysilicon 184 -238 184 -238 0 1
rlabel polysilicon 184 -244 184 -244 0 3
rlabel polysilicon 191 -238 191 -238 0 1
rlabel polysilicon 191 -244 191 -244 0 3
rlabel polysilicon 198 -238 198 -238 0 1
rlabel polysilicon 198 -244 198 -244 0 3
rlabel polysilicon 205 -238 205 -238 0 1
rlabel polysilicon 205 -244 205 -244 0 3
rlabel polysilicon 212 -238 212 -238 0 1
rlabel polysilicon 212 -244 212 -244 0 3
rlabel polysilicon 219 -238 219 -238 0 1
rlabel polysilicon 219 -244 219 -244 0 3
rlabel polysilicon 226 -238 226 -238 0 1
rlabel polysilicon 226 -244 226 -244 0 3
rlabel polysilicon 233 -238 233 -238 0 1
rlabel polysilicon 233 -244 233 -244 0 3
rlabel polysilicon 240 -238 240 -238 0 1
rlabel polysilicon 240 -244 240 -244 0 3
rlabel polysilicon 247 -238 247 -238 0 1
rlabel polysilicon 247 -244 247 -244 0 3
rlabel polysilicon 254 -238 254 -238 0 1
rlabel polysilicon 257 -238 257 -238 0 2
rlabel polysilicon 254 -244 254 -244 0 3
rlabel polysilicon 257 -244 257 -244 0 4
rlabel polysilicon 261 -238 261 -238 0 1
rlabel polysilicon 261 -244 261 -244 0 3
rlabel polysilicon 268 -238 268 -238 0 1
rlabel polysilicon 268 -244 268 -244 0 3
rlabel polysilicon 275 -238 275 -238 0 1
rlabel polysilicon 275 -244 275 -244 0 3
rlabel polysilicon 282 -238 282 -238 0 1
rlabel polysilicon 285 -238 285 -238 0 2
rlabel polysilicon 282 -244 282 -244 0 3
rlabel polysilicon 285 -244 285 -244 0 4
rlabel polysilicon 289 -238 289 -238 0 1
rlabel polysilicon 292 -238 292 -238 0 2
rlabel polysilicon 289 -244 289 -244 0 3
rlabel polysilicon 292 -244 292 -244 0 4
rlabel polysilicon 296 -238 296 -238 0 1
rlabel polysilicon 296 -244 296 -244 0 3
rlabel polysilicon 303 -238 303 -238 0 1
rlabel polysilicon 303 -244 303 -244 0 3
rlabel polysilicon 310 -238 310 -238 0 1
rlabel polysilicon 310 -244 310 -244 0 3
rlabel polysilicon 317 -238 317 -238 0 1
rlabel polysilicon 317 -244 317 -244 0 3
rlabel polysilicon 324 -238 324 -238 0 1
rlabel polysilicon 324 -244 324 -244 0 3
rlabel polysilicon 331 -238 331 -238 0 1
rlabel polysilicon 331 -244 331 -244 0 3
rlabel polysilicon 338 -238 338 -238 0 1
rlabel polysilicon 338 -244 338 -244 0 3
rlabel polysilicon 345 -238 345 -238 0 1
rlabel polysilicon 348 -238 348 -238 0 2
rlabel polysilicon 345 -244 345 -244 0 3
rlabel polysilicon 348 -244 348 -244 0 4
rlabel polysilicon 352 -238 352 -238 0 1
rlabel polysilicon 355 -238 355 -238 0 2
rlabel polysilicon 352 -244 352 -244 0 3
rlabel polysilicon 355 -244 355 -244 0 4
rlabel polysilicon 359 -238 359 -238 0 1
rlabel polysilicon 362 -238 362 -238 0 2
rlabel polysilicon 359 -244 359 -244 0 3
rlabel polysilicon 362 -244 362 -244 0 4
rlabel polysilicon 366 -238 366 -238 0 1
rlabel polysilicon 366 -244 366 -244 0 3
rlabel polysilicon 376 -238 376 -238 0 2
rlabel polysilicon 376 -244 376 -244 0 4
rlabel polysilicon 380 -238 380 -238 0 1
rlabel polysilicon 380 -244 380 -244 0 3
rlabel polysilicon 387 -238 387 -238 0 1
rlabel polysilicon 387 -244 387 -244 0 3
rlabel polysilicon 394 -238 394 -238 0 1
rlabel polysilicon 394 -244 394 -244 0 3
rlabel polysilicon 401 -238 401 -238 0 1
rlabel polysilicon 404 -238 404 -238 0 2
rlabel polysilicon 401 -244 401 -244 0 3
rlabel polysilicon 408 -238 408 -238 0 1
rlabel polysilicon 408 -244 408 -244 0 3
rlabel polysilicon 415 -238 415 -238 0 1
rlabel polysilicon 415 -244 415 -244 0 3
rlabel polysilicon 422 -238 422 -238 0 1
rlabel polysilicon 425 -238 425 -238 0 2
rlabel polysilicon 422 -244 422 -244 0 3
rlabel polysilicon 425 -244 425 -244 0 4
rlabel polysilicon 429 -238 429 -238 0 1
rlabel polysilicon 429 -244 429 -244 0 3
rlabel polysilicon 436 -238 436 -238 0 1
rlabel polysilicon 439 -238 439 -238 0 2
rlabel polysilicon 436 -244 436 -244 0 3
rlabel polysilicon 443 -238 443 -238 0 1
rlabel polysilicon 443 -244 443 -244 0 3
rlabel polysilicon 450 -238 450 -238 0 1
rlabel polysilicon 450 -244 450 -244 0 3
rlabel polysilicon 457 -238 457 -238 0 1
rlabel polysilicon 460 -238 460 -238 0 2
rlabel polysilicon 457 -244 457 -244 0 3
rlabel polysilicon 464 -238 464 -238 0 1
rlabel polysilicon 464 -244 464 -244 0 3
rlabel polysilicon 471 -238 471 -238 0 1
rlabel polysilicon 474 -238 474 -238 0 2
rlabel polysilicon 474 -244 474 -244 0 4
rlabel polysilicon 478 -238 478 -238 0 1
rlabel polysilicon 478 -244 478 -244 0 3
rlabel polysilicon 485 -238 485 -238 0 1
rlabel polysilicon 485 -244 485 -244 0 3
rlabel polysilicon 492 -238 492 -238 0 1
rlabel polysilicon 495 -238 495 -238 0 2
rlabel polysilicon 492 -244 492 -244 0 3
rlabel polysilicon 495 -244 495 -244 0 4
rlabel polysilicon 499 -238 499 -238 0 1
rlabel polysilicon 499 -244 499 -244 0 3
rlabel polysilicon 506 -238 506 -238 0 1
rlabel polysilicon 506 -244 506 -244 0 3
rlabel polysilicon 513 -238 513 -238 0 1
rlabel polysilicon 513 -244 513 -244 0 3
rlabel polysilicon 520 -238 520 -238 0 1
rlabel polysilicon 520 -244 520 -244 0 3
rlabel polysilicon 527 -238 527 -238 0 1
rlabel polysilicon 534 -238 534 -238 0 1
rlabel polysilicon 534 -244 534 -244 0 3
rlabel polysilicon 541 -238 541 -238 0 1
rlabel polysilicon 541 -244 541 -244 0 3
rlabel polysilicon 548 -238 548 -238 0 1
rlabel polysilicon 548 -244 548 -244 0 3
rlabel polysilicon 555 -238 555 -238 0 1
rlabel polysilicon 555 -244 555 -244 0 3
rlabel polysilicon 562 -238 562 -238 0 1
rlabel polysilicon 562 -244 562 -244 0 3
rlabel polysilicon 569 -238 569 -238 0 1
rlabel polysilicon 569 -244 569 -244 0 3
rlabel polysilicon 576 -238 576 -238 0 1
rlabel polysilicon 576 -244 576 -244 0 3
rlabel polysilicon 579 -244 579 -244 0 4
rlabel polysilicon 583 -238 583 -238 0 1
rlabel polysilicon 583 -244 583 -244 0 3
rlabel polysilicon 590 -238 590 -238 0 1
rlabel polysilicon 590 -244 590 -244 0 3
rlabel polysilicon 597 -238 597 -238 0 1
rlabel polysilicon 597 -244 597 -244 0 3
rlabel polysilicon 604 -238 604 -238 0 1
rlabel polysilicon 604 -244 604 -244 0 3
rlabel polysilicon 611 -238 611 -238 0 1
rlabel polysilicon 611 -244 611 -244 0 3
rlabel polysilicon 618 -238 618 -238 0 1
rlabel polysilicon 618 -244 618 -244 0 3
rlabel polysilicon 625 -238 625 -238 0 1
rlabel polysilicon 625 -244 625 -244 0 3
rlabel polysilicon 632 -238 632 -238 0 1
rlabel polysilicon 632 -244 632 -244 0 3
rlabel polysilicon 639 -238 639 -238 0 1
rlabel polysilicon 639 -244 639 -244 0 3
rlabel polysilicon 646 -238 646 -238 0 1
rlabel polysilicon 646 -244 646 -244 0 3
rlabel polysilicon 653 -238 653 -238 0 1
rlabel polysilicon 653 -244 653 -244 0 3
rlabel polysilicon 660 -238 660 -238 0 1
rlabel polysilicon 660 -244 660 -244 0 3
rlabel polysilicon 667 -238 667 -238 0 1
rlabel polysilicon 667 -244 667 -244 0 3
rlabel polysilicon 674 -238 674 -238 0 1
rlabel polysilicon 674 -244 674 -244 0 3
rlabel polysilicon 681 -238 681 -238 0 1
rlabel polysilicon 681 -244 681 -244 0 3
rlabel polysilicon 688 -238 688 -238 0 1
rlabel polysilicon 688 -244 688 -244 0 3
rlabel polysilicon 695 -238 695 -238 0 1
rlabel polysilicon 695 -244 695 -244 0 3
rlabel polysilicon 702 -238 702 -238 0 1
rlabel polysilicon 702 -244 702 -244 0 3
rlabel polysilicon 709 -238 709 -238 0 1
rlabel polysilicon 709 -244 709 -244 0 3
rlabel polysilicon 716 -238 716 -238 0 1
rlabel polysilicon 716 -244 716 -244 0 3
rlabel polysilicon 723 -238 723 -238 0 1
rlabel polysilicon 723 -244 723 -244 0 3
rlabel polysilicon 730 -238 730 -238 0 1
rlabel polysilicon 730 -244 730 -244 0 3
rlabel polysilicon 737 -238 737 -238 0 1
rlabel polysilicon 737 -244 737 -244 0 3
rlabel polysilicon 744 -238 744 -238 0 1
rlabel polysilicon 744 -244 744 -244 0 3
rlabel polysilicon 751 -238 751 -238 0 1
rlabel polysilicon 751 -244 751 -244 0 3
rlabel polysilicon 758 -238 758 -238 0 1
rlabel polysilicon 758 -244 758 -244 0 3
rlabel polysilicon 765 -238 765 -238 0 1
rlabel polysilicon 765 -244 765 -244 0 3
rlabel polysilicon 772 -238 772 -238 0 1
rlabel polysilicon 772 -244 772 -244 0 3
rlabel polysilicon 779 -238 779 -238 0 1
rlabel polysilicon 779 -244 779 -244 0 3
rlabel polysilicon 786 -238 786 -238 0 1
rlabel polysilicon 786 -244 786 -244 0 3
rlabel polysilicon 793 -238 793 -238 0 1
rlabel polysilicon 793 -244 793 -244 0 3
rlabel polysilicon 800 -238 800 -238 0 1
rlabel polysilicon 800 -244 800 -244 0 3
rlabel polysilicon 807 -238 807 -238 0 1
rlabel polysilicon 807 -244 807 -244 0 3
rlabel polysilicon 814 -238 814 -238 0 1
rlabel polysilicon 814 -244 814 -244 0 3
rlabel polysilicon 821 -238 821 -238 0 1
rlabel polysilicon 821 -244 821 -244 0 3
rlabel polysilicon 828 -238 828 -238 0 1
rlabel polysilicon 828 -244 828 -244 0 3
rlabel polysilicon 835 -238 835 -238 0 1
rlabel polysilicon 835 -244 835 -244 0 3
rlabel polysilicon 842 -238 842 -238 0 1
rlabel polysilicon 842 -244 842 -244 0 3
rlabel polysilicon 849 -238 849 -238 0 1
rlabel polysilicon 849 -244 849 -244 0 3
rlabel polysilicon 859 -238 859 -238 0 2
rlabel polysilicon 863 -238 863 -238 0 1
rlabel polysilicon 863 -244 863 -244 0 3
rlabel polysilicon 2 -327 2 -327 0 1
rlabel polysilicon 2 -333 2 -333 0 3
rlabel polysilicon 9 -327 9 -327 0 1
rlabel polysilicon 9 -333 9 -333 0 3
rlabel polysilicon 16 -327 16 -327 0 1
rlabel polysilicon 16 -333 16 -333 0 3
rlabel polysilicon 23 -327 23 -327 0 1
rlabel polysilicon 23 -333 23 -333 0 3
rlabel polysilicon 30 -327 30 -327 0 1
rlabel polysilicon 30 -333 30 -333 0 3
rlabel polysilicon 37 -327 37 -327 0 1
rlabel polysilicon 37 -333 37 -333 0 3
rlabel polysilicon 44 -327 44 -327 0 1
rlabel polysilicon 44 -333 44 -333 0 3
rlabel polysilicon 51 -327 51 -327 0 1
rlabel polysilicon 51 -333 51 -333 0 3
rlabel polysilicon 58 -327 58 -327 0 1
rlabel polysilicon 58 -333 58 -333 0 3
rlabel polysilicon 65 -327 65 -327 0 1
rlabel polysilicon 68 -327 68 -327 0 2
rlabel polysilicon 68 -333 68 -333 0 4
rlabel polysilicon 72 -327 72 -327 0 1
rlabel polysilicon 72 -333 72 -333 0 3
rlabel polysilicon 79 -327 79 -327 0 1
rlabel polysilicon 79 -333 79 -333 0 3
rlabel polysilicon 86 -327 86 -327 0 1
rlabel polysilicon 86 -333 86 -333 0 3
rlabel polysilicon 93 -327 93 -327 0 1
rlabel polysilicon 93 -333 93 -333 0 3
rlabel polysilicon 100 -327 100 -327 0 1
rlabel polysilicon 100 -333 100 -333 0 3
rlabel polysilicon 107 -327 107 -327 0 1
rlabel polysilicon 107 -333 107 -333 0 3
rlabel polysilicon 114 -327 114 -327 0 1
rlabel polysilicon 114 -333 114 -333 0 3
rlabel polysilicon 121 -327 121 -327 0 1
rlabel polysilicon 121 -333 121 -333 0 3
rlabel polysilicon 128 -333 128 -333 0 3
rlabel polysilicon 131 -333 131 -333 0 4
rlabel polysilicon 135 -327 135 -327 0 1
rlabel polysilicon 135 -333 135 -333 0 3
rlabel polysilicon 142 -327 142 -327 0 1
rlabel polysilicon 142 -333 142 -333 0 3
rlabel polysilicon 149 -327 149 -327 0 1
rlabel polysilicon 149 -333 149 -333 0 3
rlabel polysilicon 156 -327 156 -327 0 1
rlabel polysilicon 156 -333 156 -333 0 3
rlabel polysilicon 163 -327 163 -327 0 1
rlabel polysilicon 163 -333 163 -333 0 3
rlabel polysilicon 170 -327 170 -327 0 1
rlabel polysilicon 170 -333 170 -333 0 3
rlabel polysilicon 177 -327 177 -327 0 1
rlabel polysilicon 177 -333 177 -333 0 3
rlabel polysilicon 184 -327 184 -327 0 1
rlabel polysilicon 184 -333 184 -333 0 3
rlabel polysilicon 191 -327 191 -327 0 1
rlabel polysilicon 198 -327 198 -327 0 1
rlabel polysilicon 198 -333 198 -333 0 3
rlabel polysilicon 205 -327 205 -327 0 1
rlabel polysilicon 205 -333 205 -333 0 3
rlabel polysilicon 212 -327 212 -327 0 1
rlabel polysilicon 212 -333 212 -333 0 3
rlabel polysilicon 219 -327 219 -327 0 1
rlabel polysilicon 219 -333 219 -333 0 3
rlabel polysilicon 226 -327 226 -327 0 1
rlabel polysilicon 226 -333 226 -333 0 3
rlabel polysilicon 233 -327 233 -327 0 1
rlabel polysilicon 233 -333 233 -333 0 3
rlabel polysilicon 240 -327 240 -327 0 1
rlabel polysilicon 240 -333 240 -333 0 3
rlabel polysilicon 247 -327 247 -327 0 1
rlabel polysilicon 247 -333 247 -333 0 3
rlabel polysilicon 254 -327 254 -327 0 1
rlabel polysilicon 254 -333 254 -333 0 3
rlabel polysilicon 261 -327 261 -327 0 1
rlabel polysilicon 261 -333 261 -333 0 3
rlabel polysilicon 268 -327 268 -327 0 1
rlabel polysilicon 268 -333 268 -333 0 3
rlabel polysilicon 275 -327 275 -327 0 1
rlabel polysilicon 275 -333 275 -333 0 3
rlabel polysilicon 282 -327 282 -327 0 1
rlabel polysilicon 282 -333 282 -333 0 3
rlabel polysilicon 289 -327 289 -327 0 1
rlabel polysilicon 289 -333 289 -333 0 3
rlabel polysilicon 296 -327 296 -327 0 1
rlabel polysilicon 296 -333 296 -333 0 3
rlabel polysilicon 303 -327 303 -327 0 1
rlabel polysilicon 306 -327 306 -327 0 2
rlabel polysilicon 306 -333 306 -333 0 4
rlabel polysilicon 310 -327 310 -327 0 1
rlabel polysilicon 310 -333 310 -333 0 3
rlabel polysilicon 317 -327 317 -327 0 1
rlabel polysilicon 317 -333 317 -333 0 3
rlabel polysilicon 324 -327 324 -327 0 1
rlabel polysilicon 324 -333 324 -333 0 3
rlabel polysilicon 331 -327 331 -327 0 1
rlabel polysilicon 331 -333 331 -333 0 3
rlabel polysilicon 338 -327 338 -327 0 1
rlabel polysilicon 338 -333 338 -333 0 3
rlabel polysilicon 345 -327 345 -327 0 1
rlabel polysilicon 345 -333 345 -333 0 3
rlabel polysilicon 352 -327 352 -327 0 1
rlabel polysilicon 352 -333 352 -333 0 3
rlabel polysilicon 359 -327 359 -327 0 1
rlabel polysilicon 359 -333 359 -333 0 3
rlabel polysilicon 366 -327 366 -327 0 1
rlabel polysilicon 366 -333 366 -333 0 3
rlabel polysilicon 376 -327 376 -327 0 2
rlabel polysilicon 373 -333 373 -333 0 3
rlabel polysilicon 376 -333 376 -333 0 4
rlabel polysilicon 380 -327 380 -327 0 1
rlabel polysilicon 383 -327 383 -327 0 2
rlabel polysilicon 383 -333 383 -333 0 4
rlabel polysilicon 387 -327 387 -327 0 1
rlabel polysilicon 387 -333 387 -333 0 3
rlabel polysilicon 394 -327 394 -327 0 1
rlabel polysilicon 397 -327 397 -327 0 2
rlabel polysilicon 394 -333 394 -333 0 3
rlabel polysilicon 397 -333 397 -333 0 4
rlabel polysilicon 404 -327 404 -327 0 2
rlabel polysilicon 401 -333 401 -333 0 3
rlabel polysilicon 404 -333 404 -333 0 4
rlabel polysilicon 408 -327 408 -327 0 1
rlabel polysilicon 408 -333 408 -333 0 3
rlabel polysilicon 418 -327 418 -327 0 2
rlabel polysilicon 415 -333 415 -333 0 3
rlabel polysilicon 418 -333 418 -333 0 4
rlabel polysilicon 422 -327 422 -327 0 1
rlabel polysilicon 425 -327 425 -327 0 2
rlabel polysilicon 422 -333 422 -333 0 3
rlabel polysilicon 425 -333 425 -333 0 4
rlabel polysilicon 429 -327 429 -327 0 1
rlabel polysilicon 429 -333 429 -333 0 3
rlabel polysilicon 436 -327 436 -327 0 1
rlabel polysilicon 439 -327 439 -327 0 2
rlabel polysilicon 436 -333 436 -333 0 3
rlabel polysilicon 439 -333 439 -333 0 4
rlabel polysilicon 443 -327 443 -327 0 1
rlabel polysilicon 446 -327 446 -327 0 2
rlabel polysilicon 443 -333 443 -333 0 3
rlabel polysilicon 446 -333 446 -333 0 4
rlabel polysilicon 450 -327 450 -327 0 1
rlabel polysilicon 453 -327 453 -327 0 2
rlabel polysilicon 453 -333 453 -333 0 4
rlabel polysilicon 457 -327 457 -327 0 1
rlabel polysilicon 457 -333 457 -333 0 3
rlabel polysilicon 460 -333 460 -333 0 4
rlabel polysilicon 467 -327 467 -327 0 2
rlabel polysilicon 464 -333 464 -333 0 3
rlabel polysilicon 467 -333 467 -333 0 4
rlabel polysilicon 471 -327 471 -327 0 1
rlabel polysilicon 474 -327 474 -327 0 2
rlabel polysilicon 471 -333 471 -333 0 3
rlabel polysilicon 474 -333 474 -333 0 4
rlabel polysilicon 478 -327 478 -327 0 1
rlabel polysilicon 478 -333 478 -333 0 3
rlabel polysilicon 485 -327 485 -327 0 1
rlabel polysilicon 488 -327 488 -327 0 2
rlabel polysilicon 485 -333 485 -333 0 3
rlabel polysilicon 488 -333 488 -333 0 4
rlabel polysilicon 492 -327 492 -327 0 1
rlabel polysilicon 492 -333 492 -333 0 3
rlabel polysilicon 499 -327 499 -327 0 1
rlabel polysilicon 499 -333 499 -333 0 3
rlabel polysilicon 506 -327 506 -327 0 1
rlabel polysilicon 506 -333 506 -333 0 3
rlabel polysilicon 513 -327 513 -327 0 1
rlabel polysilicon 513 -333 513 -333 0 3
rlabel polysilicon 520 -327 520 -327 0 1
rlabel polysilicon 520 -333 520 -333 0 3
rlabel polysilicon 527 -333 527 -333 0 3
rlabel polysilicon 534 -327 534 -327 0 1
rlabel polysilicon 534 -333 534 -333 0 3
rlabel polysilicon 541 -327 541 -327 0 1
rlabel polysilicon 541 -333 541 -333 0 3
rlabel polysilicon 548 -327 548 -327 0 1
rlabel polysilicon 551 -327 551 -327 0 2
rlabel polysilicon 548 -333 548 -333 0 3
rlabel polysilicon 551 -333 551 -333 0 4
rlabel polysilicon 555 -327 555 -327 0 1
rlabel polysilicon 555 -333 555 -333 0 3
rlabel polysilicon 562 -327 562 -327 0 1
rlabel polysilicon 562 -333 562 -333 0 3
rlabel polysilicon 569 -327 569 -327 0 1
rlabel polysilicon 569 -333 569 -333 0 3
rlabel polysilicon 572 -333 572 -333 0 4
rlabel polysilicon 576 -327 576 -327 0 1
rlabel polysilicon 579 -327 579 -327 0 2
rlabel polysilicon 576 -333 576 -333 0 3
rlabel polysilicon 583 -327 583 -327 0 1
rlabel polysilicon 583 -333 583 -333 0 3
rlabel polysilicon 590 -327 590 -327 0 1
rlabel polysilicon 590 -333 590 -333 0 3
rlabel polysilicon 597 -327 597 -327 0 1
rlabel polysilicon 597 -333 597 -333 0 3
rlabel polysilicon 604 -327 604 -327 0 1
rlabel polysilicon 604 -333 604 -333 0 3
rlabel polysilicon 611 -327 611 -327 0 1
rlabel polysilicon 611 -333 611 -333 0 3
rlabel polysilicon 618 -327 618 -327 0 1
rlabel polysilicon 618 -333 618 -333 0 3
rlabel polysilicon 625 -327 625 -327 0 1
rlabel polysilicon 625 -333 625 -333 0 3
rlabel polysilicon 632 -327 632 -327 0 1
rlabel polysilicon 632 -333 632 -333 0 3
rlabel polysilicon 639 -327 639 -327 0 1
rlabel polysilicon 639 -333 639 -333 0 3
rlabel polysilicon 646 -327 646 -327 0 1
rlabel polysilicon 646 -333 646 -333 0 3
rlabel polysilicon 653 -327 653 -327 0 1
rlabel polysilicon 653 -333 653 -333 0 3
rlabel polysilicon 660 -327 660 -327 0 1
rlabel polysilicon 660 -333 660 -333 0 3
rlabel polysilicon 667 -327 667 -327 0 1
rlabel polysilicon 667 -333 667 -333 0 3
rlabel polysilicon 674 -327 674 -327 0 1
rlabel polysilicon 674 -333 674 -333 0 3
rlabel polysilicon 681 -327 681 -327 0 1
rlabel polysilicon 681 -333 681 -333 0 3
rlabel polysilicon 688 -327 688 -327 0 1
rlabel polysilicon 688 -333 688 -333 0 3
rlabel polysilicon 695 -327 695 -327 0 1
rlabel polysilicon 695 -333 695 -333 0 3
rlabel polysilicon 702 -327 702 -327 0 1
rlabel polysilicon 702 -333 702 -333 0 3
rlabel polysilicon 709 -327 709 -327 0 1
rlabel polysilicon 709 -333 709 -333 0 3
rlabel polysilicon 716 -327 716 -327 0 1
rlabel polysilicon 716 -333 716 -333 0 3
rlabel polysilicon 723 -327 723 -327 0 1
rlabel polysilicon 723 -333 723 -333 0 3
rlabel polysilicon 730 -327 730 -327 0 1
rlabel polysilicon 730 -333 730 -333 0 3
rlabel polysilicon 737 -327 737 -327 0 1
rlabel polysilicon 737 -333 737 -333 0 3
rlabel polysilicon 744 -327 744 -327 0 1
rlabel polysilicon 744 -333 744 -333 0 3
rlabel polysilicon 751 -327 751 -327 0 1
rlabel polysilicon 751 -333 751 -333 0 3
rlabel polysilicon 758 -327 758 -327 0 1
rlabel polysilicon 758 -333 758 -333 0 3
rlabel polysilicon 765 -327 765 -327 0 1
rlabel polysilicon 765 -333 765 -333 0 3
rlabel polysilicon 772 -327 772 -327 0 1
rlabel polysilicon 772 -333 772 -333 0 3
rlabel polysilicon 779 -327 779 -327 0 1
rlabel polysilicon 779 -333 779 -333 0 3
rlabel polysilicon 786 -327 786 -327 0 1
rlabel polysilicon 786 -333 786 -333 0 3
rlabel polysilicon 793 -327 793 -327 0 1
rlabel polysilicon 793 -333 793 -333 0 3
rlabel polysilicon 800 -327 800 -327 0 1
rlabel polysilicon 800 -333 800 -333 0 3
rlabel polysilicon 807 -327 807 -327 0 1
rlabel polysilicon 807 -333 807 -333 0 3
rlabel polysilicon 814 -327 814 -327 0 1
rlabel polysilicon 814 -333 814 -333 0 3
rlabel polysilicon 821 -327 821 -327 0 1
rlabel polysilicon 821 -333 821 -333 0 3
rlabel polysilicon 828 -327 828 -327 0 1
rlabel polysilicon 828 -333 828 -333 0 3
rlabel polysilicon 835 -327 835 -327 0 1
rlabel polysilicon 835 -333 835 -333 0 3
rlabel polysilicon 842 -327 842 -327 0 1
rlabel polysilicon 842 -333 842 -333 0 3
rlabel polysilicon 849 -327 849 -327 0 1
rlabel polysilicon 849 -333 849 -333 0 3
rlabel polysilicon 856 -327 856 -327 0 1
rlabel polysilicon 856 -333 856 -333 0 3
rlabel polysilicon 863 -327 863 -327 0 1
rlabel polysilicon 863 -333 863 -333 0 3
rlabel polysilicon 870 -327 870 -327 0 1
rlabel polysilicon 870 -333 870 -333 0 3
rlabel polysilicon 877 -327 877 -327 0 1
rlabel polysilicon 877 -333 877 -333 0 3
rlabel polysilicon 884 -327 884 -327 0 1
rlabel polysilicon 884 -333 884 -333 0 3
rlabel polysilicon 891 -327 891 -327 0 1
rlabel polysilicon 891 -333 891 -333 0 3
rlabel polysilicon 898 -327 898 -327 0 1
rlabel polysilicon 898 -333 898 -333 0 3
rlabel polysilicon 905 -327 905 -327 0 1
rlabel polysilicon 905 -333 905 -333 0 3
rlabel polysilicon 912 -327 912 -327 0 1
rlabel polysilicon 912 -333 912 -333 0 3
rlabel polysilicon 919 -327 919 -327 0 1
rlabel polysilicon 919 -333 919 -333 0 3
rlabel polysilicon 926 -327 926 -327 0 1
rlabel polysilicon 926 -333 926 -333 0 3
rlabel polysilicon 933 -327 933 -327 0 1
rlabel polysilicon 933 -333 933 -333 0 3
rlabel polysilicon 940 -327 940 -327 0 1
rlabel polysilicon 940 -333 940 -333 0 3
rlabel polysilicon 947 -327 947 -327 0 1
rlabel polysilicon 947 -333 947 -333 0 3
rlabel polysilicon 954 -327 954 -327 0 1
rlabel polysilicon 954 -333 954 -333 0 3
rlabel polysilicon 2 -414 2 -414 0 1
rlabel polysilicon 2 -420 2 -420 0 3
rlabel polysilicon 9 -414 9 -414 0 1
rlabel polysilicon 9 -420 9 -420 0 3
rlabel polysilicon 16 -414 16 -414 0 1
rlabel polysilicon 16 -420 16 -420 0 3
rlabel polysilicon 23 -414 23 -414 0 1
rlabel polysilicon 23 -420 23 -420 0 3
rlabel polysilicon 30 -414 30 -414 0 1
rlabel polysilicon 30 -420 30 -420 0 3
rlabel polysilicon 37 -414 37 -414 0 1
rlabel polysilicon 37 -420 37 -420 0 3
rlabel polysilicon 44 -414 44 -414 0 1
rlabel polysilicon 44 -420 44 -420 0 3
rlabel polysilicon 51 -414 51 -414 0 1
rlabel polysilicon 51 -420 51 -420 0 3
rlabel polysilicon 58 -414 58 -414 0 1
rlabel polysilicon 58 -420 58 -420 0 3
rlabel polysilicon 65 -414 65 -414 0 1
rlabel polysilicon 68 -414 68 -414 0 2
rlabel polysilicon 65 -420 65 -420 0 3
rlabel polysilicon 68 -420 68 -420 0 4
rlabel polysilicon 72 -414 72 -414 0 1
rlabel polysilicon 75 -414 75 -414 0 2
rlabel polysilicon 72 -420 72 -420 0 3
rlabel polysilicon 75 -420 75 -420 0 4
rlabel polysilicon 79 -414 79 -414 0 1
rlabel polysilicon 82 -414 82 -414 0 2
rlabel polysilicon 79 -420 79 -420 0 3
rlabel polysilicon 82 -420 82 -420 0 4
rlabel polysilicon 86 -414 86 -414 0 1
rlabel polysilicon 89 -414 89 -414 0 2
rlabel polysilicon 93 -414 93 -414 0 1
rlabel polysilicon 96 -414 96 -414 0 2
rlabel polysilicon 93 -420 93 -420 0 3
rlabel polysilicon 96 -420 96 -420 0 4
rlabel polysilicon 100 -414 100 -414 0 1
rlabel polysilicon 100 -420 100 -420 0 3
rlabel polysilicon 107 -414 107 -414 0 1
rlabel polysilicon 107 -420 107 -420 0 3
rlabel polysilicon 114 -414 114 -414 0 1
rlabel polysilicon 114 -420 114 -420 0 3
rlabel polysilicon 121 -414 121 -414 0 1
rlabel polysilicon 124 -414 124 -414 0 2
rlabel polysilicon 121 -420 121 -420 0 3
rlabel polysilicon 124 -420 124 -420 0 4
rlabel polysilicon 128 -414 128 -414 0 1
rlabel polysilicon 128 -420 128 -420 0 3
rlabel polysilicon 135 -414 135 -414 0 1
rlabel polysilicon 135 -420 135 -420 0 3
rlabel polysilicon 142 -414 142 -414 0 1
rlabel polysilicon 142 -420 142 -420 0 3
rlabel polysilicon 149 -414 149 -414 0 1
rlabel polysilicon 149 -420 149 -420 0 3
rlabel polysilicon 156 -414 156 -414 0 1
rlabel polysilicon 159 -414 159 -414 0 2
rlabel polysilicon 156 -420 156 -420 0 3
rlabel polysilicon 159 -420 159 -420 0 4
rlabel polysilicon 163 -414 163 -414 0 1
rlabel polysilicon 163 -420 163 -420 0 3
rlabel polysilicon 170 -414 170 -414 0 1
rlabel polysilicon 170 -420 170 -420 0 3
rlabel polysilicon 177 -414 177 -414 0 1
rlabel polysilicon 177 -420 177 -420 0 3
rlabel polysilicon 184 -414 184 -414 0 1
rlabel polysilicon 184 -420 184 -420 0 3
rlabel polysilicon 187 -420 187 -420 0 4
rlabel polysilicon 191 -414 191 -414 0 1
rlabel polysilicon 194 -414 194 -414 0 2
rlabel polysilicon 191 -420 191 -420 0 3
rlabel polysilicon 198 -414 198 -414 0 1
rlabel polysilicon 198 -420 198 -420 0 3
rlabel polysilicon 205 -414 205 -414 0 1
rlabel polysilicon 205 -420 205 -420 0 3
rlabel polysilicon 212 -414 212 -414 0 1
rlabel polysilicon 212 -420 212 -420 0 3
rlabel polysilicon 219 -414 219 -414 0 1
rlabel polysilicon 219 -420 219 -420 0 3
rlabel polysilicon 226 -414 226 -414 0 1
rlabel polysilicon 226 -420 226 -420 0 3
rlabel polysilicon 233 -414 233 -414 0 1
rlabel polysilicon 233 -420 233 -420 0 3
rlabel polysilicon 240 -414 240 -414 0 1
rlabel polysilicon 243 -414 243 -414 0 2
rlabel polysilicon 240 -420 240 -420 0 3
rlabel polysilicon 243 -420 243 -420 0 4
rlabel polysilicon 247 -414 247 -414 0 1
rlabel polysilicon 247 -420 247 -420 0 3
rlabel polysilicon 254 -414 254 -414 0 1
rlabel polysilicon 254 -420 254 -420 0 3
rlabel polysilicon 261 -414 261 -414 0 1
rlabel polysilicon 261 -420 261 -420 0 3
rlabel polysilicon 268 -414 268 -414 0 1
rlabel polysilicon 268 -420 268 -420 0 3
rlabel polysilicon 275 -414 275 -414 0 1
rlabel polysilicon 275 -420 275 -420 0 3
rlabel polysilicon 282 -414 282 -414 0 1
rlabel polysilicon 282 -420 282 -420 0 3
rlabel polysilicon 289 -414 289 -414 0 1
rlabel polysilicon 289 -420 289 -420 0 3
rlabel polysilicon 296 -414 296 -414 0 1
rlabel polysilicon 296 -420 296 -420 0 3
rlabel polysilicon 303 -414 303 -414 0 1
rlabel polysilicon 303 -420 303 -420 0 3
rlabel polysilicon 310 -414 310 -414 0 1
rlabel polysilicon 310 -420 310 -420 0 3
rlabel polysilicon 317 -414 317 -414 0 1
rlabel polysilicon 317 -420 317 -420 0 3
rlabel polysilicon 324 -414 324 -414 0 1
rlabel polysilicon 324 -420 324 -420 0 3
rlabel polysilicon 331 -414 331 -414 0 1
rlabel polysilicon 331 -420 331 -420 0 3
rlabel polysilicon 338 -414 338 -414 0 1
rlabel polysilicon 338 -420 338 -420 0 3
rlabel polysilicon 345 -414 345 -414 0 1
rlabel polysilicon 345 -420 345 -420 0 3
rlabel polysilicon 352 -414 352 -414 0 1
rlabel polysilicon 355 -414 355 -414 0 2
rlabel polysilicon 359 -414 359 -414 0 1
rlabel polysilicon 362 -414 362 -414 0 2
rlabel polysilicon 359 -420 359 -420 0 3
rlabel polysilicon 362 -420 362 -420 0 4
rlabel polysilicon 366 -414 366 -414 0 1
rlabel polysilicon 366 -420 366 -420 0 3
rlabel polysilicon 373 -414 373 -414 0 1
rlabel polysilicon 373 -420 373 -420 0 3
rlabel polysilicon 380 -414 380 -414 0 1
rlabel polysilicon 380 -420 380 -420 0 3
rlabel polysilicon 387 -414 387 -414 0 1
rlabel polysilicon 387 -420 387 -420 0 3
rlabel polysilicon 394 -414 394 -414 0 1
rlabel polysilicon 397 -414 397 -414 0 2
rlabel polysilicon 394 -420 394 -420 0 3
rlabel polysilicon 397 -420 397 -420 0 4
rlabel polysilicon 401 -414 401 -414 0 1
rlabel polysilicon 401 -420 401 -420 0 3
rlabel polysilicon 408 -414 408 -414 0 1
rlabel polysilicon 411 -414 411 -414 0 2
rlabel polysilicon 408 -420 408 -420 0 3
rlabel polysilicon 411 -420 411 -420 0 4
rlabel polysilicon 415 -414 415 -414 0 1
rlabel polysilicon 415 -420 415 -420 0 3
rlabel polysilicon 422 -414 422 -414 0 1
rlabel polysilicon 422 -420 422 -420 0 3
rlabel polysilicon 429 -414 429 -414 0 1
rlabel polysilicon 432 -414 432 -414 0 2
rlabel polysilicon 429 -420 429 -420 0 3
rlabel polysilicon 432 -420 432 -420 0 4
rlabel polysilicon 436 -414 436 -414 0 1
rlabel polysilicon 436 -420 436 -420 0 3
rlabel polysilicon 443 -414 443 -414 0 1
rlabel polysilicon 443 -420 443 -420 0 3
rlabel polysilicon 450 -414 450 -414 0 1
rlabel polysilicon 450 -420 450 -420 0 3
rlabel polysilicon 457 -414 457 -414 0 1
rlabel polysilicon 460 -414 460 -414 0 2
rlabel polysilicon 457 -420 457 -420 0 3
rlabel polysilicon 460 -420 460 -420 0 4
rlabel polysilicon 464 -414 464 -414 0 1
rlabel polysilicon 467 -414 467 -414 0 2
rlabel polysilicon 464 -420 464 -420 0 3
rlabel polysilicon 467 -420 467 -420 0 4
rlabel polysilicon 471 -414 471 -414 0 1
rlabel polysilicon 471 -420 471 -420 0 3
rlabel polysilicon 478 -414 478 -414 0 1
rlabel polysilicon 478 -420 478 -420 0 3
rlabel polysilicon 485 -414 485 -414 0 1
rlabel polysilicon 485 -420 485 -420 0 3
rlabel polysilicon 492 -414 492 -414 0 1
rlabel polysilicon 492 -420 492 -420 0 3
rlabel polysilicon 499 -414 499 -414 0 1
rlabel polysilicon 499 -420 499 -420 0 3
rlabel polysilicon 506 -414 506 -414 0 1
rlabel polysilicon 506 -420 506 -420 0 3
rlabel polysilicon 513 -414 513 -414 0 1
rlabel polysilicon 516 -414 516 -414 0 2
rlabel polysilicon 516 -420 516 -420 0 4
rlabel polysilicon 520 -414 520 -414 0 1
rlabel polysilicon 520 -420 520 -420 0 3
rlabel polysilicon 527 -414 527 -414 0 1
rlabel polysilicon 530 -414 530 -414 0 2
rlabel polysilicon 527 -420 527 -420 0 3
rlabel polysilicon 530 -420 530 -420 0 4
rlabel polysilicon 534 -414 534 -414 0 1
rlabel polysilicon 534 -420 534 -420 0 3
rlabel polysilicon 541 -414 541 -414 0 1
rlabel polysilicon 541 -420 541 -420 0 3
rlabel polysilicon 551 -414 551 -414 0 2
rlabel polysilicon 548 -420 548 -420 0 3
rlabel polysilicon 551 -420 551 -420 0 4
rlabel polysilicon 555 -414 555 -414 0 1
rlabel polysilicon 555 -420 555 -420 0 3
rlabel polysilicon 562 -414 562 -414 0 1
rlabel polysilicon 562 -420 562 -420 0 3
rlabel polysilicon 569 -414 569 -414 0 1
rlabel polysilicon 569 -420 569 -420 0 3
rlabel polysilicon 576 -414 576 -414 0 1
rlabel polysilicon 576 -420 576 -420 0 3
rlabel polysilicon 583 -414 583 -414 0 1
rlabel polysilicon 583 -420 583 -420 0 3
rlabel polysilicon 590 -414 590 -414 0 1
rlabel polysilicon 590 -420 590 -420 0 3
rlabel polysilicon 597 -414 597 -414 0 1
rlabel polysilicon 597 -420 597 -420 0 3
rlabel polysilicon 604 -414 604 -414 0 1
rlabel polysilicon 604 -420 604 -420 0 3
rlabel polysilicon 611 -414 611 -414 0 1
rlabel polysilicon 611 -420 611 -420 0 3
rlabel polysilicon 618 -414 618 -414 0 1
rlabel polysilicon 621 -414 621 -414 0 2
rlabel polysilicon 618 -420 618 -420 0 3
rlabel polysilicon 621 -420 621 -420 0 4
rlabel polysilicon 625 -414 625 -414 0 1
rlabel polysilicon 625 -420 625 -420 0 3
rlabel polysilicon 632 -414 632 -414 0 1
rlabel polysilicon 632 -420 632 -420 0 3
rlabel polysilicon 639 -414 639 -414 0 1
rlabel polysilicon 639 -420 639 -420 0 3
rlabel polysilicon 646 -414 646 -414 0 1
rlabel polysilicon 646 -420 646 -420 0 3
rlabel polysilicon 653 -414 653 -414 0 1
rlabel polysilicon 653 -420 653 -420 0 3
rlabel polysilicon 660 -414 660 -414 0 1
rlabel polysilicon 660 -420 660 -420 0 3
rlabel polysilicon 667 -414 667 -414 0 1
rlabel polysilicon 667 -420 667 -420 0 3
rlabel polysilicon 674 -414 674 -414 0 1
rlabel polysilicon 674 -420 674 -420 0 3
rlabel polysilicon 681 -414 681 -414 0 1
rlabel polysilicon 681 -420 681 -420 0 3
rlabel polysilicon 688 -414 688 -414 0 1
rlabel polysilicon 688 -420 688 -420 0 3
rlabel polysilicon 695 -414 695 -414 0 1
rlabel polysilicon 695 -420 695 -420 0 3
rlabel polysilicon 702 -414 702 -414 0 1
rlabel polysilicon 702 -420 702 -420 0 3
rlabel polysilicon 709 -414 709 -414 0 1
rlabel polysilicon 709 -420 709 -420 0 3
rlabel polysilicon 716 -414 716 -414 0 1
rlabel polysilicon 716 -420 716 -420 0 3
rlabel polysilicon 723 -414 723 -414 0 1
rlabel polysilicon 723 -420 723 -420 0 3
rlabel polysilicon 730 -414 730 -414 0 1
rlabel polysilicon 730 -420 730 -420 0 3
rlabel polysilicon 737 -414 737 -414 0 1
rlabel polysilicon 737 -420 737 -420 0 3
rlabel polysilicon 744 -414 744 -414 0 1
rlabel polysilicon 744 -420 744 -420 0 3
rlabel polysilicon 751 -414 751 -414 0 1
rlabel polysilicon 751 -420 751 -420 0 3
rlabel polysilicon 758 -414 758 -414 0 1
rlabel polysilicon 758 -420 758 -420 0 3
rlabel polysilicon 765 -414 765 -414 0 1
rlabel polysilicon 765 -420 765 -420 0 3
rlabel polysilicon 772 -414 772 -414 0 1
rlabel polysilicon 772 -420 772 -420 0 3
rlabel polysilicon 779 -414 779 -414 0 1
rlabel polysilicon 779 -420 779 -420 0 3
rlabel polysilicon 786 -414 786 -414 0 1
rlabel polysilicon 786 -420 786 -420 0 3
rlabel polysilicon 793 -414 793 -414 0 1
rlabel polysilicon 793 -420 793 -420 0 3
rlabel polysilicon 800 -414 800 -414 0 1
rlabel polysilicon 800 -420 800 -420 0 3
rlabel polysilicon 807 -414 807 -414 0 1
rlabel polysilicon 807 -420 807 -420 0 3
rlabel polysilicon 814 -414 814 -414 0 1
rlabel polysilicon 814 -420 814 -420 0 3
rlabel polysilicon 821 -414 821 -414 0 1
rlabel polysilicon 821 -420 821 -420 0 3
rlabel polysilicon 828 -414 828 -414 0 1
rlabel polysilicon 828 -420 828 -420 0 3
rlabel polysilicon 835 -414 835 -414 0 1
rlabel polysilicon 835 -420 835 -420 0 3
rlabel polysilicon 842 -414 842 -414 0 1
rlabel polysilicon 842 -420 842 -420 0 3
rlabel polysilicon 849 -414 849 -414 0 1
rlabel polysilicon 849 -420 849 -420 0 3
rlabel polysilicon 856 -414 856 -414 0 1
rlabel polysilicon 856 -420 856 -420 0 3
rlabel polysilicon 863 -414 863 -414 0 1
rlabel polysilicon 863 -420 863 -420 0 3
rlabel polysilicon 870 -414 870 -414 0 1
rlabel polysilicon 870 -420 870 -420 0 3
rlabel polysilicon 877 -414 877 -414 0 1
rlabel polysilicon 877 -420 877 -420 0 3
rlabel polysilicon 884 -414 884 -414 0 1
rlabel polysilicon 884 -420 884 -420 0 3
rlabel polysilicon 891 -414 891 -414 0 1
rlabel polysilicon 891 -420 891 -420 0 3
rlabel polysilicon 898 -414 898 -414 0 1
rlabel polysilicon 898 -420 898 -420 0 3
rlabel polysilicon 905 -414 905 -414 0 1
rlabel polysilicon 905 -420 905 -420 0 3
rlabel polysilicon 912 -414 912 -414 0 1
rlabel polysilicon 912 -420 912 -420 0 3
rlabel polysilicon 919 -414 919 -414 0 1
rlabel polysilicon 919 -420 919 -420 0 3
rlabel polysilicon 926 -414 926 -414 0 1
rlabel polysilicon 926 -420 926 -420 0 3
rlabel polysilicon 933 -414 933 -414 0 1
rlabel polysilicon 933 -420 933 -420 0 3
rlabel polysilicon 940 -414 940 -414 0 1
rlabel polysilicon 940 -420 940 -420 0 3
rlabel polysilicon 947 -414 947 -414 0 1
rlabel polysilicon 947 -420 947 -420 0 3
rlabel polysilicon 954 -414 954 -414 0 1
rlabel polysilicon 954 -420 954 -420 0 3
rlabel polysilicon 961 -414 961 -414 0 1
rlabel polysilicon 961 -420 961 -420 0 3
rlabel polysilicon 968 -414 968 -414 0 1
rlabel polysilicon 968 -420 968 -420 0 3
rlabel polysilicon 975 -414 975 -414 0 1
rlabel polysilicon 975 -420 975 -420 0 3
rlabel polysilicon 982 -414 982 -414 0 1
rlabel polysilicon 982 -420 982 -420 0 3
rlabel polysilicon 989 -414 989 -414 0 1
rlabel polysilicon 989 -420 989 -420 0 3
rlabel polysilicon 996 -414 996 -414 0 1
rlabel polysilicon 996 -420 996 -420 0 3
rlabel polysilicon 1003 -414 1003 -414 0 1
rlabel polysilicon 1003 -420 1003 -420 0 3
rlabel polysilicon 1024 -414 1024 -414 0 1
rlabel polysilicon 1024 -420 1024 -420 0 3
rlabel polysilicon 2 -509 2 -509 0 1
rlabel polysilicon 2 -515 2 -515 0 3
rlabel polysilicon 9 -509 9 -509 0 1
rlabel polysilicon 9 -515 9 -515 0 3
rlabel polysilicon 16 -509 16 -509 0 1
rlabel polysilicon 16 -515 16 -515 0 3
rlabel polysilicon 23 -509 23 -509 0 1
rlabel polysilicon 23 -515 23 -515 0 3
rlabel polysilicon 30 -509 30 -509 0 1
rlabel polysilicon 30 -515 30 -515 0 3
rlabel polysilicon 37 -509 37 -509 0 1
rlabel polysilicon 37 -515 37 -515 0 3
rlabel polysilicon 44 -509 44 -509 0 1
rlabel polysilicon 44 -515 44 -515 0 3
rlabel polysilicon 51 -509 51 -509 0 1
rlabel polysilicon 51 -515 51 -515 0 3
rlabel polysilicon 58 -509 58 -509 0 1
rlabel polysilicon 58 -515 58 -515 0 3
rlabel polysilicon 65 -509 65 -509 0 1
rlabel polysilicon 65 -515 65 -515 0 3
rlabel polysilicon 72 -509 72 -509 0 1
rlabel polysilicon 72 -515 72 -515 0 3
rlabel polysilicon 79 -509 79 -509 0 1
rlabel polysilicon 79 -515 79 -515 0 3
rlabel polysilicon 86 -509 86 -509 0 1
rlabel polysilicon 86 -515 86 -515 0 3
rlabel polysilicon 93 -509 93 -509 0 1
rlabel polysilicon 96 -509 96 -509 0 2
rlabel polysilicon 93 -515 93 -515 0 3
rlabel polysilicon 100 -509 100 -509 0 1
rlabel polysilicon 100 -515 100 -515 0 3
rlabel polysilicon 107 -509 107 -509 0 1
rlabel polysilicon 107 -515 107 -515 0 3
rlabel polysilicon 114 -509 114 -509 0 1
rlabel polysilicon 114 -515 114 -515 0 3
rlabel polysilicon 121 -509 121 -509 0 1
rlabel polysilicon 121 -515 121 -515 0 3
rlabel polysilicon 128 -509 128 -509 0 1
rlabel polysilicon 131 -509 131 -509 0 2
rlabel polysilicon 128 -515 128 -515 0 3
rlabel polysilicon 131 -515 131 -515 0 4
rlabel polysilicon 138 -509 138 -509 0 2
rlabel polysilicon 135 -515 135 -515 0 3
rlabel polysilicon 138 -515 138 -515 0 4
rlabel polysilicon 145 -515 145 -515 0 4
rlabel polysilicon 152 -509 152 -509 0 2
rlabel polysilicon 152 -515 152 -515 0 4
rlabel polysilicon 156 -509 156 -509 0 1
rlabel polysilicon 156 -515 156 -515 0 3
rlabel polysilicon 159 -515 159 -515 0 4
rlabel polysilicon 163 -509 163 -509 0 1
rlabel polysilicon 163 -515 163 -515 0 3
rlabel polysilicon 170 -509 170 -509 0 1
rlabel polysilicon 170 -515 170 -515 0 3
rlabel polysilicon 177 -509 177 -509 0 1
rlabel polysilicon 177 -515 177 -515 0 3
rlabel polysilicon 184 -509 184 -509 0 1
rlabel polysilicon 184 -515 184 -515 0 3
rlabel polysilicon 191 -509 191 -509 0 1
rlabel polysilicon 191 -515 191 -515 0 3
rlabel polysilicon 198 -509 198 -509 0 1
rlabel polysilicon 198 -515 198 -515 0 3
rlabel polysilicon 205 -509 205 -509 0 1
rlabel polysilicon 205 -515 205 -515 0 3
rlabel polysilicon 212 -509 212 -509 0 1
rlabel polysilicon 212 -515 212 -515 0 3
rlabel polysilicon 219 -509 219 -509 0 1
rlabel polysilicon 219 -515 219 -515 0 3
rlabel polysilicon 226 -509 226 -509 0 1
rlabel polysilicon 226 -515 226 -515 0 3
rlabel polysilicon 233 -509 233 -509 0 1
rlabel polysilicon 233 -515 233 -515 0 3
rlabel polysilicon 240 -509 240 -509 0 1
rlabel polysilicon 240 -515 240 -515 0 3
rlabel polysilicon 247 -509 247 -509 0 1
rlabel polysilicon 250 -509 250 -509 0 2
rlabel polysilicon 247 -515 247 -515 0 3
rlabel polysilicon 250 -515 250 -515 0 4
rlabel polysilicon 254 -509 254 -509 0 1
rlabel polysilicon 254 -515 254 -515 0 3
rlabel polysilicon 261 -509 261 -509 0 1
rlabel polysilicon 261 -515 261 -515 0 3
rlabel polysilicon 268 -509 268 -509 0 1
rlabel polysilicon 268 -515 268 -515 0 3
rlabel polysilicon 275 -509 275 -509 0 1
rlabel polysilicon 275 -515 275 -515 0 3
rlabel polysilicon 282 -509 282 -509 0 1
rlabel polysilicon 282 -515 282 -515 0 3
rlabel polysilicon 289 -509 289 -509 0 1
rlabel polysilicon 289 -515 289 -515 0 3
rlabel polysilicon 296 -509 296 -509 0 1
rlabel polysilicon 296 -515 296 -515 0 3
rlabel polysilicon 303 -509 303 -509 0 1
rlabel polysilicon 303 -515 303 -515 0 3
rlabel polysilicon 310 -509 310 -509 0 1
rlabel polysilicon 310 -515 310 -515 0 3
rlabel polysilicon 317 -509 317 -509 0 1
rlabel polysilicon 317 -515 317 -515 0 3
rlabel polysilicon 324 -509 324 -509 0 1
rlabel polysilicon 327 -509 327 -509 0 2
rlabel polysilicon 331 -509 331 -509 0 1
rlabel polysilicon 331 -515 331 -515 0 3
rlabel polysilicon 338 -509 338 -509 0 1
rlabel polysilicon 338 -515 338 -515 0 3
rlabel polysilicon 345 -509 345 -509 0 1
rlabel polysilicon 345 -515 345 -515 0 3
rlabel polysilicon 352 -509 352 -509 0 1
rlabel polysilicon 352 -515 352 -515 0 3
rlabel polysilicon 359 -509 359 -509 0 1
rlabel polysilicon 359 -515 359 -515 0 3
rlabel polysilicon 366 -509 366 -509 0 1
rlabel polysilicon 366 -515 366 -515 0 3
rlabel polysilicon 373 -509 373 -509 0 1
rlabel polysilicon 373 -515 373 -515 0 3
rlabel polysilicon 380 -509 380 -509 0 1
rlabel polysilicon 380 -515 380 -515 0 3
rlabel polysilicon 387 -509 387 -509 0 1
rlabel polysilicon 390 -509 390 -509 0 2
rlabel polysilicon 387 -515 387 -515 0 3
rlabel polysilicon 394 -509 394 -509 0 1
rlabel polysilicon 397 -509 397 -509 0 2
rlabel polysilicon 394 -515 394 -515 0 3
rlabel polysilicon 401 -509 401 -509 0 1
rlabel polysilicon 401 -515 401 -515 0 3
rlabel polysilicon 408 -509 408 -509 0 1
rlabel polysilicon 411 -509 411 -509 0 2
rlabel polysilicon 411 -515 411 -515 0 4
rlabel polysilicon 415 -509 415 -509 0 1
rlabel polysilicon 415 -515 415 -515 0 3
rlabel polysilicon 422 -509 422 -509 0 1
rlabel polysilicon 422 -515 422 -515 0 3
rlabel polysilicon 429 -509 429 -509 0 1
rlabel polysilicon 429 -515 429 -515 0 3
rlabel polysilicon 436 -509 436 -509 0 1
rlabel polysilicon 436 -515 436 -515 0 3
rlabel polysilicon 443 -509 443 -509 0 1
rlabel polysilicon 446 -509 446 -509 0 2
rlabel polysilicon 446 -515 446 -515 0 4
rlabel polysilicon 450 -509 450 -509 0 1
rlabel polysilicon 450 -515 450 -515 0 3
rlabel polysilicon 457 -509 457 -509 0 1
rlabel polysilicon 457 -515 457 -515 0 3
rlabel polysilicon 464 -509 464 -509 0 1
rlabel polysilicon 464 -515 464 -515 0 3
rlabel polysilicon 471 -509 471 -509 0 1
rlabel polysilicon 471 -515 471 -515 0 3
rlabel polysilicon 478 -509 478 -509 0 1
rlabel polysilicon 481 -509 481 -509 0 2
rlabel polysilicon 478 -515 478 -515 0 3
rlabel polysilicon 481 -515 481 -515 0 4
rlabel polysilicon 485 -509 485 -509 0 1
rlabel polysilicon 485 -515 485 -515 0 3
rlabel polysilicon 492 -509 492 -509 0 1
rlabel polysilicon 492 -515 492 -515 0 3
rlabel polysilicon 499 -509 499 -509 0 1
rlabel polysilicon 499 -515 499 -515 0 3
rlabel polysilicon 506 -509 506 -509 0 1
rlabel polysilicon 509 -509 509 -509 0 2
rlabel polysilicon 506 -515 506 -515 0 3
rlabel polysilicon 509 -515 509 -515 0 4
rlabel polysilicon 513 -509 513 -509 0 1
rlabel polysilicon 513 -515 513 -515 0 3
rlabel polysilicon 520 -509 520 -509 0 1
rlabel polysilicon 523 -509 523 -509 0 2
rlabel polysilicon 520 -515 520 -515 0 3
rlabel polysilicon 523 -515 523 -515 0 4
rlabel polysilicon 527 -509 527 -509 0 1
rlabel polysilicon 527 -515 527 -515 0 3
rlabel polysilicon 534 -509 534 -509 0 1
rlabel polysilicon 534 -515 534 -515 0 3
rlabel polysilicon 541 -509 541 -509 0 1
rlabel polysilicon 541 -515 541 -515 0 3
rlabel polysilicon 548 -509 548 -509 0 1
rlabel polysilicon 548 -515 548 -515 0 3
rlabel polysilicon 555 -509 555 -509 0 1
rlabel polysilicon 555 -515 555 -515 0 3
rlabel polysilicon 562 -509 562 -509 0 1
rlabel polysilicon 565 -509 565 -509 0 2
rlabel polysilicon 562 -515 562 -515 0 3
rlabel polysilicon 565 -515 565 -515 0 4
rlabel polysilicon 569 -509 569 -509 0 1
rlabel polysilicon 572 -509 572 -509 0 2
rlabel polysilicon 569 -515 569 -515 0 3
rlabel polysilicon 572 -515 572 -515 0 4
rlabel polysilicon 576 -509 576 -509 0 1
rlabel polysilicon 579 -509 579 -509 0 2
rlabel polysilicon 576 -515 576 -515 0 3
rlabel polysilicon 579 -515 579 -515 0 4
rlabel polysilicon 583 -509 583 -509 0 1
rlabel polysilicon 583 -515 583 -515 0 3
rlabel polysilicon 590 -509 590 -509 0 1
rlabel polysilicon 590 -515 590 -515 0 3
rlabel polysilicon 597 -509 597 -509 0 1
rlabel polysilicon 597 -515 597 -515 0 3
rlabel polysilicon 604 -509 604 -509 0 1
rlabel polysilicon 607 -509 607 -509 0 2
rlabel polysilicon 604 -515 604 -515 0 3
rlabel polysilicon 607 -515 607 -515 0 4
rlabel polysilicon 611 -509 611 -509 0 1
rlabel polysilicon 611 -515 611 -515 0 3
rlabel polysilicon 618 -509 618 -509 0 1
rlabel polysilicon 618 -515 618 -515 0 3
rlabel polysilicon 625 -509 625 -509 0 1
rlabel polysilicon 625 -515 625 -515 0 3
rlabel polysilicon 632 -509 632 -509 0 1
rlabel polysilicon 632 -515 632 -515 0 3
rlabel polysilicon 639 -509 639 -509 0 1
rlabel polysilicon 639 -515 639 -515 0 3
rlabel polysilicon 649 -509 649 -509 0 2
rlabel polysilicon 646 -515 646 -515 0 3
rlabel polysilicon 649 -515 649 -515 0 4
rlabel polysilicon 653 -509 653 -509 0 1
rlabel polysilicon 653 -515 653 -515 0 3
rlabel polysilicon 660 -509 660 -509 0 1
rlabel polysilicon 660 -515 660 -515 0 3
rlabel polysilicon 667 -509 667 -509 0 1
rlabel polysilicon 670 -509 670 -509 0 2
rlabel polysilicon 667 -515 667 -515 0 3
rlabel polysilicon 670 -515 670 -515 0 4
rlabel polysilicon 674 -509 674 -509 0 1
rlabel polysilicon 674 -515 674 -515 0 3
rlabel polysilicon 681 -509 681 -509 0 1
rlabel polysilicon 681 -515 681 -515 0 3
rlabel polysilicon 688 -509 688 -509 0 1
rlabel polysilicon 688 -515 688 -515 0 3
rlabel polysilicon 695 -509 695 -509 0 1
rlabel polysilicon 695 -515 695 -515 0 3
rlabel polysilicon 702 -509 702 -509 0 1
rlabel polysilicon 702 -515 702 -515 0 3
rlabel polysilicon 709 -509 709 -509 0 1
rlabel polysilicon 709 -515 709 -515 0 3
rlabel polysilicon 716 -509 716 -509 0 1
rlabel polysilicon 716 -515 716 -515 0 3
rlabel polysilicon 723 -509 723 -509 0 1
rlabel polysilicon 723 -515 723 -515 0 3
rlabel polysilicon 730 -509 730 -509 0 1
rlabel polysilicon 730 -515 730 -515 0 3
rlabel polysilicon 737 -509 737 -509 0 1
rlabel polysilicon 737 -515 737 -515 0 3
rlabel polysilicon 744 -509 744 -509 0 1
rlabel polysilicon 744 -515 744 -515 0 3
rlabel polysilicon 751 -509 751 -509 0 1
rlabel polysilicon 751 -515 751 -515 0 3
rlabel polysilicon 754 -515 754 -515 0 4
rlabel polysilicon 758 -509 758 -509 0 1
rlabel polysilicon 758 -515 758 -515 0 3
rlabel polysilicon 765 -509 765 -509 0 1
rlabel polysilicon 765 -515 765 -515 0 3
rlabel polysilicon 772 -509 772 -509 0 1
rlabel polysilicon 772 -515 772 -515 0 3
rlabel polysilicon 779 -509 779 -509 0 1
rlabel polysilicon 779 -515 779 -515 0 3
rlabel polysilicon 786 -509 786 -509 0 1
rlabel polysilicon 786 -515 786 -515 0 3
rlabel polysilicon 793 -509 793 -509 0 1
rlabel polysilicon 793 -515 793 -515 0 3
rlabel polysilicon 800 -509 800 -509 0 1
rlabel polysilicon 800 -515 800 -515 0 3
rlabel polysilicon 807 -509 807 -509 0 1
rlabel polysilicon 807 -515 807 -515 0 3
rlabel polysilicon 814 -509 814 -509 0 1
rlabel polysilicon 814 -515 814 -515 0 3
rlabel polysilicon 821 -509 821 -509 0 1
rlabel polysilicon 821 -515 821 -515 0 3
rlabel polysilicon 828 -509 828 -509 0 1
rlabel polysilicon 828 -515 828 -515 0 3
rlabel polysilicon 835 -509 835 -509 0 1
rlabel polysilicon 835 -515 835 -515 0 3
rlabel polysilicon 842 -509 842 -509 0 1
rlabel polysilicon 842 -515 842 -515 0 3
rlabel polysilicon 849 -509 849 -509 0 1
rlabel polysilicon 849 -515 849 -515 0 3
rlabel polysilicon 856 -509 856 -509 0 1
rlabel polysilicon 856 -515 856 -515 0 3
rlabel polysilicon 863 -509 863 -509 0 1
rlabel polysilicon 863 -515 863 -515 0 3
rlabel polysilicon 870 -509 870 -509 0 1
rlabel polysilicon 870 -515 870 -515 0 3
rlabel polysilicon 877 -509 877 -509 0 1
rlabel polysilicon 877 -515 877 -515 0 3
rlabel polysilicon 884 -509 884 -509 0 1
rlabel polysilicon 884 -515 884 -515 0 3
rlabel polysilicon 891 -509 891 -509 0 1
rlabel polysilicon 891 -515 891 -515 0 3
rlabel polysilicon 898 -509 898 -509 0 1
rlabel polysilicon 898 -515 898 -515 0 3
rlabel polysilicon 905 -509 905 -509 0 1
rlabel polysilicon 905 -515 905 -515 0 3
rlabel polysilicon 912 -509 912 -509 0 1
rlabel polysilicon 912 -515 912 -515 0 3
rlabel polysilicon 919 -509 919 -509 0 1
rlabel polysilicon 919 -515 919 -515 0 3
rlabel polysilicon 926 -509 926 -509 0 1
rlabel polysilicon 926 -515 926 -515 0 3
rlabel polysilicon 933 -509 933 -509 0 1
rlabel polysilicon 933 -515 933 -515 0 3
rlabel polysilicon 940 -509 940 -509 0 1
rlabel polysilicon 940 -515 940 -515 0 3
rlabel polysilicon 947 -509 947 -509 0 1
rlabel polysilicon 947 -515 947 -515 0 3
rlabel polysilicon 954 -509 954 -509 0 1
rlabel polysilicon 954 -515 954 -515 0 3
rlabel polysilicon 961 -509 961 -509 0 1
rlabel polysilicon 961 -515 961 -515 0 3
rlabel polysilicon 968 -509 968 -509 0 1
rlabel polysilicon 968 -515 968 -515 0 3
rlabel polysilicon 975 -509 975 -509 0 1
rlabel polysilicon 975 -515 975 -515 0 3
rlabel polysilicon 982 -509 982 -509 0 1
rlabel polysilicon 982 -515 982 -515 0 3
rlabel polysilicon 989 -509 989 -509 0 1
rlabel polysilicon 989 -515 989 -515 0 3
rlabel polysilicon 996 -509 996 -509 0 1
rlabel polysilicon 996 -515 996 -515 0 3
rlabel polysilicon 1003 -509 1003 -509 0 1
rlabel polysilicon 1003 -515 1003 -515 0 3
rlabel polysilicon 1010 -509 1010 -509 0 1
rlabel polysilicon 1010 -515 1010 -515 0 3
rlabel polysilicon 1017 -509 1017 -509 0 1
rlabel polysilicon 1017 -515 1017 -515 0 3
rlabel polysilicon 1024 -509 1024 -509 0 1
rlabel polysilicon 1024 -515 1024 -515 0 3
rlabel polysilicon 1031 -509 1031 -509 0 1
rlabel polysilicon 1031 -515 1031 -515 0 3
rlabel polysilicon 1038 -509 1038 -509 0 1
rlabel polysilicon 1038 -515 1038 -515 0 3
rlabel polysilicon 1045 -509 1045 -509 0 1
rlabel polysilicon 1045 -515 1045 -515 0 3
rlabel polysilicon 1052 -509 1052 -509 0 1
rlabel polysilicon 1052 -515 1052 -515 0 3
rlabel polysilicon 1059 -509 1059 -509 0 1
rlabel polysilicon 1059 -515 1059 -515 0 3
rlabel polysilicon 1066 -509 1066 -509 0 1
rlabel polysilicon 1066 -515 1066 -515 0 3
rlabel polysilicon 1073 -509 1073 -509 0 1
rlabel polysilicon 1073 -515 1073 -515 0 3
rlabel polysilicon 1080 -509 1080 -509 0 1
rlabel polysilicon 1080 -515 1080 -515 0 3
rlabel polysilicon 1087 -509 1087 -509 0 1
rlabel polysilicon 1087 -515 1087 -515 0 3
rlabel polysilicon 1094 -509 1094 -509 0 1
rlabel polysilicon 1094 -515 1094 -515 0 3
rlabel polysilicon 1101 -509 1101 -509 0 1
rlabel polysilicon 1101 -515 1101 -515 0 3
rlabel polysilicon 1108 -509 1108 -509 0 1
rlabel polysilicon 1108 -515 1108 -515 0 3
rlabel polysilicon 1115 -509 1115 -509 0 1
rlabel polysilicon 1115 -515 1115 -515 0 3
rlabel polysilicon 1122 -509 1122 -509 0 1
rlabel polysilicon 1122 -515 1122 -515 0 3
rlabel polysilicon 2 -608 2 -608 0 1
rlabel polysilicon 2 -614 2 -614 0 3
rlabel polysilicon 9 -608 9 -608 0 1
rlabel polysilicon 9 -614 9 -614 0 3
rlabel polysilicon 16 -608 16 -608 0 1
rlabel polysilicon 16 -614 16 -614 0 3
rlabel polysilicon 23 -608 23 -608 0 1
rlabel polysilicon 23 -614 23 -614 0 3
rlabel polysilicon 30 -608 30 -608 0 1
rlabel polysilicon 30 -614 30 -614 0 3
rlabel polysilicon 37 -608 37 -608 0 1
rlabel polysilicon 40 -614 40 -614 0 4
rlabel polysilicon 44 -608 44 -608 0 1
rlabel polysilicon 44 -614 44 -614 0 3
rlabel polysilicon 51 -608 51 -608 0 1
rlabel polysilicon 51 -614 51 -614 0 3
rlabel polysilicon 58 -608 58 -608 0 1
rlabel polysilicon 58 -614 58 -614 0 3
rlabel polysilicon 61 -614 61 -614 0 4
rlabel polysilicon 65 -608 65 -608 0 1
rlabel polysilicon 65 -614 65 -614 0 3
rlabel polysilicon 68 -614 68 -614 0 4
rlabel polysilicon 72 -608 72 -608 0 1
rlabel polysilicon 75 -608 75 -608 0 2
rlabel polysilicon 72 -614 72 -614 0 3
rlabel polysilicon 75 -614 75 -614 0 4
rlabel polysilicon 79 -608 79 -608 0 1
rlabel polysilicon 79 -614 79 -614 0 3
rlabel polysilicon 86 -608 86 -608 0 1
rlabel polysilicon 86 -614 86 -614 0 3
rlabel polysilicon 93 -608 93 -608 0 1
rlabel polysilicon 93 -614 93 -614 0 3
rlabel polysilicon 100 -608 100 -608 0 1
rlabel polysilicon 100 -614 100 -614 0 3
rlabel polysilicon 107 -608 107 -608 0 1
rlabel polysilicon 107 -614 107 -614 0 3
rlabel polysilicon 114 -608 114 -608 0 1
rlabel polysilicon 114 -614 114 -614 0 3
rlabel polysilicon 121 -608 121 -608 0 1
rlabel polysilicon 121 -614 121 -614 0 3
rlabel polysilicon 128 -608 128 -608 0 1
rlabel polysilicon 128 -614 128 -614 0 3
rlabel polysilicon 135 -608 135 -608 0 1
rlabel polysilicon 135 -614 135 -614 0 3
rlabel polysilicon 142 -608 142 -608 0 1
rlabel polysilicon 145 -608 145 -608 0 2
rlabel polysilicon 142 -614 142 -614 0 3
rlabel polysilicon 145 -614 145 -614 0 4
rlabel polysilicon 149 -608 149 -608 0 1
rlabel polysilicon 149 -614 149 -614 0 3
rlabel polysilicon 156 -608 156 -608 0 1
rlabel polysilicon 156 -614 156 -614 0 3
rlabel polysilicon 163 -608 163 -608 0 1
rlabel polysilicon 163 -614 163 -614 0 3
rlabel polysilicon 170 -608 170 -608 0 1
rlabel polysilicon 170 -614 170 -614 0 3
rlabel polysilicon 177 -608 177 -608 0 1
rlabel polysilicon 177 -614 177 -614 0 3
rlabel polysilicon 184 -608 184 -608 0 1
rlabel polysilicon 187 -608 187 -608 0 2
rlabel polysilicon 184 -614 184 -614 0 3
rlabel polysilicon 187 -614 187 -614 0 4
rlabel polysilicon 191 -608 191 -608 0 1
rlabel polysilicon 191 -614 191 -614 0 3
rlabel polysilicon 198 -608 198 -608 0 1
rlabel polysilicon 198 -614 198 -614 0 3
rlabel polysilicon 205 -608 205 -608 0 1
rlabel polysilicon 205 -614 205 -614 0 3
rlabel polysilicon 212 -608 212 -608 0 1
rlabel polysilicon 212 -614 212 -614 0 3
rlabel polysilicon 219 -608 219 -608 0 1
rlabel polysilicon 219 -614 219 -614 0 3
rlabel polysilicon 226 -608 226 -608 0 1
rlabel polysilicon 226 -614 226 -614 0 3
rlabel polysilicon 233 -608 233 -608 0 1
rlabel polysilicon 233 -614 233 -614 0 3
rlabel polysilicon 240 -608 240 -608 0 1
rlabel polysilicon 240 -614 240 -614 0 3
rlabel polysilicon 247 -608 247 -608 0 1
rlabel polysilicon 247 -614 247 -614 0 3
rlabel polysilicon 254 -608 254 -608 0 1
rlabel polysilicon 254 -614 254 -614 0 3
rlabel polysilicon 261 -608 261 -608 0 1
rlabel polysilicon 261 -614 261 -614 0 3
rlabel polysilicon 268 -608 268 -608 0 1
rlabel polysilicon 268 -614 268 -614 0 3
rlabel polysilicon 275 -608 275 -608 0 1
rlabel polysilicon 278 -608 278 -608 0 2
rlabel polysilicon 275 -614 275 -614 0 3
rlabel polysilicon 278 -614 278 -614 0 4
rlabel polysilicon 282 -608 282 -608 0 1
rlabel polysilicon 282 -614 282 -614 0 3
rlabel polysilicon 289 -608 289 -608 0 1
rlabel polysilicon 289 -614 289 -614 0 3
rlabel polysilicon 296 -608 296 -608 0 1
rlabel polysilicon 296 -614 296 -614 0 3
rlabel polysilicon 303 -608 303 -608 0 1
rlabel polysilicon 303 -614 303 -614 0 3
rlabel polysilicon 310 -608 310 -608 0 1
rlabel polysilicon 310 -614 310 -614 0 3
rlabel polysilicon 317 -608 317 -608 0 1
rlabel polysilicon 317 -614 317 -614 0 3
rlabel polysilicon 324 -608 324 -608 0 1
rlabel polysilicon 324 -614 324 -614 0 3
rlabel polysilicon 331 -608 331 -608 0 1
rlabel polysilicon 334 -608 334 -608 0 2
rlabel polysilicon 331 -614 331 -614 0 3
rlabel polysilicon 334 -614 334 -614 0 4
rlabel polysilicon 338 -608 338 -608 0 1
rlabel polysilicon 338 -614 338 -614 0 3
rlabel polysilicon 345 -608 345 -608 0 1
rlabel polysilicon 345 -614 345 -614 0 3
rlabel polysilicon 352 -608 352 -608 0 1
rlabel polysilicon 352 -614 352 -614 0 3
rlabel polysilicon 359 -608 359 -608 0 1
rlabel polysilicon 359 -614 359 -614 0 3
rlabel polysilicon 366 -608 366 -608 0 1
rlabel polysilicon 366 -614 366 -614 0 3
rlabel polysilicon 373 -608 373 -608 0 1
rlabel polysilicon 373 -614 373 -614 0 3
rlabel polysilicon 380 -608 380 -608 0 1
rlabel polysilicon 383 -608 383 -608 0 2
rlabel polysilicon 380 -614 380 -614 0 3
rlabel polysilicon 383 -614 383 -614 0 4
rlabel polysilicon 387 -608 387 -608 0 1
rlabel polysilicon 390 -608 390 -608 0 2
rlabel polysilicon 387 -614 387 -614 0 3
rlabel polysilicon 390 -614 390 -614 0 4
rlabel polysilicon 394 -608 394 -608 0 1
rlabel polysilicon 394 -614 394 -614 0 3
rlabel polysilicon 401 -608 401 -608 0 1
rlabel polysilicon 404 -608 404 -608 0 2
rlabel polysilicon 404 -614 404 -614 0 4
rlabel polysilicon 408 -608 408 -608 0 1
rlabel polysilicon 408 -614 408 -614 0 3
rlabel polysilicon 415 -608 415 -608 0 1
rlabel polysilicon 418 -614 418 -614 0 4
rlabel polysilicon 422 -608 422 -608 0 1
rlabel polysilicon 425 -608 425 -608 0 2
rlabel polysilicon 422 -614 422 -614 0 3
rlabel polysilicon 425 -614 425 -614 0 4
rlabel polysilicon 429 -608 429 -608 0 1
rlabel polysilicon 429 -614 429 -614 0 3
rlabel polysilicon 436 -608 436 -608 0 1
rlabel polysilicon 436 -614 436 -614 0 3
rlabel polysilicon 443 -608 443 -608 0 1
rlabel polysilicon 443 -614 443 -614 0 3
rlabel polysilicon 450 -608 450 -608 0 1
rlabel polysilicon 453 -608 453 -608 0 2
rlabel polysilicon 450 -614 450 -614 0 3
rlabel polysilicon 453 -614 453 -614 0 4
rlabel polysilicon 457 -608 457 -608 0 1
rlabel polysilicon 460 -608 460 -608 0 2
rlabel polysilicon 457 -614 457 -614 0 3
rlabel polysilicon 460 -614 460 -614 0 4
rlabel polysilicon 464 -608 464 -608 0 1
rlabel polysilicon 467 -608 467 -608 0 2
rlabel polysilicon 464 -614 464 -614 0 3
rlabel polysilicon 467 -614 467 -614 0 4
rlabel polysilicon 471 -608 471 -608 0 1
rlabel polysilicon 471 -614 471 -614 0 3
rlabel polysilicon 478 -608 478 -608 0 1
rlabel polysilicon 478 -614 478 -614 0 3
rlabel polysilicon 485 -608 485 -608 0 1
rlabel polysilicon 485 -614 485 -614 0 3
rlabel polysilicon 492 -608 492 -608 0 1
rlabel polysilicon 492 -614 492 -614 0 3
rlabel polysilicon 499 -608 499 -608 0 1
rlabel polysilicon 499 -614 499 -614 0 3
rlabel polysilicon 506 -608 506 -608 0 1
rlabel polysilicon 506 -614 506 -614 0 3
rlabel polysilicon 513 -608 513 -608 0 1
rlabel polysilicon 513 -614 513 -614 0 3
rlabel polysilicon 520 -608 520 -608 0 1
rlabel polysilicon 523 -608 523 -608 0 2
rlabel polysilicon 520 -614 520 -614 0 3
rlabel polysilicon 523 -614 523 -614 0 4
rlabel polysilicon 527 -608 527 -608 0 1
rlabel polysilicon 527 -614 527 -614 0 3
rlabel polysilicon 534 -608 534 -608 0 1
rlabel polysilicon 534 -614 534 -614 0 3
rlabel polysilicon 541 -608 541 -608 0 1
rlabel polysilicon 544 -608 544 -608 0 2
rlabel polysilicon 541 -614 541 -614 0 3
rlabel polysilicon 544 -614 544 -614 0 4
rlabel polysilicon 548 -608 548 -608 0 1
rlabel polysilicon 551 -608 551 -608 0 2
rlabel polysilicon 548 -614 548 -614 0 3
rlabel polysilicon 551 -614 551 -614 0 4
rlabel polysilicon 555 -608 555 -608 0 1
rlabel polysilicon 555 -614 555 -614 0 3
rlabel polysilicon 562 -608 562 -608 0 1
rlabel polysilicon 565 -608 565 -608 0 2
rlabel polysilicon 562 -614 562 -614 0 3
rlabel polysilicon 565 -614 565 -614 0 4
rlabel polysilicon 569 -608 569 -608 0 1
rlabel polysilicon 569 -614 569 -614 0 3
rlabel polysilicon 576 -608 576 -608 0 1
rlabel polysilicon 576 -614 576 -614 0 3
rlabel polysilicon 583 -608 583 -608 0 1
rlabel polysilicon 583 -614 583 -614 0 3
rlabel polysilicon 586 -614 586 -614 0 4
rlabel polysilicon 590 -608 590 -608 0 1
rlabel polysilicon 590 -614 590 -614 0 3
rlabel polysilicon 597 -608 597 -608 0 1
rlabel polysilicon 597 -614 597 -614 0 3
rlabel polysilicon 604 -608 604 -608 0 1
rlabel polysilicon 604 -614 604 -614 0 3
rlabel polysilicon 611 -608 611 -608 0 1
rlabel polysilicon 611 -614 611 -614 0 3
rlabel polysilicon 618 -608 618 -608 0 1
rlabel polysilicon 621 -608 621 -608 0 2
rlabel polysilicon 618 -614 618 -614 0 3
rlabel polysilicon 621 -614 621 -614 0 4
rlabel polysilicon 625 -608 625 -608 0 1
rlabel polysilicon 628 -608 628 -608 0 2
rlabel polysilicon 625 -614 625 -614 0 3
rlabel polysilicon 628 -614 628 -614 0 4
rlabel polysilicon 632 -608 632 -608 0 1
rlabel polysilicon 632 -614 632 -614 0 3
rlabel polysilicon 639 -608 639 -608 0 1
rlabel polysilicon 639 -614 639 -614 0 3
rlabel polysilicon 646 -608 646 -608 0 1
rlabel polysilicon 646 -614 646 -614 0 3
rlabel polysilicon 653 -608 653 -608 0 1
rlabel polysilicon 653 -614 653 -614 0 3
rlabel polysilicon 660 -608 660 -608 0 1
rlabel polysilicon 660 -614 660 -614 0 3
rlabel polysilicon 667 -608 667 -608 0 1
rlabel polysilicon 667 -614 667 -614 0 3
rlabel polysilicon 674 -608 674 -608 0 1
rlabel polysilicon 674 -614 674 -614 0 3
rlabel polysilicon 681 -608 681 -608 0 1
rlabel polysilicon 681 -614 681 -614 0 3
rlabel polysilicon 688 -608 688 -608 0 1
rlabel polysilicon 688 -614 688 -614 0 3
rlabel polysilicon 695 -608 695 -608 0 1
rlabel polysilicon 695 -614 695 -614 0 3
rlabel polysilicon 702 -608 702 -608 0 1
rlabel polysilicon 702 -614 702 -614 0 3
rlabel polysilicon 709 -608 709 -608 0 1
rlabel polysilicon 709 -614 709 -614 0 3
rlabel polysilicon 716 -608 716 -608 0 1
rlabel polysilicon 716 -614 716 -614 0 3
rlabel polysilicon 723 -608 723 -608 0 1
rlabel polysilicon 723 -614 723 -614 0 3
rlabel polysilicon 730 -608 730 -608 0 1
rlabel polysilicon 730 -614 730 -614 0 3
rlabel polysilicon 737 -608 737 -608 0 1
rlabel polysilicon 737 -614 737 -614 0 3
rlabel polysilicon 744 -608 744 -608 0 1
rlabel polysilicon 744 -614 744 -614 0 3
rlabel polysilicon 751 -608 751 -608 0 1
rlabel polysilicon 751 -614 751 -614 0 3
rlabel polysilicon 758 -608 758 -608 0 1
rlabel polysilicon 758 -614 758 -614 0 3
rlabel polysilicon 765 -608 765 -608 0 1
rlabel polysilicon 765 -614 765 -614 0 3
rlabel polysilicon 772 -608 772 -608 0 1
rlabel polysilicon 772 -614 772 -614 0 3
rlabel polysilicon 779 -608 779 -608 0 1
rlabel polysilicon 779 -614 779 -614 0 3
rlabel polysilicon 786 -608 786 -608 0 1
rlabel polysilicon 786 -614 786 -614 0 3
rlabel polysilicon 793 -608 793 -608 0 1
rlabel polysilicon 793 -614 793 -614 0 3
rlabel polysilicon 800 -608 800 -608 0 1
rlabel polysilicon 800 -614 800 -614 0 3
rlabel polysilicon 807 -608 807 -608 0 1
rlabel polysilicon 807 -614 807 -614 0 3
rlabel polysilicon 814 -608 814 -608 0 1
rlabel polysilicon 814 -614 814 -614 0 3
rlabel polysilicon 821 -608 821 -608 0 1
rlabel polysilicon 821 -614 821 -614 0 3
rlabel polysilicon 828 -608 828 -608 0 1
rlabel polysilicon 828 -614 828 -614 0 3
rlabel polysilicon 835 -608 835 -608 0 1
rlabel polysilicon 835 -614 835 -614 0 3
rlabel polysilicon 842 -608 842 -608 0 1
rlabel polysilicon 842 -614 842 -614 0 3
rlabel polysilicon 849 -608 849 -608 0 1
rlabel polysilicon 849 -614 849 -614 0 3
rlabel polysilicon 856 -608 856 -608 0 1
rlabel polysilicon 856 -614 856 -614 0 3
rlabel polysilicon 863 -608 863 -608 0 1
rlabel polysilicon 863 -614 863 -614 0 3
rlabel polysilicon 870 -608 870 -608 0 1
rlabel polysilicon 870 -614 870 -614 0 3
rlabel polysilicon 877 -608 877 -608 0 1
rlabel polysilicon 877 -614 877 -614 0 3
rlabel polysilicon 884 -608 884 -608 0 1
rlabel polysilicon 884 -614 884 -614 0 3
rlabel polysilicon 891 -608 891 -608 0 1
rlabel polysilicon 891 -614 891 -614 0 3
rlabel polysilicon 898 -608 898 -608 0 1
rlabel polysilicon 898 -614 898 -614 0 3
rlabel polysilicon 905 -608 905 -608 0 1
rlabel polysilicon 905 -614 905 -614 0 3
rlabel polysilicon 912 -608 912 -608 0 1
rlabel polysilicon 912 -614 912 -614 0 3
rlabel polysilicon 919 -608 919 -608 0 1
rlabel polysilicon 919 -614 919 -614 0 3
rlabel polysilicon 926 -608 926 -608 0 1
rlabel polysilicon 926 -614 926 -614 0 3
rlabel polysilicon 933 -608 933 -608 0 1
rlabel polysilicon 933 -614 933 -614 0 3
rlabel polysilicon 940 -608 940 -608 0 1
rlabel polysilicon 940 -614 940 -614 0 3
rlabel polysilicon 947 -608 947 -608 0 1
rlabel polysilicon 947 -614 947 -614 0 3
rlabel polysilicon 954 -608 954 -608 0 1
rlabel polysilicon 954 -614 954 -614 0 3
rlabel polysilicon 961 -608 961 -608 0 1
rlabel polysilicon 961 -614 961 -614 0 3
rlabel polysilicon 968 -608 968 -608 0 1
rlabel polysilicon 968 -614 968 -614 0 3
rlabel polysilicon 975 -608 975 -608 0 1
rlabel polysilicon 975 -614 975 -614 0 3
rlabel polysilicon 982 -608 982 -608 0 1
rlabel polysilicon 982 -614 982 -614 0 3
rlabel polysilicon 989 -608 989 -608 0 1
rlabel polysilicon 989 -614 989 -614 0 3
rlabel polysilicon 996 -608 996 -608 0 1
rlabel polysilicon 996 -614 996 -614 0 3
rlabel polysilicon 1003 -608 1003 -608 0 1
rlabel polysilicon 1003 -614 1003 -614 0 3
rlabel polysilicon 1010 -608 1010 -608 0 1
rlabel polysilicon 1010 -614 1010 -614 0 3
rlabel polysilicon 1017 -608 1017 -608 0 1
rlabel polysilicon 1017 -614 1017 -614 0 3
rlabel polysilicon 1024 -608 1024 -608 0 1
rlabel polysilicon 1024 -614 1024 -614 0 3
rlabel polysilicon 1031 -608 1031 -608 0 1
rlabel polysilicon 1031 -614 1031 -614 0 3
rlabel polysilicon 1038 -608 1038 -608 0 1
rlabel polysilicon 1038 -614 1038 -614 0 3
rlabel polysilicon 1045 -608 1045 -608 0 1
rlabel polysilicon 1045 -614 1045 -614 0 3
rlabel polysilicon 1052 -608 1052 -608 0 1
rlabel polysilicon 1052 -614 1052 -614 0 3
rlabel polysilicon 1059 -608 1059 -608 0 1
rlabel polysilicon 1059 -614 1059 -614 0 3
rlabel polysilicon 1066 -608 1066 -608 0 1
rlabel polysilicon 1066 -614 1066 -614 0 3
rlabel polysilicon 1073 -608 1073 -608 0 1
rlabel polysilicon 1073 -614 1073 -614 0 3
rlabel polysilicon 1080 -608 1080 -608 0 1
rlabel polysilicon 1083 -614 1083 -614 0 4
rlabel polysilicon 1087 -608 1087 -608 0 1
rlabel polysilicon 1087 -614 1087 -614 0 3
rlabel polysilicon 2 -717 2 -717 0 1
rlabel polysilicon 2 -723 2 -723 0 3
rlabel polysilicon 9 -717 9 -717 0 1
rlabel polysilicon 9 -723 9 -723 0 3
rlabel polysilicon 16 -717 16 -717 0 1
rlabel polysilicon 16 -723 16 -723 0 3
rlabel polysilicon 23 -717 23 -717 0 1
rlabel polysilicon 23 -723 23 -723 0 3
rlabel polysilicon 30 -717 30 -717 0 1
rlabel polysilicon 30 -723 30 -723 0 3
rlabel polysilicon 37 -717 37 -717 0 1
rlabel polysilicon 37 -723 37 -723 0 3
rlabel polysilicon 44 -717 44 -717 0 1
rlabel polysilicon 47 -717 47 -717 0 2
rlabel polysilicon 44 -723 44 -723 0 3
rlabel polysilicon 51 -717 51 -717 0 1
rlabel polysilicon 51 -723 51 -723 0 3
rlabel polysilicon 58 -717 58 -717 0 1
rlabel polysilicon 61 -717 61 -717 0 2
rlabel polysilicon 58 -723 58 -723 0 3
rlabel polysilicon 61 -723 61 -723 0 4
rlabel polysilicon 65 -717 65 -717 0 1
rlabel polysilicon 65 -723 65 -723 0 3
rlabel polysilicon 72 -717 72 -717 0 1
rlabel polysilicon 72 -723 72 -723 0 3
rlabel polysilicon 79 -717 79 -717 0 1
rlabel polysilicon 79 -723 79 -723 0 3
rlabel polysilicon 86 -717 86 -717 0 1
rlabel polysilicon 89 -717 89 -717 0 2
rlabel polysilicon 89 -723 89 -723 0 4
rlabel polysilicon 93 -717 93 -717 0 1
rlabel polysilicon 93 -723 93 -723 0 3
rlabel polysilicon 100 -717 100 -717 0 1
rlabel polysilicon 100 -723 100 -723 0 3
rlabel polysilicon 107 -717 107 -717 0 1
rlabel polysilicon 110 -717 110 -717 0 2
rlabel polysilicon 107 -723 107 -723 0 3
rlabel polysilicon 110 -723 110 -723 0 4
rlabel polysilicon 114 -717 114 -717 0 1
rlabel polysilicon 114 -723 114 -723 0 3
rlabel polysilicon 121 -717 121 -717 0 1
rlabel polysilicon 121 -723 121 -723 0 3
rlabel polysilicon 128 -717 128 -717 0 1
rlabel polysilicon 128 -723 128 -723 0 3
rlabel polysilicon 135 -717 135 -717 0 1
rlabel polysilicon 135 -723 135 -723 0 3
rlabel polysilicon 142 -717 142 -717 0 1
rlabel polysilicon 142 -723 142 -723 0 3
rlabel polysilicon 149 -717 149 -717 0 1
rlabel polysilicon 149 -723 149 -723 0 3
rlabel polysilicon 156 -717 156 -717 0 1
rlabel polysilicon 156 -723 156 -723 0 3
rlabel polysilicon 163 -717 163 -717 0 1
rlabel polysilicon 163 -723 163 -723 0 3
rlabel polysilicon 170 -717 170 -717 0 1
rlabel polysilicon 170 -723 170 -723 0 3
rlabel polysilicon 177 -717 177 -717 0 1
rlabel polysilicon 177 -723 177 -723 0 3
rlabel polysilicon 184 -717 184 -717 0 1
rlabel polysilicon 184 -723 184 -723 0 3
rlabel polysilicon 191 -717 191 -717 0 1
rlabel polysilicon 191 -723 191 -723 0 3
rlabel polysilicon 194 -723 194 -723 0 4
rlabel polysilicon 198 -717 198 -717 0 1
rlabel polysilicon 198 -723 198 -723 0 3
rlabel polysilicon 205 -717 205 -717 0 1
rlabel polysilicon 205 -723 205 -723 0 3
rlabel polysilicon 212 -717 212 -717 0 1
rlabel polysilicon 212 -723 212 -723 0 3
rlabel polysilicon 219 -717 219 -717 0 1
rlabel polysilicon 219 -723 219 -723 0 3
rlabel polysilicon 226 -717 226 -717 0 1
rlabel polysilicon 229 -717 229 -717 0 2
rlabel polysilicon 226 -723 226 -723 0 3
rlabel polysilicon 233 -717 233 -717 0 1
rlabel polysilicon 236 -717 236 -717 0 2
rlabel polysilicon 233 -723 233 -723 0 3
rlabel polysilicon 240 -717 240 -717 0 1
rlabel polysilicon 240 -723 240 -723 0 3
rlabel polysilicon 247 -717 247 -717 0 1
rlabel polysilicon 247 -723 247 -723 0 3
rlabel polysilicon 254 -717 254 -717 0 1
rlabel polysilicon 254 -723 254 -723 0 3
rlabel polysilicon 261 -717 261 -717 0 1
rlabel polysilicon 261 -723 261 -723 0 3
rlabel polysilicon 268 -717 268 -717 0 1
rlabel polysilicon 268 -723 268 -723 0 3
rlabel polysilicon 275 -717 275 -717 0 1
rlabel polysilicon 275 -723 275 -723 0 3
rlabel polysilicon 282 -717 282 -717 0 1
rlabel polysilicon 282 -723 282 -723 0 3
rlabel polysilicon 289 -717 289 -717 0 1
rlabel polysilicon 289 -723 289 -723 0 3
rlabel polysilicon 296 -717 296 -717 0 1
rlabel polysilicon 296 -723 296 -723 0 3
rlabel polysilicon 303 -717 303 -717 0 1
rlabel polysilicon 303 -723 303 -723 0 3
rlabel polysilicon 310 -717 310 -717 0 1
rlabel polysilicon 310 -723 310 -723 0 3
rlabel polysilicon 317 -717 317 -717 0 1
rlabel polysilicon 317 -723 317 -723 0 3
rlabel polysilicon 324 -717 324 -717 0 1
rlabel polysilicon 324 -723 324 -723 0 3
rlabel polysilicon 331 -717 331 -717 0 1
rlabel polysilicon 331 -723 331 -723 0 3
rlabel polysilicon 338 -717 338 -717 0 1
rlabel polysilicon 338 -723 338 -723 0 3
rlabel polysilicon 345 -717 345 -717 0 1
rlabel polysilicon 345 -723 345 -723 0 3
rlabel polysilicon 352 -717 352 -717 0 1
rlabel polysilicon 352 -723 352 -723 0 3
rlabel polysilicon 359 -717 359 -717 0 1
rlabel polysilicon 359 -723 359 -723 0 3
rlabel polysilicon 366 -717 366 -717 0 1
rlabel polysilicon 369 -717 369 -717 0 2
rlabel polysilicon 366 -723 366 -723 0 3
rlabel polysilicon 369 -723 369 -723 0 4
rlabel polysilicon 373 -717 373 -717 0 1
rlabel polysilicon 373 -723 373 -723 0 3
rlabel polysilicon 380 -717 380 -717 0 1
rlabel polysilicon 383 -717 383 -717 0 2
rlabel polysilicon 380 -723 380 -723 0 3
rlabel polysilicon 383 -723 383 -723 0 4
rlabel polysilicon 387 -717 387 -717 0 1
rlabel polysilicon 387 -723 387 -723 0 3
rlabel polysilicon 390 -723 390 -723 0 4
rlabel polysilicon 394 -717 394 -717 0 1
rlabel polysilicon 394 -723 394 -723 0 3
rlabel polysilicon 404 -717 404 -717 0 2
rlabel polysilicon 404 -723 404 -723 0 4
rlabel polysilicon 408 -717 408 -717 0 1
rlabel polysilicon 408 -723 408 -723 0 3
rlabel polysilicon 415 -717 415 -717 0 1
rlabel polysilicon 418 -717 418 -717 0 2
rlabel polysilicon 415 -723 415 -723 0 3
rlabel polysilicon 422 -717 422 -717 0 1
rlabel polysilicon 422 -723 422 -723 0 3
rlabel polysilicon 429 -717 429 -717 0 1
rlabel polysilicon 432 -717 432 -717 0 2
rlabel polysilicon 429 -723 429 -723 0 3
rlabel polysilicon 432 -723 432 -723 0 4
rlabel polysilicon 436 -717 436 -717 0 1
rlabel polysilicon 436 -723 436 -723 0 3
rlabel polysilicon 443 -717 443 -717 0 1
rlabel polysilicon 446 -717 446 -717 0 2
rlabel polysilicon 443 -723 443 -723 0 3
rlabel polysilicon 446 -723 446 -723 0 4
rlabel polysilicon 450 -717 450 -717 0 1
rlabel polysilicon 450 -723 450 -723 0 3
rlabel polysilicon 457 -717 457 -717 0 1
rlabel polysilicon 457 -723 457 -723 0 3
rlabel polysilicon 464 -717 464 -717 0 1
rlabel polysilicon 464 -723 464 -723 0 3
rlabel polysilicon 471 -717 471 -717 0 1
rlabel polysilicon 471 -723 471 -723 0 3
rlabel polysilicon 478 -717 478 -717 0 1
rlabel polysilicon 478 -723 478 -723 0 3
rlabel polysilicon 485 -717 485 -717 0 1
rlabel polysilicon 485 -723 485 -723 0 3
rlabel polysilicon 492 -717 492 -717 0 1
rlabel polysilicon 492 -723 492 -723 0 3
rlabel polysilicon 499 -717 499 -717 0 1
rlabel polysilicon 502 -717 502 -717 0 2
rlabel polysilicon 499 -723 499 -723 0 3
rlabel polysilicon 502 -723 502 -723 0 4
rlabel polysilicon 506 -717 506 -717 0 1
rlabel polysilicon 506 -723 506 -723 0 3
rlabel polysilicon 513 -717 513 -717 0 1
rlabel polysilicon 513 -723 513 -723 0 3
rlabel polysilicon 520 -717 520 -717 0 1
rlabel polysilicon 520 -723 520 -723 0 3
rlabel polysilicon 527 -717 527 -717 0 1
rlabel polysilicon 527 -723 527 -723 0 3
rlabel polysilicon 534 -717 534 -717 0 1
rlabel polysilicon 534 -723 534 -723 0 3
rlabel polysilicon 541 -717 541 -717 0 1
rlabel polysilicon 541 -723 541 -723 0 3
rlabel polysilicon 548 -717 548 -717 0 1
rlabel polysilicon 548 -723 548 -723 0 3
rlabel polysilicon 555 -717 555 -717 0 1
rlabel polysilicon 558 -717 558 -717 0 2
rlabel polysilicon 558 -723 558 -723 0 4
rlabel polysilicon 562 -717 562 -717 0 1
rlabel polysilicon 565 -717 565 -717 0 2
rlabel polysilicon 562 -723 562 -723 0 3
rlabel polysilicon 565 -723 565 -723 0 4
rlabel polysilicon 569 -717 569 -717 0 1
rlabel polysilicon 569 -723 569 -723 0 3
rlabel polysilicon 576 -717 576 -717 0 1
rlabel polysilicon 576 -723 576 -723 0 3
rlabel polysilicon 583 -717 583 -717 0 1
rlabel polysilicon 586 -717 586 -717 0 2
rlabel polysilicon 583 -723 583 -723 0 3
rlabel polysilicon 586 -723 586 -723 0 4
rlabel polysilicon 590 -717 590 -717 0 1
rlabel polysilicon 590 -723 590 -723 0 3
rlabel polysilicon 597 -717 597 -717 0 1
rlabel polysilicon 597 -723 597 -723 0 3
rlabel polysilicon 604 -717 604 -717 0 1
rlabel polysilicon 604 -723 604 -723 0 3
rlabel polysilicon 611 -717 611 -717 0 1
rlabel polysilicon 611 -723 611 -723 0 3
rlabel polysilicon 618 -717 618 -717 0 1
rlabel polysilicon 618 -723 618 -723 0 3
rlabel polysilicon 625 -717 625 -717 0 1
rlabel polysilicon 625 -723 625 -723 0 3
rlabel polysilicon 632 -717 632 -717 0 1
rlabel polysilicon 635 -717 635 -717 0 2
rlabel polysilicon 632 -723 632 -723 0 3
rlabel polysilicon 635 -723 635 -723 0 4
rlabel polysilicon 639 -717 639 -717 0 1
rlabel polysilicon 639 -723 639 -723 0 3
rlabel polysilicon 646 -717 646 -717 0 1
rlabel polysilicon 649 -717 649 -717 0 2
rlabel polysilicon 649 -723 649 -723 0 4
rlabel polysilicon 653 -717 653 -717 0 1
rlabel polysilicon 656 -717 656 -717 0 2
rlabel polysilicon 653 -723 653 -723 0 3
rlabel polysilicon 656 -723 656 -723 0 4
rlabel polysilicon 660 -717 660 -717 0 1
rlabel polysilicon 660 -723 660 -723 0 3
rlabel polysilicon 667 -717 667 -717 0 1
rlabel polysilicon 667 -723 667 -723 0 3
rlabel polysilicon 674 -717 674 -717 0 1
rlabel polysilicon 674 -723 674 -723 0 3
rlabel polysilicon 681 -717 681 -717 0 1
rlabel polysilicon 681 -723 681 -723 0 3
rlabel polysilicon 688 -717 688 -717 0 1
rlabel polysilicon 688 -723 688 -723 0 3
rlabel polysilicon 695 -717 695 -717 0 1
rlabel polysilicon 695 -723 695 -723 0 3
rlabel polysilicon 702 -717 702 -717 0 1
rlabel polysilicon 702 -723 702 -723 0 3
rlabel polysilicon 709 -717 709 -717 0 1
rlabel polysilicon 709 -723 709 -723 0 3
rlabel polysilicon 716 -717 716 -717 0 1
rlabel polysilicon 716 -723 716 -723 0 3
rlabel polysilicon 723 -717 723 -717 0 1
rlabel polysilicon 726 -717 726 -717 0 2
rlabel polysilicon 723 -723 723 -723 0 3
rlabel polysilicon 726 -723 726 -723 0 4
rlabel polysilicon 730 -717 730 -717 0 1
rlabel polysilicon 733 -717 733 -717 0 2
rlabel polysilicon 730 -723 730 -723 0 3
rlabel polysilicon 733 -723 733 -723 0 4
rlabel polysilicon 737 -717 737 -717 0 1
rlabel polysilicon 737 -723 737 -723 0 3
rlabel polysilicon 744 -717 744 -717 0 1
rlabel polysilicon 744 -723 744 -723 0 3
rlabel polysilicon 751 -717 751 -717 0 1
rlabel polysilicon 751 -723 751 -723 0 3
rlabel polysilicon 758 -717 758 -717 0 1
rlabel polysilicon 758 -723 758 -723 0 3
rlabel polysilicon 765 -717 765 -717 0 1
rlabel polysilicon 765 -723 765 -723 0 3
rlabel polysilicon 772 -717 772 -717 0 1
rlabel polysilicon 772 -723 772 -723 0 3
rlabel polysilicon 779 -717 779 -717 0 1
rlabel polysilicon 779 -723 779 -723 0 3
rlabel polysilicon 786 -717 786 -717 0 1
rlabel polysilicon 786 -723 786 -723 0 3
rlabel polysilicon 793 -717 793 -717 0 1
rlabel polysilicon 793 -723 793 -723 0 3
rlabel polysilicon 800 -717 800 -717 0 1
rlabel polysilicon 800 -723 800 -723 0 3
rlabel polysilicon 810 -717 810 -717 0 2
rlabel polysilicon 807 -723 807 -723 0 3
rlabel polysilicon 814 -717 814 -717 0 1
rlabel polysilicon 814 -723 814 -723 0 3
rlabel polysilicon 821 -717 821 -717 0 1
rlabel polysilicon 821 -723 821 -723 0 3
rlabel polysilicon 828 -717 828 -717 0 1
rlabel polysilicon 828 -723 828 -723 0 3
rlabel polysilicon 835 -717 835 -717 0 1
rlabel polysilicon 835 -723 835 -723 0 3
rlabel polysilicon 842 -717 842 -717 0 1
rlabel polysilicon 842 -723 842 -723 0 3
rlabel polysilicon 849 -717 849 -717 0 1
rlabel polysilicon 849 -723 849 -723 0 3
rlabel polysilicon 856 -717 856 -717 0 1
rlabel polysilicon 856 -723 856 -723 0 3
rlabel polysilicon 863 -717 863 -717 0 1
rlabel polysilicon 863 -723 863 -723 0 3
rlabel polysilicon 870 -717 870 -717 0 1
rlabel polysilicon 870 -723 870 -723 0 3
rlabel polysilicon 877 -717 877 -717 0 1
rlabel polysilicon 877 -723 877 -723 0 3
rlabel polysilicon 884 -717 884 -717 0 1
rlabel polysilicon 884 -723 884 -723 0 3
rlabel polysilicon 891 -717 891 -717 0 1
rlabel polysilicon 891 -723 891 -723 0 3
rlabel polysilicon 898 -717 898 -717 0 1
rlabel polysilicon 898 -723 898 -723 0 3
rlabel polysilicon 905 -717 905 -717 0 1
rlabel polysilicon 905 -723 905 -723 0 3
rlabel polysilicon 912 -717 912 -717 0 1
rlabel polysilicon 912 -723 912 -723 0 3
rlabel polysilicon 919 -717 919 -717 0 1
rlabel polysilicon 919 -723 919 -723 0 3
rlabel polysilicon 926 -717 926 -717 0 1
rlabel polysilicon 926 -723 926 -723 0 3
rlabel polysilicon 933 -717 933 -717 0 1
rlabel polysilicon 933 -723 933 -723 0 3
rlabel polysilicon 940 -717 940 -717 0 1
rlabel polysilicon 940 -723 940 -723 0 3
rlabel polysilicon 947 -717 947 -717 0 1
rlabel polysilicon 947 -723 947 -723 0 3
rlabel polysilicon 954 -717 954 -717 0 1
rlabel polysilicon 954 -723 954 -723 0 3
rlabel polysilicon 961 -717 961 -717 0 1
rlabel polysilicon 961 -723 961 -723 0 3
rlabel polysilicon 968 -717 968 -717 0 1
rlabel polysilicon 968 -723 968 -723 0 3
rlabel polysilicon 975 -717 975 -717 0 1
rlabel polysilicon 975 -723 975 -723 0 3
rlabel polysilicon 982 -717 982 -717 0 1
rlabel polysilicon 982 -723 982 -723 0 3
rlabel polysilicon 989 -717 989 -717 0 1
rlabel polysilicon 989 -723 989 -723 0 3
rlabel polysilicon 996 -717 996 -717 0 1
rlabel polysilicon 996 -723 996 -723 0 3
rlabel polysilicon 1003 -717 1003 -717 0 1
rlabel polysilicon 1003 -723 1003 -723 0 3
rlabel polysilicon 1010 -717 1010 -717 0 1
rlabel polysilicon 1010 -723 1010 -723 0 3
rlabel polysilicon 1017 -717 1017 -717 0 1
rlabel polysilicon 1017 -723 1017 -723 0 3
rlabel polysilicon 1024 -717 1024 -717 0 1
rlabel polysilicon 1024 -723 1024 -723 0 3
rlabel polysilicon 1031 -717 1031 -717 0 1
rlabel polysilicon 1031 -723 1031 -723 0 3
rlabel polysilicon 1038 -717 1038 -717 0 1
rlabel polysilicon 1038 -723 1038 -723 0 3
rlabel polysilicon 1045 -717 1045 -717 0 1
rlabel polysilicon 1045 -723 1045 -723 0 3
rlabel polysilicon 1052 -717 1052 -717 0 1
rlabel polysilicon 1052 -723 1052 -723 0 3
rlabel polysilicon 1059 -717 1059 -717 0 1
rlabel polysilicon 1059 -723 1059 -723 0 3
rlabel polysilicon 1066 -717 1066 -717 0 1
rlabel polysilicon 1066 -723 1066 -723 0 3
rlabel polysilicon 1073 -717 1073 -717 0 1
rlabel polysilicon 1073 -723 1073 -723 0 3
rlabel polysilicon 1080 -717 1080 -717 0 1
rlabel polysilicon 1080 -723 1080 -723 0 3
rlabel polysilicon 1087 -717 1087 -717 0 1
rlabel polysilicon 1087 -723 1087 -723 0 3
rlabel polysilicon 1094 -717 1094 -717 0 1
rlabel polysilicon 1094 -723 1094 -723 0 3
rlabel polysilicon 1101 -717 1101 -717 0 1
rlabel polysilicon 1101 -723 1101 -723 0 3
rlabel polysilicon 1108 -717 1108 -717 0 1
rlabel polysilicon 1108 -723 1108 -723 0 3
rlabel polysilicon 1115 -717 1115 -717 0 1
rlabel polysilicon 1115 -723 1115 -723 0 3
rlabel polysilicon 1122 -717 1122 -717 0 1
rlabel polysilicon 1122 -723 1122 -723 0 3
rlabel polysilicon 1129 -717 1129 -717 0 1
rlabel polysilicon 1129 -723 1129 -723 0 3
rlabel polysilicon 1136 -717 1136 -717 0 1
rlabel polysilicon 1136 -723 1136 -723 0 3
rlabel polysilicon 1143 -717 1143 -717 0 1
rlabel polysilicon 1143 -723 1143 -723 0 3
rlabel polysilicon 1150 -717 1150 -717 0 1
rlabel polysilicon 1150 -723 1150 -723 0 3
rlabel polysilicon 1157 -717 1157 -717 0 1
rlabel polysilicon 1157 -723 1157 -723 0 3
rlabel polysilicon 1164 -717 1164 -717 0 1
rlabel polysilicon 1164 -723 1164 -723 0 3
rlabel polysilicon 1171 -717 1171 -717 0 1
rlabel polysilicon 1171 -723 1171 -723 0 3
rlabel polysilicon 1178 -717 1178 -717 0 1
rlabel polysilicon 1178 -723 1178 -723 0 3
rlabel polysilicon 1185 -717 1185 -717 0 1
rlabel polysilicon 1185 -723 1185 -723 0 3
rlabel polysilicon 1192 -717 1192 -717 0 1
rlabel polysilicon 1192 -723 1192 -723 0 3
rlabel polysilicon 1199 -717 1199 -717 0 1
rlabel polysilicon 1199 -723 1199 -723 0 3
rlabel polysilicon 1206 -717 1206 -717 0 1
rlabel polysilicon 1206 -723 1206 -723 0 3
rlabel polysilicon 1213 -717 1213 -717 0 1
rlabel polysilicon 1216 -717 1216 -717 0 2
rlabel polysilicon 1213 -723 1213 -723 0 3
rlabel polysilicon 1360 -717 1360 -717 0 1
rlabel polysilicon 1360 -723 1360 -723 0 3
rlabel polysilicon 2 -834 2 -834 0 1
rlabel polysilicon 2 -840 2 -840 0 3
rlabel polysilicon 9 -834 9 -834 0 1
rlabel polysilicon 9 -840 9 -840 0 3
rlabel polysilicon 16 -834 16 -834 0 1
rlabel polysilicon 16 -840 16 -840 0 3
rlabel polysilicon 23 -840 23 -840 0 3
rlabel polysilicon 26 -840 26 -840 0 4
rlabel polysilicon 33 -834 33 -834 0 2
rlabel polysilicon 30 -840 30 -840 0 3
rlabel polysilicon 33 -840 33 -840 0 4
rlabel polysilicon 37 -834 37 -834 0 1
rlabel polysilicon 37 -840 37 -840 0 3
rlabel polysilicon 44 -834 44 -834 0 1
rlabel polysilicon 44 -840 44 -840 0 3
rlabel polysilicon 51 -834 51 -834 0 1
rlabel polysilicon 51 -840 51 -840 0 3
rlabel polysilicon 58 -834 58 -834 0 1
rlabel polysilicon 58 -840 58 -840 0 3
rlabel polysilicon 65 -834 65 -834 0 1
rlabel polysilicon 65 -840 65 -840 0 3
rlabel polysilicon 72 -834 72 -834 0 1
rlabel polysilicon 75 -834 75 -834 0 2
rlabel polysilicon 72 -840 72 -840 0 3
rlabel polysilicon 75 -840 75 -840 0 4
rlabel polysilicon 79 -834 79 -834 0 1
rlabel polysilicon 79 -840 79 -840 0 3
rlabel polysilicon 86 -834 86 -834 0 1
rlabel polysilicon 89 -834 89 -834 0 2
rlabel polysilicon 86 -840 86 -840 0 3
rlabel polysilicon 89 -840 89 -840 0 4
rlabel polysilicon 93 -834 93 -834 0 1
rlabel polysilicon 93 -840 93 -840 0 3
rlabel polysilicon 100 -834 100 -834 0 1
rlabel polysilicon 100 -840 100 -840 0 3
rlabel polysilicon 107 -834 107 -834 0 1
rlabel polysilicon 107 -840 107 -840 0 3
rlabel polysilicon 114 -834 114 -834 0 1
rlabel polysilicon 114 -840 114 -840 0 3
rlabel polysilicon 121 -834 121 -834 0 1
rlabel polysilicon 121 -840 121 -840 0 3
rlabel polysilicon 128 -834 128 -834 0 1
rlabel polysilicon 131 -834 131 -834 0 2
rlabel polysilicon 131 -840 131 -840 0 4
rlabel polysilicon 135 -834 135 -834 0 1
rlabel polysilicon 135 -840 135 -840 0 3
rlabel polysilicon 142 -834 142 -834 0 1
rlabel polysilicon 142 -840 142 -840 0 3
rlabel polysilicon 149 -834 149 -834 0 1
rlabel polysilicon 149 -840 149 -840 0 3
rlabel polysilicon 156 -834 156 -834 0 1
rlabel polysilicon 156 -840 156 -840 0 3
rlabel polysilicon 163 -834 163 -834 0 1
rlabel polysilicon 163 -840 163 -840 0 3
rlabel polysilicon 170 -834 170 -834 0 1
rlabel polysilicon 170 -840 170 -840 0 3
rlabel polysilicon 177 -834 177 -834 0 1
rlabel polysilicon 180 -840 180 -840 0 4
rlabel polysilicon 184 -834 184 -834 0 1
rlabel polysilicon 184 -840 184 -840 0 3
rlabel polysilicon 191 -834 191 -834 0 1
rlabel polysilicon 191 -840 191 -840 0 3
rlabel polysilicon 198 -834 198 -834 0 1
rlabel polysilicon 198 -840 198 -840 0 3
rlabel polysilicon 205 -834 205 -834 0 1
rlabel polysilicon 205 -840 205 -840 0 3
rlabel polysilicon 212 -834 212 -834 0 1
rlabel polysilicon 212 -840 212 -840 0 3
rlabel polysilicon 219 -834 219 -834 0 1
rlabel polysilicon 219 -840 219 -840 0 3
rlabel polysilicon 226 -834 226 -834 0 1
rlabel polysilicon 226 -840 226 -840 0 3
rlabel polysilicon 233 -834 233 -834 0 1
rlabel polysilicon 233 -840 233 -840 0 3
rlabel polysilicon 240 -834 240 -834 0 1
rlabel polysilicon 240 -840 240 -840 0 3
rlabel polysilicon 247 -834 247 -834 0 1
rlabel polysilicon 247 -840 247 -840 0 3
rlabel polysilicon 254 -834 254 -834 0 1
rlabel polysilicon 254 -840 254 -840 0 3
rlabel polysilicon 261 -834 261 -834 0 1
rlabel polysilicon 261 -840 261 -840 0 3
rlabel polysilicon 268 -834 268 -834 0 1
rlabel polysilicon 268 -840 268 -840 0 3
rlabel polysilicon 275 -834 275 -834 0 1
rlabel polysilicon 275 -840 275 -840 0 3
rlabel polysilicon 282 -834 282 -834 0 1
rlabel polysilicon 282 -840 282 -840 0 3
rlabel polysilicon 289 -834 289 -834 0 1
rlabel polysilicon 289 -840 289 -840 0 3
rlabel polysilicon 296 -834 296 -834 0 1
rlabel polysilicon 299 -834 299 -834 0 2
rlabel polysilicon 296 -840 296 -840 0 3
rlabel polysilicon 299 -840 299 -840 0 4
rlabel polysilicon 303 -834 303 -834 0 1
rlabel polysilicon 303 -840 303 -840 0 3
rlabel polysilicon 310 -834 310 -834 0 1
rlabel polysilicon 310 -840 310 -840 0 3
rlabel polysilicon 317 -834 317 -834 0 1
rlabel polysilicon 317 -840 317 -840 0 3
rlabel polysilicon 324 -834 324 -834 0 1
rlabel polysilicon 324 -840 324 -840 0 3
rlabel polysilicon 331 -834 331 -834 0 1
rlabel polysilicon 331 -840 331 -840 0 3
rlabel polysilicon 338 -834 338 -834 0 1
rlabel polysilicon 338 -840 338 -840 0 3
rlabel polysilicon 345 -834 345 -834 0 1
rlabel polysilicon 345 -840 345 -840 0 3
rlabel polysilicon 352 -834 352 -834 0 1
rlabel polysilicon 352 -840 352 -840 0 3
rlabel polysilicon 359 -834 359 -834 0 1
rlabel polysilicon 359 -840 359 -840 0 3
rlabel polysilicon 366 -834 366 -834 0 1
rlabel polysilicon 366 -840 366 -840 0 3
rlabel polysilicon 373 -834 373 -834 0 1
rlabel polysilicon 373 -840 373 -840 0 3
rlabel polysilicon 380 -834 380 -834 0 1
rlabel polysilicon 380 -840 380 -840 0 3
rlabel polysilicon 387 -834 387 -834 0 1
rlabel polysilicon 390 -834 390 -834 0 2
rlabel polysilicon 387 -840 387 -840 0 3
rlabel polysilicon 390 -840 390 -840 0 4
rlabel polysilicon 394 -834 394 -834 0 1
rlabel polysilicon 397 -834 397 -834 0 2
rlabel polysilicon 394 -840 394 -840 0 3
rlabel polysilicon 397 -840 397 -840 0 4
rlabel polysilicon 401 -834 401 -834 0 1
rlabel polysilicon 404 -834 404 -834 0 2
rlabel polysilicon 401 -840 401 -840 0 3
rlabel polysilicon 404 -840 404 -840 0 4
rlabel polysilicon 408 -834 408 -834 0 1
rlabel polysilicon 408 -840 408 -840 0 3
rlabel polysilicon 415 -834 415 -834 0 1
rlabel polysilicon 415 -840 415 -840 0 3
rlabel polysilicon 422 -834 422 -834 0 1
rlabel polysilicon 422 -840 422 -840 0 3
rlabel polysilicon 429 -834 429 -834 0 1
rlabel polysilicon 432 -834 432 -834 0 2
rlabel polysilicon 429 -840 429 -840 0 3
rlabel polysilicon 432 -840 432 -840 0 4
rlabel polysilicon 436 -840 436 -840 0 3
rlabel polysilicon 439 -840 439 -840 0 4
rlabel polysilicon 443 -834 443 -834 0 1
rlabel polysilicon 443 -840 443 -840 0 3
rlabel polysilicon 450 -834 450 -834 0 1
rlabel polysilicon 450 -840 450 -840 0 3
rlabel polysilicon 457 -834 457 -834 0 1
rlabel polysilicon 457 -840 457 -840 0 3
rlabel polysilicon 464 -834 464 -834 0 1
rlabel polysilicon 464 -840 464 -840 0 3
rlabel polysilicon 471 -834 471 -834 0 1
rlabel polysilicon 471 -840 471 -840 0 3
rlabel polysilicon 478 -834 478 -834 0 1
rlabel polysilicon 478 -840 478 -840 0 3
rlabel polysilicon 485 -834 485 -834 0 1
rlabel polysilicon 485 -840 485 -840 0 3
rlabel polysilicon 492 -834 492 -834 0 1
rlabel polysilicon 495 -834 495 -834 0 2
rlabel polysilicon 492 -840 492 -840 0 3
rlabel polysilicon 495 -840 495 -840 0 4
rlabel polysilicon 499 -834 499 -834 0 1
rlabel polysilicon 499 -840 499 -840 0 3
rlabel polysilicon 506 -834 506 -834 0 1
rlabel polysilicon 509 -834 509 -834 0 2
rlabel polysilicon 506 -840 506 -840 0 3
rlabel polysilicon 509 -840 509 -840 0 4
rlabel polysilicon 513 -834 513 -834 0 1
rlabel polysilicon 516 -834 516 -834 0 2
rlabel polysilicon 513 -840 513 -840 0 3
rlabel polysilicon 516 -840 516 -840 0 4
rlabel polysilicon 520 -834 520 -834 0 1
rlabel polysilicon 523 -834 523 -834 0 2
rlabel polysilicon 520 -840 520 -840 0 3
rlabel polysilicon 523 -840 523 -840 0 4
rlabel polysilicon 527 -834 527 -834 0 1
rlabel polysilicon 527 -840 527 -840 0 3
rlabel polysilicon 534 -834 534 -834 0 1
rlabel polysilicon 534 -840 534 -840 0 3
rlabel polysilicon 541 -834 541 -834 0 1
rlabel polysilicon 541 -840 541 -840 0 3
rlabel polysilicon 548 -834 548 -834 0 1
rlabel polysilicon 548 -840 548 -840 0 3
rlabel polysilicon 555 -834 555 -834 0 1
rlabel polysilicon 555 -840 555 -840 0 3
rlabel polysilicon 562 -834 562 -834 0 1
rlabel polysilicon 565 -834 565 -834 0 2
rlabel polysilicon 562 -840 562 -840 0 3
rlabel polysilicon 565 -840 565 -840 0 4
rlabel polysilicon 569 -834 569 -834 0 1
rlabel polysilicon 572 -834 572 -834 0 2
rlabel polysilicon 569 -840 569 -840 0 3
rlabel polysilicon 572 -840 572 -840 0 4
rlabel polysilicon 576 -834 576 -834 0 1
rlabel polysilicon 576 -840 576 -840 0 3
rlabel polysilicon 583 -834 583 -834 0 1
rlabel polysilicon 586 -834 586 -834 0 2
rlabel polysilicon 583 -840 583 -840 0 3
rlabel polysilicon 586 -840 586 -840 0 4
rlabel polysilicon 590 -834 590 -834 0 1
rlabel polysilicon 590 -840 590 -840 0 3
rlabel polysilicon 597 -834 597 -834 0 1
rlabel polysilicon 597 -840 597 -840 0 3
rlabel polysilicon 604 -834 604 -834 0 1
rlabel polysilicon 604 -840 604 -840 0 3
rlabel polysilicon 611 -834 611 -834 0 1
rlabel polysilicon 611 -840 611 -840 0 3
rlabel polysilicon 618 -834 618 -834 0 1
rlabel polysilicon 621 -834 621 -834 0 2
rlabel polysilicon 618 -840 618 -840 0 3
rlabel polysilicon 625 -834 625 -834 0 1
rlabel polysilicon 625 -840 625 -840 0 3
rlabel polysilicon 632 -834 632 -834 0 1
rlabel polysilicon 632 -840 632 -840 0 3
rlabel polysilicon 639 -834 639 -834 0 1
rlabel polysilicon 639 -840 639 -840 0 3
rlabel polysilicon 646 -834 646 -834 0 1
rlabel polysilicon 649 -834 649 -834 0 2
rlabel polysilicon 646 -840 646 -840 0 3
rlabel polysilicon 649 -840 649 -840 0 4
rlabel polysilicon 653 -834 653 -834 0 1
rlabel polysilicon 656 -834 656 -834 0 2
rlabel polysilicon 653 -840 653 -840 0 3
rlabel polysilicon 656 -840 656 -840 0 4
rlabel polysilicon 660 -834 660 -834 0 1
rlabel polysilicon 660 -840 660 -840 0 3
rlabel polysilicon 667 -834 667 -834 0 1
rlabel polysilicon 667 -840 667 -840 0 3
rlabel polysilicon 674 -834 674 -834 0 1
rlabel polysilicon 674 -840 674 -840 0 3
rlabel polysilicon 681 -834 681 -834 0 1
rlabel polysilicon 681 -840 681 -840 0 3
rlabel polysilicon 688 -834 688 -834 0 1
rlabel polysilicon 688 -840 688 -840 0 3
rlabel polysilicon 695 -834 695 -834 0 1
rlabel polysilicon 695 -840 695 -840 0 3
rlabel polysilicon 702 -834 702 -834 0 1
rlabel polysilicon 705 -834 705 -834 0 2
rlabel polysilicon 702 -840 702 -840 0 3
rlabel polysilicon 705 -840 705 -840 0 4
rlabel polysilicon 709 -834 709 -834 0 1
rlabel polysilicon 709 -840 709 -840 0 3
rlabel polysilicon 716 -834 716 -834 0 1
rlabel polysilicon 716 -840 716 -840 0 3
rlabel polysilicon 723 -834 723 -834 0 1
rlabel polysilicon 723 -840 723 -840 0 3
rlabel polysilicon 730 -834 730 -834 0 1
rlabel polysilicon 730 -840 730 -840 0 3
rlabel polysilicon 737 -834 737 -834 0 1
rlabel polysilicon 737 -840 737 -840 0 3
rlabel polysilicon 744 -834 744 -834 0 1
rlabel polysilicon 744 -840 744 -840 0 3
rlabel polysilicon 751 -834 751 -834 0 1
rlabel polysilicon 751 -840 751 -840 0 3
rlabel polysilicon 758 -834 758 -834 0 1
rlabel polysilicon 761 -834 761 -834 0 2
rlabel polysilicon 758 -840 758 -840 0 3
rlabel polysilicon 761 -840 761 -840 0 4
rlabel polysilicon 765 -834 765 -834 0 1
rlabel polysilicon 765 -840 765 -840 0 3
rlabel polysilicon 772 -834 772 -834 0 1
rlabel polysilicon 772 -840 772 -840 0 3
rlabel polysilicon 775 -840 775 -840 0 4
rlabel polysilicon 779 -834 779 -834 0 1
rlabel polysilicon 779 -840 779 -840 0 3
rlabel polysilicon 786 -834 786 -834 0 1
rlabel polysilicon 786 -840 786 -840 0 3
rlabel polysilicon 793 -834 793 -834 0 1
rlabel polysilicon 793 -840 793 -840 0 3
rlabel polysilicon 800 -834 800 -834 0 1
rlabel polysilicon 800 -840 800 -840 0 3
rlabel polysilicon 807 -834 807 -834 0 1
rlabel polysilicon 807 -840 807 -840 0 3
rlabel polysilicon 814 -834 814 -834 0 1
rlabel polysilicon 814 -840 814 -840 0 3
rlabel polysilicon 821 -834 821 -834 0 1
rlabel polysilicon 821 -840 821 -840 0 3
rlabel polysilicon 828 -834 828 -834 0 1
rlabel polysilicon 828 -840 828 -840 0 3
rlabel polysilicon 831 -840 831 -840 0 4
rlabel polysilicon 835 -834 835 -834 0 1
rlabel polysilicon 835 -840 835 -840 0 3
rlabel polysilicon 842 -834 842 -834 0 1
rlabel polysilicon 842 -840 842 -840 0 3
rlabel polysilicon 849 -834 849 -834 0 1
rlabel polysilicon 849 -840 849 -840 0 3
rlabel polysilicon 856 -834 856 -834 0 1
rlabel polysilicon 856 -840 856 -840 0 3
rlabel polysilicon 863 -834 863 -834 0 1
rlabel polysilicon 863 -840 863 -840 0 3
rlabel polysilicon 870 -834 870 -834 0 1
rlabel polysilicon 870 -840 870 -840 0 3
rlabel polysilicon 877 -834 877 -834 0 1
rlabel polysilicon 877 -840 877 -840 0 3
rlabel polysilicon 884 -834 884 -834 0 1
rlabel polysilicon 884 -840 884 -840 0 3
rlabel polysilicon 891 -834 891 -834 0 1
rlabel polysilicon 891 -840 891 -840 0 3
rlabel polysilicon 898 -834 898 -834 0 1
rlabel polysilicon 898 -840 898 -840 0 3
rlabel polysilicon 905 -834 905 -834 0 1
rlabel polysilicon 905 -840 905 -840 0 3
rlabel polysilicon 912 -834 912 -834 0 1
rlabel polysilicon 912 -840 912 -840 0 3
rlabel polysilicon 919 -834 919 -834 0 1
rlabel polysilicon 919 -840 919 -840 0 3
rlabel polysilicon 926 -834 926 -834 0 1
rlabel polysilicon 926 -840 926 -840 0 3
rlabel polysilicon 933 -834 933 -834 0 1
rlabel polysilicon 933 -840 933 -840 0 3
rlabel polysilicon 940 -834 940 -834 0 1
rlabel polysilicon 940 -840 940 -840 0 3
rlabel polysilicon 947 -834 947 -834 0 1
rlabel polysilicon 947 -840 947 -840 0 3
rlabel polysilicon 954 -834 954 -834 0 1
rlabel polysilicon 954 -840 954 -840 0 3
rlabel polysilicon 961 -834 961 -834 0 1
rlabel polysilicon 961 -840 961 -840 0 3
rlabel polysilicon 968 -834 968 -834 0 1
rlabel polysilicon 968 -840 968 -840 0 3
rlabel polysilicon 975 -834 975 -834 0 1
rlabel polysilicon 975 -840 975 -840 0 3
rlabel polysilicon 982 -834 982 -834 0 1
rlabel polysilicon 982 -840 982 -840 0 3
rlabel polysilicon 989 -834 989 -834 0 1
rlabel polysilicon 989 -840 989 -840 0 3
rlabel polysilicon 996 -834 996 -834 0 1
rlabel polysilicon 996 -840 996 -840 0 3
rlabel polysilicon 1003 -834 1003 -834 0 1
rlabel polysilicon 1003 -840 1003 -840 0 3
rlabel polysilicon 1010 -834 1010 -834 0 1
rlabel polysilicon 1010 -840 1010 -840 0 3
rlabel polysilicon 1017 -834 1017 -834 0 1
rlabel polysilicon 1017 -840 1017 -840 0 3
rlabel polysilicon 1024 -834 1024 -834 0 1
rlabel polysilicon 1024 -840 1024 -840 0 3
rlabel polysilicon 1031 -834 1031 -834 0 1
rlabel polysilicon 1031 -840 1031 -840 0 3
rlabel polysilicon 1038 -834 1038 -834 0 1
rlabel polysilicon 1038 -840 1038 -840 0 3
rlabel polysilicon 1045 -834 1045 -834 0 1
rlabel polysilicon 1045 -840 1045 -840 0 3
rlabel polysilicon 1052 -834 1052 -834 0 1
rlabel polysilicon 1052 -840 1052 -840 0 3
rlabel polysilicon 1059 -834 1059 -834 0 1
rlabel polysilicon 1059 -840 1059 -840 0 3
rlabel polysilicon 1066 -834 1066 -834 0 1
rlabel polysilicon 1066 -840 1066 -840 0 3
rlabel polysilicon 1073 -834 1073 -834 0 1
rlabel polysilicon 1073 -840 1073 -840 0 3
rlabel polysilicon 1080 -834 1080 -834 0 1
rlabel polysilicon 1080 -840 1080 -840 0 3
rlabel polysilicon 1087 -834 1087 -834 0 1
rlabel polysilicon 1087 -840 1087 -840 0 3
rlabel polysilicon 1094 -834 1094 -834 0 1
rlabel polysilicon 1094 -840 1094 -840 0 3
rlabel polysilicon 1101 -834 1101 -834 0 1
rlabel polysilicon 1101 -840 1101 -840 0 3
rlabel polysilicon 1108 -834 1108 -834 0 1
rlabel polysilicon 1108 -840 1108 -840 0 3
rlabel polysilicon 1115 -834 1115 -834 0 1
rlabel polysilicon 1115 -840 1115 -840 0 3
rlabel polysilicon 1122 -834 1122 -834 0 1
rlabel polysilicon 1122 -840 1122 -840 0 3
rlabel polysilicon 1129 -834 1129 -834 0 1
rlabel polysilicon 1129 -840 1129 -840 0 3
rlabel polysilicon 1136 -834 1136 -834 0 1
rlabel polysilicon 1136 -840 1136 -840 0 3
rlabel polysilicon 1143 -834 1143 -834 0 1
rlabel polysilicon 1143 -840 1143 -840 0 3
rlabel polysilicon 1150 -834 1150 -834 0 1
rlabel polysilicon 1150 -840 1150 -840 0 3
rlabel polysilicon 1157 -834 1157 -834 0 1
rlabel polysilicon 1157 -840 1157 -840 0 3
rlabel polysilicon 1164 -834 1164 -834 0 1
rlabel polysilicon 1164 -840 1164 -840 0 3
rlabel polysilicon 1171 -834 1171 -834 0 1
rlabel polysilicon 1171 -840 1171 -840 0 3
rlabel polysilicon 1178 -834 1178 -834 0 1
rlabel polysilicon 1178 -840 1178 -840 0 3
rlabel polysilicon 1185 -834 1185 -834 0 1
rlabel polysilicon 1185 -840 1185 -840 0 3
rlabel polysilicon 1192 -834 1192 -834 0 1
rlabel polysilicon 1192 -840 1192 -840 0 3
rlabel polysilicon 1199 -834 1199 -834 0 1
rlabel polysilicon 1199 -840 1199 -840 0 3
rlabel polysilicon 1206 -834 1206 -834 0 1
rlabel polysilicon 1206 -840 1206 -840 0 3
rlabel polysilicon 1213 -834 1213 -834 0 1
rlabel polysilicon 1213 -840 1213 -840 0 3
rlabel polysilicon 1220 -834 1220 -834 0 1
rlabel polysilicon 1220 -840 1220 -840 0 3
rlabel polysilicon 1227 -834 1227 -834 0 1
rlabel polysilicon 1227 -840 1227 -840 0 3
rlabel polysilicon 1234 -834 1234 -834 0 1
rlabel polysilicon 1234 -840 1234 -840 0 3
rlabel polysilicon 1241 -834 1241 -834 0 1
rlabel polysilicon 1241 -840 1241 -840 0 3
rlabel polysilicon 1248 -834 1248 -834 0 1
rlabel polysilicon 1248 -840 1248 -840 0 3
rlabel polysilicon 1255 -834 1255 -834 0 1
rlabel polysilicon 1255 -840 1255 -840 0 3
rlabel polysilicon 1262 -834 1262 -834 0 1
rlabel polysilicon 1262 -840 1262 -840 0 3
rlabel polysilicon 1416 -834 1416 -834 0 1
rlabel polysilicon 1416 -840 1416 -840 0 3
rlabel polysilicon 2 -951 2 -951 0 1
rlabel polysilicon 2 -957 2 -957 0 3
rlabel polysilicon 9 -951 9 -951 0 1
rlabel polysilicon 9 -957 9 -957 0 3
rlabel polysilicon 16 -951 16 -951 0 1
rlabel polysilicon 16 -957 16 -957 0 3
rlabel polysilicon 23 -951 23 -951 0 1
rlabel polysilicon 23 -957 23 -957 0 3
rlabel polysilicon 30 -951 30 -951 0 1
rlabel polysilicon 30 -957 30 -957 0 3
rlabel polysilicon 37 -951 37 -951 0 1
rlabel polysilicon 37 -957 37 -957 0 3
rlabel polysilicon 44 -951 44 -951 0 1
rlabel polysilicon 44 -957 44 -957 0 3
rlabel polysilicon 51 -951 51 -951 0 1
rlabel polysilicon 51 -957 51 -957 0 3
rlabel polysilicon 58 -951 58 -951 0 1
rlabel polysilicon 58 -957 58 -957 0 3
rlabel polysilicon 65 -951 65 -951 0 1
rlabel polysilicon 68 -951 68 -951 0 2
rlabel polysilicon 65 -957 65 -957 0 3
rlabel polysilicon 68 -957 68 -957 0 4
rlabel polysilicon 72 -951 72 -951 0 1
rlabel polysilicon 72 -957 72 -957 0 3
rlabel polysilicon 79 -951 79 -951 0 1
rlabel polysilicon 79 -957 79 -957 0 3
rlabel polysilicon 86 -951 86 -951 0 1
rlabel polysilicon 89 -951 89 -951 0 2
rlabel polysilicon 86 -957 86 -957 0 3
rlabel polysilicon 89 -957 89 -957 0 4
rlabel polysilicon 93 -951 93 -951 0 1
rlabel polysilicon 93 -957 93 -957 0 3
rlabel polysilicon 100 -951 100 -951 0 1
rlabel polysilicon 100 -957 100 -957 0 3
rlabel polysilicon 107 -951 107 -951 0 1
rlabel polysilicon 107 -957 107 -957 0 3
rlabel polysilicon 114 -951 114 -951 0 1
rlabel polysilicon 114 -957 114 -957 0 3
rlabel polysilicon 121 -951 121 -951 0 1
rlabel polysilicon 124 -951 124 -951 0 2
rlabel polysilicon 121 -957 121 -957 0 3
rlabel polysilicon 124 -957 124 -957 0 4
rlabel polysilicon 128 -951 128 -951 0 1
rlabel polysilicon 131 -951 131 -951 0 2
rlabel polysilicon 128 -957 128 -957 0 3
rlabel polysilicon 131 -957 131 -957 0 4
rlabel polysilicon 135 -951 135 -951 0 1
rlabel polysilicon 135 -957 135 -957 0 3
rlabel polysilicon 142 -951 142 -951 0 1
rlabel polysilicon 142 -957 142 -957 0 3
rlabel polysilicon 152 -951 152 -951 0 2
rlabel polysilicon 149 -957 149 -957 0 3
rlabel polysilicon 152 -957 152 -957 0 4
rlabel polysilicon 156 -951 156 -951 0 1
rlabel polysilicon 156 -957 156 -957 0 3
rlabel polysilicon 163 -951 163 -951 0 1
rlabel polysilicon 163 -957 163 -957 0 3
rlabel polysilicon 170 -951 170 -951 0 1
rlabel polysilicon 170 -957 170 -957 0 3
rlabel polysilicon 177 -951 177 -951 0 1
rlabel polysilicon 177 -957 177 -957 0 3
rlabel polysilicon 184 -951 184 -951 0 1
rlabel polysilicon 184 -957 184 -957 0 3
rlabel polysilicon 191 -951 191 -951 0 1
rlabel polysilicon 191 -957 191 -957 0 3
rlabel polysilicon 198 -951 198 -951 0 1
rlabel polysilicon 201 -951 201 -951 0 2
rlabel polysilicon 198 -957 198 -957 0 3
rlabel polysilicon 201 -957 201 -957 0 4
rlabel polysilicon 205 -951 205 -951 0 1
rlabel polysilicon 205 -957 205 -957 0 3
rlabel polysilicon 212 -951 212 -951 0 1
rlabel polysilicon 215 -951 215 -951 0 2
rlabel polysilicon 212 -957 212 -957 0 3
rlabel polysilicon 219 -951 219 -951 0 1
rlabel polysilicon 219 -957 219 -957 0 3
rlabel polysilicon 226 -951 226 -951 0 1
rlabel polysilicon 226 -957 226 -957 0 3
rlabel polysilicon 233 -951 233 -951 0 1
rlabel polysilicon 233 -957 233 -957 0 3
rlabel polysilicon 240 -951 240 -951 0 1
rlabel polysilicon 240 -957 240 -957 0 3
rlabel polysilicon 247 -951 247 -951 0 1
rlabel polysilicon 247 -957 247 -957 0 3
rlabel polysilicon 254 -951 254 -951 0 1
rlabel polysilicon 254 -957 254 -957 0 3
rlabel polysilicon 261 -951 261 -951 0 1
rlabel polysilicon 261 -957 261 -957 0 3
rlabel polysilicon 268 -951 268 -951 0 1
rlabel polysilicon 268 -957 268 -957 0 3
rlabel polysilicon 275 -951 275 -951 0 1
rlabel polysilicon 275 -957 275 -957 0 3
rlabel polysilicon 282 -951 282 -951 0 1
rlabel polysilicon 282 -957 282 -957 0 3
rlabel polysilicon 289 -951 289 -951 0 1
rlabel polysilicon 289 -957 289 -957 0 3
rlabel polysilicon 296 -951 296 -951 0 1
rlabel polysilicon 296 -957 296 -957 0 3
rlabel polysilicon 303 -951 303 -951 0 1
rlabel polysilicon 303 -957 303 -957 0 3
rlabel polysilicon 310 -951 310 -951 0 1
rlabel polysilicon 310 -957 310 -957 0 3
rlabel polysilicon 317 -951 317 -951 0 1
rlabel polysilicon 320 -951 320 -951 0 2
rlabel polysilicon 317 -957 317 -957 0 3
rlabel polysilicon 320 -957 320 -957 0 4
rlabel polysilicon 324 -951 324 -951 0 1
rlabel polysilicon 324 -957 324 -957 0 3
rlabel polysilicon 331 -951 331 -951 0 1
rlabel polysilicon 331 -957 331 -957 0 3
rlabel polysilicon 338 -951 338 -951 0 1
rlabel polysilicon 338 -957 338 -957 0 3
rlabel polysilicon 345 -951 345 -951 0 1
rlabel polysilicon 345 -957 345 -957 0 3
rlabel polysilicon 352 -951 352 -951 0 1
rlabel polysilicon 352 -957 352 -957 0 3
rlabel polysilicon 359 -951 359 -951 0 1
rlabel polysilicon 359 -957 359 -957 0 3
rlabel polysilicon 366 -951 366 -951 0 1
rlabel polysilicon 369 -951 369 -951 0 2
rlabel polysilicon 366 -957 366 -957 0 3
rlabel polysilicon 369 -957 369 -957 0 4
rlabel polysilicon 373 -951 373 -951 0 1
rlabel polysilicon 373 -957 373 -957 0 3
rlabel polysilicon 380 -951 380 -951 0 1
rlabel polysilicon 380 -957 380 -957 0 3
rlabel polysilicon 387 -951 387 -951 0 1
rlabel polysilicon 387 -957 387 -957 0 3
rlabel polysilicon 394 -951 394 -951 0 1
rlabel polysilicon 394 -957 394 -957 0 3
rlabel polysilicon 401 -951 401 -951 0 1
rlabel polysilicon 401 -957 401 -957 0 3
rlabel polysilicon 408 -951 408 -951 0 1
rlabel polysilicon 408 -957 408 -957 0 3
rlabel polysilicon 415 -951 415 -951 0 1
rlabel polysilicon 415 -957 415 -957 0 3
rlabel polysilicon 422 -951 422 -951 0 1
rlabel polysilicon 425 -951 425 -951 0 2
rlabel polysilicon 422 -957 422 -957 0 3
rlabel polysilicon 425 -957 425 -957 0 4
rlabel polysilicon 429 -951 429 -951 0 1
rlabel polysilicon 429 -957 429 -957 0 3
rlabel polysilicon 436 -951 436 -951 0 1
rlabel polysilicon 436 -957 436 -957 0 3
rlabel polysilicon 443 -951 443 -951 0 1
rlabel polysilicon 443 -957 443 -957 0 3
rlabel polysilicon 450 -951 450 -951 0 1
rlabel polysilicon 450 -957 450 -957 0 3
rlabel polysilicon 453 -957 453 -957 0 4
rlabel polysilicon 457 -951 457 -951 0 1
rlabel polysilicon 457 -957 457 -957 0 3
rlabel polysilicon 464 -951 464 -951 0 1
rlabel polysilicon 464 -957 464 -957 0 3
rlabel polysilicon 471 -951 471 -951 0 1
rlabel polysilicon 471 -957 471 -957 0 3
rlabel polysilicon 478 -951 478 -951 0 1
rlabel polysilicon 481 -951 481 -951 0 2
rlabel polysilicon 478 -957 478 -957 0 3
rlabel polysilicon 481 -957 481 -957 0 4
rlabel polysilicon 485 -951 485 -951 0 1
rlabel polysilicon 485 -957 485 -957 0 3
rlabel polysilicon 492 -951 492 -951 0 1
rlabel polysilicon 492 -957 492 -957 0 3
rlabel polysilicon 499 -951 499 -951 0 1
rlabel polysilicon 502 -951 502 -951 0 2
rlabel polysilicon 499 -957 499 -957 0 3
rlabel polysilicon 502 -957 502 -957 0 4
rlabel polysilicon 506 -951 506 -951 0 1
rlabel polysilicon 506 -957 506 -957 0 3
rlabel polysilicon 513 -951 513 -951 0 1
rlabel polysilicon 513 -957 513 -957 0 3
rlabel polysilicon 520 -951 520 -951 0 1
rlabel polysilicon 520 -957 520 -957 0 3
rlabel polysilicon 527 -957 527 -957 0 3
rlabel polysilicon 530 -957 530 -957 0 4
rlabel polysilicon 534 -951 534 -951 0 1
rlabel polysilicon 537 -951 537 -951 0 2
rlabel polysilicon 534 -957 534 -957 0 3
rlabel polysilicon 537 -957 537 -957 0 4
rlabel polysilicon 541 -951 541 -951 0 1
rlabel polysilicon 544 -951 544 -951 0 2
rlabel polysilicon 541 -957 541 -957 0 3
rlabel polysilicon 544 -957 544 -957 0 4
rlabel polysilicon 548 -951 548 -951 0 1
rlabel polysilicon 548 -957 548 -957 0 3
rlabel polysilicon 555 -951 555 -951 0 1
rlabel polysilicon 555 -957 555 -957 0 3
rlabel polysilicon 562 -951 562 -951 0 1
rlabel polysilicon 562 -957 562 -957 0 3
rlabel polysilicon 569 -951 569 -951 0 1
rlabel polysilicon 569 -957 569 -957 0 3
rlabel polysilicon 576 -951 576 -951 0 1
rlabel polysilicon 576 -957 576 -957 0 3
rlabel polysilicon 583 -951 583 -951 0 1
rlabel polysilicon 583 -957 583 -957 0 3
rlabel polysilicon 590 -951 590 -951 0 1
rlabel polysilicon 590 -957 590 -957 0 3
rlabel polysilicon 597 -951 597 -951 0 1
rlabel polysilicon 597 -957 597 -957 0 3
rlabel polysilicon 604 -951 604 -951 0 1
rlabel polysilicon 604 -957 604 -957 0 3
rlabel polysilicon 611 -951 611 -951 0 1
rlabel polysilicon 614 -951 614 -951 0 2
rlabel polysilicon 611 -957 611 -957 0 3
rlabel polysilicon 614 -957 614 -957 0 4
rlabel polysilicon 618 -951 618 -951 0 1
rlabel polysilicon 618 -957 618 -957 0 3
rlabel polysilicon 625 -951 625 -951 0 1
rlabel polysilicon 628 -951 628 -951 0 2
rlabel polysilicon 625 -957 625 -957 0 3
rlabel polysilicon 632 -951 632 -951 0 1
rlabel polysilicon 635 -951 635 -951 0 2
rlabel polysilicon 632 -957 632 -957 0 3
rlabel polysilicon 635 -957 635 -957 0 4
rlabel polysilicon 639 -951 639 -951 0 1
rlabel polysilicon 639 -957 639 -957 0 3
rlabel polysilicon 646 -951 646 -951 0 1
rlabel polysilicon 646 -957 646 -957 0 3
rlabel polysilicon 653 -951 653 -951 0 1
rlabel polysilicon 656 -951 656 -951 0 2
rlabel polysilicon 653 -957 653 -957 0 3
rlabel polysilicon 656 -957 656 -957 0 4
rlabel polysilicon 660 -951 660 -951 0 1
rlabel polysilicon 660 -957 660 -957 0 3
rlabel polysilicon 667 -951 667 -951 0 1
rlabel polysilicon 667 -957 667 -957 0 3
rlabel polysilicon 674 -951 674 -951 0 1
rlabel polysilicon 674 -957 674 -957 0 3
rlabel polysilicon 681 -951 681 -951 0 1
rlabel polysilicon 681 -957 681 -957 0 3
rlabel polysilicon 688 -951 688 -951 0 1
rlabel polysilicon 691 -951 691 -951 0 2
rlabel polysilicon 688 -957 688 -957 0 3
rlabel polysilicon 695 -951 695 -951 0 1
rlabel polysilicon 695 -957 695 -957 0 3
rlabel polysilicon 702 -951 702 -951 0 1
rlabel polysilicon 702 -957 702 -957 0 3
rlabel polysilicon 709 -951 709 -951 0 1
rlabel polysilicon 712 -951 712 -951 0 2
rlabel polysilicon 709 -957 709 -957 0 3
rlabel polysilicon 712 -957 712 -957 0 4
rlabel polysilicon 716 -951 716 -951 0 1
rlabel polysilicon 719 -951 719 -951 0 2
rlabel polysilicon 719 -957 719 -957 0 4
rlabel polysilicon 723 -951 723 -951 0 1
rlabel polysilicon 723 -957 723 -957 0 3
rlabel polysilicon 730 -951 730 -951 0 1
rlabel polysilicon 730 -957 730 -957 0 3
rlabel polysilicon 737 -951 737 -951 0 1
rlabel polysilicon 737 -957 737 -957 0 3
rlabel polysilicon 747 -951 747 -951 0 2
rlabel polysilicon 744 -957 744 -957 0 3
rlabel polysilicon 747 -957 747 -957 0 4
rlabel polysilicon 751 -951 751 -951 0 1
rlabel polysilicon 751 -957 751 -957 0 3
rlabel polysilicon 758 -951 758 -951 0 1
rlabel polysilicon 758 -957 758 -957 0 3
rlabel polysilicon 765 -951 765 -951 0 1
rlabel polysilicon 765 -957 765 -957 0 3
rlabel polysilicon 772 -951 772 -951 0 1
rlabel polysilicon 772 -957 772 -957 0 3
rlabel polysilicon 779 -951 779 -951 0 1
rlabel polysilicon 779 -957 779 -957 0 3
rlabel polysilicon 786 -951 786 -951 0 1
rlabel polysilicon 786 -957 786 -957 0 3
rlabel polysilicon 793 -951 793 -951 0 1
rlabel polysilicon 793 -957 793 -957 0 3
rlabel polysilicon 800 -951 800 -951 0 1
rlabel polysilicon 800 -957 800 -957 0 3
rlabel polysilicon 807 -951 807 -951 0 1
rlabel polysilicon 807 -957 807 -957 0 3
rlabel polysilicon 814 -951 814 -951 0 1
rlabel polysilicon 814 -957 814 -957 0 3
rlabel polysilicon 821 -951 821 -951 0 1
rlabel polysilicon 824 -951 824 -951 0 2
rlabel polysilicon 821 -957 821 -957 0 3
rlabel polysilicon 824 -957 824 -957 0 4
rlabel polysilicon 828 -951 828 -951 0 1
rlabel polysilicon 828 -957 828 -957 0 3
rlabel polysilicon 835 -951 835 -951 0 1
rlabel polysilicon 835 -957 835 -957 0 3
rlabel polysilicon 842 -951 842 -951 0 1
rlabel polysilicon 842 -957 842 -957 0 3
rlabel polysilicon 849 -951 849 -951 0 1
rlabel polysilicon 849 -957 849 -957 0 3
rlabel polysilicon 856 -951 856 -951 0 1
rlabel polysilicon 856 -957 856 -957 0 3
rlabel polysilicon 863 -951 863 -951 0 1
rlabel polysilicon 863 -957 863 -957 0 3
rlabel polysilicon 870 -951 870 -951 0 1
rlabel polysilicon 870 -957 870 -957 0 3
rlabel polysilicon 877 -951 877 -951 0 1
rlabel polysilicon 877 -957 877 -957 0 3
rlabel polysilicon 884 -951 884 -951 0 1
rlabel polysilicon 884 -957 884 -957 0 3
rlabel polysilicon 891 -951 891 -951 0 1
rlabel polysilicon 891 -957 891 -957 0 3
rlabel polysilicon 898 -951 898 -951 0 1
rlabel polysilicon 898 -957 898 -957 0 3
rlabel polysilicon 905 -951 905 -951 0 1
rlabel polysilicon 905 -957 905 -957 0 3
rlabel polysilicon 912 -951 912 -951 0 1
rlabel polysilicon 912 -957 912 -957 0 3
rlabel polysilicon 919 -951 919 -951 0 1
rlabel polysilicon 919 -957 919 -957 0 3
rlabel polysilicon 926 -951 926 -951 0 1
rlabel polysilicon 926 -957 926 -957 0 3
rlabel polysilicon 933 -951 933 -951 0 1
rlabel polysilicon 933 -957 933 -957 0 3
rlabel polysilicon 940 -951 940 -951 0 1
rlabel polysilicon 940 -957 940 -957 0 3
rlabel polysilicon 947 -951 947 -951 0 1
rlabel polysilicon 947 -957 947 -957 0 3
rlabel polysilicon 954 -951 954 -951 0 1
rlabel polysilicon 954 -957 954 -957 0 3
rlabel polysilicon 961 -951 961 -951 0 1
rlabel polysilicon 961 -957 961 -957 0 3
rlabel polysilicon 968 -951 968 -951 0 1
rlabel polysilicon 968 -957 968 -957 0 3
rlabel polysilicon 975 -951 975 -951 0 1
rlabel polysilicon 975 -957 975 -957 0 3
rlabel polysilicon 982 -951 982 -951 0 1
rlabel polysilicon 982 -957 982 -957 0 3
rlabel polysilicon 989 -951 989 -951 0 1
rlabel polysilicon 989 -957 989 -957 0 3
rlabel polysilicon 996 -951 996 -951 0 1
rlabel polysilicon 996 -957 996 -957 0 3
rlabel polysilicon 1003 -951 1003 -951 0 1
rlabel polysilicon 1003 -957 1003 -957 0 3
rlabel polysilicon 1010 -951 1010 -951 0 1
rlabel polysilicon 1010 -957 1010 -957 0 3
rlabel polysilicon 1017 -951 1017 -951 0 1
rlabel polysilicon 1017 -957 1017 -957 0 3
rlabel polysilicon 1024 -951 1024 -951 0 1
rlabel polysilicon 1024 -957 1024 -957 0 3
rlabel polysilicon 1031 -951 1031 -951 0 1
rlabel polysilicon 1031 -957 1031 -957 0 3
rlabel polysilicon 1038 -951 1038 -951 0 1
rlabel polysilicon 1038 -957 1038 -957 0 3
rlabel polysilicon 1045 -951 1045 -951 0 1
rlabel polysilicon 1045 -957 1045 -957 0 3
rlabel polysilicon 1052 -951 1052 -951 0 1
rlabel polysilicon 1052 -957 1052 -957 0 3
rlabel polysilicon 1059 -951 1059 -951 0 1
rlabel polysilicon 1059 -957 1059 -957 0 3
rlabel polysilicon 1066 -951 1066 -951 0 1
rlabel polysilicon 1066 -957 1066 -957 0 3
rlabel polysilicon 1073 -951 1073 -951 0 1
rlabel polysilicon 1073 -957 1073 -957 0 3
rlabel polysilicon 1080 -951 1080 -951 0 1
rlabel polysilicon 1080 -957 1080 -957 0 3
rlabel polysilicon 1087 -951 1087 -951 0 1
rlabel polysilicon 1087 -957 1087 -957 0 3
rlabel polysilicon 1094 -951 1094 -951 0 1
rlabel polysilicon 1094 -957 1094 -957 0 3
rlabel polysilicon 1101 -951 1101 -951 0 1
rlabel polysilicon 1101 -957 1101 -957 0 3
rlabel polysilicon 1108 -951 1108 -951 0 1
rlabel polysilicon 1108 -957 1108 -957 0 3
rlabel polysilicon 1115 -951 1115 -951 0 1
rlabel polysilicon 1115 -957 1115 -957 0 3
rlabel polysilicon 1122 -951 1122 -951 0 1
rlabel polysilicon 1122 -957 1122 -957 0 3
rlabel polysilicon 1129 -951 1129 -951 0 1
rlabel polysilicon 1129 -957 1129 -957 0 3
rlabel polysilicon 1136 -951 1136 -951 0 1
rlabel polysilicon 1136 -957 1136 -957 0 3
rlabel polysilicon 1143 -951 1143 -951 0 1
rlabel polysilicon 1143 -957 1143 -957 0 3
rlabel polysilicon 1150 -951 1150 -951 0 1
rlabel polysilicon 1150 -957 1150 -957 0 3
rlabel polysilicon 1157 -951 1157 -951 0 1
rlabel polysilicon 1157 -957 1157 -957 0 3
rlabel polysilicon 1164 -951 1164 -951 0 1
rlabel polysilicon 1164 -957 1164 -957 0 3
rlabel polysilicon 1171 -951 1171 -951 0 1
rlabel polysilicon 1171 -957 1171 -957 0 3
rlabel polysilicon 1178 -951 1178 -951 0 1
rlabel polysilicon 1178 -957 1178 -957 0 3
rlabel polysilicon 1185 -951 1185 -951 0 1
rlabel polysilicon 1185 -957 1185 -957 0 3
rlabel polysilicon 1192 -951 1192 -951 0 1
rlabel polysilicon 1192 -957 1192 -957 0 3
rlabel polysilicon 1195 -957 1195 -957 0 4
rlabel polysilicon 1199 -951 1199 -951 0 1
rlabel polysilicon 1202 -951 1202 -951 0 2
rlabel polysilicon 1199 -957 1199 -957 0 3
rlabel polysilicon 1206 -951 1206 -951 0 1
rlabel polysilicon 1206 -957 1206 -957 0 3
rlabel polysilicon 1437 -951 1437 -951 0 1
rlabel polysilicon 1437 -957 1437 -957 0 3
rlabel polysilicon 2 -1080 2 -1080 0 1
rlabel polysilicon 5 -1080 5 -1080 0 2
rlabel polysilicon 5 -1086 5 -1086 0 4
rlabel polysilicon 9 -1080 9 -1080 0 1
rlabel polysilicon 9 -1086 9 -1086 0 3
rlabel polysilicon 16 -1080 16 -1080 0 1
rlabel polysilicon 16 -1086 16 -1086 0 3
rlabel polysilicon 23 -1080 23 -1080 0 1
rlabel polysilicon 23 -1086 23 -1086 0 3
rlabel polysilicon 30 -1080 30 -1080 0 1
rlabel polysilicon 33 -1080 33 -1080 0 2
rlabel polysilicon 33 -1086 33 -1086 0 4
rlabel polysilicon 37 -1080 37 -1080 0 1
rlabel polysilicon 40 -1080 40 -1080 0 2
rlabel polysilicon 40 -1086 40 -1086 0 4
rlabel polysilicon 44 -1080 44 -1080 0 1
rlabel polysilicon 44 -1086 44 -1086 0 3
rlabel polysilicon 51 -1080 51 -1080 0 1
rlabel polysilicon 54 -1080 54 -1080 0 2
rlabel polysilicon 51 -1086 51 -1086 0 3
rlabel polysilicon 54 -1086 54 -1086 0 4
rlabel polysilicon 58 -1080 58 -1080 0 1
rlabel polysilicon 58 -1086 58 -1086 0 3
rlabel polysilicon 65 -1080 65 -1080 0 1
rlabel polysilicon 65 -1086 65 -1086 0 3
rlabel polysilicon 72 -1080 72 -1080 0 1
rlabel polysilicon 75 -1080 75 -1080 0 2
rlabel polysilicon 72 -1086 72 -1086 0 3
rlabel polysilicon 75 -1086 75 -1086 0 4
rlabel polysilicon 79 -1080 79 -1080 0 1
rlabel polysilicon 79 -1086 79 -1086 0 3
rlabel polysilicon 86 -1080 86 -1080 0 1
rlabel polysilicon 86 -1086 86 -1086 0 3
rlabel polysilicon 93 -1080 93 -1080 0 1
rlabel polysilicon 96 -1080 96 -1080 0 2
rlabel polysilicon 93 -1086 93 -1086 0 3
rlabel polysilicon 96 -1086 96 -1086 0 4
rlabel polysilicon 100 -1080 100 -1080 0 1
rlabel polysilicon 103 -1080 103 -1080 0 2
rlabel polysilicon 100 -1086 100 -1086 0 3
rlabel polysilicon 103 -1086 103 -1086 0 4
rlabel polysilicon 107 -1080 107 -1080 0 1
rlabel polysilicon 107 -1086 107 -1086 0 3
rlabel polysilicon 114 -1080 114 -1080 0 1
rlabel polysilicon 114 -1086 114 -1086 0 3
rlabel polysilicon 121 -1080 121 -1080 0 1
rlabel polysilicon 121 -1086 121 -1086 0 3
rlabel polysilicon 128 -1080 128 -1080 0 1
rlabel polysilicon 128 -1086 128 -1086 0 3
rlabel polysilicon 135 -1080 135 -1080 0 1
rlabel polysilicon 135 -1086 135 -1086 0 3
rlabel polysilicon 142 -1080 142 -1080 0 1
rlabel polysilicon 142 -1086 142 -1086 0 3
rlabel polysilicon 149 -1080 149 -1080 0 1
rlabel polysilicon 149 -1086 149 -1086 0 3
rlabel polysilicon 152 -1086 152 -1086 0 4
rlabel polysilicon 156 -1080 156 -1080 0 1
rlabel polysilicon 156 -1086 156 -1086 0 3
rlabel polysilicon 163 -1080 163 -1080 0 1
rlabel polysilicon 163 -1086 163 -1086 0 3
rlabel polysilicon 170 -1080 170 -1080 0 1
rlabel polysilicon 170 -1086 170 -1086 0 3
rlabel polysilicon 177 -1080 177 -1080 0 1
rlabel polysilicon 177 -1086 177 -1086 0 3
rlabel polysilicon 184 -1080 184 -1080 0 1
rlabel polysilicon 184 -1086 184 -1086 0 3
rlabel polysilicon 191 -1080 191 -1080 0 1
rlabel polysilicon 191 -1086 191 -1086 0 3
rlabel polysilicon 198 -1080 198 -1080 0 1
rlabel polysilicon 198 -1086 198 -1086 0 3
rlabel polysilicon 205 -1080 205 -1080 0 1
rlabel polysilicon 205 -1086 205 -1086 0 3
rlabel polysilicon 212 -1080 212 -1080 0 1
rlabel polysilicon 212 -1086 212 -1086 0 3
rlabel polysilicon 219 -1080 219 -1080 0 1
rlabel polysilicon 219 -1086 219 -1086 0 3
rlabel polysilicon 226 -1080 226 -1080 0 1
rlabel polysilicon 226 -1086 226 -1086 0 3
rlabel polysilicon 233 -1080 233 -1080 0 1
rlabel polysilicon 233 -1086 233 -1086 0 3
rlabel polysilicon 240 -1080 240 -1080 0 1
rlabel polysilicon 240 -1086 240 -1086 0 3
rlabel polysilicon 247 -1080 247 -1080 0 1
rlabel polysilicon 247 -1086 247 -1086 0 3
rlabel polysilicon 254 -1080 254 -1080 0 1
rlabel polysilicon 254 -1086 254 -1086 0 3
rlabel polysilicon 261 -1080 261 -1080 0 1
rlabel polysilicon 264 -1080 264 -1080 0 2
rlabel polysilicon 261 -1086 261 -1086 0 3
rlabel polysilicon 264 -1086 264 -1086 0 4
rlabel polysilicon 268 -1080 268 -1080 0 1
rlabel polysilicon 268 -1086 268 -1086 0 3
rlabel polysilicon 275 -1080 275 -1080 0 1
rlabel polysilicon 275 -1086 275 -1086 0 3
rlabel polysilicon 282 -1080 282 -1080 0 1
rlabel polysilicon 282 -1086 282 -1086 0 3
rlabel polysilicon 289 -1080 289 -1080 0 1
rlabel polysilicon 289 -1086 289 -1086 0 3
rlabel polysilicon 296 -1080 296 -1080 0 1
rlabel polysilicon 296 -1086 296 -1086 0 3
rlabel polysilicon 303 -1080 303 -1080 0 1
rlabel polysilicon 306 -1080 306 -1080 0 2
rlabel polysilicon 303 -1086 303 -1086 0 3
rlabel polysilicon 310 -1080 310 -1080 0 1
rlabel polysilicon 310 -1086 310 -1086 0 3
rlabel polysilicon 317 -1080 317 -1080 0 1
rlabel polysilicon 317 -1086 317 -1086 0 3
rlabel polysilicon 324 -1080 324 -1080 0 1
rlabel polysilicon 324 -1086 324 -1086 0 3
rlabel polysilicon 331 -1080 331 -1080 0 1
rlabel polysilicon 331 -1086 331 -1086 0 3
rlabel polysilicon 338 -1080 338 -1080 0 1
rlabel polysilicon 341 -1080 341 -1080 0 2
rlabel polysilicon 341 -1086 341 -1086 0 4
rlabel polysilicon 345 -1080 345 -1080 0 1
rlabel polysilicon 345 -1086 345 -1086 0 3
rlabel polysilicon 352 -1080 352 -1080 0 1
rlabel polysilicon 352 -1086 352 -1086 0 3
rlabel polysilicon 359 -1080 359 -1080 0 1
rlabel polysilicon 359 -1086 359 -1086 0 3
rlabel polysilicon 366 -1080 366 -1080 0 1
rlabel polysilicon 366 -1086 366 -1086 0 3
rlabel polysilicon 373 -1080 373 -1080 0 1
rlabel polysilicon 376 -1080 376 -1080 0 2
rlabel polysilicon 373 -1086 373 -1086 0 3
rlabel polysilicon 376 -1086 376 -1086 0 4
rlabel polysilicon 380 -1080 380 -1080 0 1
rlabel polysilicon 380 -1086 380 -1086 0 3
rlabel polysilicon 387 -1080 387 -1080 0 1
rlabel polysilicon 387 -1086 387 -1086 0 3
rlabel polysilicon 394 -1080 394 -1080 0 1
rlabel polysilicon 394 -1086 394 -1086 0 3
rlabel polysilicon 401 -1080 401 -1080 0 1
rlabel polysilicon 401 -1086 401 -1086 0 3
rlabel polysilicon 408 -1080 408 -1080 0 1
rlabel polysilicon 408 -1086 408 -1086 0 3
rlabel polysilicon 415 -1080 415 -1080 0 1
rlabel polysilicon 415 -1086 415 -1086 0 3
rlabel polysilicon 422 -1080 422 -1080 0 1
rlabel polysilicon 422 -1086 422 -1086 0 3
rlabel polysilicon 429 -1080 429 -1080 0 1
rlabel polysilicon 429 -1086 429 -1086 0 3
rlabel polysilicon 436 -1080 436 -1080 0 1
rlabel polysilicon 439 -1080 439 -1080 0 2
rlabel polysilicon 436 -1086 436 -1086 0 3
rlabel polysilicon 439 -1086 439 -1086 0 4
rlabel polysilicon 443 -1080 443 -1080 0 1
rlabel polysilicon 443 -1086 443 -1086 0 3
rlabel polysilicon 450 -1080 450 -1080 0 1
rlabel polysilicon 450 -1086 450 -1086 0 3
rlabel polysilicon 457 -1080 457 -1080 0 1
rlabel polysilicon 457 -1086 457 -1086 0 3
rlabel polysilicon 464 -1080 464 -1080 0 1
rlabel polysilicon 464 -1086 464 -1086 0 3
rlabel polysilicon 471 -1080 471 -1080 0 1
rlabel polysilicon 471 -1086 471 -1086 0 3
rlabel polysilicon 478 -1080 478 -1080 0 1
rlabel polysilicon 481 -1080 481 -1080 0 2
rlabel polysilicon 478 -1086 478 -1086 0 3
rlabel polysilicon 481 -1086 481 -1086 0 4
rlabel polysilicon 485 -1080 485 -1080 0 1
rlabel polysilicon 485 -1086 485 -1086 0 3
rlabel polysilicon 492 -1080 492 -1080 0 1
rlabel polysilicon 495 -1080 495 -1080 0 2
rlabel polysilicon 492 -1086 492 -1086 0 3
rlabel polysilicon 495 -1086 495 -1086 0 4
rlabel polysilicon 499 -1080 499 -1080 0 1
rlabel polysilicon 502 -1080 502 -1080 0 2
rlabel polysilicon 499 -1086 499 -1086 0 3
rlabel polysilicon 502 -1086 502 -1086 0 4
rlabel polysilicon 506 -1080 506 -1080 0 1
rlabel polysilicon 506 -1086 506 -1086 0 3
rlabel polysilicon 513 -1080 513 -1080 0 1
rlabel polysilicon 516 -1080 516 -1080 0 2
rlabel polysilicon 513 -1086 513 -1086 0 3
rlabel polysilicon 516 -1086 516 -1086 0 4
rlabel polysilicon 520 -1080 520 -1080 0 1
rlabel polysilicon 520 -1086 520 -1086 0 3
rlabel polysilicon 527 -1080 527 -1080 0 1
rlabel polysilicon 530 -1080 530 -1080 0 2
rlabel polysilicon 527 -1086 527 -1086 0 3
rlabel polysilicon 530 -1086 530 -1086 0 4
rlabel polysilicon 534 -1080 534 -1080 0 1
rlabel polysilicon 534 -1086 534 -1086 0 3
rlabel polysilicon 541 -1080 541 -1080 0 1
rlabel polysilicon 541 -1086 541 -1086 0 3
rlabel polysilicon 548 -1080 548 -1080 0 1
rlabel polysilicon 548 -1086 548 -1086 0 3
rlabel polysilicon 558 -1080 558 -1080 0 2
rlabel polysilicon 555 -1086 555 -1086 0 3
rlabel polysilicon 558 -1086 558 -1086 0 4
rlabel polysilicon 565 -1080 565 -1080 0 2
rlabel polysilicon 562 -1086 562 -1086 0 3
rlabel polysilicon 565 -1086 565 -1086 0 4
rlabel polysilicon 569 -1080 569 -1080 0 1
rlabel polysilicon 572 -1080 572 -1080 0 2
rlabel polysilicon 569 -1086 569 -1086 0 3
rlabel polysilicon 572 -1086 572 -1086 0 4
rlabel polysilicon 576 -1080 576 -1080 0 1
rlabel polysilicon 576 -1086 576 -1086 0 3
rlabel polysilicon 583 -1080 583 -1080 0 1
rlabel polysilicon 583 -1086 583 -1086 0 3
rlabel polysilicon 590 -1080 590 -1080 0 1
rlabel polysilicon 590 -1086 590 -1086 0 3
rlabel polysilicon 597 -1080 597 -1080 0 1
rlabel polysilicon 597 -1086 597 -1086 0 3
rlabel polysilicon 604 -1080 604 -1080 0 1
rlabel polysilicon 604 -1086 604 -1086 0 3
rlabel polysilicon 611 -1080 611 -1080 0 1
rlabel polysilicon 611 -1086 611 -1086 0 3
rlabel polysilicon 618 -1080 618 -1080 0 1
rlabel polysilicon 618 -1086 618 -1086 0 3
rlabel polysilicon 625 -1080 625 -1080 0 1
rlabel polysilicon 628 -1080 628 -1080 0 2
rlabel polysilicon 625 -1086 625 -1086 0 3
rlabel polysilicon 635 -1080 635 -1080 0 2
rlabel polysilicon 632 -1086 632 -1086 0 3
rlabel polysilicon 635 -1086 635 -1086 0 4
rlabel polysilicon 639 -1080 639 -1080 0 1
rlabel polysilicon 639 -1086 639 -1086 0 3
rlabel polysilicon 646 -1080 646 -1080 0 1
rlabel polysilicon 646 -1086 646 -1086 0 3
rlabel polysilicon 653 -1080 653 -1080 0 1
rlabel polysilicon 653 -1086 653 -1086 0 3
rlabel polysilicon 660 -1080 660 -1080 0 1
rlabel polysilicon 660 -1086 660 -1086 0 3
rlabel polysilicon 667 -1080 667 -1080 0 1
rlabel polysilicon 667 -1086 667 -1086 0 3
rlabel polysilicon 674 -1080 674 -1080 0 1
rlabel polysilicon 677 -1080 677 -1080 0 2
rlabel polysilicon 674 -1086 674 -1086 0 3
rlabel polysilicon 677 -1086 677 -1086 0 4
rlabel polysilicon 681 -1080 681 -1080 0 1
rlabel polysilicon 681 -1086 681 -1086 0 3
rlabel polysilicon 688 -1080 688 -1080 0 1
rlabel polysilicon 688 -1086 688 -1086 0 3
rlabel polysilicon 695 -1080 695 -1080 0 1
rlabel polysilicon 695 -1086 695 -1086 0 3
rlabel polysilicon 702 -1080 702 -1080 0 1
rlabel polysilicon 702 -1086 702 -1086 0 3
rlabel polysilicon 709 -1080 709 -1080 0 1
rlabel polysilicon 709 -1086 709 -1086 0 3
rlabel polysilicon 716 -1080 716 -1080 0 1
rlabel polysilicon 716 -1086 716 -1086 0 3
rlabel polysilicon 723 -1080 723 -1080 0 1
rlabel polysilicon 726 -1080 726 -1080 0 2
rlabel polysilicon 723 -1086 723 -1086 0 3
rlabel polysilicon 726 -1086 726 -1086 0 4
rlabel polysilicon 730 -1080 730 -1080 0 1
rlabel polysilicon 730 -1086 730 -1086 0 3
rlabel polysilicon 737 -1080 737 -1080 0 1
rlabel polysilicon 737 -1086 737 -1086 0 3
rlabel polysilicon 744 -1080 744 -1080 0 1
rlabel polysilicon 747 -1080 747 -1080 0 2
rlabel polysilicon 744 -1086 744 -1086 0 3
rlabel polysilicon 747 -1086 747 -1086 0 4
rlabel polysilicon 751 -1080 751 -1080 0 1
rlabel polysilicon 751 -1086 751 -1086 0 3
rlabel polysilicon 758 -1080 758 -1080 0 1
rlabel polysilicon 758 -1086 758 -1086 0 3
rlabel polysilicon 765 -1080 765 -1080 0 1
rlabel polysilicon 765 -1086 765 -1086 0 3
rlabel polysilicon 772 -1080 772 -1080 0 1
rlabel polysilicon 772 -1086 772 -1086 0 3
rlabel polysilicon 779 -1080 779 -1080 0 1
rlabel polysilicon 779 -1086 779 -1086 0 3
rlabel polysilicon 786 -1080 786 -1080 0 1
rlabel polysilicon 786 -1086 786 -1086 0 3
rlabel polysilicon 793 -1080 793 -1080 0 1
rlabel polysilicon 793 -1086 793 -1086 0 3
rlabel polysilicon 800 -1080 800 -1080 0 1
rlabel polysilicon 800 -1086 800 -1086 0 3
rlabel polysilicon 807 -1080 807 -1080 0 1
rlabel polysilicon 807 -1086 807 -1086 0 3
rlabel polysilicon 814 -1080 814 -1080 0 1
rlabel polysilicon 814 -1086 814 -1086 0 3
rlabel polysilicon 821 -1080 821 -1080 0 1
rlabel polysilicon 821 -1086 821 -1086 0 3
rlabel polysilicon 828 -1080 828 -1080 0 1
rlabel polysilicon 828 -1086 828 -1086 0 3
rlabel polysilicon 835 -1080 835 -1080 0 1
rlabel polysilicon 835 -1086 835 -1086 0 3
rlabel polysilicon 842 -1080 842 -1080 0 1
rlabel polysilicon 842 -1086 842 -1086 0 3
rlabel polysilicon 849 -1080 849 -1080 0 1
rlabel polysilicon 849 -1086 849 -1086 0 3
rlabel polysilicon 856 -1080 856 -1080 0 1
rlabel polysilicon 856 -1086 856 -1086 0 3
rlabel polysilicon 863 -1080 863 -1080 0 1
rlabel polysilicon 866 -1080 866 -1080 0 2
rlabel polysilicon 863 -1086 863 -1086 0 3
rlabel polysilicon 866 -1086 866 -1086 0 4
rlabel polysilicon 870 -1080 870 -1080 0 1
rlabel polysilicon 870 -1086 870 -1086 0 3
rlabel polysilicon 877 -1080 877 -1080 0 1
rlabel polysilicon 877 -1086 877 -1086 0 3
rlabel polysilicon 884 -1080 884 -1080 0 1
rlabel polysilicon 884 -1086 884 -1086 0 3
rlabel polysilicon 891 -1080 891 -1080 0 1
rlabel polysilicon 891 -1086 891 -1086 0 3
rlabel polysilicon 898 -1080 898 -1080 0 1
rlabel polysilicon 898 -1086 898 -1086 0 3
rlabel polysilicon 905 -1080 905 -1080 0 1
rlabel polysilicon 905 -1086 905 -1086 0 3
rlabel polysilicon 912 -1080 912 -1080 0 1
rlabel polysilicon 912 -1086 912 -1086 0 3
rlabel polysilicon 919 -1080 919 -1080 0 1
rlabel polysilicon 919 -1086 919 -1086 0 3
rlabel polysilicon 926 -1080 926 -1080 0 1
rlabel polysilicon 929 -1080 929 -1080 0 2
rlabel polysilicon 929 -1086 929 -1086 0 4
rlabel polysilicon 933 -1080 933 -1080 0 1
rlabel polysilicon 933 -1086 933 -1086 0 3
rlabel polysilicon 940 -1080 940 -1080 0 1
rlabel polysilicon 940 -1086 940 -1086 0 3
rlabel polysilicon 947 -1080 947 -1080 0 1
rlabel polysilicon 947 -1086 947 -1086 0 3
rlabel polysilicon 954 -1080 954 -1080 0 1
rlabel polysilicon 954 -1086 954 -1086 0 3
rlabel polysilicon 961 -1080 961 -1080 0 1
rlabel polysilicon 961 -1086 961 -1086 0 3
rlabel polysilicon 968 -1080 968 -1080 0 1
rlabel polysilicon 968 -1086 968 -1086 0 3
rlabel polysilicon 975 -1080 975 -1080 0 1
rlabel polysilicon 975 -1086 975 -1086 0 3
rlabel polysilicon 982 -1080 982 -1080 0 1
rlabel polysilicon 982 -1086 982 -1086 0 3
rlabel polysilicon 989 -1080 989 -1080 0 1
rlabel polysilicon 989 -1086 989 -1086 0 3
rlabel polysilicon 996 -1080 996 -1080 0 1
rlabel polysilicon 996 -1086 996 -1086 0 3
rlabel polysilicon 1003 -1080 1003 -1080 0 1
rlabel polysilicon 1003 -1086 1003 -1086 0 3
rlabel polysilicon 1010 -1080 1010 -1080 0 1
rlabel polysilicon 1010 -1086 1010 -1086 0 3
rlabel polysilicon 1017 -1080 1017 -1080 0 1
rlabel polysilicon 1017 -1086 1017 -1086 0 3
rlabel polysilicon 1024 -1080 1024 -1080 0 1
rlabel polysilicon 1024 -1086 1024 -1086 0 3
rlabel polysilicon 1031 -1080 1031 -1080 0 1
rlabel polysilicon 1031 -1086 1031 -1086 0 3
rlabel polysilicon 1038 -1080 1038 -1080 0 1
rlabel polysilicon 1038 -1086 1038 -1086 0 3
rlabel polysilicon 1045 -1080 1045 -1080 0 1
rlabel polysilicon 1045 -1086 1045 -1086 0 3
rlabel polysilicon 1052 -1080 1052 -1080 0 1
rlabel polysilicon 1052 -1086 1052 -1086 0 3
rlabel polysilicon 1059 -1080 1059 -1080 0 1
rlabel polysilicon 1059 -1086 1059 -1086 0 3
rlabel polysilicon 1066 -1080 1066 -1080 0 1
rlabel polysilicon 1066 -1086 1066 -1086 0 3
rlabel polysilicon 1073 -1080 1073 -1080 0 1
rlabel polysilicon 1073 -1086 1073 -1086 0 3
rlabel polysilicon 1080 -1080 1080 -1080 0 1
rlabel polysilicon 1080 -1086 1080 -1086 0 3
rlabel polysilicon 1087 -1080 1087 -1080 0 1
rlabel polysilicon 1087 -1086 1087 -1086 0 3
rlabel polysilicon 1094 -1080 1094 -1080 0 1
rlabel polysilicon 1094 -1086 1094 -1086 0 3
rlabel polysilicon 1101 -1080 1101 -1080 0 1
rlabel polysilicon 1101 -1086 1101 -1086 0 3
rlabel polysilicon 1108 -1080 1108 -1080 0 1
rlabel polysilicon 1108 -1086 1108 -1086 0 3
rlabel polysilicon 1115 -1080 1115 -1080 0 1
rlabel polysilicon 1115 -1086 1115 -1086 0 3
rlabel polysilicon 1122 -1080 1122 -1080 0 1
rlabel polysilicon 1122 -1086 1122 -1086 0 3
rlabel polysilicon 1129 -1080 1129 -1080 0 1
rlabel polysilicon 1129 -1086 1129 -1086 0 3
rlabel polysilicon 1136 -1080 1136 -1080 0 1
rlabel polysilicon 1136 -1086 1136 -1086 0 3
rlabel polysilicon 1143 -1080 1143 -1080 0 1
rlabel polysilicon 1143 -1086 1143 -1086 0 3
rlabel polysilicon 1150 -1080 1150 -1080 0 1
rlabel polysilicon 1150 -1086 1150 -1086 0 3
rlabel polysilicon 1157 -1080 1157 -1080 0 1
rlabel polysilicon 1157 -1086 1157 -1086 0 3
rlabel polysilicon 1164 -1080 1164 -1080 0 1
rlabel polysilicon 1164 -1086 1164 -1086 0 3
rlabel polysilicon 1171 -1080 1171 -1080 0 1
rlabel polysilicon 1171 -1086 1171 -1086 0 3
rlabel polysilicon 1178 -1080 1178 -1080 0 1
rlabel polysilicon 1178 -1086 1178 -1086 0 3
rlabel polysilicon 1185 -1080 1185 -1080 0 1
rlabel polysilicon 1185 -1086 1185 -1086 0 3
rlabel polysilicon 1192 -1080 1192 -1080 0 1
rlabel polysilicon 1192 -1086 1192 -1086 0 3
rlabel polysilicon 1199 -1080 1199 -1080 0 1
rlabel polysilicon 1199 -1086 1199 -1086 0 3
rlabel polysilicon 1206 -1080 1206 -1080 0 1
rlabel polysilicon 1206 -1086 1206 -1086 0 3
rlabel polysilicon 1213 -1080 1213 -1080 0 1
rlabel polysilicon 1213 -1086 1213 -1086 0 3
rlabel polysilicon 1220 -1080 1220 -1080 0 1
rlabel polysilicon 1220 -1086 1220 -1086 0 3
rlabel polysilicon 1227 -1080 1227 -1080 0 1
rlabel polysilicon 1227 -1086 1227 -1086 0 3
rlabel polysilicon 1234 -1080 1234 -1080 0 1
rlabel polysilicon 1234 -1086 1234 -1086 0 3
rlabel polysilicon 1241 -1080 1241 -1080 0 1
rlabel polysilicon 1241 -1086 1241 -1086 0 3
rlabel polysilicon 1248 -1080 1248 -1080 0 1
rlabel polysilicon 1248 -1086 1248 -1086 0 3
rlabel polysilicon 1255 -1080 1255 -1080 0 1
rlabel polysilicon 1255 -1086 1255 -1086 0 3
rlabel polysilicon 1262 -1080 1262 -1080 0 1
rlabel polysilicon 1262 -1086 1262 -1086 0 3
rlabel polysilicon 1269 -1080 1269 -1080 0 1
rlabel polysilicon 1269 -1086 1269 -1086 0 3
rlabel polysilicon 1276 -1080 1276 -1080 0 1
rlabel polysilicon 1276 -1086 1276 -1086 0 3
rlabel polysilicon 1283 -1080 1283 -1080 0 1
rlabel polysilicon 1283 -1086 1283 -1086 0 3
rlabel polysilicon 1290 -1080 1290 -1080 0 1
rlabel polysilicon 1290 -1086 1290 -1086 0 3
rlabel polysilicon 1297 -1080 1297 -1080 0 1
rlabel polysilicon 1297 -1086 1297 -1086 0 3
rlabel polysilicon 1304 -1080 1304 -1080 0 1
rlabel polysilicon 1304 -1086 1304 -1086 0 3
rlabel polysilicon 1311 -1080 1311 -1080 0 1
rlabel polysilicon 1311 -1086 1311 -1086 0 3
rlabel polysilicon 1318 -1080 1318 -1080 0 1
rlabel polysilicon 1318 -1086 1318 -1086 0 3
rlabel polysilicon 1325 -1080 1325 -1080 0 1
rlabel polysilicon 1325 -1086 1325 -1086 0 3
rlabel polysilicon 1332 -1080 1332 -1080 0 1
rlabel polysilicon 1332 -1086 1332 -1086 0 3
rlabel polysilicon 1339 -1080 1339 -1080 0 1
rlabel polysilicon 1339 -1086 1339 -1086 0 3
rlabel polysilicon 1346 -1080 1346 -1080 0 1
rlabel polysilicon 1346 -1086 1346 -1086 0 3
rlabel polysilicon 1444 -1080 1444 -1080 0 1
rlabel polysilicon 1444 -1086 1444 -1086 0 3
rlabel polysilicon 2 -1205 2 -1205 0 1
rlabel polysilicon 5 -1205 5 -1205 0 2
rlabel polysilicon 5 -1211 5 -1211 0 4
rlabel polysilicon 9 -1205 9 -1205 0 1
rlabel polysilicon 9 -1211 9 -1211 0 3
rlabel polysilicon 16 -1205 16 -1205 0 1
rlabel polysilicon 16 -1211 16 -1211 0 3
rlabel polysilicon 23 -1205 23 -1205 0 1
rlabel polysilicon 23 -1211 23 -1211 0 3
rlabel polysilicon 30 -1205 30 -1205 0 1
rlabel polysilicon 30 -1211 30 -1211 0 3
rlabel polysilicon 37 -1205 37 -1205 0 1
rlabel polysilicon 37 -1211 37 -1211 0 3
rlabel polysilicon 44 -1205 44 -1205 0 1
rlabel polysilicon 44 -1211 44 -1211 0 3
rlabel polysilicon 51 -1205 51 -1205 0 1
rlabel polysilicon 51 -1211 51 -1211 0 3
rlabel polysilicon 58 -1205 58 -1205 0 1
rlabel polysilicon 58 -1211 58 -1211 0 3
rlabel polysilicon 65 -1205 65 -1205 0 1
rlabel polysilicon 65 -1211 65 -1211 0 3
rlabel polysilicon 72 -1205 72 -1205 0 1
rlabel polysilicon 75 -1205 75 -1205 0 2
rlabel polysilicon 75 -1211 75 -1211 0 4
rlabel polysilicon 79 -1205 79 -1205 0 1
rlabel polysilicon 79 -1211 79 -1211 0 3
rlabel polysilicon 86 -1205 86 -1205 0 1
rlabel polysilicon 86 -1211 86 -1211 0 3
rlabel polysilicon 93 -1205 93 -1205 0 1
rlabel polysilicon 93 -1211 93 -1211 0 3
rlabel polysilicon 100 -1205 100 -1205 0 1
rlabel polysilicon 103 -1205 103 -1205 0 2
rlabel polysilicon 103 -1211 103 -1211 0 4
rlabel polysilicon 107 -1205 107 -1205 0 1
rlabel polysilicon 107 -1211 107 -1211 0 3
rlabel polysilicon 114 -1205 114 -1205 0 1
rlabel polysilicon 117 -1205 117 -1205 0 2
rlabel polysilicon 114 -1211 114 -1211 0 3
rlabel polysilicon 117 -1211 117 -1211 0 4
rlabel polysilicon 121 -1205 121 -1205 0 1
rlabel polysilicon 121 -1211 121 -1211 0 3
rlabel polysilicon 128 -1205 128 -1205 0 1
rlabel polysilicon 128 -1211 128 -1211 0 3
rlabel polysilicon 135 -1205 135 -1205 0 1
rlabel polysilicon 135 -1211 135 -1211 0 3
rlabel polysilicon 142 -1205 142 -1205 0 1
rlabel polysilicon 142 -1211 142 -1211 0 3
rlabel polysilicon 149 -1205 149 -1205 0 1
rlabel polysilicon 149 -1211 149 -1211 0 3
rlabel polysilicon 156 -1205 156 -1205 0 1
rlabel polysilicon 156 -1211 156 -1211 0 3
rlabel polysilicon 163 -1205 163 -1205 0 1
rlabel polysilicon 163 -1211 163 -1211 0 3
rlabel polysilicon 170 -1205 170 -1205 0 1
rlabel polysilicon 170 -1211 170 -1211 0 3
rlabel polysilicon 177 -1205 177 -1205 0 1
rlabel polysilicon 180 -1205 180 -1205 0 2
rlabel polysilicon 184 -1205 184 -1205 0 1
rlabel polysilicon 184 -1211 184 -1211 0 3
rlabel polysilicon 191 -1205 191 -1205 0 1
rlabel polysilicon 191 -1211 191 -1211 0 3
rlabel polysilicon 198 -1205 198 -1205 0 1
rlabel polysilicon 198 -1211 198 -1211 0 3
rlabel polysilicon 205 -1205 205 -1205 0 1
rlabel polysilicon 205 -1211 205 -1211 0 3
rlabel polysilicon 212 -1205 212 -1205 0 1
rlabel polysilicon 215 -1205 215 -1205 0 2
rlabel polysilicon 212 -1211 212 -1211 0 3
rlabel polysilicon 219 -1205 219 -1205 0 1
rlabel polysilicon 219 -1211 219 -1211 0 3
rlabel polysilicon 226 -1205 226 -1205 0 1
rlabel polysilicon 226 -1211 226 -1211 0 3
rlabel polysilicon 233 -1205 233 -1205 0 1
rlabel polysilicon 233 -1211 233 -1211 0 3
rlabel polysilicon 240 -1205 240 -1205 0 1
rlabel polysilicon 240 -1211 240 -1211 0 3
rlabel polysilicon 247 -1205 247 -1205 0 1
rlabel polysilicon 247 -1211 247 -1211 0 3
rlabel polysilicon 254 -1205 254 -1205 0 1
rlabel polysilicon 254 -1211 254 -1211 0 3
rlabel polysilicon 261 -1205 261 -1205 0 1
rlabel polysilicon 261 -1211 261 -1211 0 3
rlabel polysilicon 268 -1205 268 -1205 0 1
rlabel polysilicon 268 -1211 268 -1211 0 3
rlabel polysilicon 275 -1205 275 -1205 0 1
rlabel polysilicon 275 -1211 275 -1211 0 3
rlabel polysilicon 282 -1205 282 -1205 0 1
rlabel polysilicon 282 -1211 282 -1211 0 3
rlabel polysilicon 289 -1205 289 -1205 0 1
rlabel polysilicon 289 -1211 289 -1211 0 3
rlabel polysilicon 296 -1205 296 -1205 0 1
rlabel polysilicon 296 -1211 296 -1211 0 3
rlabel polysilicon 303 -1205 303 -1205 0 1
rlabel polysilicon 303 -1211 303 -1211 0 3
rlabel polysilicon 310 -1205 310 -1205 0 1
rlabel polysilicon 310 -1211 310 -1211 0 3
rlabel polysilicon 317 -1205 317 -1205 0 1
rlabel polysilicon 317 -1211 317 -1211 0 3
rlabel polysilicon 324 -1205 324 -1205 0 1
rlabel polysilicon 324 -1211 324 -1211 0 3
rlabel polysilicon 331 -1205 331 -1205 0 1
rlabel polysilicon 331 -1211 331 -1211 0 3
rlabel polysilicon 338 -1205 338 -1205 0 1
rlabel polysilicon 338 -1211 338 -1211 0 3
rlabel polysilicon 345 -1205 345 -1205 0 1
rlabel polysilicon 345 -1211 345 -1211 0 3
rlabel polysilicon 352 -1205 352 -1205 0 1
rlabel polysilicon 352 -1211 352 -1211 0 3
rlabel polysilicon 359 -1205 359 -1205 0 1
rlabel polysilicon 359 -1211 359 -1211 0 3
rlabel polysilicon 366 -1205 366 -1205 0 1
rlabel polysilicon 366 -1211 366 -1211 0 3
rlabel polysilicon 373 -1205 373 -1205 0 1
rlabel polysilicon 373 -1211 373 -1211 0 3
rlabel polysilicon 380 -1205 380 -1205 0 1
rlabel polysilicon 380 -1211 380 -1211 0 3
rlabel polysilicon 387 -1205 387 -1205 0 1
rlabel polysilicon 387 -1211 387 -1211 0 3
rlabel polysilicon 394 -1205 394 -1205 0 1
rlabel polysilicon 394 -1211 394 -1211 0 3
rlabel polysilicon 401 -1205 401 -1205 0 1
rlabel polysilicon 404 -1205 404 -1205 0 2
rlabel polysilicon 401 -1211 401 -1211 0 3
rlabel polysilicon 404 -1211 404 -1211 0 4
rlabel polysilicon 408 -1205 408 -1205 0 1
rlabel polysilicon 408 -1211 408 -1211 0 3
rlabel polysilicon 415 -1205 415 -1205 0 1
rlabel polysilicon 415 -1211 415 -1211 0 3
rlabel polysilicon 422 -1205 422 -1205 0 1
rlabel polysilicon 422 -1211 422 -1211 0 3
rlabel polysilicon 429 -1205 429 -1205 0 1
rlabel polysilicon 429 -1211 429 -1211 0 3
rlabel polysilicon 436 -1205 436 -1205 0 1
rlabel polysilicon 436 -1211 436 -1211 0 3
rlabel polysilicon 443 -1205 443 -1205 0 1
rlabel polysilicon 443 -1211 443 -1211 0 3
rlabel polysilicon 450 -1205 450 -1205 0 1
rlabel polysilicon 450 -1211 450 -1211 0 3
rlabel polysilicon 457 -1205 457 -1205 0 1
rlabel polysilicon 457 -1211 457 -1211 0 3
rlabel polysilicon 464 -1205 464 -1205 0 1
rlabel polysilicon 467 -1205 467 -1205 0 2
rlabel polysilicon 464 -1211 464 -1211 0 3
rlabel polysilicon 467 -1211 467 -1211 0 4
rlabel polysilicon 471 -1205 471 -1205 0 1
rlabel polysilicon 471 -1211 471 -1211 0 3
rlabel polysilicon 478 -1205 478 -1205 0 1
rlabel polysilicon 478 -1211 478 -1211 0 3
rlabel polysilicon 485 -1205 485 -1205 0 1
rlabel polysilicon 485 -1211 485 -1211 0 3
rlabel polysilicon 492 -1205 492 -1205 0 1
rlabel polysilicon 495 -1205 495 -1205 0 2
rlabel polysilicon 492 -1211 492 -1211 0 3
rlabel polysilicon 495 -1211 495 -1211 0 4
rlabel polysilicon 499 -1205 499 -1205 0 1
rlabel polysilicon 499 -1211 499 -1211 0 3
rlabel polysilicon 506 -1205 506 -1205 0 1
rlabel polysilicon 506 -1211 506 -1211 0 3
rlabel polysilicon 513 -1205 513 -1205 0 1
rlabel polysilicon 513 -1211 513 -1211 0 3
rlabel polysilicon 523 -1205 523 -1205 0 2
rlabel polysilicon 520 -1211 520 -1211 0 3
rlabel polysilicon 523 -1211 523 -1211 0 4
rlabel polysilicon 527 -1205 527 -1205 0 1
rlabel polysilicon 530 -1205 530 -1205 0 2
rlabel polysilicon 527 -1211 527 -1211 0 3
rlabel polysilicon 530 -1211 530 -1211 0 4
rlabel polysilicon 534 -1205 534 -1205 0 1
rlabel polysilicon 534 -1211 534 -1211 0 3
rlabel polysilicon 541 -1205 541 -1205 0 1
rlabel polysilicon 544 -1205 544 -1205 0 2
rlabel polysilicon 541 -1211 541 -1211 0 3
rlabel polysilicon 544 -1211 544 -1211 0 4
rlabel polysilicon 551 -1205 551 -1205 0 2
rlabel polysilicon 548 -1211 548 -1211 0 3
rlabel polysilicon 551 -1211 551 -1211 0 4
rlabel polysilicon 555 -1205 555 -1205 0 1
rlabel polysilicon 558 -1205 558 -1205 0 2
rlabel polysilicon 555 -1211 555 -1211 0 3
rlabel polysilicon 558 -1211 558 -1211 0 4
rlabel polysilicon 562 -1205 562 -1205 0 1
rlabel polysilicon 562 -1211 562 -1211 0 3
rlabel polysilicon 569 -1205 569 -1205 0 1
rlabel polysilicon 569 -1211 569 -1211 0 3
rlabel polysilicon 576 -1205 576 -1205 0 1
rlabel polysilicon 576 -1211 576 -1211 0 3
rlabel polysilicon 583 -1205 583 -1205 0 1
rlabel polysilicon 583 -1211 583 -1211 0 3
rlabel polysilicon 590 -1205 590 -1205 0 1
rlabel polysilicon 590 -1211 590 -1211 0 3
rlabel polysilicon 597 -1205 597 -1205 0 1
rlabel polysilicon 600 -1205 600 -1205 0 2
rlabel polysilicon 597 -1211 597 -1211 0 3
rlabel polysilicon 600 -1211 600 -1211 0 4
rlabel polysilicon 607 -1205 607 -1205 0 2
rlabel polysilicon 604 -1211 604 -1211 0 3
rlabel polysilicon 607 -1211 607 -1211 0 4
rlabel polysilicon 611 -1205 611 -1205 0 1
rlabel polysilicon 611 -1211 611 -1211 0 3
rlabel polysilicon 618 -1205 618 -1205 0 1
rlabel polysilicon 618 -1211 618 -1211 0 3
rlabel polysilicon 625 -1205 625 -1205 0 1
rlabel polysilicon 628 -1205 628 -1205 0 2
rlabel polysilicon 625 -1211 625 -1211 0 3
rlabel polysilicon 628 -1211 628 -1211 0 4
rlabel polysilicon 632 -1205 632 -1205 0 1
rlabel polysilicon 635 -1205 635 -1205 0 2
rlabel polysilicon 632 -1211 632 -1211 0 3
rlabel polysilicon 639 -1205 639 -1205 0 1
rlabel polysilicon 639 -1211 639 -1211 0 3
rlabel polysilicon 646 -1205 646 -1205 0 1
rlabel polysilicon 649 -1205 649 -1205 0 2
rlabel polysilicon 646 -1211 646 -1211 0 3
rlabel polysilicon 649 -1211 649 -1211 0 4
rlabel polysilicon 653 -1205 653 -1205 0 1
rlabel polysilicon 653 -1211 653 -1211 0 3
rlabel polysilicon 660 -1205 660 -1205 0 1
rlabel polysilicon 660 -1211 660 -1211 0 3
rlabel polysilicon 667 -1205 667 -1205 0 1
rlabel polysilicon 667 -1211 667 -1211 0 3
rlabel polysilicon 674 -1205 674 -1205 0 1
rlabel polysilicon 674 -1211 674 -1211 0 3
rlabel polysilicon 681 -1205 681 -1205 0 1
rlabel polysilicon 684 -1205 684 -1205 0 2
rlabel polysilicon 681 -1211 681 -1211 0 3
rlabel polysilicon 688 -1205 688 -1205 0 1
rlabel polysilicon 688 -1211 688 -1211 0 3
rlabel polysilicon 695 -1205 695 -1205 0 1
rlabel polysilicon 695 -1211 695 -1211 0 3
rlabel polysilicon 702 -1205 702 -1205 0 1
rlabel polysilicon 702 -1211 702 -1211 0 3
rlabel polysilicon 709 -1205 709 -1205 0 1
rlabel polysilicon 712 -1205 712 -1205 0 2
rlabel polysilicon 709 -1211 709 -1211 0 3
rlabel polysilicon 712 -1211 712 -1211 0 4
rlabel polysilicon 716 -1205 716 -1205 0 1
rlabel polysilicon 716 -1211 716 -1211 0 3
rlabel polysilicon 723 -1205 723 -1205 0 1
rlabel polysilicon 723 -1211 723 -1211 0 3
rlabel polysilicon 730 -1205 730 -1205 0 1
rlabel polysilicon 733 -1205 733 -1205 0 2
rlabel polysilicon 730 -1211 730 -1211 0 3
rlabel polysilicon 733 -1211 733 -1211 0 4
rlabel polysilicon 737 -1205 737 -1205 0 1
rlabel polysilicon 737 -1211 737 -1211 0 3
rlabel polysilicon 744 -1205 744 -1205 0 1
rlabel polysilicon 747 -1205 747 -1205 0 2
rlabel polysilicon 744 -1211 744 -1211 0 3
rlabel polysilicon 747 -1211 747 -1211 0 4
rlabel polysilicon 751 -1205 751 -1205 0 1
rlabel polysilicon 754 -1205 754 -1205 0 2
rlabel polysilicon 751 -1211 751 -1211 0 3
rlabel polysilicon 754 -1211 754 -1211 0 4
rlabel polysilicon 758 -1205 758 -1205 0 1
rlabel polysilicon 761 -1205 761 -1205 0 2
rlabel polysilicon 758 -1211 758 -1211 0 3
rlabel polysilicon 761 -1211 761 -1211 0 4
rlabel polysilicon 765 -1205 765 -1205 0 1
rlabel polysilicon 765 -1211 765 -1211 0 3
rlabel polysilicon 768 -1211 768 -1211 0 4
rlabel polysilicon 772 -1205 772 -1205 0 1
rlabel polysilicon 772 -1211 772 -1211 0 3
rlabel polysilicon 779 -1205 779 -1205 0 1
rlabel polysilicon 779 -1211 779 -1211 0 3
rlabel polysilicon 786 -1205 786 -1205 0 1
rlabel polysilicon 786 -1211 786 -1211 0 3
rlabel polysilicon 793 -1205 793 -1205 0 1
rlabel polysilicon 796 -1205 796 -1205 0 2
rlabel polysilicon 796 -1211 796 -1211 0 4
rlabel polysilicon 800 -1205 800 -1205 0 1
rlabel polysilicon 800 -1211 800 -1211 0 3
rlabel polysilicon 807 -1205 807 -1205 0 1
rlabel polysilicon 807 -1211 807 -1211 0 3
rlabel polysilicon 814 -1205 814 -1205 0 1
rlabel polysilicon 814 -1211 814 -1211 0 3
rlabel polysilicon 821 -1205 821 -1205 0 1
rlabel polysilicon 821 -1211 821 -1211 0 3
rlabel polysilicon 828 -1205 828 -1205 0 1
rlabel polysilicon 828 -1211 828 -1211 0 3
rlabel polysilicon 835 -1205 835 -1205 0 1
rlabel polysilicon 835 -1211 835 -1211 0 3
rlabel polysilicon 845 -1205 845 -1205 0 2
rlabel polysilicon 842 -1211 842 -1211 0 3
rlabel polysilicon 845 -1211 845 -1211 0 4
rlabel polysilicon 849 -1205 849 -1205 0 1
rlabel polysilicon 849 -1211 849 -1211 0 3
rlabel polysilicon 856 -1205 856 -1205 0 1
rlabel polysilicon 856 -1211 856 -1211 0 3
rlabel polysilicon 863 -1205 863 -1205 0 1
rlabel polysilicon 863 -1211 863 -1211 0 3
rlabel polysilicon 870 -1205 870 -1205 0 1
rlabel polysilicon 870 -1211 870 -1211 0 3
rlabel polysilicon 877 -1205 877 -1205 0 1
rlabel polysilicon 877 -1211 877 -1211 0 3
rlabel polysilicon 884 -1205 884 -1205 0 1
rlabel polysilicon 884 -1211 884 -1211 0 3
rlabel polysilicon 891 -1205 891 -1205 0 1
rlabel polysilicon 891 -1211 891 -1211 0 3
rlabel polysilicon 898 -1205 898 -1205 0 1
rlabel polysilicon 898 -1211 898 -1211 0 3
rlabel polysilicon 905 -1205 905 -1205 0 1
rlabel polysilicon 905 -1211 905 -1211 0 3
rlabel polysilicon 912 -1205 912 -1205 0 1
rlabel polysilicon 912 -1211 912 -1211 0 3
rlabel polysilicon 919 -1205 919 -1205 0 1
rlabel polysilicon 919 -1211 919 -1211 0 3
rlabel polysilicon 926 -1205 926 -1205 0 1
rlabel polysilicon 926 -1211 926 -1211 0 3
rlabel polysilicon 933 -1205 933 -1205 0 1
rlabel polysilicon 933 -1211 933 -1211 0 3
rlabel polysilicon 940 -1205 940 -1205 0 1
rlabel polysilicon 940 -1211 940 -1211 0 3
rlabel polysilicon 947 -1205 947 -1205 0 1
rlabel polysilicon 947 -1211 947 -1211 0 3
rlabel polysilicon 954 -1205 954 -1205 0 1
rlabel polysilicon 954 -1211 954 -1211 0 3
rlabel polysilicon 961 -1205 961 -1205 0 1
rlabel polysilicon 961 -1211 961 -1211 0 3
rlabel polysilicon 968 -1205 968 -1205 0 1
rlabel polysilicon 968 -1211 968 -1211 0 3
rlabel polysilicon 975 -1205 975 -1205 0 1
rlabel polysilicon 975 -1211 975 -1211 0 3
rlabel polysilicon 982 -1205 982 -1205 0 1
rlabel polysilicon 982 -1211 982 -1211 0 3
rlabel polysilicon 989 -1205 989 -1205 0 1
rlabel polysilicon 989 -1211 989 -1211 0 3
rlabel polysilicon 996 -1205 996 -1205 0 1
rlabel polysilicon 996 -1211 996 -1211 0 3
rlabel polysilicon 1003 -1205 1003 -1205 0 1
rlabel polysilicon 1003 -1211 1003 -1211 0 3
rlabel polysilicon 1010 -1205 1010 -1205 0 1
rlabel polysilicon 1010 -1211 1010 -1211 0 3
rlabel polysilicon 1017 -1205 1017 -1205 0 1
rlabel polysilicon 1017 -1211 1017 -1211 0 3
rlabel polysilicon 1024 -1205 1024 -1205 0 1
rlabel polysilicon 1024 -1211 1024 -1211 0 3
rlabel polysilicon 1031 -1205 1031 -1205 0 1
rlabel polysilicon 1031 -1211 1031 -1211 0 3
rlabel polysilicon 1038 -1205 1038 -1205 0 1
rlabel polysilicon 1038 -1211 1038 -1211 0 3
rlabel polysilicon 1045 -1205 1045 -1205 0 1
rlabel polysilicon 1045 -1211 1045 -1211 0 3
rlabel polysilicon 1052 -1205 1052 -1205 0 1
rlabel polysilicon 1052 -1211 1052 -1211 0 3
rlabel polysilicon 1059 -1205 1059 -1205 0 1
rlabel polysilicon 1059 -1211 1059 -1211 0 3
rlabel polysilicon 1066 -1205 1066 -1205 0 1
rlabel polysilicon 1066 -1211 1066 -1211 0 3
rlabel polysilicon 1073 -1205 1073 -1205 0 1
rlabel polysilicon 1073 -1211 1073 -1211 0 3
rlabel polysilicon 1080 -1205 1080 -1205 0 1
rlabel polysilicon 1080 -1211 1080 -1211 0 3
rlabel polysilicon 1087 -1205 1087 -1205 0 1
rlabel polysilicon 1087 -1211 1087 -1211 0 3
rlabel polysilicon 1094 -1205 1094 -1205 0 1
rlabel polysilicon 1094 -1211 1094 -1211 0 3
rlabel polysilicon 1101 -1205 1101 -1205 0 1
rlabel polysilicon 1101 -1211 1101 -1211 0 3
rlabel polysilicon 1108 -1205 1108 -1205 0 1
rlabel polysilicon 1108 -1211 1108 -1211 0 3
rlabel polysilicon 1115 -1205 1115 -1205 0 1
rlabel polysilicon 1122 -1205 1122 -1205 0 1
rlabel polysilicon 1122 -1211 1122 -1211 0 3
rlabel polysilicon 1129 -1205 1129 -1205 0 1
rlabel polysilicon 1129 -1211 1129 -1211 0 3
rlabel polysilicon 1136 -1205 1136 -1205 0 1
rlabel polysilicon 1136 -1211 1136 -1211 0 3
rlabel polysilicon 1143 -1205 1143 -1205 0 1
rlabel polysilicon 1143 -1211 1143 -1211 0 3
rlabel polysilicon 1150 -1205 1150 -1205 0 1
rlabel polysilicon 1150 -1211 1150 -1211 0 3
rlabel polysilicon 1157 -1205 1157 -1205 0 1
rlabel polysilicon 1157 -1211 1157 -1211 0 3
rlabel polysilicon 1164 -1205 1164 -1205 0 1
rlabel polysilicon 1164 -1211 1164 -1211 0 3
rlabel polysilicon 1171 -1205 1171 -1205 0 1
rlabel polysilicon 1171 -1211 1171 -1211 0 3
rlabel polysilicon 1178 -1205 1178 -1205 0 1
rlabel polysilicon 1178 -1211 1178 -1211 0 3
rlabel polysilicon 1185 -1205 1185 -1205 0 1
rlabel polysilicon 1185 -1211 1185 -1211 0 3
rlabel polysilicon 1192 -1205 1192 -1205 0 1
rlabel polysilicon 1192 -1211 1192 -1211 0 3
rlabel polysilicon 1199 -1205 1199 -1205 0 1
rlabel polysilicon 1199 -1211 1199 -1211 0 3
rlabel polysilicon 1206 -1205 1206 -1205 0 1
rlabel polysilicon 1206 -1211 1206 -1211 0 3
rlabel polysilicon 1213 -1205 1213 -1205 0 1
rlabel polysilicon 1213 -1211 1213 -1211 0 3
rlabel polysilicon 1220 -1205 1220 -1205 0 1
rlabel polysilicon 1220 -1211 1220 -1211 0 3
rlabel polysilicon 1227 -1205 1227 -1205 0 1
rlabel polysilicon 1227 -1211 1227 -1211 0 3
rlabel polysilicon 1234 -1205 1234 -1205 0 1
rlabel polysilicon 1234 -1211 1234 -1211 0 3
rlabel polysilicon 1241 -1205 1241 -1205 0 1
rlabel polysilicon 1241 -1211 1241 -1211 0 3
rlabel polysilicon 1248 -1205 1248 -1205 0 1
rlabel polysilicon 1248 -1211 1248 -1211 0 3
rlabel polysilicon 1255 -1205 1255 -1205 0 1
rlabel polysilicon 1255 -1211 1255 -1211 0 3
rlabel polysilicon 1262 -1205 1262 -1205 0 1
rlabel polysilicon 1262 -1211 1262 -1211 0 3
rlabel polysilicon 1269 -1205 1269 -1205 0 1
rlabel polysilicon 1269 -1211 1269 -1211 0 3
rlabel polysilicon 1272 -1211 1272 -1211 0 4
rlabel polysilicon 1276 -1205 1276 -1205 0 1
rlabel polysilicon 1276 -1211 1276 -1211 0 3
rlabel polysilicon 1283 -1205 1283 -1205 0 1
rlabel polysilicon 1283 -1211 1283 -1211 0 3
rlabel polysilicon 1290 -1205 1290 -1205 0 1
rlabel polysilicon 1290 -1211 1290 -1211 0 3
rlabel polysilicon 1297 -1205 1297 -1205 0 1
rlabel polysilicon 1297 -1211 1297 -1211 0 3
rlabel polysilicon 1304 -1205 1304 -1205 0 1
rlabel polysilicon 1304 -1211 1304 -1211 0 3
rlabel polysilicon 1311 -1205 1311 -1205 0 1
rlabel polysilicon 1311 -1211 1311 -1211 0 3
rlabel polysilicon 1318 -1205 1318 -1205 0 1
rlabel polysilicon 1318 -1211 1318 -1211 0 3
rlabel polysilicon 1325 -1205 1325 -1205 0 1
rlabel polysilicon 1325 -1211 1325 -1211 0 3
rlabel polysilicon 1332 -1205 1332 -1205 0 1
rlabel polysilicon 1332 -1211 1332 -1211 0 3
rlabel polysilicon 1339 -1205 1339 -1205 0 1
rlabel polysilicon 1339 -1211 1339 -1211 0 3
rlabel polysilicon 1346 -1205 1346 -1205 0 1
rlabel polysilicon 1346 -1211 1346 -1211 0 3
rlabel polysilicon 1353 -1205 1353 -1205 0 1
rlabel polysilicon 1353 -1211 1353 -1211 0 3
rlabel polysilicon 1360 -1205 1360 -1205 0 1
rlabel polysilicon 1360 -1211 1360 -1211 0 3
rlabel polysilicon 1367 -1205 1367 -1205 0 1
rlabel polysilicon 1367 -1211 1367 -1211 0 3
rlabel polysilicon 1374 -1205 1374 -1205 0 1
rlabel polysilicon 1374 -1211 1374 -1211 0 3
rlabel polysilicon 1451 -1205 1451 -1205 0 1
rlabel polysilicon 1451 -1211 1451 -1211 0 3
rlabel polysilicon 2 -1326 2 -1326 0 1
rlabel polysilicon 2 -1332 2 -1332 0 3
rlabel polysilicon 9 -1326 9 -1326 0 1
rlabel polysilicon 9 -1332 9 -1332 0 3
rlabel polysilicon 16 -1326 16 -1326 0 1
rlabel polysilicon 16 -1332 16 -1332 0 3
rlabel polysilicon 23 -1326 23 -1326 0 1
rlabel polysilicon 23 -1332 23 -1332 0 3
rlabel polysilicon 30 -1326 30 -1326 0 1
rlabel polysilicon 30 -1332 30 -1332 0 3
rlabel polysilicon 37 -1326 37 -1326 0 1
rlabel polysilicon 37 -1332 37 -1332 0 3
rlabel polysilicon 44 -1326 44 -1326 0 1
rlabel polysilicon 44 -1332 44 -1332 0 3
rlabel polysilicon 51 -1326 51 -1326 0 1
rlabel polysilicon 51 -1332 51 -1332 0 3
rlabel polysilicon 58 -1326 58 -1326 0 1
rlabel polysilicon 61 -1326 61 -1326 0 2
rlabel polysilicon 58 -1332 58 -1332 0 3
rlabel polysilicon 61 -1332 61 -1332 0 4
rlabel polysilicon 68 -1326 68 -1326 0 2
rlabel polysilicon 65 -1332 65 -1332 0 3
rlabel polysilicon 68 -1332 68 -1332 0 4
rlabel polysilicon 72 -1326 72 -1326 0 1
rlabel polysilicon 72 -1332 72 -1332 0 3
rlabel polysilicon 79 -1326 79 -1326 0 1
rlabel polysilicon 79 -1332 79 -1332 0 3
rlabel polysilicon 82 -1332 82 -1332 0 4
rlabel polysilicon 86 -1326 86 -1326 0 1
rlabel polysilicon 89 -1326 89 -1326 0 2
rlabel polysilicon 86 -1332 86 -1332 0 3
rlabel polysilicon 89 -1332 89 -1332 0 4
rlabel polysilicon 93 -1326 93 -1326 0 1
rlabel polysilicon 93 -1332 93 -1332 0 3
rlabel polysilicon 100 -1326 100 -1326 0 1
rlabel polysilicon 100 -1332 100 -1332 0 3
rlabel polysilicon 107 -1326 107 -1326 0 1
rlabel polysilicon 107 -1332 107 -1332 0 3
rlabel polysilicon 114 -1326 114 -1326 0 1
rlabel polysilicon 114 -1332 114 -1332 0 3
rlabel polysilicon 121 -1326 121 -1326 0 1
rlabel polysilicon 124 -1326 124 -1326 0 2
rlabel polysilicon 121 -1332 121 -1332 0 3
rlabel polysilicon 124 -1332 124 -1332 0 4
rlabel polysilicon 128 -1326 128 -1326 0 1
rlabel polysilicon 128 -1332 128 -1332 0 3
rlabel polysilicon 135 -1326 135 -1326 0 1
rlabel polysilicon 138 -1326 138 -1326 0 2
rlabel polysilicon 135 -1332 135 -1332 0 3
rlabel polysilicon 138 -1332 138 -1332 0 4
rlabel polysilicon 142 -1326 142 -1326 0 1
rlabel polysilicon 142 -1332 142 -1332 0 3
rlabel polysilicon 149 -1326 149 -1326 0 1
rlabel polysilicon 149 -1332 149 -1332 0 3
rlabel polysilicon 156 -1326 156 -1326 0 1
rlabel polysilicon 156 -1332 156 -1332 0 3
rlabel polysilicon 163 -1326 163 -1326 0 1
rlabel polysilicon 163 -1332 163 -1332 0 3
rlabel polysilicon 166 -1332 166 -1332 0 4
rlabel polysilicon 170 -1326 170 -1326 0 1
rlabel polysilicon 173 -1326 173 -1326 0 2
rlabel polysilicon 170 -1332 170 -1332 0 3
rlabel polysilicon 173 -1332 173 -1332 0 4
rlabel polysilicon 177 -1326 177 -1326 0 1
rlabel polysilicon 177 -1332 177 -1332 0 3
rlabel polysilicon 184 -1326 184 -1326 0 1
rlabel polysilicon 184 -1332 184 -1332 0 3
rlabel polysilicon 191 -1326 191 -1326 0 1
rlabel polysilicon 191 -1332 191 -1332 0 3
rlabel polysilicon 198 -1326 198 -1326 0 1
rlabel polysilicon 198 -1332 198 -1332 0 3
rlabel polysilicon 205 -1326 205 -1326 0 1
rlabel polysilicon 205 -1332 205 -1332 0 3
rlabel polysilicon 212 -1326 212 -1326 0 1
rlabel polysilicon 212 -1332 212 -1332 0 3
rlabel polysilicon 219 -1326 219 -1326 0 1
rlabel polysilicon 219 -1332 219 -1332 0 3
rlabel polysilicon 226 -1326 226 -1326 0 1
rlabel polysilicon 226 -1332 226 -1332 0 3
rlabel polysilicon 233 -1326 233 -1326 0 1
rlabel polysilicon 233 -1332 233 -1332 0 3
rlabel polysilicon 240 -1326 240 -1326 0 1
rlabel polysilicon 240 -1332 240 -1332 0 3
rlabel polysilicon 247 -1326 247 -1326 0 1
rlabel polysilicon 247 -1332 247 -1332 0 3
rlabel polysilicon 254 -1326 254 -1326 0 1
rlabel polysilicon 254 -1332 254 -1332 0 3
rlabel polysilicon 261 -1326 261 -1326 0 1
rlabel polysilicon 261 -1332 261 -1332 0 3
rlabel polysilicon 268 -1326 268 -1326 0 1
rlabel polysilicon 268 -1332 268 -1332 0 3
rlabel polysilicon 275 -1326 275 -1326 0 1
rlabel polysilicon 275 -1332 275 -1332 0 3
rlabel polysilicon 282 -1326 282 -1326 0 1
rlabel polysilicon 282 -1332 282 -1332 0 3
rlabel polysilicon 289 -1326 289 -1326 0 1
rlabel polysilicon 289 -1332 289 -1332 0 3
rlabel polysilicon 296 -1326 296 -1326 0 1
rlabel polysilicon 296 -1332 296 -1332 0 3
rlabel polysilicon 303 -1326 303 -1326 0 1
rlabel polysilicon 303 -1332 303 -1332 0 3
rlabel polysilicon 310 -1326 310 -1326 0 1
rlabel polysilicon 310 -1332 310 -1332 0 3
rlabel polysilicon 317 -1326 317 -1326 0 1
rlabel polysilicon 317 -1332 317 -1332 0 3
rlabel polysilicon 324 -1326 324 -1326 0 1
rlabel polysilicon 324 -1332 324 -1332 0 3
rlabel polysilicon 331 -1326 331 -1326 0 1
rlabel polysilicon 331 -1332 331 -1332 0 3
rlabel polysilicon 338 -1326 338 -1326 0 1
rlabel polysilicon 338 -1332 338 -1332 0 3
rlabel polysilicon 345 -1326 345 -1326 0 1
rlabel polysilicon 345 -1332 345 -1332 0 3
rlabel polysilicon 352 -1326 352 -1326 0 1
rlabel polysilicon 352 -1332 352 -1332 0 3
rlabel polysilicon 359 -1326 359 -1326 0 1
rlabel polysilicon 359 -1332 359 -1332 0 3
rlabel polysilicon 366 -1326 366 -1326 0 1
rlabel polysilicon 369 -1326 369 -1326 0 2
rlabel polysilicon 366 -1332 366 -1332 0 3
rlabel polysilicon 369 -1332 369 -1332 0 4
rlabel polysilicon 376 -1326 376 -1326 0 2
rlabel polysilicon 373 -1332 373 -1332 0 3
rlabel polysilicon 376 -1332 376 -1332 0 4
rlabel polysilicon 380 -1326 380 -1326 0 1
rlabel polysilicon 380 -1332 380 -1332 0 3
rlabel polysilicon 387 -1326 387 -1326 0 1
rlabel polysilicon 390 -1326 390 -1326 0 2
rlabel polysilicon 387 -1332 387 -1332 0 3
rlabel polysilicon 390 -1332 390 -1332 0 4
rlabel polysilicon 394 -1326 394 -1326 0 1
rlabel polysilicon 394 -1332 394 -1332 0 3
rlabel polysilicon 401 -1326 401 -1326 0 1
rlabel polysilicon 401 -1332 401 -1332 0 3
rlabel polysilicon 408 -1326 408 -1326 0 1
rlabel polysilicon 408 -1332 408 -1332 0 3
rlabel polysilicon 415 -1326 415 -1326 0 1
rlabel polysilicon 418 -1326 418 -1326 0 2
rlabel polysilicon 415 -1332 415 -1332 0 3
rlabel polysilicon 418 -1332 418 -1332 0 4
rlabel polysilicon 422 -1326 422 -1326 0 1
rlabel polysilicon 422 -1332 422 -1332 0 3
rlabel polysilicon 432 -1326 432 -1326 0 2
rlabel polysilicon 429 -1332 429 -1332 0 3
rlabel polysilicon 436 -1326 436 -1326 0 1
rlabel polysilicon 436 -1332 436 -1332 0 3
rlabel polysilicon 443 -1326 443 -1326 0 1
rlabel polysilicon 446 -1326 446 -1326 0 2
rlabel polysilicon 443 -1332 443 -1332 0 3
rlabel polysilicon 446 -1332 446 -1332 0 4
rlabel polysilicon 450 -1326 450 -1326 0 1
rlabel polysilicon 450 -1332 450 -1332 0 3
rlabel polysilicon 457 -1326 457 -1326 0 1
rlabel polysilicon 457 -1332 457 -1332 0 3
rlabel polysilicon 464 -1326 464 -1326 0 1
rlabel polysilicon 464 -1332 464 -1332 0 3
rlabel polysilicon 471 -1326 471 -1326 0 1
rlabel polysilicon 471 -1332 471 -1332 0 3
rlabel polysilicon 478 -1326 478 -1326 0 1
rlabel polysilicon 478 -1332 478 -1332 0 3
rlabel polysilicon 485 -1326 485 -1326 0 1
rlabel polysilicon 485 -1332 485 -1332 0 3
rlabel polysilicon 492 -1326 492 -1326 0 1
rlabel polysilicon 492 -1332 492 -1332 0 3
rlabel polysilicon 499 -1326 499 -1326 0 1
rlabel polysilicon 499 -1332 499 -1332 0 3
rlabel polysilicon 506 -1326 506 -1326 0 1
rlabel polysilicon 506 -1332 506 -1332 0 3
rlabel polysilicon 513 -1326 513 -1326 0 1
rlabel polysilicon 513 -1332 513 -1332 0 3
rlabel polysilicon 520 -1326 520 -1326 0 1
rlabel polysilicon 520 -1332 520 -1332 0 3
rlabel polysilicon 527 -1326 527 -1326 0 1
rlabel polysilicon 527 -1332 527 -1332 0 3
rlabel polysilicon 534 -1326 534 -1326 0 1
rlabel polysilicon 534 -1332 534 -1332 0 3
rlabel polysilicon 541 -1326 541 -1326 0 1
rlabel polysilicon 544 -1326 544 -1326 0 2
rlabel polysilicon 541 -1332 541 -1332 0 3
rlabel polysilicon 544 -1332 544 -1332 0 4
rlabel polysilicon 548 -1326 548 -1326 0 1
rlabel polysilicon 548 -1332 548 -1332 0 3
rlabel polysilicon 555 -1326 555 -1326 0 1
rlabel polysilicon 555 -1332 555 -1332 0 3
rlabel polysilicon 562 -1326 562 -1326 0 1
rlabel polysilicon 562 -1332 562 -1332 0 3
rlabel polysilicon 569 -1326 569 -1326 0 1
rlabel polysilicon 572 -1326 572 -1326 0 2
rlabel polysilicon 569 -1332 569 -1332 0 3
rlabel polysilicon 572 -1332 572 -1332 0 4
rlabel polysilicon 576 -1326 576 -1326 0 1
rlabel polysilicon 576 -1332 576 -1332 0 3
rlabel polysilicon 583 -1326 583 -1326 0 1
rlabel polysilicon 583 -1332 583 -1332 0 3
rlabel polysilicon 590 -1326 590 -1326 0 1
rlabel polysilicon 590 -1332 590 -1332 0 3
rlabel polysilicon 597 -1326 597 -1326 0 1
rlabel polysilicon 597 -1332 597 -1332 0 3
rlabel polysilicon 604 -1326 604 -1326 0 1
rlabel polysilicon 604 -1332 604 -1332 0 3
rlabel polysilicon 611 -1326 611 -1326 0 1
rlabel polysilicon 614 -1326 614 -1326 0 2
rlabel polysilicon 611 -1332 611 -1332 0 3
rlabel polysilicon 614 -1332 614 -1332 0 4
rlabel polysilicon 618 -1326 618 -1326 0 1
rlabel polysilicon 621 -1326 621 -1326 0 2
rlabel polysilicon 625 -1326 625 -1326 0 1
rlabel polysilicon 625 -1332 625 -1332 0 3
rlabel polysilicon 632 -1326 632 -1326 0 1
rlabel polysilicon 635 -1326 635 -1326 0 2
rlabel polysilicon 632 -1332 632 -1332 0 3
rlabel polysilicon 635 -1332 635 -1332 0 4
rlabel polysilicon 639 -1326 639 -1326 0 1
rlabel polysilicon 639 -1332 639 -1332 0 3
rlabel polysilicon 646 -1326 646 -1326 0 1
rlabel polysilicon 646 -1332 646 -1332 0 3
rlabel polysilicon 653 -1326 653 -1326 0 1
rlabel polysilicon 653 -1332 653 -1332 0 3
rlabel polysilicon 660 -1326 660 -1326 0 1
rlabel polysilicon 660 -1332 660 -1332 0 3
rlabel polysilicon 667 -1326 667 -1326 0 1
rlabel polysilicon 667 -1332 667 -1332 0 3
rlabel polysilicon 674 -1326 674 -1326 0 1
rlabel polysilicon 674 -1332 674 -1332 0 3
rlabel polysilicon 681 -1326 681 -1326 0 1
rlabel polysilicon 684 -1326 684 -1326 0 2
rlabel polysilicon 681 -1332 681 -1332 0 3
rlabel polysilicon 684 -1332 684 -1332 0 4
rlabel polysilicon 688 -1326 688 -1326 0 1
rlabel polysilicon 688 -1332 688 -1332 0 3
rlabel polysilicon 695 -1326 695 -1326 0 1
rlabel polysilicon 698 -1326 698 -1326 0 2
rlabel polysilicon 695 -1332 695 -1332 0 3
rlabel polysilicon 698 -1332 698 -1332 0 4
rlabel polysilicon 702 -1326 702 -1326 0 1
rlabel polysilicon 705 -1326 705 -1326 0 2
rlabel polysilicon 702 -1332 702 -1332 0 3
rlabel polysilicon 705 -1332 705 -1332 0 4
rlabel polysilicon 709 -1326 709 -1326 0 1
rlabel polysilicon 709 -1332 709 -1332 0 3
rlabel polysilicon 719 -1326 719 -1326 0 2
rlabel polysilicon 716 -1332 716 -1332 0 3
rlabel polysilicon 719 -1332 719 -1332 0 4
rlabel polysilicon 723 -1326 723 -1326 0 1
rlabel polysilicon 723 -1332 723 -1332 0 3
rlabel polysilicon 730 -1326 730 -1326 0 1
rlabel polysilicon 733 -1326 733 -1326 0 2
rlabel polysilicon 730 -1332 730 -1332 0 3
rlabel polysilicon 737 -1326 737 -1326 0 1
rlabel polysilicon 737 -1332 737 -1332 0 3
rlabel polysilicon 744 -1326 744 -1326 0 1
rlabel polysilicon 744 -1332 744 -1332 0 3
rlabel polysilicon 751 -1326 751 -1326 0 1
rlabel polysilicon 751 -1332 751 -1332 0 3
rlabel polysilicon 758 -1326 758 -1326 0 1
rlabel polysilicon 758 -1332 758 -1332 0 3
rlabel polysilicon 765 -1326 765 -1326 0 1
rlabel polysilicon 765 -1332 765 -1332 0 3
rlabel polysilicon 772 -1326 772 -1326 0 1
rlabel polysilicon 772 -1332 772 -1332 0 3
rlabel polysilicon 779 -1326 779 -1326 0 1
rlabel polysilicon 779 -1332 779 -1332 0 3
rlabel polysilicon 786 -1326 786 -1326 0 1
rlabel polysilicon 786 -1332 786 -1332 0 3
rlabel polysilicon 793 -1326 793 -1326 0 1
rlabel polysilicon 793 -1332 793 -1332 0 3
rlabel polysilicon 800 -1326 800 -1326 0 1
rlabel polysilicon 800 -1332 800 -1332 0 3
rlabel polysilicon 807 -1326 807 -1326 0 1
rlabel polysilicon 807 -1332 807 -1332 0 3
rlabel polysilicon 814 -1326 814 -1326 0 1
rlabel polysilicon 817 -1326 817 -1326 0 2
rlabel polysilicon 814 -1332 814 -1332 0 3
rlabel polysilicon 821 -1326 821 -1326 0 1
rlabel polysilicon 821 -1332 821 -1332 0 3
rlabel polysilicon 828 -1326 828 -1326 0 1
rlabel polysilicon 828 -1332 828 -1332 0 3
rlabel polysilicon 835 -1326 835 -1326 0 1
rlabel polysilicon 835 -1332 835 -1332 0 3
rlabel polysilicon 842 -1326 842 -1326 0 1
rlabel polysilicon 842 -1332 842 -1332 0 3
rlabel polysilicon 849 -1326 849 -1326 0 1
rlabel polysilicon 849 -1332 849 -1332 0 3
rlabel polysilicon 856 -1326 856 -1326 0 1
rlabel polysilicon 856 -1332 856 -1332 0 3
rlabel polysilicon 863 -1326 863 -1326 0 1
rlabel polysilicon 866 -1326 866 -1326 0 2
rlabel polysilicon 866 -1332 866 -1332 0 4
rlabel polysilicon 870 -1326 870 -1326 0 1
rlabel polysilicon 870 -1332 870 -1332 0 3
rlabel polysilicon 877 -1326 877 -1326 0 1
rlabel polysilicon 877 -1332 877 -1332 0 3
rlabel polysilicon 884 -1326 884 -1326 0 1
rlabel polysilicon 884 -1332 884 -1332 0 3
rlabel polysilicon 891 -1326 891 -1326 0 1
rlabel polysilicon 891 -1332 891 -1332 0 3
rlabel polysilicon 898 -1326 898 -1326 0 1
rlabel polysilicon 898 -1332 898 -1332 0 3
rlabel polysilicon 905 -1326 905 -1326 0 1
rlabel polysilicon 905 -1332 905 -1332 0 3
rlabel polysilicon 912 -1326 912 -1326 0 1
rlabel polysilicon 915 -1326 915 -1326 0 2
rlabel polysilicon 912 -1332 912 -1332 0 3
rlabel polysilicon 915 -1332 915 -1332 0 4
rlabel polysilicon 919 -1326 919 -1326 0 1
rlabel polysilicon 919 -1332 919 -1332 0 3
rlabel polysilicon 926 -1326 926 -1326 0 1
rlabel polysilicon 926 -1332 926 -1332 0 3
rlabel polysilicon 933 -1326 933 -1326 0 1
rlabel polysilicon 933 -1332 933 -1332 0 3
rlabel polysilicon 940 -1326 940 -1326 0 1
rlabel polysilicon 940 -1332 940 -1332 0 3
rlabel polysilicon 947 -1326 947 -1326 0 1
rlabel polysilicon 947 -1332 947 -1332 0 3
rlabel polysilicon 954 -1326 954 -1326 0 1
rlabel polysilicon 954 -1332 954 -1332 0 3
rlabel polysilicon 961 -1326 961 -1326 0 1
rlabel polysilicon 961 -1332 961 -1332 0 3
rlabel polysilicon 968 -1326 968 -1326 0 1
rlabel polysilicon 968 -1332 968 -1332 0 3
rlabel polysilicon 975 -1326 975 -1326 0 1
rlabel polysilicon 975 -1332 975 -1332 0 3
rlabel polysilicon 982 -1326 982 -1326 0 1
rlabel polysilicon 982 -1332 982 -1332 0 3
rlabel polysilicon 989 -1326 989 -1326 0 1
rlabel polysilicon 989 -1332 989 -1332 0 3
rlabel polysilicon 996 -1326 996 -1326 0 1
rlabel polysilicon 996 -1332 996 -1332 0 3
rlabel polysilicon 1003 -1326 1003 -1326 0 1
rlabel polysilicon 1003 -1332 1003 -1332 0 3
rlabel polysilicon 1010 -1326 1010 -1326 0 1
rlabel polysilicon 1010 -1332 1010 -1332 0 3
rlabel polysilicon 1017 -1326 1017 -1326 0 1
rlabel polysilicon 1017 -1332 1017 -1332 0 3
rlabel polysilicon 1024 -1326 1024 -1326 0 1
rlabel polysilicon 1024 -1332 1024 -1332 0 3
rlabel polysilicon 1031 -1326 1031 -1326 0 1
rlabel polysilicon 1031 -1332 1031 -1332 0 3
rlabel polysilicon 1038 -1326 1038 -1326 0 1
rlabel polysilicon 1038 -1332 1038 -1332 0 3
rlabel polysilicon 1045 -1326 1045 -1326 0 1
rlabel polysilicon 1045 -1332 1045 -1332 0 3
rlabel polysilicon 1052 -1326 1052 -1326 0 1
rlabel polysilicon 1052 -1332 1052 -1332 0 3
rlabel polysilicon 1059 -1326 1059 -1326 0 1
rlabel polysilicon 1059 -1332 1059 -1332 0 3
rlabel polysilicon 1066 -1326 1066 -1326 0 1
rlabel polysilicon 1066 -1332 1066 -1332 0 3
rlabel polysilicon 1073 -1326 1073 -1326 0 1
rlabel polysilicon 1073 -1332 1073 -1332 0 3
rlabel polysilicon 1080 -1326 1080 -1326 0 1
rlabel polysilicon 1080 -1332 1080 -1332 0 3
rlabel polysilicon 1087 -1326 1087 -1326 0 1
rlabel polysilicon 1087 -1332 1087 -1332 0 3
rlabel polysilicon 1094 -1326 1094 -1326 0 1
rlabel polysilicon 1094 -1332 1094 -1332 0 3
rlabel polysilicon 1101 -1326 1101 -1326 0 1
rlabel polysilicon 1101 -1332 1101 -1332 0 3
rlabel polysilicon 1108 -1326 1108 -1326 0 1
rlabel polysilicon 1108 -1332 1108 -1332 0 3
rlabel polysilicon 1115 -1332 1115 -1332 0 3
rlabel polysilicon 1122 -1326 1122 -1326 0 1
rlabel polysilicon 1122 -1332 1122 -1332 0 3
rlabel polysilicon 1129 -1326 1129 -1326 0 1
rlabel polysilicon 1129 -1332 1129 -1332 0 3
rlabel polysilicon 1136 -1326 1136 -1326 0 1
rlabel polysilicon 1136 -1332 1136 -1332 0 3
rlabel polysilicon 1143 -1326 1143 -1326 0 1
rlabel polysilicon 1143 -1332 1143 -1332 0 3
rlabel polysilicon 1150 -1326 1150 -1326 0 1
rlabel polysilicon 1150 -1332 1150 -1332 0 3
rlabel polysilicon 1157 -1326 1157 -1326 0 1
rlabel polysilicon 1157 -1332 1157 -1332 0 3
rlabel polysilicon 1164 -1326 1164 -1326 0 1
rlabel polysilicon 1164 -1332 1164 -1332 0 3
rlabel polysilicon 1171 -1326 1171 -1326 0 1
rlabel polysilicon 1171 -1332 1171 -1332 0 3
rlabel polysilicon 1178 -1326 1178 -1326 0 1
rlabel polysilicon 1178 -1332 1178 -1332 0 3
rlabel polysilicon 1185 -1326 1185 -1326 0 1
rlabel polysilicon 1185 -1332 1185 -1332 0 3
rlabel polysilicon 1192 -1326 1192 -1326 0 1
rlabel polysilicon 1192 -1332 1192 -1332 0 3
rlabel polysilicon 1199 -1326 1199 -1326 0 1
rlabel polysilicon 1199 -1332 1199 -1332 0 3
rlabel polysilicon 1206 -1326 1206 -1326 0 1
rlabel polysilicon 1206 -1332 1206 -1332 0 3
rlabel polysilicon 1213 -1326 1213 -1326 0 1
rlabel polysilicon 1213 -1332 1213 -1332 0 3
rlabel polysilicon 1220 -1326 1220 -1326 0 1
rlabel polysilicon 1220 -1332 1220 -1332 0 3
rlabel polysilicon 1227 -1326 1227 -1326 0 1
rlabel polysilicon 1227 -1332 1227 -1332 0 3
rlabel polysilicon 1234 -1326 1234 -1326 0 1
rlabel polysilicon 1234 -1332 1234 -1332 0 3
rlabel polysilicon 1241 -1326 1241 -1326 0 1
rlabel polysilicon 1241 -1332 1241 -1332 0 3
rlabel polysilicon 1248 -1326 1248 -1326 0 1
rlabel polysilicon 1248 -1332 1248 -1332 0 3
rlabel polysilicon 1255 -1326 1255 -1326 0 1
rlabel polysilicon 1255 -1332 1255 -1332 0 3
rlabel polysilicon 1262 -1326 1262 -1326 0 1
rlabel polysilicon 1262 -1332 1262 -1332 0 3
rlabel polysilicon 1269 -1326 1269 -1326 0 1
rlabel polysilicon 1272 -1326 1272 -1326 0 2
rlabel polysilicon 1269 -1332 1269 -1332 0 3
rlabel polysilicon 1276 -1326 1276 -1326 0 1
rlabel polysilicon 1276 -1332 1276 -1332 0 3
rlabel polysilicon 1283 -1326 1283 -1326 0 1
rlabel polysilicon 1283 -1332 1283 -1332 0 3
rlabel polysilicon 1290 -1326 1290 -1326 0 1
rlabel polysilicon 1290 -1332 1290 -1332 0 3
rlabel polysilicon 1297 -1326 1297 -1326 0 1
rlabel polysilicon 1297 -1332 1297 -1332 0 3
rlabel polysilicon 1304 -1326 1304 -1326 0 1
rlabel polysilicon 1304 -1332 1304 -1332 0 3
rlabel polysilicon 1311 -1326 1311 -1326 0 1
rlabel polysilicon 1311 -1332 1311 -1332 0 3
rlabel polysilicon 1318 -1326 1318 -1326 0 1
rlabel polysilicon 1318 -1332 1318 -1332 0 3
rlabel polysilicon 1325 -1326 1325 -1326 0 1
rlabel polysilicon 1325 -1332 1325 -1332 0 3
rlabel polysilicon 1332 -1326 1332 -1326 0 1
rlabel polysilicon 1332 -1332 1332 -1332 0 3
rlabel polysilicon 1339 -1326 1339 -1326 0 1
rlabel polysilicon 1339 -1332 1339 -1332 0 3
rlabel polysilicon 1346 -1326 1346 -1326 0 1
rlabel polysilicon 1346 -1332 1346 -1332 0 3
rlabel polysilicon 1353 -1326 1353 -1326 0 1
rlabel polysilicon 1353 -1332 1353 -1332 0 3
rlabel polysilicon 1360 -1326 1360 -1326 0 1
rlabel polysilicon 1360 -1332 1360 -1332 0 3
rlabel polysilicon 1367 -1326 1367 -1326 0 1
rlabel polysilicon 1367 -1332 1367 -1332 0 3
rlabel polysilicon 1374 -1326 1374 -1326 0 1
rlabel polysilicon 1374 -1332 1374 -1332 0 3
rlabel polysilicon 1381 -1326 1381 -1326 0 1
rlabel polysilicon 1381 -1332 1381 -1332 0 3
rlabel polysilicon 1388 -1326 1388 -1326 0 1
rlabel polysilicon 1388 -1332 1388 -1332 0 3
rlabel polysilicon 1458 -1326 1458 -1326 0 1
rlabel polysilicon 1458 -1332 1458 -1332 0 3
rlabel polysilicon 2 -1451 2 -1451 0 1
rlabel polysilicon 2 -1457 2 -1457 0 3
rlabel polysilicon 9 -1451 9 -1451 0 1
rlabel polysilicon 9 -1457 9 -1457 0 3
rlabel polysilicon 16 -1451 16 -1451 0 1
rlabel polysilicon 16 -1457 16 -1457 0 3
rlabel polysilicon 23 -1451 23 -1451 0 1
rlabel polysilicon 23 -1457 23 -1457 0 3
rlabel polysilicon 33 -1451 33 -1451 0 2
rlabel polysilicon 30 -1457 30 -1457 0 3
rlabel polysilicon 33 -1457 33 -1457 0 4
rlabel polysilicon 37 -1451 37 -1451 0 1
rlabel polysilicon 37 -1457 37 -1457 0 3
rlabel polysilicon 44 -1451 44 -1451 0 1
rlabel polysilicon 44 -1457 44 -1457 0 3
rlabel polysilicon 51 -1451 51 -1451 0 1
rlabel polysilicon 51 -1457 51 -1457 0 3
rlabel polysilicon 58 -1451 58 -1451 0 1
rlabel polysilicon 58 -1457 58 -1457 0 3
rlabel polysilicon 65 -1451 65 -1451 0 1
rlabel polysilicon 65 -1457 65 -1457 0 3
rlabel polysilicon 72 -1451 72 -1451 0 1
rlabel polysilicon 72 -1457 72 -1457 0 3
rlabel polysilicon 79 -1451 79 -1451 0 1
rlabel polysilicon 82 -1451 82 -1451 0 2
rlabel polysilicon 79 -1457 79 -1457 0 3
rlabel polysilicon 82 -1457 82 -1457 0 4
rlabel polysilicon 86 -1451 86 -1451 0 1
rlabel polysilicon 86 -1457 86 -1457 0 3
rlabel polysilicon 93 -1451 93 -1451 0 1
rlabel polysilicon 93 -1457 93 -1457 0 3
rlabel polysilicon 100 -1451 100 -1451 0 1
rlabel polysilicon 100 -1457 100 -1457 0 3
rlabel polysilicon 107 -1451 107 -1451 0 1
rlabel polysilicon 107 -1457 107 -1457 0 3
rlabel polysilicon 114 -1451 114 -1451 0 1
rlabel polysilicon 114 -1457 114 -1457 0 3
rlabel polysilicon 121 -1451 121 -1451 0 1
rlabel polysilicon 121 -1457 121 -1457 0 3
rlabel polysilicon 128 -1451 128 -1451 0 1
rlabel polysilicon 131 -1451 131 -1451 0 2
rlabel polysilicon 128 -1457 128 -1457 0 3
rlabel polysilicon 131 -1457 131 -1457 0 4
rlabel polysilicon 135 -1451 135 -1451 0 1
rlabel polysilicon 135 -1457 135 -1457 0 3
rlabel polysilicon 142 -1451 142 -1451 0 1
rlabel polysilicon 142 -1457 142 -1457 0 3
rlabel polysilicon 149 -1451 149 -1451 0 1
rlabel polysilicon 152 -1451 152 -1451 0 2
rlabel polysilicon 149 -1457 149 -1457 0 3
rlabel polysilicon 152 -1457 152 -1457 0 4
rlabel polysilicon 156 -1451 156 -1451 0 1
rlabel polysilicon 156 -1457 156 -1457 0 3
rlabel polysilicon 163 -1451 163 -1451 0 1
rlabel polysilicon 163 -1457 163 -1457 0 3
rlabel polysilicon 170 -1451 170 -1451 0 1
rlabel polysilicon 170 -1457 170 -1457 0 3
rlabel polysilicon 177 -1451 177 -1451 0 1
rlabel polysilicon 177 -1457 177 -1457 0 3
rlabel polysilicon 184 -1451 184 -1451 0 1
rlabel polysilicon 184 -1457 184 -1457 0 3
rlabel polysilicon 191 -1451 191 -1451 0 1
rlabel polysilicon 191 -1457 191 -1457 0 3
rlabel polysilicon 198 -1451 198 -1451 0 1
rlabel polysilicon 198 -1457 198 -1457 0 3
rlabel polysilicon 205 -1451 205 -1451 0 1
rlabel polysilicon 205 -1457 205 -1457 0 3
rlabel polysilicon 212 -1451 212 -1451 0 1
rlabel polysilicon 212 -1457 212 -1457 0 3
rlabel polysilicon 219 -1451 219 -1451 0 1
rlabel polysilicon 219 -1457 219 -1457 0 3
rlabel polysilicon 226 -1451 226 -1451 0 1
rlabel polysilicon 226 -1457 226 -1457 0 3
rlabel polysilicon 233 -1451 233 -1451 0 1
rlabel polysilicon 233 -1457 233 -1457 0 3
rlabel polysilicon 240 -1451 240 -1451 0 1
rlabel polysilicon 240 -1457 240 -1457 0 3
rlabel polysilicon 247 -1451 247 -1451 0 1
rlabel polysilicon 247 -1457 247 -1457 0 3
rlabel polysilicon 254 -1451 254 -1451 0 1
rlabel polysilicon 254 -1457 254 -1457 0 3
rlabel polysilicon 261 -1451 261 -1451 0 1
rlabel polysilicon 261 -1457 261 -1457 0 3
rlabel polysilicon 268 -1451 268 -1451 0 1
rlabel polysilicon 268 -1457 268 -1457 0 3
rlabel polysilicon 275 -1451 275 -1451 0 1
rlabel polysilicon 275 -1457 275 -1457 0 3
rlabel polysilicon 282 -1451 282 -1451 0 1
rlabel polysilicon 282 -1457 282 -1457 0 3
rlabel polysilicon 289 -1451 289 -1451 0 1
rlabel polysilicon 289 -1457 289 -1457 0 3
rlabel polysilicon 296 -1451 296 -1451 0 1
rlabel polysilicon 296 -1457 296 -1457 0 3
rlabel polysilicon 303 -1451 303 -1451 0 1
rlabel polysilicon 303 -1457 303 -1457 0 3
rlabel polysilicon 310 -1451 310 -1451 0 1
rlabel polysilicon 310 -1457 310 -1457 0 3
rlabel polysilicon 317 -1451 317 -1451 0 1
rlabel polysilicon 320 -1451 320 -1451 0 2
rlabel polysilicon 317 -1457 317 -1457 0 3
rlabel polysilicon 324 -1451 324 -1451 0 1
rlabel polysilicon 324 -1457 324 -1457 0 3
rlabel polysilicon 331 -1451 331 -1451 0 1
rlabel polysilicon 331 -1457 331 -1457 0 3
rlabel polysilicon 338 -1451 338 -1451 0 1
rlabel polysilicon 338 -1457 338 -1457 0 3
rlabel polysilicon 345 -1451 345 -1451 0 1
rlabel polysilicon 345 -1457 345 -1457 0 3
rlabel polysilicon 352 -1451 352 -1451 0 1
rlabel polysilicon 352 -1457 352 -1457 0 3
rlabel polysilicon 359 -1451 359 -1451 0 1
rlabel polysilicon 359 -1457 359 -1457 0 3
rlabel polysilicon 366 -1451 366 -1451 0 1
rlabel polysilicon 366 -1457 366 -1457 0 3
rlabel polysilicon 373 -1451 373 -1451 0 1
rlabel polysilicon 373 -1457 373 -1457 0 3
rlabel polysilicon 380 -1451 380 -1451 0 1
rlabel polysilicon 380 -1457 380 -1457 0 3
rlabel polysilicon 387 -1451 387 -1451 0 1
rlabel polysilicon 387 -1457 387 -1457 0 3
rlabel polysilicon 394 -1451 394 -1451 0 1
rlabel polysilicon 397 -1451 397 -1451 0 2
rlabel polysilicon 394 -1457 394 -1457 0 3
rlabel polysilicon 397 -1457 397 -1457 0 4
rlabel polysilicon 401 -1451 401 -1451 0 1
rlabel polysilicon 401 -1457 401 -1457 0 3
rlabel polysilicon 408 -1451 408 -1451 0 1
rlabel polysilicon 411 -1451 411 -1451 0 2
rlabel polysilicon 408 -1457 408 -1457 0 3
rlabel polysilicon 415 -1451 415 -1451 0 1
rlabel polysilicon 415 -1457 415 -1457 0 3
rlabel polysilicon 422 -1451 422 -1451 0 1
rlabel polysilicon 422 -1457 422 -1457 0 3
rlabel polysilicon 429 -1451 429 -1451 0 1
rlabel polysilicon 429 -1457 429 -1457 0 3
rlabel polysilicon 436 -1451 436 -1451 0 1
rlabel polysilicon 436 -1457 436 -1457 0 3
rlabel polysilicon 446 -1451 446 -1451 0 2
rlabel polysilicon 443 -1457 443 -1457 0 3
rlabel polysilicon 446 -1457 446 -1457 0 4
rlabel polysilicon 450 -1451 450 -1451 0 1
rlabel polysilicon 450 -1457 450 -1457 0 3
rlabel polysilicon 457 -1451 457 -1451 0 1
rlabel polysilicon 460 -1451 460 -1451 0 2
rlabel polysilicon 457 -1457 457 -1457 0 3
rlabel polysilicon 464 -1451 464 -1451 0 1
rlabel polysilicon 464 -1457 464 -1457 0 3
rlabel polysilicon 471 -1451 471 -1451 0 1
rlabel polysilicon 471 -1457 471 -1457 0 3
rlabel polysilicon 478 -1451 478 -1451 0 1
rlabel polysilicon 478 -1457 478 -1457 0 3
rlabel polysilicon 485 -1451 485 -1451 0 1
rlabel polysilicon 485 -1457 485 -1457 0 3
rlabel polysilicon 492 -1451 492 -1451 0 1
rlabel polysilicon 492 -1457 492 -1457 0 3
rlabel polysilicon 499 -1451 499 -1451 0 1
rlabel polysilicon 499 -1457 499 -1457 0 3
rlabel polysilicon 506 -1451 506 -1451 0 1
rlabel polysilicon 509 -1451 509 -1451 0 2
rlabel polysilicon 506 -1457 506 -1457 0 3
rlabel polysilicon 509 -1457 509 -1457 0 4
rlabel polysilicon 513 -1451 513 -1451 0 1
rlabel polysilicon 513 -1457 513 -1457 0 3
rlabel polysilicon 520 -1451 520 -1451 0 1
rlabel polysilicon 520 -1457 520 -1457 0 3
rlabel polysilicon 527 -1451 527 -1451 0 1
rlabel polysilicon 527 -1457 527 -1457 0 3
rlabel polysilicon 534 -1451 534 -1451 0 1
rlabel polysilicon 534 -1457 534 -1457 0 3
rlabel polysilicon 537 -1457 537 -1457 0 4
rlabel polysilicon 541 -1451 541 -1451 0 1
rlabel polysilicon 541 -1457 541 -1457 0 3
rlabel polysilicon 548 -1451 548 -1451 0 1
rlabel polysilicon 551 -1451 551 -1451 0 2
rlabel polysilicon 548 -1457 548 -1457 0 3
rlabel polysilicon 551 -1457 551 -1457 0 4
rlabel polysilicon 555 -1451 555 -1451 0 1
rlabel polysilicon 555 -1457 555 -1457 0 3
rlabel polysilicon 562 -1451 562 -1451 0 1
rlabel polysilicon 565 -1451 565 -1451 0 2
rlabel polysilicon 562 -1457 562 -1457 0 3
rlabel polysilicon 565 -1457 565 -1457 0 4
rlabel polysilicon 569 -1451 569 -1451 0 1
rlabel polysilicon 569 -1457 569 -1457 0 3
rlabel polysilicon 576 -1451 576 -1451 0 1
rlabel polysilicon 576 -1457 576 -1457 0 3
rlabel polysilicon 583 -1451 583 -1451 0 1
rlabel polysilicon 583 -1457 583 -1457 0 3
rlabel polysilicon 590 -1451 590 -1451 0 1
rlabel polysilicon 590 -1457 590 -1457 0 3
rlabel polysilicon 597 -1451 597 -1451 0 1
rlabel polysilicon 597 -1457 597 -1457 0 3
rlabel polysilicon 604 -1451 604 -1451 0 1
rlabel polysilicon 604 -1457 604 -1457 0 3
rlabel polysilicon 611 -1451 611 -1451 0 1
rlabel polysilicon 611 -1457 611 -1457 0 3
rlabel polysilicon 618 -1451 618 -1451 0 1
rlabel polysilicon 618 -1457 618 -1457 0 3
rlabel polysilicon 625 -1451 625 -1451 0 1
rlabel polysilicon 625 -1457 625 -1457 0 3
rlabel polysilicon 632 -1451 632 -1451 0 1
rlabel polysilicon 632 -1457 632 -1457 0 3
rlabel polysilicon 639 -1451 639 -1451 0 1
rlabel polysilicon 642 -1451 642 -1451 0 2
rlabel polysilicon 639 -1457 639 -1457 0 3
rlabel polysilicon 642 -1457 642 -1457 0 4
rlabel polysilicon 646 -1451 646 -1451 0 1
rlabel polysilicon 649 -1451 649 -1451 0 2
rlabel polysilicon 646 -1457 646 -1457 0 3
rlabel polysilicon 649 -1457 649 -1457 0 4
rlabel polysilicon 653 -1451 653 -1451 0 1
rlabel polysilicon 653 -1457 653 -1457 0 3
rlabel polysilicon 660 -1451 660 -1451 0 1
rlabel polysilicon 660 -1457 660 -1457 0 3
rlabel polysilicon 667 -1451 667 -1451 0 1
rlabel polysilicon 667 -1457 667 -1457 0 3
rlabel polysilicon 674 -1451 674 -1451 0 1
rlabel polysilicon 674 -1457 674 -1457 0 3
rlabel polysilicon 681 -1451 681 -1451 0 1
rlabel polysilicon 681 -1457 681 -1457 0 3
rlabel polysilicon 688 -1451 688 -1451 0 1
rlabel polysilicon 688 -1457 688 -1457 0 3
rlabel polysilicon 695 -1451 695 -1451 0 1
rlabel polysilicon 695 -1457 695 -1457 0 3
rlabel polysilicon 702 -1451 702 -1451 0 1
rlabel polysilicon 702 -1457 702 -1457 0 3
rlabel polysilicon 709 -1451 709 -1451 0 1
rlabel polysilicon 709 -1457 709 -1457 0 3
rlabel polysilicon 716 -1451 716 -1451 0 1
rlabel polysilicon 716 -1457 716 -1457 0 3
rlabel polysilicon 723 -1451 723 -1451 0 1
rlabel polysilicon 726 -1451 726 -1451 0 2
rlabel polysilicon 723 -1457 723 -1457 0 3
rlabel polysilicon 730 -1451 730 -1451 0 1
rlabel polysilicon 730 -1457 730 -1457 0 3
rlabel polysilicon 737 -1451 737 -1451 0 1
rlabel polysilicon 737 -1457 737 -1457 0 3
rlabel polysilicon 744 -1451 744 -1451 0 1
rlabel polysilicon 747 -1451 747 -1451 0 2
rlabel polysilicon 744 -1457 744 -1457 0 3
rlabel polysilicon 747 -1457 747 -1457 0 4
rlabel polysilicon 751 -1451 751 -1451 0 1
rlabel polysilicon 751 -1457 751 -1457 0 3
rlabel polysilicon 758 -1451 758 -1451 0 1
rlabel polysilicon 758 -1457 758 -1457 0 3
rlabel polysilicon 765 -1451 765 -1451 0 1
rlabel polysilicon 765 -1457 765 -1457 0 3
rlabel polysilicon 772 -1451 772 -1451 0 1
rlabel polysilicon 772 -1457 772 -1457 0 3
rlabel polysilicon 779 -1451 779 -1451 0 1
rlabel polysilicon 782 -1451 782 -1451 0 2
rlabel polysilicon 779 -1457 779 -1457 0 3
rlabel polysilicon 782 -1457 782 -1457 0 4
rlabel polysilicon 786 -1451 786 -1451 0 1
rlabel polysilicon 786 -1457 786 -1457 0 3
rlabel polysilicon 793 -1451 793 -1451 0 1
rlabel polysilicon 796 -1451 796 -1451 0 2
rlabel polysilicon 793 -1457 793 -1457 0 3
rlabel polysilicon 796 -1457 796 -1457 0 4
rlabel polysilicon 800 -1451 800 -1451 0 1
rlabel polysilicon 800 -1457 800 -1457 0 3
rlabel polysilicon 807 -1451 807 -1451 0 1
rlabel polysilicon 807 -1457 807 -1457 0 3
rlabel polysilicon 814 -1451 814 -1451 0 1
rlabel polysilicon 817 -1451 817 -1451 0 2
rlabel polysilicon 814 -1457 814 -1457 0 3
rlabel polysilicon 817 -1457 817 -1457 0 4
rlabel polysilicon 821 -1451 821 -1451 0 1
rlabel polysilicon 824 -1451 824 -1451 0 2
rlabel polysilicon 824 -1457 824 -1457 0 4
rlabel polysilicon 828 -1451 828 -1451 0 1
rlabel polysilicon 831 -1451 831 -1451 0 2
rlabel polysilicon 831 -1457 831 -1457 0 4
rlabel polysilicon 835 -1451 835 -1451 0 1
rlabel polysilicon 835 -1457 835 -1457 0 3
rlabel polysilicon 842 -1451 842 -1451 0 1
rlabel polysilicon 842 -1457 842 -1457 0 3
rlabel polysilicon 849 -1451 849 -1451 0 1
rlabel polysilicon 852 -1451 852 -1451 0 2
rlabel polysilicon 849 -1457 849 -1457 0 3
rlabel polysilicon 852 -1457 852 -1457 0 4
rlabel polysilicon 856 -1451 856 -1451 0 1
rlabel polysilicon 859 -1451 859 -1451 0 2
rlabel polysilicon 856 -1457 856 -1457 0 3
rlabel polysilicon 859 -1457 859 -1457 0 4
rlabel polysilicon 866 -1451 866 -1451 0 2
rlabel polysilicon 863 -1457 863 -1457 0 3
rlabel polysilicon 866 -1457 866 -1457 0 4
rlabel polysilicon 870 -1451 870 -1451 0 1
rlabel polysilicon 870 -1457 870 -1457 0 3
rlabel polysilicon 877 -1451 877 -1451 0 1
rlabel polysilicon 877 -1457 877 -1457 0 3
rlabel polysilicon 887 -1451 887 -1451 0 2
rlabel polysilicon 887 -1457 887 -1457 0 4
rlabel polysilicon 891 -1451 891 -1451 0 1
rlabel polysilicon 891 -1457 891 -1457 0 3
rlabel polysilicon 898 -1451 898 -1451 0 1
rlabel polysilicon 898 -1457 898 -1457 0 3
rlabel polysilicon 905 -1451 905 -1451 0 1
rlabel polysilicon 905 -1457 905 -1457 0 3
rlabel polysilicon 912 -1451 912 -1451 0 1
rlabel polysilicon 912 -1457 912 -1457 0 3
rlabel polysilicon 919 -1451 919 -1451 0 1
rlabel polysilicon 919 -1457 919 -1457 0 3
rlabel polysilicon 926 -1451 926 -1451 0 1
rlabel polysilicon 926 -1457 926 -1457 0 3
rlabel polysilicon 933 -1451 933 -1451 0 1
rlabel polysilicon 933 -1457 933 -1457 0 3
rlabel polysilicon 940 -1451 940 -1451 0 1
rlabel polysilicon 940 -1457 940 -1457 0 3
rlabel polysilicon 947 -1451 947 -1451 0 1
rlabel polysilicon 947 -1457 947 -1457 0 3
rlabel polysilicon 954 -1451 954 -1451 0 1
rlabel polysilicon 954 -1457 954 -1457 0 3
rlabel polysilicon 961 -1451 961 -1451 0 1
rlabel polysilicon 961 -1457 961 -1457 0 3
rlabel polysilicon 968 -1451 968 -1451 0 1
rlabel polysilicon 968 -1457 968 -1457 0 3
rlabel polysilicon 975 -1451 975 -1451 0 1
rlabel polysilicon 975 -1457 975 -1457 0 3
rlabel polysilicon 982 -1451 982 -1451 0 1
rlabel polysilicon 982 -1457 982 -1457 0 3
rlabel polysilicon 989 -1451 989 -1451 0 1
rlabel polysilicon 989 -1457 989 -1457 0 3
rlabel polysilicon 996 -1451 996 -1451 0 1
rlabel polysilicon 996 -1457 996 -1457 0 3
rlabel polysilicon 1003 -1451 1003 -1451 0 1
rlabel polysilicon 1003 -1457 1003 -1457 0 3
rlabel polysilicon 1010 -1451 1010 -1451 0 1
rlabel polysilicon 1010 -1457 1010 -1457 0 3
rlabel polysilicon 1017 -1451 1017 -1451 0 1
rlabel polysilicon 1017 -1457 1017 -1457 0 3
rlabel polysilicon 1024 -1451 1024 -1451 0 1
rlabel polysilicon 1024 -1457 1024 -1457 0 3
rlabel polysilicon 1031 -1451 1031 -1451 0 1
rlabel polysilicon 1031 -1457 1031 -1457 0 3
rlabel polysilicon 1038 -1451 1038 -1451 0 1
rlabel polysilicon 1038 -1457 1038 -1457 0 3
rlabel polysilicon 1045 -1451 1045 -1451 0 1
rlabel polysilicon 1045 -1457 1045 -1457 0 3
rlabel polysilicon 1052 -1451 1052 -1451 0 1
rlabel polysilicon 1052 -1457 1052 -1457 0 3
rlabel polysilicon 1059 -1451 1059 -1451 0 1
rlabel polysilicon 1059 -1457 1059 -1457 0 3
rlabel polysilicon 1066 -1451 1066 -1451 0 1
rlabel polysilicon 1066 -1457 1066 -1457 0 3
rlabel polysilicon 1073 -1451 1073 -1451 0 1
rlabel polysilicon 1073 -1457 1073 -1457 0 3
rlabel polysilicon 1080 -1451 1080 -1451 0 1
rlabel polysilicon 1080 -1457 1080 -1457 0 3
rlabel polysilicon 1087 -1451 1087 -1451 0 1
rlabel polysilicon 1087 -1457 1087 -1457 0 3
rlabel polysilicon 1094 -1451 1094 -1451 0 1
rlabel polysilicon 1094 -1457 1094 -1457 0 3
rlabel polysilicon 1101 -1451 1101 -1451 0 1
rlabel polysilicon 1101 -1457 1101 -1457 0 3
rlabel polysilicon 1108 -1451 1108 -1451 0 1
rlabel polysilicon 1108 -1457 1108 -1457 0 3
rlabel polysilicon 1115 -1451 1115 -1451 0 1
rlabel polysilicon 1115 -1457 1115 -1457 0 3
rlabel polysilicon 1122 -1451 1122 -1451 0 1
rlabel polysilicon 1122 -1457 1122 -1457 0 3
rlabel polysilicon 1129 -1451 1129 -1451 0 1
rlabel polysilicon 1129 -1457 1129 -1457 0 3
rlabel polysilicon 1136 -1451 1136 -1451 0 1
rlabel polysilicon 1136 -1457 1136 -1457 0 3
rlabel polysilicon 1143 -1451 1143 -1451 0 1
rlabel polysilicon 1143 -1457 1143 -1457 0 3
rlabel polysilicon 1150 -1451 1150 -1451 0 1
rlabel polysilicon 1150 -1457 1150 -1457 0 3
rlabel polysilicon 1157 -1451 1157 -1451 0 1
rlabel polysilicon 1157 -1457 1157 -1457 0 3
rlabel polysilicon 1164 -1451 1164 -1451 0 1
rlabel polysilicon 1164 -1457 1164 -1457 0 3
rlabel polysilicon 1171 -1451 1171 -1451 0 1
rlabel polysilicon 1171 -1457 1171 -1457 0 3
rlabel polysilicon 1178 -1451 1178 -1451 0 1
rlabel polysilicon 1178 -1457 1178 -1457 0 3
rlabel polysilicon 1185 -1451 1185 -1451 0 1
rlabel polysilicon 1185 -1457 1185 -1457 0 3
rlabel polysilicon 1192 -1451 1192 -1451 0 1
rlabel polysilicon 1192 -1457 1192 -1457 0 3
rlabel polysilicon 1199 -1451 1199 -1451 0 1
rlabel polysilicon 1199 -1457 1199 -1457 0 3
rlabel polysilicon 1206 -1451 1206 -1451 0 1
rlabel polysilicon 1206 -1457 1206 -1457 0 3
rlabel polysilicon 1213 -1451 1213 -1451 0 1
rlabel polysilicon 1213 -1457 1213 -1457 0 3
rlabel polysilicon 1220 -1451 1220 -1451 0 1
rlabel polysilicon 1220 -1457 1220 -1457 0 3
rlabel polysilicon 1227 -1451 1227 -1451 0 1
rlabel polysilicon 1227 -1457 1227 -1457 0 3
rlabel polysilicon 1234 -1451 1234 -1451 0 1
rlabel polysilicon 1234 -1457 1234 -1457 0 3
rlabel polysilicon 1241 -1451 1241 -1451 0 1
rlabel polysilicon 1241 -1457 1241 -1457 0 3
rlabel polysilicon 1248 -1451 1248 -1451 0 1
rlabel polysilicon 1248 -1457 1248 -1457 0 3
rlabel polysilicon 1255 -1451 1255 -1451 0 1
rlabel polysilicon 1255 -1457 1255 -1457 0 3
rlabel polysilicon 1262 -1451 1262 -1451 0 1
rlabel polysilicon 1262 -1457 1262 -1457 0 3
rlabel polysilicon 1269 -1451 1269 -1451 0 1
rlabel polysilicon 1269 -1457 1269 -1457 0 3
rlabel polysilicon 1276 -1451 1276 -1451 0 1
rlabel polysilicon 1276 -1457 1276 -1457 0 3
rlabel polysilicon 1283 -1451 1283 -1451 0 1
rlabel polysilicon 1283 -1457 1283 -1457 0 3
rlabel polysilicon 1290 -1451 1290 -1451 0 1
rlabel polysilicon 1290 -1457 1290 -1457 0 3
rlabel polysilicon 1297 -1451 1297 -1451 0 1
rlabel polysilicon 1297 -1457 1297 -1457 0 3
rlabel polysilicon 1304 -1451 1304 -1451 0 1
rlabel polysilicon 1304 -1457 1304 -1457 0 3
rlabel polysilicon 1311 -1451 1311 -1451 0 1
rlabel polysilicon 1311 -1457 1311 -1457 0 3
rlabel polysilicon 1318 -1451 1318 -1451 0 1
rlabel polysilicon 1318 -1457 1318 -1457 0 3
rlabel polysilicon 1325 -1451 1325 -1451 0 1
rlabel polysilicon 1325 -1457 1325 -1457 0 3
rlabel polysilicon 1332 -1451 1332 -1451 0 1
rlabel polysilicon 1332 -1457 1332 -1457 0 3
rlabel polysilicon 1339 -1451 1339 -1451 0 1
rlabel polysilicon 1339 -1457 1339 -1457 0 3
rlabel polysilicon 1346 -1451 1346 -1451 0 1
rlabel polysilicon 1346 -1457 1346 -1457 0 3
rlabel polysilicon 1353 -1451 1353 -1451 0 1
rlabel polysilicon 1353 -1457 1353 -1457 0 3
rlabel polysilicon 1360 -1451 1360 -1451 0 1
rlabel polysilicon 1360 -1457 1360 -1457 0 3
rlabel polysilicon 1367 -1451 1367 -1451 0 1
rlabel polysilicon 1367 -1457 1367 -1457 0 3
rlabel polysilicon 1374 -1451 1374 -1451 0 1
rlabel polysilicon 1374 -1457 1374 -1457 0 3
rlabel polysilicon 1381 -1451 1381 -1451 0 1
rlabel polysilicon 1381 -1457 1381 -1457 0 3
rlabel polysilicon 1388 -1451 1388 -1451 0 1
rlabel polysilicon 1388 -1457 1388 -1457 0 3
rlabel polysilicon 1395 -1451 1395 -1451 0 1
rlabel polysilicon 1395 -1457 1395 -1457 0 3
rlabel polysilicon 1402 -1451 1402 -1451 0 1
rlabel polysilicon 1402 -1457 1402 -1457 0 3
rlabel polysilicon 1409 -1451 1409 -1451 0 1
rlabel polysilicon 1409 -1457 1409 -1457 0 3
rlabel polysilicon 1416 -1451 1416 -1451 0 1
rlabel polysilicon 1416 -1457 1416 -1457 0 3
rlabel polysilicon 1423 -1451 1423 -1451 0 1
rlabel polysilicon 1423 -1457 1423 -1457 0 3
rlabel polysilicon 1430 -1451 1430 -1451 0 1
rlabel polysilicon 1430 -1457 1430 -1457 0 3
rlabel polysilicon 1437 -1451 1437 -1451 0 1
rlabel polysilicon 1437 -1457 1437 -1457 0 3
rlabel polysilicon 1444 -1451 1444 -1451 0 1
rlabel polysilicon 1444 -1457 1444 -1457 0 3
rlabel polysilicon 1451 -1451 1451 -1451 0 1
rlabel polysilicon 1451 -1457 1451 -1457 0 3
rlabel polysilicon 1454 -1457 1454 -1457 0 4
rlabel polysilicon 1458 -1451 1458 -1451 0 1
rlabel polysilicon 1458 -1457 1458 -1457 0 3
rlabel polysilicon 1465 -1451 1465 -1451 0 1
rlabel polysilicon 1465 -1457 1465 -1457 0 3
rlabel polysilicon 2 -1588 2 -1588 0 1
rlabel polysilicon 2 -1594 2 -1594 0 3
rlabel polysilicon 9 -1588 9 -1588 0 1
rlabel polysilicon 12 -1588 12 -1588 0 2
rlabel polysilicon 12 -1594 12 -1594 0 4
rlabel polysilicon 16 -1588 16 -1588 0 1
rlabel polysilicon 19 -1588 19 -1588 0 2
rlabel polysilicon 16 -1594 16 -1594 0 3
rlabel polysilicon 23 -1588 23 -1588 0 1
rlabel polysilicon 23 -1594 23 -1594 0 3
rlabel polysilicon 30 -1588 30 -1588 0 1
rlabel polysilicon 30 -1594 30 -1594 0 3
rlabel polysilicon 37 -1588 37 -1588 0 1
rlabel polysilicon 40 -1588 40 -1588 0 2
rlabel polysilicon 37 -1594 37 -1594 0 3
rlabel polysilicon 40 -1594 40 -1594 0 4
rlabel polysilicon 44 -1588 44 -1588 0 1
rlabel polysilicon 44 -1594 44 -1594 0 3
rlabel polysilicon 51 -1588 51 -1588 0 1
rlabel polysilicon 54 -1588 54 -1588 0 2
rlabel polysilicon 51 -1594 51 -1594 0 3
rlabel polysilicon 54 -1594 54 -1594 0 4
rlabel polysilicon 58 -1588 58 -1588 0 1
rlabel polysilicon 58 -1594 58 -1594 0 3
rlabel polysilicon 65 -1588 65 -1588 0 1
rlabel polysilicon 65 -1594 65 -1594 0 3
rlabel polysilicon 72 -1588 72 -1588 0 1
rlabel polysilicon 72 -1594 72 -1594 0 3
rlabel polysilicon 79 -1588 79 -1588 0 1
rlabel polysilicon 79 -1594 79 -1594 0 3
rlabel polysilicon 86 -1588 86 -1588 0 1
rlabel polysilicon 89 -1588 89 -1588 0 2
rlabel polysilicon 86 -1594 86 -1594 0 3
rlabel polysilicon 89 -1594 89 -1594 0 4
rlabel polysilicon 93 -1588 93 -1588 0 1
rlabel polysilicon 93 -1594 93 -1594 0 3
rlabel polysilicon 100 -1588 100 -1588 0 1
rlabel polysilicon 103 -1588 103 -1588 0 2
rlabel polysilicon 100 -1594 100 -1594 0 3
rlabel polysilicon 103 -1594 103 -1594 0 4
rlabel polysilicon 107 -1588 107 -1588 0 1
rlabel polysilicon 107 -1594 107 -1594 0 3
rlabel polysilicon 114 -1588 114 -1588 0 1
rlabel polysilicon 117 -1588 117 -1588 0 2
rlabel polysilicon 114 -1594 114 -1594 0 3
rlabel polysilicon 117 -1594 117 -1594 0 4
rlabel polysilicon 121 -1588 121 -1588 0 1
rlabel polysilicon 121 -1594 121 -1594 0 3
rlabel polysilicon 128 -1588 128 -1588 0 1
rlabel polysilicon 128 -1594 128 -1594 0 3
rlabel polysilicon 135 -1588 135 -1588 0 1
rlabel polysilicon 138 -1588 138 -1588 0 2
rlabel polysilicon 135 -1594 135 -1594 0 3
rlabel polysilicon 138 -1594 138 -1594 0 4
rlabel polysilicon 142 -1588 142 -1588 0 1
rlabel polysilicon 145 -1588 145 -1588 0 2
rlabel polysilicon 142 -1594 142 -1594 0 3
rlabel polysilicon 145 -1594 145 -1594 0 4
rlabel polysilicon 149 -1588 149 -1588 0 1
rlabel polysilicon 149 -1594 149 -1594 0 3
rlabel polysilicon 156 -1588 156 -1588 0 1
rlabel polysilicon 156 -1594 156 -1594 0 3
rlabel polysilicon 163 -1588 163 -1588 0 1
rlabel polysilicon 163 -1594 163 -1594 0 3
rlabel polysilicon 170 -1588 170 -1588 0 1
rlabel polysilicon 170 -1594 170 -1594 0 3
rlabel polysilicon 180 -1588 180 -1588 0 2
rlabel polysilicon 177 -1594 177 -1594 0 3
rlabel polysilicon 180 -1594 180 -1594 0 4
rlabel polysilicon 184 -1588 184 -1588 0 1
rlabel polysilicon 184 -1594 184 -1594 0 3
rlabel polysilicon 191 -1588 191 -1588 0 1
rlabel polysilicon 191 -1594 191 -1594 0 3
rlabel polysilicon 198 -1588 198 -1588 0 1
rlabel polysilicon 198 -1594 198 -1594 0 3
rlabel polysilicon 205 -1588 205 -1588 0 1
rlabel polysilicon 205 -1594 205 -1594 0 3
rlabel polysilicon 212 -1588 212 -1588 0 1
rlabel polysilicon 212 -1594 212 -1594 0 3
rlabel polysilicon 219 -1588 219 -1588 0 1
rlabel polysilicon 219 -1594 219 -1594 0 3
rlabel polysilicon 226 -1588 226 -1588 0 1
rlabel polysilicon 226 -1594 226 -1594 0 3
rlabel polysilicon 233 -1588 233 -1588 0 1
rlabel polysilicon 233 -1594 233 -1594 0 3
rlabel polysilicon 240 -1588 240 -1588 0 1
rlabel polysilicon 240 -1594 240 -1594 0 3
rlabel polysilicon 247 -1588 247 -1588 0 1
rlabel polysilicon 247 -1594 247 -1594 0 3
rlabel polysilicon 254 -1588 254 -1588 0 1
rlabel polysilicon 254 -1594 254 -1594 0 3
rlabel polysilicon 261 -1588 261 -1588 0 1
rlabel polysilicon 261 -1594 261 -1594 0 3
rlabel polysilicon 268 -1588 268 -1588 0 1
rlabel polysilicon 268 -1594 268 -1594 0 3
rlabel polysilicon 275 -1588 275 -1588 0 1
rlabel polysilicon 275 -1594 275 -1594 0 3
rlabel polysilicon 282 -1588 282 -1588 0 1
rlabel polysilicon 282 -1594 282 -1594 0 3
rlabel polysilicon 289 -1588 289 -1588 0 1
rlabel polysilicon 289 -1594 289 -1594 0 3
rlabel polysilicon 296 -1588 296 -1588 0 1
rlabel polysilicon 296 -1594 296 -1594 0 3
rlabel polysilicon 303 -1588 303 -1588 0 1
rlabel polysilicon 303 -1594 303 -1594 0 3
rlabel polysilicon 310 -1588 310 -1588 0 1
rlabel polysilicon 310 -1594 310 -1594 0 3
rlabel polysilicon 317 -1588 317 -1588 0 1
rlabel polysilicon 317 -1594 317 -1594 0 3
rlabel polysilicon 324 -1588 324 -1588 0 1
rlabel polysilicon 324 -1594 324 -1594 0 3
rlabel polysilicon 331 -1588 331 -1588 0 1
rlabel polysilicon 331 -1594 331 -1594 0 3
rlabel polysilicon 338 -1588 338 -1588 0 1
rlabel polysilicon 338 -1594 338 -1594 0 3
rlabel polysilicon 345 -1588 345 -1588 0 1
rlabel polysilicon 345 -1594 345 -1594 0 3
rlabel polysilicon 352 -1588 352 -1588 0 1
rlabel polysilicon 352 -1594 352 -1594 0 3
rlabel polysilicon 359 -1588 359 -1588 0 1
rlabel polysilicon 359 -1594 359 -1594 0 3
rlabel polysilicon 366 -1588 366 -1588 0 1
rlabel polysilicon 366 -1594 366 -1594 0 3
rlabel polysilicon 373 -1588 373 -1588 0 1
rlabel polysilicon 373 -1594 373 -1594 0 3
rlabel polysilicon 380 -1588 380 -1588 0 1
rlabel polysilicon 380 -1594 380 -1594 0 3
rlabel polysilicon 387 -1588 387 -1588 0 1
rlabel polysilicon 387 -1594 387 -1594 0 3
rlabel polysilicon 394 -1588 394 -1588 0 1
rlabel polysilicon 394 -1594 394 -1594 0 3
rlabel polysilicon 401 -1588 401 -1588 0 1
rlabel polysilicon 404 -1588 404 -1588 0 2
rlabel polysilicon 404 -1594 404 -1594 0 4
rlabel polysilicon 408 -1588 408 -1588 0 1
rlabel polysilicon 408 -1594 408 -1594 0 3
rlabel polysilicon 415 -1588 415 -1588 0 1
rlabel polysilicon 415 -1594 415 -1594 0 3
rlabel polysilicon 422 -1588 422 -1588 0 1
rlabel polysilicon 422 -1594 422 -1594 0 3
rlabel polysilicon 429 -1588 429 -1588 0 1
rlabel polysilicon 432 -1588 432 -1588 0 2
rlabel polysilicon 429 -1594 429 -1594 0 3
rlabel polysilicon 432 -1594 432 -1594 0 4
rlabel polysilicon 436 -1588 436 -1588 0 1
rlabel polysilicon 436 -1594 436 -1594 0 3
rlabel polysilicon 443 -1588 443 -1588 0 1
rlabel polysilicon 443 -1594 443 -1594 0 3
rlabel polysilicon 450 -1588 450 -1588 0 1
rlabel polysilicon 450 -1594 450 -1594 0 3
rlabel polysilicon 457 -1588 457 -1588 0 1
rlabel polysilicon 460 -1588 460 -1588 0 2
rlabel polysilicon 457 -1594 457 -1594 0 3
rlabel polysilicon 460 -1594 460 -1594 0 4
rlabel polysilicon 464 -1588 464 -1588 0 1
rlabel polysilicon 464 -1594 464 -1594 0 3
rlabel polysilicon 471 -1588 471 -1588 0 1
rlabel polysilicon 471 -1594 471 -1594 0 3
rlabel polysilicon 478 -1588 478 -1588 0 1
rlabel polysilicon 478 -1594 478 -1594 0 3
rlabel polysilicon 485 -1588 485 -1588 0 1
rlabel polysilicon 488 -1588 488 -1588 0 2
rlabel polysilicon 485 -1594 485 -1594 0 3
rlabel polysilicon 492 -1588 492 -1588 0 1
rlabel polysilicon 492 -1594 492 -1594 0 3
rlabel polysilicon 495 -1594 495 -1594 0 4
rlabel polysilicon 499 -1588 499 -1588 0 1
rlabel polysilicon 499 -1594 499 -1594 0 3
rlabel polysilicon 506 -1588 506 -1588 0 1
rlabel polysilicon 506 -1594 506 -1594 0 3
rlabel polysilicon 513 -1588 513 -1588 0 1
rlabel polysilicon 513 -1594 513 -1594 0 3
rlabel polysilicon 520 -1588 520 -1588 0 1
rlabel polysilicon 523 -1588 523 -1588 0 2
rlabel polysilicon 520 -1594 520 -1594 0 3
rlabel polysilicon 523 -1594 523 -1594 0 4
rlabel polysilicon 527 -1588 527 -1588 0 1
rlabel polysilicon 527 -1594 527 -1594 0 3
rlabel polysilicon 534 -1588 534 -1588 0 1
rlabel polysilicon 537 -1588 537 -1588 0 2
rlabel polysilicon 534 -1594 534 -1594 0 3
rlabel polysilicon 537 -1594 537 -1594 0 4
rlabel polysilicon 541 -1588 541 -1588 0 1
rlabel polysilicon 541 -1594 541 -1594 0 3
rlabel polysilicon 548 -1588 548 -1588 0 1
rlabel polysilicon 548 -1594 548 -1594 0 3
rlabel polysilicon 555 -1588 555 -1588 0 1
rlabel polysilicon 558 -1588 558 -1588 0 2
rlabel polysilicon 555 -1594 555 -1594 0 3
rlabel polysilicon 558 -1594 558 -1594 0 4
rlabel polysilicon 562 -1588 562 -1588 0 1
rlabel polysilicon 562 -1594 562 -1594 0 3
rlabel polysilicon 569 -1588 569 -1588 0 1
rlabel polysilicon 572 -1588 572 -1588 0 2
rlabel polysilicon 569 -1594 569 -1594 0 3
rlabel polysilicon 572 -1594 572 -1594 0 4
rlabel polysilicon 576 -1588 576 -1588 0 1
rlabel polysilicon 576 -1594 576 -1594 0 3
rlabel polysilicon 583 -1588 583 -1588 0 1
rlabel polysilicon 583 -1594 583 -1594 0 3
rlabel polysilicon 590 -1588 590 -1588 0 1
rlabel polysilicon 590 -1594 590 -1594 0 3
rlabel polysilicon 597 -1588 597 -1588 0 1
rlabel polysilicon 597 -1594 597 -1594 0 3
rlabel polysilicon 604 -1588 604 -1588 0 1
rlabel polysilicon 604 -1594 604 -1594 0 3
rlabel polysilicon 611 -1588 611 -1588 0 1
rlabel polysilicon 611 -1594 611 -1594 0 3
rlabel polysilicon 618 -1588 618 -1588 0 1
rlabel polysilicon 621 -1588 621 -1588 0 2
rlabel polysilicon 618 -1594 618 -1594 0 3
rlabel polysilicon 621 -1594 621 -1594 0 4
rlabel polysilicon 625 -1588 625 -1588 0 1
rlabel polysilicon 625 -1594 625 -1594 0 3
rlabel polysilicon 632 -1588 632 -1588 0 1
rlabel polysilicon 632 -1594 632 -1594 0 3
rlabel polysilicon 639 -1588 639 -1588 0 1
rlabel polysilicon 639 -1594 639 -1594 0 3
rlabel polysilicon 646 -1588 646 -1588 0 1
rlabel polysilicon 646 -1594 646 -1594 0 3
rlabel polysilicon 653 -1588 653 -1588 0 1
rlabel polysilicon 653 -1594 653 -1594 0 3
rlabel polysilicon 663 -1588 663 -1588 0 2
rlabel polysilicon 660 -1594 660 -1594 0 3
rlabel polysilicon 663 -1594 663 -1594 0 4
rlabel polysilicon 667 -1588 667 -1588 0 1
rlabel polysilicon 667 -1594 667 -1594 0 3
rlabel polysilicon 674 -1588 674 -1588 0 1
rlabel polysilicon 674 -1594 674 -1594 0 3
rlabel polysilicon 681 -1588 681 -1588 0 1
rlabel polysilicon 681 -1594 681 -1594 0 3
rlabel polysilicon 688 -1588 688 -1588 0 1
rlabel polysilicon 688 -1594 688 -1594 0 3
rlabel polysilicon 695 -1588 695 -1588 0 1
rlabel polysilicon 695 -1594 695 -1594 0 3
rlabel polysilicon 702 -1588 702 -1588 0 1
rlabel polysilicon 705 -1588 705 -1588 0 2
rlabel polysilicon 702 -1594 702 -1594 0 3
rlabel polysilicon 705 -1594 705 -1594 0 4
rlabel polysilicon 709 -1588 709 -1588 0 1
rlabel polysilicon 709 -1594 709 -1594 0 3
rlabel polysilicon 716 -1588 716 -1588 0 1
rlabel polysilicon 716 -1594 716 -1594 0 3
rlabel polysilicon 723 -1588 723 -1588 0 1
rlabel polysilicon 723 -1594 723 -1594 0 3
rlabel polysilicon 730 -1588 730 -1588 0 1
rlabel polysilicon 730 -1594 730 -1594 0 3
rlabel polysilicon 737 -1588 737 -1588 0 1
rlabel polysilicon 737 -1594 737 -1594 0 3
rlabel polysilicon 744 -1588 744 -1588 0 1
rlabel polysilicon 744 -1594 744 -1594 0 3
rlabel polysilicon 751 -1588 751 -1588 0 1
rlabel polysilicon 751 -1594 751 -1594 0 3
rlabel polysilicon 758 -1588 758 -1588 0 1
rlabel polysilicon 758 -1594 758 -1594 0 3
rlabel polysilicon 765 -1588 765 -1588 0 1
rlabel polysilicon 765 -1594 765 -1594 0 3
rlabel polysilicon 772 -1588 772 -1588 0 1
rlabel polysilicon 772 -1594 772 -1594 0 3
rlabel polysilicon 779 -1588 779 -1588 0 1
rlabel polysilicon 779 -1594 779 -1594 0 3
rlabel polysilicon 786 -1588 786 -1588 0 1
rlabel polysilicon 786 -1594 786 -1594 0 3
rlabel polysilicon 793 -1588 793 -1588 0 1
rlabel polysilicon 793 -1594 793 -1594 0 3
rlabel polysilicon 800 -1588 800 -1588 0 1
rlabel polysilicon 803 -1588 803 -1588 0 2
rlabel polysilicon 800 -1594 800 -1594 0 3
rlabel polysilicon 803 -1594 803 -1594 0 4
rlabel polysilicon 807 -1588 807 -1588 0 1
rlabel polysilicon 807 -1594 807 -1594 0 3
rlabel polysilicon 814 -1588 814 -1588 0 1
rlabel polysilicon 814 -1594 814 -1594 0 3
rlabel polysilicon 821 -1588 821 -1588 0 1
rlabel polysilicon 821 -1594 821 -1594 0 3
rlabel polysilicon 828 -1588 828 -1588 0 1
rlabel polysilicon 831 -1588 831 -1588 0 2
rlabel polysilicon 828 -1594 828 -1594 0 3
rlabel polysilicon 831 -1594 831 -1594 0 4
rlabel polysilicon 835 -1588 835 -1588 0 1
rlabel polysilicon 835 -1594 835 -1594 0 3
rlabel polysilicon 842 -1588 842 -1588 0 1
rlabel polysilicon 842 -1594 842 -1594 0 3
rlabel polysilicon 849 -1588 849 -1588 0 1
rlabel polysilicon 849 -1594 849 -1594 0 3
rlabel polysilicon 856 -1588 856 -1588 0 1
rlabel polysilicon 859 -1588 859 -1588 0 2
rlabel polysilicon 856 -1594 856 -1594 0 3
rlabel polysilicon 859 -1594 859 -1594 0 4
rlabel polysilicon 863 -1588 863 -1588 0 1
rlabel polysilicon 863 -1594 863 -1594 0 3
rlabel polysilicon 870 -1588 870 -1588 0 1
rlabel polysilicon 870 -1594 870 -1594 0 3
rlabel polysilicon 877 -1588 877 -1588 0 1
rlabel polysilicon 877 -1594 877 -1594 0 3
rlabel polysilicon 884 -1588 884 -1588 0 1
rlabel polysilicon 884 -1594 884 -1594 0 3
rlabel polysilicon 891 -1588 891 -1588 0 1
rlabel polysilicon 894 -1588 894 -1588 0 2
rlabel polysilicon 898 -1588 898 -1588 0 1
rlabel polysilicon 898 -1594 898 -1594 0 3
rlabel polysilicon 905 -1588 905 -1588 0 1
rlabel polysilicon 905 -1594 905 -1594 0 3
rlabel polysilicon 912 -1588 912 -1588 0 1
rlabel polysilicon 912 -1594 912 -1594 0 3
rlabel polysilicon 919 -1588 919 -1588 0 1
rlabel polysilicon 919 -1594 919 -1594 0 3
rlabel polysilicon 926 -1588 926 -1588 0 1
rlabel polysilicon 926 -1594 926 -1594 0 3
rlabel polysilicon 933 -1588 933 -1588 0 1
rlabel polysilicon 933 -1594 933 -1594 0 3
rlabel polysilicon 940 -1588 940 -1588 0 1
rlabel polysilicon 940 -1594 940 -1594 0 3
rlabel polysilicon 947 -1588 947 -1588 0 1
rlabel polysilicon 947 -1594 947 -1594 0 3
rlabel polysilicon 954 -1588 954 -1588 0 1
rlabel polysilicon 954 -1594 954 -1594 0 3
rlabel polysilicon 961 -1588 961 -1588 0 1
rlabel polysilicon 961 -1594 961 -1594 0 3
rlabel polysilicon 968 -1588 968 -1588 0 1
rlabel polysilicon 968 -1594 968 -1594 0 3
rlabel polysilicon 975 -1588 975 -1588 0 1
rlabel polysilicon 975 -1594 975 -1594 0 3
rlabel polysilicon 982 -1588 982 -1588 0 1
rlabel polysilicon 982 -1594 982 -1594 0 3
rlabel polysilicon 989 -1588 989 -1588 0 1
rlabel polysilicon 989 -1594 989 -1594 0 3
rlabel polysilicon 996 -1588 996 -1588 0 1
rlabel polysilicon 996 -1594 996 -1594 0 3
rlabel polysilicon 1003 -1588 1003 -1588 0 1
rlabel polysilicon 1003 -1594 1003 -1594 0 3
rlabel polysilicon 1010 -1588 1010 -1588 0 1
rlabel polysilicon 1010 -1594 1010 -1594 0 3
rlabel polysilicon 1017 -1588 1017 -1588 0 1
rlabel polysilicon 1017 -1594 1017 -1594 0 3
rlabel polysilicon 1024 -1588 1024 -1588 0 1
rlabel polysilicon 1024 -1594 1024 -1594 0 3
rlabel polysilicon 1031 -1588 1031 -1588 0 1
rlabel polysilicon 1031 -1594 1031 -1594 0 3
rlabel polysilicon 1038 -1588 1038 -1588 0 1
rlabel polysilicon 1038 -1594 1038 -1594 0 3
rlabel polysilicon 1045 -1588 1045 -1588 0 1
rlabel polysilicon 1048 -1588 1048 -1588 0 2
rlabel polysilicon 1045 -1594 1045 -1594 0 3
rlabel polysilicon 1052 -1588 1052 -1588 0 1
rlabel polysilicon 1052 -1594 1052 -1594 0 3
rlabel polysilicon 1059 -1588 1059 -1588 0 1
rlabel polysilicon 1059 -1594 1059 -1594 0 3
rlabel polysilicon 1066 -1588 1066 -1588 0 1
rlabel polysilicon 1066 -1594 1066 -1594 0 3
rlabel polysilicon 1073 -1588 1073 -1588 0 1
rlabel polysilicon 1073 -1594 1073 -1594 0 3
rlabel polysilicon 1080 -1588 1080 -1588 0 1
rlabel polysilicon 1080 -1594 1080 -1594 0 3
rlabel polysilicon 1087 -1588 1087 -1588 0 1
rlabel polysilicon 1087 -1594 1087 -1594 0 3
rlabel polysilicon 1094 -1588 1094 -1588 0 1
rlabel polysilicon 1094 -1594 1094 -1594 0 3
rlabel polysilicon 1101 -1588 1101 -1588 0 1
rlabel polysilicon 1101 -1594 1101 -1594 0 3
rlabel polysilicon 1108 -1588 1108 -1588 0 1
rlabel polysilicon 1108 -1594 1108 -1594 0 3
rlabel polysilicon 1115 -1588 1115 -1588 0 1
rlabel polysilicon 1115 -1594 1115 -1594 0 3
rlabel polysilicon 1122 -1588 1122 -1588 0 1
rlabel polysilicon 1122 -1594 1122 -1594 0 3
rlabel polysilicon 1129 -1588 1129 -1588 0 1
rlabel polysilicon 1129 -1594 1129 -1594 0 3
rlabel polysilicon 1136 -1588 1136 -1588 0 1
rlabel polysilicon 1136 -1594 1136 -1594 0 3
rlabel polysilicon 1143 -1588 1143 -1588 0 1
rlabel polysilicon 1143 -1594 1143 -1594 0 3
rlabel polysilicon 1150 -1588 1150 -1588 0 1
rlabel polysilicon 1157 -1588 1157 -1588 0 1
rlabel polysilicon 1157 -1594 1157 -1594 0 3
rlabel polysilicon 1164 -1588 1164 -1588 0 1
rlabel polysilicon 1164 -1594 1164 -1594 0 3
rlabel polysilicon 1171 -1588 1171 -1588 0 1
rlabel polysilicon 1171 -1594 1171 -1594 0 3
rlabel polysilicon 1178 -1588 1178 -1588 0 1
rlabel polysilicon 1178 -1594 1178 -1594 0 3
rlabel polysilicon 1185 -1588 1185 -1588 0 1
rlabel polysilicon 1185 -1594 1185 -1594 0 3
rlabel polysilicon 1192 -1588 1192 -1588 0 1
rlabel polysilicon 1192 -1594 1192 -1594 0 3
rlabel polysilicon 1199 -1588 1199 -1588 0 1
rlabel polysilicon 1199 -1594 1199 -1594 0 3
rlabel polysilicon 1206 -1588 1206 -1588 0 1
rlabel polysilicon 1206 -1594 1206 -1594 0 3
rlabel polysilicon 1213 -1588 1213 -1588 0 1
rlabel polysilicon 1213 -1594 1213 -1594 0 3
rlabel polysilicon 1220 -1588 1220 -1588 0 1
rlabel polysilicon 1220 -1594 1220 -1594 0 3
rlabel polysilicon 1227 -1588 1227 -1588 0 1
rlabel polysilicon 1227 -1594 1227 -1594 0 3
rlabel polysilicon 1234 -1588 1234 -1588 0 1
rlabel polysilicon 1234 -1594 1234 -1594 0 3
rlabel polysilicon 1241 -1588 1241 -1588 0 1
rlabel polysilicon 1241 -1594 1241 -1594 0 3
rlabel polysilicon 1248 -1588 1248 -1588 0 1
rlabel polysilicon 1248 -1594 1248 -1594 0 3
rlabel polysilicon 1255 -1588 1255 -1588 0 1
rlabel polysilicon 1255 -1594 1255 -1594 0 3
rlabel polysilicon 1258 -1594 1258 -1594 0 4
rlabel polysilicon 1262 -1588 1262 -1588 0 1
rlabel polysilicon 1262 -1594 1262 -1594 0 3
rlabel polysilicon 1269 -1588 1269 -1588 0 1
rlabel polysilicon 1269 -1594 1269 -1594 0 3
rlabel polysilicon 1276 -1588 1276 -1588 0 1
rlabel polysilicon 1276 -1594 1276 -1594 0 3
rlabel polysilicon 1283 -1588 1283 -1588 0 1
rlabel polysilicon 1283 -1594 1283 -1594 0 3
rlabel polysilicon 1290 -1588 1290 -1588 0 1
rlabel polysilicon 1290 -1594 1290 -1594 0 3
rlabel polysilicon 1297 -1588 1297 -1588 0 1
rlabel polysilicon 1297 -1594 1297 -1594 0 3
rlabel polysilicon 1304 -1588 1304 -1588 0 1
rlabel polysilicon 1304 -1594 1304 -1594 0 3
rlabel polysilicon 1311 -1588 1311 -1588 0 1
rlabel polysilicon 1311 -1594 1311 -1594 0 3
rlabel polysilicon 1318 -1588 1318 -1588 0 1
rlabel polysilicon 1318 -1594 1318 -1594 0 3
rlabel polysilicon 1325 -1588 1325 -1588 0 1
rlabel polysilicon 1325 -1594 1325 -1594 0 3
rlabel polysilicon 1332 -1588 1332 -1588 0 1
rlabel polysilicon 1332 -1594 1332 -1594 0 3
rlabel polysilicon 1339 -1588 1339 -1588 0 1
rlabel polysilicon 1339 -1594 1339 -1594 0 3
rlabel polysilicon 1346 -1588 1346 -1588 0 1
rlabel polysilicon 1346 -1594 1346 -1594 0 3
rlabel polysilicon 1353 -1588 1353 -1588 0 1
rlabel polysilicon 1353 -1594 1353 -1594 0 3
rlabel polysilicon 2 -1719 2 -1719 0 1
rlabel polysilicon 2 -1725 2 -1725 0 3
rlabel polysilicon 9 -1719 9 -1719 0 1
rlabel polysilicon 9 -1725 9 -1725 0 3
rlabel polysilicon 16 -1725 16 -1725 0 3
rlabel polysilicon 19 -1725 19 -1725 0 4
rlabel polysilicon 23 -1725 23 -1725 0 3
rlabel polysilicon 26 -1725 26 -1725 0 4
rlabel polysilicon 30 -1719 30 -1719 0 1
rlabel polysilicon 30 -1725 30 -1725 0 3
rlabel polysilicon 33 -1725 33 -1725 0 4
rlabel polysilicon 37 -1719 37 -1719 0 1
rlabel polysilicon 37 -1725 37 -1725 0 3
rlabel polysilicon 44 -1719 44 -1719 0 1
rlabel polysilicon 47 -1719 47 -1719 0 2
rlabel polysilicon 44 -1725 44 -1725 0 3
rlabel polysilicon 51 -1719 51 -1719 0 1
rlabel polysilicon 54 -1719 54 -1719 0 2
rlabel polysilicon 51 -1725 51 -1725 0 3
rlabel polysilicon 54 -1725 54 -1725 0 4
rlabel polysilicon 58 -1719 58 -1719 0 1
rlabel polysilicon 58 -1725 58 -1725 0 3
rlabel polysilicon 65 -1719 65 -1719 0 1
rlabel polysilicon 65 -1725 65 -1725 0 3
rlabel polysilicon 72 -1719 72 -1719 0 1
rlabel polysilicon 72 -1725 72 -1725 0 3
rlabel polysilicon 79 -1719 79 -1719 0 1
rlabel polysilicon 79 -1725 79 -1725 0 3
rlabel polysilicon 86 -1719 86 -1719 0 1
rlabel polysilicon 86 -1725 86 -1725 0 3
rlabel polysilicon 93 -1719 93 -1719 0 1
rlabel polysilicon 96 -1719 96 -1719 0 2
rlabel polysilicon 93 -1725 93 -1725 0 3
rlabel polysilicon 96 -1725 96 -1725 0 4
rlabel polysilicon 100 -1719 100 -1719 0 1
rlabel polysilicon 100 -1725 100 -1725 0 3
rlabel polysilicon 107 -1719 107 -1719 0 1
rlabel polysilicon 110 -1719 110 -1719 0 2
rlabel polysilicon 107 -1725 107 -1725 0 3
rlabel polysilicon 110 -1725 110 -1725 0 4
rlabel polysilicon 114 -1719 114 -1719 0 1
rlabel polysilicon 114 -1725 114 -1725 0 3
rlabel polysilicon 121 -1719 121 -1719 0 1
rlabel polysilicon 121 -1725 121 -1725 0 3
rlabel polysilicon 128 -1719 128 -1719 0 1
rlabel polysilicon 128 -1725 128 -1725 0 3
rlabel polysilicon 135 -1719 135 -1719 0 1
rlabel polysilicon 135 -1725 135 -1725 0 3
rlabel polysilicon 142 -1719 142 -1719 0 1
rlabel polysilicon 142 -1725 142 -1725 0 3
rlabel polysilicon 149 -1719 149 -1719 0 1
rlabel polysilicon 152 -1719 152 -1719 0 2
rlabel polysilicon 149 -1725 149 -1725 0 3
rlabel polysilicon 152 -1725 152 -1725 0 4
rlabel polysilicon 159 -1719 159 -1719 0 2
rlabel polysilicon 156 -1725 156 -1725 0 3
rlabel polysilicon 159 -1725 159 -1725 0 4
rlabel polysilicon 163 -1719 163 -1719 0 1
rlabel polysilicon 163 -1725 163 -1725 0 3
rlabel polysilicon 170 -1719 170 -1719 0 1
rlabel polysilicon 170 -1725 170 -1725 0 3
rlabel polysilicon 177 -1719 177 -1719 0 1
rlabel polysilicon 177 -1725 177 -1725 0 3
rlabel polysilicon 184 -1719 184 -1719 0 1
rlabel polysilicon 184 -1725 184 -1725 0 3
rlabel polysilicon 191 -1719 191 -1719 0 1
rlabel polysilicon 194 -1719 194 -1719 0 2
rlabel polysilicon 191 -1725 191 -1725 0 3
rlabel polysilicon 194 -1725 194 -1725 0 4
rlabel polysilicon 198 -1719 198 -1719 0 1
rlabel polysilicon 198 -1725 198 -1725 0 3
rlabel polysilicon 205 -1719 205 -1719 0 1
rlabel polysilicon 205 -1725 205 -1725 0 3
rlabel polysilicon 212 -1719 212 -1719 0 1
rlabel polysilicon 212 -1725 212 -1725 0 3
rlabel polysilicon 219 -1719 219 -1719 0 1
rlabel polysilicon 219 -1725 219 -1725 0 3
rlabel polysilicon 226 -1719 226 -1719 0 1
rlabel polysilicon 226 -1725 226 -1725 0 3
rlabel polysilicon 233 -1719 233 -1719 0 1
rlabel polysilicon 233 -1725 233 -1725 0 3
rlabel polysilicon 240 -1719 240 -1719 0 1
rlabel polysilicon 240 -1725 240 -1725 0 3
rlabel polysilicon 247 -1719 247 -1719 0 1
rlabel polysilicon 247 -1725 247 -1725 0 3
rlabel polysilicon 254 -1719 254 -1719 0 1
rlabel polysilicon 254 -1725 254 -1725 0 3
rlabel polysilicon 261 -1719 261 -1719 0 1
rlabel polysilicon 261 -1725 261 -1725 0 3
rlabel polysilicon 268 -1719 268 -1719 0 1
rlabel polysilicon 268 -1725 268 -1725 0 3
rlabel polysilicon 275 -1719 275 -1719 0 1
rlabel polysilicon 275 -1725 275 -1725 0 3
rlabel polysilicon 282 -1719 282 -1719 0 1
rlabel polysilicon 282 -1725 282 -1725 0 3
rlabel polysilicon 289 -1719 289 -1719 0 1
rlabel polysilicon 289 -1725 289 -1725 0 3
rlabel polysilicon 296 -1719 296 -1719 0 1
rlabel polysilicon 296 -1725 296 -1725 0 3
rlabel polysilicon 303 -1719 303 -1719 0 1
rlabel polysilicon 303 -1725 303 -1725 0 3
rlabel polysilicon 310 -1719 310 -1719 0 1
rlabel polysilicon 310 -1725 310 -1725 0 3
rlabel polysilicon 317 -1719 317 -1719 0 1
rlabel polysilicon 320 -1719 320 -1719 0 2
rlabel polysilicon 317 -1725 317 -1725 0 3
rlabel polysilicon 320 -1725 320 -1725 0 4
rlabel polysilicon 324 -1719 324 -1719 0 1
rlabel polysilicon 324 -1725 324 -1725 0 3
rlabel polysilicon 331 -1719 331 -1719 0 1
rlabel polysilicon 331 -1725 331 -1725 0 3
rlabel polysilicon 338 -1719 338 -1719 0 1
rlabel polysilicon 338 -1725 338 -1725 0 3
rlabel polysilicon 345 -1719 345 -1719 0 1
rlabel polysilicon 345 -1725 345 -1725 0 3
rlabel polysilicon 352 -1719 352 -1719 0 1
rlabel polysilicon 352 -1725 352 -1725 0 3
rlabel polysilicon 359 -1719 359 -1719 0 1
rlabel polysilicon 359 -1725 359 -1725 0 3
rlabel polysilicon 366 -1719 366 -1719 0 1
rlabel polysilicon 366 -1725 366 -1725 0 3
rlabel polysilicon 373 -1719 373 -1719 0 1
rlabel polysilicon 376 -1719 376 -1719 0 2
rlabel polysilicon 373 -1725 373 -1725 0 3
rlabel polysilicon 376 -1725 376 -1725 0 4
rlabel polysilicon 380 -1719 380 -1719 0 1
rlabel polysilicon 380 -1725 380 -1725 0 3
rlabel polysilicon 387 -1719 387 -1719 0 1
rlabel polysilicon 387 -1725 387 -1725 0 3
rlabel polysilicon 394 -1719 394 -1719 0 1
rlabel polysilicon 394 -1725 394 -1725 0 3
rlabel polysilicon 401 -1719 401 -1719 0 1
rlabel polysilicon 404 -1719 404 -1719 0 2
rlabel polysilicon 401 -1725 401 -1725 0 3
rlabel polysilicon 404 -1725 404 -1725 0 4
rlabel polysilicon 408 -1719 408 -1719 0 1
rlabel polysilicon 408 -1725 408 -1725 0 3
rlabel polysilicon 415 -1719 415 -1719 0 1
rlabel polysilicon 415 -1725 415 -1725 0 3
rlabel polysilicon 422 -1719 422 -1719 0 1
rlabel polysilicon 422 -1725 422 -1725 0 3
rlabel polysilicon 429 -1719 429 -1719 0 1
rlabel polysilicon 429 -1725 429 -1725 0 3
rlabel polysilicon 436 -1719 436 -1719 0 1
rlabel polysilicon 436 -1725 436 -1725 0 3
rlabel polysilicon 443 -1719 443 -1719 0 1
rlabel polysilicon 443 -1725 443 -1725 0 3
rlabel polysilicon 450 -1719 450 -1719 0 1
rlabel polysilicon 450 -1725 450 -1725 0 3
rlabel polysilicon 457 -1719 457 -1719 0 1
rlabel polysilicon 460 -1719 460 -1719 0 2
rlabel polysilicon 457 -1725 457 -1725 0 3
rlabel polysilicon 460 -1725 460 -1725 0 4
rlabel polysilicon 464 -1719 464 -1719 0 1
rlabel polysilicon 464 -1725 464 -1725 0 3
rlabel polysilicon 471 -1719 471 -1719 0 1
rlabel polysilicon 471 -1725 471 -1725 0 3
rlabel polysilicon 478 -1719 478 -1719 0 1
rlabel polysilicon 478 -1725 478 -1725 0 3
rlabel polysilicon 485 -1719 485 -1719 0 1
rlabel polysilicon 488 -1719 488 -1719 0 2
rlabel polysilicon 485 -1725 485 -1725 0 3
rlabel polysilicon 488 -1725 488 -1725 0 4
rlabel polysilicon 492 -1719 492 -1719 0 1
rlabel polysilicon 492 -1725 492 -1725 0 3
rlabel polysilicon 499 -1719 499 -1719 0 1
rlabel polysilicon 499 -1725 499 -1725 0 3
rlabel polysilicon 506 -1719 506 -1719 0 1
rlabel polysilicon 506 -1725 506 -1725 0 3
rlabel polysilicon 513 -1719 513 -1719 0 1
rlabel polysilicon 513 -1725 513 -1725 0 3
rlabel polysilicon 520 -1719 520 -1719 0 1
rlabel polysilicon 523 -1719 523 -1719 0 2
rlabel polysilicon 520 -1725 520 -1725 0 3
rlabel polysilicon 523 -1725 523 -1725 0 4
rlabel polysilicon 527 -1719 527 -1719 0 1
rlabel polysilicon 527 -1725 527 -1725 0 3
rlabel polysilicon 534 -1719 534 -1719 0 1
rlabel polysilicon 534 -1725 534 -1725 0 3
rlabel polysilicon 541 -1719 541 -1719 0 1
rlabel polysilicon 541 -1725 541 -1725 0 3
rlabel polysilicon 551 -1719 551 -1719 0 2
rlabel polysilicon 548 -1725 548 -1725 0 3
rlabel polysilicon 551 -1725 551 -1725 0 4
rlabel polysilicon 555 -1719 555 -1719 0 1
rlabel polysilicon 555 -1725 555 -1725 0 3
rlabel polysilicon 558 -1725 558 -1725 0 4
rlabel polysilicon 562 -1719 562 -1719 0 1
rlabel polysilicon 562 -1725 562 -1725 0 3
rlabel polysilicon 569 -1719 569 -1719 0 1
rlabel polysilicon 569 -1725 569 -1725 0 3
rlabel polysilicon 576 -1719 576 -1719 0 1
rlabel polysilicon 576 -1725 576 -1725 0 3
rlabel polysilicon 583 -1719 583 -1719 0 1
rlabel polysilicon 583 -1725 583 -1725 0 3
rlabel polysilicon 590 -1719 590 -1719 0 1
rlabel polysilicon 590 -1725 590 -1725 0 3
rlabel polysilicon 597 -1719 597 -1719 0 1
rlabel polysilicon 597 -1725 597 -1725 0 3
rlabel polysilicon 604 -1719 604 -1719 0 1
rlabel polysilicon 604 -1725 604 -1725 0 3
rlabel polysilicon 611 -1719 611 -1719 0 1
rlabel polysilicon 611 -1725 611 -1725 0 3
rlabel polysilicon 618 -1719 618 -1719 0 1
rlabel polysilicon 618 -1725 618 -1725 0 3
rlabel polysilicon 625 -1719 625 -1719 0 1
rlabel polysilicon 625 -1725 625 -1725 0 3
rlabel polysilicon 632 -1719 632 -1719 0 1
rlabel polysilicon 632 -1725 632 -1725 0 3
rlabel polysilicon 639 -1719 639 -1719 0 1
rlabel polysilicon 639 -1725 639 -1725 0 3
rlabel polysilicon 646 -1719 646 -1719 0 1
rlabel polysilicon 646 -1725 646 -1725 0 3
rlabel polysilicon 653 -1719 653 -1719 0 1
rlabel polysilicon 653 -1725 653 -1725 0 3
rlabel polysilicon 660 -1719 660 -1719 0 1
rlabel polysilicon 660 -1725 660 -1725 0 3
rlabel polysilicon 667 -1719 667 -1719 0 1
rlabel polysilicon 670 -1719 670 -1719 0 2
rlabel polysilicon 667 -1725 667 -1725 0 3
rlabel polysilicon 674 -1719 674 -1719 0 1
rlabel polysilicon 674 -1725 674 -1725 0 3
rlabel polysilicon 681 -1719 681 -1719 0 1
rlabel polysilicon 681 -1725 681 -1725 0 3
rlabel polysilicon 688 -1719 688 -1719 0 1
rlabel polysilicon 688 -1725 688 -1725 0 3
rlabel polysilicon 695 -1719 695 -1719 0 1
rlabel polysilicon 695 -1725 695 -1725 0 3
rlabel polysilicon 702 -1719 702 -1719 0 1
rlabel polysilicon 702 -1725 702 -1725 0 3
rlabel polysilicon 709 -1719 709 -1719 0 1
rlabel polysilicon 709 -1725 709 -1725 0 3
rlabel polysilicon 716 -1719 716 -1719 0 1
rlabel polysilicon 716 -1725 716 -1725 0 3
rlabel polysilicon 723 -1719 723 -1719 0 1
rlabel polysilicon 723 -1725 723 -1725 0 3
rlabel polysilicon 730 -1719 730 -1719 0 1
rlabel polysilicon 730 -1725 730 -1725 0 3
rlabel polysilicon 737 -1719 737 -1719 0 1
rlabel polysilicon 737 -1725 737 -1725 0 3
rlabel polysilicon 744 -1719 744 -1719 0 1
rlabel polysilicon 747 -1719 747 -1719 0 2
rlabel polysilicon 744 -1725 744 -1725 0 3
rlabel polysilicon 747 -1725 747 -1725 0 4
rlabel polysilicon 751 -1719 751 -1719 0 1
rlabel polysilicon 754 -1719 754 -1719 0 2
rlabel polysilicon 751 -1725 751 -1725 0 3
rlabel polysilicon 754 -1725 754 -1725 0 4
rlabel polysilicon 758 -1719 758 -1719 0 1
rlabel polysilicon 758 -1725 758 -1725 0 3
rlabel polysilicon 765 -1719 765 -1719 0 1
rlabel polysilicon 765 -1725 765 -1725 0 3
rlabel polysilicon 772 -1719 772 -1719 0 1
rlabel polysilicon 775 -1719 775 -1719 0 2
rlabel polysilicon 772 -1725 772 -1725 0 3
rlabel polysilicon 775 -1725 775 -1725 0 4
rlabel polysilicon 779 -1719 779 -1719 0 1
rlabel polysilicon 779 -1725 779 -1725 0 3
rlabel polysilicon 786 -1719 786 -1719 0 1
rlabel polysilicon 786 -1725 786 -1725 0 3
rlabel polysilicon 793 -1719 793 -1719 0 1
rlabel polysilicon 793 -1725 793 -1725 0 3
rlabel polysilicon 800 -1719 800 -1719 0 1
rlabel polysilicon 800 -1725 800 -1725 0 3
rlabel polysilicon 807 -1719 807 -1719 0 1
rlabel polysilicon 807 -1725 807 -1725 0 3
rlabel polysilicon 814 -1719 814 -1719 0 1
rlabel polysilicon 814 -1725 814 -1725 0 3
rlabel polysilicon 821 -1719 821 -1719 0 1
rlabel polysilicon 821 -1725 821 -1725 0 3
rlabel polysilicon 828 -1719 828 -1719 0 1
rlabel polysilicon 828 -1725 828 -1725 0 3
rlabel polysilicon 835 -1719 835 -1719 0 1
rlabel polysilicon 835 -1725 835 -1725 0 3
rlabel polysilicon 842 -1719 842 -1719 0 1
rlabel polysilicon 842 -1725 842 -1725 0 3
rlabel polysilicon 849 -1719 849 -1719 0 1
rlabel polysilicon 849 -1725 849 -1725 0 3
rlabel polysilicon 856 -1719 856 -1719 0 1
rlabel polysilicon 856 -1725 856 -1725 0 3
rlabel polysilicon 863 -1719 863 -1719 0 1
rlabel polysilicon 863 -1725 863 -1725 0 3
rlabel polysilicon 870 -1719 870 -1719 0 1
rlabel polysilicon 870 -1725 870 -1725 0 3
rlabel polysilicon 877 -1719 877 -1719 0 1
rlabel polysilicon 877 -1725 877 -1725 0 3
rlabel polysilicon 884 -1719 884 -1719 0 1
rlabel polysilicon 884 -1725 884 -1725 0 3
rlabel polysilicon 891 -1719 891 -1719 0 1
rlabel polysilicon 894 -1719 894 -1719 0 2
rlabel polysilicon 894 -1725 894 -1725 0 4
rlabel polysilicon 898 -1719 898 -1719 0 1
rlabel polysilicon 901 -1719 901 -1719 0 2
rlabel polysilicon 898 -1725 898 -1725 0 3
rlabel polysilicon 901 -1725 901 -1725 0 4
rlabel polysilicon 905 -1719 905 -1719 0 1
rlabel polysilicon 905 -1725 905 -1725 0 3
rlabel polysilicon 912 -1719 912 -1719 0 1
rlabel polysilicon 912 -1725 912 -1725 0 3
rlabel polysilicon 919 -1719 919 -1719 0 1
rlabel polysilicon 919 -1725 919 -1725 0 3
rlabel polysilicon 926 -1719 926 -1719 0 1
rlabel polysilicon 926 -1725 926 -1725 0 3
rlabel polysilicon 933 -1719 933 -1719 0 1
rlabel polysilicon 933 -1725 933 -1725 0 3
rlabel polysilicon 940 -1719 940 -1719 0 1
rlabel polysilicon 940 -1725 940 -1725 0 3
rlabel polysilicon 943 -1725 943 -1725 0 4
rlabel polysilicon 947 -1719 947 -1719 0 1
rlabel polysilicon 947 -1725 947 -1725 0 3
rlabel polysilicon 954 -1719 954 -1719 0 1
rlabel polysilicon 954 -1725 954 -1725 0 3
rlabel polysilicon 961 -1719 961 -1719 0 1
rlabel polysilicon 961 -1725 961 -1725 0 3
rlabel polysilicon 968 -1719 968 -1719 0 1
rlabel polysilicon 968 -1725 968 -1725 0 3
rlabel polysilicon 975 -1719 975 -1719 0 1
rlabel polysilicon 975 -1725 975 -1725 0 3
rlabel polysilicon 982 -1719 982 -1719 0 1
rlabel polysilicon 982 -1725 982 -1725 0 3
rlabel polysilicon 989 -1719 989 -1719 0 1
rlabel polysilicon 989 -1725 989 -1725 0 3
rlabel polysilicon 996 -1719 996 -1719 0 1
rlabel polysilicon 996 -1725 996 -1725 0 3
rlabel polysilicon 1003 -1719 1003 -1719 0 1
rlabel polysilicon 1003 -1725 1003 -1725 0 3
rlabel polysilicon 1010 -1719 1010 -1719 0 1
rlabel polysilicon 1010 -1725 1010 -1725 0 3
rlabel polysilicon 1017 -1719 1017 -1719 0 1
rlabel polysilicon 1017 -1725 1017 -1725 0 3
rlabel polysilicon 1024 -1719 1024 -1719 0 1
rlabel polysilicon 1024 -1725 1024 -1725 0 3
rlabel polysilicon 1031 -1719 1031 -1719 0 1
rlabel polysilicon 1031 -1725 1031 -1725 0 3
rlabel polysilicon 1038 -1719 1038 -1719 0 1
rlabel polysilicon 1038 -1725 1038 -1725 0 3
rlabel polysilicon 1045 -1719 1045 -1719 0 1
rlabel polysilicon 1045 -1725 1045 -1725 0 3
rlabel polysilicon 1052 -1719 1052 -1719 0 1
rlabel polysilicon 1052 -1725 1052 -1725 0 3
rlabel polysilicon 1059 -1719 1059 -1719 0 1
rlabel polysilicon 1059 -1725 1059 -1725 0 3
rlabel polysilicon 1066 -1719 1066 -1719 0 1
rlabel polysilicon 1066 -1725 1066 -1725 0 3
rlabel polysilicon 1069 -1725 1069 -1725 0 4
rlabel polysilicon 1073 -1719 1073 -1719 0 1
rlabel polysilicon 1073 -1725 1073 -1725 0 3
rlabel polysilicon 1080 -1719 1080 -1719 0 1
rlabel polysilicon 1080 -1725 1080 -1725 0 3
rlabel polysilicon 1087 -1719 1087 -1719 0 1
rlabel polysilicon 1087 -1725 1087 -1725 0 3
rlabel polysilicon 1094 -1719 1094 -1719 0 1
rlabel polysilicon 1094 -1725 1094 -1725 0 3
rlabel polysilicon 1101 -1719 1101 -1719 0 1
rlabel polysilicon 1101 -1725 1101 -1725 0 3
rlabel polysilicon 1108 -1719 1108 -1719 0 1
rlabel polysilicon 1108 -1725 1108 -1725 0 3
rlabel polysilicon 1115 -1719 1115 -1719 0 1
rlabel polysilicon 1115 -1725 1115 -1725 0 3
rlabel polysilicon 1122 -1725 1122 -1725 0 3
rlabel polysilicon 1125 -1725 1125 -1725 0 4
rlabel polysilicon 1129 -1719 1129 -1719 0 1
rlabel polysilicon 1129 -1725 1129 -1725 0 3
rlabel polysilicon 1136 -1719 1136 -1719 0 1
rlabel polysilicon 1136 -1725 1136 -1725 0 3
rlabel polysilicon 1143 -1719 1143 -1719 0 1
rlabel polysilicon 1143 -1725 1143 -1725 0 3
rlabel polysilicon 1150 -1725 1150 -1725 0 3
rlabel polysilicon 1157 -1719 1157 -1719 0 1
rlabel polysilicon 1157 -1725 1157 -1725 0 3
rlabel polysilicon 1164 -1719 1164 -1719 0 1
rlabel polysilicon 1164 -1725 1164 -1725 0 3
rlabel polysilicon 1171 -1719 1171 -1719 0 1
rlabel polysilicon 1171 -1725 1171 -1725 0 3
rlabel polysilicon 1178 -1719 1178 -1719 0 1
rlabel polysilicon 1178 -1725 1178 -1725 0 3
rlabel polysilicon 1185 -1719 1185 -1719 0 1
rlabel polysilicon 1185 -1725 1185 -1725 0 3
rlabel polysilicon 1192 -1719 1192 -1719 0 1
rlabel polysilicon 1192 -1725 1192 -1725 0 3
rlabel polysilicon 1199 -1719 1199 -1719 0 1
rlabel polysilicon 1199 -1725 1199 -1725 0 3
rlabel polysilicon 1206 -1719 1206 -1719 0 1
rlabel polysilicon 1206 -1725 1206 -1725 0 3
rlabel polysilicon 1213 -1719 1213 -1719 0 1
rlabel polysilicon 1213 -1725 1213 -1725 0 3
rlabel polysilicon 1220 -1719 1220 -1719 0 1
rlabel polysilicon 1220 -1725 1220 -1725 0 3
rlabel polysilicon 1227 -1719 1227 -1719 0 1
rlabel polysilicon 1227 -1725 1227 -1725 0 3
rlabel polysilicon 1234 -1719 1234 -1719 0 1
rlabel polysilicon 1234 -1725 1234 -1725 0 3
rlabel polysilicon 1241 -1719 1241 -1719 0 1
rlabel polysilicon 1241 -1725 1241 -1725 0 3
rlabel polysilicon 1248 -1719 1248 -1719 0 1
rlabel polysilicon 1248 -1725 1248 -1725 0 3
rlabel polysilicon 1255 -1719 1255 -1719 0 1
rlabel polysilicon 1258 -1719 1258 -1719 0 2
rlabel polysilicon 1255 -1725 1255 -1725 0 3
rlabel polysilicon 1262 -1719 1262 -1719 0 1
rlabel polysilicon 1262 -1725 1262 -1725 0 3
rlabel polysilicon 1269 -1719 1269 -1719 0 1
rlabel polysilicon 1269 -1725 1269 -1725 0 3
rlabel polysilicon 1276 -1719 1276 -1719 0 1
rlabel polysilicon 1276 -1725 1276 -1725 0 3
rlabel polysilicon 1283 -1719 1283 -1719 0 1
rlabel polysilicon 1283 -1725 1283 -1725 0 3
rlabel polysilicon 1290 -1719 1290 -1719 0 1
rlabel polysilicon 1290 -1725 1290 -1725 0 3
rlabel polysilicon 1297 -1719 1297 -1719 0 1
rlabel polysilicon 1297 -1725 1297 -1725 0 3
rlabel polysilicon 1304 -1719 1304 -1719 0 1
rlabel polysilicon 1304 -1725 1304 -1725 0 3
rlabel polysilicon 1311 -1719 1311 -1719 0 1
rlabel polysilicon 1311 -1725 1311 -1725 0 3
rlabel polysilicon 1318 -1719 1318 -1719 0 1
rlabel polysilicon 1318 -1725 1318 -1725 0 3
rlabel polysilicon 1325 -1719 1325 -1719 0 1
rlabel polysilicon 1328 -1719 1328 -1719 0 2
rlabel polysilicon 1328 -1725 1328 -1725 0 4
rlabel polysilicon 2 -1838 2 -1838 0 1
rlabel polysilicon 2 -1844 2 -1844 0 3
rlabel polysilicon 9 -1838 9 -1838 0 1
rlabel polysilicon 9 -1844 9 -1844 0 3
rlabel polysilicon 16 -1838 16 -1838 0 1
rlabel polysilicon 16 -1844 16 -1844 0 3
rlabel polysilicon 23 -1838 23 -1838 0 1
rlabel polysilicon 26 -1838 26 -1838 0 2
rlabel polysilicon 23 -1844 23 -1844 0 3
rlabel polysilicon 30 -1838 30 -1838 0 1
rlabel polysilicon 30 -1844 30 -1844 0 3
rlabel polysilicon 40 -1838 40 -1838 0 2
rlabel polysilicon 37 -1844 37 -1844 0 3
rlabel polysilicon 40 -1844 40 -1844 0 4
rlabel polysilicon 44 -1838 44 -1838 0 1
rlabel polysilicon 47 -1838 47 -1838 0 2
rlabel polysilicon 44 -1844 44 -1844 0 3
rlabel polysilicon 47 -1844 47 -1844 0 4
rlabel polysilicon 51 -1838 51 -1838 0 1
rlabel polysilicon 54 -1838 54 -1838 0 2
rlabel polysilicon 51 -1844 51 -1844 0 3
rlabel polysilicon 54 -1844 54 -1844 0 4
rlabel polysilicon 58 -1838 58 -1838 0 1
rlabel polysilicon 58 -1844 58 -1844 0 3
rlabel polysilicon 65 -1838 65 -1838 0 1
rlabel polysilicon 68 -1838 68 -1838 0 2
rlabel polysilicon 68 -1844 68 -1844 0 4
rlabel polysilicon 72 -1838 72 -1838 0 1
rlabel polysilicon 72 -1844 72 -1844 0 3
rlabel polysilicon 79 -1838 79 -1838 0 1
rlabel polysilicon 79 -1844 79 -1844 0 3
rlabel polysilicon 86 -1838 86 -1838 0 1
rlabel polysilicon 86 -1844 86 -1844 0 3
rlabel polysilicon 93 -1838 93 -1838 0 1
rlabel polysilicon 93 -1844 93 -1844 0 3
rlabel polysilicon 100 -1838 100 -1838 0 1
rlabel polysilicon 100 -1844 100 -1844 0 3
rlabel polysilicon 107 -1838 107 -1838 0 1
rlabel polysilicon 107 -1844 107 -1844 0 3
rlabel polysilicon 114 -1838 114 -1838 0 1
rlabel polysilicon 117 -1838 117 -1838 0 2
rlabel polysilicon 114 -1844 114 -1844 0 3
rlabel polysilicon 121 -1838 121 -1838 0 1
rlabel polysilicon 121 -1844 121 -1844 0 3
rlabel polysilicon 128 -1838 128 -1838 0 1
rlabel polysilicon 128 -1844 128 -1844 0 3
rlabel polysilicon 135 -1838 135 -1838 0 1
rlabel polysilicon 138 -1838 138 -1838 0 2
rlabel polysilicon 135 -1844 135 -1844 0 3
rlabel polysilicon 138 -1844 138 -1844 0 4
rlabel polysilicon 142 -1838 142 -1838 0 1
rlabel polysilicon 142 -1844 142 -1844 0 3
rlabel polysilicon 149 -1838 149 -1838 0 1
rlabel polysilicon 152 -1838 152 -1838 0 2
rlabel polysilicon 149 -1844 149 -1844 0 3
rlabel polysilicon 152 -1844 152 -1844 0 4
rlabel polysilicon 156 -1838 156 -1838 0 1
rlabel polysilicon 156 -1844 156 -1844 0 3
rlabel polysilicon 163 -1838 163 -1838 0 1
rlabel polysilicon 163 -1844 163 -1844 0 3
rlabel polysilicon 170 -1838 170 -1838 0 1
rlabel polysilicon 170 -1844 170 -1844 0 3
rlabel polysilicon 177 -1838 177 -1838 0 1
rlabel polysilicon 177 -1844 177 -1844 0 3
rlabel polysilicon 184 -1838 184 -1838 0 1
rlabel polysilicon 184 -1844 184 -1844 0 3
rlabel polysilicon 191 -1838 191 -1838 0 1
rlabel polysilicon 191 -1844 191 -1844 0 3
rlabel polysilicon 198 -1838 198 -1838 0 1
rlabel polysilicon 198 -1844 198 -1844 0 3
rlabel polysilicon 205 -1838 205 -1838 0 1
rlabel polysilicon 205 -1844 205 -1844 0 3
rlabel polysilicon 212 -1838 212 -1838 0 1
rlabel polysilicon 212 -1844 212 -1844 0 3
rlabel polysilicon 219 -1838 219 -1838 0 1
rlabel polysilicon 219 -1844 219 -1844 0 3
rlabel polysilicon 226 -1838 226 -1838 0 1
rlabel polysilicon 226 -1844 226 -1844 0 3
rlabel polysilicon 233 -1838 233 -1838 0 1
rlabel polysilicon 233 -1844 233 -1844 0 3
rlabel polysilicon 240 -1838 240 -1838 0 1
rlabel polysilicon 240 -1844 240 -1844 0 3
rlabel polysilicon 247 -1838 247 -1838 0 1
rlabel polysilicon 247 -1844 247 -1844 0 3
rlabel polysilicon 254 -1838 254 -1838 0 1
rlabel polysilicon 254 -1844 254 -1844 0 3
rlabel polysilicon 261 -1838 261 -1838 0 1
rlabel polysilicon 261 -1844 261 -1844 0 3
rlabel polysilicon 268 -1838 268 -1838 0 1
rlabel polysilicon 268 -1844 268 -1844 0 3
rlabel polysilicon 275 -1838 275 -1838 0 1
rlabel polysilicon 275 -1844 275 -1844 0 3
rlabel polysilicon 282 -1838 282 -1838 0 1
rlabel polysilicon 282 -1844 282 -1844 0 3
rlabel polysilicon 289 -1838 289 -1838 0 1
rlabel polysilicon 289 -1844 289 -1844 0 3
rlabel polysilicon 296 -1838 296 -1838 0 1
rlabel polysilicon 299 -1838 299 -1838 0 2
rlabel polysilicon 296 -1844 296 -1844 0 3
rlabel polysilicon 299 -1844 299 -1844 0 4
rlabel polysilicon 303 -1838 303 -1838 0 1
rlabel polysilicon 303 -1844 303 -1844 0 3
rlabel polysilicon 310 -1838 310 -1838 0 1
rlabel polysilicon 310 -1844 310 -1844 0 3
rlabel polysilicon 317 -1838 317 -1838 0 1
rlabel polysilicon 317 -1844 317 -1844 0 3
rlabel polysilicon 324 -1838 324 -1838 0 1
rlabel polysilicon 324 -1844 324 -1844 0 3
rlabel polysilicon 331 -1838 331 -1838 0 1
rlabel polysilicon 331 -1844 331 -1844 0 3
rlabel polysilicon 338 -1838 338 -1838 0 1
rlabel polysilicon 338 -1844 338 -1844 0 3
rlabel polysilicon 345 -1838 345 -1838 0 1
rlabel polysilicon 345 -1844 345 -1844 0 3
rlabel polysilicon 352 -1838 352 -1838 0 1
rlabel polysilicon 355 -1838 355 -1838 0 2
rlabel polysilicon 352 -1844 352 -1844 0 3
rlabel polysilicon 355 -1844 355 -1844 0 4
rlabel polysilicon 359 -1838 359 -1838 0 1
rlabel polysilicon 359 -1844 359 -1844 0 3
rlabel polysilicon 366 -1838 366 -1838 0 1
rlabel polysilicon 369 -1838 369 -1838 0 2
rlabel polysilicon 366 -1844 366 -1844 0 3
rlabel polysilicon 369 -1844 369 -1844 0 4
rlabel polysilicon 373 -1838 373 -1838 0 1
rlabel polysilicon 373 -1844 373 -1844 0 3
rlabel polysilicon 380 -1838 380 -1838 0 1
rlabel polysilicon 380 -1844 380 -1844 0 3
rlabel polysilicon 387 -1838 387 -1838 0 1
rlabel polysilicon 390 -1838 390 -1838 0 2
rlabel polysilicon 387 -1844 387 -1844 0 3
rlabel polysilicon 394 -1838 394 -1838 0 1
rlabel polysilicon 394 -1844 394 -1844 0 3
rlabel polysilicon 401 -1838 401 -1838 0 1
rlabel polysilicon 401 -1844 401 -1844 0 3
rlabel polysilicon 408 -1838 408 -1838 0 1
rlabel polysilicon 408 -1844 408 -1844 0 3
rlabel polysilicon 415 -1838 415 -1838 0 1
rlabel polysilicon 415 -1844 415 -1844 0 3
rlabel polysilicon 422 -1838 422 -1838 0 1
rlabel polysilicon 422 -1844 422 -1844 0 3
rlabel polysilicon 429 -1838 429 -1838 0 1
rlabel polysilicon 429 -1844 429 -1844 0 3
rlabel polysilicon 436 -1838 436 -1838 0 1
rlabel polysilicon 436 -1844 436 -1844 0 3
rlabel polysilicon 443 -1838 443 -1838 0 1
rlabel polysilicon 443 -1844 443 -1844 0 3
rlabel polysilicon 450 -1838 450 -1838 0 1
rlabel polysilicon 450 -1844 450 -1844 0 3
rlabel polysilicon 457 -1838 457 -1838 0 1
rlabel polysilicon 457 -1844 457 -1844 0 3
rlabel polysilicon 464 -1838 464 -1838 0 1
rlabel polysilicon 467 -1838 467 -1838 0 2
rlabel polysilicon 464 -1844 464 -1844 0 3
rlabel polysilicon 467 -1844 467 -1844 0 4
rlabel polysilicon 471 -1838 471 -1838 0 1
rlabel polysilicon 471 -1844 471 -1844 0 3
rlabel polysilicon 478 -1838 478 -1838 0 1
rlabel polysilicon 481 -1838 481 -1838 0 2
rlabel polysilicon 478 -1844 478 -1844 0 3
rlabel polysilicon 481 -1844 481 -1844 0 4
rlabel polysilicon 485 -1838 485 -1838 0 1
rlabel polysilicon 485 -1844 485 -1844 0 3
rlabel polysilicon 492 -1838 492 -1838 0 1
rlabel polysilicon 492 -1844 492 -1844 0 3
rlabel polysilicon 499 -1838 499 -1838 0 1
rlabel polysilicon 499 -1844 499 -1844 0 3
rlabel polysilicon 506 -1838 506 -1838 0 1
rlabel polysilicon 506 -1844 506 -1844 0 3
rlabel polysilicon 513 -1838 513 -1838 0 1
rlabel polysilicon 516 -1844 516 -1844 0 4
rlabel polysilicon 520 -1838 520 -1838 0 1
rlabel polysilicon 520 -1844 520 -1844 0 3
rlabel polysilicon 527 -1838 527 -1838 0 1
rlabel polysilicon 527 -1844 527 -1844 0 3
rlabel polysilicon 534 -1838 534 -1838 0 1
rlabel polysilicon 534 -1844 534 -1844 0 3
rlabel polysilicon 541 -1838 541 -1838 0 1
rlabel polysilicon 541 -1844 541 -1844 0 3
rlabel polysilicon 548 -1838 548 -1838 0 1
rlabel polysilicon 548 -1844 548 -1844 0 3
rlabel polysilicon 555 -1838 555 -1838 0 1
rlabel polysilicon 555 -1844 555 -1844 0 3
rlabel polysilicon 562 -1838 562 -1838 0 1
rlabel polysilicon 562 -1844 562 -1844 0 3
rlabel polysilicon 569 -1838 569 -1838 0 1
rlabel polysilicon 569 -1844 569 -1844 0 3
rlabel polysilicon 576 -1838 576 -1838 0 1
rlabel polysilicon 576 -1844 576 -1844 0 3
rlabel polysilicon 583 -1838 583 -1838 0 1
rlabel polysilicon 586 -1838 586 -1838 0 2
rlabel polysilicon 583 -1844 583 -1844 0 3
rlabel polysilicon 586 -1844 586 -1844 0 4
rlabel polysilicon 590 -1838 590 -1838 0 1
rlabel polysilicon 590 -1844 590 -1844 0 3
rlabel polysilicon 597 -1838 597 -1838 0 1
rlabel polysilicon 597 -1844 597 -1844 0 3
rlabel polysilicon 604 -1838 604 -1838 0 1
rlabel polysilicon 607 -1838 607 -1838 0 2
rlabel polysilicon 604 -1844 604 -1844 0 3
rlabel polysilicon 607 -1844 607 -1844 0 4
rlabel polysilicon 611 -1838 611 -1838 0 1
rlabel polysilicon 614 -1838 614 -1838 0 2
rlabel polysilicon 611 -1844 611 -1844 0 3
rlabel polysilicon 614 -1844 614 -1844 0 4
rlabel polysilicon 618 -1838 618 -1838 0 1
rlabel polysilicon 618 -1844 618 -1844 0 3
rlabel polysilicon 625 -1838 625 -1838 0 1
rlabel polysilicon 628 -1838 628 -1838 0 2
rlabel polysilicon 625 -1844 625 -1844 0 3
rlabel polysilicon 628 -1844 628 -1844 0 4
rlabel polysilicon 632 -1838 632 -1838 0 1
rlabel polysilicon 632 -1844 632 -1844 0 3
rlabel polysilicon 639 -1838 639 -1838 0 1
rlabel polysilicon 642 -1838 642 -1838 0 2
rlabel polysilicon 639 -1844 639 -1844 0 3
rlabel polysilicon 642 -1844 642 -1844 0 4
rlabel polysilicon 646 -1838 646 -1838 0 1
rlabel polysilicon 646 -1844 646 -1844 0 3
rlabel polysilicon 653 -1838 653 -1838 0 1
rlabel polysilicon 653 -1844 653 -1844 0 3
rlabel polysilicon 656 -1844 656 -1844 0 4
rlabel polysilicon 660 -1838 660 -1838 0 1
rlabel polysilicon 660 -1844 660 -1844 0 3
rlabel polysilicon 667 -1838 667 -1838 0 1
rlabel polysilicon 667 -1844 667 -1844 0 3
rlabel polysilicon 674 -1838 674 -1838 0 1
rlabel polysilicon 674 -1844 674 -1844 0 3
rlabel polysilicon 681 -1838 681 -1838 0 1
rlabel polysilicon 681 -1844 681 -1844 0 3
rlabel polysilicon 688 -1838 688 -1838 0 1
rlabel polysilicon 688 -1844 688 -1844 0 3
rlabel polysilicon 695 -1838 695 -1838 0 1
rlabel polysilicon 695 -1844 695 -1844 0 3
rlabel polysilicon 702 -1838 702 -1838 0 1
rlabel polysilicon 702 -1844 702 -1844 0 3
rlabel polysilicon 709 -1838 709 -1838 0 1
rlabel polysilicon 712 -1838 712 -1838 0 2
rlabel polysilicon 709 -1844 709 -1844 0 3
rlabel polysilicon 712 -1844 712 -1844 0 4
rlabel polysilicon 716 -1838 716 -1838 0 1
rlabel polysilicon 719 -1838 719 -1838 0 2
rlabel polysilicon 716 -1844 716 -1844 0 3
rlabel polysilicon 719 -1844 719 -1844 0 4
rlabel polysilicon 723 -1838 723 -1838 0 1
rlabel polysilicon 723 -1844 723 -1844 0 3
rlabel polysilicon 730 -1838 730 -1838 0 1
rlabel polysilicon 733 -1838 733 -1838 0 2
rlabel polysilicon 737 -1838 737 -1838 0 1
rlabel polysilicon 737 -1844 737 -1844 0 3
rlabel polysilicon 744 -1838 744 -1838 0 1
rlabel polysilicon 744 -1844 744 -1844 0 3
rlabel polysilicon 751 -1838 751 -1838 0 1
rlabel polysilicon 754 -1838 754 -1838 0 2
rlabel polysilicon 751 -1844 751 -1844 0 3
rlabel polysilicon 754 -1844 754 -1844 0 4
rlabel polysilicon 758 -1838 758 -1838 0 1
rlabel polysilicon 761 -1838 761 -1838 0 2
rlabel polysilicon 758 -1844 758 -1844 0 3
rlabel polysilicon 761 -1844 761 -1844 0 4
rlabel polysilicon 765 -1838 765 -1838 0 1
rlabel polysilicon 765 -1844 765 -1844 0 3
rlabel polysilicon 772 -1838 772 -1838 0 1
rlabel polysilicon 772 -1844 772 -1844 0 3
rlabel polysilicon 779 -1838 779 -1838 0 1
rlabel polysilicon 779 -1844 779 -1844 0 3
rlabel polysilicon 786 -1838 786 -1838 0 1
rlabel polysilicon 786 -1844 786 -1844 0 3
rlabel polysilicon 793 -1838 793 -1838 0 1
rlabel polysilicon 793 -1844 793 -1844 0 3
rlabel polysilicon 800 -1838 800 -1838 0 1
rlabel polysilicon 800 -1844 800 -1844 0 3
rlabel polysilicon 807 -1838 807 -1838 0 1
rlabel polysilicon 807 -1844 807 -1844 0 3
rlabel polysilicon 814 -1838 814 -1838 0 1
rlabel polysilicon 814 -1844 814 -1844 0 3
rlabel polysilicon 821 -1838 821 -1838 0 1
rlabel polysilicon 821 -1844 821 -1844 0 3
rlabel polysilicon 828 -1838 828 -1838 0 1
rlabel polysilicon 828 -1844 828 -1844 0 3
rlabel polysilicon 835 -1838 835 -1838 0 1
rlabel polysilicon 835 -1844 835 -1844 0 3
rlabel polysilicon 842 -1838 842 -1838 0 1
rlabel polysilicon 842 -1844 842 -1844 0 3
rlabel polysilicon 849 -1838 849 -1838 0 1
rlabel polysilicon 849 -1844 849 -1844 0 3
rlabel polysilicon 856 -1838 856 -1838 0 1
rlabel polysilicon 856 -1844 856 -1844 0 3
rlabel polysilicon 863 -1838 863 -1838 0 1
rlabel polysilicon 863 -1844 863 -1844 0 3
rlabel polysilicon 870 -1838 870 -1838 0 1
rlabel polysilicon 870 -1844 870 -1844 0 3
rlabel polysilicon 877 -1838 877 -1838 0 1
rlabel polysilicon 877 -1844 877 -1844 0 3
rlabel polysilicon 884 -1838 884 -1838 0 1
rlabel polysilicon 884 -1844 884 -1844 0 3
rlabel polysilicon 891 -1838 891 -1838 0 1
rlabel polysilicon 891 -1844 891 -1844 0 3
rlabel polysilicon 898 -1838 898 -1838 0 1
rlabel polysilicon 898 -1844 898 -1844 0 3
rlabel polysilicon 905 -1838 905 -1838 0 1
rlabel polysilicon 905 -1844 905 -1844 0 3
rlabel polysilicon 912 -1838 912 -1838 0 1
rlabel polysilicon 912 -1844 912 -1844 0 3
rlabel polysilicon 919 -1838 919 -1838 0 1
rlabel polysilicon 919 -1844 919 -1844 0 3
rlabel polysilicon 926 -1838 926 -1838 0 1
rlabel polysilicon 926 -1844 926 -1844 0 3
rlabel polysilicon 933 -1838 933 -1838 0 1
rlabel polysilicon 933 -1844 933 -1844 0 3
rlabel polysilicon 940 -1838 940 -1838 0 1
rlabel polysilicon 940 -1844 940 -1844 0 3
rlabel polysilicon 947 -1838 947 -1838 0 1
rlabel polysilicon 947 -1844 947 -1844 0 3
rlabel polysilicon 954 -1838 954 -1838 0 1
rlabel polysilicon 954 -1844 954 -1844 0 3
rlabel polysilicon 961 -1838 961 -1838 0 1
rlabel polysilicon 961 -1844 961 -1844 0 3
rlabel polysilicon 968 -1838 968 -1838 0 1
rlabel polysilicon 968 -1844 968 -1844 0 3
rlabel polysilicon 975 -1838 975 -1838 0 1
rlabel polysilicon 975 -1844 975 -1844 0 3
rlabel polysilicon 982 -1838 982 -1838 0 1
rlabel polysilicon 982 -1844 982 -1844 0 3
rlabel polysilicon 989 -1838 989 -1838 0 1
rlabel polysilicon 989 -1844 989 -1844 0 3
rlabel polysilicon 996 -1838 996 -1838 0 1
rlabel polysilicon 996 -1844 996 -1844 0 3
rlabel polysilicon 1003 -1838 1003 -1838 0 1
rlabel polysilicon 1003 -1844 1003 -1844 0 3
rlabel polysilicon 1010 -1838 1010 -1838 0 1
rlabel polysilicon 1010 -1844 1010 -1844 0 3
rlabel polysilicon 1017 -1838 1017 -1838 0 1
rlabel polysilicon 1017 -1844 1017 -1844 0 3
rlabel polysilicon 1024 -1838 1024 -1838 0 1
rlabel polysilicon 1024 -1844 1024 -1844 0 3
rlabel polysilicon 1031 -1838 1031 -1838 0 1
rlabel polysilicon 1031 -1844 1031 -1844 0 3
rlabel polysilicon 1038 -1838 1038 -1838 0 1
rlabel polysilicon 1038 -1844 1038 -1844 0 3
rlabel polysilicon 1045 -1838 1045 -1838 0 1
rlabel polysilicon 1045 -1844 1045 -1844 0 3
rlabel polysilicon 1052 -1838 1052 -1838 0 1
rlabel polysilicon 1052 -1844 1052 -1844 0 3
rlabel polysilicon 1059 -1838 1059 -1838 0 1
rlabel polysilicon 1059 -1844 1059 -1844 0 3
rlabel polysilicon 1066 -1838 1066 -1838 0 1
rlabel polysilicon 1066 -1844 1066 -1844 0 3
rlabel polysilicon 1073 -1838 1073 -1838 0 1
rlabel polysilicon 1073 -1844 1073 -1844 0 3
rlabel polysilicon 1080 -1838 1080 -1838 0 1
rlabel polysilicon 1080 -1844 1080 -1844 0 3
rlabel polysilicon 1087 -1838 1087 -1838 0 1
rlabel polysilicon 1087 -1844 1087 -1844 0 3
rlabel polysilicon 1094 -1838 1094 -1838 0 1
rlabel polysilicon 1094 -1844 1094 -1844 0 3
rlabel polysilicon 1101 -1838 1101 -1838 0 1
rlabel polysilicon 1101 -1844 1101 -1844 0 3
rlabel polysilicon 1108 -1838 1108 -1838 0 1
rlabel polysilicon 1108 -1844 1108 -1844 0 3
rlabel polysilicon 1115 -1838 1115 -1838 0 1
rlabel polysilicon 1115 -1844 1115 -1844 0 3
rlabel polysilicon 1122 -1838 1122 -1838 0 1
rlabel polysilicon 1122 -1844 1122 -1844 0 3
rlabel polysilicon 1129 -1838 1129 -1838 0 1
rlabel polysilicon 1129 -1844 1129 -1844 0 3
rlabel polysilicon 1136 -1838 1136 -1838 0 1
rlabel polysilicon 1136 -1844 1136 -1844 0 3
rlabel polysilicon 1143 -1838 1143 -1838 0 1
rlabel polysilicon 1143 -1844 1143 -1844 0 3
rlabel polysilicon 1150 -1838 1150 -1838 0 1
rlabel polysilicon 1150 -1844 1150 -1844 0 3
rlabel polysilicon 1157 -1838 1157 -1838 0 1
rlabel polysilicon 1157 -1844 1157 -1844 0 3
rlabel polysilicon 1164 -1838 1164 -1838 0 1
rlabel polysilicon 1164 -1844 1164 -1844 0 3
rlabel polysilicon 1171 -1838 1171 -1838 0 1
rlabel polysilicon 1171 -1844 1171 -1844 0 3
rlabel polysilicon 1178 -1838 1178 -1838 0 1
rlabel polysilicon 1178 -1844 1178 -1844 0 3
rlabel polysilicon 1185 -1838 1185 -1838 0 1
rlabel polysilicon 1185 -1844 1185 -1844 0 3
rlabel polysilicon 1192 -1838 1192 -1838 0 1
rlabel polysilicon 1192 -1844 1192 -1844 0 3
rlabel polysilicon 1199 -1838 1199 -1838 0 1
rlabel polysilicon 1199 -1844 1199 -1844 0 3
rlabel polysilicon 1206 -1838 1206 -1838 0 1
rlabel polysilicon 1206 -1844 1206 -1844 0 3
rlabel polysilicon 1213 -1838 1213 -1838 0 1
rlabel polysilicon 1213 -1844 1213 -1844 0 3
rlabel polysilicon 1220 -1838 1220 -1838 0 1
rlabel polysilicon 1220 -1844 1220 -1844 0 3
rlabel polysilicon 1227 -1838 1227 -1838 0 1
rlabel polysilicon 1227 -1844 1227 -1844 0 3
rlabel polysilicon 1234 -1838 1234 -1838 0 1
rlabel polysilicon 1234 -1844 1234 -1844 0 3
rlabel polysilicon 1241 -1838 1241 -1838 0 1
rlabel polysilicon 1241 -1844 1241 -1844 0 3
rlabel polysilicon 1248 -1838 1248 -1838 0 1
rlabel polysilicon 1248 -1844 1248 -1844 0 3
rlabel polysilicon 1255 -1838 1255 -1838 0 1
rlabel polysilicon 1255 -1844 1255 -1844 0 3
rlabel polysilicon 1262 -1838 1262 -1838 0 1
rlabel polysilicon 1262 -1844 1262 -1844 0 3
rlabel polysilicon 1269 -1838 1269 -1838 0 1
rlabel polysilicon 1269 -1844 1269 -1844 0 3
rlabel polysilicon 1276 -1838 1276 -1838 0 1
rlabel polysilicon 1276 -1844 1276 -1844 0 3
rlabel polysilicon 1283 -1838 1283 -1838 0 1
rlabel polysilicon 1286 -1838 1286 -1838 0 2
rlabel polysilicon 9 -1961 9 -1961 0 1
rlabel polysilicon 9 -1967 9 -1967 0 3
rlabel polysilicon 16 -1961 16 -1961 0 1
rlabel polysilicon 16 -1967 16 -1967 0 3
rlabel polysilicon 23 -1961 23 -1961 0 1
rlabel polysilicon 23 -1967 23 -1967 0 3
rlabel polysilicon 30 -1961 30 -1961 0 1
rlabel polysilicon 30 -1967 30 -1967 0 3
rlabel polysilicon 37 -1961 37 -1961 0 1
rlabel polysilicon 37 -1967 37 -1967 0 3
rlabel polysilicon 44 -1961 44 -1961 0 1
rlabel polysilicon 44 -1967 44 -1967 0 3
rlabel polysilicon 51 -1961 51 -1961 0 1
rlabel polysilicon 51 -1967 51 -1967 0 3
rlabel polysilicon 54 -1967 54 -1967 0 4
rlabel polysilicon 58 -1961 58 -1961 0 1
rlabel polysilicon 58 -1967 58 -1967 0 3
rlabel polysilicon 65 -1961 65 -1961 0 1
rlabel polysilicon 68 -1961 68 -1961 0 2
rlabel polysilicon 65 -1967 65 -1967 0 3
rlabel polysilicon 68 -1967 68 -1967 0 4
rlabel polysilicon 72 -1961 72 -1961 0 1
rlabel polysilicon 72 -1967 72 -1967 0 3
rlabel polysilicon 79 -1961 79 -1961 0 1
rlabel polysilicon 79 -1967 79 -1967 0 3
rlabel polysilicon 86 -1961 86 -1961 0 1
rlabel polysilicon 89 -1961 89 -1961 0 2
rlabel polysilicon 86 -1967 86 -1967 0 3
rlabel polysilicon 89 -1967 89 -1967 0 4
rlabel polysilicon 93 -1961 93 -1961 0 1
rlabel polysilicon 96 -1961 96 -1961 0 2
rlabel polysilicon 93 -1967 93 -1967 0 3
rlabel polysilicon 96 -1967 96 -1967 0 4
rlabel polysilicon 100 -1961 100 -1961 0 1
rlabel polysilicon 103 -1961 103 -1961 0 2
rlabel polysilicon 103 -1967 103 -1967 0 4
rlabel polysilicon 107 -1961 107 -1961 0 1
rlabel polysilicon 107 -1967 107 -1967 0 3
rlabel polysilicon 114 -1961 114 -1961 0 1
rlabel polysilicon 114 -1967 114 -1967 0 3
rlabel polysilicon 121 -1961 121 -1961 0 1
rlabel polysilicon 121 -1967 121 -1967 0 3
rlabel polysilicon 128 -1961 128 -1961 0 1
rlabel polysilicon 128 -1967 128 -1967 0 3
rlabel polysilicon 135 -1961 135 -1961 0 1
rlabel polysilicon 138 -1961 138 -1961 0 2
rlabel polysilicon 135 -1967 135 -1967 0 3
rlabel polysilicon 138 -1967 138 -1967 0 4
rlabel polysilicon 142 -1961 142 -1961 0 1
rlabel polysilicon 142 -1967 142 -1967 0 3
rlabel polysilicon 149 -1961 149 -1961 0 1
rlabel polysilicon 149 -1967 149 -1967 0 3
rlabel polysilicon 156 -1961 156 -1961 0 1
rlabel polysilicon 156 -1967 156 -1967 0 3
rlabel polysilicon 163 -1961 163 -1961 0 1
rlabel polysilicon 163 -1967 163 -1967 0 3
rlabel polysilicon 170 -1961 170 -1961 0 1
rlabel polysilicon 170 -1967 170 -1967 0 3
rlabel polysilicon 173 -1967 173 -1967 0 4
rlabel polysilicon 177 -1961 177 -1961 0 1
rlabel polysilicon 177 -1967 177 -1967 0 3
rlabel polysilicon 184 -1961 184 -1961 0 1
rlabel polysilicon 184 -1967 184 -1967 0 3
rlabel polysilicon 191 -1961 191 -1961 0 1
rlabel polysilicon 191 -1967 191 -1967 0 3
rlabel polysilicon 198 -1961 198 -1961 0 1
rlabel polysilicon 198 -1967 198 -1967 0 3
rlabel polysilicon 205 -1961 205 -1961 0 1
rlabel polysilicon 205 -1967 205 -1967 0 3
rlabel polysilicon 212 -1961 212 -1961 0 1
rlabel polysilicon 212 -1967 212 -1967 0 3
rlabel polysilicon 219 -1961 219 -1961 0 1
rlabel polysilicon 219 -1967 219 -1967 0 3
rlabel polysilicon 226 -1961 226 -1961 0 1
rlabel polysilicon 226 -1967 226 -1967 0 3
rlabel polysilicon 233 -1961 233 -1961 0 1
rlabel polysilicon 233 -1967 233 -1967 0 3
rlabel polysilicon 240 -1961 240 -1961 0 1
rlabel polysilicon 240 -1967 240 -1967 0 3
rlabel polysilicon 247 -1961 247 -1961 0 1
rlabel polysilicon 247 -1967 247 -1967 0 3
rlabel polysilicon 254 -1961 254 -1961 0 1
rlabel polysilicon 254 -1967 254 -1967 0 3
rlabel polysilicon 261 -1961 261 -1961 0 1
rlabel polysilicon 264 -1961 264 -1961 0 2
rlabel polysilicon 261 -1967 261 -1967 0 3
rlabel polysilicon 268 -1961 268 -1961 0 1
rlabel polysilicon 268 -1967 268 -1967 0 3
rlabel polysilicon 275 -1961 275 -1961 0 1
rlabel polysilicon 275 -1967 275 -1967 0 3
rlabel polysilicon 282 -1961 282 -1961 0 1
rlabel polysilicon 285 -1961 285 -1961 0 2
rlabel polysilicon 282 -1967 282 -1967 0 3
rlabel polysilicon 285 -1967 285 -1967 0 4
rlabel polysilicon 289 -1961 289 -1961 0 1
rlabel polysilicon 289 -1967 289 -1967 0 3
rlabel polysilicon 296 -1961 296 -1961 0 1
rlabel polysilicon 296 -1967 296 -1967 0 3
rlabel polysilicon 303 -1961 303 -1961 0 1
rlabel polysilicon 303 -1967 303 -1967 0 3
rlabel polysilicon 310 -1961 310 -1961 0 1
rlabel polysilicon 310 -1967 310 -1967 0 3
rlabel polysilicon 317 -1961 317 -1961 0 1
rlabel polysilicon 320 -1961 320 -1961 0 2
rlabel polysilicon 317 -1967 317 -1967 0 3
rlabel polysilicon 320 -1967 320 -1967 0 4
rlabel polysilicon 324 -1961 324 -1961 0 1
rlabel polysilicon 324 -1967 324 -1967 0 3
rlabel polysilicon 331 -1961 331 -1961 0 1
rlabel polysilicon 331 -1967 331 -1967 0 3
rlabel polysilicon 338 -1961 338 -1961 0 1
rlabel polysilicon 338 -1967 338 -1967 0 3
rlabel polysilicon 345 -1961 345 -1961 0 1
rlabel polysilicon 345 -1967 345 -1967 0 3
rlabel polysilicon 352 -1961 352 -1961 0 1
rlabel polysilicon 352 -1967 352 -1967 0 3
rlabel polysilicon 359 -1961 359 -1961 0 1
rlabel polysilicon 359 -1967 359 -1967 0 3
rlabel polysilicon 366 -1961 366 -1961 0 1
rlabel polysilicon 369 -1961 369 -1961 0 2
rlabel polysilicon 366 -1967 366 -1967 0 3
rlabel polysilicon 369 -1967 369 -1967 0 4
rlabel polysilicon 373 -1961 373 -1961 0 1
rlabel polysilicon 373 -1967 373 -1967 0 3
rlabel polysilicon 380 -1961 380 -1961 0 1
rlabel polysilicon 387 -1961 387 -1961 0 1
rlabel polysilicon 387 -1967 387 -1967 0 3
rlabel polysilicon 394 -1961 394 -1961 0 1
rlabel polysilicon 394 -1967 394 -1967 0 3
rlabel polysilicon 401 -1961 401 -1961 0 1
rlabel polysilicon 401 -1967 401 -1967 0 3
rlabel polysilicon 408 -1961 408 -1961 0 1
rlabel polysilicon 408 -1967 408 -1967 0 3
rlabel polysilicon 415 -1961 415 -1961 0 1
rlabel polysilicon 415 -1967 415 -1967 0 3
rlabel polysilicon 422 -1961 422 -1961 0 1
rlabel polysilicon 422 -1967 422 -1967 0 3
rlabel polysilicon 429 -1961 429 -1961 0 1
rlabel polysilicon 432 -1961 432 -1961 0 2
rlabel polysilicon 429 -1967 429 -1967 0 3
rlabel polysilicon 432 -1967 432 -1967 0 4
rlabel polysilicon 436 -1961 436 -1961 0 1
rlabel polysilicon 436 -1967 436 -1967 0 3
rlabel polysilicon 443 -1961 443 -1961 0 1
rlabel polysilicon 443 -1967 443 -1967 0 3
rlabel polysilicon 450 -1961 450 -1961 0 1
rlabel polysilicon 450 -1967 450 -1967 0 3
rlabel polysilicon 457 -1961 457 -1961 0 1
rlabel polysilicon 460 -1961 460 -1961 0 2
rlabel polysilicon 457 -1967 457 -1967 0 3
rlabel polysilicon 460 -1967 460 -1967 0 4
rlabel polysilicon 464 -1961 464 -1961 0 1
rlabel polysilicon 464 -1967 464 -1967 0 3
rlabel polysilicon 471 -1961 471 -1961 0 1
rlabel polysilicon 471 -1967 471 -1967 0 3
rlabel polysilicon 478 -1961 478 -1961 0 1
rlabel polysilicon 478 -1967 478 -1967 0 3
rlabel polysilicon 485 -1961 485 -1961 0 1
rlabel polysilicon 485 -1967 485 -1967 0 3
rlabel polysilicon 492 -1961 492 -1961 0 1
rlabel polysilicon 495 -1961 495 -1961 0 2
rlabel polysilicon 492 -1967 492 -1967 0 3
rlabel polysilicon 499 -1961 499 -1961 0 1
rlabel polysilicon 499 -1967 499 -1967 0 3
rlabel polysilicon 506 -1961 506 -1961 0 1
rlabel polysilicon 506 -1967 506 -1967 0 3
rlabel polysilicon 513 -1961 513 -1961 0 1
rlabel polysilicon 513 -1967 513 -1967 0 3
rlabel polysilicon 520 -1961 520 -1961 0 1
rlabel polysilicon 523 -1961 523 -1961 0 2
rlabel polysilicon 520 -1967 520 -1967 0 3
rlabel polysilicon 523 -1967 523 -1967 0 4
rlabel polysilicon 527 -1961 527 -1961 0 1
rlabel polysilicon 527 -1967 527 -1967 0 3
rlabel polysilicon 534 -1961 534 -1961 0 1
rlabel polysilicon 534 -1967 534 -1967 0 3
rlabel polysilicon 541 -1961 541 -1961 0 1
rlabel polysilicon 541 -1967 541 -1967 0 3
rlabel polysilicon 548 -1961 548 -1961 0 1
rlabel polysilicon 548 -1967 548 -1967 0 3
rlabel polysilicon 555 -1961 555 -1961 0 1
rlabel polysilicon 558 -1961 558 -1961 0 2
rlabel polysilicon 555 -1967 555 -1967 0 3
rlabel polysilicon 558 -1967 558 -1967 0 4
rlabel polysilicon 562 -1961 562 -1961 0 1
rlabel polysilicon 562 -1967 562 -1967 0 3
rlabel polysilicon 569 -1961 569 -1961 0 1
rlabel polysilicon 572 -1961 572 -1961 0 2
rlabel polysilicon 569 -1967 569 -1967 0 3
rlabel polysilicon 572 -1967 572 -1967 0 4
rlabel polysilicon 576 -1961 576 -1961 0 1
rlabel polysilicon 576 -1967 576 -1967 0 3
rlabel polysilicon 583 -1961 583 -1961 0 1
rlabel polysilicon 583 -1967 583 -1967 0 3
rlabel polysilicon 590 -1961 590 -1961 0 1
rlabel polysilicon 590 -1967 590 -1967 0 3
rlabel polysilicon 597 -1961 597 -1961 0 1
rlabel polysilicon 597 -1967 597 -1967 0 3
rlabel polysilicon 604 -1961 604 -1961 0 1
rlabel polysilicon 607 -1961 607 -1961 0 2
rlabel polysilicon 604 -1967 604 -1967 0 3
rlabel polysilicon 607 -1967 607 -1967 0 4
rlabel polysilicon 611 -1961 611 -1961 0 1
rlabel polysilicon 611 -1967 611 -1967 0 3
rlabel polysilicon 618 -1961 618 -1961 0 1
rlabel polysilicon 618 -1967 618 -1967 0 3
rlabel polysilicon 625 -1961 625 -1961 0 1
rlabel polysilicon 625 -1967 625 -1967 0 3
rlabel polysilicon 632 -1961 632 -1961 0 1
rlabel polysilicon 632 -1967 632 -1967 0 3
rlabel polysilicon 639 -1961 639 -1961 0 1
rlabel polysilicon 639 -1967 639 -1967 0 3
rlabel polysilicon 646 -1961 646 -1961 0 1
rlabel polysilicon 646 -1967 646 -1967 0 3
rlabel polysilicon 653 -1961 653 -1961 0 1
rlabel polysilicon 653 -1967 653 -1967 0 3
rlabel polysilicon 660 -1961 660 -1961 0 1
rlabel polysilicon 660 -1967 660 -1967 0 3
rlabel polysilicon 667 -1961 667 -1961 0 1
rlabel polysilicon 667 -1967 667 -1967 0 3
rlabel polysilicon 677 -1961 677 -1961 0 2
rlabel polysilicon 674 -1967 674 -1967 0 3
rlabel polysilicon 677 -1967 677 -1967 0 4
rlabel polysilicon 681 -1961 681 -1961 0 1
rlabel polysilicon 681 -1967 681 -1967 0 3
rlabel polysilicon 688 -1961 688 -1961 0 1
rlabel polysilicon 688 -1967 688 -1967 0 3
rlabel polysilicon 695 -1961 695 -1961 0 1
rlabel polysilicon 695 -1967 695 -1967 0 3
rlabel polysilicon 702 -1961 702 -1961 0 1
rlabel polysilicon 705 -1961 705 -1961 0 2
rlabel polysilicon 702 -1967 702 -1967 0 3
rlabel polysilicon 709 -1961 709 -1961 0 1
rlabel polysilicon 709 -1967 709 -1967 0 3
rlabel polysilicon 716 -1961 716 -1961 0 1
rlabel polysilicon 716 -1967 716 -1967 0 3
rlabel polysilicon 723 -1961 723 -1961 0 1
rlabel polysilicon 723 -1967 723 -1967 0 3
rlabel polysilicon 730 -1961 730 -1961 0 1
rlabel polysilicon 730 -1967 730 -1967 0 3
rlabel polysilicon 737 -1961 737 -1961 0 1
rlabel polysilicon 737 -1967 737 -1967 0 3
rlabel polysilicon 744 -1961 744 -1961 0 1
rlabel polysilicon 744 -1967 744 -1967 0 3
rlabel polysilicon 751 -1961 751 -1961 0 1
rlabel polysilicon 751 -1967 751 -1967 0 3
rlabel polysilicon 758 -1961 758 -1961 0 1
rlabel polysilicon 761 -1961 761 -1961 0 2
rlabel polysilicon 758 -1967 758 -1967 0 3
rlabel polysilicon 761 -1967 761 -1967 0 4
rlabel polysilicon 765 -1961 765 -1961 0 1
rlabel polysilicon 765 -1967 765 -1967 0 3
rlabel polysilicon 772 -1961 772 -1961 0 1
rlabel polysilicon 772 -1967 772 -1967 0 3
rlabel polysilicon 779 -1961 779 -1961 0 1
rlabel polysilicon 779 -1967 779 -1967 0 3
rlabel polysilicon 786 -1961 786 -1961 0 1
rlabel polysilicon 786 -1967 786 -1967 0 3
rlabel polysilicon 793 -1961 793 -1961 0 1
rlabel polysilicon 793 -1967 793 -1967 0 3
rlabel polysilicon 800 -1961 800 -1961 0 1
rlabel polysilicon 800 -1967 800 -1967 0 3
rlabel polysilicon 807 -1961 807 -1961 0 1
rlabel polysilicon 807 -1967 807 -1967 0 3
rlabel polysilicon 814 -1961 814 -1961 0 1
rlabel polysilicon 814 -1967 814 -1967 0 3
rlabel polysilicon 821 -1961 821 -1961 0 1
rlabel polysilicon 821 -1967 821 -1967 0 3
rlabel polysilicon 828 -1961 828 -1961 0 1
rlabel polysilicon 828 -1967 828 -1967 0 3
rlabel polysilicon 835 -1961 835 -1961 0 1
rlabel polysilicon 838 -1961 838 -1961 0 2
rlabel polysilicon 835 -1967 835 -1967 0 3
rlabel polysilicon 838 -1967 838 -1967 0 4
rlabel polysilicon 842 -1961 842 -1961 0 1
rlabel polysilicon 842 -1967 842 -1967 0 3
rlabel polysilicon 849 -1961 849 -1961 0 1
rlabel polysilicon 849 -1967 849 -1967 0 3
rlabel polysilicon 856 -1961 856 -1961 0 1
rlabel polysilicon 856 -1967 856 -1967 0 3
rlabel polysilicon 863 -1961 863 -1961 0 1
rlabel polysilicon 863 -1967 863 -1967 0 3
rlabel polysilicon 870 -1961 870 -1961 0 1
rlabel polysilicon 870 -1967 870 -1967 0 3
rlabel polysilicon 877 -1961 877 -1961 0 1
rlabel polysilicon 877 -1967 877 -1967 0 3
rlabel polysilicon 884 -1961 884 -1961 0 1
rlabel polysilicon 884 -1967 884 -1967 0 3
rlabel polysilicon 891 -1961 891 -1961 0 1
rlabel polysilicon 891 -1967 891 -1967 0 3
rlabel polysilicon 898 -1961 898 -1961 0 1
rlabel polysilicon 898 -1967 898 -1967 0 3
rlabel polysilicon 905 -1961 905 -1961 0 1
rlabel polysilicon 905 -1967 905 -1967 0 3
rlabel polysilicon 912 -1961 912 -1961 0 1
rlabel polysilicon 912 -1967 912 -1967 0 3
rlabel polysilicon 919 -1961 919 -1961 0 1
rlabel polysilicon 922 -1961 922 -1961 0 2
rlabel polysilicon 919 -1967 919 -1967 0 3
rlabel polysilicon 926 -1961 926 -1961 0 1
rlabel polysilicon 926 -1967 926 -1967 0 3
rlabel polysilicon 933 -1961 933 -1961 0 1
rlabel polysilicon 933 -1967 933 -1967 0 3
rlabel polysilicon 940 -1961 940 -1961 0 1
rlabel polysilicon 940 -1967 940 -1967 0 3
rlabel polysilicon 947 -1961 947 -1961 0 1
rlabel polysilicon 947 -1967 947 -1967 0 3
rlabel polysilicon 954 -1961 954 -1961 0 1
rlabel polysilicon 954 -1967 954 -1967 0 3
rlabel polysilicon 961 -1961 961 -1961 0 1
rlabel polysilicon 961 -1967 961 -1967 0 3
rlabel polysilicon 964 -1967 964 -1967 0 4
rlabel polysilicon 968 -1961 968 -1961 0 1
rlabel polysilicon 968 -1967 968 -1967 0 3
rlabel polysilicon 971 -1967 971 -1967 0 4
rlabel polysilicon 975 -1961 975 -1961 0 1
rlabel polysilicon 975 -1967 975 -1967 0 3
rlabel polysilicon 982 -1961 982 -1961 0 1
rlabel polysilicon 982 -1967 982 -1967 0 3
rlabel polysilicon 989 -1961 989 -1961 0 1
rlabel polysilicon 989 -1967 989 -1967 0 3
rlabel polysilicon 996 -1961 996 -1961 0 1
rlabel polysilicon 996 -1967 996 -1967 0 3
rlabel polysilicon 1003 -1961 1003 -1961 0 1
rlabel polysilicon 1003 -1967 1003 -1967 0 3
rlabel polysilicon 1010 -1961 1010 -1961 0 1
rlabel polysilicon 1010 -1967 1010 -1967 0 3
rlabel polysilicon 1017 -1961 1017 -1961 0 1
rlabel polysilicon 1017 -1967 1017 -1967 0 3
rlabel polysilicon 1024 -1961 1024 -1961 0 1
rlabel polysilicon 1024 -1967 1024 -1967 0 3
rlabel polysilicon 1031 -1961 1031 -1961 0 1
rlabel polysilicon 1031 -1967 1031 -1967 0 3
rlabel polysilicon 1038 -1961 1038 -1961 0 1
rlabel polysilicon 1038 -1967 1038 -1967 0 3
rlabel polysilicon 1045 -1961 1045 -1961 0 1
rlabel polysilicon 1045 -1967 1045 -1967 0 3
rlabel polysilicon 1052 -1961 1052 -1961 0 1
rlabel polysilicon 1052 -1967 1052 -1967 0 3
rlabel polysilicon 1059 -1961 1059 -1961 0 1
rlabel polysilicon 1059 -1967 1059 -1967 0 3
rlabel polysilicon 1066 -1961 1066 -1961 0 1
rlabel polysilicon 1066 -1967 1066 -1967 0 3
rlabel polysilicon 1073 -1961 1073 -1961 0 1
rlabel polysilicon 1073 -1967 1073 -1967 0 3
rlabel polysilicon 1080 -1961 1080 -1961 0 1
rlabel polysilicon 1080 -1967 1080 -1967 0 3
rlabel polysilicon 1087 -1961 1087 -1961 0 1
rlabel polysilicon 1087 -1967 1087 -1967 0 3
rlabel polysilicon 1094 -1961 1094 -1961 0 1
rlabel polysilicon 1094 -1967 1094 -1967 0 3
rlabel polysilicon 1101 -1961 1101 -1961 0 1
rlabel polysilicon 1101 -1967 1101 -1967 0 3
rlabel polysilicon 1108 -1961 1108 -1961 0 1
rlabel polysilicon 1108 -1967 1108 -1967 0 3
rlabel polysilicon 1115 -1961 1115 -1961 0 1
rlabel polysilicon 1115 -1967 1115 -1967 0 3
rlabel polysilicon 1122 -1961 1122 -1961 0 1
rlabel polysilicon 1122 -1967 1122 -1967 0 3
rlabel polysilicon 1129 -1961 1129 -1961 0 1
rlabel polysilicon 1129 -1967 1129 -1967 0 3
rlabel polysilicon 1136 -1961 1136 -1961 0 1
rlabel polysilicon 1136 -1967 1136 -1967 0 3
rlabel polysilicon 1143 -1961 1143 -1961 0 1
rlabel polysilicon 1143 -1967 1143 -1967 0 3
rlabel polysilicon 1150 -1961 1150 -1961 0 1
rlabel polysilicon 1150 -1967 1150 -1967 0 3
rlabel polysilicon 1157 -1961 1157 -1961 0 1
rlabel polysilicon 1157 -1967 1157 -1967 0 3
rlabel polysilicon 1164 -1961 1164 -1961 0 1
rlabel polysilicon 1164 -1967 1164 -1967 0 3
rlabel polysilicon 1171 -1961 1171 -1961 0 1
rlabel polysilicon 1171 -1967 1171 -1967 0 3
rlabel polysilicon 1178 -1961 1178 -1961 0 1
rlabel polysilicon 1178 -1967 1178 -1967 0 3
rlabel polysilicon 1185 -1961 1185 -1961 0 1
rlabel polysilicon 1185 -1967 1185 -1967 0 3
rlabel polysilicon 1192 -1961 1192 -1961 0 1
rlabel polysilicon 1192 -1967 1192 -1967 0 3
rlabel polysilicon 1199 -1961 1199 -1961 0 1
rlabel polysilicon 1199 -1967 1199 -1967 0 3
rlabel polysilicon 1206 -1961 1206 -1961 0 1
rlabel polysilicon 1206 -1967 1206 -1967 0 3
rlabel polysilicon 1213 -1961 1213 -1961 0 1
rlabel polysilicon 1213 -1967 1213 -1967 0 3
rlabel polysilicon 1223 -1961 1223 -1961 0 2
rlabel polysilicon 1220 -1967 1220 -1967 0 3
rlabel polysilicon 1223 -1967 1223 -1967 0 4
rlabel polysilicon 1227 -1961 1227 -1961 0 1
rlabel polysilicon 1227 -1967 1227 -1967 0 3
rlabel polysilicon 1234 -1961 1234 -1961 0 1
rlabel polysilicon 1234 -1967 1234 -1967 0 3
rlabel polysilicon 2 -2064 2 -2064 0 1
rlabel polysilicon 2 -2070 2 -2070 0 3
rlabel polysilicon 9 -2064 9 -2064 0 1
rlabel polysilicon 9 -2070 9 -2070 0 3
rlabel polysilicon 16 -2064 16 -2064 0 1
rlabel polysilicon 16 -2070 16 -2070 0 3
rlabel polysilicon 23 -2064 23 -2064 0 1
rlabel polysilicon 23 -2070 23 -2070 0 3
rlabel polysilicon 30 -2064 30 -2064 0 1
rlabel polysilicon 30 -2070 30 -2070 0 3
rlabel polysilicon 37 -2064 37 -2064 0 1
rlabel polysilicon 37 -2070 37 -2070 0 3
rlabel polysilicon 44 -2064 44 -2064 0 1
rlabel polysilicon 44 -2070 44 -2070 0 3
rlabel polysilicon 51 -2064 51 -2064 0 1
rlabel polysilicon 51 -2070 51 -2070 0 3
rlabel polysilicon 58 -2064 58 -2064 0 1
rlabel polysilicon 58 -2070 58 -2070 0 3
rlabel polysilicon 65 -2064 65 -2064 0 1
rlabel polysilicon 65 -2070 65 -2070 0 3
rlabel polysilicon 72 -2064 72 -2064 0 1
rlabel polysilicon 72 -2070 72 -2070 0 3
rlabel polysilicon 79 -2064 79 -2064 0 1
rlabel polysilicon 79 -2070 79 -2070 0 3
rlabel polysilicon 86 -2064 86 -2064 0 1
rlabel polysilicon 89 -2064 89 -2064 0 2
rlabel polysilicon 86 -2070 86 -2070 0 3
rlabel polysilicon 89 -2070 89 -2070 0 4
rlabel polysilicon 93 -2064 93 -2064 0 1
rlabel polysilicon 96 -2064 96 -2064 0 2
rlabel polysilicon 93 -2070 93 -2070 0 3
rlabel polysilicon 100 -2064 100 -2064 0 1
rlabel polysilicon 100 -2070 100 -2070 0 3
rlabel polysilicon 107 -2064 107 -2064 0 1
rlabel polysilicon 110 -2064 110 -2064 0 2
rlabel polysilicon 107 -2070 107 -2070 0 3
rlabel polysilicon 110 -2070 110 -2070 0 4
rlabel polysilicon 114 -2064 114 -2064 0 1
rlabel polysilicon 117 -2064 117 -2064 0 2
rlabel polysilicon 114 -2070 114 -2070 0 3
rlabel polysilicon 117 -2070 117 -2070 0 4
rlabel polysilicon 121 -2064 121 -2064 0 1
rlabel polysilicon 121 -2070 121 -2070 0 3
rlabel polysilicon 128 -2064 128 -2064 0 1
rlabel polysilicon 128 -2070 128 -2070 0 3
rlabel polysilicon 135 -2064 135 -2064 0 1
rlabel polysilicon 135 -2070 135 -2070 0 3
rlabel polysilicon 142 -2064 142 -2064 0 1
rlabel polysilicon 142 -2070 142 -2070 0 3
rlabel polysilicon 149 -2064 149 -2064 0 1
rlabel polysilicon 152 -2064 152 -2064 0 2
rlabel polysilicon 149 -2070 149 -2070 0 3
rlabel polysilicon 152 -2070 152 -2070 0 4
rlabel polysilicon 156 -2064 156 -2064 0 1
rlabel polysilicon 156 -2070 156 -2070 0 3
rlabel polysilicon 163 -2064 163 -2064 0 1
rlabel polysilicon 166 -2064 166 -2064 0 2
rlabel polysilicon 163 -2070 163 -2070 0 3
rlabel polysilicon 166 -2070 166 -2070 0 4
rlabel polysilicon 170 -2064 170 -2064 0 1
rlabel polysilicon 170 -2070 170 -2070 0 3
rlabel polysilicon 177 -2064 177 -2064 0 1
rlabel polysilicon 177 -2070 177 -2070 0 3
rlabel polysilicon 184 -2064 184 -2064 0 1
rlabel polysilicon 184 -2070 184 -2070 0 3
rlabel polysilicon 191 -2064 191 -2064 0 1
rlabel polysilicon 191 -2070 191 -2070 0 3
rlabel polysilicon 198 -2064 198 -2064 0 1
rlabel polysilicon 198 -2070 198 -2070 0 3
rlabel polysilicon 205 -2064 205 -2064 0 1
rlabel polysilicon 205 -2070 205 -2070 0 3
rlabel polysilicon 212 -2064 212 -2064 0 1
rlabel polysilicon 212 -2070 212 -2070 0 3
rlabel polysilicon 219 -2064 219 -2064 0 1
rlabel polysilicon 219 -2070 219 -2070 0 3
rlabel polysilicon 226 -2064 226 -2064 0 1
rlabel polysilicon 226 -2070 226 -2070 0 3
rlabel polysilicon 233 -2064 233 -2064 0 1
rlabel polysilicon 233 -2070 233 -2070 0 3
rlabel polysilicon 240 -2064 240 -2064 0 1
rlabel polysilicon 243 -2064 243 -2064 0 2
rlabel polysilicon 240 -2070 240 -2070 0 3
rlabel polysilicon 243 -2070 243 -2070 0 4
rlabel polysilicon 247 -2064 247 -2064 0 1
rlabel polysilicon 247 -2070 247 -2070 0 3
rlabel polysilicon 254 -2064 254 -2064 0 1
rlabel polysilicon 254 -2070 254 -2070 0 3
rlabel polysilicon 261 -2064 261 -2064 0 1
rlabel polysilicon 261 -2070 261 -2070 0 3
rlabel polysilicon 268 -2064 268 -2064 0 1
rlabel polysilicon 268 -2070 268 -2070 0 3
rlabel polysilicon 275 -2064 275 -2064 0 1
rlabel polysilicon 278 -2064 278 -2064 0 2
rlabel polysilicon 278 -2070 278 -2070 0 4
rlabel polysilicon 282 -2064 282 -2064 0 1
rlabel polysilicon 282 -2070 282 -2070 0 3
rlabel polysilicon 289 -2064 289 -2064 0 1
rlabel polysilicon 289 -2070 289 -2070 0 3
rlabel polysilicon 296 -2064 296 -2064 0 1
rlabel polysilicon 296 -2070 296 -2070 0 3
rlabel polysilicon 303 -2064 303 -2064 0 1
rlabel polysilicon 303 -2070 303 -2070 0 3
rlabel polysilicon 310 -2064 310 -2064 0 1
rlabel polysilicon 310 -2070 310 -2070 0 3
rlabel polysilicon 317 -2064 317 -2064 0 1
rlabel polysilicon 317 -2070 317 -2070 0 3
rlabel polysilicon 324 -2070 324 -2070 0 3
rlabel polysilicon 327 -2070 327 -2070 0 4
rlabel polysilicon 331 -2064 331 -2064 0 1
rlabel polysilicon 334 -2064 334 -2064 0 2
rlabel polysilicon 331 -2070 331 -2070 0 3
rlabel polysilicon 334 -2070 334 -2070 0 4
rlabel polysilicon 338 -2064 338 -2064 0 1
rlabel polysilicon 338 -2070 338 -2070 0 3
rlabel polysilicon 345 -2064 345 -2064 0 1
rlabel polysilicon 345 -2070 345 -2070 0 3
rlabel polysilicon 352 -2064 352 -2064 0 1
rlabel polysilicon 352 -2070 352 -2070 0 3
rlabel polysilicon 359 -2064 359 -2064 0 1
rlabel polysilicon 359 -2070 359 -2070 0 3
rlabel polysilicon 366 -2064 366 -2064 0 1
rlabel polysilicon 366 -2070 366 -2070 0 3
rlabel polysilicon 373 -2064 373 -2064 0 1
rlabel polysilicon 373 -2070 373 -2070 0 3
rlabel polysilicon 380 -2070 380 -2070 0 3
rlabel polysilicon 387 -2064 387 -2064 0 1
rlabel polysilicon 387 -2070 387 -2070 0 3
rlabel polysilicon 394 -2064 394 -2064 0 1
rlabel polysilicon 394 -2070 394 -2070 0 3
rlabel polysilicon 401 -2064 401 -2064 0 1
rlabel polysilicon 401 -2070 401 -2070 0 3
rlabel polysilicon 408 -2064 408 -2064 0 1
rlabel polysilicon 408 -2070 408 -2070 0 3
rlabel polysilicon 415 -2064 415 -2064 0 1
rlabel polysilicon 415 -2070 415 -2070 0 3
rlabel polysilicon 422 -2064 422 -2064 0 1
rlabel polysilicon 422 -2070 422 -2070 0 3
rlabel polysilicon 429 -2064 429 -2064 0 1
rlabel polysilicon 429 -2070 429 -2070 0 3
rlabel polysilicon 436 -2064 436 -2064 0 1
rlabel polysilicon 436 -2070 436 -2070 0 3
rlabel polysilicon 443 -2064 443 -2064 0 1
rlabel polysilicon 443 -2070 443 -2070 0 3
rlabel polysilicon 450 -2064 450 -2064 0 1
rlabel polysilicon 450 -2070 450 -2070 0 3
rlabel polysilicon 457 -2064 457 -2064 0 1
rlabel polysilicon 457 -2070 457 -2070 0 3
rlabel polysilicon 464 -2064 464 -2064 0 1
rlabel polysilicon 464 -2070 464 -2070 0 3
rlabel polysilicon 471 -2064 471 -2064 0 1
rlabel polysilicon 471 -2070 471 -2070 0 3
rlabel polysilicon 478 -2064 478 -2064 0 1
rlabel polysilicon 481 -2064 481 -2064 0 2
rlabel polysilicon 478 -2070 478 -2070 0 3
rlabel polysilicon 481 -2070 481 -2070 0 4
rlabel polysilicon 488 -2064 488 -2064 0 2
rlabel polysilicon 485 -2070 485 -2070 0 3
rlabel polysilicon 488 -2070 488 -2070 0 4
rlabel polysilicon 492 -2064 492 -2064 0 1
rlabel polysilicon 492 -2070 492 -2070 0 3
rlabel polysilicon 499 -2064 499 -2064 0 1
rlabel polysilicon 502 -2064 502 -2064 0 2
rlabel polysilicon 499 -2070 499 -2070 0 3
rlabel polysilicon 502 -2070 502 -2070 0 4
rlabel polysilicon 506 -2064 506 -2064 0 1
rlabel polysilicon 506 -2070 506 -2070 0 3
rlabel polysilicon 513 -2064 513 -2064 0 1
rlabel polysilicon 513 -2070 513 -2070 0 3
rlabel polysilicon 520 -2064 520 -2064 0 1
rlabel polysilicon 520 -2070 520 -2070 0 3
rlabel polysilicon 527 -2064 527 -2064 0 1
rlabel polysilicon 527 -2070 527 -2070 0 3
rlabel polysilicon 534 -2064 534 -2064 0 1
rlabel polysilicon 534 -2070 534 -2070 0 3
rlabel polysilicon 541 -2064 541 -2064 0 1
rlabel polysilicon 541 -2070 541 -2070 0 3
rlabel polysilicon 548 -2064 548 -2064 0 1
rlabel polysilicon 548 -2070 548 -2070 0 3
rlabel polysilicon 555 -2064 555 -2064 0 1
rlabel polysilicon 555 -2070 555 -2070 0 3
rlabel polysilicon 562 -2064 562 -2064 0 1
rlabel polysilicon 562 -2070 562 -2070 0 3
rlabel polysilicon 569 -2064 569 -2064 0 1
rlabel polysilicon 569 -2070 569 -2070 0 3
rlabel polysilicon 576 -2064 576 -2064 0 1
rlabel polysilicon 579 -2064 579 -2064 0 2
rlabel polysilicon 576 -2070 576 -2070 0 3
rlabel polysilicon 579 -2070 579 -2070 0 4
rlabel polysilicon 583 -2064 583 -2064 0 1
rlabel polysilicon 583 -2070 583 -2070 0 3
rlabel polysilicon 590 -2064 590 -2064 0 1
rlabel polysilicon 590 -2070 590 -2070 0 3
rlabel polysilicon 597 -2064 597 -2064 0 1
rlabel polysilicon 597 -2070 597 -2070 0 3
rlabel polysilicon 604 -2064 604 -2064 0 1
rlabel polysilicon 604 -2070 604 -2070 0 3
rlabel polysilicon 611 -2064 611 -2064 0 1
rlabel polysilicon 611 -2070 611 -2070 0 3
rlabel polysilicon 618 -2064 618 -2064 0 1
rlabel polysilicon 621 -2064 621 -2064 0 2
rlabel polysilicon 618 -2070 618 -2070 0 3
rlabel polysilicon 621 -2070 621 -2070 0 4
rlabel polysilicon 625 -2064 625 -2064 0 1
rlabel polysilicon 625 -2070 625 -2070 0 3
rlabel polysilicon 632 -2064 632 -2064 0 1
rlabel polysilicon 632 -2070 632 -2070 0 3
rlabel polysilicon 639 -2064 639 -2064 0 1
rlabel polysilicon 639 -2070 639 -2070 0 3
rlabel polysilicon 646 -2064 646 -2064 0 1
rlabel polysilicon 646 -2070 646 -2070 0 3
rlabel polysilicon 653 -2064 653 -2064 0 1
rlabel polysilicon 660 -2064 660 -2064 0 1
rlabel polysilicon 663 -2064 663 -2064 0 2
rlabel polysilicon 660 -2070 660 -2070 0 3
rlabel polysilicon 663 -2070 663 -2070 0 4
rlabel polysilicon 667 -2064 667 -2064 0 1
rlabel polysilicon 667 -2070 667 -2070 0 3
rlabel polysilicon 674 -2064 674 -2064 0 1
rlabel polysilicon 674 -2070 674 -2070 0 3
rlabel polysilicon 681 -2064 681 -2064 0 1
rlabel polysilicon 681 -2070 681 -2070 0 3
rlabel polysilicon 688 -2064 688 -2064 0 1
rlabel polysilicon 688 -2070 688 -2070 0 3
rlabel polysilicon 695 -2064 695 -2064 0 1
rlabel polysilicon 698 -2064 698 -2064 0 2
rlabel polysilicon 695 -2070 695 -2070 0 3
rlabel polysilicon 698 -2070 698 -2070 0 4
rlabel polysilicon 702 -2064 702 -2064 0 1
rlabel polysilicon 702 -2070 702 -2070 0 3
rlabel polysilicon 709 -2064 709 -2064 0 1
rlabel polysilicon 709 -2070 709 -2070 0 3
rlabel polysilicon 716 -2064 716 -2064 0 1
rlabel polysilicon 716 -2070 716 -2070 0 3
rlabel polysilicon 723 -2064 723 -2064 0 1
rlabel polysilicon 723 -2070 723 -2070 0 3
rlabel polysilicon 730 -2064 730 -2064 0 1
rlabel polysilicon 730 -2070 730 -2070 0 3
rlabel polysilicon 737 -2064 737 -2064 0 1
rlabel polysilicon 737 -2070 737 -2070 0 3
rlabel polysilicon 744 -2064 744 -2064 0 1
rlabel polysilicon 744 -2070 744 -2070 0 3
rlabel polysilicon 751 -2064 751 -2064 0 1
rlabel polysilicon 751 -2070 751 -2070 0 3
rlabel polysilicon 758 -2064 758 -2064 0 1
rlabel polysilicon 758 -2070 758 -2070 0 3
rlabel polysilicon 765 -2064 765 -2064 0 1
rlabel polysilicon 765 -2070 765 -2070 0 3
rlabel polysilicon 772 -2064 772 -2064 0 1
rlabel polysilicon 772 -2070 772 -2070 0 3
rlabel polysilicon 779 -2064 779 -2064 0 1
rlabel polysilicon 779 -2070 779 -2070 0 3
rlabel polysilicon 786 -2064 786 -2064 0 1
rlabel polysilicon 786 -2070 786 -2070 0 3
rlabel polysilicon 793 -2064 793 -2064 0 1
rlabel polysilicon 793 -2070 793 -2070 0 3
rlabel polysilicon 800 -2064 800 -2064 0 1
rlabel polysilicon 800 -2070 800 -2070 0 3
rlabel polysilicon 807 -2064 807 -2064 0 1
rlabel polysilicon 807 -2070 807 -2070 0 3
rlabel polysilicon 814 -2064 814 -2064 0 1
rlabel polysilicon 814 -2070 814 -2070 0 3
rlabel polysilicon 817 -2070 817 -2070 0 4
rlabel polysilicon 821 -2064 821 -2064 0 1
rlabel polysilicon 821 -2070 821 -2070 0 3
rlabel polysilicon 828 -2064 828 -2064 0 1
rlabel polysilicon 828 -2070 828 -2070 0 3
rlabel polysilicon 835 -2064 835 -2064 0 1
rlabel polysilicon 835 -2070 835 -2070 0 3
rlabel polysilicon 842 -2064 842 -2064 0 1
rlabel polysilicon 842 -2070 842 -2070 0 3
rlabel polysilicon 849 -2064 849 -2064 0 1
rlabel polysilicon 849 -2070 849 -2070 0 3
rlabel polysilicon 856 -2064 856 -2064 0 1
rlabel polysilicon 856 -2070 856 -2070 0 3
rlabel polysilicon 863 -2064 863 -2064 0 1
rlabel polysilicon 863 -2070 863 -2070 0 3
rlabel polysilicon 866 -2070 866 -2070 0 4
rlabel polysilicon 870 -2064 870 -2064 0 1
rlabel polysilicon 870 -2070 870 -2070 0 3
rlabel polysilicon 877 -2064 877 -2064 0 1
rlabel polysilicon 877 -2070 877 -2070 0 3
rlabel polysilicon 884 -2064 884 -2064 0 1
rlabel polysilicon 884 -2070 884 -2070 0 3
rlabel polysilicon 891 -2064 891 -2064 0 1
rlabel polysilicon 891 -2070 891 -2070 0 3
rlabel polysilicon 898 -2064 898 -2064 0 1
rlabel polysilicon 898 -2070 898 -2070 0 3
rlabel polysilicon 905 -2064 905 -2064 0 1
rlabel polysilicon 905 -2070 905 -2070 0 3
rlabel polysilicon 912 -2064 912 -2064 0 1
rlabel polysilicon 912 -2070 912 -2070 0 3
rlabel polysilicon 919 -2064 919 -2064 0 1
rlabel polysilicon 919 -2070 919 -2070 0 3
rlabel polysilicon 926 -2064 926 -2064 0 1
rlabel polysilicon 926 -2070 926 -2070 0 3
rlabel polysilicon 933 -2064 933 -2064 0 1
rlabel polysilicon 933 -2070 933 -2070 0 3
rlabel polysilicon 940 -2064 940 -2064 0 1
rlabel polysilicon 940 -2070 940 -2070 0 3
rlabel polysilicon 947 -2064 947 -2064 0 1
rlabel polysilicon 947 -2070 947 -2070 0 3
rlabel polysilicon 954 -2064 954 -2064 0 1
rlabel polysilicon 954 -2070 954 -2070 0 3
rlabel polysilicon 961 -2064 961 -2064 0 1
rlabel polysilicon 961 -2070 961 -2070 0 3
rlabel polysilicon 968 -2064 968 -2064 0 1
rlabel polysilicon 971 -2064 971 -2064 0 2
rlabel polysilicon 968 -2070 968 -2070 0 3
rlabel polysilicon 975 -2064 975 -2064 0 1
rlabel polysilicon 975 -2070 975 -2070 0 3
rlabel polysilicon 982 -2064 982 -2064 0 1
rlabel polysilicon 982 -2070 982 -2070 0 3
rlabel polysilicon 989 -2064 989 -2064 0 1
rlabel polysilicon 989 -2070 989 -2070 0 3
rlabel polysilicon 996 -2064 996 -2064 0 1
rlabel polysilicon 996 -2070 996 -2070 0 3
rlabel polysilicon 1003 -2064 1003 -2064 0 1
rlabel polysilicon 1003 -2070 1003 -2070 0 3
rlabel polysilicon 1010 -2064 1010 -2064 0 1
rlabel polysilicon 1010 -2070 1010 -2070 0 3
rlabel polysilicon 1017 -2064 1017 -2064 0 1
rlabel polysilicon 1017 -2070 1017 -2070 0 3
rlabel polysilicon 1024 -2064 1024 -2064 0 1
rlabel polysilicon 1027 -2064 1027 -2064 0 2
rlabel polysilicon 1031 -2064 1031 -2064 0 1
rlabel polysilicon 1031 -2070 1031 -2070 0 3
rlabel polysilicon 1038 -2064 1038 -2064 0 1
rlabel polysilicon 1038 -2070 1038 -2070 0 3
rlabel polysilicon 1045 -2064 1045 -2064 0 1
rlabel polysilicon 1045 -2070 1045 -2070 0 3
rlabel polysilicon 1052 -2064 1052 -2064 0 1
rlabel polysilicon 1052 -2070 1052 -2070 0 3
rlabel polysilicon 1059 -2064 1059 -2064 0 1
rlabel polysilicon 1059 -2070 1059 -2070 0 3
rlabel polysilicon 1066 -2064 1066 -2064 0 1
rlabel polysilicon 1066 -2070 1066 -2070 0 3
rlabel polysilicon 1073 -2064 1073 -2064 0 1
rlabel polysilicon 1073 -2070 1073 -2070 0 3
rlabel polysilicon 1080 -2064 1080 -2064 0 1
rlabel polysilicon 1080 -2070 1080 -2070 0 3
rlabel polysilicon 1087 -2064 1087 -2064 0 1
rlabel polysilicon 1087 -2070 1087 -2070 0 3
rlabel polysilicon 1094 -2064 1094 -2064 0 1
rlabel polysilicon 1094 -2070 1094 -2070 0 3
rlabel polysilicon 1101 -2064 1101 -2064 0 1
rlabel polysilicon 1101 -2070 1101 -2070 0 3
rlabel polysilicon 1108 -2064 1108 -2064 0 1
rlabel polysilicon 1108 -2070 1108 -2070 0 3
rlabel polysilicon 1115 -2064 1115 -2064 0 1
rlabel polysilicon 1115 -2070 1115 -2070 0 3
rlabel polysilicon 1122 -2064 1122 -2064 0 1
rlabel polysilicon 1122 -2070 1122 -2070 0 3
rlabel polysilicon 1129 -2064 1129 -2064 0 1
rlabel polysilicon 1129 -2070 1129 -2070 0 3
rlabel polysilicon 1136 -2064 1136 -2064 0 1
rlabel polysilicon 1136 -2070 1136 -2070 0 3
rlabel polysilicon 1139 -2070 1139 -2070 0 4
rlabel polysilicon 1143 -2064 1143 -2064 0 1
rlabel polysilicon 1143 -2070 1143 -2070 0 3
rlabel polysilicon 1150 -2064 1150 -2064 0 1
rlabel polysilicon 1150 -2070 1150 -2070 0 3
rlabel polysilicon 1157 -2064 1157 -2064 0 1
rlabel polysilicon 1157 -2070 1157 -2070 0 3
rlabel polysilicon 1185 -2064 1185 -2064 0 1
rlabel polysilicon 1185 -2070 1185 -2070 0 3
rlabel polysilicon 23 -2149 23 -2149 0 1
rlabel polysilicon 23 -2155 23 -2155 0 3
rlabel polysilicon 30 -2149 30 -2149 0 1
rlabel polysilicon 30 -2155 30 -2155 0 3
rlabel polysilicon 37 -2149 37 -2149 0 1
rlabel polysilicon 37 -2155 37 -2155 0 3
rlabel polysilicon 44 -2149 44 -2149 0 1
rlabel polysilicon 44 -2155 44 -2155 0 3
rlabel polysilicon 51 -2149 51 -2149 0 1
rlabel polysilicon 51 -2155 51 -2155 0 3
rlabel polysilicon 58 -2149 58 -2149 0 1
rlabel polysilicon 58 -2155 58 -2155 0 3
rlabel polysilicon 65 -2149 65 -2149 0 1
rlabel polysilicon 65 -2155 65 -2155 0 3
rlabel polysilicon 72 -2149 72 -2149 0 1
rlabel polysilicon 72 -2155 72 -2155 0 3
rlabel polysilicon 79 -2149 79 -2149 0 1
rlabel polysilicon 79 -2155 79 -2155 0 3
rlabel polysilicon 86 -2149 86 -2149 0 1
rlabel polysilicon 86 -2155 86 -2155 0 3
rlabel polysilicon 93 -2149 93 -2149 0 1
rlabel polysilicon 96 -2149 96 -2149 0 2
rlabel polysilicon 93 -2155 93 -2155 0 3
rlabel polysilicon 96 -2155 96 -2155 0 4
rlabel polysilicon 100 -2149 100 -2149 0 1
rlabel polysilicon 103 -2149 103 -2149 0 2
rlabel polysilicon 100 -2155 100 -2155 0 3
rlabel polysilicon 103 -2155 103 -2155 0 4
rlabel polysilicon 107 -2149 107 -2149 0 1
rlabel polysilicon 107 -2155 107 -2155 0 3
rlabel polysilicon 114 -2149 114 -2149 0 1
rlabel polysilicon 117 -2149 117 -2149 0 2
rlabel polysilicon 114 -2155 114 -2155 0 3
rlabel polysilicon 117 -2155 117 -2155 0 4
rlabel polysilicon 121 -2149 121 -2149 0 1
rlabel polysilicon 121 -2155 121 -2155 0 3
rlabel polysilicon 128 -2149 128 -2149 0 1
rlabel polysilicon 128 -2155 128 -2155 0 3
rlabel polysilicon 135 -2149 135 -2149 0 1
rlabel polysilicon 138 -2149 138 -2149 0 2
rlabel polysilicon 135 -2155 135 -2155 0 3
rlabel polysilicon 138 -2155 138 -2155 0 4
rlabel polysilicon 142 -2149 142 -2149 0 1
rlabel polysilicon 142 -2155 142 -2155 0 3
rlabel polysilicon 149 -2149 149 -2149 0 1
rlabel polysilicon 149 -2155 149 -2155 0 3
rlabel polysilicon 156 -2149 156 -2149 0 1
rlabel polysilicon 156 -2155 156 -2155 0 3
rlabel polysilicon 163 -2149 163 -2149 0 1
rlabel polysilicon 163 -2155 163 -2155 0 3
rlabel polysilicon 173 -2149 173 -2149 0 2
rlabel polysilicon 170 -2155 170 -2155 0 3
rlabel polysilicon 177 -2149 177 -2149 0 1
rlabel polysilicon 177 -2155 177 -2155 0 3
rlabel polysilicon 184 -2149 184 -2149 0 1
rlabel polysilicon 184 -2155 184 -2155 0 3
rlabel polysilicon 191 -2149 191 -2149 0 1
rlabel polysilicon 191 -2155 191 -2155 0 3
rlabel polysilicon 198 -2149 198 -2149 0 1
rlabel polysilicon 198 -2155 198 -2155 0 3
rlabel polysilicon 205 -2149 205 -2149 0 1
rlabel polysilicon 205 -2155 205 -2155 0 3
rlabel polysilicon 212 -2149 212 -2149 0 1
rlabel polysilicon 212 -2155 212 -2155 0 3
rlabel polysilicon 219 -2149 219 -2149 0 1
rlabel polysilicon 219 -2155 219 -2155 0 3
rlabel polysilicon 226 -2149 226 -2149 0 1
rlabel polysilicon 226 -2155 226 -2155 0 3
rlabel polysilicon 233 -2149 233 -2149 0 1
rlabel polysilicon 233 -2155 233 -2155 0 3
rlabel polysilicon 240 -2149 240 -2149 0 1
rlabel polysilicon 240 -2155 240 -2155 0 3
rlabel polysilicon 247 -2149 247 -2149 0 1
rlabel polysilicon 247 -2155 247 -2155 0 3
rlabel polysilicon 254 -2149 254 -2149 0 1
rlabel polysilicon 254 -2155 254 -2155 0 3
rlabel polysilicon 261 -2149 261 -2149 0 1
rlabel polysilicon 261 -2155 261 -2155 0 3
rlabel polysilicon 268 -2149 268 -2149 0 1
rlabel polysilicon 268 -2155 268 -2155 0 3
rlabel polysilicon 275 -2149 275 -2149 0 1
rlabel polysilicon 275 -2155 275 -2155 0 3
rlabel polysilicon 282 -2149 282 -2149 0 1
rlabel polysilicon 282 -2155 282 -2155 0 3
rlabel polysilicon 289 -2149 289 -2149 0 1
rlabel polysilicon 289 -2155 289 -2155 0 3
rlabel polysilicon 299 -2149 299 -2149 0 2
rlabel polysilicon 296 -2155 296 -2155 0 3
rlabel polysilicon 299 -2155 299 -2155 0 4
rlabel polysilicon 303 -2149 303 -2149 0 1
rlabel polysilicon 303 -2155 303 -2155 0 3
rlabel polysilicon 310 -2149 310 -2149 0 1
rlabel polysilicon 310 -2155 310 -2155 0 3
rlabel polysilicon 317 -2149 317 -2149 0 1
rlabel polysilicon 320 -2149 320 -2149 0 2
rlabel polysilicon 320 -2155 320 -2155 0 4
rlabel polysilicon 324 -2149 324 -2149 0 1
rlabel polysilicon 324 -2155 324 -2155 0 3
rlabel polysilicon 331 -2149 331 -2149 0 1
rlabel polysilicon 331 -2155 331 -2155 0 3
rlabel polysilicon 338 -2149 338 -2149 0 1
rlabel polysilicon 338 -2155 338 -2155 0 3
rlabel polysilicon 345 -2149 345 -2149 0 1
rlabel polysilicon 345 -2155 345 -2155 0 3
rlabel polysilicon 352 -2149 352 -2149 0 1
rlabel polysilicon 352 -2155 352 -2155 0 3
rlabel polysilicon 359 -2149 359 -2149 0 1
rlabel polysilicon 359 -2155 359 -2155 0 3
rlabel polysilicon 366 -2149 366 -2149 0 1
rlabel polysilicon 366 -2155 366 -2155 0 3
rlabel polysilicon 373 -2149 373 -2149 0 1
rlabel polysilicon 373 -2155 373 -2155 0 3
rlabel polysilicon 380 -2149 380 -2149 0 1
rlabel polysilicon 380 -2155 380 -2155 0 3
rlabel polysilicon 387 -2149 387 -2149 0 1
rlabel polysilicon 387 -2155 387 -2155 0 3
rlabel polysilicon 394 -2149 394 -2149 0 1
rlabel polysilicon 394 -2155 394 -2155 0 3
rlabel polysilicon 401 -2149 401 -2149 0 1
rlabel polysilicon 401 -2155 401 -2155 0 3
rlabel polysilicon 408 -2149 408 -2149 0 1
rlabel polysilicon 408 -2155 408 -2155 0 3
rlabel polysilicon 415 -2149 415 -2149 0 1
rlabel polysilicon 415 -2155 415 -2155 0 3
rlabel polysilicon 422 -2149 422 -2149 0 1
rlabel polysilicon 422 -2155 422 -2155 0 3
rlabel polysilicon 429 -2149 429 -2149 0 1
rlabel polysilicon 429 -2155 429 -2155 0 3
rlabel polysilicon 436 -2149 436 -2149 0 1
rlabel polysilicon 436 -2155 436 -2155 0 3
rlabel polysilicon 443 -2149 443 -2149 0 1
rlabel polysilicon 443 -2155 443 -2155 0 3
rlabel polysilicon 450 -2149 450 -2149 0 1
rlabel polysilicon 450 -2155 450 -2155 0 3
rlabel polysilicon 457 -2149 457 -2149 0 1
rlabel polysilicon 457 -2155 457 -2155 0 3
rlabel polysilicon 464 -2149 464 -2149 0 1
rlabel polysilicon 467 -2149 467 -2149 0 2
rlabel polysilicon 464 -2155 464 -2155 0 3
rlabel polysilicon 467 -2155 467 -2155 0 4
rlabel polysilicon 471 -2149 471 -2149 0 1
rlabel polysilicon 471 -2155 471 -2155 0 3
rlabel polysilicon 478 -2149 478 -2149 0 1
rlabel polysilicon 481 -2149 481 -2149 0 2
rlabel polysilicon 478 -2155 478 -2155 0 3
rlabel polysilicon 485 -2149 485 -2149 0 1
rlabel polysilicon 485 -2155 485 -2155 0 3
rlabel polysilicon 488 -2155 488 -2155 0 4
rlabel polysilicon 492 -2149 492 -2149 0 1
rlabel polysilicon 492 -2155 492 -2155 0 3
rlabel polysilicon 499 -2149 499 -2149 0 1
rlabel polysilicon 499 -2155 499 -2155 0 3
rlabel polysilicon 509 -2149 509 -2149 0 2
rlabel polysilicon 506 -2155 506 -2155 0 3
rlabel polysilicon 509 -2155 509 -2155 0 4
rlabel polysilicon 513 -2149 513 -2149 0 1
rlabel polysilicon 516 -2149 516 -2149 0 2
rlabel polysilicon 513 -2155 513 -2155 0 3
rlabel polysilicon 516 -2155 516 -2155 0 4
rlabel polysilicon 520 -2149 520 -2149 0 1
rlabel polysilicon 520 -2155 520 -2155 0 3
rlabel polysilicon 527 -2149 527 -2149 0 1
rlabel polysilicon 530 -2149 530 -2149 0 2
rlabel polysilicon 527 -2155 527 -2155 0 3
rlabel polysilicon 534 -2149 534 -2149 0 1
rlabel polysilicon 534 -2155 534 -2155 0 3
rlabel polysilicon 541 -2149 541 -2149 0 1
rlabel polysilicon 541 -2155 541 -2155 0 3
rlabel polysilicon 548 -2149 548 -2149 0 1
rlabel polysilicon 548 -2155 548 -2155 0 3
rlabel polysilicon 555 -2149 555 -2149 0 1
rlabel polysilicon 555 -2155 555 -2155 0 3
rlabel polysilicon 562 -2149 562 -2149 0 1
rlabel polysilicon 562 -2155 562 -2155 0 3
rlabel polysilicon 569 -2149 569 -2149 0 1
rlabel polysilicon 569 -2155 569 -2155 0 3
rlabel polysilicon 576 -2149 576 -2149 0 1
rlabel polysilicon 576 -2155 576 -2155 0 3
rlabel polysilicon 583 -2149 583 -2149 0 1
rlabel polysilicon 583 -2155 583 -2155 0 3
rlabel polysilicon 590 -2149 590 -2149 0 1
rlabel polysilicon 590 -2155 590 -2155 0 3
rlabel polysilicon 597 -2149 597 -2149 0 1
rlabel polysilicon 600 -2149 600 -2149 0 2
rlabel polysilicon 597 -2155 597 -2155 0 3
rlabel polysilicon 600 -2155 600 -2155 0 4
rlabel polysilicon 604 -2149 604 -2149 0 1
rlabel polysilicon 604 -2155 604 -2155 0 3
rlabel polysilicon 611 -2149 611 -2149 0 1
rlabel polysilicon 614 -2149 614 -2149 0 2
rlabel polysilicon 611 -2155 611 -2155 0 3
rlabel polysilicon 614 -2155 614 -2155 0 4
rlabel polysilicon 618 -2149 618 -2149 0 1
rlabel polysilicon 618 -2155 618 -2155 0 3
rlabel polysilicon 625 -2149 625 -2149 0 1
rlabel polysilicon 625 -2155 625 -2155 0 3
rlabel polysilicon 632 -2149 632 -2149 0 1
rlabel polysilicon 632 -2155 632 -2155 0 3
rlabel polysilicon 639 -2149 639 -2149 0 1
rlabel polysilicon 642 -2149 642 -2149 0 2
rlabel polysilicon 646 -2149 646 -2149 0 1
rlabel polysilicon 646 -2155 646 -2155 0 3
rlabel polysilicon 653 -2149 653 -2149 0 1
rlabel polysilicon 656 -2149 656 -2149 0 2
rlabel polysilicon 653 -2155 653 -2155 0 3
rlabel polysilicon 656 -2155 656 -2155 0 4
rlabel polysilicon 660 -2149 660 -2149 0 1
rlabel polysilicon 660 -2155 660 -2155 0 3
rlabel polysilicon 667 -2149 667 -2149 0 1
rlabel polysilicon 667 -2155 667 -2155 0 3
rlabel polysilicon 674 -2149 674 -2149 0 1
rlabel polysilicon 674 -2155 674 -2155 0 3
rlabel polysilicon 681 -2149 681 -2149 0 1
rlabel polysilicon 681 -2155 681 -2155 0 3
rlabel polysilicon 688 -2149 688 -2149 0 1
rlabel polysilicon 691 -2149 691 -2149 0 2
rlabel polysilicon 688 -2155 688 -2155 0 3
rlabel polysilicon 691 -2155 691 -2155 0 4
rlabel polysilicon 695 -2149 695 -2149 0 1
rlabel polysilicon 695 -2155 695 -2155 0 3
rlabel polysilicon 702 -2149 702 -2149 0 1
rlabel polysilicon 702 -2155 702 -2155 0 3
rlabel polysilicon 709 -2149 709 -2149 0 1
rlabel polysilicon 709 -2155 709 -2155 0 3
rlabel polysilicon 716 -2149 716 -2149 0 1
rlabel polysilicon 716 -2155 716 -2155 0 3
rlabel polysilicon 723 -2149 723 -2149 0 1
rlabel polysilicon 723 -2155 723 -2155 0 3
rlabel polysilicon 730 -2149 730 -2149 0 1
rlabel polysilicon 730 -2155 730 -2155 0 3
rlabel polysilicon 737 -2149 737 -2149 0 1
rlabel polysilicon 737 -2155 737 -2155 0 3
rlabel polysilicon 744 -2149 744 -2149 0 1
rlabel polysilicon 744 -2155 744 -2155 0 3
rlabel polysilicon 751 -2149 751 -2149 0 1
rlabel polysilicon 751 -2155 751 -2155 0 3
rlabel polysilicon 758 -2149 758 -2149 0 1
rlabel polysilicon 758 -2155 758 -2155 0 3
rlabel polysilicon 765 -2149 765 -2149 0 1
rlabel polysilicon 765 -2155 765 -2155 0 3
rlabel polysilicon 772 -2149 772 -2149 0 1
rlabel polysilicon 772 -2155 772 -2155 0 3
rlabel polysilicon 779 -2149 779 -2149 0 1
rlabel polysilicon 779 -2155 779 -2155 0 3
rlabel polysilicon 786 -2149 786 -2149 0 1
rlabel polysilicon 789 -2149 789 -2149 0 2
rlabel polysilicon 786 -2155 786 -2155 0 3
rlabel polysilicon 789 -2155 789 -2155 0 4
rlabel polysilicon 793 -2149 793 -2149 0 1
rlabel polysilicon 793 -2155 793 -2155 0 3
rlabel polysilicon 800 -2149 800 -2149 0 1
rlabel polysilicon 800 -2155 800 -2155 0 3
rlabel polysilicon 807 -2149 807 -2149 0 1
rlabel polysilicon 807 -2155 807 -2155 0 3
rlabel polysilicon 814 -2149 814 -2149 0 1
rlabel polysilicon 814 -2155 814 -2155 0 3
rlabel polysilicon 821 -2149 821 -2149 0 1
rlabel polysilicon 821 -2155 821 -2155 0 3
rlabel polysilicon 828 -2149 828 -2149 0 1
rlabel polysilicon 828 -2155 828 -2155 0 3
rlabel polysilicon 835 -2149 835 -2149 0 1
rlabel polysilicon 835 -2155 835 -2155 0 3
rlabel polysilicon 842 -2149 842 -2149 0 1
rlabel polysilicon 842 -2155 842 -2155 0 3
rlabel polysilicon 849 -2149 849 -2149 0 1
rlabel polysilicon 849 -2155 849 -2155 0 3
rlabel polysilicon 856 -2149 856 -2149 0 1
rlabel polysilicon 856 -2155 856 -2155 0 3
rlabel polysilicon 863 -2149 863 -2149 0 1
rlabel polysilicon 863 -2155 863 -2155 0 3
rlabel polysilicon 870 -2149 870 -2149 0 1
rlabel polysilicon 870 -2155 870 -2155 0 3
rlabel polysilicon 877 -2149 877 -2149 0 1
rlabel polysilicon 877 -2155 877 -2155 0 3
rlabel polysilicon 884 -2149 884 -2149 0 1
rlabel polysilicon 884 -2155 884 -2155 0 3
rlabel polysilicon 891 -2149 891 -2149 0 1
rlabel polysilicon 891 -2155 891 -2155 0 3
rlabel polysilicon 898 -2149 898 -2149 0 1
rlabel polysilicon 898 -2155 898 -2155 0 3
rlabel polysilicon 905 -2149 905 -2149 0 1
rlabel polysilicon 905 -2155 905 -2155 0 3
rlabel polysilicon 912 -2149 912 -2149 0 1
rlabel polysilicon 912 -2155 912 -2155 0 3
rlabel polysilicon 919 -2149 919 -2149 0 1
rlabel polysilicon 919 -2155 919 -2155 0 3
rlabel polysilicon 926 -2149 926 -2149 0 1
rlabel polysilicon 926 -2155 926 -2155 0 3
rlabel polysilicon 933 -2149 933 -2149 0 1
rlabel polysilicon 933 -2155 933 -2155 0 3
rlabel polysilicon 940 -2149 940 -2149 0 1
rlabel polysilicon 940 -2155 940 -2155 0 3
rlabel polysilicon 947 -2149 947 -2149 0 1
rlabel polysilicon 947 -2155 947 -2155 0 3
rlabel polysilicon 954 -2149 954 -2149 0 1
rlabel polysilicon 954 -2155 954 -2155 0 3
rlabel polysilicon 961 -2149 961 -2149 0 1
rlabel polysilicon 961 -2155 961 -2155 0 3
rlabel polysilicon 968 -2149 968 -2149 0 1
rlabel polysilicon 971 -2155 971 -2155 0 4
rlabel polysilicon 975 -2149 975 -2149 0 1
rlabel polysilicon 975 -2155 975 -2155 0 3
rlabel polysilicon 982 -2149 982 -2149 0 1
rlabel polysilicon 982 -2155 982 -2155 0 3
rlabel polysilicon 989 -2149 989 -2149 0 1
rlabel polysilicon 989 -2155 989 -2155 0 3
rlabel polysilicon 996 -2149 996 -2149 0 1
rlabel polysilicon 996 -2155 996 -2155 0 3
rlabel polysilicon 1003 -2149 1003 -2149 0 1
rlabel polysilicon 1003 -2155 1003 -2155 0 3
rlabel polysilicon 1010 -2149 1010 -2149 0 1
rlabel polysilicon 1010 -2155 1010 -2155 0 3
rlabel polysilicon 1017 -2149 1017 -2149 0 1
rlabel polysilicon 1017 -2155 1017 -2155 0 3
rlabel polysilicon 1024 -2149 1024 -2149 0 1
rlabel polysilicon 1024 -2155 1024 -2155 0 3
rlabel polysilicon 1031 -2149 1031 -2149 0 1
rlabel polysilicon 1031 -2155 1031 -2155 0 3
rlabel polysilicon 1038 -2149 1038 -2149 0 1
rlabel polysilicon 1038 -2155 1038 -2155 0 3
rlabel polysilicon 1045 -2149 1045 -2149 0 1
rlabel polysilicon 1045 -2155 1045 -2155 0 3
rlabel polysilicon 1052 -2149 1052 -2149 0 1
rlabel polysilicon 1052 -2155 1052 -2155 0 3
rlabel polysilicon 1059 -2149 1059 -2149 0 1
rlabel polysilicon 1059 -2155 1059 -2155 0 3
rlabel polysilicon 1066 -2149 1066 -2149 0 1
rlabel polysilicon 1066 -2155 1066 -2155 0 3
rlabel polysilicon 1101 -2149 1101 -2149 0 1
rlabel polysilicon 1104 -2149 1104 -2149 0 2
rlabel polysilicon 1101 -2155 1101 -2155 0 3
rlabel polysilicon 1104 -2155 1104 -2155 0 4
rlabel polysilicon 1108 -2149 1108 -2149 0 1
rlabel polysilicon 1108 -2155 1108 -2155 0 3
rlabel polysilicon 1122 -2149 1122 -2149 0 1
rlabel polysilicon 1122 -2155 1122 -2155 0 3
rlabel polysilicon 30 -2230 30 -2230 0 1
rlabel polysilicon 30 -2236 30 -2236 0 3
rlabel polysilicon 37 -2230 37 -2230 0 1
rlabel polysilicon 37 -2236 37 -2236 0 3
rlabel polysilicon 44 -2230 44 -2230 0 1
rlabel polysilicon 44 -2236 44 -2236 0 3
rlabel polysilicon 51 -2230 51 -2230 0 1
rlabel polysilicon 51 -2236 51 -2236 0 3
rlabel polysilicon 58 -2230 58 -2230 0 1
rlabel polysilicon 65 -2230 65 -2230 0 1
rlabel polysilicon 65 -2236 65 -2236 0 3
rlabel polysilicon 72 -2230 72 -2230 0 1
rlabel polysilicon 72 -2236 72 -2236 0 3
rlabel polysilicon 79 -2230 79 -2230 0 1
rlabel polysilicon 86 -2230 86 -2230 0 1
rlabel polysilicon 89 -2236 89 -2236 0 4
rlabel polysilicon 93 -2230 93 -2230 0 1
rlabel polysilicon 96 -2230 96 -2230 0 2
rlabel polysilicon 93 -2236 93 -2236 0 3
rlabel polysilicon 96 -2236 96 -2236 0 4
rlabel polysilicon 100 -2230 100 -2230 0 1
rlabel polysilicon 100 -2236 100 -2236 0 3
rlabel polysilicon 107 -2230 107 -2230 0 1
rlabel polysilicon 107 -2236 107 -2236 0 3
rlabel polysilicon 114 -2230 114 -2230 0 1
rlabel polysilicon 114 -2236 114 -2236 0 3
rlabel polysilicon 121 -2230 121 -2230 0 1
rlabel polysilicon 124 -2230 124 -2230 0 2
rlabel polysilicon 121 -2236 121 -2236 0 3
rlabel polysilicon 124 -2236 124 -2236 0 4
rlabel polysilicon 128 -2230 128 -2230 0 1
rlabel polysilicon 131 -2230 131 -2230 0 2
rlabel polysilicon 128 -2236 128 -2236 0 3
rlabel polysilicon 131 -2236 131 -2236 0 4
rlabel polysilicon 135 -2230 135 -2230 0 1
rlabel polysilicon 135 -2236 135 -2236 0 3
rlabel polysilicon 142 -2230 142 -2230 0 1
rlabel polysilicon 142 -2236 142 -2236 0 3
rlabel polysilicon 149 -2230 149 -2230 0 1
rlabel polysilicon 149 -2236 149 -2236 0 3
rlabel polysilicon 156 -2230 156 -2230 0 1
rlabel polysilicon 156 -2236 156 -2236 0 3
rlabel polysilicon 163 -2230 163 -2230 0 1
rlabel polysilicon 163 -2236 163 -2236 0 3
rlabel polysilicon 170 -2230 170 -2230 0 1
rlabel polysilicon 170 -2236 170 -2236 0 3
rlabel polysilicon 177 -2230 177 -2230 0 1
rlabel polysilicon 180 -2230 180 -2230 0 2
rlabel polysilicon 177 -2236 177 -2236 0 3
rlabel polysilicon 180 -2236 180 -2236 0 4
rlabel polysilicon 184 -2230 184 -2230 0 1
rlabel polysilicon 184 -2236 184 -2236 0 3
rlabel polysilicon 191 -2230 191 -2230 0 1
rlabel polysilicon 191 -2236 191 -2236 0 3
rlabel polysilicon 198 -2230 198 -2230 0 1
rlabel polysilicon 198 -2236 198 -2236 0 3
rlabel polysilicon 205 -2230 205 -2230 0 1
rlabel polysilicon 205 -2236 205 -2236 0 3
rlabel polysilicon 212 -2230 212 -2230 0 1
rlabel polysilicon 212 -2236 212 -2236 0 3
rlabel polysilicon 219 -2230 219 -2230 0 1
rlabel polysilicon 219 -2236 219 -2236 0 3
rlabel polysilicon 226 -2230 226 -2230 0 1
rlabel polysilicon 226 -2236 226 -2236 0 3
rlabel polysilicon 233 -2230 233 -2230 0 1
rlabel polysilicon 233 -2236 233 -2236 0 3
rlabel polysilicon 240 -2230 240 -2230 0 1
rlabel polysilicon 240 -2236 240 -2236 0 3
rlabel polysilicon 247 -2230 247 -2230 0 1
rlabel polysilicon 247 -2236 247 -2236 0 3
rlabel polysilicon 254 -2230 254 -2230 0 1
rlabel polysilicon 254 -2236 254 -2236 0 3
rlabel polysilicon 261 -2230 261 -2230 0 1
rlabel polysilicon 261 -2236 261 -2236 0 3
rlabel polysilicon 268 -2230 268 -2230 0 1
rlabel polysilicon 268 -2236 268 -2236 0 3
rlabel polysilicon 275 -2230 275 -2230 0 1
rlabel polysilicon 275 -2236 275 -2236 0 3
rlabel polysilicon 282 -2230 282 -2230 0 1
rlabel polysilicon 282 -2236 282 -2236 0 3
rlabel polysilicon 289 -2230 289 -2230 0 1
rlabel polysilicon 289 -2236 289 -2236 0 3
rlabel polysilicon 296 -2230 296 -2230 0 1
rlabel polysilicon 296 -2236 296 -2236 0 3
rlabel polysilicon 303 -2230 303 -2230 0 1
rlabel polysilicon 303 -2236 303 -2236 0 3
rlabel polysilicon 310 -2230 310 -2230 0 1
rlabel polysilicon 310 -2236 310 -2236 0 3
rlabel polysilicon 317 -2230 317 -2230 0 1
rlabel polysilicon 317 -2236 317 -2236 0 3
rlabel polysilicon 324 -2230 324 -2230 0 1
rlabel polysilicon 324 -2236 324 -2236 0 3
rlabel polysilicon 331 -2230 331 -2230 0 1
rlabel polysilicon 331 -2236 331 -2236 0 3
rlabel polysilicon 338 -2230 338 -2230 0 1
rlabel polysilicon 338 -2236 338 -2236 0 3
rlabel polysilicon 345 -2230 345 -2230 0 1
rlabel polysilicon 345 -2236 345 -2236 0 3
rlabel polysilicon 355 -2230 355 -2230 0 2
rlabel polysilicon 352 -2236 352 -2236 0 3
rlabel polysilicon 355 -2236 355 -2236 0 4
rlabel polysilicon 359 -2230 359 -2230 0 1
rlabel polysilicon 359 -2236 359 -2236 0 3
rlabel polysilicon 366 -2230 366 -2230 0 1
rlabel polysilicon 366 -2236 366 -2236 0 3
rlabel polysilicon 373 -2230 373 -2230 0 1
rlabel polysilicon 373 -2236 373 -2236 0 3
rlabel polysilicon 380 -2230 380 -2230 0 1
rlabel polysilicon 380 -2236 380 -2236 0 3
rlabel polysilicon 387 -2230 387 -2230 0 1
rlabel polysilicon 387 -2236 387 -2236 0 3
rlabel polysilicon 394 -2230 394 -2230 0 1
rlabel polysilicon 397 -2230 397 -2230 0 2
rlabel polysilicon 394 -2236 394 -2236 0 3
rlabel polysilicon 397 -2236 397 -2236 0 4
rlabel polysilicon 401 -2230 401 -2230 0 1
rlabel polysilicon 401 -2236 401 -2236 0 3
rlabel polysilicon 408 -2230 408 -2230 0 1
rlabel polysilicon 408 -2236 408 -2236 0 3
rlabel polysilicon 415 -2230 415 -2230 0 1
rlabel polysilicon 415 -2236 415 -2236 0 3
rlabel polysilicon 422 -2230 422 -2230 0 1
rlabel polysilicon 422 -2236 422 -2236 0 3
rlabel polysilicon 429 -2230 429 -2230 0 1
rlabel polysilicon 429 -2236 429 -2236 0 3
rlabel polysilicon 436 -2230 436 -2230 0 1
rlabel polysilicon 436 -2236 436 -2236 0 3
rlabel polysilicon 443 -2230 443 -2230 0 1
rlabel polysilicon 443 -2236 443 -2236 0 3
rlabel polysilicon 446 -2236 446 -2236 0 4
rlabel polysilicon 450 -2230 450 -2230 0 1
rlabel polysilicon 453 -2230 453 -2230 0 2
rlabel polysilicon 450 -2236 450 -2236 0 3
rlabel polysilicon 453 -2236 453 -2236 0 4
rlabel polysilicon 457 -2230 457 -2230 0 1
rlabel polysilicon 457 -2236 457 -2236 0 3
rlabel polysilicon 464 -2230 464 -2230 0 1
rlabel polysilicon 464 -2236 464 -2236 0 3
rlabel polysilicon 471 -2230 471 -2230 0 1
rlabel polysilicon 471 -2236 471 -2236 0 3
rlabel polysilicon 481 -2230 481 -2230 0 2
rlabel polysilicon 478 -2236 478 -2236 0 3
rlabel polysilicon 481 -2236 481 -2236 0 4
rlabel polysilicon 485 -2230 485 -2230 0 1
rlabel polysilicon 488 -2230 488 -2230 0 2
rlabel polysilicon 485 -2236 485 -2236 0 3
rlabel polysilicon 492 -2230 492 -2230 0 1
rlabel polysilicon 492 -2236 492 -2236 0 3
rlabel polysilicon 499 -2230 499 -2230 0 1
rlabel polysilicon 499 -2236 499 -2236 0 3
rlabel polysilicon 506 -2230 506 -2230 0 1
rlabel polysilicon 506 -2236 506 -2236 0 3
rlabel polysilicon 513 -2230 513 -2230 0 1
rlabel polysilicon 513 -2236 513 -2236 0 3
rlabel polysilicon 520 -2230 520 -2230 0 1
rlabel polysilicon 520 -2236 520 -2236 0 3
rlabel polysilicon 527 -2230 527 -2230 0 1
rlabel polysilicon 530 -2230 530 -2230 0 2
rlabel polysilicon 527 -2236 527 -2236 0 3
rlabel polysilicon 530 -2236 530 -2236 0 4
rlabel polysilicon 534 -2230 534 -2230 0 1
rlabel polysilicon 534 -2236 534 -2236 0 3
rlabel polysilicon 541 -2230 541 -2230 0 1
rlabel polysilicon 541 -2236 541 -2236 0 3
rlabel polysilicon 548 -2230 548 -2230 0 1
rlabel polysilicon 548 -2236 548 -2236 0 3
rlabel polysilicon 555 -2230 555 -2230 0 1
rlabel polysilicon 555 -2236 555 -2236 0 3
rlabel polysilicon 562 -2230 562 -2230 0 1
rlabel polysilicon 562 -2236 562 -2236 0 3
rlabel polysilicon 569 -2230 569 -2230 0 1
rlabel polysilicon 569 -2236 569 -2236 0 3
rlabel polysilicon 576 -2230 576 -2230 0 1
rlabel polysilicon 576 -2236 576 -2236 0 3
rlabel polysilicon 583 -2230 583 -2230 0 1
rlabel polysilicon 583 -2236 583 -2236 0 3
rlabel polysilicon 590 -2230 590 -2230 0 1
rlabel polysilicon 590 -2236 590 -2236 0 3
rlabel polysilicon 597 -2230 597 -2230 0 1
rlabel polysilicon 604 -2230 604 -2230 0 1
rlabel polysilicon 604 -2236 604 -2236 0 3
rlabel polysilicon 611 -2230 611 -2230 0 1
rlabel polysilicon 611 -2236 611 -2236 0 3
rlabel polysilicon 618 -2230 618 -2230 0 1
rlabel polysilicon 618 -2236 618 -2236 0 3
rlabel polysilicon 625 -2230 625 -2230 0 1
rlabel polysilicon 625 -2236 625 -2236 0 3
rlabel polysilicon 632 -2230 632 -2230 0 1
rlabel polysilicon 632 -2236 632 -2236 0 3
rlabel polysilicon 639 -2230 639 -2230 0 1
rlabel polysilicon 639 -2236 639 -2236 0 3
rlabel polysilicon 646 -2230 646 -2230 0 1
rlabel polysilicon 646 -2236 646 -2236 0 3
rlabel polysilicon 653 -2230 653 -2230 0 1
rlabel polysilicon 656 -2230 656 -2230 0 2
rlabel polysilicon 653 -2236 653 -2236 0 3
rlabel polysilicon 656 -2236 656 -2236 0 4
rlabel polysilicon 660 -2230 660 -2230 0 1
rlabel polysilicon 660 -2236 660 -2236 0 3
rlabel polysilicon 667 -2230 667 -2230 0 1
rlabel polysilicon 670 -2230 670 -2230 0 2
rlabel polysilicon 667 -2236 667 -2236 0 3
rlabel polysilicon 670 -2236 670 -2236 0 4
rlabel polysilicon 674 -2230 674 -2230 0 1
rlabel polysilicon 674 -2236 674 -2236 0 3
rlabel polysilicon 681 -2230 681 -2230 0 1
rlabel polysilicon 681 -2236 681 -2236 0 3
rlabel polysilicon 684 -2236 684 -2236 0 4
rlabel polysilicon 688 -2230 688 -2230 0 1
rlabel polysilicon 688 -2236 688 -2236 0 3
rlabel polysilicon 695 -2230 695 -2230 0 1
rlabel polysilicon 698 -2230 698 -2230 0 2
rlabel polysilicon 698 -2236 698 -2236 0 4
rlabel polysilicon 702 -2230 702 -2230 0 1
rlabel polysilicon 702 -2236 702 -2236 0 3
rlabel polysilicon 709 -2230 709 -2230 0 1
rlabel polysilicon 709 -2236 709 -2236 0 3
rlabel polysilicon 716 -2230 716 -2230 0 1
rlabel polysilicon 716 -2236 716 -2236 0 3
rlabel polysilicon 723 -2230 723 -2230 0 1
rlabel polysilicon 723 -2236 723 -2236 0 3
rlabel polysilicon 730 -2230 730 -2230 0 1
rlabel polysilicon 730 -2236 730 -2236 0 3
rlabel polysilicon 740 -2230 740 -2230 0 2
rlabel polysilicon 737 -2236 737 -2236 0 3
rlabel polysilicon 740 -2236 740 -2236 0 4
rlabel polysilicon 747 -2230 747 -2230 0 2
rlabel polysilicon 744 -2236 744 -2236 0 3
rlabel polysilicon 747 -2236 747 -2236 0 4
rlabel polysilicon 751 -2230 751 -2230 0 1
rlabel polysilicon 751 -2236 751 -2236 0 3
rlabel polysilicon 758 -2230 758 -2230 0 1
rlabel polysilicon 758 -2236 758 -2236 0 3
rlabel polysilicon 765 -2230 765 -2230 0 1
rlabel polysilicon 765 -2236 765 -2236 0 3
rlabel polysilicon 772 -2230 772 -2230 0 1
rlabel polysilicon 772 -2236 772 -2236 0 3
rlabel polysilicon 779 -2230 779 -2230 0 1
rlabel polysilicon 779 -2236 779 -2236 0 3
rlabel polysilicon 786 -2230 786 -2230 0 1
rlabel polysilicon 786 -2236 786 -2236 0 3
rlabel polysilicon 793 -2230 793 -2230 0 1
rlabel polysilicon 793 -2236 793 -2236 0 3
rlabel polysilicon 800 -2230 800 -2230 0 1
rlabel polysilicon 800 -2236 800 -2236 0 3
rlabel polysilicon 807 -2230 807 -2230 0 1
rlabel polysilicon 807 -2236 807 -2236 0 3
rlabel polysilicon 810 -2236 810 -2236 0 4
rlabel polysilicon 814 -2230 814 -2230 0 1
rlabel polysilicon 814 -2236 814 -2236 0 3
rlabel polysilicon 821 -2230 821 -2230 0 1
rlabel polysilicon 821 -2236 821 -2236 0 3
rlabel polysilicon 828 -2230 828 -2230 0 1
rlabel polysilicon 828 -2236 828 -2236 0 3
rlabel polysilicon 835 -2230 835 -2230 0 1
rlabel polysilicon 835 -2236 835 -2236 0 3
rlabel polysilicon 842 -2230 842 -2230 0 1
rlabel polysilicon 842 -2236 842 -2236 0 3
rlabel polysilicon 849 -2230 849 -2230 0 1
rlabel polysilicon 849 -2236 849 -2236 0 3
rlabel polysilicon 856 -2230 856 -2230 0 1
rlabel polysilicon 856 -2236 856 -2236 0 3
rlabel polysilicon 863 -2230 863 -2230 0 1
rlabel polysilicon 863 -2236 863 -2236 0 3
rlabel polysilicon 870 -2230 870 -2230 0 1
rlabel polysilicon 870 -2236 870 -2236 0 3
rlabel polysilicon 877 -2230 877 -2230 0 1
rlabel polysilicon 877 -2236 877 -2236 0 3
rlabel polysilicon 884 -2230 884 -2230 0 1
rlabel polysilicon 884 -2236 884 -2236 0 3
rlabel polysilicon 891 -2230 891 -2230 0 1
rlabel polysilicon 891 -2236 891 -2236 0 3
rlabel polysilicon 898 -2230 898 -2230 0 1
rlabel polysilicon 898 -2236 898 -2236 0 3
rlabel polysilicon 905 -2230 905 -2230 0 1
rlabel polysilicon 905 -2236 905 -2236 0 3
rlabel polysilicon 912 -2230 912 -2230 0 1
rlabel polysilicon 912 -2236 912 -2236 0 3
rlabel polysilicon 919 -2230 919 -2230 0 1
rlabel polysilicon 919 -2236 919 -2236 0 3
rlabel polysilicon 926 -2230 926 -2230 0 1
rlabel polysilicon 926 -2236 926 -2236 0 3
rlabel polysilicon 933 -2230 933 -2230 0 1
rlabel polysilicon 933 -2236 933 -2236 0 3
rlabel polysilicon 940 -2230 940 -2230 0 1
rlabel polysilicon 943 -2230 943 -2230 0 2
rlabel polysilicon 940 -2236 940 -2236 0 3
rlabel polysilicon 943 -2236 943 -2236 0 4
rlabel polysilicon 947 -2230 947 -2230 0 1
rlabel polysilicon 947 -2236 947 -2236 0 3
rlabel polysilicon 954 -2230 954 -2230 0 1
rlabel polysilicon 954 -2236 954 -2236 0 3
rlabel polysilicon 957 -2236 957 -2236 0 4
rlabel polysilicon 961 -2230 961 -2230 0 1
rlabel polysilicon 961 -2236 961 -2236 0 3
rlabel polysilicon 968 -2230 968 -2230 0 1
rlabel polysilicon 968 -2236 968 -2236 0 3
rlabel polysilicon 975 -2230 975 -2230 0 1
rlabel polysilicon 975 -2236 975 -2236 0 3
rlabel polysilicon 982 -2230 982 -2230 0 1
rlabel polysilicon 982 -2236 982 -2236 0 3
rlabel polysilicon 996 -2230 996 -2230 0 1
rlabel polysilicon 996 -2236 996 -2236 0 3
rlabel polysilicon 1003 -2230 1003 -2230 0 1
rlabel polysilicon 1003 -2236 1003 -2236 0 3
rlabel polysilicon 1017 -2230 1017 -2230 0 1
rlabel polysilicon 1017 -2236 1017 -2236 0 3
rlabel polysilicon 1066 -2230 1066 -2230 0 1
rlabel polysilicon 1066 -2236 1066 -2236 0 3
rlabel polysilicon 44 -2313 44 -2313 0 1
rlabel polysilicon 44 -2319 44 -2319 0 3
rlabel polysilicon 51 -2313 51 -2313 0 1
rlabel polysilicon 51 -2319 51 -2319 0 3
rlabel polysilicon 58 -2319 58 -2319 0 3
rlabel polysilicon 65 -2313 65 -2313 0 1
rlabel polysilicon 65 -2319 65 -2319 0 3
rlabel polysilicon 72 -2313 72 -2313 0 1
rlabel polysilicon 72 -2319 72 -2319 0 3
rlabel polysilicon 79 -2313 79 -2313 0 1
rlabel polysilicon 79 -2319 79 -2319 0 3
rlabel polysilicon 89 -2313 89 -2313 0 2
rlabel polysilicon 86 -2319 86 -2319 0 3
rlabel polysilicon 89 -2319 89 -2319 0 4
rlabel polysilicon 93 -2313 93 -2313 0 1
rlabel polysilicon 93 -2319 93 -2319 0 3
rlabel polysilicon 100 -2313 100 -2313 0 1
rlabel polysilicon 100 -2319 100 -2319 0 3
rlabel polysilicon 107 -2313 107 -2313 0 1
rlabel polysilicon 107 -2319 107 -2319 0 3
rlabel polysilicon 114 -2313 114 -2313 0 1
rlabel polysilicon 114 -2319 114 -2319 0 3
rlabel polysilicon 121 -2313 121 -2313 0 1
rlabel polysilicon 121 -2319 121 -2319 0 3
rlabel polysilicon 128 -2313 128 -2313 0 1
rlabel polysilicon 128 -2319 128 -2319 0 3
rlabel polysilicon 135 -2313 135 -2313 0 1
rlabel polysilicon 138 -2313 138 -2313 0 2
rlabel polysilicon 138 -2319 138 -2319 0 4
rlabel polysilicon 142 -2313 142 -2313 0 1
rlabel polysilicon 142 -2319 142 -2319 0 3
rlabel polysilicon 149 -2313 149 -2313 0 1
rlabel polysilicon 149 -2319 149 -2319 0 3
rlabel polysilicon 156 -2313 156 -2313 0 1
rlabel polysilicon 156 -2319 156 -2319 0 3
rlabel polysilicon 163 -2313 163 -2313 0 1
rlabel polysilicon 163 -2319 163 -2319 0 3
rlabel polysilicon 170 -2313 170 -2313 0 1
rlabel polysilicon 170 -2319 170 -2319 0 3
rlabel polysilicon 177 -2313 177 -2313 0 1
rlabel polysilicon 177 -2319 177 -2319 0 3
rlabel polysilicon 184 -2313 184 -2313 0 1
rlabel polysilicon 187 -2313 187 -2313 0 2
rlabel polysilicon 184 -2319 184 -2319 0 3
rlabel polysilicon 191 -2313 191 -2313 0 1
rlabel polysilicon 191 -2319 191 -2319 0 3
rlabel polysilicon 198 -2313 198 -2313 0 1
rlabel polysilicon 198 -2319 198 -2319 0 3
rlabel polysilicon 205 -2313 205 -2313 0 1
rlabel polysilicon 205 -2319 205 -2319 0 3
rlabel polysilicon 212 -2313 212 -2313 0 1
rlabel polysilicon 212 -2319 212 -2319 0 3
rlabel polysilicon 219 -2313 219 -2313 0 1
rlabel polysilicon 219 -2319 219 -2319 0 3
rlabel polysilicon 226 -2313 226 -2313 0 1
rlabel polysilicon 226 -2319 226 -2319 0 3
rlabel polysilicon 233 -2313 233 -2313 0 1
rlabel polysilicon 233 -2319 233 -2319 0 3
rlabel polysilicon 240 -2313 240 -2313 0 1
rlabel polysilicon 240 -2319 240 -2319 0 3
rlabel polysilicon 247 -2313 247 -2313 0 1
rlabel polysilicon 247 -2319 247 -2319 0 3
rlabel polysilicon 254 -2313 254 -2313 0 1
rlabel polysilicon 254 -2319 254 -2319 0 3
rlabel polysilicon 261 -2313 261 -2313 0 1
rlabel polysilicon 261 -2319 261 -2319 0 3
rlabel polysilicon 268 -2313 268 -2313 0 1
rlabel polysilicon 268 -2319 268 -2319 0 3
rlabel polysilicon 275 -2313 275 -2313 0 1
rlabel polysilicon 275 -2319 275 -2319 0 3
rlabel polysilicon 282 -2313 282 -2313 0 1
rlabel polysilicon 282 -2319 282 -2319 0 3
rlabel polysilicon 292 -2313 292 -2313 0 2
rlabel polysilicon 289 -2319 289 -2319 0 3
rlabel polysilicon 292 -2319 292 -2319 0 4
rlabel polysilicon 296 -2313 296 -2313 0 1
rlabel polysilicon 296 -2319 296 -2319 0 3
rlabel polysilicon 303 -2313 303 -2313 0 1
rlabel polysilicon 303 -2319 303 -2319 0 3
rlabel polysilicon 310 -2313 310 -2313 0 1
rlabel polysilicon 310 -2319 310 -2319 0 3
rlabel polysilicon 317 -2313 317 -2313 0 1
rlabel polysilicon 317 -2319 317 -2319 0 3
rlabel polysilicon 324 -2313 324 -2313 0 1
rlabel polysilicon 324 -2319 324 -2319 0 3
rlabel polysilicon 331 -2313 331 -2313 0 1
rlabel polysilicon 331 -2319 331 -2319 0 3
rlabel polysilicon 338 -2313 338 -2313 0 1
rlabel polysilicon 338 -2319 338 -2319 0 3
rlabel polysilicon 345 -2313 345 -2313 0 1
rlabel polysilicon 348 -2313 348 -2313 0 2
rlabel polysilicon 345 -2319 345 -2319 0 3
rlabel polysilicon 348 -2319 348 -2319 0 4
rlabel polysilicon 352 -2313 352 -2313 0 1
rlabel polysilicon 352 -2319 352 -2319 0 3
rlabel polysilicon 359 -2313 359 -2313 0 1
rlabel polysilicon 359 -2319 359 -2319 0 3
rlabel polysilicon 366 -2313 366 -2313 0 1
rlabel polysilicon 366 -2319 366 -2319 0 3
rlabel polysilicon 373 -2313 373 -2313 0 1
rlabel polysilicon 376 -2313 376 -2313 0 2
rlabel polysilicon 373 -2319 373 -2319 0 3
rlabel polysilicon 376 -2319 376 -2319 0 4
rlabel polysilicon 380 -2313 380 -2313 0 1
rlabel polysilicon 380 -2319 380 -2319 0 3
rlabel polysilicon 387 -2313 387 -2313 0 1
rlabel polysilicon 387 -2319 387 -2319 0 3
rlabel polysilicon 394 -2313 394 -2313 0 1
rlabel polysilicon 394 -2319 394 -2319 0 3
rlabel polysilicon 401 -2313 401 -2313 0 1
rlabel polysilicon 401 -2319 401 -2319 0 3
rlabel polysilicon 408 -2313 408 -2313 0 1
rlabel polysilicon 408 -2319 408 -2319 0 3
rlabel polysilicon 415 -2313 415 -2313 0 1
rlabel polysilicon 415 -2319 415 -2319 0 3
rlabel polysilicon 422 -2313 422 -2313 0 1
rlabel polysilicon 422 -2319 422 -2319 0 3
rlabel polysilicon 425 -2319 425 -2319 0 4
rlabel polysilicon 429 -2313 429 -2313 0 1
rlabel polysilicon 429 -2319 429 -2319 0 3
rlabel polysilicon 436 -2313 436 -2313 0 1
rlabel polysilicon 436 -2319 436 -2319 0 3
rlabel polysilicon 443 -2313 443 -2313 0 1
rlabel polysilicon 446 -2313 446 -2313 0 2
rlabel polysilicon 443 -2319 443 -2319 0 3
rlabel polysilicon 446 -2319 446 -2319 0 4
rlabel polysilicon 453 -2313 453 -2313 0 2
rlabel polysilicon 450 -2319 450 -2319 0 3
rlabel polysilicon 453 -2319 453 -2319 0 4
rlabel polysilicon 457 -2313 457 -2313 0 1
rlabel polysilicon 457 -2319 457 -2319 0 3
rlabel polysilicon 464 -2313 464 -2313 0 1
rlabel polysilicon 464 -2319 464 -2319 0 3
rlabel polysilicon 471 -2313 471 -2313 0 1
rlabel polysilicon 471 -2319 471 -2319 0 3
rlabel polysilicon 478 -2313 478 -2313 0 1
rlabel polysilicon 478 -2319 478 -2319 0 3
rlabel polysilicon 485 -2313 485 -2313 0 1
rlabel polysilicon 485 -2319 485 -2319 0 3
rlabel polysilicon 492 -2313 492 -2313 0 1
rlabel polysilicon 492 -2319 492 -2319 0 3
rlabel polysilicon 495 -2319 495 -2319 0 4
rlabel polysilicon 499 -2313 499 -2313 0 1
rlabel polysilicon 499 -2319 499 -2319 0 3
rlabel polysilicon 506 -2313 506 -2313 0 1
rlabel polysilicon 506 -2319 506 -2319 0 3
rlabel polysilicon 513 -2313 513 -2313 0 1
rlabel polysilicon 513 -2319 513 -2319 0 3
rlabel polysilicon 520 -2313 520 -2313 0 1
rlabel polysilicon 520 -2319 520 -2319 0 3
rlabel polysilicon 527 -2313 527 -2313 0 1
rlabel polysilicon 527 -2319 527 -2319 0 3
rlabel polysilicon 534 -2313 534 -2313 0 1
rlabel polysilicon 537 -2313 537 -2313 0 2
rlabel polysilicon 534 -2319 534 -2319 0 3
rlabel polysilicon 541 -2313 541 -2313 0 1
rlabel polysilicon 541 -2319 541 -2319 0 3
rlabel polysilicon 548 -2313 548 -2313 0 1
rlabel polysilicon 548 -2319 548 -2319 0 3
rlabel polysilicon 555 -2313 555 -2313 0 1
rlabel polysilicon 555 -2319 555 -2319 0 3
rlabel polysilicon 562 -2313 562 -2313 0 1
rlabel polysilicon 565 -2313 565 -2313 0 2
rlabel polysilicon 562 -2319 562 -2319 0 3
rlabel polysilicon 565 -2319 565 -2319 0 4
rlabel polysilicon 569 -2313 569 -2313 0 1
rlabel polysilicon 572 -2313 572 -2313 0 2
rlabel polysilicon 569 -2319 569 -2319 0 3
rlabel polysilicon 572 -2319 572 -2319 0 4
rlabel polysilicon 576 -2313 576 -2313 0 1
rlabel polysilicon 579 -2313 579 -2313 0 2
rlabel polysilicon 576 -2319 576 -2319 0 3
rlabel polysilicon 583 -2313 583 -2313 0 1
rlabel polysilicon 583 -2319 583 -2319 0 3
rlabel polysilicon 590 -2313 590 -2313 0 1
rlabel polysilicon 590 -2319 590 -2319 0 3
rlabel polysilicon 597 -2319 597 -2319 0 3
rlabel polysilicon 604 -2313 604 -2313 0 1
rlabel polysilicon 604 -2319 604 -2319 0 3
rlabel polysilicon 611 -2313 611 -2313 0 1
rlabel polysilicon 611 -2319 611 -2319 0 3
rlabel polysilicon 618 -2313 618 -2313 0 1
rlabel polysilicon 621 -2313 621 -2313 0 2
rlabel polysilicon 618 -2319 618 -2319 0 3
rlabel polysilicon 621 -2319 621 -2319 0 4
rlabel polysilicon 625 -2313 625 -2313 0 1
rlabel polysilicon 625 -2319 625 -2319 0 3
rlabel polysilicon 632 -2313 632 -2313 0 1
rlabel polysilicon 632 -2319 632 -2319 0 3
rlabel polysilicon 639 -2313 639 -2313 0 1
rlabel polysilicon 639 -2319 639 -2319 0 3
rlabel polysilicon 646 -2313 646 -2313 0 1
rlabel polysilicon 653 -2313 653 -2313 0 1
rlabel polysilicon 656 -2313 656 -2313 0 2
rlabel polysilicon 653 -2319 653 -2319 0 3
rlabel polysilicon 656 -2319 656 -2319 0 4
rlabel polysilicon 660 -2313 660 -2313 0 1
rlabel polysilicon 660 -2319 660 -2319 0 3
rlabel polysilicon 667 -2313 667 -2313 0 1
rlabel polysilicon 667 -2319 667 -2319 0 3
rlabel polysilicon 674 -2313 674 -2313 0 1
rlabel polysilicon 674 -2319 674 -2319 0 3
rlabel polysilicon 681 -2313 681 -2313 0 1
rlabel polysilicon 684 -2313 684 -2313 0 2
rlabel polysilicon 681 -2319 681 -2319 0 3
rlabel polysilicon 688 -2313 688 -2313 0 1
rlabel polysilicon 688 -2319 688 -2319 0 3
rlabel polysilicon 695 -2313 695 -2313 0 1
rlabel polysilicon 695 -2319 695 -2319 0 3
rlabel polysilicon 702 -2313 702 -2313 0 1
rlabel polysilicon 702 -2319 702 -2319 0 3
rlabel polysilicon 709 -2313 709 -2313 0 1
rlabel polysilicon 709 -2319 709 -2319 0 3
rlabel polysilicon 716 -2313 716 -2313 0 1
rlabel polysilicon 716 -2319 716 -2319 0 3
rlabel polysilicon 719 -2319 719 -2319 0 4
rlabel polysilicon 723 -2313 723 -2313 0 1
rlabel polysilicon 723 -2319 723 -2319 0 3
rlabel polysilicon 730 -2313 730 -2313 0 1
rlabel polysilicon 730 -2319 730 -2319 0 3
rlabel polysilicon 737 -2313 737 -2313 0 1
rlabel polysilicon 737 -2319 737 -2319 0 3
rlabel polysilicon 744 -2313 744 -2313 0 1
rlabel polysilicon 744 -2319 744 -2319 0 3
rlabel polysilicon 751 -2313 751 -2313 0 1
rlabel polysilicon 751 -2319 751 -2319 0 3
rlabel polysilicon 758 -2313 758 -2313 0 1
rlabel polysilicon 758 -2319 758 -2319 0 3
rlabel polysilicon 765 -2313 765 -2313 0 1
rlabel polysilicon 765 -2319 765 -2319 0 3
rlabel polysilicon 772 -2313 772 -2313 0 1
rlabel polysilicon 772 -2319 772 -2319 0 3
rlabel polysilicon 779 -2313 779 -2313 0 1
rlabel polysilicon 779 -2319 779 -2319 0 3
rlabel polysilicon 786 -2313 786 -2313 0 1
rlabel polysilicon 786 -2319 786 -2319 0 3
rlabel polysilicon 793 -2313 793 -2313 0 1
rlabel polysilicon 793 -2319 793 -2319 0 3
rlabel polysilicon 800 -2313 800 -2313 0 1
rlabel polysilicon 803 -2313 803 -2313 0 2
rlabel polysilicon 803 -2319 803 -2319 0 4
rlabel polysilicon 807 -2313 807 -2313 0 1
rlabel polysilicon 810 -2313 810 -2313 0 2
rlabel polysilicon 807 -2319 807 -2319 0 3
rlabel polysilicon 814 -2313 814 -2313 0 1
rlabel polysilicon 814 -2319 814 -2319 0 3
rlabel polysilicon 821 -2313 821 -2313 0 1
rlabel polysilicon 821 -2319 821 -2319 0 3
rlabel polysilicon 828 -2313 828 -2313 0 1
rlabel polysilicon 828 -2319 828 -2319 0 3
rlabel polysilicon 835 -2313 835 -2313 0 1
rlabel polysilicon 835 -2319 835 -2319 0 3
rlabel polysilicon 842 -2313 842 -2313 0 1
rlabel polysilicon 842 -2319 842 -2319 0 3
rlabel polysilicon 849 -2313 849 -2313 0 1
rlabel polysilicon 849 -2319 849 -2319 0 3
rlabel polysilicon 856 -2313 856 -2313 0 1
rlabel polysilicon 856 -2319 856 -2319 0 3
rlabel polysilicon 863 -2313 863 -2313 0 1
rlabel polysilicon 863 -2319 863 -2319 0 3
rlabel polysilicon 870 -2313 870 -2313 0 1
rlabel polysilicon 870 -2319 870 -2319 0 3
rlabel polysilicon 877 -2313 877 -2313 0 1
rlabel polysilicon 877 -2319 877 -2319 0 3
rlabel polysilicon 884 -2313 884 -2313 0 1
rlabel polysilicon 884 -2319 884 -2319 0 3
rlabel polysilicon 891 -2313 891 -2313 0 1
rlabel polysilicon 891 -2319 891 -2319 0 3
rlabel polysilicon 898 -2313 898 -2313 0 1
rlabel polysilicon 898 -2319 898 -2319 0 3
rlabel polysilicon 968 -2313 968 -2313 0 1
rlabel polysilicon 968 -2319 968 -2319 0 3
rlabel polysilicon 989 -2313 989 -2313 0 1
rlabel polysilicon 989 -2319 989 -2319 0 3
rlabel polysilicon 996 -2313 996 -2313 0 1
rlabel polysilicon 996 -2319 996 -2319 0 3
rlabel polysilicon 1038 -2313 1038 -2313 0 1
rlabel polysilicon 1038 -2319 1038 -2319 0 3
rlabel polysilicon 1059 -2313 1059 -2313 0 1
rlabel polysilicon 1059 -2319 1059 -2319 0 3
rlabel polysilicon 72 -2378 72 -2378 0 1
rlabel polysilicon 72 -2384 72 -2384 0 3
rlabel polysilicon 79 -2378 79 -2378 0 1
rlabel polysilicon 79 -2384 79 -2384 0 3
rlabel polysilicon 86 -2378 86 -2378 0 1
rlabel polysilicon 86 -2384 86 -2384 0 3
rlabel polysilicon 93 -2378 93 -2378 0 1
rlabel polysilicon 93 -2384 93 -2384 0 3
rlabel polysilicon 100 -2378 100 -2378 0 1
rlabel polysilicon 100 -2384 100 -2384 0 3
rlabel polysilicon 107 -2378 107 -2378 0 1
rlabel polysilicon 107 -2384 107 -2384 0 3
rlabel polysilicon 114 -2378 114 -2378 0 1
rlabel polysilicon 114 -2384 114 -2384 0 3
rlabel polysilicon 121 -2378 121 -2378 0 1
rlabel polysilicon 121 -2384 121 -2384 0 3
rlabel polysilicon 128 -2378 128 -2378 0 1
rlabel polysilicon 128 -2384 128 -2384 0 3
rlabel polysilicon 135 -2378 135 -2378 0 1
rlabel polysilicon 135 -2384 135 -2384 0 3
rlabel polysilicon 142 -2378 142 -2378 0 1
rlabel polysilicon 142 -2384 142 -2384 0 3
rlabel polysilicon 149 -2378 149 -2378 0 1
rlabel polysilicon 152 -2378 152 -2378 0 2
rlabel polysilicon 149 -2384 149 -2384 0 3
rlabel polysilicon 156 -2378 156 -2378 0 1
rlabel polysilicon 156 -2384 156 -2384 0 3
rlabel polysilicon 163 -2378 163 -2378 0 1
rlabel polysilicon 163 -2384 163 -2384 0 3
rlabel polysilicon 166 -2384 166 -2384 0 4
rlabel polysilicon 170 -2378 170 -2378 0 1
rlabel polysilicon 173 -2384 173 -2384 0 4
rlabel polysilicon 177 -2384 177 -2384 0 3
rlabel polysilicon 184 -2378 184 -2378 0 1
rlabel polysilicon 187 -2378 187 -2378 0 2
rlabel polysilicon 184 -2384 184 -2384 0 3
rlabel polysilicon 187 -2384 187 -2384 0 4
rlabel polysilicon 191 -2378 191 -2378 0 1
rlabel polysilicon 191 -2384 191 -2384 0 3
rlabel polysilicon 198 -2378 198 -2378 0 1
rlabel polysilicon 198 -2384 198 -2384 0 3
rlabel polysilicon 205 -2378 205 -2378 0 1
rlabel polysilicon 205 -2384 205 -2384 0 3
rlabel polysilicon 212 -2378 212 -2378 0 1
rlabel polysilicon 212 -2384 212 -2384 0 3
rlabel polysilicon 219 -2378 219 -2378 0 1
rlabel polysilicon 219 -2384 219 -2384 0 3
rlabel polysilicon 226 -2378 226 -2378 0 1
rlabel polysilicon 226 -2384 226 -2384 0 3
rlabel polysilicon 233 -2378 233 -2378 0 1
rlabel polysilicon 236 -2378 236 -2378 0 2
rlabel polysilicon 233 -2384 233 -2384 0 3
rlabel polysilicon 236 -2384 236 -2384 0 4
rlabel polysilicon 240 -2378 240 -2378 0 1
rlabel polysilicon 240 -2384 240 -2384 0 3
rlabel polysilicon 247 -2378 247 -2378 0 1
rlabel polysilicon 247 -2384 247 -2384 0 3
rlabel polysilicon 254 -2378 254 -2378 0 1
rlabel polysilicon 254 -2384 254 -2384 0 3
rlabel polysilicon 261 -2378 261 -2378 0 1
rlabel polysilicon 261 -2384 261 -2384 0 3
rlabel polysilicon 271 -2378 271 -2378 0 2
rlabel polysilicon 268 -2384 268 -2384 0 3
rlabel polysilicon 275 -2378 275 -2378 0 1
rlabel polysilicon 275 -2384 275 -2384 0 3
rlabel polysilicon 282 -2378 282 -2378 0 1
rlabel polysilicon 282 -2384 282 -2384 0 3
rlabel polysilicon 289 -2378 289 -2378 0 1
rlabel polysilicon 289 -2384 289 -2384 0 3
rlabel polysilicon 296 -2378 296 -2378 0 1
rlabel polysilicon 296 -2384 296 -2384 0 3
rlabel polysilicon 303 -2378 303 -2378 0 1
rlabel polysilicon 306 -2378 306 -2378 0 2
rlabel polysilicon 303 -2384 303 -2384 0 3
rlabel polysilicon 306 -2384 306 -2384 0 4
rlabel polysilicon 310 -2378 310 -2378 0 1
rlabel polysilicon 310 -2384 310 -2384 0 3
rlabel polysilicon 317 -2378 317 -2378 0 1
rlabel polysilicon 317 -2384 317 -2384 0 3
rlabel polysilicon 324 -2378 324 -2378 0 1
rlabel polysilicon 324 -2384 324 -2384 0 3
rlabel polysilicon 331 -2378 331 -2378 0 1
rlabel polysilicon 331 -2384 331 -2384 0 3
rlabel polysilicon 338 -2378 338 -2378 0 1
rlabel polysilicon 338 -2384 338 -2384 0 3
rlabel polysilicon 345 -2378 345 -2378 0 1
rlabel polysilicon 345 -2384 345 -2384 0 3
rlabel polysilicon 352 -2378 352 -2378 0 1
rlabel polysilicon 352 -2384 352 -2384 0 3
rlabel polysilicon 359 -2378 359 -2378 0 1
rlabel polysilicon 359 -2384 359 -2384 0 3
rlabel polysilicon 366 -2378 366 -2378 0 1
rlabel polysilicon 366 -2384 366 -2384 0 3
rlabel polysilicon 373 -2378 373 -2378 0 1
rlabel polysilicon 373 -2384 373 -2384 0 3
rlabel polysilicon 383 -2378 383 -2378 0 2
rlabel polysilicon 380 -2384 380 -2384 0 3
rlabel polysilicon 383 -2384 383 -2384 0 4
rlabel polysilicon 387 -2378 387 -2378 0 1
rlabel polysilicon 387 -2384 387 -2384 0 3
rlabel polysilicon 394 -2378 394 -2378 0 1
rlabel polysilicon 394 -2384 394 -2384 0 3
rlabel polysilicon 401 -2378 401 -2378 0 1
rlabel polysilicon 401 -2384 401 -2384 0 3
rlabel polysilicon 408 -2378 408 -2378 0 1
rlabel polysilicon 408 -2384 408 -2384 0 3
rlabel polysilicon 415 -2378 415 -2378 0 1
rlabel polysilicon 415 -2384 415 -2384 0 3
rlabel polysilicon 422 -2378 422 -2378 0 1
rlabel polysilicon 422 -2384 422 -2384 0 3
rlabel polysilicon 429 -2378 429 -2378 0 1
rlabel polysilicon 429 -2384 429 -2384 0 3
rlabel polysilicon 436 -2378 436 -2378 0 1
rlabel polysilicon 436 -2384 436 -2384 0 3
rlabel polysilicon 443 -2378 443 -2378 0 1
rlabel polysilicon 443 -2384 443 -2384 0 3
rlabel polysilicon 450 -2378 450 -2378 0 1
rlabel polysilicon 450 -2384 450 -2384 0 3
rlabel polysilicon 453 -2384 453 -2384 0 4
rlabel polysilicon 457 -2378 457 -2378 0 1
rlabel polysilicon 457 -2384 457 -2384 0 3
rlabel polysilicon 464 -2378 464 -2378 0 1
rlabel polysilicon 464 -2384 464 -2384 0 3
rlabel polysilicon 471 -2378 471 -2378 0 1
rlabel polysilicon 471 -2384 471 -2384 0 3
rlabel polysilicon 478 -2378 478 -2378 0 1
rlabel polysilicon 478 -2384 478 -2384 0 3
rlabel polysilicon 485 -2378 485 -2378 0 1
rlabel polysilicon 485 -2384 485 -2384 0 3
rlabel polysilicon 492 -2378 492 -2378 0 1
rlabel polysilicon 492 -2384 492 -2384 0 3
rlabel polysilicon 499 -2378 499 -2378 0 1
rlabel polysilicon 499 -2384 499 -2384 0 3
rlabel polysilicon 506 -2378 506 -2378 0 1
rlabel polysilicon 506 -2384 506 -2384 0 3
rlabel polysilicon 513 -2378 513 -2378 0 1
rlabel polysilicon 516 -2378 516 -2378 0 2
rlabel polysilicon 513 -2384 513 -2384 0 3
rlabel polysilicon 516 -2384 516 -2384 0 4
rlabel polysilicon 520 -2378 520 -2378 0 1
rlabel polysilicon 520 -2384 520 -2384 0 3
rlabel polysilicon 527 -2378 527 -2378 0 1
rlabel polysilicon 530 -2378 530 -2378 0 2
rlabel polysilicon 530 -2384 530 -2384 0 4
rlabel polysilicon 534 -2378 534 -2378 0 1
rlabel polysilicon 534 -2384 534 -2384 0 3
rlabel polysilicon 541 -2378 541 -2378 0 1
rlabel polysilicon 541 -2384 541 -2384 0 3
rlabel polysilicon 548 -2378 548 -2378 0 1
rlabel polysilicon 548 -2384 548 -2384 0 3
rlabel polysilicon 555 -2378 555 -2378 0 1
rlabel polysilicon 558 -2378 558 -2378 0 2
rlabel polysilicon 555 -2384 555 -2384 0 3
rlabel polysilicon 558 -2384 558 -2384 0 4
rlabel polysilicon 562 -2378 562 -2378 0 1
rlabel polysilicon 562 -2384 562 -2384 0 3
rlabel polysilicon 569 -2378 569 -2378 0 1
rlabel polysilicon 569 -2384 569 -2384 0 3
rlabel polysilicon 576 -2378 576 -2378 0 1
rlabel polysilicon 576 -2384 576 -2384 0 3
rlabel polysilicon 583 -2378 583 -2378 0 1
rlabel polysilicon 583 -2384 583 -2384 0 3
rlabel polysilicon 590 -2378 590 -2378 0 1
rlabel polysilicon 590 -2384 590 -2384 0 3
rlabel polysilicon 597 -2378 597 -2378 0 1
rlabel polysilicon 597 -2384 597 -2384 0 3
rlabel polysilicon 604 -2378 604 -2378 0 1
rlabel polysilicon 604 -2384 604 -2384 0 3
rlabel polysilicon 611 -2378 611 -2378 0 1
rlabel polysilicon 614 -2378 614 -2378 0 2
rlabel polysilicon 611 -2384 611 -2384 0 3
rlabel polysilicon 614 -2384 614 -2384 0 4
rlabel polysilicon 618 -2378 618 -2378 0 1
rlabel polysilicon 618 -2384 618 -2384 0 3
rlabel polysilicon 625 -2378 625 -2378 0 1
rlabel polysilicon 625 -2384 625 -2384 0 3
rlabel polysilicon 632 -2378 632 -2378 0 1
rlabel polysilicon 632 -2384 632 -2384 0 3
rlabel polysilicon 639 -2378 639 -2378 0 1
rlabel polysilicon 639 -2384 639 -2384 0 3
rlabel polysilicon 646 -2384 646 -2384 0 3
rlabel polysilicon 653 -2378 653 -2378 0 1
rlabel polysilicon 653 -2384 653 -2384 0 3
rlabel polysilicon 660 -2378 660 -2378 0 1
rlabel polysilicon 660 -2384 660 -2384 0 3
rlabel polysilicon 667 -2378 667 -2378 0 1
rlabel polysilicon 667 -2384 667 -2384 0 3
rlabel polysilicon 674 -2378 674 -2378 0 1
rlabel polysilicon 674 -2384 674 -2384 0 3
rlabel polysilicon 681 -2378 681 -2378 0 1
rlabel polysilicon 681 -2384 681 -2384 0 3
rlabel polysilicon 688 -2378 688 -2378 0 1
rlabel polysilicon 688 -2384 688 -2384 0 3
rlabel polysilicon 695 -2378 695 -2378 0 1
rlabel polysilicon 698 -2378 698 -2378 0 2
rlabel polysilicon 698 -2384 698 -2384 0 4
rlabel polysilicon 702 -2378 702 -2378 0 1
rlabel polysilicon 702 -2384 702 -2384 0 3
rlabel polysilicon 709 -2378 709 -2378 0 1
rlabel polysilicon 709 -2384 709 -2384 0 3
rlabel polysilicon 716 -2378 716 -2378 0 1
rlabel polysilicon 719 -2378 719 -2378 0 2
rlabel polysilicon 716 -2384 716 -2384 0 3
rlabel polysilicon 730 -2378 730 -2378 0 1
rlabel polysilicon 730 -2384 730 -2384 0 3
rlabel polysilicon 737 -2378 737 -2378 0 1
rlabel polysilicon 737 -2384 737 -2384 0 3
rlabel polysilicon 744 -2378 744 -2378 0 1
rlabel polysilicon 744 -2384 744 -2384 0 3
rlabel polysilicon 751 -2378 751 -2378 0 1
rlabel polysilicon 751 -2384 751 -2384 0 3
rlabel polysilicon 758 -2378 758 -2378 0 1
rlabel polysilicon 758 -2384 758 -2384 0 3
rlabel polysilicon 765 -2378 765 -2378 0 1
rlabel polysilicon 765 -2384 765 -2384 0 3
rlabel polysilicon 772 -2378 772 -2378 0 1
rlabel polysilicon 772 -2384 772 -2384 0 3
rlabel polysilicon 779 -2378 779 -2378 0 1
rlabel polysilicon 779 -2384 779 -2384 0 3
rlabel polysilicon 793 -2378 793 -2378 0 1
rlabel polysilicon 793 -2384 793 -2384 0 3
rlabel polysilicon 800 -2378 800 -2378 0 1
rlabel polysilicon 800 -2384 800 -2384 0 3
rlabel polysilicon 814 -2378 814 -2378 0 1
rlabel polysilicon 814 -2384 814 -2384 0 3
rlabel polysilicon 898 -2378 898 -2378 0 1
rlabel polysilicon 898 -2384 898 -2384 0 3
rlabel polysilicon 905 -2378 905 -2378 0 1
rlabel polysilicon 905 -2384 905 -2384 0 3
rlabel polysilicon 940 -2378 940 -2378 0 1
rlabel polysilicon 940 -2384 940 -2384 0 3
rlabel polysilicon 978 -2378 978 -2378 0 2
rlabel polysilicon 975 -2384 975 -2384 0 3
rlabel polysilicon 978 -2384 978 -2384 0 4
rlabel polysilicon 982 -2378 982 -2378 0 1
rlabel polysilicon 982 -2384 982 -2384 0 3
rlabel polysilicon 989 -2378 989 -2378 0 1
rlabel polysilicon 989 -2384 989 -2384 0 3
rlabel polysilicon 1003 -2378 1003 -2378 0 1
rlabel polysilicon 1006 -2378 1006 -2378 0 2
rlabel polysilicon 1006 -2384 1006 -2384 0 4
rlabel polysilicon 198 -2429 198 -2429 0 1
rlabel polysilicon 198 -2435 198 -2435 0 3
rlabel polysilicon 219 -2429 219 -2429 0 1
rlabel polysilicon 219 -2435 219 -2435 0 3
rlabel polysilicon 226 -2429 226 -2429 0 1
rlabel polysilicon 226 -2435 226 -2435 0 3
rlabel polysilicon 233 -2429 233 -2429 0 1
rlabel polysilicon 233 -2435 233 -2435 0 3
rlabel polysilicon 240 -2429 240 -2429 0 1
rlabel polysilicon 240 -2435 240 -2435 0 3
rlabel polysilicon 247 -2429 247 -2429 0 1
rlabel polysilicon 254 -2429 254 -2429 0 1
rlabel polysilicon 254 -2435 254 -2435 0 3
rlabel polysilicon 261 -2429 261 -2429 0 1
rlabel polysilicon 261 -2435 261 -2435 0 3
rlabel polysilicon 268 -2429 268 -2429 0 1
rlabel polysilicon 268 -2435 268 -2435 0 3
rlabel polysilicon 275 -2429 275 -2429 0 1
rlabel polysilicon 275 -2435 275 -2435 0 3
rlabel polysilicon 282 -2429 282 -2429 0 1
rlabel polysilicon 282 -2435 282 -2435 0 3
rlabel polysilicon 289 -2429 289 -2429 0 1
rlabel polysilicon 289 -2435 289 -2435 0 3
rlabel polysilicon 296 -2429 296 -2429 0 1
rlabel polysilicon 296 -2435 296 -2435 0 3
rlabel polysilicon 303 -2429 303 -2429 0 1
rlabel polysilicon 303 -2435 303 -2435 0 3
rlabel polysilicon 310 -2429 310 -2429 0 1
rlabel polysilicon 310 -2435 310 -2435 0 3
rlabel polysilicon 317 -2429 317 -2429 0 1
rlabel polysilicon 317 -2435 317 -2435 0 3
rlabel polysilicon 324 -2429 324 -2429 0 1
rlabel polysilicon 327 -2435 327 -2435 0 4
rlabel polysilicon 331 -2429 331 -2429 0 1
rlabel polysilicon 331 -2435 331 -2435 0 3
rlabel polysilicon 338 -2429 338 -2429 0 1
rlabel polysilicon 338 -2435 338 -2435 0 3
rlabel polysilicon 345 -2429 345 -2429 0 1
rlabel polysilicon 345 -2435 345 -2435 0 3
rlabel polysilicon 355 -2429 355 -2429 0 2
rlabel polysilicon 352 -2435 352 -2435 0 3
rlabel polysilicon 359 -2429 359 -2429 0 1
rlabel polysilicon 359 -2435 359 -2435 0 3
rlabel polysilicon 369 -2429 369 -2429 0 2
rlabel polysilicon 366 -2435 366 -2435 0 3
rlabel polysilicon 369 -2435 369 -2435 0 4
rlabel polysilicon 373 -2429 373 -2429 0 1
rlabel polysilicon 373 -2435 373 -2435 0 3
rlabel polysilicon 380 -2429 380 -2429 0 1
rlabel polysilicon 383 -2429 383 -2429 0 2
rlabel polysilicon 380 -2435 380 -2435 0 3
rlabel polysilicon 387 -2429 387 -2429 0 1
rlabel polysilicon 387 -2435 387 -2435 0 3
rlabel polysilicon 394 -2429 394 -2429 0 1
rlabel polysilicon 394 -2435 394 -2435 0 3
rlabel polysilicon 401 -2429 401 -2429 0 1
rlabel polysilicon 401 -2435 401 -2435 0 3
rlabel polysilicon 408 -2429 408 -2429 0 1
rlabel polysilicon 408 -2435 408 -2435 0 3
rlabel polysilicon 418 -2429 418 -2429 0 2
rlabel polysilicon 415 -2435 415 -2435 0 3
rlabel polysilicon 418 -2435 418 -2435 0 4
rlabel polysilicon 422 -2429 422 -2429 0 1
rlabel polysilicon 422 -2435 422 -2435 0 3
rlabel polysilicon 429 -2429 429 -2429 0 1
rlabel polysilicon 429 -2435 429 -2435 0 3
rlabel polysilicon 436 -2429 436 -2429 0 1
rlabel polysilicon 436 -2435 436 -2435 0 3
rlabel polysilicon 443 -2429 443 -2429 0 1
rlabel polysilicon 443 -2435 443 -2435 0 3
rlabel polysilicon 450 -2429 450 -2429 0 1
rlabel polysilicon 450 -2435 450 -2435 0 3
rlabel polysilicon 453 -2435 453 -2435 0 4
rlabel polysilicon 460 -2429 460 -2429 0 2
rlabel polysilicon 457 -2435 457 -2435 0 3
rlabel polysilicon 460 -2435 460 -2435 0 4
rlabel polysilicon 464 -2429 464 -2429 0 1
rlabel polysilicon 464 -2435 464 -2435 0 3
rlabel polysilicon 471 -2429 471 -2429 0 1
rlabel polysilicon 471 -2435 471 -2435 0 3
rlabel polysilicon 478 -2429 478 -2429 0 1
rlabel polysilicon 478 -2435 478 -2435 0 3
rlabel polysilicon 488 -2429 488 -2429 0 2
rlabel polysilicon 485 -2435 485 -2435 0 3
rlabel polysilicon 492 -2429 492 -2429 0 1
rlabel polysilicon 492 -2435 492 -2435 0 3
rlabel polysilicon 499 -2429 499 -2429 0 1
rlabel polysilicon 499 -2435 499 -2435 0 3
rlabel polysilicon 506 -2429 506 -2429 0 1
rlabel polysilicon 509 -2429 509 -2429 0 2
rlabel polysilicon 506 -2435 506 -2435 0 3
rlabel polysilicon 509 -2435 509 -2435 0 4
rlabel polysilicon 513 -2429 513 -2429 0 1
rlabel polysilicon 516 -2429 516 -2429 0 2
rlabel polysilicon 516 -2435 516 -2435 0 4
rlabel polysilicon 520 -2429 520 -2429 0 1
rlabel polysilicon 523 -2429 523 -2429 0 2
rlabel polysilicon 523 -2435 523 -2435 0 4
rlabel polysilicon 527 -2429 527 -2429 0 1
rlabel polysilicon 527 -2435 527 -2435 0 3
rlabel polysilicon 534 -2429 534 -2429 0 1
rlabel polysilicon 534 -2435 534 -2435 0 3
rlabel polysilicon 541 -2429 541 -2429 0 1
rlabel polysilicon 541 -2435 541 -2435 0 3
rlabel polysilicon 548 -2429 548 -2429 0 1
rlabel polysilicon 548 -2435 548 -2435 0 3
rlabel polysilicon 555 -2429 555 -2429 0 1
rlabel polysilicon 555 -2435 555 -2435 0 3
rlabel polysilicon 562 -2429 562 -2429 0 1
rlabel polysilicon 562 -2435 562 -2435 0 3
rlabel polysilicon 569 -2429 569 -2429 0 1
rlabel polysilicon 569 -2435 569 -2435 0 3
rlabel polysilicon 572 -2435 572 -2435 0 4
rlabel polysilicon 576 -2429 576 -2429 0 1
rlabel polysilicon 576 -2435 576 -2435 0 3
rlabel polysilicon 583 -2429 583 -2429 0 1
rlabel polysilicon 583 -2435 583 -2435 0 3
rlabel polysilicon 590 -2429 590 -2429 0 1
rlabel polysilicon 590 -2435 590 -2435 0 3
rlabel polysilicon 597 -2429 597 -2429 0 1
rlabel polysilicon 597 -2435 597 -2435 0 3
rlabel polysilicon 604 -2429 604 -2429 0 1
rlabel polysilicon 604 -2435 604 -2435 0 3
rlabel polysilicon 611 -2429 611 -2429 0 1
rlabel polysilicon 611 -2435 611 -2435 0 3
rlabel polysilicon 618 -2429 618 -2429 0 1
rlabel polysilicon 618 -2435 618 -2435 0 3
rlabel polysilicon 625 -2429 625 -2429 0 1
rlabel polysilicon 625 -2435 625 -2435 0 3
rlabel polysilicon 632 -2429 632 -2429 0 1
rlabel polysilicon 632 -2435 632 -2435 0 3
rlabel polysilicon 646 -2429 646 -2429 0 1
rlabel polysilicon 646 -2435 646 -2435 0 3
rlabel polysilicon 653 -2429 653 -2429 0 1
rlabel polysilicon 653 -2435 653 -2435 0 3
rlabel polysilicon 660 -2429 660 -2429 0 1
rlabel polysilicon 660 -2435 660 -2435 0 3
rlabel polysilicon 663 -2435 663 -2435 0 4
rlabel polysilicon 667 -2429 667 -2429 0 1
rlabel polysilicon 667 -2435 667 -2435 0 3
rlabel polysilicon 674 -2429 674 -2429 0 1
rlabel polysilicon 674 -2435 674 -2435 0 3
rlabel polysilicon 681 -2429 681 -2429 0 1
rlabel polysilicon 684 -2429 684 -2429 0 2
rlabel polysilicon 688 -2429 688 -2429 0 1
rlabel polysilicon 691 -2429 691 -2429 0 2
rlabel polysilicon 688 -2435 688 -2435 0 3
rlabel polysilicon 691 -2435 691 -2435 0 4
rlabel polysilicon 716 -2429 716 -2429 0 1
rlabel polysilicon 716 -2435 716 -2435 0 3
rlabel polysilicon 723 -2429 723 -2429 0 1
rlabel polysilicon 723 -2435 723 -2435 0 3
rlabel polysilicon 730 -2429 730 -2429 0 1
rlabel polysilicon 730 -2435 730 -2435 0 3
rlabel polysilicon 737 -2429 737 -2429 0 1
rlabel polysilicon 737 -2435 737 -2435 0 3
rlabel polysilicon 744 -2429 744 -2429 0 1
rlabel polysilicon 744 -2435 744 -2435 0 3
rlabel polysilicon 747 -2435 747 -2435 0 4
rlabel polysilicon 751 -2429 751 -2429 0 1
rlabel polysilicon 751 -2435 751 -2435 0 3
rlabel polysilicon 758 -2429 758 -2429 0 1
rlabel polysilicon 758 -2435 758 -2435 0 3
rlabel polysilicon 765 -2429 765 -2429 0 1
rlabel polysilicon 765 -2435 765 -2435 0 3
rlabel polysilicon 772 -2429 772 -2429 0 1
rlabel polysilicon 772 -2435 772 -2435 0 3
rlabel polysilicon 800 -2429 800 -2429 0 1
rlabel polysilicon 800 -2435 800 -2435 0 3
rlabel polysilicon 807 -2429 807 -2429 0 1
rlabel polysilicon 807 -2435 807 -2435 0 3
rlabel polysilicon 828 -2429 828 -2429 0 1
rlabel polysilicon 828 -2435 828 -2435 0 3
rlabel polysilicon 891 -2429 891 -2429 0 1
rlabel polysilicon 891 -2435 891 -2435 0 3
rlabel polysilicon 898 -2429 898 -2429 0 1
rlabel polysilicon 898 -2435 898 -2435 0 3
rlabel polysilicon 905 -2429 905 -2429 0 1
rlabel polysilicon 905 -2435 905 -2435 0 3
rlabel polysilicon 908 -2435 908 -2435 0 4
rlabel polysilicon 226 -2470 226 -2470 0 1
rlabel polysilicon 226 -2476 226 -2476 0 3
rlabel polysilicon 233 -2470 233 -2470 0 1
rlabel polysilicon 236 -2470 236 -2470 0 2
rlabel polysilicon 240 -2470 240 -2470 0 1
rlabel polysilicon 240 -2476 240 -2476 0 3
rlabel polysilicon 247 -2476 247 -2476 0 3
rlabel polysilicon 254 -2470 254 -2470 0 1
rlabel polysilicon 254 -2476 254 -2476 0 3
rlabel polysilicon 296 -2470 296 -2470 0 1
rlabel polysilicon 296 -2476 296 -2476 0 3
rlabel polysilicon 310 -2470 310 -2470 0 1
rlabel polysilicon 310 -2476 310 -2476 0 3
rlabel polysilicon 331 -2470 331 -2470 0 1
rlabel polysilicon 331 -2476 331 -2476 0 3
rlabel polysilicon 341 -2470 341 -2470 0 2
rlabel polysilicon 341 -2476 341 -2476 0 4
rlabel polysilicon 345 -2470 345 -2470 0 1
rlabel polysilicon 348 -2470 348 -2470 0 2
rlabel polysilicon 348 -2476 348 -2476 0 4
rlabel polysilicon 352 -2470 352 -2470 0 1
rlabel polysilicon 352 -2476 352 -2476 0 3
rlabel polysilicon 359 -2470 359 -2470 0 1
rlabel polysilicon 359 -2476 359 -2476 0 3
rlabel polysilicon 366 -2470 366 -2470 0 1
rlabel polysilicon 366 -2476 366 -2476 0 3
rlabel polysilicon 373 -2470 373 -2470 0 1
rlabel polysilicon 373 -2476 373 -2476 0 3
rlabel polysilicon 387 -2470 387 -2470 0 1
rlabel polysilicon 387 -2476 387 -2476 0 3
rlabel polysilicon 394 -2470 394 -2470 0 1
rlabel polysilicon 394 -2476 394 -2476 0 3
rlabel polysilicon 401 -2470 401 -2470 0 1
rlabel polysilicon 401 -2476 401 -2476 0 3
rlabel polysilicon 408 -2470 408 -2470 0 1
rlabel polysilicon 408 -2476 408 -2476 0 3
rlabel polysilicon 422 -2470 422 -2470 0 1
rlabel polysilicon 422 -2476 422 -2476 0 3
rlabel polysilicon 432 -2470 432 -2470 0 2
rlabel polysilicon 429 -2476 429 -2476 0 3
rlabel polysilicon 432 -2476 432 -2476 0 4
rlabel polysilicon 436 -2470 436 -2470 0 1
rlabel polysilicon 436 -2476 436 -2476 0 3
rlabel polysilicon 443 -2470 443 -2470 0 1
rlabel polysilicon 443 -2476 443 -2476 0 3
rlabel polysilicon 446 -2476 446 -2476 0 4
rlabel polysilicon 450 -2470 450 -2470 0 1
rlabel polysilicon 453 -2470 453 -2470 0 2
rlabel polysilicon 453 -2476 453 -2476 0 4
rlabel polysilicon 457 -2470 457 -2470 0 1
rlabel polysilicon 457 -2476 457 -2476 0 3
rlabel polysilicon 464 -2470 464 -2470 0 1
rlabel polysilicon 464 -2476 464 -2476 0 3
rlabel polysilicon 471 -2470 471 -2470 0 1
rlabel polysilicon 471 -2476 471 -2476 0 3
rlabel polysilicon 478 -2470 478 -2470 0 1
rlabel polysilicon 478 -2476 478 -2476 0 3
rlabel polysilicon 485 -2470 485 -2470 0 1
rlabel polysilicon 485 -2476 485 -2476 0 3
rlabel polysilicon 492 -2470 492 -2470 0 1
rlabel polysilicon 492 -2476 492 -2476 0 3
rlabel polysilicon 499 -2470 499 -2470 0 1
rlabel polysilicon 499 -2476 499 -2476 0 3
rlabel polysilicon 509 -2470 509 -2470 0 2
rlabel polysilicon 509 -2476 509 -2476 0 4
rlabel polysilicon 513 -2470 513 -2470 0 1
rlabel polysilicon 513 -2476 513 -2476 0 3
rlabel polysilicon 527 -2470 527 -2470 0 1
rlabel polysilicon 527 -2476 527 -2476 0 3
rlabel polysilicon 541 -2470 541 -2470 0 1
rlabel polysilicon 541 -2476 541 -2476 0 3
rlabel polysilicon 548 -2470 548 -2470 0 1
rlabel polysilicon 548 -2476 548 -2476 0 3
rlabel polysilicon 576 -2470 576 -2470 0 1
rlabel polysilicon 576 -2476 576 -2476 0 3
rlabel polysilicon 597 -2470 597 -2470 0 1
rlabel polysilicon 597 -2476 597 -2476 0 3
rlabel polysilicon 607 -2470 607 -2470 0 2
rlabel polysilicon 604 -2476 604 -2476 0 3
rlabel polysilicon 611 -2470 611 -2470 0 1
rlabel polysilicon 614 -2470 614 -2470 0 2
rlabel polysilicon 614 -2476 614 -2476 0 4
rlabel polysilicon 618 -2470 618 -2470 0 1
rlabel polysilicon 618 -2476 618 -2476 0 3
rlabel polysilicon 625 -2470 625 -2470 0 1
rlabel polysilicon 625 -2476 625 -2476 0 3
rlabel polysilicon 632 -2470 632 -2470 0 1
rlabel polysilicon 632 -2476 632 -2476 0 3
rlabel polysilicon 639 -2470 639 -2470 0 1
rlabel polysilicon 639 -2476 639 -2476 0 3
rlabel polysilicon 646 -2470 646 -2470 0 1
rlabel polysilicon 649 -2470 649 -2470 0 2
rlabel polysilicon 649 -2476 649 -2476 0 4
rlabel polysilicon 653 -2470 653 -2470 0 1
rlabel polysilicon 653 -2476 653 -2476 0 3
rlabel polysilicon 660 -2470 660 -2470 0 1
rlabel polysilicon 663 -2470 663 -2470 0 2
rlabel polysilicon 660 -2476 660 -2476 0 3
rlabel polysilicon 674 -2470 674 -2470 0 1
rlabel polysilicon 674 -2476 674 -2476 0 3
rlabel polysilicon 688 -2470 688 -2470 0 1
rlabel polysilicon 688 -2476 688 -2476 0 3
rlabel polysilicon 702 -2470 702 -2470 0 1
rlabel polysilicon 702 -2476 702 -2476 0 3
rlabel polysilicon 723 -2470 723 -2470 0 1
rlabel polysilicon 723 -2476 723 -2476 0 3
rlabel polysilicon 744 -2470 744 -2470 0 1
rlabel polysilicon 744 -2476 744 -2476 0 3
rlabel polysilicon 751 -2470 751 -2470 0 1
rlabel polysilicon 754 -2470 754 -2470 0 2
rlabel polysilicon 751 -2476 751 -2476 0 3
rlabel polysilicon 807 -2470 807 -2470 0 1
rlabel polysilicon 807 -2476 807 -2476 0 3
rlabel polysilicon 817 -2470 817 -2470 0 2
rlabel polysilicon 817 -2476 817 -2476 0 4
rlabel polysilicon 828 -2470 828 -2470 0 1
rlabel polysilicon 828 -2476 828 -2476 0 3
rlabel polysilicon 838 -2470 838 -2470 0 2
rlabel polysilicon 835 -2476 835 -2476 0 3
rlabel polysilicon 898 -2470 898 -2470 0 1
rlabel polysilicon 898 -2476 898 -2476 0 3
rlabel polysilicon 226 -2491 226 -2491 0 1
rlabel polysilicon 226 -2497 226 -2497 0 3
rlabel polysilicon 233 -2497 233 -2497 0 3
rlabel polysilicon 236 -2497 236 -2497 0 4
rlabel polysilicon 240 -2491 240 -2491 0 1
rlabel polysilicon 240 -2497 240 -2497 0 3
rlabel polysilicon 359 -2491 359 -2491 0 1
rlabel polysilicon 359 -2497 359 -2497 0 3
rlabel polysilicon 366 -2491 366 -2491 0 1
rlabel polysilicon 369 -2491 369 -2491 0 2
rlabel polysilicon 366 -2497 366 -2497 0 3
rlabel polysilicon 373 -2491 373 -2491 0 1
rlabel polysilicon 373 -2497 373 -2497 0 3
rlabel polysilicon 380 -2491 380 -2491 0 1
rlabel polysilicon 380 -2497 380 -2497 0 3
rlabel polysilicon 387 -2491 387 -2491 0 1
rlabel polysilicon 390 -2491 390 -2491 0 2
rlabel polysilicon 394 -2491 394 -2491 0 1
rlabel polysilicon 394 -2497 394 -2497 0 3
rlabel polysilicon 397 -2497 397 -2497 0 4
rlabel polysilicon 401 -2491 401 -2491 0 1
rlabel polysilicon 404 -2491 404 -2491 0 2
rlabel polysilicon 401 -2497 401 -2497 0 3
rlabel polysilicon 408 -2491 408 -2491 0 1
rlabel polysilicon 408 -2497 408 -2497 0 3
rlabel polysilicon 534 -2491 534 -2491 0 1
rlabel polysilicon 534 -2497 534 -2497 0 3
rlabel polysilicon 548 -2491 548 -2491 0 1
rlabel polysilicon 551 -2491 551 -2491 0 2
rlabel polysilicon 548 -2497 548 -2497 0 3
rlabel polysilicon 555 -2491 555 -2491 0 1
rlabel polysilicon 558 -2497 558 -2497 0 4
rlabel polysilicon 604 -2491 604 -2491 0 1
rlabel polysilicon 604 -2497 604 -2497 0 3
rlabel polysilicon 611 -2491 611 -2491 0 1
rlabel polysilicon 614 -2491 614 -2491 0 2
rlabel polysilicon 611 -2497 611 -2497 0 3
rlabel polysilicon 632 -2491 632 -2491 0 1
rlabel polysilicon 632 -2497 632 -2497 0 3
rlabel polysilicon 653 -2491 653 -2491 0 1
rlabel polysilicon 653 -2497 653 -2497 0 3
rlabel polysilicon 660 -2491 660 -2491 0 1
rlabel polysilicon 660 -2497 660 -2497 0 3
rlabel polysilicon 688 -2491 688 -2491 0 1
rlabel polysilicon 691 -2491 691 -2491 0 2
rlabel polysilicon 691 -2497 691 -2497 0 4
rlabel polysilicon 702 -2491 702 -2491 0 1
rlabel polysilicon 702 -2497 702 -2497 0 3
rlabel polysilicon 723 -2491 723 -2491 0 1
rlabel polysilicon 726 -2491 726 -2491 0 2
rlabel polysilicon 726 -2497 726 -2497 0 4
rlabel polysilicon 901 -2491 901 -2491 0 2
rlabel polysilicon 898 -2497 898 -2497 0 3
rlabel polysilicon 901 -2497 901 -2497 0 4
rlabel polysilicon 905 -2491 905 -2491 0 1
rlabel polysilicon 905 -2497 905 -2497 0 3
rlabel metal2 152 1 152 1 0 net=880
rlabel metal2 338 1 338 1 0 net=3491
rlabel metal2 366 1 366 1 0 net=3885
rlabel metal2 432 1 432 1 0 net=4941
rlabel metal2 341 -1 341 -1 0 net=2923
rlabel metal2 394 -1 394 -1 0 net=6307
rlabel metal2 492 -1 492 -1 0 net=6759
rlabel metal2 345 -3 345 -3 0 net=2921
rlabel metal2 408 -3 408 -3 0 net=4303
rlabel metal2 464 -3 464 -3 0 net=7397
rlabel metal2 128 -14 128 -14 0 net=5909
rlabel metal2 198 -14 198 -14 0 net=1177
rlabel metal2 292 -14 292 -14 0 net=1679
rlabel metal2 320 -14 320 -14 0 net=3589
rlabel metal2 464 -14 464 -14 0 net=7399
rlabel metal2 502 -14 502 -14 0 net=7285
rlabel metal2 576 -14 576 -14 0 net=6761
rlabel metal2 208 -16 208 -16 0 net=1513
rlabel metal2 243 -16 243 -16 0 net=7149
rlabel metal2 282 -16 282 -16 0 net=2741
rlabel metal2 352 -16 352 -16 0 net=3493
rlabel metal2 415 -16 415 -16 0 net=5501
rlabel metal2 513 -16 513 -16 0 net=4943
rlabel metal2 593 -16 593 -16 0 net=5609
rlabel metal2 296 -18 296 -18 0 net=3505
rlabel metal2 450 -18 450 -18 0 net=4305
rlabel metal2 474 -18 474 -18 0 net=7217
rlabel metal2 303 -20 303 -20 0 net=1361
rlabel metal2 450 -20 450 -20 0 net=3447
rlabel metal2 324 -22 324 -22 0 net=2922
rlabel metal2 352 -22 352 -22 0 net=2341
rlabel metal2 436 -22 436 -22 0 net=4903
rlabel metal2 327 -24 327 -24 0 net=6645
rlabel metal2 429 -24 429 -24 0 net=3775
rlabel metal2 331 -26 331 -26 0 net=3887
rlabel metal2 376 -26 376 -26 0 net=2907
rlabel metal2 401 -26 401 -26 0 net=2969
rlabel metal2 464 -26 464 -26 0 net=5923
rlabel metal2 338 -28 338 -28 0 net=6309
rlabel metal2 401 -28 401 -28 0 net=2719
rlabel metal2 345 -30 345 -30 0 net=2383
rlabel metal2 359 -32 359 -32 0 net=2925
rlabel metal2 359 -32 359 -32 0 net=2925
rlabel metal2 366 -32 366 -32 0 net=2185
rlabel metal2 394 -32 394 -32 0 net=4423
rlabel metal2 373 -34 373 -34 0 net=3637
rlabel metal2 114 -45 114 -45 0 net=5910
rlabel metal2 142 -45 142 -45 0 net=1179
rlabel metal2 205 -45 205 -45 0 net=1515
rlabel metal2 233 -45 233 -45 0 net=1111
rlabel metal2 247 -45 247 -45 0 net=4439
rlabel metal2 415 -45 415 -45 0 net=5503
rlabel metal2 432 -45 432 -45 0 net=6895
rlabel metal2 593 -45 593 -45 0 net=7577
rlabel metal2 170 -47 170 -47 0 net=2477
rlabel metal2 254 -47 254 -47 0 net=7150
rlabel metal2 317 -47 317 -47 0 net=2909
rlabel metal2 443 -47 443 -47 0 net=4547
rlabel metal2 593 -47 593 -47 0 net=2805
rlabel metal2 618 -47 618 -47 0 net=5611
rlabel metal2 653 -47 653 -47 0 net=6491
rlabel metal2 191 -49 191 -49 0 net=3507
rlabel metal2 331 -49 331 -49 0 net=3889
rlabel metal2 443 -49 443 -49 0 net=4375
rlabel metal2 495 -49 495 -49 0 net=4595
rlabel metal2 625 -49 625 -49 0 net=6763
rlabel metal2 674 -49 674 -49 0 net=6793
rlabel metal2 198 -51 198 -51 0 net=1021
rlabel metal2 338 -51 338 -51 0 net=6310
rlabel metal2 394 -51 394 -51 0 net=6351
rlabel metal2 502 -51 502 -51 0 net=7041
rlabel metal2 212 -53 212 -53 0 net=1363
rlabel metal2 338 -53 338 -53 0 net=3495
rlabel metal2 478 -53 478 -53 0 net=4905
rlabel metal2 219 -55 219 -55 0 net=1681
rlabel metal2 359 -55 359 -55 0 net=2927
rlabel metal2 359 -55 359 -55 0 net=2927
rlabel metal2 369 -55 369 -55 0 net=5341
rlabel metal2 527 -55 527 -55 0 net=7218
rlabel metal2 534 -55 534 -55 0 net=6975
rlabel metal2 240 -57 240 -57 0 net=1183
rlabel metal2 380 -57 380 -57 0 net=5935
rlabel metal2 254 -59 254 -59 0 net=3449
rlabel metal2 478 -59 478 -59 0 net=6433
rlabel metal2 177 -61 177 -61 0 net=2165
rlabel metal2 485 -61 485 -61 0 net=7401
rlabel metal2 261 -63 261 -63 0 net=2187
rlabel metal2 408 -63 408 -63 0 net=6647
rlabel metal2 499 -63 499 -63 0 net=6909
rlabel metal2 541 -63 541 -63 0 net=4945
rlabel metal2 541 -63 541 -63 0 net=4945
rlabel metal2 548 -63 548 -63 0 net=7287
rlabel metal2 226 -65 226 -65 0 net=1921
rlabel metal2 387 -65 387 -65 0 net=6539
rlabel metal2 268 -67 268 -67 0 net=2235
rlabel metal2 408 -67 408 -67 0 net=3591
rlabel metal2 506 -67 506 -67 0 net=3639
rlabel metal2 282 -69 282 -69 0 net=2743
rlabel metal2 436 -69 436 -69 0 net=2971
rlabel metal2 474 -69 474 -69 0 net=4321
rlabel metal2 513 -69 513 -69 0 net=3777
rlabel metal2 282 -71 282 -71 0 net=2385
rlabel metal2 422 -71 422 -71 0 net=4425
rlabel metal2 446 -71 446 -71 0 net=5333
rlabel metal2 527 -71 527 -71 0 net=5633
rlabel metal2 163 -73 163 -73 0 net=2527
rlabel metal2 422 -73 422 -73 0 net=4307
rlabel metal2 289 -75 289 -75 0 net=2839
rlabel metal2 464 -75 464 -75 0 net=5925
rlabel metal2 289 -77 289 -77 0 net=2721
rlabel metal2 296 -79 296 -79 0 net=3563
rlabel metal2 184 -81 184 -81 0 net=4855
rlabel metal2 303 -83 303 -83 0 net=2343
rlabel metal2 373 -83 373 -83 0 net=3715
rlabel metal2 348 -85 348 -85 0 net=5425
rlabel metal2 352 -87 352 -87 0 net=2845
rlabel metal2 51 -98 51 -98 0 net=5015
rlabel metal2 464 -98 464 -98 0 net=5427
rlabel metal2 58 -100 58 -100 0 net=6401
rlabel metal2 471 -100 471 -100 0 net=7553
rlabel metal2 65 -102 65 -102 0 net=1181
rlabel metal2 145 -102 145 -102 0 net=4856
rlabel metal2 198 -102 198 -102 0 net=1023
rlabel metal2 275 -102 275 -102 0 net=697
rlabel metal2 394 -102 394 -102 0 net=7273
rlabel metal2 72 -104 72 -104 0 net=4517
rlabel metal2 86 -104 86 -104 0 net=2567
rlabel metal2 121 -104 121 -104 0 net=2893
rlabel metal2 198 -104 198 -104 0 net=2236
rlabel metal2 275 -104 275 -104 0 net=2009
rlabel metal2 485 -104 485 -104 0 net=6649
rlabel metal2 93 -106 93 -106 0 net=3565
rlabel metal2 331 -106 331 -106 0 net=195
rlabel metal2 485 -106 485 -106 0 net=3779
rlabel metal2 632 -106 632 -106 0 net=7289
rlabel metal2 107 -108 107 -108 0 net=4441
rlabel metal2 268 -108 268 -108 0 net=3497
rlabel metal2 345 -108 345 -108 0 net=5504
rlabel metal2 492 -108 492 -108 0 net=6353
rlabel metal2 114 -110 114 -110 0 net=3125
rlabel metal2 156 -110 156 -110 0 net=2723
rlabel metal2 359 -110 359 -110 0 net=2929
rlabel metal2 418 -110 418 -110 0 net=5121
rlabel metal2 639 -110 639 -110 0 net=4907
rlabel metal2 114 -112 114 -112 0 net=3537
rlabel metal2 324 -112 324 -112 0 net=2841
rlabel metal2 366 -112 366 -112 0 net=1245
rlabel metal2 450 -112 450 -112 0 net=4197
rlabel metal2 653 -112 653 -112 0 net=6493
rlabel metal2 128 -114 128 -114 0 net=3451
rlabel metal2 261 -114 261 -114 0 net=2189
rlabel metal2 310 -114 310 -114 0 net=2745
rlabel metal2 369 -114 369 -114 0 net=2987
rlabel metal2 495 -114 495 -114 0 net=6129
rlabel metal2 152 -116 152 -116 0 net=1769
rlabel metal2 303 -116 303 -116 0 net=2345
rlabel metal2 387 -116 387 -116 0 net=3717
rlabel metal2 520 -116 520 -116 0 net=5343
rlabel metal2 660 -116 660 -116 0 net=6765
rlabel metal2 170 -118 170 -118 0 net=2479
rlabel metal2 303 -118 303 -118 0 net=2241
rlabel metal2 478 -118 478 -118 0 net=5349
rlabel metal2 667 -118 667 -118 0 net=6977
rlabel metal2 170 -120 170 -120 0 net=1923
rlabel metal2 247 -120 247 -120 0 net=1551
rlabel metal2 534 -120 534 -120 0 net=6911
rlabel metal2 100 -122 100 -122 0 net=2773
rlabel metal2 254 -122 254 -122 0 net=2231
rlabel metal2 534 -122 534 -122 0 net=3803
rlabel metal2 583 -122 583 -122 0 net=7043
rlabel metal2 646 -122 646 -122 0 net=5613
rlabel metal2 674 -122 674 -122 0 net=6795
rlabel metal2 184 -124 184 -124 0 net=387
rlabel metal2 201 -124 201 -124 0 net=4301
rlabel metal2 380 -124 380 -124 0 net=2829
rlabel metal2 499 -124 499 -124 0 net=5335
rlabel metal2 681 -124 681 -124 0 net=7579
rlabel metal2 219 -126 219 -126 0 net=1683
rlabel metal2 436 -126 436 -126 0 net=4427
rlabel metal2 513 -126 513 -126 0 net=5927
rlabel metal2 688 -126 688 -126 0 net=7091
rlabel metal2 191 -128 191 -128 0 net=3509
rlabel metal2 467 -128 467 -128 0 net=4567
rlabel metal2 590 -128 590 -128 0 net=4597
rlabel metal2 625 -128 625 -128 0 net=6435
rlabel metal2 219 -130 219 -130 0 net=1185
rlabel metal2 317 -130 317 -130 0 net=2911
rlabel metal2 453 -130 453 -130 0 net=5149
rlabel metal2 205 -132 205 -132 0 net=1517
rlabel metal2 282 -132 282 -132 0 net=2387
rlabel metal2 481 -132 481 -132 0 net=4191
rlabel metal2 527 -132 527 -132 0 net=5635
rlabel metal2 177 -134 177 -134 0 net=2167
rlabel metal2 506 -134 506 -134 0 net=4323
rlabel metal2 548 -134 548 -134 0 net=6541
rlabel metal2 177 -136 177 -136 0 net=1365
rlabel metal2 373 -136 373 -136 0 net=4887
rlabel metal2 562 -136 562 -136 0 net=7403
rlabel metal2 163 -138 163 -138 0 net=2529
rlabel metal2 334 -138 334 -138 0 net=4459
rlabel metal2 569 -138 569 -138 0 net=6897
rlabel metal2 163 -140 163 -140 0 net=2847
rlabel metal2 373 -140 373 -140 0 net=2807
rlabel metal2 205 -142 205 -142 0 net=1113
rlabel metal2 352 -142 352 -142 0 net=5429
rlabel metal2 415 -144 415 -144 0 net=3891
rlabel metal2 541 -144 541 -144 0 net=4947
rlabel metal2 576 -144 576 -144 0 net=5937
rlabel metal2 345 -146 345 -146 0 net=2659
rlabel metal2 422 -146 422 -146 0 net=4309
rlabel metal2 555 -146 555 -146 0 net=4549
rlabel metal2 422 -148 422 -148 0 net=2973
rlabel metal2 520 -148 520 -148 0 net=4041
rlabel metal2 443 -150 443 -150 0 net=4377
rlabel metal2 408 -152 408 -152 0 net=3593
rlabel metal2 457 -152 457 -152 0 net=3641
rlabel metal2 593 -154 593 -154 0 net=4719
rlabel metal2 44 -165 44 -165 0 net=5537
rlabel metal2 191 -165 191 -165 0 net=2530
rlabel metal2 240 -165 240 -165 0 net=1519
rlabel metal2 240 -165 240 -165 0 net=1519
rlabel metal2 268 -165 268 -165 0 net=3498
rlabel metal2 362 -165 362 -165 0 net=6912
rlabel metal2 793 -165 793 -165 0 net=7093
rlabel metal2 65 -167 65 -167 0 net=1182
rlabel metal2 184 -167 184 -167 0 net=2347
rlabel metal2 348 -167 348 -167 0 net=6354
rlabel metal2 751 -167 751 -167 0 net=6979
rlabel metal2 800 -167 800 -167 0 net=7405
rlabel metal2 65 -169 65 -169 0 net=4519
rlabel metal2 79 -169 79 -169 0 net=2569
rlabel metal2 100 -169 100 -169 0 net=272
rlabel metal2 310 -169 310 -169 0 net=2747
rlabel metal2 352 -169 352 -169 0 net=792
rlabel metal2 464 -169 464 -169 0 net=6650
rlabel metal2 814 -169 814 -169 0 net=7555
rlabel metal2 72 -171 72 -171 0 net=2843
rlabel metal2 408 -171 408 -171 0 net=4908
rlabel metal2 821 -171 821 -171 0 net=7581
rlabel metal2 86 -173 86 -173 0 net=1839
rlabel metal2 198 -173 198 -173 0 net=1025
rlabel metal2 324 -173 324 -173 0 net=2975
rlabel metal2 471 -173 471 -173 0 net=7125
rlabel metal2 103 -175 103 -175 0 net=551
rlabel metal2 411 -175 411 -175 0 net=5428
rlabel metal2 730 -175 730 -175 0 net=6797
rlabel metal2 117 -177 117 -177 0 net=6377
rlabel metal2 772 -177 772 -177 0 net=7275
rlabel metal2 121 -179 121 -179 0 net=2894
rlabel metal2 212 -179 212 -179 0 net=2011
rlabel metal2 285 -179 285 -179 0 net=913
rlabel metal2 492 -179 492 -179 0 net=4888
rlabel metal2 576 -179 576 -179 0 net=7315
rlabel metal2 121 -181 121 -181 0 net=467
rlabel metal2 128 -181 128 -181 0 net=3453
rlabel metal2 495 -181 495 -181 0 net=6542
rlabel metal2 779 -181 779 -181 0 net=7291
rlabel metal2 128 -183 128 -183 0 net=2775
rlabel metal2 275 -183 275 -183 0 net=2389
rlabel metal2 415 -183 415 -183 0 net=6898
rlabel metal2 138 -185 138 -185 0 net=417
rlabel metal2 460 -185 460 -185 0 net=6365
rlabel metal2 145 -187 145 -187 0 net=1246
rlabel metal2 415 -187 415 -187 0 net=2871
rlabel metal2 495 -187 495 -187 0 net=6494
rlabel metal2 163 -189 163 -189 0 net=2849
rlabel metal2 443 -189 443 -189 0 net=3595
rlabel metal2 499 -189 499 -189 0 net=4429
rlabel metal2 632 -189 632 -189 0 net=7045
rlabel metal2 58 -191 58 -191 0 net=6402
rlabel metal2 177 -191 177 -191 0 net=1367
rlabel metal2 296 -191 296 -191 0 net=2481
rlabel metal2 359 -191 359 -191 0 net=6095
rlabel metal2 51 -193 51 -193 0 net=5017
rlabel metal2 177 -193 177 -193 0 net=1553
rlabel metal2 282 -193 282 -193 0 net=2169
rlabel metal2 366 -193 366 -193 0 net=2913
rlabel metal2 443 -193 443 -193 0 net=2979
rlabel metal2 520 -193 520 -193 0 net=4043
rlabel metal2 548 -193 548 -193 0 net=4461
rlabel metal2 660 -193 660 -193 0 net=5351
rlabel metal2 730 -193 730 -193 0 net=5931
rlabel metal2 51 -195 51 -195 0 net=3719
rlabel metal2 450 -195 450 -195 0 net=4889
rlabel metal2 667 -195 667 -195 0 net=5615
rlabel metal2 709 -195 709 -195 0 net=6131
rlabel metal2 191 -197 191 -197 0 net=1187
rlabel metal2 247 -197 247 -197 0 net=2831
rlabel metal2 429 -197 429 -197 0 net=2989
rlabel metal2 457 -197 457 -197 0 net=3643
rlabel metal2 520 -197 520 -197 0 net=3805
rlabel metal2 618 -197 618 -197 0 net=5151
rlabel metal2 681 -197 681 -197 0 net=5929
rlabel metal2 205 -199 205 -199 0 net=1115
rlabel metal2 226 -199 226 -199 0 net=2653
rlabel metal2 474 -199 474 -199 0 net=5385
rlabel metal2 688 -199 688 -199 0 net=6437
rlabel metal2 205 -201 205 -201 0 net=2233
rlabel metal2 303 -201 303 -201 0 net=2243
rlabel metal2 394 -201 394 -201 0 net=2931
rlabel metal2 439 -201 439 -201 0 net=4821
rlabel metal2 646 -201 646 -201 0 net=5337
rlabel metal2 702 -201 702 -201 0 net=5939
rlabel metal2 716 -201 716 -201 0 net=6767
rlabel metal2 156 -203 156 -203 0 net=2725
rlabel metal2 474 -203 474 -203 0 net=4310
rlabel metal2 653 -203 653 -203 0 net=5345
rlabel metal2 114 -205 114 -205 0 net=3539
rlabel metal2 254 -205 254 -205 0 net=1907
rlabel metal2 289 -205 289 -205 0 net=2191
rlabel metal2 331 -205 331 -205 0 net=4302
rlabel metal2 404 -205 404 -205 0 net=4061
rlabel metal2 639 -205 639 -205 0 net=4199
rlabel metal2 674 -205 674 -205 0 net=5637
rlabel metal2 289 -207 289 -207 0 net=5045
rlabel metal2 331 -209 331 -209 0 net=3511
rlabel metal2 492 -209 492 -209 0 net=6083
rlabel metal2 338 -211 338 -211 0 net=1684
rlabel metal2 569 -211 569 -211 0 net=4949
rlabel metal2 261 -213 261 -213 0 net=1771
rlabel metal2 373 -213 373 -213 0 net=2809
rlabel metal2 527 -213 527 -213 0 net=4325
rlabel metal2 611 -213 611 -213 0 net=5123
rlabel metal2 261 -215 261 -215 0 net=2661
rlabel metal2 506 -215 506 -215 0 net=3893
rlabel metal2 555 -215 555 -215 0 net=4379
rlabel metal2 583 -215 583 -215 0 net=4569
rlabel metal2 107 -217 107 -217 0 net=4443
rlabel metal2 107 -219 107 -219 0 net=2135
rlabel metal2 345 -219 345 -219 0 net=5430
rlabel metal2 142 -221 142 -221 0 net=5733
rlabel metal2 597 -221 597 -221 0 net=4551
rlabel metal2 142 -223 142 -223 0 net=1283
rlabel metal2 597 -223 597 -223 0 net=4721
rlabel metal2 149 -225 149 -225 0 net=4999
rlabel metal2 590 -225 590 -225 0 net=4599
rlabel metal2 149 -227 149 -227 0 net=1925
rlabel metal2 513 -227 513 -227 0 net=4193
rlabel metal2 135 -229 135 -229 0 net=3127
rlabel metal2 485 -229 485 -229 0 net=3781
rlabel metal2 93 -231 93 -231 0 net=3567
rlabel metal2 93 -233 93 -233 0 net=1285
rlabel metal2 135 -235 135 -235 0 net=157
rlabel metal2 2 -246 2 -246 0 net=3835
rlabel metal2 72 -246 72 -246 0 net=2844
rlabel metal2 352 -246 352 -246 0 net=5930
rlabel metal2 807 -246 807 -246 0 net=7127
rlabel metal2 9 -248 9 -248 0 net=6579
rlabel metal2 289 -248 289 -248 0 net=2748
rlabel metal2 352 -248 352 -248 0 net=4045
rlabel metal2 569 -248 569 -248 0 net=4381
rlabel metal2 16 -250 16 -250 0 net=5431
rlabel metal2 383 -250 383 -250 0 net=5124
rlabel metal2 681 -250 681 -250 0 net=5347
rlabel metal2 23 -252 23 -252 0 net=5019
rlabel metal2 72 -252 72 -252 0 net=1909
rlabel metal2 289 -252 289 -252 0 net=2991
rlabel metal2 471 -252 471 -252 0 net=6917
rlabel metal2 30 -254 30 -254 0 net=6065
rlabel metal2 492 -254 492 -254 0 net=4570
rlabel metal2 730 -254 730 -254 0 net=5933
rlabel metal2 37 -256 37 -256 0 net=4521
rlabel metal2 86 -256 86 -256 0 net=1840
rlabel metal2 303 -256 303 -256 0 net=2193
rlabel metal2 359 -256 359 -256 0 net=2583
rlabel metal2 513 -256 513 -256 0 net=3783
rlabel metal2 513 -256 513 -256 0 net=3783
rlabel metal2 520 -256 520 -256 0 net=3807
rlabel metal2 548 -256 548 -256 0 net=4463
rlabel metal2 667 -256 667 -256 0 net=5387
rlabel metal2 744 -256 744 -256 0 net=6439
rlabel metal2 814 -256 814 -256 0 net=7277
rlabel metal2 51 -258 51 -258 0 net=3720
rlabel metal2 268 -258 268 -258 0 net=1773
rlabel metal2 401 -258 401 -258 0 net=4194
rlabel metal2 597 -258 597 -258 0 net=4723
rlabel metal2 758 -258 758 -258 0 net=6367
rlabel metal2 51 -260 51 -260 0 net=2727
rlabel metal2 418 -260 418 -260 0 net=5815
rlabel metal2 821 -260 821 -260 0 net=7293
rlabel metal2 58 -262 58 -262 0 net=3645
rlabel metal2 506 -262 506 -262 0 net=5735
rlabel metal2 758 -262 758 -262 0 net=7047
rlabel metal2 828 -262 828 -262 0 net=7317
rlabel metal2 65 -264 65 -264 0 net=7255
rlabel metal2 79 -266 79 -266 0 net=2571
rlabel metal2 93 -266 93 -266 0 net=1286
rlabel metal2 303 -266 303 -266 0 net=544
rlabel metal2 376 -266 376 -266 0 net=4015
rlabel metal2 520 -266 520 -266 0 net=3895
rlabel metal2 555 -266 555 -266 0 net=5001
rlabel metal2 751 -266 751 -266 0 net=6133
rlabel metal2 835 -266 835 -266 0 net=7557
rlabel metal2 79 -268 79 -268 0 net=2981
rlabel metal2 464 -268 464 -268 0 net=3455
rlabel metal2 541 -268 541 -268 0 net=4063
rlabel metal2 569 -268 569 -268 0 net=4327
rlabel metal2 653 -268 653 -268 0 net=4201
rlabel metal2 723 -268 723 -268 0 net=5353
rlabel metal2 765 -268 765 -268 0 net=6379
rlabel metal2 842 -268 842 -268 0 net=7583
rlabel metal2 93 -270 93 -270 0 net=5041
rlabel metal2 103 -270 103 -270 0 net=4237
rlabel metal2 632 -270 632 -270 0 net=4891
rlabel metal2 709 -270 709 -270 0 net=5941
rlabel metal2 793 -270 793 -270 0 net=6981
rlabel metal2 849 -270 849 -270 0 net=7095
rlabel metal2 100 -272 100 -272 0 net=2873
rlabel metal2 425 -272 425 -272 0 net=7406
rlabel metal2 121 -274 121 -274 0 net=409
rlabel metal2 170 -274 170 -274 0 net=3129
rlabel metal2 338 -274 338 -274 0 net=3417
rlabel metal2 387 -274 387 -274 0 net=2810
rlabel metal2 450 -274 450 -274 0 net=6711
rlabel metal2 121 -276 121 -276 0 net=2915
rlabel metal2 394 -276 394 -276 0 net=5338
rlabel metal2 702 -276 702 -276 0 net=5639
rlabel metal2 142 -278 142 -278 0 net=1284
rlabel metal2 366 -278 366 -278 0 net=2195
rlabel metal2 576 -278 576 -278 0 net=4431
rlabel metal2 583 -278 583 -278 0 net=4445
rlabel metal2 646 -278 646 -278 0 net=5047
rlabel metal2 772 -278 772 -278 0 net=6769
rlabel metal2 142 -280 142 -280 0 net=1271
rlabel metal2 474 -280 474 -280 0 net=3899
rlabel metal2 576 -280 576 -280 0 net=4601
rlabel metal2 625 -280 625 -280 0 net=4553
rlabel metal2 660 -280 660 -280 0 net=5153
rlabel metal2 716 -280 716 -280 0 net=6085
rlabel metal2 786 -280 786 -280 0 net=6799
rlabel metal2 149 -282 149 -282 0 net=1927
rlabel metal2 149 -282 149 -282 0 net=1927
rlabel metal2 156 -282 156 -282 0 net=3541
rlabel metal2 397 -282 397 -282 0 net=6355
rlabel metal2 156 -284 156 -284 0 net=2391
rlabel metal2 425 -284 425 -284 0 net=4027
rlabel metal2 551 -284 551 -284 0 net=5299
rlabel metal2 737 -284 737 -284 0 net=6097
rlabel metal2 163 -286 163 -286 0 net=2663
rlabel metal2 275 -286 275 -286 0 net=1197
rlabel metal2 436 -286 436 -286 0 net=6403
rlabel metal2 44 -288 44 -288 0 net=5538
rlabel metal2 439 -288 439 -288 0 net=5959
rlabel metal2 170 -290 170 -290 0 net=3513
rlabel metal2 457 -290 457 -290 0 net=4067
rlabel metal2 639 -290 639 -290 0 net=4951
rlabel metal2 688 -290 688 -290 0 net=7253
rlabel metal2 128 -292 128 -292 0 net=2777
rlabel metal2 457 -292 457 -292 0 net=4677
rlabel metal2 695 -292 695 -292 0 net=5617
rlabel metal2 177 -294 177 -294 0 net=1555
rlabel metal2 177 -294 177 -294 0 net=1555
rlabel metal2 184 -294 184 -294 0 net=2348
rlabel metal2 478 -294 478 -294 0 net=3597
rlabel metal2 579 -294 579 -294 0 net=1
rlabel metal2 618 -294 618 -294 0 net=4823
rlabel metal2 166 -296 166 -296 0 net=7533
rlabel metal2 184 -298 184 -298 0 net=1189
rlabel metal2 205 -298 205 -298 0 net=2234
rlabel metal2 478 -298 478 -298 0 net=3569
rlabel metal2 488 -298 488 -298 0 net=4531
rlabel metal2 107 -300 107 -300 0 net=2136
rlabel metal2 205 -300 205 -300 0 net=1117
rlabel metal2 240 -300 240 -300 0 net=1521
rlabel metal2 240 -300 240 -300 0 net=1521
rlabel metal2 254 -300 254 -300 0 net=1731
rlabel metal2 485 -300 485 -300 0 net=4326
rlabel metal2 107 -302 107 -302 0 net=4797
rlabel metal2 219 -302 219 -302 0 net=1369
rlabel metal2 261 -302 261 -302 0 net=1733
rlabel metal2 446 -302 446 -302 0 net=4187
rlabel metal2 198 -304 198 -304 0 net=1027
rlabel metal2 247 -304 247 -304 0 net=2832
rlabel metal2 114 -306 114 -306 0 net=2433
rlabel metal2 317 -306 317 -306 0 net=2483
rlabel metal2 114 -308 114 -308 0 net=2933
rlabel metal2 198 -310 198 -310 0 net=2171
rlabel metal2 380 -310 380 -310 0 net=2245
rlabel metal2 44 -312 44 -312 0 net=3651
rlabel metal2 135 -314 135 -314 0 net=2103
rlabel metal2 135 -316 135 -316 0 net=2013
rlabel metal2 226 -316 226 -316 0 net=2655
rlabel metal2 212 -318 212 -318 0 net=2977
rlabel metal2 226 -320 226 -320 0 net=2851
rlabel metal2 117 -322 117 -322 0 net=3653
rlabel metal2 324 -324 324 -324 0 net=3909
rlabel metal2 16 -335 16 -335 0 net=5432
rlabel metal2 436 -335 436 -335 0 net=4724
rlabel metal2 905 -335 905 -335 0 net=7129
rlabel metal2 16 -337 16 -337 0 net=4799
rlabel metal2 124 -337 124 -337 0 net=3130
rlabel metal2 289 -337 289 -337 0 net=2992
rlabel metal2 401 -337 401 -337 0 net=4824
rlabel metal2 758 -337 758 -337 0 net=7049
rlabel metal2 912 -337 912 -337 0 net=7257
rlabel metal2 44 -339 44 -339 0 net=3652
rlabel metal2 79 -339 79 -339 0 net=2983
rlabel metal2 439 -339 439 -339 0 net=225
rlabel metal2 618 -339 618 -339 0 net=7535
rlabel metal2 37 -341 37 -341 0 net=4522
rlabel metal2 96 -341 96 -341 0 net=4691
rlabel metal2 730 -341 730 -341 0 net=5389
rlabel metal2 779 -341 779 -341 0 net=6441
rlabel metal2 919 -341 919 -341 0 net=7295
rlabel metal2 2 -343 2 -343 0 net=3837
rlabel metal2 44 -343 44 -343 0 net=5043
rlabel metal2 100 -343 100 -343 0 net=2875
rlabel metal2 296 -343 296 -343 0 net=2105
rlabel metal2 310 -343 310 -343 0 net=2194
rlabel metal2 467 -343 467 -343 0 net=5934
rlabel metal2 926 -343 926 -343 0 net=7319
rlabel metal2 2 -345 2 -345 0 net=2485
rlabel metal2 355 -345 355 -345 0 net=3299
rlabel metal2 443 -345 443 -345 0 net=7453
rlabel metal2 51 -347 51 -347 0 net=2728
rlabel metal2 467 -347 467 -347 0 net=7254
rlabel metal2 933 -347 933 -347 0 net=7559
rlabel metal2 51 -349 51 -349 0 net=4863
rlabel metal2 548 -349 548 -349 0 net=7263
rlabel metal2 65 -351 65 -351 0 net=2664
rlabel metal2 191 -351 191 -351 0 net=1983
rlabel metal2 331 -351 331 -351 0 net=2779
rlabel metal2 411 -351 411 -351 0 net=4382
rlabel metal2 947 -351 947 -351 0 net=7585
rlabel metal2 947 -351 947 -351 0 net=7585
rlabel metal2 93 -353 93 -353 0 net=2172
rlabel metal2 205 -353 205 -353 0 net=1119
rlabel metal2 205 -353 205 -353 0 net=1119
rlabel metal2 212 -353 212 -353 0 net=2978
rlabel metal2 457 -353 457 -353 0 net=7278
rlabel metal2 100 -355 100 -355 0 net=1273
rlabel metal2 149 -355 149 -355 0 net=1929
rlabel metal2 198 -355 198 -355 0 net=1029
rlabel metal2 243 -355 243 -355 0 net=2025
rlabel metal2 296 -355 296 -355 0 net=3037
rlabel metal2 583 -355 583 -355 0 net=4068
rlabel metal2 621 -355 621 -355 0 net=6165
rlabel metal2 793 -355 793 -355 0 net=6801
rlabel metal2 107 -357 107 -357 0 net=3575
rlabel metal2 142 -357 142 -357 0 net=1371
rlabel metal2 226 -357 226 -357 0 net=2852
rlabel metal2 422 -357 422 -357 0 net=6369
rlabel metal2 72 -359 72 -359 0 net=1911
rlabel metal2 233 -359 233 -359 0 net=1261
rlabel metal2 380 -359 380 -359 0 net=3131
rlabel metal2 667 -359 667 -359 0 net=4203
rlabel metal2 751 -359 751 -359 0 net=5355
rlabel metal2 800 -359 800 -359 0 net=6135
rlabel metal2 114 -361 114 -361 0 net=2934
rlabel metal2 446 -361 446 -361 0 net=4446
rlabel metal2 744 -361 744 -361 0 net=5737
rlabel metal2 842 -361 842 -361 0 net=6713
rlabel metal2 86 -363 86 -363 0 net=2573
rlabel metal2 177 -363 177 -363 0 net=1557
rlabel metal2 254 -363 254 -363 0 net=1732
rlabel metal2 387 -363 387 -363 0 net=3543
rlabel metal2 457 -363 457 -363 0 net=4602
rlabel metal2 597 -363 597 -363 0 net=4329
rlabel metal2 702 -363 702 -363 0 net=5049
rlabel metal2 786 -363 786 -363 0 net=6099
rlabel metal2 849 -363 849 -363 0 net=6771
rlabel metal2 177 -365 177 -365 0 net=1191
rlabel metal2 194 -365 194 -365 0 net=4801
rlabel metal2 737 -365 737 -365 0 net=5619
rlabel metal2 814 -365 814 -365 0 net=6983
rlabel metal2 856 -365 856 -365 0 net=6919
rlabel metal2 128 -367 128 -367 0 net=88
rlabel metal2 254 -367 254 -367 0 net=1199
rlabel metal2 338 -367 338 -367 0 net=3419
rlabel metal2 464 -367 464 -367 0 net=6151
rlabel metal2 877 -367 877 -367 0 net=7097
rlabel metal2 128 -369 128 -369 0 net=2015
rlabel metal2 156 -369 156 -369 0 net=2393
rlabel metal2 352 -369 352 -369 0 net=4047
rlabel metal2 632 -369 632 -369 0 net=4679
rlabel metal2 660 -369 660 -369 0 net=4953
rlabel metal2 835 -369 835 -369 0 net=6405
rlabel metal2 86 -371 86 -371 0 net=3287
rlabel metal2 156 -371 156 -371 0 net=2656
rlabel metal2 359 -371 359 -371 0 net=2584
rlabel metal2 485 -371 485 -371 0 net=6899
rlabel metal2 772 -371 772 -371 0 net=6087
rlabel metal2 170 -373 170 -373 0 net=3514
rlabel metal2 373 -373 373 -373 0 net=6368
rlabel metal2 82 -375 82 -375 0 net=2737
rlabel metal2 212 -375 212 -375 0 net=3617
rlabel metal2 387 -375 387 -375 0 net=2247
rlabel metal2 464 -375 464 -375 0 net=3553
rlabel metal2 516 -375 516 -375 0 net=4263
rlabel metal2 646 -375 646 -375 0 net=4555
rlabel metal2 709 -375 709 -375 0 net=5155
rlabel metal2 261 -377 261 -377 0 net=1735
rlabel metal2 425 -377 425 -377 0 net=3997
rlabel metal2 653 -377 653 -377 0 net=4893
rlabel metal2 723 -377 723 -377 0 net=5943
rlabel metal2 247 -379 247 -379 0 net=2435
rlabel metal2 268 -379 268 -379 0 net=1775
rlabel metal2 429 -379 429 -379 0 net=3277
rlabel metal2 471 -379 471 -379 0 net=5640
rlabel metal2 72 -381 72 -381 0 net=3525
rlabel metal2 541 -381 541 -381 0 net=3901
rlabel metal2 625 -381 625 -381 0 net=4533
rlabel metal2 674 -381 674 -381 0 net=5003
rlabel metal2 821 -381 821 -381 0 net=6357
rlabel metal2 121 -383 121 -383 0 net=2917
rlabel metal2 275 -383 275 -383 0 net=3169
rlabel metal2 506 -383 506 -383 0 net=3457
rlabel metal2 551 -383 551 -383 0 net=5539
rlabel metal2 23 -385 23 -385 0 net=5020
rlabel metal2 240 -385 240 -385 0 net=1523
rlabel metal2 306 -385 306 -385 0 net=4267
rlabel metal2 765 -385 765 -385 0 net=5961
rlabel metal2 23 -387 23 -387 0 net=6067
rlabel metal2 58 -387 58 -387 0 net=3647
rlabel metal2 520 -387 520 -387 0 net=3897
rlabel metal2 716 -387 716 -387 0 net=5301
rlabel metal2 30 -389 30 -389 0 net=2349
rlabel metal2 149 -389 149 -389 0 net=2379
rlabel metal2 317 -389 317 -389 0 net=2197
rlabel metal2 394 -389 394 -389 0 net=5816
rlabel metal2 58 -391 58 -391 0 net=3911
rlabel metal2 362 -391 362 -391 0 net=5721
rlabel metal2 688 -391 688 -391 0 net=6199
rlabel metal2 68 -393 68 -393 0 net=2455
rlabel metal2 366 -393 366 -393 0 net=2317
rlabel metal2 513 -393 513 -393 0 net=3785
rlabel metal2 562 -393 562 -393 0 net=4189
rlabel metal2 324 -395 324 -395 0 net=4065
rlabel metal2 569 -395 569 -395 0 net=5143
rlabel metal2 499 -397 499 -397 0 net=4017
rlabel metal2 569 -397 569 -397 0 net=4465
rlabel metal2 478 -399 478 -399 0 net=3571
rlabel metal2 513 -399 513 -399 0 net=5348
rlabel metal2 478 -401 478 -401 0 net=3599
rlabel metal2 527 -401 527 -401 0 net=3809
rlabel metal2 590 -401 590 -401 0 net=4239
rlabel metal2 828 -401 828 -401 0 net=6381
rlabel metal2 9 -403 9 -403 0 net=6580
rlabel metal2 534 -403 534 -403 0 net=4029
rlabel metal2 604 -403 604 -403 0 net=4433
rlabel metal2 9 -405 9 -405 0 net=6181
rlabel metal2 159 -405 159 -405 0 net=6071
rlabel metal2 404 -407 404 -407 0 net=4159
rlabel metal2 408 -409 408 -409 0 net=3655
rlabel metal2 408 -411 408 -411 0 net=3017
rlabel metal2 9 -422 9 -422 0 net=6182
rlabel metal2 142 -422 142 -422 0 net=1372
rlabel metal2 275 -422 275 -422 0 net=3171
rlabel metal2 362 -422 362 -422 0 net=3898
rlabel metal2 695 -422 695 -422 0 net=4205
rlabel metal2 695 -422 695 -422 0 net=4205
rlabel metal2 814 -422 814 -422 0 net=5945
rlabel metal2 9 -424 9 -424 0 net=4265
rlabel metal2 849 -424 849 -424 0 net=6985
rlabel metal2 16 -426 16 -426 0 net=4800
rlabel metal2 114 -426 114 -426 0 net=2575
rlabel metal2 114 -426 114 -426 0 net=2575
rlabel metal2 156 -426 156 -426 0 net=2876
rlabel metal2 324 -426 324 -426 0 net=4066
rlabel metal2 415 -426 415 -426 0 net=2985
rlabel metal2 912 -426 912 -426 0 net=6443
rlabel metal2 16 -428 16 -428 0 net=4535
rlabel metal2 765 -428 765 -428 0 net=5303
rlabel metal2 926 -428 926 -428 0 net=6773
rlabel metal2 23 -430 23 -430 0 net=6068
rlabel metal2 191 -430 191 -430 0 net=3544
rlabel metal2 429 -430 429 -430 0 net=4434
rlabel metal2 828 -430 828 -430 0 net=6073
rlabel metal2 933 -430 933 -430 0 net=6803
rlabel metal2 1024 -430 1024 -430 0 net=7259
rlabel metal2 23 -432 23 -432 0 net=4077
rlabel metal2 394 -432 394 -432 0 net=7323
rlabel metal2 828 -432 828 -432 0 net=6383
rlabel metal2 940 -432 940 -432 0 net=6921
rlabel metal2 30 -434 30 -434 0 net=2350
rlabel metal2 198 -434 198 -434 0 net=1031
rlabel metal2 198 -434 198 -434 0 net=1031
rlabel metal2 226 -434 226 -434 0 net=1912
rlabel metal2 373 -434 373 -434 0 net=1776
rlabel metal2 513 -434 513 -434 0 net=3657
rlabel metal2 548 -434 548 -434 0 net=6136
rlabel metal2 940 -434 940 -434 0 net=7537
rlabel metal2 30 -436 30 -436 0 net=3913
rlabel metal2 65 -436 65 -436 0 net=378
rlabel metal2 397 -436 397 -436 0 net=4330
rlabel metal2 670 -436 670 -436 0 net=6697
rlabel metal2 37 -438 37 -438 0 net=3838
rlabel metal2 86 -438 86 -438 0 net=1275
rlabel metal2 163 -438 163 -438 0 net=1931
rlabel metal2 219 -438 219 -438 0 net=1559
rlabel metal2 275 -438 275 -438 0 net=1883
rlabel metal2 401 -438 401 -438 0 net=2781
rlabel metal2 432 -438 432 -438 0 net=6200
rlabel metal2 730 -438 730 -438 0 net=6901
rlabel metal2 37 -440 37 -440 0 net=2881
rlabel metal2 100 -440 100 -440 0 net=3577
rlabel metal2 184 -440 184 -440 0 net=2199
rlabel metal2 324 -440 324 -440 0 net=3731
rlabel metal2 450 -440 450 -440 0 net=3279
rlabel metal2 467 -440 467 -440 0 net=3600
rlabel metal2 523 -440 523 -440 0 net=7211
rlabel metal2 44 -442 44 -442 0 net=5044
rlabel metal2 187 -442 187 -442 0 net=2181
rlabel metal2 296 -442 296 -442 0 net=3039
rlabel metal2 450 -442 450 -442 0 net=5005
rlabel metal2 730 -442 730 -442 0 net=5145
rlabel metal2 786 -442 786 -442 0 net=5621
rlabel metal2 954 -442 954 -442 0 net=7099
rlabel metal2 44 -444 44 -444 0 net=3371
rlabel metal2 310 -444 310 -444 0 net=1985
rlabel metal2 331 -444 331 -444 0 net=2457
rlabel metal2 401 -444 401 -444 0 net=2749
rlabel metal2 478 -444 478 -444 0 net=7050
rlabel metal2 961 -444 961 -444 0 net=7131
rlabel metal2 51 -446 51 -446 0 net=4864
rlabel metal2 247 -446 247 -446 0 net=1525
rlabel metal2 331 -446 331 -446 0 net=2319
rlabel metal2 460 -446 460 -446 0 net=6263
rlabel metal2 968 -446 968 -446 0 net=7265
rlabel metal2 51 -448 51 -448 0 net=3555
rlabel metal2 530 -448 530 -448 0 net=5156
rlabel metal2 975 -448 975 -448 0 net=7561
rlabel metal2 58 -450 58 -450 0 net=3353
rlabel metal2 555 -450 555 -450 0 net=3811
rlabel metal2 555 -450 555 -450 0 net=3811
rlabel metal2 562 -450 562 -450 0 net=4019
rlabel metal2 649 -450 649 -450 0 net=4759
rlabel metal2 772 -450 772 -450 0 net=5541
rlabel metal2 884 -450 884 -450 0 net=6371
rlabel metal2 982 -450 982 -450 0 net=7297
rlabel metal2 65 -452 65 -452 0 net=2249
rlabel metal2 408 -452 408 -452 0 net=505
rlabel metal2 576 -452 576 -452 0 net=3999
rlabel metal2 674 -452 674 -452 0 net=5723
rlabel metal2 989 -452 989 -452 0 net=7321
rlabel metal2 68 -454 68 -454 0 net=4243
rlabel metal2 737 -454 737 -454 0 net=4955
rlabel metal2 996 -454 996 -454 0 net=7455
rlabel metal2 72 -456 72 -456 0 net=3561
rlabel metal2 709 -456 709 -456 0 net=4895
rlabel metal2 800 -456 800 -456 0 net=5739
rlabel metal2 75 -458 75 -458 0 net=1699
rlabel metal2 121 -458 121 -458 0 net=5603
rlabel metal2 79 -460 79 -460 0 net=2739
rlabel metal2 205 -460 205 -460 0 net=1120
rlabel metal2 261 -460 261 -460 0 net=2437
rlabel metal2 387 -460 387 -460 0 net=6845
rlabel metal2 82 -462 82 -462 0 net=4785
rlabel metal2 779 -462 779 -462 0 net=6167
rlabel metal2 121 -464 121 -464 0 net=1193
rlabel metal2 233 -464 233 -464 0 net=1262
rlabel metal2 485 -464 485 -464 0 net=3205
rlabel metal2 597 -464 597 -464 0 net=4049
rlabel metal2 702 -464 702 -464 0 net=4803
rlabel metal2 744 -464 744 -464 0 net=5051
rlabel metal2 821 -464 821 -464 0 net=5963
rlabel metal2 128 -466 128 -466 0 net=2017
rlabel metal2 177 -466 177 -466 0 net=3133
rlabel metal2 520 -466 520 -466 0 net=3787
rlabel metal2 604 -466 604 -466 0 net=4161
rlabel metal2 681 -466 681 -466 0 net=4693
rlabel metal2 835 -466 835 -466 0 net=6089
rlabel metal2 96 -468 96 -468 0 net=475
rlabel metal2 135 -468 135 -468 0 net=3289
rlabel metal2 338 -468 338 -468 0 net=2395
rlabel metal2 464 -468 464 -468 0 net=5125
rlabel metal2 856 -468 856 -468 0 net=6153
rlabel metal2 96 -470 96 -470 0 net=1647
rlabel metal2 212 -470 212 -470 0 net=3619
rlabel metal2 464 -470 464 -470 0 net=2855
rlabel metal2 534 -470 534 -470 0 net=1657
rlabel metal2 607 -470 607 -470 0 net=4417
rlabel metal2 793 -470 793 -470 0 net=5357
rlabel metal2 863 -470 863 -470 0 net=6359
rlabel metal2 156 -472 156 -472 0 net=2789
rlabel metal2 471 -472 471 -472 0 net=3527
rlabel metal2 548 -472 548 -472 0 net=2683
rlabel metal2 758 -472 758 -472 0 net=5391
rlabel metal2 877 -472 877 -472 0 net=6407
rlabel metal2 149 -474 149 -474 0 net=2381
rlabel metal2 509 -474 509 -474 0 net=4923
rlabel metal2 212 -476 212 -476 0 net=2107
rlabel metal2 516 -476 516 -476 0 net=5557
rlabel metal2 2 -478 2 -478 0 net=2487
rlabel metal2 520 -478 520 -478 0 net=4190
rlabel metal2 2 -480 2 -480 0 net=4843
rlabel metal2 233 -480 233 -480 0 net=1201
rlabel metal2 261 -480 261 -480 0 net=2919
rlabel metal2 572 -480 572 -480 0 net=6139
rlabel metal2 124 -482 124 -482 0 net=3825
rlabel metal2 604 -482 604 -482 0 net=4367
rlabel metal2 240 -484 240 -484 0 net=2027
rlabel metal2 611 -484 611 -484 0 net=4241
rlabel metal2 254 -486 254 -486 0 net=3421
rlabel metal2 618 -486 618 -486 0 net=6487
rlabel metal2 205 -488 205 -488 0 net=3989
rlabel metal2 569 -488 569 -488 0 net=4467
rlabel metal2 621 -488 621 -488 0 net=7586
rlabel metal2 289 -490 289 -490 0 net=3573
rlabel metal2 569 -490 569 -490 0 net=6714
rlabel metal2 345 -492 345 -492 0 net=1737
rlabel metal2 632 -492 632 -492 0 net=4681
rlabel metal2 842 -492 842 -492 0 net=6101
rlabel metal2 159 -494 159 -494 0 net=2329
rlabel metal2 436 -494 436 -494 0 net=3301
rlabel metal2 583 -494 583 -494 0 net=3903
rlabel metal2 394 -496 394 -496 0 net=3115
rlabel metal2 446 -496 446 -496 0 net=5283
rlabel metal2 646 -496 646 -496 0 net=4269
rlabel metal2 457 -498 457 -498 0 net=5641
rlabel metal2 457 -500 457 -500 0 net=3459
rlabel metal2 583 -500 583 -500 0 net=4031
rlabel metal2 660 -500 660 -500 0 net=4557
rlabel metal2 492 -502 492 -502 0 net=3019
rlabel metal2 565 -502 565 -502 0 net=4151
rlabel metal2 506 -504 506 -504 0 net=3649
rlabel metal2 282 -506 282 -506 0 net=1561
rlabel metal2 2 -517 2 -517 0 net=4844
rlabel metal2 149 -517 149 -517 0 net=3663
rlabel metal2 390 -517 390 -517 0 net=2635
rlabel metal2 411 -517 411 -517 0 net=4270
rlabel metal2 1087 -517 1087 -517 0 net=7261
rlabel metal2 1087 -517 1087 -517 0 net=7261
rlabel metal2 2 -519 2 -519 0 net=5655
rlabel metal2 425 -519 425 -519 0 net=93
rlabel metal2 509 -519 509 -519 0 net=7298
rlabel metal2 9 -521 9 -521 0 net=4266
rlabel metal2 159 -521 159 -521 0 net=5006
rlabel metal2 544 -521 544 -521 0 net=7266
rlabel metal2 9 -523 9 -523 0 net=4897
rlabel metal2 821 -523 821 -523 0 net=5305
rlabel metal2 16 -525 16 -525 0 net=4536
rlabel metal2 107 -525 107 -525 0 net=1700
rlabel metal2 177 -525 177 -525 0 net=3135
rlabel metal2 572 -525 572 -525 0 net=4956
rlabel metal2 58 -527 58 -527 0 net=3354
rlabel metal2 576 -527 576 -527 0 net=3904
rlabel metal2 989 -527 989 -527 0 net=6847
rlabel metal2 72 -529 72 -529 0 net=3562
rlabel metal2 177 -529 177 -529 0 net=1877
rlabel metal2 212 -529 212 -529 0 net=2108
rlabel metal2 579 -529 579 -529 0 net=7322
rlabel metal2 75 -531 75 -531 0 net=3620
rlabel metal2 429 -531 429 -531 0 net=3040
rlabel metal2 628 -531 628 -531 0 net=5946
rlabel metal2 79 -533 79 -533 0 net=2740
rlabel metal2 415 -533 415 -533 0 net=2783
rlabel metal2 443 -533 443 -533 0 net=2857
rlabel metal2 555 -533 555 -533 0 net=3813
rlabel metal2 646 -533 646 -533 0 net=6444
rlabel metal2 58 -535 58 -535 0 net=1913
rlabel metal2 86 -535 86 -535 0 net=1277
rlabel metal2 128 -535 128 -535 0 net=2489
rlabel metal2 317 -535 317 -535 0 net=1986
rlabel metal2 464 -535 464 -535 0 net=4242
rlabel metal2 786 -535 786 -535 0 net=6103
rlabel metal2 1017 -535 1017 -535 0 net=6923
rlabel metal2 86 -537 86 -537 0 net=3701
rlabel metal2 145 -537 145 -537 0 net=2089
rlabel metal2 240 -537 240 -537 0 net=2029
rlabel metal2 331 -537 331 -537 0 net=2320
rlabel metal2 331 -537 331 -537 0 net=2320
rlabel metal2 387 -537 387 -537 0 net=3650
rlabel metal2 667 -537 667 -537 0 net=7132
rlabel metal2 51 -539 51 -539 0 net=3557
rlabel metal2 674 -539 674 -539 0 net=4163
rlabel metal2 947 -539 947 -539 0 net=6409
rlabel metal2 1031 -539 1031 -539 0 net=6987
rlabel metal2 51 -541 51 -541 0 net=3789
rlabel metal2 674 -541 674 -541 0 net=5147
rlabel metal2 754 -541 754 -541 0 net=7212
rlabel metal2 121 -543 121 -543 0 net=1195
rlabel metal2 446 -543 446 -543 0 net=2986
rlabel metal2 828 -543 828 -543 0 net=6385
rlabel metal2 72 -545 72 -545 0 net=1375
rlabel metal2 135 -545 135 -545 0 net=1433
rlabel metal2 247 -545 247 -545 0 net=1526
rlabel metal2 481 -545 481 -545 0 net=4245
rlabel metal2 695 -545 695 -545 0 net=4207
rlabel metal2 730 -545 730 -545 0 net=4787
rlabel metal2 807 -545 807 -545 0 net=7325
rlabel metal2 135 -547 135 -547 0 net=3991
rlabel metal2 247 -547 247 -547 0 net=1463
rlabel metal2 520 -547 520 -547 0 net=4079
rlabel metal2 695 -547 695 -547 0 net=4419
rlabel metal2 772 -547 772 -547 0 net=5605
rlabel metal2 996 -547 996 -547 0 net=6903
rlabel metal2 1038 -547 1038 -547 0 net=7101
rlabel metal2 145 -549 145 -549 0 net=1560
rlabel metal2 250 -549 250 -549 0 net=1995
rlabel metal2 471 -549 471 -549 0 net=2382
rlabel metal2 551 -549 551 -549 0 net=5771
rlabel metal2 1059 -549 1059 -549 0 net=7457
rlabel metal2 37 -551 37 -551 0 net=2883
rlabel metal2 261 -551 261 -551 0 net=2920
rlabel metal2 555 -551 555 -551 0 net=3721
rlabel metal2 597 -551 597 -551 0 net=4021
rlabel metal2 723 -551 723 -551 0 net=6489
rlabel metal2 44 -553 44 -553 0 net=3373
rlabel metal2 632 -553 632 -553 0 net=5285
rlabel metal2 814 -553 814 -553 0 net=5623
rlabel metal2 940 -553 940 -553 0 net=7539
rlabel metal2 44 -555 44 -555 0 net=3733
rlabel metal2 436 -555 436 -555 0 net=3117
rlabel metal2 492 -555 492 -555 0 net=3281
rlabel metal2 583 -555 583 -555 0 net=4033
rlabel metal2 639 -555 639 -555 0 net=4051
rlabel metal2 723 -555 723 -555 0 net=5053
rlabel metal2 828 -555 828 -555 0 net=5359
rlabel metal2 940 -555 940 -555 0 net=6361
rlabel metal2 156 -557 156 -557 0 net=1933
rlabel metal2 205 -557 205 -557 0 net=1885
rlabel metal2 289 -557 289 -557 0 net=3574
rlabel metal2 422 -557 422 -557 0 net=5693
rlabel metal2 800 -557 800 -557 0 net=5393
rlabel metal2 114 -559 114 -559 0 net=2577
rlabel metal2 296 -559 296 -559 0 net=2751
rlabel metal2 492 -559 492 -559 0 net=3303
rlabel metal2 583 -559 583 -559 0 net=435
rlabel metal2 653 -559 653 -559 0 net=4153
rlabel metal2 835 -559 835 -559 0 net=5127
rlabel metal2 100 -561 100 -561 0 net=3579
rlabel metal2 152 -561 152 -561 0 net=305
rlabel metal2 338 -561 338 -561 0 net=2791
rlabel metal2 499 -561 499 -561 0 net=3529
rlabel metal2 604 -561 604 -561 0 net=5861
rlabel metal2 30 -563 30 -563 0 net=3915
rlabel metal2 401 -563 401 -563 0 net=1738
rlabel metal2 660 -563 660 -563 0 net=4369
rlabel metal2 835 -563 835 -563 0 net=5543
rlabel metal2 30 -565 30 -565 0 net=3207
rlabel metal2 513 -565 513 -565 0 net=3659
rlabel metal2 604 -565 604 -565 0 net=4001
rlabel metal2 842 -565 842 -565 0 net=5559
rlabel metal2 16 -567 16 -567 0 net=5105
rlabel metal2 856 -567 856 -567 0 net=6169
rlabel metal2 100 -569 100 -569 0 net=2183
rlabel metal2 261 -569 261 -569 0 net=1609
rlabel metal2 352 -569 352 -569 0 net=3173
rlabel metal2 513 -569 513 -569 0 net=3021
rlabel metal2 863 -569 863 -569 0 net=5643
rlabel metal2 954 -569 954 -569 0 net=6699
rlabel metal2 37 -571 37 -571 0 net=1251
rlabel metal2 254 -571 254 -571 0 net=3423
rlabel metal2 394 -571 394 -571 0 net=4383
rlabel metal2 870 -571 870 -571 0 net=5725
rlabel metal2 975 -571 975 -571 0 net=6373
rlabel metal2 191 -573 191 -573 0 net=1203
rlabel metal2 254 -573 254 -573 0 net=1563
rlabel metal2 394 -573 394 -573 0 net=1659
rlabel metal2 541 -573 541 -573 0 net=4244
rlabel metal2 877 -573 877 -573 0 net=5741
rlabel metal2 975 -573 975 -573 0 net=6805
rlabel metal2 233 -575 233 -575 0 net=2997
rlabel metal2 716 -575 716 -575 0 net=4683
rlabel metal2 898 -575 898 -575 0 net=5965
rlabel metal2 1010 -575 1010 -575 0 net=7563
rlabel metal2 107 -577 107 -577 0 net=2173
rlabel metal2 268 -579 268 -579 0 net=3827
rlabel metal2 268 -579 268 -579 0 net=3827
rlabel metal2 282 -579 282 -579 0 net=2439
rlabel metal2 457 -579 457 -579 0 net=3461
rlabel metal2 565 -579 565 -579 0 net=6027
rlabel metal2 919 -579 919 -579 0 net=6075
rlabel metal2 65 -581 65 -581 0 net=2251
rlabel metal2 457 -581 457 -581 0 net=6154
rlabel metal2 65 -583 65 -583 0 net=3290
rlabel metal2 523 -583 523 -583 0 net=3801
rlabel metal2 709 -583 709 -583 0 net=4805
rlabel metal2 751 -583 751 -583 0 net=5059
rlabel metal2 170 -585 170 -585 0 net=2019
rlabel metal2 373 -585 373 -585 0 net=2458
rlabel metal2 565 -585 565 -585 0 net=5493
rlabel metal2 170 -587 170 -587 0 net=1033
rlabel metal2 345 -587 345 -587 0 net=2331
rlabel metal2 681 -587 681 -587 0 net=4559
rlabel metal2 751 -587 751 -587 0 net=4761
rlabel metal2 198 -589 198 -589 0 net=2159
rlabel metal2 618 -589 618 -589 0 net=4469
rlabel metal2 345 -591 345 -591 0 net=2397
rlabel metal2 453 -591 453 -591 0 net=4275
rlabel metal2 758 -591 758 -591 0 net=6141
rlabel metal2 184 -593 184 -593 0 net=2201
rlabel metal2 618 -593 618 -593 0 net=6774
rlabel metal2 23 -595 23 -595 0 net=4078
rlabel metal2 744 -595 744 -595 0 net=4695
rlabel metal2 933 -595 933 -595 0 net=6091
rlabel metal2 23 -597 23 -597 0 net=1649
rlabel metal2 744 -597 744 -597 0 net=4925
rlabel metal2 933 -597 933 -597 0 net=6265
rlabel metal2 163 -599 163 -599 0 net=2685
rlabel metal2 334 -601 334 -601 0 net=5205
rlabel metal2 467 -603 467 -603 0 net=7181
rlabel metal2 548 -605 548 -605 0 net=703
rlabel metal2 23 -616 23 -616 0 net=1650
rlabel metal2 415 -616 415 -616 0 net=2792
rlabel metal2 453 -616 453 -616 0 net=4470
rlabel metal2 905 -616 905 -616 0 net=5494
rlabel metal2 1216 -616 1216 -616 0 net=6201
rlabel metal2 30 -618 30 -618 0 net=3209
rlabel metal2 30 -618 30 -618 0 net=3209
rlabel metal2 40 -618 40 -618 0 net=257
rlabel metal2 618 -618 618 -618 0 net=5148
rlabel metal2 716 -618 716 -618 0 net=4685
rlabel metal2 814 -618 814 -618 0 net=5625
rlabel metal2 961 -618 961 -618 0 net=7183
rlabel metal2 2 -620 2 -620 0 net=5657
rlabel metal2 702 -620 702 -620 0 net=4209
rlabel metal2 723 -620 723 -620 0 net=5055
rlabel metal2 961 -620 961 -620 0 net=5061
rlabel metal2 989 -620 989 -620 0 net=6849
rlabel metal2 2 -622 2 -622 0 net=6363
rlabel metal2 975 -622 975 -622 0 net=6807
rlabel metal2 44 -624 44 -624 0 net=3735
rlabel metal2 621 -624 621 -624 0 net=5887
rlabel metal2 996 -624 996 -624 0 net=6905
rlabel metal2 44 -626 44 -626 0 net=3916
rlabel metal2 352 -626 352 -626 0 net=3425
rlabel metal2 352 -626 352 -626 0 net=3425
rlabel metal2 380 -626 380 -626 0 net=3802
rlabel metal2 635 -626 635 -626 0 net=6092
rlabel metal2 1059 -626 1059 -626 0 net=7459
rlabel metal2 47 -628 47 -628 0 net=1886
rlabel metal2 229 -628 229 -628 0 net=1196
rlabel metal2 324 -628 324 -628 0 net=2031
rlabel metal2 387 -628 387 -628 0 net=852
rlabel metal2 726 -628 726 -628 0 net=6170
rlabel metal2 884 -628 884 -628 0 net=5773
rlabel metal2 1010 -628 1010 -628 0 net=7565
rlabel metal2 51 -630 51 -630 0 net=3790
rlabel metal2 460 -630 460 -630 0 net=279
rlabel metal2 649 -630 649 -630 0 net=6485
rlabel metal2 58 -632 58 -632 0 net=6104
rlabel metal2 821 -632 821 -632 0 net=5307
rlabel metal2 870 -632 870 -632 0 net=5727
rlabel metal2 891 -632 891 -632 0 net=5863
rlabel metal2 1031 -632 1031 -632 0 net=6989
rlabel metal2 51 -634 51 -634 0 net=2099
rlabel metal2 65 -634 65 -634 0 net=526
rlabel metal2 551 -634 551 -634 0 net=4164
rlabel metal2 898 -634 898 -634 0 net=5967
rlabel metal2 1038 -634 1038 -634 0 net=7103
rlabel metal2 65 -636 65 -636 0 net=2175
rlabel metal2 121 -636 121 -636 0 net=1377
rlabel metal2 331 -636 331 -636 0 net=2398
rlabel metal2 404 -636 404 -636 0 net=6635
rlabel metal2 1066 -636 1066 -636 0 net=7541
rlabel metal2 16 -638 16 -638 0 net=5106
rlabel metal2 121 -638 121 -638 0 net=1287
rlabel metal2 667 -638 667 -638 0 net=4247
rlabel metal2 730 -638 730 -638 0 net=4789
rlabel metal2 1045 -638 1045 -638 0 net=7327
rlabel metal2 1083 -638 1083 -638 0 net=7262
rlabel metal2 16 -640 16 -640 0 net=1337
rlabel metal2 226 -640 226 -640 0 net=2884
rlabel metal2 418 -640 418 -640 0 net=573
rlabel metal2 464 -640 464 -640 0 net=7213
rlabel metal2 75 -642 75 -642 0 net=6374
rlabel metal2 86 -644 86 -644 0 net=3703
rlabel metal2 247 -644 247 -644 0 net=1465
rlabel metal2 422 -644 422 -644 0 net=2858
rlabel metal2 464 -644 464 -644 0 net=3023
rlabel metal2 523 -644 523 -644 0 net=6490
rlabel metal2 37 -646 37 -646 0 net=4271
rlabel metal2 89 -646 89 -646 0 net=7495
rlabel metal2 100 -648 100 -648 0 net=2184
rlabel metal2 492 -648 492 -648 0 net=3305
rlabel metal2 541 -648 541 -648 0 net=4857
rlabel metal2 800 -648 800 -648 0 net=5395
rlabel metal2 912 -648 912 -648 0 net=6029
rlabel metal2 100 -650 100 -650 0 net=2399
rlabel metal2 408 -650 408 -650 0 net=2637
rlabel metal2 478 -650 478 -650 0 net=3137
rlabel metal2 544 -650 544 -650 0 net=4762
rlabel metal2 779 -650 779 -650 0 net=5695
rlabel metal2 947 -650 947 -650 0 net=6411
rlabel metal2 128 -652 128 -652 0 net=2490
rlabel metal2 289 -652 289 -652 0 net=2579
rlabel metal2 492 -652 492 -652 0 net=4371
rlabel metal2 709 -652 709 -652 0 net=4561
rlabel metal2 807 -652 807 -652 0 net=5287
rlabel metal2 912 -652 912 -652 0 net=6143
rlabel metal2 947 -652 947 -652 0 net=6925
rlabel metal2 93 -654 93 -654 0 net=1279
rlabel metal2 142 -654 142 -654 0 net=7177
rlabel metal2 61 -656 61 -656 0 net=3105
rlabel metal2 240 -656 240 -656 0 net=1434
rlabel metal2 502 -656 502 -656 0 net=6325
rlabel metal2 9 -658 9 -658 0 net=4898
rlabel metal2 93 -658 93 -658 0 net=2161
rlabel metal2 247 -658 247 -658 0 net=2441
rlabel metal2 289 -658 289 -658 0 net=2253
rlabel metal2 394 -658 394 -658 0 net=1661
rlabel metal2 520 -658 520 -658 0 net=5029
rlabel metal2 810 -658 810 -658 0 net=6853
rlabel metal2 9 -660 9 -660 0 net=5681
rlabel metal2 418 -660 418 -660 0 net=3233
rlabel metal2 548 -660 548 -660 0 net=3375
rlabel metal2 590 -660 590 -660 0 net=3559
rlabel metal2 632 -660 632 -660 0 net=4035
rlabel metal2 709 -660 709 -660 0 net=4927
rlabel metal2 821 -660 821 -660 0 net=6077
rlabel metal2 933 -660 933 -660 0 net=6267
rlabel metal2 23 -662 23 -662 0 net=5567
rlabel metal2 534 -662 534 -662 0 net=3463
rlabel metal2 576 -662 576 -662 0 net=3815
rlabel metal2 597 -662 597 -662 0 net=4023
rlabel metal2 632 -662 632 -662 0 net=7051
rlabel metal2 110 -664 110 -664 0 net=2415
rlabel metal2 534 -664 534 -664 0 net=3723
rlabel metal2 558 -664 558 -664 0 net=6317
rlabel metal2 145 -666 145 -666 0 net=4357
rlabel metal2 261 -666 261 -666 0 net=1611
rlabel metal2 296 -666 296 -666 0 net=2753
rlabel metal2 555 -666 555 -666 0 net=3385
rlabel metal2 597 -666 597 -666 0 net=3355
rlabel metal2 733 -666 733 -666 0 net=6565
rlabel metal2 198 -668 198 -668 0 net=1587
rlabel metal2 254 -668 254 -668 0 net=1565
rlabel metal2 275 -668 275 -668 0 net=3003
rlabel metal2 562 -668 562 -668 0 net=6386
rlabel metal2 278 -670 278 -670 0 net=2613
rlabel metal2 303 -670 303 -670 0 net=2021
rlabel metal2 317 -670 317 -670 0 net=1997
rlabel metal2 334 -670 334 -670 0 net=5415
rlabel metal2 954 -670 954 -670 0 net=6701
rlabel metal2 163 -672 163 -672 0 net=2687
rlabel metal2 457 -672 457 -672 0 net=6537
rlabel metal2 163 -674 163 -674 0 net=2091
rlabel metal2 268 -674 268 -674 0 net=3829
rlabel metal2 562 -674 562 -674 0 net=4696
rlabel metal2 772 -674 772 -674 0 net=5607
rlabel metal2 968 -674 968 -674 0 net=5129
rlabel metal2 191 -676 191 -676 0 net=1205
rlabel metal2 219 -676 219 -676 0 net=1253
rlabel metal2 310 -676 310 -676 0 net=3175
rlabel metal2 565 -676 565 -676 0 net=7165
rlabel metal2 177 -678 177 -678 0 net=1878
rlabel metal2 383 -678 383 -678 0 net=5747
rlabel metal2 177 -680 177 -680 0 net=3531
rlabel metal2 565 -680 565 -680 0 net=7225
rlabel metal2 149 -682 149 -682 0 net=3664
rlabel metal2 583 -682 583 -682 0 net=5919
rlabel metal2 842 -682 842 -682 0 net=5561
rlabel metal2 149 -684 149 -684 0 net=1935
rlabel metal2 184 -684 184 -684 0 net=1009
rlabel metal2 485 -684 485 -684 0 net=3661
rlabel metal2 583 -684 583 -684 0 net=7597
rlabel metal2 156 -686 156 -686 0 net=2785
rlabel metal2 506 -686 506 -686 0 net=3283
rlabel metal2 586 -686 586 -686 0 net=5399
rlabel metal2 863 -686 863 -686 0 net=5645
rlabel metal2 72 -688 72 -688 0 net=3193
rlabel metal2 628 -688 628 -688 0 net=5223
rlabel metal2 877 -688 877 -688 0 net=5743
rlabel metal2 72 -690 72 -690 0 net=1915
rlabel metal2 170 -690 170 -690 0 net=1035
rlabel metal2 429 -690 429 -690 0 net=4873
rlabel metal2 695 -690 695 -690 0 net=4421
rlabel metal2 828 -690 828 -690 0 net=5361
rlabel metal2 68 -692 68 -692 0 net=1959
rlabel metal2 114 -692 114 -692 0 net=3581
rlabel metal2 646 -692 646 -692 0 net=4081
rlabel metal2 114 -694 114 -694 0 net=2333
rlabel metal2 681 -694 681 -694 0 net=4277
rlabel metal2 737 -694 737 -694 0 net=4807
rlabel metal2 835 -694 835 -694 0 net=5545
rlabel metal2 373 -696 373 -696 0 net=3119
rlabel metal2 688 -696 688 -696 0 net=4385
rlabel metal2 233 -698 233 -698 0 net=2999
rlabel metal2 653 -698 653 -698 0 net=4155
rlabel metal2 793 -698 793 -698 0 net=5207
rlabel metal2 233 -700 233 -700 0 net=2202
rlabel metal2 383 -700 383 -700 0 net=4629
rlabel metal2 226 -702 226 -702 0 net=3177
rlabel metal2 446 -702 446 -702 0 net=4109
rlabel metal2 254 -704 254 -704 0 net=1591
rlabel metal2 639 -706 639 -706 0 net=4053
rlabel metal2 135 -708 135 -708 0 net=3993
rlabel metal2 135 -710 135 -710 0 net=4003
rlabel metal2 450 -712 450 -712 0 net=5021
rlabel metal2 450 -714 450 -714 0 net=1755
rlabel metal2 2 -725 2 -725 0 net=6364
rlabel metal2 131 -725 131 -725 0 net=3176
rlabel metal2 338 -725 338 -725 0 net=2032
rlabel metal2 464 -725 464 -725 0 net=3025
rlabel metal2 569 -725 569 -725 0 net=3464
rlabel metal2 586 -725 586 -725 0 net=4082
rlabel metal2 1136 -725 1136 -725 0 net=7167
rlabel metal2 1360 -725 1360 -725 0 net=6203
rlabel metal2 2 -727 2 -727 0 net=1961
rlabel metal2 89 -727 89 -727 0 net=282
rlabel metal2 198 -727 198 -727 0 net=1589
rlabel metal2 254 -727 254 -727 0 net=1592
rlabel metal2 737 -727 737 -727 0 net=4631
rlabel metal2 737 -727 737 -727 0 net=4631
rlabel metal2 828 -727 828 -727 0 net=4387
rlabel metal2 9 -729 9 -729 0 net=5682
rlabel metal2 726 -729 726 -729 0 net=6854
rlabel metal2 1143 -729 1143 -729 0 net=7179
rlabel metal2 9 -731 9 -731 0 net=2101
rlabel metal2 79 -731 79 -731 0 net=4359
rlabel metal2 254 -731 254 -731 0 net=3121
rlabel metal2 390 -731 390 -731 0 net=7598
rlabel metal2 16 -733 16 -733 0 net=1338
rlabel metal2 89 -733 89 -733 0 net=4278
rlabel metal2 705 -733 705 -733 0 net=7542
rlabel metal2 16 -735 16 -735 0 net=2951
rlabel metal2 401 -735 401 -735 0 net=5864
rlabel metal2 1017 -735 1017 -735 0 net=6269
rlabel metal2 1164 -735 1164 -735 0 net=7215
rlabel metal2 30 -737 30 -737 0 net=3210
rlabel metal2 156 -737 156 -737 0 net=2787
rlabel metal2 338 -737 338 -737 0 net=2581
rlabel metal2 422 -737 422 -737 0 net=2639
rlabel metal2 485 -737 485 -737 0 net=3662
rlabel metal2 611 -737 611 -737 0 net=3560
rlabel metal2 635 -737 635 -737 0 net=7226
rlabel metal2 1178 -737 1178 -737 0 net=7497
rlabel metal2 37 -739 37 -739 0 net=4272
rlabel metal2 390 -739 390 -739 0 net=5417
rlabel metal2 436 -739 436 -739 0 net=2755
rlabel metal2 495 -739 495 -739 0 net=3724
rlabel metal2 576 -739 576 -739 0 net=3387
rlabel metal2 646 -739 646 -739 0 net=4422
rlabel metal2 828 -739 828 -739 0 net=7351
rlabel metal2 37 -741 37 -741 0 net=2163
rlabel metal2 100 -741 100 -741 0 net=2400
rlabel metal2 576 -741 576 -741 0 net=4025
rlabel metal2 649 -741 649 -741 0 net=6078
rlabel metal2 905 -741 905 -741 0 net=5627
rlabel metal2 975 -741 975 -741 0 net=5775
rlabel metal2 1017 -741 1017 -741 0 net=6567
rlabel metal2 1080 -741 1080 -741 0 net=7329
rlabel metal2 51 -743 51 -743 0 net=1493
rlabel metal2 65 -745 65 -745 0 net=2177
rlabel metal2 100 -745 100 -745 0 net=1281
rlabel metal2 142 -745 142 -745 0 net=3107
rlabel metal2 163 -745 163 -745 0 net=2092
rlabel metal2 380 -745 380 -745 0 net=2595
rlabel metal2 443 -745 443 -745 0 net=7611
rlabel metal2 65 -747 65 -747 0 net=2589
rlabel metal2 289 -747 289 -747 0 net=2255
rlabel metal2 457 -747 457 -747 0 net=3831
rlabel metal2 649 -747 649 -747 0 net=6486
rlabel metal2 1185 -747 1185 -747 0 net=7567
rlabel metal2 86 -749 86 -749 0 net=6451
rlabel metal2 1094 -749 1094 -749 0 net=6809
rlabel metal2 1157 -749 1157 -749 0 net=7185
rlabel metal2 107 -751 107 -751 0 net=1937
rlabel metal2 170 -751 170 -751 0 net=3583
rlabel metal2 177 -751 177 -751 0 net=3533
rlabel metal2 590 -751 590 -751 0 net=3817
rlabel metal2 1101 -751 1101 -751 0 net=6851
rlabel metal2 142 -753 142 -753 0 net=1901
rlabel metal2 408 -753 408 -753 0 net=1663
rlabel metal2 502 -753 502 -753 0 net=4790
rlabel metal2 1108 -753 1108 -753 0 net=6907
rlabel metal2 149 -755 149 -755 0 net=3307
rlabel metal2 516 -755 516 -755 0 net=4137
rlabel metal2 709 -755 709 -755 0 net=4929
rlabel metal2 856 -755 856 -755 0 net=5309
rlabel metal2 912 -755 912 -755 0 net=6145
rlabel metal2 1115 -755 1115 -755 0 net=7053
rlabel metal2 170 -757 170 -757 0 net=3705
rlabel metal2 212 -757 212 -757 0 net=1207
rlabel metal2 299 -757 299 -757 0 net=5067
rlabel metal2 856 -757 856 -757 0 net=5749
rlabel metal2 1059 -757 1059 -757 0 net=6703
rlabel metal2 1122 -757 1122 -757 0 net=7105
rlabel metal2 44 -759 44 -759 0 net=5667
rlabel metal2 44 -761 44 -761 0 net=2119
rlabel metal2 415 -761 415 -761 0 net=4111
rlabel metal2 709 -761 709 -761 0 net=4211
rlabel metal2 723 -761 723 -761 0 net=4563
rlabel metal2 765 -761 765 -761 0 net=4687
rlabel metal2 961 -761 961 -761 0 net=5063
rlabel metal2 33 -763 33 -763 0 net=4771
rlabel metal2 765 -763 765 -763 0 net=6637
rlabel metal2 114 -765 114 -765 0 net=2335
rlabel metal2 702 -765 702 -765 0 net=4249
rlabel metal2 730 -765 730 -765 0 net=5968
rlabel metal2 114 -767 114 -767 0 net=1887
rlabel metal2 506 -767 506 -767 0 net=3195
rlabel metal2 639 -767 639 -767 0 net=3995
rlabel metal2 128 -769 128 -769 0 net=7485
rlabel metal2 135 -771 135 -771 0 net=4005
rlabel metal2 653 -771 653 -771 0 net=6593
rlabel metal2 75 -773 75 -773 0 net=1487
rlabel metal2 191 -773 191 -773 0 net=2225
rlabel metal2 352 -773 352 -773 0 net=3426
rlabel metal2 457 -773 457 -773 0 net=3075
rlabel metal2 513 -773 513 -773 0 net=7460
rlabel metal2 121 -775 121 -775 0 net=1289
rlabel metal2 198 -775 198 -775 0 net=1011
rlabel metal2 359 -775 359 -775 0 net=3179
rlabel metal2 478 -775 478 -775 0 net=3357
rlabel metal2 656 -775 656 -775 0 net=6990
rlabel metal2 121 -777 121 -777 0 net=2767
rlabel metal2 870 -777 870 -777 0 net=5397
rlabel metal2 1024 -777 1024 -777 0 net=5131
rlabel metal2 177 -779 177 -779 0 net=2401
rlabel metal2 359 -779 359 -779 0 net=4221
rlabel metal2 432 -779 432 -779 0 net=6043
rlabel metal2 205 -781 205 -781 0 net=1467
rlabel metal2 366 -781 366 -781 0 net=1757
rlabel metal2 492 -781 492 -781 0 net=4373
rlabel metal2 184 -783 184 -783 0 net=1037
rlabel metal2 492 -783 492 -783 0 net=4054
rlabel metal2 870 -783 870 -783 0 net=5697
rlabel metal2 947 -783 947 -783 0 net=6927
rlabel metal2 184 -785 184 -785 0 net=2023
rlabel metal2 520 -785 520 -785 0 net=3234
rlabel metal2 569 -785 569 -785 0 net=6529
rlabel metal2 23 -787 23 -787 0 net=5568
rlabel metal2 523 -787 523 -787 0 net=5608
rlabel metal2 926 -787 926 -787 0 net=5647
rlabel metal2 954 -787 954 -787 0 net=5745
rlabel metal2 219 -789 219 -789 0 net=1567
rlabel metal2 275 -789 275 -789 0 net=3005
rlabel metal2 527 -789 527 -789 0 net=3285
rlabel metal2 961 -789 961 -789 0 net=6031
rlabel metal2 261 -791 261 -791 0 net=1613
rlabel metal2 527 -791 527 -791 0 net=4859
rlabel metal2 877 -791 877 -791 0 net=5547
rlabel metal2 583 -793 583 -793 0 net=5511
rlabel metal2 268 -795 268 -795 0 net=1255
rlabel metal2 499 -795 499 -795 0 net=3519
rlabel metal2 586 -795 586 -795 0 net=6747
rlabel metal2 268 -797 268 -797 0 net=2417
rlabel metal2 590 -797 590 -797 0 net=3737
rlabel metal2 653 -797 653 -797 0 net=5455
rlabel metal2 849 -797 849 -797 0 net=5289
rlabel metal2 898 -797 898 -797 0 net=5563
rlabel metal2 163 -799 163 -799 0 net=1319
rlabel metal2 656 -799 656 -799 0 net=6187
rlabel metal2 387 -801 387 -801 0 net=327
rlabel metal2 429 -801 429 -801 0 net=2337
rlabel metal2 919 -801 919 -801 0 net=5889
rlabel metal2 429 -803 429 -803 0 net=6591
rlabel metal2 597 -805 597 -805 0 net=5659
rlabel metal2 688 -805 688 -805 0 net=4157
rlabel metal2 814 -805 814 -805 0 net=5057
rlabel metal2 884 -805 884 -805 0 net=5729
rlabel metal2 58 -807 58 -807 0 net=6963
rlabel metal2 702 -807 702 -807 0 net=5416
rlabel metal2 58 -809 58 -809 0 net=1917
rlabel metal2 404 -809 404 -809 0 net=6297
rlabel metal2 779 -809 779 -809 0 net=4809
rlabel metal2 72 -811 72 -811 0 net=1895
rlabel metal2 471 -811 471 -811 0 net=3001
rlabel metal2 800 -811 800 -811 0 net=5031
rlabel metal2 863 -811 863 -811 0 net=5363
rlabel metal2 317 -813 317 -813 0 net=2689
rlabel metal2 604 -813 604 -813 0 net=5023
rlabel metal2 842 -813 842 -813 0 net=5225
rlabel metal2 226 -815 226 -815 0 net=2151
rlabel metal2 548 -815 548 -815 0 net=3377
rlabel metal2 667 -815 667 -815 0 net=4875
rlabel metal2 835 -815 835 -815 0 net=5209
rlabel metal2 226 -817 226 -817 0 net=2443
rlabel metal2 541 -817 541 -817 0 net=3139
rlabel metal2 660 -817 660 -817 0 net=4037
rlabel metal2 807 -817 807 -817 0 net=5187
rlabel metal2 247 -819 247 -819 0 net=1379
rlabel metal2 509 -819 509 -819 0 net=3011
rlabel metal2 562 -819 562 -819 0 net=3729
rlabel metal2 758 -819 758 -819 0 net=5401
rlabel metal2 324 -821 324 -821 0 net=1999
rlabel metal2 562 -821 562 -821 0 net=455
rlabel metal2 758 -821 758 -821 0 net=6412
rlabel metal2 296 -823 296 -823 0 net=2615
rlabel metal2 1031 -823 1031 -823 0 net=6319
rlabel metal2 296 -825 296 -825 0 net=6538
rlabel metal2 432 -827 432 -827 0 net=6079
rlabel metal2 1038 -827 1038 -827 0 net=6327
rlabel metal2 772 -829 772 -829 0 net=5921
rlabel metal2 310 -831 310 -831 0 net=2697
rlabel metal2 16 -842 16 -842 0 net=2952
rlabel metal2 649 -842 649 -842 0 net=3002
rlabel metal2 824 -842 824 -842 0 net=7498
rlabel metal2 1416 -842 1416 -842 0 net=6205
rlabel metal2 16 -844 16 -844 0 net=1919
rlabel metal2 68 -844 68 -844 0 net=2582
rlabel metal2 390 -844 390 -844 0 net=2338
rlabel metal2 961 -844 961 -844 0 net=6033
rlabel metal2 26 -846 26 -846 0 net=2120
rlabel metal2 58 -846 58 -846 0 net=1321
rlabel metal2 170 -846 170 -846 0 net=3706
rlabel metal2 439 -846 439 -846 0 net=6592
rlabel metal2 30 -848 30 -848 0 net=2178
rlabel metal2 124 -848 124 -848 0 net=6594
rlabel metal2 30 -850 30 -850 0 net=4113
rlabel metal2 425 -850 425 -850 0 net=4158
rlabel metal2 828 -850 828 -850 0 net=7168
rlabel metal2 33 -852 33 -852 0 net=5512
rlabel metal2 961 -852 961 -852 0 net=5777
rlabel metal2 1143 -852 1143 -852 0 net=7331
rlabel metal2 37 -854 37 -854 0 net=2164
rlabel metal2 537 -854 537 -854 0 net=4026
rlabel metal2 586 -854 586 -854 0 net=5746
rlabel metal2 1129 -854 1129 -854 0 net=5132
rlabel metal2 37 -856 37 -856 0 net=1495
rlabel metal2 72 -856 72 -856 0 net=2024
rlabel metal2 198 -856 198 -856 0 net=1012
rlabel metal2 443 -856 443 -856 0 net=2256
rlabel metal2 544 -856 544 -856 0 net=3196
rlabel metal2 653 -856 653 -856 0 net=4810
rlabel metal2 898 -856 898 -856 0 net=5649
rlabel metal2 947 -856 947 -856 0 net=5669
rlabel metal2 1010 -856 1010 -856 0 net=6189
rlabel metal2 44 -858 44 -858 0 net=4633
rlabel metal2 758 -858 758 -858 0 net=7180
rlabel metal2 51 -860 51 -860 0 net=3201
rlabel metal2 205 -860 205 -860 0 net=1468
rlabel metal2 618 -860 618 -860 0 net=5564
rlabel metal2 1052 -860 1052 -860 0 net=5969
rlabel metal2 65 -862 65 -862 0 net=2591
rlabel metal2 79 -862 79 -862 0 net=4361
rlabel metal2 611 -862 611 -862 0 net=3389
rlabel metal2 625 -862 625 -862 0 net=6908
rlabel metal2 65 -864 65 -864 0 net=1282
rlabel metal2 121 -864 121 -864 0 net=2769
rlabel metal2 443 -864 443 -864 0 net=4139
rlabel metal2 702 -864 702 -864 0 net=5922
rlabel metal2 1164 -864 1164 -864 0 net=7055
rlabel metal2 79 -866 79 -866 0 net=3359
rlabel metal2 485 -866 485 -866 0 net=2757
rlabel metal2 565 -866 565 -866 0 net=6270
rlabel metal2 86 -868 86 -868 0 net=5277
rlabel metal2 856 -868 856 -868 0 net=5751
rlabel metal2 1003 -868 1003 -868 0 net=6147
rlabel metal2 1059 -868 1059 -868 0 net=7487
rlabel metal2 9 -870 9 -870 0 net=2102
rlabel metal2 89 -870 89 -870 0 net=3584
rlabel metal2 380 -870 380 -870 0 net=2597
rlabel metal2 471 -870 471 -870 0 net=2691
rlabel metal2 506 -870 506 -870 0 net=3286
rlabel metal2 968 -870 968 -870 0 net=6329
rlabel metal2 1087 -870 1087 -870 0 net=6749
rlabel metal2 2 -872 2 -872 0 net=1963
rlabel metal2 331 -872 331 -872 0 net=2617
rlabel metal2 397 -872 397 -872 0 net=3996
rlabel metal2 23 -874 23 -874 0 net=5507
rlabel metal2 982 -874 982 -874 0 net=5731
rlabel metal2 23 -876 23 -876 0 net=3095
rlabel metal2 509 -876 509 -876 0 net=3730
rlabel metal2 674 -876 674 -876 0 net=6299
rlabel metal2 93 -878 93 -878 0 net=2123
rlabel metal2 233 -878 233 -878 0 net=1209
rlabel metal2 233 -878 233 -878 0 net=1209
rlabel metal2 240 -878 240 -878 0 net=2788
rlabel metal2 408 -878 408 -878 0 net=1665
rlabel metal2 569 -878 569 -878 0 net=6852
rlabel metal2 100 -880 100 -880 0 net=3521
rlabel metal2 572 -880 572 -880 0 net=5517
rlabel metal2 761 -880 761 -880 0 net=5759
rlabel metal2 1017 -880 1017 -880 0 net=6569
rlabel metal2 121 -882 121 -882 0 net=4711
rlabel metal2 688 -882 688 -882 0 net=6965
rlabel metal2 131 -884 131 -884 0 net=7569
rlabel metal2 152 -886 152 -886 0 net=6215
rlabel metal2 1017 -886 1017 -886 0 net=6321
rlabel metal2 156 -888 156 -888 0 net=3109
rlabel metal2 369 -888 369 -888 0 net=2095
rlabel metal2 422 -888 422 -888 0 net=5419
rlabel metal2 478 -888 478 -888 0 net=4688
rlabel metal2 1031 -888 1031 -888 0 net=6081
rlabel metal2 2 -890 2 -890 0 net=2599
rlabel metal2 499 -890 499 -890 0 net=3818
rlabel metal2 1031 -890 1031 -890 0 net=6453
rlabel metal2 156 -892 156 -892 0 net=1425
rlabel metal2 723 -892 723 -892 0 net=4565
rlabel metal2 765 -892 765 -892 0 net=6639
rlabel metal2 1080 -892 1080 -892 0 net=6705
rlabel metal2 89 -894 89 -894 0 net=6943
rlabel metal2 131 -896 131 -896 0 net=4851
rlabel metal2 730 -896 730 -896 0 net=4877
rlabel metal2 786 -896 786 -896 0 net=5227
rlabel metal2 919 -896 919 -896 0 net=5891
rlabel metal2 163 -898 163 -898 0 net=1291
rlabel metal2 198 -898 198 -898 0 net=1301
rlabel metal2 254 -898 254 -898 0 net=3122
rlabel metal2 611 -898 611 -898 0 net=6928
rlabel metal2 114 -900 114 -900 0 net=1889
rlabel metal2 205 -900 205 -900 0 net=1897
rlabel metal2 296 -900 296 -900 0 net=1038
rlabel metal2 632 -900 632 -900 0 net=3833
rlabel metal2 695 -900 695 -900 0 net=4251
rlabel metal2 765 -900 765 -900 0 net=5025
rlabel metal2 807 -900 807 -900 0 net=5403
rlabel metal2 919 -900 919 -900 0 net=5549
rlabel metal2 1094 -900 1094 -900 0 net=5064
rlabel metal2 107 -902 107 -902 0 net=1939
rlabel metal2 170 -902 170 -902 0 net=2445
rlabel metal2 569 -902 569 -902 0 net=4011
rlabel metal2 646 -902 646 -902 0 net=6949
rlabel metal2 1094 -902 1094 -902 0 net=6811
rlabel metal2 107 -904 107 -904 0 net=4223
rlabel metal2 590 -904 590 -904 0 net=3739
rlabel metal2 653 -904 653 -904 0 net=5398
rlabel metal2 1150 -904 1150 -904 0 net=7353
rlabel metal2 177 -906 177 -906 0 net=1257
rlabel metal2 282 -906 282 -906 0 net=1590
rlabel metal2 345 -906 345 -906 0 net=3465
rlabel metal2 614 -906 614 -906 0 net=5683
rlabel metal2 996 -906 996 -906 0 net=6045
rlabel metal2 1185 -906 1185 -906 0 net=7187
rlabel metal2 180 -908 180 -908 0 net=2336
rlabel metal2 702 -908 702 -908 0 net=5211
rlabel metal2 863 -908 863 -908 0 net=5629
rlabel metal2 1024 -908 1024 -908 0 net=6531
rlabel metal2 1185 -908 1185 -908 0 net=7613
rlabel metal2 184 -910 184 -910 0 net=2459
rlabel metal2 709 -910 709 -910 0 net=4213
rlabel metal2 751 -910 751 -910 0 net=4773
rlabel metal2 807 -910 807 -910 0 net=5033
rlabel metal2 870 -910 870 -910 0 net=5699
rlabel metal2 212 -912 212 -912 0 net=2227
rlabel metal2 513 -912 513 -912 0 net=5251
rlabel metal2 870 -912 870 -912 0 net=4389
rlabel metal2 212 -914 212 -914 0 net=135
rlabel metal2 555 -914 555 -914 0 net=3027
rlabel metal2 656 -914 656 -914 0 net=5310
rlabel metal2 219 -916 219 -916 0 net=1569
rlabel metal2 299 -916 299 -916 0 net=1767
rlabel metal2 450 -916 450 -916 0 net=3007
rlabel metal2 562 -916 562 -916 0 net=2053
rlabel metal2 772 -916 772 -916 0 net=7216
rlabel metal2 219 -918 219 -918 0 net=1247
rlabel metal2 527 -918 527 -918 0 net=4861
rlabel metal2 775 -918 775 -918 0 net=5095
rlabel metal2 247 -920 247 -920 0 net=1381
rlabel metal2 261 -920 261 -920 0 net=1615
rlabel metal2 282 -920 282 -920 0 net=1717
rlabel metal2 450 -920 450 -920 0 net=7019
rlabel metal2 247 -922 247 -922 0 net=1039
rlabel metal2 261 -924 261 -924 0 net=1759
rlabel metal2 373 -924 373 -924 0 net=3181
rlabel metal2 576 -924 576 -924 0 net=5157
rlabel metal2 667 -924 667 -924 0 net=4039
rlabel metal2 709 -924 709 -924 0 net=7568
rlabel metal2 226 -926 226 -926 0 net=2444
rlabel metal2 436 -926 436 -926 0 net=3013
rlabel metal2 597 -926 597 -926 0 net=5661
rlabel metal2 135 -928 135 -928 0 net=1489
rlabel metal2 268 -928 268 -928 0 net=2419
rlabel metal2 352 -928 352 -928 0 net=2403
rlabel metal2 541 -928 541 -928 0 net=5058
rlabel metal2 135 -930 135 -930 0 net=2261
rlabel metal2 548 -930 548 -930 0 net=3141
rlabel metal2 639 -930 639 -930 0 net=4007
rlabel metal2 716 -930 716 -930 0 net=4374
rlabel metal2 142 -932 142 -932 0 net=1903
rlabel metal2 457 -932 457 -932 0 net=3077
rlabel metal2 604 -932 604 -932 0 net=3379
rlabel metal2 688 -932 688 -932 0 net=6685
rlabel metal2 142 -934 142 -934 0 net=1535
rlabel metal2 719 -934 719 -934 0 net=6913
rlabel metal2 149 -936 149 -936 0 net=3309
rlabel metal2 534 -936 534 -936 0 net=3535
rlabel metal2 744 -936 744 -936 0 net=4931
rlabel metal2 793 -936 793 -936 0 net=5457
rlabel metal2 268 -938 268 -938 0 net=1443
rlabel metal2 534 -938 534 -938 0 net=7429
rlabel metal2 289 -940 289 -940 0 net=2001
rlabel metal2 457 -940 457 -940 0 net=2641
rlabel metal2 793 -940 793 -940 0 net=5189
rlabel metal2 849 -940 849 -940 0 net=5291
rlabel metal2 310 -942 310 -942 0 net=2699
rlabel metal2 464 -942 464 -942 0 net=3755
rlabel metal2 821 -942 821 -942 0 net=5069
rlabel metal2 877 -942 877 -942 0 net=5365
rlabel metal2 75 -944 75 -944 0 net=2735
rlabel metal2 317 -944 317 -944 0 net=2153
rlabel metal2 821 -944 821 -944 0 net=7106
rlabel metal2 9 -946 9 -946 0 net=3147
rlabel metal2 324 -946 324 -946 0 net=1233
rlabel metal2 128 -948 128 -948 0 net=5467
rlabel metal2 2 -959 2 -959 0 net=2600
rlabel metal2 152 -959 152 -959 0 net=529
rlabel metal2 485 -959 485 -959 0 net=2693
rlabel metal2 485 -959 485 -959 0 net=2693
rlabel metal2 502 -959 502 -959 0 net=4040
rlabel metal2 688 -959 688 -959 0 net=5550
rlabel metal2 929 -959 929 -959 0 net=7547
rlabel metal2 1437 -959 1437 -959 0 net=6207
rlabel metal2 5 -961 5 -961 0 net=2154
rlabel metal2 541 -961 541 -961 0 net=6991
rlabel metal2 9 -963 9 -963 0 net=3148
rlabel metal2 548 -963 548 -963 0 net=3078
rlabel metal2 719 -963 719 -963 0 net=7189
rlabel metal2 16 -965 16 -965 0 net=1920
rlabel metal2 103 -965 103 -965 0 net=3545
rlabel metal2 744 -965 744 -965 0 net=5732
rlabel metal2 1136 -965 1136 -965 0 net=7021
rlabel metal2 16 -967 16 -967 0 net=1941
rlabel metal2 558 -967 558 -967 0 net=5228
rlabel metal2 863 -967 863 -967 0 net=5631
rlabel metal2 1143 -967 1143 -967 0 net=7333
rlabel metal2 30 -969 30 -969 0 net=4114
rlabel metal2 565 -969 565 -969 0 net=6300
rlabel metal2 1073 -969 1073 -969 0 net=6951
rlabel metal2 2 -971 2 -971 0 net=131
rlabel metal2 33 -971 33 -971 0 net=4862
rlabel metal2 866 -971 866 -971 0 net=6330
rlabel metal2 1087 -971 1087 -971 0 net=6751
rlabel metal2 44 -973 44 -973 0 net=4634
rlabel metal2 320 -973 320 -973 0 net=1847
rlabel metal2 502 -973 502 -973 0 net=7279
rlabel metal2 877 -973 877 -973 0 net=5367
rlabel metal2 1157 -973 1157 -973 0 net=7431
rlabel metal2 44 -975 44 -975 0 net=2447
rlabel metal2 198 -975 198 -975 0 net=2155
rlabel metal2 198 -975 198 -975 0 net=2155
rlabel metal2 201 -975 201 -975 0 net=1768
rlabel metal2 611 -975 611 -975 0 net=6515
rlabel metal2 37 -977 37 -977 0 net=1497
rlabel metal2 212 -977 212 -977 0 net=713
rlabel metal2 744 -977 744 -977 0 net=351
rlabel metal2 870 -977 870 -977 0 net=4391
rlabel metal2 912 -977 912 -977 0 net=5459
rlabel metal2 954 -977 954 -977 0 net=5761
rlabel metal2 1094 -977 1094 -977 0 net=6813
rlabel metal2 75 -979 75 -979 0 net=3834
rlabel metal2 667 -979 667 -979 0 net=4009
rlabel metal2 849 -979 849 -979 0 net=5293
rlabel metal2 961 -979 961 -979 0 net=5779
rlabel metal2 51 -981 51 -981 0 net=3203
rlabel metal2 695 -981 695 -981 0 net=4253
rlabel metal2 51 -983 51 -983 0 net=5468
rlabel metal2 968 -983 968 -983 0 net=6191
rlabel metal2 1052 -983 1052 -983 0 net=5971
rlabel metal2 1101 -983 1101 -983 0 net=6915
rlabel metal2 79 -985 79 -985 0 net=3360
rlabel metal2 572 -985 572 -985 0 net=6271
rlabel metal2 884 -985 884 -985 0 net=5753
rlabel metal2 975 -985 975 -985 0 net=5893
rlabel metal2 1115 -985 1115 -985 0 net=6945
rlabel metal2 23 -987 23 -987 0 net=3097
rlabel metal2 576 -987 576 -987 0 net=5159
rlabel metal2 933 -987 933 -987 0 net=5701
rlabel metal2 1150 -987 1150 -987 0 net=7355
rlabel metal2 1164 -987 1164 -987 0 net=7489
rlabel metal2 23 -989 23 -989 0 net=1445
rlabel metal2 282 -989 282 -989 0 net=1718
rlabel metal2 436 -989 436 -989 0 net=3015
rlabel metal2 702 -989 702 -989 0 net=5213
rlabel metal2 1003 -989 1003 -989 0 net=6149
rlabel metal2 1171 -989 1171 -989 0 net=7057
rlabel metal2 1171 -989 1171 -989 0 net=7057
rlabel metal2 1185 -989 1185 -989 0 net=7615
rlabel metal2 79 -991 79 -991 0 net=1249
rlabel metal2 254 -991 254 -991 0 net=1382
rlabel metal2 618 -991 618 -991 0 net=3391
rlabel metal2 709 -991 709 -991 0 net=5705
rlabel metal2 1192 -991 1192 -991 0 net=7188
rlabel metal2 114 -993 114 -993 0 net=1940
rlabel metal2 149 -993 149 -993 0 net=2601
rlabel metal2 436 -993 436 -993 0 net=5065
rlabel metal2 611 -993 611 -993 0 net=3433
rlabel metal2 856 -993 856 -993 0 net=5509
rlabel metal2 96 -995 96 -995 0 net=1685
rlabel metal2 121 -995 121 -995 0 net=1005
rlabel metal2 121 -995 121 -995 0 net=1005
rlabel metal2 124 -995 124 -995 0 net=715
rlabel metal2 723 -995 723 -995 0 net=4853
rlabel metal2 1017 -995 1017 -995 0 net=6323
rlabel metal2 156 -997 156 -997 0 net=1427
rlabel metal2 156 -997 156 -997 0 net=1427
rlabel metal2 177 -997 177 -997 0 net=1259
rlabel metal2 264 -997 264 -997 0 net=266
rlabel metal2 499 -997 499 -997 0 net=4911
rlabel metal2 891 -997 891 -997 0 net=5405
rlabel metal2 982 -997 982 -997 0 net=6217
rlabel metal2 1045 -997 1045 -997 0 net=6571
rlabel metal2 177 -999 177 -999 0 net=1303
rlabel metal2 268 -999 268 -999 0 net=1099
rlabel metal2 471 -999 471 -999 0 net=5421
rlabel metal2 1066 -999 1066 -999 0 net=6641
rlabel metal2 205 -1001 205 -1001 0 net=1899
rlabel metal2 219 -1001 219 -1001 0 net=1385
rlabel metal2 240 -1003 240 -1003 0 net=1235
rlabel metal2 331 -1003 331 -1003 0 net=3111
rlabel metal2 331 -1003 331 -1003 0 net=3111
rlabel metal2 338 -1003 338 -1003 0 net=2421
rlabel metal2 471 -1003 471 -1003 0 net=1667
rlabel metal2 513 -1003 513 -1003 0 net=3183
rlabel metal2 723 -1003 723 -1003 0 net=5325
rlabel metal2 1080 -1003 1080 -1003 0 net=6707
rlabel metal2 282 -1005 282 -1005 0 net=2771
rlabel metal2 478 -1005 478 -1005 0 net=6686
rlabel metal2 289 -1007 289 -1007 0 net=2003
rlabel metal2 341 -1007 341 -1007 0 net=2598
rlabel metal2 499 -1007 499 -1007 0 net=2629
rlabel metal2 555 -1007 555 -1007 0 net=3009
rlabel metal2 628 -1007 628 -1007 0 net=4566
rlabel metal2 747 -1007 747 -1007 0 net=4878
rlabel metal2 800 -1007 800 -1007 0 net=4775
rlabel metal2 835 -1007 835 -1007 0 net=5071
rlabel metal2 926 -1007 926 -1007 0 net=5685
rlabel metal2 1080 -1007 1080 -1007 0 net=6967
rlabel metal2 128 -1009 128 -1009 0 net=3793
rlabel metal2 747 -1009 747 -1009 0 net=6815
rlabel metal2 37 -1011 37 -1011 0 net=3881
rlabel metal2 142 -1011 142 -1011 0 net=1537
rlabel metal2 303 -1011 303 -1011 0 net=1965
rlabel metal2 506 -1011 506 -1011 0 net=2055
rlabel metal2 632 -1011 632 -1011 0 net=7587
rlabel metal2 86 -1013 86 -1013 0 net=310
rlabel metal2 306 -1013 306 -1013 0 net=2736
rlabel metal2 317 -1013 317 -1013 0 net=1573
rlabel metal2 513 -1013 513 -1013 0 net=3740
rlabel metal2 656 -1013 656 -1013 0 net=4331
rlabel metal2 814 -1013 814 -1013 0 net=5253
rlabel metal2 996 -1013 996 -1013 0 net=6047
rlabel metal2 86 -1015 86 -1015 0 net=2491
rlabel metal2 597 -1015 597 -1015 0 net=3143
rlabel metal2 751 -1015 751 -1015 0 net=4933
rlabel metal2 807 -1015 807 -1015 0 net=5035
rlabel metal2 989 -1015 989 -1015 0 net=6035
rlabel metal2 1031 -1015 1031 -1015 0 net=6455
rlabel metal2 40 -1017 40 -1017 0 net=2947
rlabel metal2 635 -1017 635 -1017 0 net=7607
rlabel metal2 310 -1019 310 -1019 0 net=2887
rlabel metal2 345 -1019 345 -1019 0 net=3467
rlabel metal2 730 -1019 730 -1019 0 net=4215
rlabel metal2 758 -1019 758 -1019 0 net=5519
rlabel metal2 345 -1021 345 -1021 0 net=2701
rlabel metal2 376 -1021 376 -1021 0 net=7570
rlabel metal2 352 -1023 352 -1023 0 net=1904
rlabel metal2 569 -1023 569 -1023 0 net=4013
rlabel metal2 765 -1023 765 -1023 0 net=5027
rlabel metal2 9 -1025 9 -1025 0 net=2217
rlabel metal2 569 -1025 569 -1025 0 net=3536
rlabel metal2 639 -1025 639 -1025 0 net=3381
rlabel metal2 793 -1025 793 -1025 0 net=5191
rlabel metal2 1024 -1025 1024 -1025 0 net=6533
rlabel metal2 261 -1027 261 -1027 0 net=1761
rlabel metal2 359 -1027 359 -1027 0 net=2229
rlabel metal2 677 -1027 677 -1027 0 net=4117
rlabel metal2 793 -1027 793 -1027 0 net=4279
rlabel metal2 898 -1027 898 -1027 0 net=5651
rlabel metal2 68 -1029 68 -1029 0 net=5083
rlabel metal2 905 -1029 905 -1029 0 net=5663
rlabel metal2 107 -1031 107 -1031 0 net=4225
rlabel metal2 366 -1031 366 -1031 0 net=5551
rlabel metal2 107 -1033 107 -1033 0 net=1071
rlabel metal2 842 -1033 842 -1033 0 net=5097
rlabel metal2 100 -1035 100 -1035 0 net=3523
rlabel metal2 100 -1037 100 -1037 0 net=6082
rlabel metal2 296 -1039 296 -1039 0 net=1571
rlabel metal2 947 -1039 947 -1039 0 net=5671
rlabel metal2 135 -1041 135 -1041 0 net=2263
rlabel metal2 366 -1041 366 -1041 0 net=1749
rlabel metal2 65 -1043 65 -1043 0 net=1435
rlabel metal2 369 -1043 369 -1043 0 net=7145
rlabel metal2 65 -1045 65 -1045 0 net=3633
rlabel metal2 520 -1045 520 -1045 0 net=2759
rlabel metal2 373 -1047 373 -1047 0 net=2096
rlabel metal2 401 -1047 401 -1047 0 net=2643
rlabel metal2 464 -1047 464 -1047 0 net=3757
rlabel metal2 828 -1047 828 -1047 0 net=5279
rlabel metal2 191 -1049 191 -1049 0 net=1891
rlabel metal2 429 -1049 429 -1049 0 net=2405
rlabel metal2 481 -1049 481 -1049 0 net=6687
rlabel metal2 163 -1051 163 -1051 0 net=1293
rlabel metal2 261 -1051 261 -1051 0 net=3291
rlabel metal2 492 -1051 492 -1051 0 net=3311
rlabel metal2 527 -1051 527 -1051 0 net=6483
rlabel metal2 163 -1053 163 -1053 0 net=2547
rlabel metal2 184 -1055 184 -1055 0 net=2461
rlabel metal2 492 -1055 492 -1055 0 net=4501
rlabel metal2 184 -1057 184 -1057 0 net=1041
rlabel metal2 380 -1057 380 -1057 0 net=2619
rlabel metal2 583 -1057 583 -1057 0 net=4363
rlabel metal2 233 -1059 233 -1059 0 net=1211
rlabel metal2 380 -1059 380 -1059 0 net=1821
rlabel metal2 527 -1059 527 -1059 0 net=4811
rlabel metal2 54 -1061 54 -1061 0 net=3059
rlabel metal2 534 -1061 534 -1061 0 net=5193
rlabel metal2 674 -1061 674 -1061 0 net=4713
rlabel metal2 443 -1063 443 -1063 0 net=4140
rlabel metal2 93 -1065 93 -1065 0 net=2125
rlabel metal2 583 -1065 583 -1065 0 net=2269
rlabel metal2 93 -1067 93 -1067 0 net=1045
rlabel metal2 590 -1067 590 -1067 0 net=3029
rlabel metal2 226 -1069 226 -1069 0 net=1491
rlabel metal2 226 -1071 226 -1071 0 net=1617
rlabel metal2 58 -1073 58 -1073 0 net=1323
rlabel metal2 58 -1075 58 -1075 0 net=2593
rlabel metal2 72 -1077 72 -1077 0 net=2083
rlabel metal2 2 -1088 2 -1088 0 net=5422
rlabel metal2 1241 -1088 1241 -1088 0 net=6947
rlabel metal2 1444 -1088 1444 -1088 0 net=6209
rlabel metal2 9 -1090 9 -1090 0 net=2219
rlabel metal2 404 -1090 404 -1090 0 net=2230
rlabel metal2 674 -1090 674 -1090 0 net=7022
rlabel metal2 1318 -1090 1318 -1090 0 net=7491
rlabel metal2 9 -1092 9 -1092 0 net=2665
rlabel metal2 37 -1092 37 -1092 0 net=1007
rlabel metal2 149 -1092 149 -1092 0 net=1618
rlabel metal2 247 -1092 247 -1092 0 net=1212
rlabel metal2 439 -1092 439 -1092 0 net=3312
rlabel metal2 527 -1092 527 -1092 0 net=5028
rlabel metal2 1213 -1092 1213 -1092 0 net=6753
rlabel metal2 1325 -1092 1325 -1092 0 net=7549
rlabel metal2 16 -1094 16 -1094 0 net=1943
rlabel metal2 16 -1094 16 -1094 0 net=1943
rlabel metal2 30 -1094 30 -1094 0 net=1373
rlabel metal2 569 -1094 569 -1094 0 net=7299
rlabel metal2 1339 -1094 1339 -1094 0 net=7617
rlabel metal2 54 -1096 54 -1096 0 net=3524
rlabel metal2 845 -1096 845 -1096 0 net=5235
rlabel metal2 1220 -1096 1220 -1096 0 net=6953
rlabel metal2 1311 -1096 1311 -1096 0 net=7433
rlabel metal2 58 -1098 58 -1098 0 net=2594
rlabel metal2 121 -1098 121 -1098 0 net=1539
rlabel metal2 408 -1098 408 -1098 0 net=2603
rlabel metal2 572 -1098 572 -1098 0 net=4010
rlabel metal2 786 -1098 786 -1098 0 net=7281
rlabel metal2 58 -1100 58 -1100 0 net=1305
rlabel metal2 212 -1100 212 -1100 0 net=1900
rlabel metal2 530 -1100 530 -1100 0 net=3010
rlabel metal2 628 -1100 628 -1100 0 net=5632
rlabel metal2 1192 -1100 1192 -1100 0 net=6643
rlabel metal2 75 -1102 75 -1102 0 net=5510
rlabel metal2 75 -1104 75 -1104 0 net=3204
rlabel metal2 667 -1104 667 -1104 0 net=3759
rlabel metal2 733 -1104 733 -1104 0 net=5339
rlabel metal2 79 -1106 79 -1106 0 net=1250
rlabel metal2 558 -1106 558 -1106 0 net=4118
rlabel metal2 863 -1106 863 -1106 0 net=7335
rlabel metal2 79 -1108 79 -1108 0 net=2127
rlabel metal2 471 -1108 471 -1108 0 net=1668
rlabel metal2 653 -1108 653 -1108 0 net=3185
rlabel metal2 684 -1108 684 -1108 0 net=6708
rlabel metal2 93 -1110 93 -1110 0 net=586
rlabel metal2 541 -1110 541 -1110 0 net=2621
rlabel metal2 576 -1110 576 -1110 0 net=5066
rlabel metal2 726 -1110 726 -1110 0 net=6324
rlabel metal2 1178 -1110 1178 -1110 0 net=6535
rlabel metal2 93 -1112 93 -1112 0 net=1499
rlabel metal2 177 -1112 177 -1112 0 net=2264
rlabel metal2 310 -1112 310 -1112 0 net=2889
rlabel metal2 450 -1112 450 -1112 0 net=3099
rlabel metal2 660 -1112 660 -1112 0 net=4093
rlabel metal2 765 -1112 765 -1112 0 net=6916
rlabel metal2 72 -1114 72 -1114 0 net=1345
rlabel metal2 205 -1114 205 -1114 0 net=2085
rlabel metal2 478 -1114 478 -1114 0 net=2694
rlabel metal2 492 -1114 492 -1114 0 net=5192
rlabel metal2 1087 -1114 1087 -1114 0 net=5895
rlabel metal2 1150 -1114 1150 -1114 0 net=7357
rlabel metal2 44 -1116 44 -1116 0 net=2449
rlabel metal2 499 -1116 499 -1116 0 net=4392
rlabel metal2 929 -1116 929 -1116 0 net=7334
rlabel metal2 44 -1118 44 -1118 0 net=1823
rlabel metal2 408 -1118 408 -1118 0 net=1849
rlabel metal2 457 -1118 457 -1118 0 net=2407
rlabel metal2 499 -1118 499 -1118 0 net=3435
rlabel metal2 632 -1118 632 -1118 0 net=6814
rlabel metal2 1290 -1118 1290 -1118 0 net=7191
rlabel metal2 23 -1120 23 -1120 0 net=1447
rlabel metal2 394 -1120 394 -1120 0 net=1893
rlabel metal2 457 -1120 457 -1120 0 net=2057
rlabel metal2 541 -1120 541 -1120 0 net=4254
rlabel metal2 23 -1122 23 -1122 0 net=1751
rlabel metal2 464 -1122 464 -1122 0 net=3293
rlabel metal2 695 -1122 695 -1122 0 net=3016
rlabel metal2 828 -1122 828 -1122 0 net=4715
rlabel metal2 954 -1122 954 -1122 0 net=5295
rlabel metal2 1227 -1122 1227 -1122 0 net=6817
rlabel metal2 1283 -1122 1283 -1122 0 net=7147
rlabel metal2 72 -1124 72 -1124 0 net=4014
rlabel metal2 821 -1124 821 -1124 0 net=4777
rlabel metal2 849 -1124 849 -1124 0 net=5255
rlabel metal2 1045 -1124 1045 -1124 0 net=5687
rlabel metal2 1171 -1124 1171 -1124 0 net=7059
rlabel metal2 96 -1126 96 -1126 0 net=1572
rlabel metal2 681 -1126 681 -1126 0 net=3383
rlabel metal2 712 -1126 712 -1126 0 net=6331
rlabel metal2 1199 -1126 1199 -1126 0 net=6689
rlabel metal2 100 -1128 100 -1128 0 net=4447
rlabel metal2 866 -1128 866 -1128 0 net=6572
rlabel metal2 117 -1130 117 -1130 0 net=6301
rlabel metal2 128 -1132 128 -1132 0 net=3883
rlabel metal2 464 -1132 464 -1132 0 net=6516
rlabel metal2 128 -1134 128 -1134 0 net=1411
rlabel metal2 716 -1134 716 -1134 0 net=3547
rlabel metal2 730 -1134 730 -1134 0 net=6150
rlabel metal2 1262 -1134 1262 -1134 0 net=6993
rlabel metal2 149 -1136 149 -1136 0 net=3145
rlabel metal2 702 -1136 702 -1136 0 net=3469
rlabel metal2 744 -1136 744 -1136 0 net=4502
rlabel metal2 870 -1136 870 -1136 0 net=6273
rlabel metal2 163 -1138 163 -1138 0 net=2549
rlabel metal2 212 -1138 212 -1138 0 net=994
rlabel metal2 688 -1138 688 -1138 0 net=3393
rlabel metal2 744 -1138 744 -1138 0 net=5368
rlabel metal2 163 -1140 163 -1140 0 net=4195
rlabel metal2 502 -1140 502 -1140 0 net=2760
rlabel metal2 1073 -1140 1073 -1140 0 net=5763
rlabel metal2 226 -1142 226 -1142 0 net=1325
rlabel metal2 282 -1142 282 -1142 0 net=2772
rlabel metal2 548 -1142 548 -1142 0 net=2631
rlabel metal2 600 -1142 600 -1142 0 net=5780
rlabel metal2 152 -1144 152 -1144 0 net=1309
rlabel metal2 289 -1144 289 -1144 0 net=3709
rlabel metal2 495 -1144 495 -1144 0 net=4623
rlabel metal2 905 -1144 905 -1144 0 net=5099
rlabel metal2 968 -1144 968 -1144 0 net=6193
rlabel metal2 1255 -1144 1255 -1144 0 net=7589
rlabel metal2 184 -1146 184 -1146 0 net=1043
rlabel metal2 296 -1146 296 -1146 0 net=1763
rlabel metal2 373 -1146 373 -1146 0 net=3047
rlabel metal2 649 -1146 649 -1146 0 net=3313
rlabel metal2 747 -1146 747 -1146 0 net=4854
rlabel metal2 1010 -1146 1010 -1146 0 net=5553
rlabel metal2 1066 -1146 1066 -1146 0 net=6457
rlabel metal2 103 -1148 103 -1148 0 net=1701
rlabel metal2 506 -1148 506 -1148 0 net=1161
rlabel metal2 800 -1148 800 -1148 0 net=4333
rlabel metal2 856 -1148 856 -1148 0 net=4913
rlabel metal2 933 -1148 933 -1148 0 net=5215
rlabel metal2 1080 -1148 1080 -1148 0 net=6969
rlabel metal2 5 -1150 5 -1150 0 net=4489
rlabel metal2 891 -1150 891 -1150 0 net=5073
rlabel metal2 961 -1150 961 -1150 0 net=5327
rlabel metal2 1017 -1150 1017 -1150 0 net=6219
rlabel metal2 5 -1152 5 -1152 0 net=7107
rlabel metal2 103 -1154 103 -1154 0 net=198
rlabel metal2 233 -1154 233 -1154 0 net=3061
rlabel metal2 534 -1154 534 -1154 0 net=5195
rlabel metal2 1017 -1154 1017 -1154 0 net=5973
rlabel metal2 1108 -1154 1108 -1154 0 net=6049
rlabel metal2 135 -1156 135 -1156 0 net=1437
rlabel metal2 240 -1156 240 -1156 0 net=1237
rlabel metal2 254 -1156 254 -1156 0 net=1260
rlabel metal2 534 -1156 534 -1156 0 net=2121
rlabel metal2 709 -1156 709 -1156 0 net=4813
rlabel metal2 912 -1156 912 -1156 0 net=5161
rlabel metal2 1031 -1156 1031 -1156 0 net=5665
rlabel metal2 40 -1158 40 -1158 0 net=1469
rlabel metal2 156 -1158 156 -1158 0 net=1429
rlabel metal2 240 -1158 240 -1158 0 net=2271
rlabel metal2 604 -1158 604 -1158 0 net=3031
rlabel metal2 747 -1158 747 -1158 0 net=5679
rlabel metal2 156 -1160 156 -1160 0 net=1133
rlabel metal2 481 -1160 481 -1160 0 net=2303
rlabel metal2 607 -1160 607 -1160 0 net=6484
rlabel metal2 261 -1162 261 -1162 0 net=4177
rlabel metal2 814 -1162 814 -1162 0 net=5037
rlabel metal2 1052 -1162 1052 -1162 0 net=5703
rlabel metal2 191 -1164 191 -1164 0 net=1295
rlabel metal2 303 -1164 303 -1164 0 net=4401
rlabel metal2 884 -1164 884 -1164 0 net=5755
rlabel metal2 142 -1166 142 -1166 0 net=1047
rlabel metal2 219 -1166 219 -1166 0 net=1387
rlabel metal2 310 -1166 310 -1166 0 net=2949
rlabel metal2 751 -1166 751 -1166 0 net=4217
rlabel metal2 807 -1166 807 -1166 0 net=4365
rlabel metal2 919 -1166 919 -1166 0 net=5461
rlabel metal2 1059 -1166 1059 -1166 0 net=5707
rlabel metal2 107 -1168 107 -1168 0 net=1073
rlabel metal2 219 -1168 219 -1168 0 net=2895
rlabel metal2 558 -1168 558 -1168 0 net=5787
rlabel metal2 107 -1170 107 -1170 0 net=2157
rlabel metal2 317 -1170 317 -1170 0 net=1575
rlabel metal2 401 -1170 401 -1170 0 net=2645
rlabel metal2 513 -1170 513 -1170 0 net=5569
rlabel metal2 180 -1172 180 -1172 0 net=4435
rlabel metal2 530 -1172 530 -1172 0 net=7527
rlabel metal2 198 -1174 198 -1174 0 net=1101
rlabel metal2 317 -1174 317 -1174 0 net=2005
rlabel metal2 341 -1174 341 -1174 0 net=1905
rlabel metal2 359 -1174 359 -1174 0 net=4227
rlabel metal2 1024 -1174 1024 -1174 0 net=5653
rlabel metal2 254 -1176 254 -1176 0 net=1263
rlabel metal2 555 -1176 555 -1176 0 net=6631
rlabel metal2 268 -1178 268 -1178 0 net=2463
rlabel metal2 565 -1178 565 -1178 0 net=4055
rlabel metal2 779 -1178 779 -1178 0 net=4935
rlabel metal2 975 -1178 975 -1178 0 net=5407
rlabel metal2 324 -1180 324 -1180 0 net=2703
rlabel metal2 359 -1180 359 -1180 0 net=2033
rlabel metal2 751 -1180 751 -1180 0 net=4985
rlabel metal2 975 -1180 975 -1180 0 net=5673
rlabel metal2 331 -1182 331 -1182 0 net=3113
rlabel metal2 793 -1182 793 -1182 0 net=4281
rlabel metal2 1003 -1182 1003 -1182 0 net=5521
rlabel metal2 331 -1184 331 -1184 0 net=1967
rlabel metal2 429 -1184 429 -1184 0 net=1527
rlabel metal2 758 -1184 758 -1184 0 net=7608
rlabel metal2 51 -1186 51 -1186 0 net=7435
rlabel metal2 345 -1188 345 -1188 0 net=3795
rlabel metal2 793 -1188 793 -1188 0 net=4603
rlabel metal2 996 -1188 996 -1188 0 net=6037
rlabel metal2 65 -1190 65 -1190 0 net=3635
rlabel metal2 947 -1190 947 -1190 0 net=5281
rlabel metal2 65 -1192 65 -1192 0 net=2493
rlabel metal2 387 -1192 387 -1192 0 net=2423
rlabel metal2 597 -1192 597 -1192 0 net=6709
rlabel metal2 86 -1194 86 -1194 0 net=1687
rlabel metal2 387 -1194 387 -1194 0 net=1593
rlabel metal2 625 -1194 625 -1194 0 net=4957
rlabel metal2 51 -1196 51 -1196 0 net=3621
rlabel metal2 898 -1196 898 -1196 0 net=5085
rlabel metal2 114 -1198 114 -1198 0 net=1492
rlabel metal2 551 -1200 551 -1200 0 net=4867
rlabel metal2 590 -1202 590 -1202 0 net=2797
rlabel metal2 2 -1213 2 -1213 0 net=1389
rlabel metal2 366 -1213 366 -1213 0 net=1576
rlabel metal2 607 -1213 607 -1213 0 net=5196
rlabel metal2 982 -1213 982 -1213 0 net=5237
rlabel metal2 982 -1213 982 -1213 0 net=5237
rlabel metal2 1017 -1213 1017 -1213 0 net=5975
rlabel metal2 1269 -1213 1269 -1213 0 net=6955
rlabel metal2 1304 -1213 1304 -1213 0 net=7193
rlabel metal2 1304 -1213 1304 -1213 0 net=7193
rlabel metal2 1360 -1213 1360 -1213 0 net=7551
rlabel metal2 1451 -1213 1451 -1213 0 net=6211
rlabel metal2 5 -1215 5 -1215 0 net=3114
rlabel metal2 793 -1215 793 -1215 0 net=4449
rlabel metal2 870 -1215 870 -1215 0 net=4625
rlabel metal2 1017 -1215 1017 -1215 0 net=5765
rlabel metal2 1269 -1215 1269 -1215 0 net=7061
rlabel metal2 30 -1217 30 -1217 0 net=1374
rlabel metal2 614 -1217 614 -1217 0 net=3032
rlabel metal2 628 -1217 628 -1217 0 net=3384
rlabel metal2 698 -1217 698 -1217 0 net=5216
rlabel metal2 1283 -1217 1283 -1217 0 net=7301
rlabel metal2 30 -1219 30 -1219 0 net=2605
rlabel metal2 632 -1219 632 -1219 0 net=5296
rlabel metal2 1272 -1219 1272 -1219 0 net=1
rlabel metal2 37 -1221 37 -1221 0 net=1008
rlabel metal2 261 -1221 261 -1221 0 net=1297
rlabel metal2 261 -1221 261 -1221 0 net=1297
rlabel metal2 289 -1221 289 -1221 0 net=3711
rlabel metal2 646 -1221 646 -1221 0 net=7618
rlabel metal2 37 -1223 37 -1223 0 net=1307
rlabel metal2 72 -1223 72 -1223 0 net=1541
rlabel metal2 124 -1223 124 -1223 0 net=1906
rlabel metal2 366 -1223 366 -1223 0 net=567
rlabel metal2 653 -1223 653 -1223 0 net=3101
rlabel metal2 44 -1225 44 -1225 0 net=1824
rlabel metal2 653 -1225 653 -1225 0 net=3471
rlabel metal2 719 -1225 719 -1225 0 net=6105
rlabel metal2 44 -1227 44 -1227 0 net=1501
rlabel metal2 100 -1227 100 -1227 0 net=1001
rlabel metal2 121 -1227 121 -1227 0 net=447
rlabel metal2 600 -1227 600 -1227 0 net=2957
rlabel metal2 667 -1227 667 -1227 0 net=3761
rlabel metal2 667 -1227 667 -1227 0 net=3761
rlabel metal2 684 -1227 684 -1227 0 net=7148
rlabel metal2 51 -1229 51 -1229 0 net=3623
rlabel metal2 138 -1229 138 -1229 0 net=2622
rlabel metal2 709 -1229 709 -1229 0 net=3636
rlabel metal2 751 -1229 751 -1229 0 net=4607
rlabel metal2 51 -1231 51 -1231 0 net=2265
rlabel metal2 432 -1231 432 -1231 0 net=2122
rlabel metal2 544 -1231 544 -1231 0 net=7599
rlabel metal2 58 -1233 58 -1233 0 net=2450
rlabel metal2 492 -1233 492 -1233 0 net=4366
rlabel metal2 915 -1233 915 -1233 0 net=5680
rlabel metal2 1150 -1233 1150 -1233 0 net=7359
rlabel metal2 75 -1235 75 -1235 0 net=1894
rlabel metal2 436 -1235 436 -1235 0 net=2646
rlabel metal2 520 -1235 520 -1235 0 net=3665
rlabel metal2 712 -1235 712 -1235 0 net=5704
rlabel metal2 1150 -1235 1150 -1235 0 net=6195
rlabel metal2 89 -1237 89 -1237 0 net=1326
rlabel metal2 289 -1237 289 -1237 0 net=1703
rlabel metal2 394 -1237 394 -1237 0 net=3884
rlabel metal2 534 -1237 534 -1237 0 net=2499
rlabel metal2 754 -1237 754 -1237 0 net=7434
rlabel metal2 142 -1239 142 -1239 0 net=1075
rlabel metal2 142 -1239 142 -1239 0 net=1075
rlabel metal2 149 -1239 149 -1239 0 net=3146
rlabel metal2 604 -1239 604 -1239 0 net=4825
rlabel metal2 940 -1239 940 -1239 0 net=5075
rlabel metal2 940 -1239 940 -1239 0 net=5075
rlabel metal2 1010 -1239 1010 -1239 0 net=5329
rlabel metal2 1080 -1239 1080 -1239 0 net=5757
rlabel metal2 1157 -1239 1157 -1239 0 net=6221
rlabel metal2 149 -1241 149 -1241 0 net=3797
rlabel metal2 352 -1241 352 -1241 0 net=1595
rlabel metal2 436 -1241 436 -1241 0 net=3601
rlabel metal2 548 -1241 548 -1241 0 net=5282
rlabel metal2 1010 -1241 1010 -1241 0 net=5523
rlabel metal2 1094 -1241 1094 -1241 0 net=6275
rlabel metal2 163 -1243 163 -1243 0 net=4196
rlabel metal2 163 -1243 163 -1243 0 net=4196
rlabel metal2 173 -1243 173 -1243 0 net=5666
rlabel metal2 177 -1245 177 -1245 0 net=1265
rlabel metal2 282 -1245 282 -1245 0 net=1044
rlabel metal2 446 -1245 446 -1245 0 net=6445
rlabel metal2 191 -1247 191 -1247 0 net=1049
rlabel metal2 310 -1247 310 -1247 0 net=2950
rlabel metal2 660 -1247 660 -1247 0 net=4095
rlabel metal2 765 -1247 765 -1247 0 net=5408
rlabel metal2 1038 -1247 1038 -1247 0 net=5555
rlabel metal2 1129 -1247 1129 -1247 0 net=5709
rlabel metal2 1178 -1247 1178 -1247 0 net=6333
rlabel metal2 170 -1249 170 -1249 0 net=1347
rlabel metal2 198 -1249 198 -1249 0 net=1102
rlabel metal2 695 -1249 695 -1249 0 net=3839
rlabel metal2 758 -1249 758 -1249 0 net=5831
rlabel metal2 1164 -1249 1164 -1249 0 net=7529
rlabel metal2 198 -1251 198 -1251 0 net=1765
rlabel metal2 310 -1251 310 -1251 0 net=4529
rlabel metal2 520 -1251 520 -1251 0 net=2321
rlabel metal2 604 -1251 604 -1251 0 net=3295
rlabel metal2 660 -1251 660 -1251 0 net=3395
rlabel metal2 758 -1251 758 -1251 0 net=4179
rlabel metal2 796 -1251 796 -1251 0 net=6536
rlabel metal2 205 -1253 205 -1253 0 net=2551
rlabel metal2 450 -1253 450 -1253 0 net=3063
rlabel metal2 527 -1253 527 -1253 0 net=6710
rlabel metal2 135 -1255 135 -1255 0 net=1471
rlabel metal2 212 -1255 212 -1255 0 net=2007
rlabel metal2 331 -1255 331 -1255 0 net=1969
rlabel metal2 464 -1255 464 -1255 0 net=2087
rlabel metal2 527 -1255 527 -1255 0 net=4337
rlabel metal2 548 -1255 548 -1255 0 net=1637
rlabel metal2 765 -1255 765 -1255 0 net=4229
rlabel metal2 842 -1255 842 -1255 0 net=6970
rlabel metal2 135 -1257 135 -1257 0 net=6644
rlabel metal2 1234 -1257 1234 -1257 0 net=6819
rlabel metal2 219 -1259 219 -1259 0 net=2897
rlabel metal2 621 -1259 621 -1259 0 net=7271
rlabel metal2 156 -1261 156 -1261 0 net=1135
rlabel metal2 226 -1261 226 -1261 0 net=2289
rlabel metal2 555 -1261 555 -1261 0 net=2633
rlabel metal2 681 -1261 681 -1261 0 net=6948
rlabel metal2 103 -1263 103 -1263 0 net=2993
rlabel metal2 233 -1263 233 -1263 0 net=1439
rlabel metal2 296 -1263 296 -1263 0 net=1851
rlabel metal2 457 -1263 457 -1263 0 net=2059
rlabel metal2 569 -1263 569 -1263 0 net=6050
rlabel metal2 1353 -1263 1353 -1263 0 net=7493
rlabel metal2 16 -1265 16 -1265 0 net=1945
rlabel metal2 576 -1265 576 -1265 0 net=2799
rlabel metal2 779 -1265 779 -1265 0 net=4219
rlabel metal2 807 -1265 807 -1265 0 net=4335
rlabel metal2 828 -1265 828 -1265 0 net=4779
rlabel metal2 845 -1265 845 -1265 0 net=5100
rlabel metal2 989 -1265 989 -1265 0 net=5257
rlabel metal2 1003 -1265 1003 -1265 0 net=6039
rlabel metal2 1164 -1265 1164 -1265 0 net=6303
rlabel metal2 1332 -1265 1332 -1265 0 net=7437
rlabel metal2 16 -1267 16 -1267 0 net=3049
rlabel metal2 786 -1267 786 -1267 0 net=4403
rlabel metal2 849 -1267 849 -1267 0 net=4815
rlabel metal2 961 -1267 961 -1267 0 net=5163
rlabel metal2 1003 -1267 1003 -1267 0 net=5463
rlabel metal2 1066 -1267 1066 -1267 0 net=6459
rlabel metal2 1255 -1267 1255 -1267 0 net=7591
rlabel metal2 61 -1269 61 -1269 0 net=7427
rlabel metal2 170 -1271 170 -1271 0 net=5691
rlabel metal2 1087 -1271 1087 -1271 0 net=5689
rlabel metal2 1255 -1271 1255 -1271 0 net=6995
rlabel metal2 233 -1273 233 -1273 0 net=1163
rlabel metal2 625 -1273 625 -1273 0 net=4733
rlabel metal2 866 -1273 866 -1273 0 net=7001
rlabel metal2 1276 -1273 1276 -1273 0 net=7109
rlabel metal2 240 -1275 240 -1275 0 net=2273
rlabel metal2 485 -1275 485 -1275 0 net=2409
rlabel metal2 583 -1275 583 -1275 0 net=2305
rlabel metal2 639 -1275 639 -1275 0 net=3187
rlabel metal2 800 -1275 800 -1275 0 net=4869
rlabel metal2 933 -1275 933 -1275 0 net=5039
rlabel metal2 975 -1275 975 -1275 0 net=5675
rlabel metal2 1087 -1275 1087 -1275 0 net=5897
rlabel metal2 1122 -1275 1122 -1275 0 net=5789
rlabel metal2 1290 -1275 1290 -1275 0 net=7337
rlabel metal2 68 -1277 68 -1277 0 net=5983
rlabel metal2 1311 -1277 1311 -1277 0 net=7283
rlabel metal2 114 -1279 114 -1279 0 net=5903
rlabel metal2 65 -1281 65 -1281 0 net=2495
rlabel metal2 240 -1281 240 -1281 0 net=1215
rlabel metal2 744 -1281 744 -1281 0 net=4977
rlabel metal2 1024 -1281 1024 -1281 0 net=5571
rlabel metal2 247 -1283 247 -1283 0 net=1239
rlabel metal2 324 -1283 324 -1283 0 net=2705
rlabel metal2 499 -1283 499 -1283 0 net=3437
rlabel metal2 730 -1283 730 -1283 0 net=7089
rlabel metal2 79 -1285 79 -1285 0 net=2129
rlabel metal2 583 -1285 583 -1285 0 net=2859
rlabel metal2 821 -1285 821 -1285 0 net=4491
rlabel metal2 870 -1285 870 -1285 0 net=5087
rlabel metal2 79 -1287 79 -1287 0 net=1809
rlabel metal2 331 -1287 331 -1287 0 net=1529
rlabel metal2 443 -1287 443 -1287 0 net=2891
rlabel metal2 730 -1287 730 -1287 0 net=5654
rlabel metal2 107 -1289 107 -1289 0 net=2158
rlabel metal2 513 -1289 513 -1289 0 net=4437
rlabel metal2 1059 -1289 1059 -1289 0 net=6691
rlabel metal2 86 -1291 86 -1291 0 net=1689
rlabel metal2 184 -1291 184 -1291 0 net=1431
rlabel metal2 338 -1291 338 -1291 0 net=2221
rlabel metal2 513 -1291 513 -1291 0 net=3315
rlabel metal2 744 -1291 744 -1291 0 net=3939
rlabel metal2 828 -1291 828 -1291 0 net=4987
rlabel metal2 1213 -1291 1213 -1291 0 net=6633
rlabel metal2 86 -1293 86 -1293 0 net=5947
rlabel metal2 1213 -1293 1213 -1293 0 net=6755
rlabel metal2 184 -1295 184 -1295 0 net=1147
rlabel metal2 747 -1295 747 -1295 0 net=5197
rlabel metal2 247 -1297 247 -1297 0 net=4291
rlabel metal2 688 -1297 688 -1297 0 net=3549
rlabel metal2 856 -1297 856 -1297 0 net=4605
rlabel metal2 877 -1297 877 -1297 0 net=4717
rlabel metal2 877 -1297 877 -1297 0 net=4717
rlabel metal2 891 -1297 891 -1297 0 net=4915
rlabel metal2 338 -1299 338 -1299 0 net=1879
rlabel metal2 523 -1299 523 -1299 0 net=6971
rlabel metal2 9 -1301 9 -1301 0 net=2667
rlabel metal2 702 -1301 702 -1301 0 net=4969
rlabel metal2 9 -1303 9 -1303 0 net=4057
rlabel metal2 863 -1303 863 -1303 0 net=7251
rlabel metal2 345 -1305 345 -1305 0 net=2425
rlabel metal2 772 -1305 772 -1305 0 net=4283
rlabel metal2 898 -1305 898 -1305 0 net=5133
rlabel metal2 268 -1307 268 -1307 0 net=2464
rlabel metal2 814 -1307 814 -1307 0 net=5340
rlabel metal2 268 -1309 268 -1309 0 net=2035
rlabel metal2 369 -1309 369 -1309 0 net=6413
rlabel metal2 359 -1311 359 -1311 0 net=2465
rlabel metal2 905 -1311 905 -1311 0 net=4959
rlabel metal2 376 -1313 376 -1313 0 net=3397
rlabel metal2 912 -1313 912 -1313 0 net=4937
rlabel metal2 380 -1315 380 -1315 0 net=1449
rlabel metal2 761 -1315 761 -1315 0 net=411
rlabel metal2 23 -1317 23 -1317 0 net=1753
rlabel metal2 404 -1317 404 -1317 0 net=6061
rlabel metal2 23 -1319 23 -1319 0 net=1413
rlabel metal2 128 -1321 128 -1321 0 net=1311
rlabel metal2 275 -1323 275 -1323 0 net=3905
rlabel metal2 9 -1334 9 -1334 0 net=4059
rlabel metal2 9 -1334 9 -1334 0 net=4059
rlabel metal2 33 -1334 33 -1334 0 net=1690
rlabel metal2 121 -1334 121 -1334 0 net=7428
rlabel metal2 1423 -1334 1423 -1334 0 net=7373
rlabel metal2 1458 -1334 1458 -1334 0 net=6213
rlabel metal2 44 -1336 44 -1336 0 net=1502
rlabel metal2 387 -1336 387 -1336 0 net=5692
rlabel metal2 1122 -1336 1122 -1336 0 net=5985
rlabel metal2 44 -1338 44 -1338 0 net=4097
rlabel metal2 814 -1338 814 -1338 0 net=6634
rlabel metal2 1255 -1338 1255 -1338 0 net=6997
rlabel metal2 1360 -1338 1360 -1338 0 net=7601
rlabel metal2 65 -1340 65 -1340 0 net=2634
rlabel metal2 583 -1340 583 -1340 0 net=2861
rlabel metal2 635 -1340 635 -1340 0 net=4718
rlabel metal2 887 -1340 887 -1340 0 net=4608
rlabel metal2 65 -1342 65 -1342 0 net=3503
rlabel metal2 135 -1342 135 -1342 0 net=7385
rlabel metal2 61 -1344 61 -1344 0 net=1397
rlabel metal2 163 -1344 163 -1344 0 net=769
rlabel metal2 793 -1344 793 -1344 0 net=4451
rlabel metal2 898 -1344 898 -1344 0 net=5330
rlabel metal2 1129 -1344 1129 -1344 0 net=6041
rlabel metal2 68 -1346 68 -1346 0 net=109
rlabel metal2 464 -1346 464 -1346 0 net=2088
rlabel metal2 614 -1346 614 -1346 0 net=5758
rlabel metal2 1136 -1346 1136 -1346 0 net=6063
rlabel metal2 1136 -1346 1136 -1346 0 net=6063
rlabel metal2 1150 -1346 1150 -1346 0 net=6197
rlabel metal2 1262 -1346 1262 -1346 0 net=7003
rlabel metal2 30 -1348 30 -1348 0 net=2607
rlabel metal2 646 -1348 646 -1348 0 net=2958
rlabel metal2 821 -1348 821 -1348 0 net=4493
rlabel metal2 912 -1348 912 -1348 0 net=7494
rlabel metal2 79 -1350 79 -1350 0 net=1432
rlabel metal2 380 -1350 380 -1350 0 net=1754
rlabel metal2 478 -1350 478 -1350 0 net=2223
rlabel metal2 478 -1350 478 -1350 0 net=2223
rlabel metal2 509 -1350 509 -1350 0 net=7194
rlabel metal2 1332 -1350 1332 -1350 0 net=7439
rlabel metal2 82 -1352 82 -1352 0 net=5690
rlabel metal2 1234 -1352 1234 -1352 0 net=6821
rlabel metal2 1339 -1352 1339 -1352 0 net=7531
rlabel metal2 82 -1354 82 -1354 0 net=707
rlabel metal2 821 -1354 821 -1354 0 net=7272
rlabel metal2 1269 -1354 1269 -1354 0 net=7063
rlabel metal2 86 -1356 86 -1356 0 net=1002
rlabel metal2 107 -1356 107 -1356 0 net=3707
rlabel metal2 380 -1356 380 -1356 0 net=3321
rlabel metal2 695 -1356 695 -1356 0 net=3398
rlabel metal2 852 -1356 852 -1356 0 net=7090
rlabel metal2 1094 -1356 1094 -1356 0 net=6277
rlabel metal2 1297 -1356 1297 -1356 0 net=7361
rlabel metal2 86 -1358 86 -1358 0 net=1137
rlabel metal2 254 -1358 254 -1358 0 net=1811
rlabel metal2 376 -1358 376 -1358 0 net=5179
rlabel metal2 1059 -1358 1059 -1358 0 net=6693
rlabel metal2 1318 -1358 1318 -1358 0 net=6957
rlabel metal2 1346 -1358 1346 -1358 0 net=7593
rlabel metal2 100 -1360 100 -1360 0 net=1853
rlabel metal2 317 -1360 317 -1360 0 net=1241
rlabel metal2 415 -1360 415 -1360 0 net=7252
rlabel metal2 23 -1362 23 -1362 0 net=1415
rlabel metal2 324 -1362 324 -1362 0 net=1531
rlabel metal2 418 -1362 418 -1362 0 net=4606
rlabel metal2 866 -1362 866 -1362 0 net=4626
rlabel metal2 982 -1362 982 -1362 0 net=5239
rlabel metal2 1157 -1362 1157 -1362 0 net=6223
rlabel metal2 1241 -1362 1241 -1362 0 net=6973
rlabel metal2 23 -1364 23 -1364 0 net=4293
rlabel metal2 429 -1364 429 -1364 0 net=937
rlabel metal2 968 -1364 968 -1364 0 net=5199
rlabel metal2 996 -1364 996 -1364 0 net=5259
rlabel metal2 1164 -1364 1164 -1364 0 net=6305
rlabel metal2 37 -1366 37 -1366 0 net=1308
rlabel metal2 429 -1366 429 -1366 0 net=1975
rlabel metal2 583 -1366 583 -1366 0 net=1801
rlabel metal2 649 -1366 649 -1366 0 net=5556
rlabel metal2 1045 -1366 1045 -1366 0 net=5833
rlabel metal2 1164 -1366 1164 -1366 0 net=5711
rlabel metal2 1178 -1366 1178 -1366 0 net=6335
rlabel metal2 37 -1368 37 -1368 0 net=2501
rlabel metal2 541 -1368 541 -1368 0 net=4438
rlabel metal2 954 -1368 954 -1368 0 net=5135
rlabel metal2 1045 -1368 1045 -1368 0 net=3103
rlabel metal2 93 -1370 93 -1370 0 net=3625
rlabel metal2 436 -1370 436 -1370 0 net=3603
rlabel metal2 698 -1370 698 -1370 0 net=4833
rlabel metal2 1017 -1370 1017 -1370 0 net=5767
rlabel metal2 1192 -1370 1192 -1370 0 net=6415
rlabel metal2 1276 -1370 1276 -1370 0 net=7111
rlabel metal2 93 -1372 93 -1372 0 net=1213
rlabel metal2 534 -1372 534 -1372 0 net=2935
rlabel metal2 632 -1372 632 -1372 0 net=6543
rlabel metal2 121 -1374 121 -1374 0 net=3799
rlabel metal2 152 -1374 152 -1374 0 net=2531
rlabel metal2 436 -1374 436 -1374 0 net=1947
rlabel metal2 541 -1374 541 -1374 0 net=4405
rlabel metal2 793 -1374 793 -1374 0 net=7069
rlabel metal2 1024 -1374 1024 -1374 0 net=5573
rlabel metal2 1101 -1374 1101 -1374 0 net=5905
rlabel metal2 1192 -1374 1192 -1374 0 net=7303
rlabel metal2 128 -1376 128 -1376 0 net=1313
rlabel metal2 443 -1376 443 -1376 0 net=4515
rlabel metal2 1199 -1376 1199 -1376 0 net=6447
rlabel metal2 128 -1378 128 -1378 0 net=4530
rlabel metal2 457 -1378 457 -1378 0 net=6785
rlabel metal2 131 -1380 131 -1380 0 net=6375
rlabel metal2 149 -1382 149 -1382 0 net=2892
rlabel metal2 632 -1382 632 -1382 0 net=2093
rlabel metal2 870 -1382 870 -1382 0 net=5089
rlabel metal2 1031 -1382 1031 -1382 0 net=5677
rlabel metal2 1199 -1382 1199 -1382 0 net=7339
rlabel metal2 163 -1384 163 -1384 0 net=1087
rlabel metal2 527 -1384 527 -1384 0 net=4339
rlabel metal2 884 -1384 884 -1384 0 net=4827
rlabel metal2 1010 -1384 1010 -1384 0 net=5525
rlabel metal2 1206 -1384 1206 -1384 0 net=6461
rlabel metal2 170 -1386 170 -1386 0 net=4725
rlabel metal2 933 -1386 933 -1386 0 net=4979
rlabel metal2 1143 -1386 1143 -1386 0 net=6107
rlabel metal2 170 -1388 170 -1388 0 net=1987
rlabel metal2 702 -1388 702 -1388 0 net=5164
rlabel metal2 198 -1390 198 -1390 0 net=1766
rlabel metal2 513 -1390 513 -1390 0 net=3317
rlabel metal2 705 -1390 705 -1390 0 net=5040
rlabel metal2 184 -1392 184 -1392 0 net=1149
rlabel metal2 205 -1392 205 -1392 0 net=1473
rlabel metal2 205 -1392 205 -1392 0 net=1473
rlabel metal2 212 -1392 212 -1392 0 net=2008
rlabel metal2 394 -1392 394 -1392 0 net=2553
rlabel metal2 544 -1392 544 -1392 0 net=3396
rlabel metal2 667 -1392 667 -1392 0 net=3763
rlabel metal2 758 -1392 758 -1392 0 net=4181
rlabel metal2 814 -1392 814 -1392 0 net=6473
rlabel metal2 184 -1394 184 -1394 0 net=1217
rlabel metal2 247 -1394 247 -1394 0 net=1787
rlabel metal2 590 -1394 590 -1394 0 net=3473
rlabel metal2 667 -1394 667 -1394 0 net=4871
rlabel metal2 828 -1394 828 -1394 0 net=4989
rlabel metal2 191 -1396 191 -1396 0 net=1349
rlabel metal2 219 -1396 219 -1396 0 net=1627
rlabel metal2 401 -1396 401 -1396 0 net=2669
rlabel metal2 551 -1396 551 -1396 0 net=5495
rlabel metal2 2 -1398 2 -1398 0 net=1391
rlabel metal2 240 -1398 240 -1398 0 net=2707
rlabel metal2 492 -1398 492 -1398 0 net=3065
rlabel metal2 716 -1398 716 -1398 0 net=4220
rlabel metal2 831 -1398 831 -1398 0 net=6051
rlabel metal2 2 -1400 2 -1400 0 net=2267
rlabel metal2 275 -1400 275 -1400 0 net=3907
rlabel metal2 842 -1400 842 -1400 0 net=4781
rlabel metal2 940 -1400 940 -1400 0 net=5077
rlabel metal2 51 -1402 51 -1402 0 net=1299
rlabel metal2 275 -1402 275 -1402 0 net=1639
rlabel metal2 625 -1402 625 -1402 0 net=2307
rlabel metal2 716 -1402 716 -1402 0 net=3941
rlabel metal2 758 -1402 758 -1402 0 net=4285
rlabel metal2 779 -1402 779 -1402 0 net=5845
rlabel metal2 79 -1404 79 -1404 0 net=2959
rlabel metal2 303 -1404 303 -1404 0 net=1050
rlabel metal2 450 -1404 450 -1404 0 net=2275
rlabel metal2 492 -1404 492 -1404 0 net=2323
rlabel metal2 548 -1404 548 -1404 0 net=7284
rlabel metal2 89 -1406 89 -1406 0 net=3937
rlabel metal2 1213 -1406 1213 -1406 0 net=6757
rlabel metal2 138 -1408 138 -1408 0 net=4311
rlabel metal2 866 -1408 866 -1408 0 net=5109
rlabel metal2 1185 -1408 1185 -1408 0 net=5791
rlabel metal2 282 -1410 282 -1410 0 net=1441
rlabel metal2 464 -1410 464 -1410 0 net=1339
rlabel metal2 891 -1410 891 -1410 0 net=4917
rlabel metal2 1115 -1410 1115 -1410 0 net=5977
rlabel metal2 282 -1412 282 -1412 0 net=1705
rlabel metal2 303 -1412 303 -1412 0 net=1597
rlabel metal2 520 -1412 520 -1412 0 net=7247
rlabel metal2 289 -1414 289 -1414 0 net=4231
rlabel metal2 796 -1414 796 -1414 0 net=5513
rlabel metal2 310 -1416 310 -1416 0 net=2143
rlabel metal2 730 -1416 730 -1416 0 net=5229
rlabel metal2 352 -1418 352 -1418 0 net=2467
rlabel metal2 562 -1418 562 -1418 0 net=3713
rlabel metal2 905 -1418 905 -1418 0 net=4961
rlabel metal2 338 -1420 338 -1420 0 net=1880
rlabel metal2 597 -1420 597 -1420 0 net=2899
rlabel metal2 639 -1420 639 -1420 0 net=3189
rlabel metal2 688 -1420 688 -1420 0 net=3551
rlabel metal2 737 -1420 737 -1420 0 net=3841
rlabel metal2 905 -1420 905 -1420 0 net=5949
rlabel metal2 166 -1422 166 -1422 0 net=2793
rlabel metal2 604 -1422 604 -1422 0 net=3297
rlabel metal2 709 -1422 709 -1422 0 net=3667
rlabel metal2 926 -1422 926 -1422 0 net=4971
rlabel metal2 1087 -1422 1087 -1422 0 net=5899
rlabel metal2 268 -1424 268 -1424 0 net=2037
rlabel metal2 359 -1424 359 -1424 0 net=2131
rlabel metal2 576 -1424 576 -1424 0 net=2801
rlabel metal2 642 -1424 642 -1424 0 net=4585
rlabel metal2 915 -1424 915 -1424 0 net=4749
rlabel metal2 1003 -1424 1003 -1424 0 net=5465
rlabel metal2 58 -1426 58 -1426 0 net=5011
rlabel metal2 58 -1428 58 -1428 0 net=1543
rlabel metal2 114 -1428 114 -1428 0 net=2497
rlabel metal2 387 -1428 387 -1428 0 net=1803
rlabel metal2 674 -1428 674 -1428 0 net=3439
rlabel metal2 719 -1428 719 -1428 0 net=7552
rlabel metal2 72 -1430 72 -1430 0 net=2291
rlabel metal2 499 -1430 499 -1430 0 net=2411
rlabel metal2 611 -1430 611 -1430 0 net=3261
rlabel metal2 723 -1430 723 -1430 0 net=6517
rlabel metal2 16 -1432 16 -1432 0 net=3051
rlabel metal2 919 -1432 919 -1432 0 net=4939
rlabel metal2 16 -1434 16 -1434 0 net=1451
rlabel metal2 506 -1434 506 -1434 0 net=6229
rlabel metal2 114 -1436 114 -1436 0 net=2427
rlabel metal2 408 -1436 408 -1436 0 net=4336
rlabel metal2 835 -1436 835 -1436 0 net=4735
rlabel metal2 173 -1438 173 -1438 0 net=2709
rlabel metal2 807 -1438 807 -1438 0 net=4817
rlabel metal2 226 -1440 226 -1440 0 net=1165
rlabel metal2 345 -1440 345 -1440 0 net=1971
rlabel metal2 828 -1440 828 -1440 0 net=4115
rlabel metal2 156 -1442 156 -1442 0 net=2995
rlabel metal2 401 -1442 401 -1442 0 net=1825
rlabel metal2 156 -1444 156 -1444 0 net=1267
rlabel metal2 422 -1444 422 -1444 0 net=2061
rlabel metal2 142 -1446 142 -1446 0 net=1077
rlabel metal2 390 -1446 390 -1446 0 net=2257
rlabel metal2 142 -1448 142 -1448 0 net=3857
rlabel metal2 9 -1459 9 -1459 0 net=4060
rlabel metal2 44 -1459 44 -1459 0 net=4098
rlabel metal2 460 -1459 460 -1459 0 net=3938
rlabel metal2 1454 -1459 1454 -1459 0 net=6214
rlabel metal2 12 -1461 12 -1461 0 net=2498
rlabel metal2 282 -1461 282 -1461 0 net=1706
rlabel metal2 523 -1461 523 -1461 0 net=3440
rlabel metal2 723 -1461 723 -1461 0 net=4116
rlabel metal2 852 -1461 852 -1461 0 net=6462
rlabel metal2 19 -1463 19 -1463 0 net=5986
rlabel metal2 44 -1465 44 -1465 0 net=2277
rlabel metal2 520 -1465 520 -1465 0 net=3298
rlabel metal2 702 -1465 702 -1465 0 net=2308
rlabel metal2 793 -1465 793 -1465 0 net=6376
rlabel metal2 51 -1467 51 -1467 0 net=1300
rlabel metal2 527 -1467 527 -1467 0 net=2555
rlabel metal2 527 -1467 527 -1467 0 net=2555
rlabel metal2 534 -1467 534 -1467 0 net=3474
rlabel metal2 621 -1467 621 -1467 0 net=6694
rlabel metal2 51 -1469 51 -1469 0 net=3552
rlabel metal2 744 -1469 744 -1469 0 net=6198
rlabel metal2 1269 -1469 1269 -1469 0 net=7065
rlabel metal2 65 -1471 65 -1471 0 net=3504
rlabel metal2 558 -1471 558 -1471 0 net=4990
rlabel metal2 1297 -1471 1297 -1471 0 net=7249
rlabel metal2 65 -1473 65 -1473 0 net=4341
rlabel metal2 884 -1473 884 -1473 0 net=5137
rlabel metal2 93 -1475 93 -1475 0 net=1214
rlabel metal2 534 -1475 534 -1475 0 net=4872
rlabel metal2 688 -1475 688 -1475 0 net=3605
rlabel metal2 705 -1475 705 -1475 0 net=5180
rlabel metal2 37 -1477 37 -1477 0 net=2503
rlabel metal2 100 -1477 100 -1477 0 net=1854
rlabel metal2 562 -1477 562 -1477 0 net=6306
rlabel metal2 37 -1479 37 -1479 0 net=4494
rlabel metal2 940 -1479 940 -1479 0 net=4981
rlabel metal2 1010 -1479 1010 -1479 0 net=5261
rlabel metal2 1234 -1479 1234 -1479 0 net=6787
rlabel metal2 103 -1481 103 -1481 0 net=1442
rlabel metal2 548 -1481 548 -1481 0 net=2803
rlabel metal2 639 -1481 639 -1481 0 net=4940
rlabel metal2 107 -1483 107 -1483 0 net=3708
rlabel metal2 121 -1483 121 -1483 0 net=3800
rlabel metal2 180 -1483 180 -1483 0 net=5311
rlabel metal2 779 -1483 779 -1483 0 net=6822
rlabel metal2 100 -1485 100 -1485 0 net=3409
rlabel metal2 121 -1485 121 -1485 0 net=2533
rlabel metal2 443 -1485 443 -1485 0 net=3714
rlabel metal2 793 -1485 793 -1485 0 net=4313
rlabel metal2 859 -1485 859 -1485 0 net=6758
rlabel metal2 1332 -1485 1332 -1485 0 net=7387
rlabel metal2 128 -1487 128 -1487 0 net=5906
rlabel metal2 1318 -1487 1318 -1487 0 net=7363
rlabel metal2 128 -1489 128 -1489 0 net=2063
rlabel metal2 446 -1489 446 -1489 0 net=6781
rlabel metal2 1325 -1489 1325 -1489 0 net=7375
rlabel metal2 131 -1491 131 -1491 0 net=363
rlabel metal2 450 -1491 450 -1491 0 net=3067
rlabel metal2 663 -1491 663 -1491 0 net=77
rlabel metal2 138 -1493 138 -1493 0 net=3908
rlabel metal2 814 -1493 814 -1493 0 net=4516
rlabel metal2 1171 -1493 1171 -1493 0 net=6417
rlabel metal2 149 -1495 149 -1495 0 net=738
rlabel metal2 863 -1495 863 -1495 0 net=6042
rlabel metal2 149 -1497 149 -1497 0 net=1989
rlabel metal2 226 -1497 226 -1497 0 net=1167
rlabel metal2 226 -1497 226 -1497 0 net=1167
rlabel metal2 240 -1497 240 -1497 0 net=2708
rlabel metal2 562 -1497 562 -1497 0 net=2863
rlabel metal2 639 -1497 639 -1497 0 net=3191
rlabel metal2 667 -1497 667 -1497 0 net=3669
rlabel metal2 758 -1497 758 -1497 0 net=4287
rlabel metal2 796 -1497 796 -1497 0 net=3104
rlabel metal2 1052 -1497 1052 -1497 0 net=5527
rlabel metal2 1157 -1497 1157 -1497 0 net=5793
rlabel metal2 72 -1499 72 -1499 0 net=2293
rlabel metal2 191 -1499 191 -1499 0 net=1393
rlabel metal2 261 -1499 261 -1499 0 net=2961
rlabel metal2 653 -1499 653 -1499 0 net=3319
rlabel metal2 702 -1499 702 -1499 0 net=6555
rlabel metal2 58 -1501 58 -1501 0 net=1545
rlabel metal2 86 -1501 86 -1501 0 net=1139
rlabel metal2 254 -1501 254 -1501 0 net=1315
rlabel metal2 268 -1501 268 -1501 0 net=1331
rlabel metal2 415 -1501 415 -1501 0 net=3053
rlabel metal2 709 -1501 709 -1501 0 net=3727
rlabel metal2 765 -1501 765 -1501 0 net=4183
rlabel metal2 800 -1501 800 -1501 0 net=6974
rlabel metal2 23 -1503 23 -1503 0 net=4295
rlabel metal2 814 -1503 814 -1503 0 net=4453
rlabel metal2 898 -1503 898 -1503 0 net=5575
rlabel metal2 1192 -1503 1192 -1503 0 net=7305
rlabel metal2 1346 -1503 1346 -1503 0 net=7595
rlabel metal2 23 -1505 23 -1505 0 net=2585
rlabel metal2 58 -1505 58 -1505 0 net=2145
rlabel metal2 331 -1505 331 -1505 0 net=3627
rlabel metal2 716 -1505 716 -1505 0 net=3943
rlabel metal2 817 -1505 817 -1505 0 net=5466
rlabel metal2 1094 -1505 1094 -1505 0 net=6545
rlabel metal2 16 -1507 16 -1507 0 net=1453
rlabel metal2 338 -1507 338 -1507 0 net=2039
rlabel metal2 478 -1507 478 -1507 0 net=2224
rlabel metal2 716 -1507 716 -1507 0 net=3765
rlabel metal2 821 -1507 821 -1507 0 net=4471
rlabel metal2 982 -1507 982 -1507 0 net=7071
rlabel metal2 16 -1509 16 -1509 0 net=3515
rlabel metal2 723 -1509 723 -1509 0 net=3843
rlabel metal2 824 -1509 824 -1509 0 net=7532
rlabel metal2 219 -1511 219 -1511 0 net=1629
rlabel metal2 338 -1511 338 -1511 0 net=2413
rlabel metal2 565 -1511 565 -1511 0 net=3949
rlabel metal2 828 -1511 828 -1511 0 net=5978
rlabel metal2 1192 -1511 1192 -1511 0 net=6475
rlabel metal2 2 -1513 2 -1513 0 net=2268
rlabel metal2 247 -1513 247 -1513 0 net=1789
rlabel metal2 282 -1513 282 -1513 0 net=1973
rlabel metal2 380 -1513 380 -1513 0 net=3323
rlabel metal2 478 -1513 478 -1513 0 net=2325
rlabel metal2 572 -1513 572 -1513 0 net=212
rlabel metal2 870 -1513 870 -1513 0 net=5079
rlabel metal2 1038 -1513 1038 -1513 0 net=5497
rlabel metal2 1185 -1513 1185 -1513 0 net=6449
rlabel metal2 2 -1515 2 -1515 0 net=1641
rlabel metal2 289 -1515 289 -1515 0 net=4233
rlabel metal2 831 -1515 831 -1515 0 net=5678
rlabel metal2 1199 -1515 1199 -1515 0 net=7341
rlabel metal2 9 -1517 9 -1517 0 net=2075
rlabel metal2 289 -1517 289 -1517 0 net=1719
rlabel metal2 485 -1517 485 -1517 0 net=4125
rlabel metal2 831 -1517 831 -1517 0 net=7004
rlabel metal2 114 -1519 114 -1519 0 net=2429
rlabel metal2 583 -1519 583 -1519 0 net=1802
rlabel metal2 835 -1519 835 -1519 0 net=4587
rlabel metal2 905 -1519 905 -1519 0 net=5951
rlabel metal2 1129 -1519 1129 -1519 0 net=5769
rlabel metal2 1283 -1519 1283 -1519 0 net=7113
rlabel metal2 40 -1521 40 -1521 0 net=2869
rlabel metal2 590 -1521 590 -1521 0 net=3263
rlabel metal2 842 -1521 842 -1521 0 net=4727
rlabel metal2 954 -1521 954 -1521 0 net=4835
rlabel metal2 996 -1521 996 -1521 0 net=5847
rlabel metal2 89 -1523 89 -1523 0 net=4909
rlabel metal2 1059 -1523 1059 -1523 0 net=5231
rlabel metal2 1129 -1523 1129 -1523 0 net=6053
rlabel metal2 30 -1525 30 -1525 0 net=5119
rlabel metal2 30 -1527 30 -1527 0 net=2133
rlabel metal2 380 -1527 380 -1527 0 net=2795
rlabel metal2 611 -1527 611 -1527 0 net=3041
rlabel metal2 649 -1527 649 -1527 0 net=3427
rlabel metal2 807 -1527 807 -1527 0 net=4819
rlabel metal2 1073 -1527 1073 -1527 0 net=6519
rlabel metal2 114 -1529 114 -1529 0 net=3917
rlabel metal2 849 -1529 849 -1529 0 net=4737
rlabel metal2 1080 -1529 1080 -1529 0 net=6225
rlabel metal2 1304 -1529 1304 -1529 0 net=6959
rlabel metal2 142 -1531 142 -1531 0 net=3859
rlabel metal2 1115 -1531 1115 -1531 0 net=5515
rlabel metal2 1339 -1531 1339 -1531 0 net=7441
rlabel metal2 142 -1533 142 -1533 0 net=2996
rlabel metal2 317 -1533 317 -1533 0 net=4865
rlabel metal2 1108 -1533 1108 -1533 0 net=5901
rlabel metal2 1150 -1533 1150 -1533 0 net=6231
rlabel metal2 198 -1535 198 -1535 0 net=1151
rlabel metal2 324 -1535 324 -1535 0 net=1533
rlabel metal2 919 -1535 919 -1535 0 net=4919
rlabel metal2 82 -1537 82 -1537 0 net=4879
rlabel metal2 345 -1537 345 -1537 0 net=1813
rlabel metal2 397 -1537 397 -1537 0 net=6064
rlabel metal2 198 -1539 198 -1539 0 net=1351
rlabel metal2 233 -1539 233 -1539 0 net=1599
rlabel metal2 352 -1539 352 -1539 0 net=2469
rlabel metal2 366 -1539 366 -1539 0 net=2711
rlabel metal2 625 -1539 625 -1539 0 net=2901
rlabel metal2 859 -1539 859 -1539 0 net=5447
rlabel metal2 177 -1541 177 -1541 0 net=1079
rlabel metal2 296 -1541 296 -1541 0 net=1417
rlabel metal2 352 -1541 352 -1541 0 net=1243
rlabel metal2 404 -1541 404 -1541 0 net=2094
rlabel metal2 863 -1541 863 -1541 0 net=4783
rlabel metal2 961 -1541 961 -1541 0 net=5091
rlabel metal2 135 -1543 135 -1543 0 net=1399
rlabel metal2 373 -1543 373 -1543 0 net=1805
rlabel metal2 408 -1543 408 -1543 0 net=3071
rlabel metal2 513 -1543 513 -1543 0 net=2671
rlabel metal2 625 -1543 625 -1543 0 net=4751
rlabel metal2 933 -1543 933 -1543 0 net=4973
rlabel metal2 1024 -1543 1024 -1543 0 net=6109
rlabel metal2 79 -1545 79 -1545 0 net=4845
rlabel metal2 541 -1545 541 -1545 0 net=4407
rlabel metal2 877 -1545 877 -1545 0 net=4829
rlabel metal2 968 -1545 968 -1545 0 net=5201
rlabel metal2 1143 -1545 1143 -1545 0 net=5835
rlabel metal2 79 -1547 79 -1547 0 net=4523
rlabel metal2 135 -1547 135 -1547 0 net=6823
rlabel metal2 205 -1549 205 -1549 0 net=1475
rlabel metal2 387 -1549 387 -1549 0 net=1341
rlabel metal2 541 -1549 541 -1549 0 net=2609
rlabel metal2 891 -1549 891 -1549 0 net=6336
rlabel metal2 205 -1551 205 -1551 0 net=1051
rlabel metal2 555 -1551 555 -1551 0 net=2937
rlabel metal2 926 -1551 926 -1551 0 net=4963
rlabel metal2 1143 -1551 1143 -1551 0 net=5713
rlabel metal2 1262 -1551 1262 -1551 0 net=6999
rlabel metal2 394 -1553 394 -1553 0 net=2351
rlabel metal2 555 -1553 555 -1553 0 net=607
rlabel metal2 1353 -1553 1353 -1553 0 net=7603
rlabel metal2 394 -1555 394 -1555 0 net=1949
rlabel metal2 569 -1555 569 -1555 0 net=7151
rlabel metal2 401 -1557 401 -1557 0 net=1827
rlabel metal2 856 -1557 856 -1557 0 net=6425
rlabel metal2 163 -1559 163 -1559 0 net=1088
rlabel metal2 429 -1559 429 -1559 0 net=1977
rlabel metal2 856 -1559 856 -1559 0 net=5877
rlabel metal2 163 -1561 163 -1561 0 net=5013
rlabel metal2 429 -1563 429 -1563 0 net=5817
rlabel metal2 887 -1565 887 -1565 0 net=6311
rlabel metal2 947 -1567 947 -1567 0 net=6715
rlabel metal2 968 -1569 968 -1569 0 net=5111
rlabel metal2 145 -1571 145 -1571 0 net=5469
rlabel metal2 1003 -1573 1003 -1573 0 net=5241
rlabel metal2 1066 -1575 1066 -1575 0 net=6279
rlabel metal2 506 -1577 506 -1577 0 net=6869
rlabel metal2 471 -1579 471 -1579 0 net=2259
rlabel metal2 184 -1581 184 -1581 0 net=1219
rlabel metal2 156 -1583 156 -1583 0 net=1269
rlabel metal2 156 -1585 156 -1585 0 net=1013
rlabel metal2 2 -1596 2 -1596 0 net=1642
rlabel metal2 569 -1596 569 -1596 0 net=4738
rlabel metal2 856 -1596 856 -1596 0 net=6280
rlabel metal2 1094 -1596 1094 -1596 0 net=6547
rlabel metal2 1255 -1596 1255 -1596 0 net=7307
rlabel metal2 2 -1598 2 -1598 0 net=2049
rlabel metal2 415 -1598 415 -1598 0 net=3055
rlabel metal2 572 -1598 572 -1598 0 net=2672
rlabel metal2 632 -1598 632 -1598 0 net=1978
rlabel metal2 705 -1598 705 -1598 0 net=4820
rlabel metal2 1045 -1598 1045 -1598 0 net=7596
rlabel metal2 9 -1600 9 -1600 0 net=4983
rlabel metal2 954 -1600 954 -1600 0 net=6055
rlabel metal2 1255 -1600 1255 -1600 0 net=7115
rlabel metal2 12 -1602 12 -1602 0 net=5014
rlabel metal2 177 -1602 177 -1602 0 net=1080
rlabel metal2 233 -1602 233 -1602 0 net=1601
rlabel metal2 233 -1602 233 -1602 0 net=1601
rlabel metal2 320 -1602 320 -1602 0 net=1534
rlabel metal2 940 -1602 940 -1602 0 net=7364
rlabel metal2 51 -1604 51 -1604 0 net=2870
rlabel metal2 632 -1604 632 -1604 0 net=3767
rlabel metal2 754 -1604 754 -1604 0 net=5448
rlabel metal2 1304 -1604 1304 -1604 0 net=6961
rlabel metal2 58 -1606 58 -1606 0 net=2147
rlabel metal2 464 -1606 464 -1606 0 net=2353
rlabel metal2 464 -1606 464 -1606 0 net=2353
rlabel metal2 478 -1606 478 -1606 0 net=2327
rlabel metal2 478 -1606 478 -1606 0 net=2327
rlabel metal2 485 -1606 485 -1606 0 net=3192
rlabel metal2 660 -1606 660 -1606 0 net=3606
rlabel metal2 716 -1606 716 -1606 0 net=3919
rlabel metal2 775 -1606 775 -1606 0 net=4784
rlabel metal2 884 -1606 884 -1606 0 net=5139
rlabel metal2 975 -1606 975 -1606 0 net=6427
rlabel metal2 1304 -1606 1304 -1606 0 net=7389
rlabel metal2 58 -1608 58 -1608 0 net=4847
rlabel metal2 534 -1608 534 -1608 0 net=4836
rlabel metal2 1045 -1608 1045 -1608 0 net=5879
rlabel metal2 1129 -1608 1129 -1608 0 net=6419
rlabel metal2 65 -1610 65 -1610 0 net=4342
rlabel metal2 639 -1610 639 -1610 0 net=3429
rlabel metal2 688 -1610 688 -1610 0 net=4185
rlabel metal2 800 -1610 800 -1610 0 net=5770
rlabel metal2 65 -1612 65 -1612 0 net=1081
rlabel metal2 765 -1612 765 -1612 0 net=4289
rlabel metal2 803 -1612 803 -1612 0 net=6387
rlabel metal2 1199 -1612 1199 -1612 0 net=6789
rlabel metal2 79 -1614 79 -1614 0 net=4525
rlabel metal2 849 -1614 849 -1614 0 net=5081
rlabel metal2 884 -1614 884 -1614 0 net=5577
rlabel metal2 975 -1614 975 -1614 0 net=5529
rlabel metal2 1094 -1614 1094 -1614 0 net=6233
rlabel metal2 1234 -1614 1234 -1614 0 net=7377
rlabel metal2 86 -1616 86 -1616 0 net=943
rlabel metal2 495 -1616 495 -1616 0 net=2804
rlabel metal2 625 -1616 625 -1616 0 net=4753
rlabel metal2 779 -1616 779 -1616 0 net=4455
rlabel metal2 856 -1616 856 -1616 0 net=3725
rlabel metal2 86 -1618 86 -1618 0 net=3411
rlabel metal2 110 -1618 110 -1618 0 net=3331
rlabel metal2 621 -1618 621 -1618 0 net=4651
rlabel metal2 660 -1618 660 -1618 0 net=5243
rlabel metal2 1052 -1618 1052 -1618 0 net=5953
rlabel metal2 1220 -1618 1220 -1618 0 net=5516
rlabel metal2 40 -1620 40 -1620 0 net=5595
rlabel metal2 1220 -1620 1220 -1620 0 net=7073
rlabel metal2 89 -1622 89 -1622 0 net=3728
rlabel metal2 814 -1622 814 -1622 0 net=4729
rlabel metal2 859 -1622 859 -1622 0 net=4866
rlabel metal2 1258 -1622 1258 -1622 0 net=1
rlabel metal2 100 -1624 100 -1624 0 net=6450
rlabel metal2 1276 -1624 1276 -1624 0 net=7605
rlabel metal2 23 -1626 23 -1626 0 net=2587
rlabel metal2 107 -1626 107 -1626 0 net=5797
rlabel metal2 709 -1626 709 -1626 0 net=3945
rlabel metal2 842 -1626 842 -1626 0 net=4831
rlabel metal2 891 -1626 891 -1626 0 net=7000
rlabel metal2 117 -1628 117 -1628 0 net=1270
rlabel metal2 194 -1628 194 -1628 0 net=2796
rlabel metal2 499 -1628 499 -1628 0 net=2431
rlabel metal2 537 -1628 537 -1628 0 net=3861
rlabel metal2 737 -1628 737 -1628 0 net=5181
rlabel metal2 863 -1628 863 -1628 0 net=4921
rlabel metal2 947 -1628 947 -1628 0 net=6717
rlabel metal2 1262 -1628 1262 -1628 0 net=7153
rlabel metal2 138 -1630 138 -1630 0 net=1220
rlabel metal2 485 -1630 485 -1630 0 net=2877
rlabel metal2 506 -1630 506 -1630 0 net=2260
rlabel metal2 730 -1630 730 -1630 0 net=5313
rlabel metal2 982 -1630 982 -1630 0 net=5499
rlabel metal2 1290 -1630 1290 -1630 0 net=7343
rlabel metal2 142 -1632 142 -1632 0 net=5232
rlabel metal2 1311 -1632 1311 -1632 0 net=7443
rlabel metal2 47 -1634 47 -1634 0 net=2471
rlabel metal2 145 -1634 145 -1634 0 net=1790
rlabel metal2 338 -1634 338 -1634 0 net=2414
rlabel metal2 471 -1634 471 -1634 0 net=3043
rlabel metal2 730 -1634 730 -1634 0 net=5979
rlabel metal2 870 -1634 870 -1634 0 net=5113
rlabel metal2 996 -1634 996 -1634 0 net=5849
rlabel metal2 1080 -1634 1080 -1634 0 net=6227
rlabel metal2 93 -1636 93 -1636 0 net=2505
rlabel metal2 345 -1636 345 -1636 0 net=1815
rlabel metal2 345 -1636 345 -1636 0 net=1815
rlabel metal2 352 -1636 352 -1636 0 net=1244
rlabel metal2 506 -1636 506 -1636 0 net=5093
rlabel metal2 968 -1636 968 -1636 0 net=5203
rlabel metal2 996 -1636 996 -1636 0 net=6313
rlabel metal2 93 -1638 93 -1638 0 net=5836
rlabel metal2 103 -1640 103 -1640 0 net=5583
rlabel metal2 1164 -1640 1164 -1640 0 net=6557
rlabel metal2 135 -1642 135 -1642 0 net=6855
rlabel metal2 135 -1644 135 -1644 0 net=1353
rlabel metal2 212 -1644 212 -1644 0 net=1153
rlabel metal2 254 -1644 254 -1644 0 net=1221
rlabel metal2 443 -1644 443 -1644 0 net=3325
rlabel metal2 877 -1644 877 -1644 0 net=4975
rlabel metal2 961 -1644 961 -1644 0 net=5471
rlabel metal2 1206 -1644 1206 -1644 0 net=6783
rlabel metal2 121 -1646 121 -1646 0 net=2535
rlabel metal2 460 -1646 460 -1646 0 net=5423
rlabel metal2 1031 -1646 1031 -1646 0 net=5819
rlabel metal2 1157 -1646 1157 -1646 0 net=5795
rlabel metal2 114 -1648 114 -1648 0 net=6183
rlabel metal2 96 -1650 96 -1650 0 net=1707
rlabel metal2 121 -1650 121 -1650 0 net=1395
rlabel metal2 247 -1650 247 -1650 0 net=2077
rlabel metal2 352 -1650 352 -1650 0 net=2211
rlabel metal2 513 -1650 513 -1650 0 net=4127
rlabel metal2 894 -1650 894 -1650 0 net=5120
rlabel metal2 152 -1652 152 -1652 0 net=1974
rlabel metal2 366 -1652 366 -1652 0 net=2712
rlabel metal2 492 -1652 492 -1652 0 net=2557
rlabel metal2 758 -1652 758 -1652 0 net=4235
rlabel metal2 1066 -1652 1066 -1652 0 net=6651
rlabel metal2 159 -1654 159 -1654 0 net=5297
rlabel metal2 1073 -1654 1073 -1654 0 net=6521
rlabel metal2 163 -1656 163 -1656 0 net=3235
rlabel metal2 1024 -1656 1024 -1656 0 net=6111
rlabel metal2 177 -1658 177 -1658 0 net=3951
rlabel metal2 772 -1658 772 -1658 0 net=5902
rlabel metal2 180 -1660 180 -1660 0 net=2470
rlabel metal2 366 -1660 366 -1660 0 net=2865
rlabel metal2 751 -1660 751 -1660 0 net=4089
rlabel metal2 1024 -1660 1024 -1660 0 net=6825
rlabel metal2 44 -1662 44 -1662 0 net=2279
rlabel metal2 373 -1662 373 -1662 0 net=1807
rlabel metal2 523 -1662 523 -1662 0 net=6581
rlabel metal2 1241 -1662 1241 -1662 0 net=7067
rlabel metal2 44 -1664 44 -1664 0 net=869
rlabel metal2 184 -1664 184 -1664 0 net=1053
rlabel metal2 240 -1664 240 -1664 0 net=1401
rlabel metal2 376 -1664 376 -1664 0 net=3860
rlabel metal2 1115 -1664 1115 -1664 0 net=5715
rlabel metal2 54 -1666 54 -1666 0 net=1845
rlabel metal2 198 -1666 198 -1666 0 net=1631
rlabel metal2 380 -1666 380 -1666 0 net=2041
rlabel metal2 450 -1666 450 -1666 0 net=3069
rlabel metal2 1143 -1666 1143 -1666 0 net=6477
rlabel metal2 51 -1668 51 -1668 0 net=6775
rlabel metal2 205 -1670 205 -1670 0 net=2885
rlabel metal2 422 -1670 422 -1670 0 net=1829
rlabel metal2 450 -1670 450 -1670 0 net=3629
rlabel metal2 828 -1670 828 -1670 0 net=7227
rlabel metal2 226 -1672 226 -1672 0 net=1169
rlabel metal2 324 -1672 324 -1672 0 net=4881
rlabel metal2 226 -1674 226 -1674 0 net=1455
rlabel metal2 324 -1674 324 -1674 0 net=1343
rlabel metal2 394 -1674 394 -1674 0 net=1951
rlabel metal2 527 -1674 527 -1674 0 net=2611
rlabel metal2 562 -1674 562 -1674 0 net=2713
rlabel metal2 695 -1674 695 -1674 0 net=3741
rlabel metal2 128 -1676 128 -1676 0 net=2065
rlabel metal2 394 -1676 394 -1676 0 net=2939
rlabel metal2 72 -1678 72 -1678 0 net=1547
rlabel metal2 275 -1678 275 -1678 0 net=1721
rlabel metal2 303 -1678 303 -1678 0 net=1419
rlabel metal2 331 -1678 331 -1678 0 net=1691
rlabel metal2 541 -1678 541 -1678 0 net=4297
rlabel metal2 72 -1680 72 -1680 0 net=1317
rlabel metal2 282 -1680 282 -1680 0 net=3607
rlabel metal2 786 -1680 786 -1680 0 net=4473
rlabel metal2 156 -1682 156 -1682 0 net=1015
rlabel metal2 404 -1682 404 -1682 0 net=751
rlabel metal2 555 -1682 555 -1682 0 net=3341
rlabel metal2 821 -1682 821 -1682 0 net=3823
rlabel metal2 30 -1684 30 -1684 0 net=2134
rlabel metal2 590 -1684 590 -1684 0 net=3265
rlabel metal2 16 -1686 16 -1686 0 net=402
rlabel metal2 170 -1686 170 -1686 0 net=2295
rlabel metal2 408 -1686 408 -1686 0 net=3073
rlabel metal2 170 -1688 170 -1688 0 net=1333
rlabel metal2 408 -1688 408 -1688 0 net=2963
rlabel metal2 149 -1690 149 -1690 0 net=1991
rlabel metal2 604 -1690 604 -1690 0 net=2903
rlabel metal2 149 -1692 149 -1692 0 net=4910
rlabel metal2 219 -1694 219 -1694 0 net=1791
rlabel metal2 520 -1694 520 -1694 0 net=5165
rlabel metal2 191 -1696 191 -1696 0 net=1141
rlabel metal2 646 -1696 646 -1696 0 net=3517
rlabel metal2 191 -1698 191 -1698 0 net=3320
rlabel metal2 681 -1698 681 -1698 0 net=3845
rlabel metal2 653 -1700 653 -1700 0 net=3671
rlabel metal2 723 -1700 723 -1700 0 net=4315
rlabel metal2 667 -1702 667 -1702 0 net=7250
rlabel metal2 793 -1704 793 -1704 0 net=4409
rlabel metal2 1248 -1704 1248 -1704 0 net=6871
rlabel metal2 37 -1706 37 -1706 0 net=7169
rlabel metal2 37 -1708 37 -1708 0 net=1477
rlabel metal2 807 -1708 807 -1708 0 net=4589
rlabel metal2 317 -1710 317 -1710 0 net=6155
rlabel metal2 835 -1712 835 -1712 0 net=4965
rlabel metal2 926 -1714 926 -1714 0 net=5263
rlabel metal2 373 -1716 373 -1716 0 net=6245
rlabel metal2 9 -1727 9 -1727 0 net=4984
rlabel metal2 117 -1727 117 -1727 0 net=3518
rlabel metal2 667 -1727 667 -1727 0 net=5424
rlabel metal2 940 -1727 940 -1727 0 net=5204
rlabel metal2 1069 -1727 1069 -1727 0 net=7068
rlabel metal2 1318 -1727 1318 -1727 0 net=6962
rlabel metal2 16 -1729 16 -1729 0 net=666
rlabel metal2 33 -1729 33 -1729 0 net=229
rlabel metal2 72 -1729 72 -1729 0 net=1318
rlabel metal2 390 -1729 390 -1729 0 net=3726
rlabel metal2 898 -1729 898 -1729 0 net=6228
rlabel metal2 1122 -1729 1122 -1729 0 net=7606
rlabel metal2 16 -1731 16 -1731 0 net=3259
rlabel metal2 152 -1731 152 -1731 0 net=6503
rlabel metal2 1122 -1731 1122 -1731 0 net=6583
rlabel metal2 1227 -1731 1227 -1731 0 net=5796
rlabel metal2 9 -1733 9 -1733 0 net=3249
rlabel metal2 205 -1733 205 -1733 0 net=2886
rlabel metal2 359 -1733 359 -1733 0 net=2281
rlabel metal2 667 -1733 667 -1733 0 net=3863
rlabel metal2 712 -1733 712 -1733 0 net=4290
rlabel metal2 814 -1733 814 -1733 0 net=4731
rlabel metal2 898 -1733 898 -1733 0 net=5531
rlabel metal2 1171 -1733 1171 -1733 0 net=6857
rlabel metal2 1241 -1733 1241 -1733 0 net=7345
rlabel metal2 19 -1735 19 -1735 0 net=4410
rlabel metal2 828 -1735 828 -1735 0 net=4883
rlabel metal2 828 -1735 828 -1735 0 net=4883
rlabel metal2 835 -1735 835 -1735 0 net=4967
rlabel metal2 901 -1735 901 -1735 0 net=7543
rlabel metal2 23 -1737 23 -1737 0 net=3326
rlabel metal2 702 -1737 702 -1737 0 net=4317
rlabel metal2 744 -1737 744 -1737 0 net=5082
rlabel metal2 933 -1737 933 -1737 0 net=5315
rlabel metal2 968 -1737 968 -1737 0 net=5881
rlabel metal2 1213 -1737 1213 -1737 0 net=7117
rlabel metal2 26 -1739 26 -1739 0 net=2588
rlabel metal2 107 -1739 107 -1739 0 net=3070
rlabel metal2 1255 -1739 1255 -1739 0 net=7391
rlabel metal2 26 -1741 26 -1741 0 net=5500
rlabel metal2 1010 -1741 1010 -1741 0 net=6247
rlabel metal2 30 -1743 30 -1743 0 net=1993
rlabel metal2 324 -1743 324 -1743 0 net=1344
rlabel metal2 404 -1743 404 -1743 0 net=2432
rlabel metal2 548 -1743 548 -1743 0 net=4627
rlabel metal2 835 -1743 835 -1743 0 net=5115
rlabel metal2 940 -1743 940 -1743 0 net=6315
rlabel metal2 1017 -1743 1017 -1743 0 net=6113
rlabel metal2 37 -1745 37 -1745 0 net=1478
rlabel metal2 205 -1745 205 -1745 0 net=1421
rlabel metal2 359 -1745 359 -1745 0 net=2067
rlabel metal2 457 -1745 457 -1745 0 net=6872
rlabel metal2 44 -1747 44 -1747 0 net=1402
rlabel metal2 268 -1747 268 -1747 0 net=2149
rlabel metal2 457 -1747 457 -1747 0 net=4083
rlabel metal2 555 -1747 555 -1747 0 net=3768
rlabel metal2 719 -1747 719 -1747 0 net=5578
rlabel metal2 975 -1747 975 -1747 0 net=5821
rlabel metal2 1073 -1747 1073 -1747 0 net=5717
rlabel metal2 44 -1749 44 -1749 0 net=5298
rlabel metal2 1115 -1749 1115 -1749 0 net=6559
rlabel metal2 47 -1751 47 -1751 0 net=5987
rlabel metal2 1031 -1751 1031 -1751 0 net=6235
rlabel metal2 1164 -1751 1164 -1751 0 net=6777
rlabel metal2 54 -1753 54 -1753 0 net=7170
rlabel metal2 72 -1755 72 -1755 0 net=3699
rlabel metal2 100 -1755 100 -1755 0 net=3369
rlabel metal2 478 -1755 478 -1755 0 net=2328
rlabel metal2 478 -1755 478 -1755 0 net=2328
rlabel metal2 485 -1755 485 -1755 0 net=6137
rlabel metal2 1234 -1755 1234 -1755 0 net=7379
rlabel metal2 51 -1757 51 -1757 0 net=1229
rlabel metal2 107 -1757 107 -1757 0 net=1793
rlabel metal2 369 -1757 369 -1757 0 net=4613
rlabel metal2 747 -1757 747 -1757 0 net=3824
rlabel metal2 849 -1757 849 -1757 0 net=5167
rlabel metal2 1059 -1757 1059 -1757 0 net=6389
rlabel metal2 1192 -1757 1192 -1757 0 net=7075
rlabel metal2 1234 -1757 1234 -1757 0 net=7309
rlabel metal2 51 -1759 51 -1759 0 net=4832
rlabel metal2 912 -1759 912 -1759 0 net=5585
rlabel metal2 1108 -1759 1108 -1759 0 net=6549
rlabel metal2 1220 -1759 1220 -1759 0 net=7229
rlabel metal2 58 -1761 58 -1761 0 net=4849
rlabel metal2 989 -1761 989 -1761 0 net=5955
rlabel metal2 1269 -1761 1269 -1761 0 net=7445
rlabel metal2 58 -1763 58 -1763 0 net=1055
rlabel metal2 212 -1763 212 -1763 0 net=1155
rlabel metal2 212 -1763 212 -1763 0 net=1155
rlabel metal2 226 -1763 226 -1763 0 net=1456
rlabel metal2 534 -1763 534 -1763 0 net=4591
rlabel metal2 821 -1763 821 -1763 0 net=5265
rlabel metal2 1052 -1763 1052 -1763 0 net=6185
rlabel metal2 2 -1765 2 -1765 0 net=2051
rlabel metal2 233 -1765 233 -1765 0 net=1603
rlabel metal2 275 -1765 275 -1765 0 net=1723
rlabel metal2 373 -1765 373 -1765 0 net=2283
rlabel metal2 625 -1765 625 -1765 0 net=4653
rlabel metal2 926 -1765 926 -1765 0 net=5597
rlabel metal2 1087 -1765 1087 -1765 0 net=6479
rlabel metal2 2 -1767 2 -1767 0 net=2967
rlabel metal2 79 -1767 79 -1767 0 net=1846
rlabel metal2 604 -1767 604 -1767 0 net=2905
rlabel metal2 1143 -1767 1143 -1767 0 net=6719
rlabel metal2 79 -1769 79 -1769 0 net=3413
rlabel metal2 121 -1769 121 -1769 0 net=1396
rlabel metal2 401 -1769 401 -1769 0 net=7009
rlabel metal2 86 -1771 86 -1771 0 net=1003
rlabel metal2 317 -1771 317 -1771 0 net=1693
rlabel metal2 401 -1771 401 -1771 0 net=1831
rlabel metal2 488 -1771 488 -1771 0 net=579
rlabel metal2 114 -1773 114 -1773 0 net=1709
rlabel metal2 128 -1773 128 -1773 0 net=1549
rlabel metal2 331 -1773 331 -1773 0 net=1817
rlabel metal2 415 -1773 415 -1773 0 net=1953
rlabel metal2 506 -1773 506 -1773 0 net=5094
rlabel metal2 660 -1773 660 -1773 0 net=5245
rlabel metal2 128 -1775 128 -1775 0 net=1017
rlabel metal2 345 -1775 345 -1775 0 net=2043
rlabel metal2 436 -1775 436 -1775 0 net=3045
rlabel metal2 506 -1775 506 -1775 0 net=4299
rlabel metal2 555 -1775 555 -1775 0 net=2815
rlabel metal2 138 -1777 138 -1777 0 net=2296
rlabel metal2 464 -1777 464 -1777 0 net=2355
rlabel metal2 513 -1777 513 -1777 0 net=4129
rlabel metal2 576 -1777 576 -1777 0 net=3333
rlabel metal2 142 -1779 142 -1779 0 net=2472
rlabel metal2 142 -1781 142 -1781 0 net=2375
rlabel metal2 513 -1781 513 -1781 0 net=2612
rlabel metal2 541 -1781 541 -1781 0 net=2715
rlabel metal2 576 -1781 576 -1781 0 net=3267
rlabel metal2 611 -1781 611 -1781 0 net=4186
rlabel metal2 723 -1781 723 -1781 0 net=4571
rlabel metal2 149 -1783 149 -1783 0 net=3074
rlabel metal2 597 -1783 597 -1783 0 net=3431
rlabel metal2 660 -1783 660 -1783 0 net=3847
rlabel metal2 730 -1783 730 -1783 0 net=5981
rlabel metal2 156 -1785 156 -1785 0 net=6495
rlabel metal2 625 -1785 625 -1785 0 net=4922
rlabel metal2 156 -1787 156 -1787 0 net=1335
rlabel metal2 177 -1787 177 -1787 0 net=3953
rlabel metal2 730 -1787 730 -1787 0 net=4090
rlabel metal2 96 -1789 96 -1789 0 net=5331
rlabel metal2 163 -1791 163 -1791 0 net=3237
rlabel metal2 408 -1791 408 -1791 0 net=2965
rlabel metal2 562 -1791 562 -1791 0 net=3343
rlabel metal2 628 -1791 628 -1791 0 net=5101
rlabel metal2 170 -1793 170 -1793 0 net=3609
rlabel metal2 394 -1793 394 -1793 0 net=2941
rlabel metal2 464 -1793 464 -1793 0 net=5911
rlabel metal2 177 -1795 177 -1795 0 net=1171
rlabel metal2 394 -1795 394 -1795 0 net=1855
rlabel metal2 520 -1795 520 -1795 0 net=6784
rlabel metal2 184 -1797 184 -1797 0 net=1143
rlabel metal2 233 -1797 233 -1797 0 net=3631
rlabel metal2 520 -1797 520 -1797 0 net=3149
rlabel metal2 65 -1799 65 -1799 0 net=1083
rlabel metal2 247 -1799 247 -1799 0 net=2079
rlabel metal2 282 -1799 282 -1799 0 net=2879
rlabel metal2 569 -1799 569 -1799 0 net=3057
rlabel metal2 733 -1799 733 -1799 0 net=4635
rlabel metal2 863 -1799 863 -1799 0 net=6057
rlabel metal2 40 -1801 40 -1801 0 net=898
rlabel metal2 191 -1801 191 -1801 0 net=7171
rlabel metal2 114 -1803 114 -1803 0 net=2953
rlabel metal2 198 -1803 198 -1803 0 net=1633
rlabel metal2 338 -1803 338 -1803 0 net=2507
rlabel metal2 569 -1803 569 -1803 0 net=3743
rlabel metal2 737 -1803 737 -1803 0 net=5183
rlabel metal2 135 -1805 135 -1805 0 net=1355
rlabel metal2 247 -1805 247 -1805 0 net=1223
rlabel metal2 261 -1805 261 -1805 0 net=2559
rlabel metal2 583 -1805 583 -1805 0 net=5799
rlabel metal2 135 -1807 135 -1807 0 net=1503
rlabel metal2 254 -1807 254 -1807 0 net=3585
rlabel metal2 443 -1807 443 -1807 0 net=2537
rlabel metal2 583 -1807 583 -1807 0 net=4236
rlabel metal2 761 -1807 761 -1807 0 net=4976
rlabel metal2 296 -1809 296 -1809 0 net=3920
rlabel metal2 751 -1809 751 -1809 0 net=6522
rlabel metal2 310 -1811 310 -1811 0 net=1669
rlabel metal2 765 -1811 765 -1811 0 net=4527
rlabel metal2 877 -1811 877 -1811 0 net=5141
rlabel metal2 1024 -1811 1024 -1811 0 net=6827
rlabel metal2 338 -1813 338 -1813 0 net=2213
rlabel metal2 366 -1813 366 -1813 0 net=2867
rlabel metal2 618 -1813 618 -1813 0 net=3673
rlabel metal2 674 -1813 674 -1813 0 net=4755
rlabel metal2 905 -1813 905 -1813 0 net=5473
rlabel metal2 1024 -1813 1024 -1813 0 net=6157
rlabel metal2 320 -1815 320 -1815 0 net=3929
rlabel metal2 695 -1815 695 -1815 0 net=3947
rlabel metal2 716 -1815 716 -1815 0 net=6737
rlabel metal2 352 -1817 352 -1817 0 net=394
rlabel metal2 961 -1817 961 -1817 0 net=5851
rlabel metal2 1080 -1817 1080 -1817 0 net=6429
rlabel metal2 366 -1819 366 -1819 0 net=1808
rlabel metal2 443 -1819 443 -1819 0 net=3965
rlabel metal2 607 -1819 607 -1819 0 net=6659
rlabel metal2 23 -1821 23 -1821 0 net=4255
rlabel metal2 485 -1821 485 -1821 0 net=2833
rlabel metal2 1038 -1821 1038 -1821 0 net=7267
rlabel metal2 422 -1823 422 -1823 0 net=3769
rlabel metal2 737 -1823 737 -1823 0 net=5781
rlabel metal2 1066 -1823 1066 -1823 0 net=6421
rlabel metal2 632 -1825 632 -1825 0 net=4457
rlabel metal2 1129 -1825 1129 -1825 0 net=6653
rlabel metal2 639 -1827 639 -1827 0 net=927
rlabel metal2 1178 -1827 1178 -1827 0 net=6791
rlabel metal2 653 -1829 653 -1829 0 net=4791
rlabel metal2 1199 -1829 1199 -1829 0 net=7155
rlabel metal2 558 -1831 558 -1831 0 net=7407
rlabel metal2 779 -1833 779 -1833 0 net=4475
rlabel metal2 194 -1835 194 -1835 0 net=4671
rlabel metal2 2 -1846 2 -1846 0 net=2968
rlabel metal2 604 -1846 604 -1846 0 net=2282
rlabel metal2 653 -1846 653 -1846 0 net=3948
rlabel metal2 712 -1846 712 -1846 0 net=5142
rlabel metal2 16 -1848 16 -1848 0 net=3260
rlabel metal2 432 -1848 432 -1848 0 net=5982
rlabel metal2 9 -1850 9 -1850 0 net=3251
rlabel metal2 23 -1850 23 -1850 0 net=1994
rlabel metal2 37 -1850 37 -1850 0 net=6792
rlabel metal2 9 -1852 9 -1852 0 net=3415
rlabel metal2 89 -1852 89 -1852 0 net=1224
rlabel metal2 254 -1852 254 -1852 0 net=3586
rlabel metal2 373 -1852 373 -1852 0 net=2285
rlabel metal2 373 -1852 373 -1852 0 net=2285
rlabel metal2 387 -1852 387 -1852 0 net=2817
rlabel metal2 558 -1852 558 -1852 0 net=4411
rlabel metal2 656 -1852 656 -1852 0 net=4732
rlabel metal2 1178 -1852 1178 -1852 0 net=7447
rlabel metal2 23 -1854 23 -1854 0 net=1231
rlabel metal2 103 -1854 103 -1854 0 net=3334
rlabel metal2 30 -1856 30 -1856 0 net=3151
rlabel metal2 555 -1856 555 -1856 0 net=6186
rlabel metal2 1094 -1856 1094 -1856 0 net=7347
rlabel metal2 37 -1858 37 -1858 0 net=2215
rlabel metal2 366 -1858 366 -1858 0 net=3046
rlabel metal2 464 -1858 464 -1858 0 net=4300
rlabel metal2 513 -1858 513 -1858 0 net=2717
rlabel metal2 607 -1858 607 -1858 0 net=4968
rlabel metal2 877 -1858 877 -1858 0 net=5989
rlabel metal2 1052 -1858 1052 -1858 0 net=6829
rlabel metal2 40 -1860 40 -1860 0 net=1550
rlabel metal2 296 -1860 296 -1860 0 net=983
rlabel metal2 478 -1860 478 -1860 0 net=4458
rlabel metal2 639 -1860 639 -1860 0 net=4528
rlabel metal2 856 -1860 856 -1860 0 net=6391
rlabel metal2 1157 -1860 1157 -1860 0 net=7311
rlabel metal2 44 -1862 44 -1862 0 net=5102
rlabel metal2 1115 -1862 1115 -1862 0 net=6561
rlabel metal2 44 -1864 44 -1864 0 net=1979
rlabel metal2 114 -1864 114 -1864 0 net=3632
rlabel metal2 254 -1864 254 -1864 0 net=1725
rlabel metal2 331 -1864 331 -1864 0 net=1819
rlabel metal2 331 -1864 331 -1864 0 net=1819
rlabel metal2 408 -1864 408 -1864 0 net=2943
rlabel metal2 471 -1864 471 -1864 0 net=2357
rlabel metal2 485 -1864 485 -1864 0 net=2835
rlabel metal2 485 -1864 485 -1864 0 net=2835
rlabel metal2 492 -1864 492 -1864 0 net=2868
rlabel metal2 719 -1864 719 -1864 0 net=2906
rlabel metal2 996 -1864 996 -1864 0 net=6431
rlabel metal2 1115 -1864 1115 -1864 0 net=7157
rlabel metal2 47 -1866 47 -1866 0 net=5332
rlabel metal2 933 -1866 933 -1866 0 net=5317
rlabel metal2 1080 -1866 1080 -1866 0 net=7077
rlabel metal2 79 -1868 79 -1868 0 net=1955
rlabel metal2 429 -1868 429 -1868 0 net=4257
rlabel metal2 646 -1868 646 -1868 0 net=5599
rlabel metal2 933 -1868 933 -1868 0 net=6237
rlabel metal2 1143 -1868 1143 -1868 0 net=6721
rlabel metal2 93 -1870 93 -1870 0 net=3370
rlabel metal2 114 -1870 114 -1870 0 net=3345
rlabel metal2 597 -1870 597 -1870 0 net=3432
rlabel metal2 614 -1870 614 -1870 0 net=4850
rlabel metal2 891 -1870 891 -1870 0 net=6171
rlabel metal2 926 -1870 926 -1870 0 net=7011
rlabel metal2 100 -1872 100 -1872 0 net=2966
rlabel metal2 534 -1872 534 -1872 0 net=4593
rlabel metal2 597 -1872 597 -1872 0 net=3675
rlabel metal2 628 -1872 628 -1872 0 net=6679
rlabel metal2 1038 -1872 1038 -1872 0 net=7269
rlabel metal2 135 -1874 135 -1874 0 net=4654
rlabel metal2 842 -1874 842 -1874 0 net=5883
rlabel metal2 1164 -1874 1164 -1874 0 net=6779
rlabel metal2 135 -1876 135 -1876 0 net=7365
rlabel metal2 149 -1878 149 -1878 0 net=2137
rlabel metal2 264 -1878 264 -1878 0 net=2880
rlabel metal2 289 -1878 289 -1878 0 net=1671
rlabel metal2 324 -1878 324 -1878 0 net=1857
rlabel metal2 408 -1878 408 -1878 0 net=3931
rlabel metal2 677 -1878 677 -1878 0 net=3058
rlabel metal2 695 -1878 695 -1878 0 net=4673
rlabel metal2 919 -1878 919 -1878 0 net=6589
rlabel metal2 1073 -1878 1073 -1878 0 net=5719
rlabel metal2 86 -1880 86 -1880 0 net=1004
rlabel metal2 299 -1880 299 -1880 0 net=231
rlabel metal2 688 -1880 688 -1880 0 net=4637
rlabel metal2 786 -1880 786 -1880 0 net=5533
rlabel metal2 947 -1880 947 -1880 0 net=6505
rlabel metal2 86 -1882 86 -1882 0 net=6138
rlabel metal2 149 -1884 149 -1884 0 net=1357
rlabel metal2 226 -1884 226 -1884 0 net=2052
rlabel metal2 730 -1884 730 -1884 0 net=4885
rlabel metal2 863 -1884 863 -1884 0 net=6059
rlabel metal2 152 -1886 152 -1886 0 net=2150
rlabel metal2 275 -1886 275 -1886 0 net=2081
rlabel metal2 436 -1886 436 -1886 0 net=2509
rlabel metal2 457 -1886 457 -1886 0 net=4085
rlabel metal2 709 -1886 709 -1886 0 net=5823
rlabel metal2 863 -1886 863 -1886 0 net=5853
rlabel metal2 968 -1886 968 -1886 0 net=6551
rlabel metal2 163 -1888 163 -1888 0 net=1505
rlabel metal2 303 -1888 303 -1888 0 net=1635
rlabel metal2 352 -1888 352 -1888 0 net=514
rlabel metal2 1073 -1888 1073 -1888 0 net=7393
rlabel metal2 163 -1890 163 -1890 0 net=3197
rlabel metal2 422 -1890 422 -1890 0 net=3771
rlabel metal2 471 -1890 471 -1890 0 net=2761
rlabel metal2 898 -1890 898 -1890 0 net=6481
rlabel metal2 177 -1892 177 -1892 0 net=1173
rlabel metal2 275 -1892 275 -1892 0 net=1619
rlabel metal2 177 -1894 177 -1894 0 net=1157
rlabel metal2 285 -1894 285 -1894 0 net=7133
rlabel metal2 184 -1896 184 -1896 0 net=1145
rlabel metal2 303 -1896 303 -1896 0 net=4091
rlabel metal2 527 -1896 527 -1896 0 net=3269
rlabel metal2 709 -1896 709 -1896 0 net=4615
rlabel metal2 751 -1896 751 -1896 0 net=5822
rlabel metal2 1066 -1896 1066 -1896 0 net=6423
rlabel metal2 128 -1898 128 -1898 0 net=1019
rlabel metal2 198 -1898 198 -1898 0 net=1423
rlabel metal2 212 -1898 212 -1898 0 net=1085
rlabel metal2 345 -1898 345 -1898 0 net=2045
rlabel metal2 380 -1898 380 -1898 0 net=3239
rlabel metal2 443 -1898 443 -1898 0 net=3967
rlabel metal2 737 -1898 737 -1898 0 net=5783
rlabel metal2 912 -1898 912 -1898 0 net=5587
rlabel metal2 128 -1900 128 -1900 0 net=2377
rlabel metal2 205 -1900 205 -1900 0 net=1605
rlabel metal2 345 -1900 345 -1900 0 net=1833
rlabel metal2 495 -1900 495 -1900 0 net=4628
rlabel metal2 912 -1900 912 -1900 0 net=6249
rlabel metal2 1066 -1900 1066 -1900 0 net=6859
rlabel metal2 51 -1902 51 -1902 0 net=4763
rlabel metal2 506 -1902 506 -1902 0 net=4573
rlabel metal2 737 -1902 737 -1902 0 net=5169
rlabel metal2 975 -1902 975 -1902 0 net=6661
rlabel metal2 1171 -1902 1171 -1902 0 net=7409
rlabel metal2 51 -1904 51 -1904 0 net=699
rlabel metal2 516 -1904 516 -1904 0 net=6573
rlabel metal2 1045 -1904 1045 -1904 0 net=6739
rlabel metal2 58 -1906 58 -1906 0 net=1057
rlabel metal2 219 -1906 219 -1906 0 net=1695
rlabel metal2 359 -1906 359 -1906 0 net=2069
rlabel metal2 534 -1906 534 -1906 0 net=6497
rlabel metal2 744 -1906 744 -1906 0 net=5117
rlabel metal2 849 -1906 849 -1906 0 net=6159
rlabel metal2 1150 -1906 1150 -1906 0 net=7381
rlabel metal2 58 -1908 58 -1908 0 net=2539
rlabel metal2 541 -1908 541 -1908 0 net=3865
rlabel metal2 751 -1908 751 -1908 0 net=6023
rlabel metal2 765 -1908 765 -1908 0 net=5247
rlabel metal2 1024 -1908 1024 -1908 0 net=6655
rlabel metal2 65 -1910 65 -1910 0 net=5481
rlabel metal2 835 -1910 835 -1910 0 net=7118
rlabel metal2 138 -1912 138 -1912 0 net=4739
rlabel metal2 754 -1912 754 -1912 0 net=6316
rlabel metal2 1213 -1912 1213 -1912 0 net=7545
rlabel metal2 138 -1914 138 -1914 0 net=1336
rlabel metal2 191 -1914 191 -1914 0 net=2955
rlabel metal2 548 -1914 548 -1914 0 net=4131
rlabel metal2 667 -1914 667 -1914 0 net=4319
rlabel metal2 758 -1914 758 -1914 0 net=4476
rlabel metal2 156 -1916 156 -1916 0 net=1121
rlabel metal2 548 -1916 548 -1916 0 net=3475
rlabel metal2 702 -1916 702 -1916 0 net=6723
rlabel metal2 191 -1918 191 -1918 0 net=1383
rlabel metal2 380 -1918 380 -1918 0 net=3211
rlabel metal2 761 -1918 761 -1918 0 net=6011
rlabel metal2 72 -1920 72 -1920 0 net=3700
rlabel metal2 429 -1920 429 -1920 0 net=7241
rlabel metal2 68 -1922 68 -1922 0 net=2657
rlabel metal2 240 -1922 240 -1922 0 net=2561
rlabel metal2 317 -1922 317 -1922 0 net=4343
rlabel metal2 359 -1922 359 -1922 0 net=1509
rlabel metal2 590 -1922 590 -1922 0 net=3849
rlabel metal2 772 -1922 772 -1922 0 net=5957
rlabel metal2 54 -1924 54 -1924 0 net=291
rlabel metal2 107 -1924 107 -1924 0 net=1794
rlabel metal2 320 -1924 320 -1924 0 net=4477
rlabel metal2 779 -1924 779 -1924 0 net=5267
rlabel metal2 107 -1926 107 -1926 0 net=1711
rlabel metal2 247 -1926 247 -1926 0 net=3399
rlabel metal2 821 -1926 821 -1926 0 net=5801
rlabel metal2 121 -1928 121 -1928 0 net=3611
rlabel metal2 460 -1928 460 -1928 0 net=7195
rlabel metal2 170 -1930 170 -1930 0 net=2097
rlabel metal2 492 -1930 492 -1930 0 net=7509
rlabel metal2 569 -1932 569 -1932 0 net=3745
rlabel metal2 954 -1932 954 -1932 0 net=7231
rlabel metal2 569 -1934 569 -1934 0 net=6281
rlabel metal2 576 -1936 576 -1936 0 net=4793
rlabel metal2 814 -1938 814 -1938 0 net=5185
rlabel metal2 870 -1940 870 -1940 0 net=5913
rlabel metal2 611 -1942 611 -1942 0 net=7033
rlabel metal2 611 -1944 611 -1944 0 net=3955
rlabel metal2 681 -1946 681 -1946 0 net=4503
rlabel metal2 716 -1948 716 -1948 0 net=4757
rlabel metal2 800 -1950 800 -1950 0 net=5475
rlabel metal2 905 -1952 905 -1952 0 net=6115
rlabel metal2 1017 -1954 1017 -1954 0 net=6585
rlabel metal2 1122 -1956 1122 -1956 0 net=7173
rlabel metal2 586 -1958 586 -1958 0 net=7461
rlabel metal2 2 -1969 2 -1969 0 net=5601
rlabel metal2 674 -1969 674 -1969 0 net=7232
rlabel metal2 964 -1969 964 -1969 0 net=7348
rlabel metal2 1157 -1969 1157 -1969 0 net=7313
rlabel metal2 1157 -1969 1157 -1969 0 net=7313
rlabel metal2 1164 -1969 1164 -1969 0 net=5720
rlabel metal2 9 -1971 9 -1971 0 net=3416
rlabel metal2 142 -1971 142 -1971 0 net=1058
rlabel metal2 310 -1971 310 -1971 0 net=1636
rlabel metal2 320 -1971 320 -1971 0 net=1820
rlabel metal2 373 -1971 373 -1971 0 net=2287
rlabel metal2 401 -1971 401 -1971 0 net=4765
rlabel metal2 702 -1971 702 -1971 0 net=6060
rlabel metal2 9 -1973 9 -1973 0 net=5413
rlabel metal2 184 -1973 184 -1973 0 net=1020
rlabel metal2 499 -1973 499 -1973 0 net=2956
rlabel metal2 702 -1973 702 -1973 0 net=5171
rlabel metal2 758 -1973 758 -1973 0 net=6424
rlabel metal2 1094 -1973 1094 -1973 0 net=7243
rlabel metal2 16 -1975 16 -1975 0 net=3252
rlabel metal2 282 -1975 282 -1975 0 net=464
rlabel metal2 464 -1975 464 -1975 0 net=2945
rlabel metal2 499 -1975 499 -1975 0 net=7546
rlabel metal2 37 -1977 37 -1977 0 net=2216
rlabel metal2 184 -1977 184 -1977 0 net=1859
rlabel metal2 331 -1977 331 -1977 0 net=2098
rlabel metal2 408 -1977 408 -1977 0 net=3933
rlabel metal2 464 -1977 464 -1977 0 net=3867
rlabel metal2 569 -1977 569 -1977 0 net=4758
rlabel metal2 737 -1977 737 -1977 0 net=6173
rlabel metal2 919 -1977 919 -1977 0 net=6432
rlabel metal2 1027 -1977 1027 -1977 0 net=6780
rlabel metal2 37 -1979 37 -1979 0 net=3199
rlabel metal2 191 -1979 191 -1979 0 net=1384
rlabel metal2 373 -1979 373 -1979 0 net=3213
rlabel metal2 394 -1979 394 -1979 0 net=4639
rlabel metal2 716 -1979 716 -1979 0 net=5477
rlabel metal2 891 -1979 891 -1979 0 net=6239
rlabel metal2 954 -1979 954 -1979 0 net=6595
rlabel metal2 968 -1979 968 -1979 0 net=6553
rlabel metal2 996 -1979 996 -1979 0 net=7175
rlabel metal2 16 -1981 16 -1981 0 net=4837
rlabel metal2 198 -1981 198 -1981 0 net=1424
rlabel metal2 481 -1981 481 -1981 0 net=6590
rlabel metal2 1073 -1981 1073 -1981 0 net=7395
rlabel metal2 51 -1983 51 -1983 0 net=2562
rlabel metal2 243 -1983 243 -1983 0 net=5369
rlabel metal2 758 -1983 758 -1983 0 net=5535
rlabel metal2 800 -1983 800 -1983 0 net=5885
rlabel metal2 919 -1983 919 -1983 0 net=6283
rlabel metal2 968 -1983 968 -1983 0 net=6663
rlabel metal2 1010 -1983 1010 -1983 0 net=7367
rlabel metal2 54 -1985 54 -1985 0 net=5118
rlabel metal2 761 -1985 761 -1985 0 net=7510
rlabel metal2 1059 -1985 1059 -1985 0 net=5319
rlabel metal2 58 -1987 58 -1987 0 net=2541
rlabel metal2 488 -1987 488 -1987 0 net=5958
rlabel metal2 786 -1987 786 -1987 0 net=5915
rlabel metal2 940 -1987 940 -1987 0 net=6507
rlabel metal2 982 -1987 982 -1987 0 net=7035
rlabel metal2 1073 -1987 1073 -1987 0 net=7135
rlabel metal2 58 -1989 58 -1989 0 net=4119
rlabel metal2 408 -1989 408 -1989 0 net=2082
rlabel metal2 429 -1989 429 -1989 0 net=2359
rlabel metal2 502 -1989 502 -1989 0 net=4537
rlabel metal2 677 -1989 677 -1989 0 net=6615
rlabel metal2 982 -1989 982 -1989 0 net=6741
rlabel metal2 1087 -1989 1087 -1989 0 net=5589
rlabel metal2 65 -1991 65 -1991 0 net=812
rlabel metal2 100 -1991 100 -1991 0 net=1673
rlabel metal2 310 -1991 310 -1991 0 net=3677
rlabel metal2 604 -1991 604 -1991 0 net=6722
rlabel metal2 23 -1993 23 -1993 0 net=1232
rlabel metal2 110 -1993 110 -1993 0 net=2836
rlabel metal2 513 -1993 513 -1993 0 net=2718
rlabel metal2 569 -1993 569 -1993 0 net=3957
rlabel metal2 744 -1993 744 -1993 0 net=4689
rlabel metal2 842 -1993 842 -1993 0 net=6587
rlabel metal2 1101 -1993 1101 -1993 0 net=7411
rlabel metal2 23 -1995 23 -1995 0 net=4575
rlabel metal2 520 -1995 520 -1995 0 net=6482
rlabel metal2 947 -1995 947 -1995 0 net=6575
rlabel metal2 1017 -1995 1017 -1995 0 net=6861
rlabel metal2 1108 -1995 1108 -1995 0 net=7449
rlabel metal2 44 -1997 44 -1997 0 net=1981
rlabel metal2 68 -1997 68 -1997 0 net=4886
rlabel metal2 772 -1997 772 -1997 0 net=5871
rlabel metal2 849 -1997 849 -1997 0 net=6161
rlabel metal2 898 -1997 898 -1997 0 net=6725
rlabel metal2 1066 -1997 1066 -1997 0 net=7079
rlabel metal2 72 -1999 72 -1999 0 net=2658
rlabel metal2 835 -1999 835 -1999 0 net=5991
rlabel metal2 971 -1999 971 -1999 0 net=1
rlabel metal2 989 -1999 989 -1999 0 net=6657
rlabel metal2 1031 -1999 1031 -1999 0 net=6681
rlabel metal2 1080 -1999 1080 -1999 0 net=7159
rlabel metal2 72 -2001 72 -2001 0 net=1713
rlabel metal2 114 -2001 114 -2001 0 net=3347
rlabel metal2 478 -2001 478 -2001 0 net=6337
rlabel metal2 877 -2001 877 -2001 0 net=6013
rlabel metal2 1003 -2001 1003 -2001 0 net=6831
rlabel metal2 1115 -2001 1115 -2001 0 net=7463
rlabel metal2 86 -2003 86 -2003 0 net=1739
rlabel metal2 142 -2003 142 -2003 0 net=1175
rlabel metal2 282 -2003 282 -2003 0 net=3773
rlabel metal2 506 -2003 506 -2003 0 net=3335
rlabel metal2 926 -2003 926 -2003 0 net=7013
rlabel metal2 86 -2005 86 -2005 0 net=4594
rlabel metal2 576 -2005 576 -2005 0 net=4795
rlabel metal2 1031 -2005 1031 -2005 0 net=7383
rlabel metal2 44 -2007 44 -2007 0 net=2515
rlabel metal2 579 -2007 579 -2007 0 net=5186
rlabel metal2 856 -2007 856 -2007 0 net=6393
rlabel metal2 1136 -2007 1136 -2007 0 net=5591
rlabel metal2 51 -2009 51 -2009 0 net=4393
rlabel metal2 856 -2009 856 -2009 0 net=6117
rlabel metal2 89 -2011 89 -2011 0 net=905
rlabel metal2 117 -2011 117 -2011 0 net=1086
rlabel metal2 226 -2011 226 -2011 0 net=1146
rlabel metal2 317 -2011 317 -2011 0 net=1835
rlabel metal2 450 -2011 450 -2011 0 net=2763
rlabel metal2 534 -2011 534 -2011 0 net=6499
rlabel metal2 93 -2013 93 -2013 0 net=4616
rlabel metal2 905 -2013 905 -2013 0 net=6251
rlabel metal2 93 -2015 93 -2015 0 net=4092
rlabel metal2 338 -2015 338 -2015 0 net=4345
rlabel metal2 611 -2015 611 -2015 0 net=4087
rlabel metal2 709 -2015 709 -2015 0 net=5249
rlabel metal2 30 -2017 30 -2017 0 net=3153
rlabel metal2 471 -2017 471 -2017 0 net=3477
rlabel metal2 562 -2017 562 -2017 0 net=4505
rlabel metal2 751 -2017 751 -2017 0 net=6025
rlabel metal2 30 -2019 30 -2019 0 net=1511
rlabel metal2 534 -2019 534 -2019 0 net=3851
rlabel metal2 597 -2019 597 -2019 0 net=4133
rlabel metal2 681 -2019 681 -2019 0 net=4675
rlabel metal2 751 -2019 751 -2019 0 net=5269
rlabel metal2 114 -2021 114 -2021 0 net=7023
rlabel metal2 432 -2021 432 -2021 0 net=3977
rlabel metal2 625 -2021 625 -2021 0 net=4479
rlabel metal2 765 -2021 765 -2021 0 net=5803
rlabel metal2 121 -2023 121 -2023 0 net=3613
rlabel metal2 541 -2023 541 -2023 0 net=3747
rlabel metal2 632 -2023 632 -2023 0 net=4259
rlabel metal2 660 -2023 660 -2023 0 net=4320
rlabel metal2 821 -2023 821 -2023 0 net=5855
rlabel metal2 103 -2025 103 -2025 0 net=4697
rlabel metal2 863 -2025 863 -2025 0 net=7270
rlabel metal2 121 -2027 121 -2027 0 net=4413
rlabel metal2 1185 -2027 1185 -2027 0 net=6563
rlabel metal2 128 -2029 128 -2029 0 net=2378
rlabel metal2 583 -2029 583 -2029 0 net=5217
rlabel metal2 152 -2031 152 -2031 0 net=6015
rlabel metal2 170 -2033 170 -2033 0 net=2811
rlabel metal2 548 -2033 548 -2033 0 net=3969
rlabel metal2 639 -2033 639 -2033 0 net=4273
rlabel metal2 149 -2035 149 -2035 0 net=1359
rlabel metal2 177 -2035 177 -2035 0 net=1159
rlabel metal2 226 -2035 226 -2035 0 net=1621
rlabel metal2 618 -2035 618 -2035 0 net=6873
rlabel metal2 128 -2037 128 -2037 0 net=2237
rlabel metal2 177 -2037 177 -2037 0 net=3327
rlabel metal2 191 -2039 191 -2039 0 net=1059
rlabel metal2 247 -2039 247 -2039 0 net=3401
rlabel metal2 653 -2039 653 -2039 0 net=5784
rlabel metal2 198 -2041 198 -2041 0 net=2819
rlabel metal2 807 -2041 807 -2041 0 net=5825
rlabel metal2 205 -2043 205 -2043 0 net=1607
rlabel metal2 268 -2043 268 -2043 0 net=2047
rlabel metal2 828 -2043 828 -2043 0 net=7197
rlabel metal2 156 -2045 156 -2045 0 net=1123
rlabel metal2 233 -2045 233 -2045 0 net=2139
rlabel metal2 723 -2045 723 -2045 0 net=4741
rlabel metal2 79 -2047 79 -2047 0 net=1957
rlabel metal2 233 -2047 233 -2047 0 net=1403
rlabel metal2 723 -2047 723 -2047 0 net=5483
rlabel metal2 79 -2049 79 -2049 0 net=1457
rlabel metal2 352 -2049 352 -2049 0 net=3241
rlabel metal2 555 -2049 555 -2049 0 net=5441
rlabel metal2 247 -2051 247 -2051 0 net=2339
rlabel metal2 555 -2051 555 -2051 0 net=1745
rlabel metal2 254 -2053 254 -2053 0 net=1727
rlabel metal2 296 -2053 296 -2053 0 net=1507
rlabel metal2 422 -2053 422 -2053 0 net=3271
rlabel metal2 138 -2055 138 -2055 0 net=2113
rlabel metal2 436 -2055 436 -2055 0 net=2511
rlabel metal2 219 -2057 219 -2057 0 net=1697
rlabel metal2 275 -2057 275 -2057 0 net=3693
rlabel metal2 436 -2057 436 -2057 0 net=2071
rlabel metal2 89 -2059 89 -2059 0 net=2837
rlabel metal2 219 -2061 219 -2061 0 net=3033
rlabel metal2 2 -2072 2 -2072 0 net=5602
rlabel metal2 103 -2072 103 -2072 0 net=4690
rlabel metal2 789 -2072 789 -2072 0 net=7396
rlabel metal2 1136 -2072 1136 -2072 0 net=6564
rlabel metal2 30 -2074 30 -2074 0 net=1512
rlabel metal2 247 -2074 247 -2074 0 net=2340
rlabel metal2 394 -2074 394 -2074 0 net=4640
rlabel metal2 621 -2074 621 -2074 0 net=5886
rlabel metal2 817 -2074 817 -2074 0 net=6554
rlabel metal2 1010 -2074 1010 -2074 0 net=7369
rlabel metal2 1010 -2074 1010 -2074 0 net=7369
rlabel metal2 1108 -2074 1108 -2074 0 net=7451
rlabel metal2 1108 -2074 1108 -2074 0 net=7451
rlabel metal2 1122 -2074 1122 -2074 0 net=5593
rlabel metal2 30 -2076 30 -2076 0 net=5107
rlabel metal2 93 -2076 93 -2076 0 net=182
rlabel metal2 166 -2076 166 -2076 0 net=7176
rlabel metal2 1139 -2076 1139 -2076 0 net=7314
rlabel metal2 37 -2078 37 -2078 0 net=3200
rlabel metal2 394 -2078 394 -2078 0 net=3479
rlabel metal2 481 -2078 481 -2078 0 net=2512
rlabel metal2 562 -2078 562 -2078 0 net=4507
rlabel metal2 576 -2078 576 -2078 0 net=6014
rlabel metal2 975 -2078 975 -2078 0 net=6683
rlabel metal2 65 -2080 65 -2080 0 net=1982
rlabel metal2 156 -2080 156 -2080 0 net=1958
rlabel metal2 509 -2080 509 -2080 0 net=4274
rlabel metal2 653 -2080 653 -2080 0 net=7511
rlabel metal2 65 -2082 65 -2082 0 net=2115
rlabel metal2 387 -2082 387 -2082 0 net=1508
rlabel metal2 492 -2082 492 -2082 0 net=2946
rlabel metal2 562 -2082 562 -2082 0 net=3979
rlabel metal2 600 -2082 600 -2082 0 net=4260
rlabel metal2 639 -2082 639 -2082 0 net=4796
rlabel metal2 72 -2084 72 -2084 0 net=1715
rlabel metal2 72 -2084 72 -2084 0 net=1715
rlabel metal2 86 -2084 86 -2084 0 net=1741
rlabel metal2 138 -2084 138 -2084 0 net=5442
rlabel metal2 863 -2084 863 -2084 0 net=5590
rlabel metal2 37 -2086 37 -2086 0 net=5103
rlabel metal2 142 -2086 142 -2086 0 net=1176
rlabel metal2 614 -2086 614 -2086 0 net=619
rlabel metal2 100 -2088 100 -2088 0 net=1675
rlabel metal2 254 -2088 254 -2088 0 net=1698
rlabel metal2 387 -2088 387 -2088 0 net=2765
rlabel metal2 457 -2088 457 -2088 0 net=2543
rlabel metal2 576 -2088 576 -2088 0 net=4481
rlabel metal2 632 -2088 632 -2088 0 net=4699
rlabel metal2 695 -2088 695 -2088 0 net=5536
rlabel metal2 793 -2088 793 -2088 0 net=4743
rlabel metal2 100 -2090 100 -2090 0 net=4655
rlabel metal2 170 -2090 170 -2090 0 net=1360
rlabel metal2 254 -2090 254 -2090 0 net=1729
rlabel metal2 401 -2090 401 -2090 0 net=3695
rlabel metal2 579 -2090 579 -2090 0 net=4088
rlabel metal2 618 -2090 618 -2090 0 net=4767
rlabel metal2 695 -2090 695 -2090 0 net=6577
rlabel metal2 107 -2092 107 -2092 0 net=2
rlabel metal2 117 -2092 117 -2092 0 net=3774
rlabel metal2 289 -2092 289 -2092 0 net=3155
rlabel metal2 401 -2092 401 -2092 0 net=3869
rlabel metal2 467 -2092 467 -2092 0 net=7571
rlabel metal2 58 -2094 58 -2094 0 net=4121
rlabel metal2 114 -2094 114 -2094 0 net=2288
rlabel metal2 429 -2094 429 -2094 0 net=2361
rlabel metal2 457 -2094 457 -2094 0 net=4539
rlabel metal2 656 -2094 656 -2094 0 net=5250
rlabel metal2 716 -2094 716 -2094 0 net=5479
rlabel metal2 863 -2094 863 -2094 0 net=6395
rlabel metal2 947 -2094 947 -2094 0 net=7413
rlabel metal2 23 -2096 23 -2096 0 net=4577
rlabel metal2 142 -2096 142 -2096 0 net=1405
rlabel metal2 240 -2096 240 -2096 0 net=1651
rlabel metal2 373 -2096 373 -2096 0 net=3215
rlabel metal2 408 -2096 408 -2096 0 net=5443
rlabel metal2 660 -2096 660 -2096 0 net=6588
rlabel metal2 877 -2096 877 -2096 0 net=6597
rlabel metal2 23 -2098 23 -2098 0 net=7017
rlabel metal2 96 -2098 96 -2098 0 net=2731
rlabel metal2 429 -2098 429 -2098 0 net=2073
rlabel metal2 443 -2098 443 -2098 0 net=2838
rlabel metal2 625 -2098 625 -2098 0 net=5371
rlabel metal2 709 -2098 709 -2098 0 net=5827
rlabel metal2 842 -2098 842 -2098 0 net=6241
rlabel metal2 926 -2098 926 -2098 0 net=6743
rlabel metal2 149 -2100 149 -2100 0 net=601
rlabel metal2 583 -2100 583 -2100 0 net=6026
rlabel metal2 933 -2100 933 -2100 0 net=6501
rlabel metal2 982 -2100 982 -2100 0 net=7081
rlabel metal2 44 -2102 44 -2102 0 net=2517
rlabel metal2 156 -2102 156 -2102 0 net=3035
rlabel metal2 233 -2102 233 -2102 0 net=1837
rlabel metal2 345 -2102 345 -2102 0 net=2813
rlabel metal2 443 -2102 443 -2102 0 net=3123
rlabel metal2 716 -2102 716 -2102 0 net=5873
rlabel metal2 807 -2102 807 -2102 0 net=5857
rlabel metal2 884 -2102 884 -2102 0 net=6617
rlabel metal2 1066 -2102 1066 -2102 0 net=7161
rlabel metal2 44 -2104 44 -2104 0 net=5409
rlabel metal2 737 -2104 737 -2104 0 net=6175
rlabel metal2 772 -2104 772 -2104 0 net=5917
rlabel metal2 821 -2104 821 -2104 0 net=6253
rlabel metal2 933 -2104 933 -2104 0 net=6863
rlabel metal2 51 -2106 51 -2106 0 net=4395
rlabel metal2 261 -2106 261 -2106 0 net=1608
rlabel metal2 338 -2106 338 -2106 0 net=7025
rlabel metal2 1017 -2106 1017 -2106 0 net=7465
rlabel metal2 16 -2108 16 -2108 0 net=4839
rlabel metal2 173 -2108 173 -2108 0 net=4676
rlabel metal2 737 -2108 737 -2108 0 net=5805
rlabel metal2 891 -2108 891 -2108 0 net=6665
rlabel metal2 110 -2110 110 -2110 0 net=5997
rlabel metal2 898 -2110 898 -2110 0 net=6727
rlabel metal2 968 -2110 968 -2110 0 net=7384
rlabel metal2 184 -2112 184 -2112 0 net=1861
rlabel metal2 303 -2112 303 -2112 0 net=5009
rlabel metal2 583 -2112 583 -2112 0 net=4135
rlabel metal2 660 -2112 660 -2112 0 net=3085
rlabel metal2 667 -2112 667 -2112 0 net=5173
rlabel metal2 744 -2112 744 -2112 0 net=5271
rlabel metal2 814 -2112 814 -2112 0 net=6093
rlabel metal2 905 -2112 905 -2112 0 net=7037
rlabel metal2 184 -2114 184 -2114 0 net=3853
rlabel metal2 674 -2114 674 -2114 0 net=5485
rlabel metal2 751 -2114 751 -2114 0 net=5219
rlabel metal2 814 -2114 814 -2114 0 net=6119
rlabel metal2 866 -2114 866 -2114 0 net=3587
rlabel metal2 205 -2116 205 -2116 0 net=1125
rlabel metal2 338 -2116 338 -2116 0 net=6463
rlabel metal2 681 -2116 681 -2116 0 net=6017
rlabel metal2 856 -2116 856 -2116 0 net=6833
rlabel metal2 1031 -2116 1031 -2116 0 net=7517
rlabel metal2 205 -2118 205 -2118 0 net=1623
rlabel metal2 261 -2118 261 -2118 0 net=7349
rlabel metal2 702 -2118 702 -2118 0 net=6163
rlabel metal2 1003 -2118 1003 -2118 0 net=5321
rlabel metal2 79 -2120 79 -2120 0 net=1459
rlabel metal2 268 -2120 268 -2120 0 net=2048
rlabel metal2 345 -2120 345 -2120 0 net=3273
rlabel metal2 471 -2120 471 -2120 0 net=3971
rlabel metal2 723 -2120 723 -2120 0 net=5993
rlabel metal2 849 -2120 849 -2120 0 net=7015
rlabel metal2 79 -2122 79 -2122 0 net=1795
rlabel metal2 548 -2122 548 -2122 0 net=2563
rlabel metal2 730 -2122 730 -2122 0 net=6339
rlabel metal2 835 -2122 835 -2122 0 net=6875
rlabel metal2 1052 -2122 1052 -2122 0 net=2309
rlabel metal2 128 -2124 128 -2124 0 net=2239
rlabel metal2 352 -2124 352 -2124 0 net=3243
rlabel metal2 478 -2124 478 -2124 0 net=6658
rlabel metal2 128 -2126 128 -2126 0 net=3329
rlabel metal2 212 -2126 212 -2126 0 net=1160
rlabel metal2 352 -2126 352 -2126 0 net=3403
rlabel metal2 597 -2126 597 -2126 0 net=1069
rlabel metal2 9 -2128 9 -2128 0 net=5414
rlabel metal2 730 -2128 730 -2128 0 net=7199
rlabel metal2 870 -2128 870 -2128 0 net=6509
rlabel metal2 989 -2128 989 -2128 0 net=7137
rlabel metal2 177 -2130 177 -2130 0 net=1061
rlabel metal2 212 -2130 212 -2130 0 net=2141
rlabel metal2 366 -2130 366 -2130 0 net=3349
rlabel metal2 485 -2130 485 -2130 0 net=6885
rlabel metal2 121 -2132 121 -2132 0 net=4415
rlabel metal2 268 -2132 268 -2132 0 net=3337
rlabel metal2 828 -2132 828 -2132 0 net=6285
rlabel metal2 117 -2134 117 -2134 0 net=1871
rlabel metal2 275 -2134 275 -2134 0 net=1747
rlabel metal2 919 -2134 919 -2134 0 net=7245
rlabel metal2 310 -2136 310 -2136 0 net=3679
rlabel metal2 555 -2136 555 -2136 0 net=3959
rlabel metal2 198 -2138 198 -2138 0 net=2821
rlabel metal2 359 -2138 359 -2138 0 net=3935
rlabel metal2 464 -2138 464 -2138 0 net=4165
rlabel metal2 198 -2140 198 -2140 0 net=2473
rlabel metal2 366 -2140 366 -2140 0 net=3615
rlabel metal2 415 -2142 415 -2142 0 net=4347
rlabel metal2 520 -2144 520 -2144 0 net=3749
rlabel metal2 604 -2144 604 -2144 0 net=5007
rlabel metal2 541 -2146 541 -2146 0 net=3921
rlabel metal2 23 -2157 23 -2157 0 net=7018
rlabel metal2 124 -2157 124 -2157 0 net=5010
rlabel metal2 317 -2157 317 -2157 0 net=1127
rlabel metal2 331 -2157 331 -2157 0 net=2240
rlabel metal2 975 -2157 975 -2157 0 net=6684
rlabel metal2 1066 -2157 1066 -2157 0 net=7163
rlabel metal2 1066 -2157 1066 -2157 0 net=7163
rlabel metal2 1101 -2157 1101 -2157 0 net=7452
rlabel metal2 37 -2159 37 -2159 0 net=5104
rlabel metal2 103 -2159 103 -2159 0 net=3036
rlabel metal2 198 -2159 198 -2159 0 net=2475
rlabel metal2 324 -2159 324 -2159 0 net=3217
rlabel metal2 387 -2159 387 -2159 0 net=2766
rlabel metal2 509 -2159 509 -2159 0 net=7016
rlabel metal2 933 -2159 933 -2159 0 net=6865
rlabel metal2 982 -2159 982 -2159 0 net=7083
rlabel metal2 1104 -2159 1104 -2159 0 net=5594
rlabel metal2 37 -2161 37 -2161 0 net=1743
rlabel metal2 93 -2161 93 -2161 0 net=7350
rlabel metal2 275 -2161 275 -2161 0 net=1748
rlabel metal2 485 -2161 485 -2161 0 net=4136
rlabel metal2 597 -2161 597 -2161 0 net=6164
rlabel metal2 786 -2161 786 -2161 0 net=6094
rlabel metal2 933 -2161 933 -2161 0 net=7573
rlabel metal2 30 -2163 30 -2163 0 net=5108
rlabel metal2 100 -2163 100 -2163 0 net=1407
rlabel metal2 198 -2163 198 -2163 0 net=1677
rlabel metal2 254 -2163 254 -2163 0 net=1730
rlabel metal2 513 -2163 513 -2163 0 net=6578
rlabel metal2 702 -2163 702 -2163 0 net=5807
rlabel metal2 786 -2163 786 -2163 0 net=6619
rlabel metal2 943 -2163 943 -2163 0 net=3588
rlabel metal2 30 -2165 30 -2165 0 net=7609
rlabel metal2 597 -2165 597 -2165 0 net=4701
rlabel metal2 639 -2165 639 -2165 0 net=5487
rlabel metal2 688 -2165 688 -2165 0 net=7246
rlabel metal2 982 -2165 982 -2165 0 net=5323
rlabel metal2 51 -2167 51 -2167 0 net=4841
rlabel metal2 226 -2167 226 -2167 0 net=1461
rlabel metal2 226 -2167 226 -2167 0 net=1461
rlabel metal2 233 -2167 233 -2167 0 net=1838
rlabel metal2 513 -2167 513 -2167 0 net=3923
rlabel metal2 611 -2167 611 -2167 0 net=6502
rlabel metal2 1003 -2167 1003 -2167 0 net=2311
rlabel metal2 44 -2169 44 -2169 0 net=5411
rlabel metal2 65 -2169 65 -2169 0 net=2117
rlabel metal2 289 -2169 289 -2169 0 net=3156
rlabel metal2 541 -2169 541 -2169 0 net=4167
rlabel metal2 611 -2169 611 -2169 0 net=5433
rlabel metal2 842 -2169 842 -2169 0 net=6243
rlabel metal2 58 -2171 58 -2171 0 net=4579
rlabel metal2 72 -2171 72 -2171 0 net=1716
rlabel metal2 138 -2171 138 -2171 0 net=4991
rlabel metal2 614 -2171 614 -2171 0 net=7499
rlabel metal2 919 -2171 919 -2171 0 net=7519
rlabel metal2 58 -2173 58 -2173 0 net=5449
rlabel metal2 408 -2173 408 -2173 0 net=2814
rlabel metal2 632 -2173 632 -2173 0 net=5829
rlabel metal2 842 -2173 842 -2173 0 net=7027
rlabel metal2 72 -2175 72 -2175 0 net=3855
rlabel metal2 240 -2175 240 -2175 0 net=1653
rlabel metal2 254 -2175 254 -2175 0 net=3339
rlabel metal2 289 -2175 289 -2175 0 net=3481
rlabel metal2 401 -2175 401 -2175 0 net=3871
rlabel metal2 429 -2175 429 -2175 0 net=2074
rlabel metal2 646 -2175 646 -2175 0 net=5445
rlabel metal2 96 -2177 96 -2177 0 net=6629
rlabel metal2 205 -2177 205 -2177 0 net=1625
rlabel metal2 268 -2177 268 -2177 0 net=1777
rlabel metal2 96 -2179 96 -2179 0 net=248
rlabel metal2 674 -2179 674 -2179 0 net=6019
rlabel metal2 688 -2179 688 -2179 0 net=5999
rlabel metal2 114 -2181 114 -2181 0 net=1881
rlabel metal2 296 -2181 296 -2181 0 net=3079
rlabel metal2 355 -2181 355 -2181 0 net=5008
rlabel metal2 646 -2181 646 -2181 0 net=5175
rlabel metal2 681 -2181 681 -2181 0 net=6177
rlabel metal2 114 -2183 114 -2183 0 net=1873
rlabel metal2 131 -2183 131 -2183 0 net=3936
rlabel metal2 366 -2183 366 -2183 0 net=3616
rlabel metal2 401 -2183 401 -2183 0 net=2363
rlabel metal2 464 -2183 464 -2183 0 net=2545
rlabel metal2 506 -2183 506 -2183 0 net=3961
rlabel metal2 604 -2183 604 -2183 0 net=4665
rlabel metal2 751 -2183 751 -2183 0 net=5221
rlabel metal2 121 -2185 121 -2185 0 net=3124
rlabel metal2 457 -2185 457 -2185 0 net=4541
rlabel metal2 656 -2185 656 -2185 0 net=6834
rlabel metal2 135 -2187 135 -2187 0 net=4397
rlabel metal2 282 -2187 282 -2187 0 net=1863
rlabel metal2 310 -2187 310 -2187 0 net=2823
rlabel metal2 373 -2187 373 -2187 0 net=2733
rlabel metal2 443 -2187 443 -2187 0 net=3696
rlabel metal2 499 -2187 499 -2187 0 net=4141
rlabel metal2 691 -2187 691 -2187 0 net=5480
rlabel metal2 856 -2187 856 -2187 0 net=7039
rlabel metal2 79 -2189 79 -2189 0 net=1797
rlabel metal2 310 -2189 310 -2189 0 net=3405
rlabel metal2 359 -2189 359 -2189 0 net=2565
rlabel metal2 695 -2189 695 -2189 0 net=1070
rlabel metal2 79 -2191 79 -2191 0 net=3330
rlabel metal2 142 -2191 142 -2191 0 net=2519
rlabel metal2 163 -2191 163 -2191 0 net=4657
rlabel metal2 709 -2191 709 -2191 0 net=6341
rlabel metal2 800 -2191 800 -2191 0 net=5859
rlabel metal2 905 -2191 905 -2191 0 net=7513
rlabel metal2 44 -2193 44 -2193 0 net=6933
rlabel metal2 163 -2193 163 -2193 0 net=2451
rlabel metal2 751 -2193 751 -2193 0 net=6511
rlabel metal2 86 -2195 86 -2195 0 net=2369
rlabel metal2 170 -2195 170 -2195 0 net=1481
rlabel metal2 320 -2195 320 -2195 0 net=7141
rlabel metal2 870 -2195 870 -2195 0 net=7467
rlabel metal2 170 -2197 170 -2197 0 net=1063
rlabel metal2 180 -2197 180 -2197 0 net=6835
rlabel metal2 548 -2197 548 -2197 0 net=4509
rlabel metal2 653 -2197 653 -2197 0 net=5918
rlabel metal2 779 -2197 779 -2197 0 net=6255
rlabel metal2 954 -2197 954 -2197 0 net=6611
rlabel metal2 177 -2199 177 -2199 0 net=2142
rlabel metal2 219 -2199 219 -2199 0 net=3275
rlabel metal2 373 -2199 373 -2199 0 net=3973
rlabel metal2 590 -2199 590 -2199 0 net=5373
rlabel metal2 758 -2199 758 -2199 0 net=6599
rlabel metal2 107 -2201 107 -2201 0 net=4123
rlabel metal2 380 -2201 380 -2201 0 net=4483
rlabel metal2 618 -2201 618 -2201 0 net=4769
rlabel metal2 772 -2201 772 -2201 0 net=6287
rlabel metal2 877 -2201 877 -2201 0 net=7415
rlabel metal2 107 -2203 107 -2203 0 net=1327
rlabel metal2 387 -2203 387 -2203 0 net=3245
rlabel metal2 450 -2203 450 -2203 0 net=4617
rlabel metal2 618 -2203 618 -2203 0 net=4745
rlabel metal2 807 -2203 807 -2203 0 net=6121
rlabel metal2 821 -2203 821 -2203 0 net=6667
rlabel metal2 191 -2205 191 -2205 0 net=4416
rlabel metal2 670 -2205 670 -2205 0 net=7477
rlabel metal2 191 -2207 191 -2207 0 net=3981
rlabel metal2 793 -2207 793 -2207 0 net=6877
rlabel metal2 205 -2209 205 -2209 0 net=3087
rlabel metal2 814 -2209 814 -2209 0 net=6729
rlabel metal2 212 -2211 212 -2211 0 net=3819
rlabel metal2 471 -2211 471 -2211 0 net=3751
rlabel metal2 660 -2211 660 -2211 0 net=5875
rlabel metal2 828 -2211 828 -2211 0 net=6887
rlabel metal2 338 -2213 338 -2213 0 net=6465
rlabel metal2 765 -2213 765 -2213 0 net=6523
rlabel metal2 338 -2215 338 -2215 0 net=7483
rlabel metal2 835 -2215 835 -2215 0 net=6745
rlabel metal2 422 -2217 422 -2217 0 net=3351
rlabel metal2 485 -2217 485 -2217 0 net=7619
rlabel metal2 415 -2219 415 -2219 0 net=4349
rlabel metal2 436 -2219 436 -2219 0 net=5995
rlabel metal2 912 -2219 912 -2219 0 net=7139
rlabel metal2 415 -2221 415 -2221 0 net=3157
rlabel metal2 723 -2221 723 -2221 0 net=6397
rlabel metal2 926 -2221 926 -2221 0 net=7371
rlabel metal2 516 -2223 516 -2223 0 net=2729
rlabel metal2 730 -2223 730 -2223 0 net=7201
rlabel metal2 520 -2225 520 -2225 0 net=3681
rlabel metal2 730 -2225 730 -2225 0 net=5273
rlabel metal2 534 -2227 534 -2227 0 net=3225
rlabel metal2 30 -2238 30 -2238 0 net=7610
rlabel metal2 131 -2238 131 -2238 0 net=7484
rlabel metal2 345 -2238 345 -2238 0 net=4124
rlabel metal2 359 -2238 359 -2238 0 net=2566
rlabel metal2 667 -2238 667 -2238 0 net=6746
rlabel metal2 940 -2238 940 -2238 0 net=5222
rlabel metal2 968 -2238 968 -2238 0 net=6867
rlabel metal2 968 -2238 968 -2238 0 net=6867
rlabel metal2 989 -2238 989 -2238 0 net=2313
rlabel metal2 1017 -2238 1017 -2238 0 net=6613
rlabel metal2 1059 -2238 1059 -2238 0 net=7164
rlabel metal2 44 -2240 44 -2240 0 net=6935
rlabel metal2 51 -2240 51 -2240 0 net=5412
rlabel metal2 93 -2240 93 -2240 0 net=361
rlabel metal2 481 -2240 481 -2240 0 net=5830
rlabel metal2 667 -2240 667 -2240 0 net=6001
rlabel metal2 695 -2240 695 -2240 0 net=6513
rlabel metal2 800 -2240 800 -2240 0 net=5860
rlabel metal2 807 -2240 807 -2240 0 net=6123
rlabel metal2 835 -2240 835 -2240 0 net=7469
rlabel metal2 943 -2240 943 -2240 0 net=5324
rlabel metal2 996 -2240 996 -2240 0 net=7085
rlabel metal2 996 -2240 996 -2240 0 net=7085
rlabel metal2 37 -2242 37 -2242 0 net=1744
rlabel metal2 135 -2242 135 -2242 0 net=4399
rlabel metal2 359 -2242 359 -2242 0 net=3975
rlabel metal2 429 -2242 429 -2242 0 net=2734
rlabel metal2 520 -2242 520 -2242 0 net=3683
rlabel metal2 520 -2242 520 -2242 0 net=3683
rlabel metal2 527 -2242 527 -2242 0 net=5876
rlabel metal2 674 -2242 674 -2242 0 net=6021
rlabel metal2 681 -2242 681 -2242 0 net=6179
rlabel metal2 688 -2242 688 -2242 0 net=6525
rlabel metal2 800 -2242 800 -2242 0 net=7372
rlabel metal2 957 -2242 957 -2242 0 net=6244
rlabel metal2 44 -2244 44 -2244 0 net=5451
rlabel metal2 65 -2244 65 -2244 0 net=4581
rlabel metal2 135 -2244 135 -2244 0 net=4842
rlabel metal2 177 -2244 177 -2244 0 net=1626
rlabel metal2 261 -2244 261 -2244 0 net=2118
rlabel metal2 429 -2244 429 -2244 0 net=3963
rlabel metal2 527 -2244 527 -2244 0 net=4511
rlabel metal2 583 -2244 583 -2244 0 net=4993
rlabel metal2 632 -2244 632 -2244 0 net=5177
rlabel metal2 674 -2244 674 -2244 0 net=6601
rlabel metal2 765 -2244 765 -2244 0 net=6731
rlabel metal2 870 -2244 870 -2244 0 net=7223
rlabel metal2 51 -2246 51 -2246 0 net=1875
rlabel metal2 138 -2246 138 -2246 0 net=283
rlabel metal2 583 -2246 583 -2246 0 net=4703
rlabel metal2 621 -2246 621 -2246 0 net=5865
rlabel metal2 681 -2246 681 -2246 0 net=6467
rlabel metal2 723 -2246 723 -2246 0 net=6399
rlabel metal2 807 -2246 807 -2246 0 net=7029
rlabel metal2 65 -2248 65 -2248 0 net=1409
rlabel metal2 114 -2248 114 -2248 0 net=2521
rlabel metal2 170 -2248 170 -2248 0 net=1065
rlabel metal2 180 -2248 180 -2248 0 net=4099
rlabel metal2 247 -2248 247 -2248 0 net=1655
rlabel metal2 303 -2248 303 -2248 0 net=2476
rlabel metal2 436 -2248 436 -2248 0 net=5996
rlabel metal2 478 -2248 478 -2248 0 net=4495
rlabel metal2 639 -2248 639 -2248 0 net=5489
rlabel metal2 698 -2248 698 -2248 0 net=7140
rlabel metal2 72 -2250 72 -2250 0 net=3856
rlabel metal2 534 -2250 534 -2250 0 net=3227
rlabel metal2 611 -2250 611 -2250 0 net=5435
rlabel metal2 702 -2250 702 -2250 0 net=5809
rlabel metal2 730 -2250 730 -2250 0 net=5274
rlabel metal2 747 -2250 747 -2250 0 net=5446
rlabel metal2 72 -2252 72 -2252 0 net=2453
rlabel metal2 184 -2252 184 -2252 0 net=6630
rlabel metal2 408 -2252 408 -2252 0 net=3873
rlabel metal2 446 -2252 446 -2252 0 net=3352
rlabel metal2 499 -2252 499 -2252 0 net=4143
rlabel metal2 604 -2252 604 -2252 0 net=4667
rlabel metal2 656 -2252 656 -2252 0 net=5579
rlabel metal2 79 -2254 79 -2254 0 net=3821
rlabel metal2 226 -2254 226 -2254 0 net=1462
rlabel metal2 709 -2254 709 -2254 0 net=6343
rlabel metal2 730 -2254 730 -2254 0 net=6289
rlabel metal2 814 -2254 814 -2254 0 net=7203
rlabel metal2 96 -2256 96 -2256 0 net=3253
rlabel metal2 247 -2256 247 -2256 0 net=3247
rlabel metal2 408 -2256 408 -2256 0 net=4169
rlabel metal2 576 -2256 576 -2256 0 net=4619
rlabel metal2 737 -2256 737 -2256 0 net=5785
rlabel metal2 772 -2256 772 -2256 0 net=6257
rlabel metal2 842 -2256 842 -2256 0 net=7479
rlabel metal2 100 -2258 100 -2258 0 net=3483
rlabel metal2 303 -2258 303 -2258 0 net=2109
rlabel metal2 387 -2258 387 -2258 0 net=6069
rlabel metal2 737 -2258 737 -2258 0 net=6621
rlabel metal2 810 -2258 810 -2258 0 net=1
rlabel metal2 107 -2260 107 -2260 0 net=1329
rlabel metal2 156 -2260 156 -2260 0 net=1103
rlabel metal2 471 -2260 471 -2260 0 net=3753
rlabel metal2 740 -2260 740 -2260 0 net=7040
rlabel metal2 863 -2260 863 -2260 0 net=7621
rlabel metal2 107 -2262 107 -2262 0 net=3983
rlabel metal2 198 -2262 198 -2262 0 net=1678
rlabel metal2 310 -2262 310 -2262 0 net=3407
rlabel metal2 366 -2262 366 -2262 0 net=2825
rlabel metal2 492 -2262 492 -2262 0 net=6837
rlabel metal2 744 -2262 744 -2262 0 net=6879
rlabel metal2 856 -2262 856 -2262 0 net=7521
rlabel metal2 124 -2264 124 -2264 0 net=1643
rlabel metal2 198 -2264 198 -2264 0 net=1779
rlabel metal2 275 -2264 275 -2264 0 net=1882
rlabel metal2 779 -2264 779 -2264 0 net=6669
rlabel metal2 149 -2266 149 -2266 0 net=2371
rlabel metal2 205 -2266 205 -2266 0 net=3089
rlabel metal2 205 -2266 205 -2266 0 net=3089
rlabel metal2 212 -2266 212 -2266 0 net=1483
rlabel metal2 254 -2266 254 -2266 0 net=3340
rlabel metal2 653 -2266 653 -2266 0 net=7219
rlabel metal2 149 -2268 149 -2268 0 net=1841
rlabel metal2 219 -2268 219 -2268 0 net=3276
rlabel metal2 786 -2268 786 -2268 0 net=6889
rlabel metal2 163 -2270 163 -2270 0 net=1577
rlabel metal2 793 -2270 793 -2270 0 net=7515
rlabel metal2 184 -2272 184 -2272 0 net=4609
rlabel metal2 268 -2272 268 -2272 0 net=2203
rlabel metal2 828 -2272 828 -2272 0 net=7143
rlabel metal2 219 -2274 219 -2274 0 net=4069
rlabel metal2 443 -2274 443 -2274 0 net=5837
rlabel metal2 849 -2274 849 -2274 0 net=7501
rlabel metal2 93 -2276 93 -2276 0 net=1089
rlabel metal2 877 -2276 877 -2276 0 net=7417
rlabel metal2 233 -2278 233 -2278 0 net=1865
rlabel metal2 310 -2278 310 -2278 0 net=4485
rlabel metal2 877 -2278 877 -2278 0 net=7575
rlabel metal2 275 -2280 275 -2280 0 net=1799
rlabel metal2 296 -2280 296 -2280 0 net=2695
rlabel metal2 282 -2282 282 -2282 0 net=1129
rlabel metal2 324 -2282 324 -2282 0 net=3219
rlabel metal2 317 -2284 317 -2284 0 net=7005
rlabel metal2 324 -2286 324 -2286 0 net=2365
rlabel metal2 331 -2288 331 -2288 0 net=3081
rlabel metal2 331 -2288 331 -2288 0 net=3081
rlabel metal2 345 -2288 345 -2288 0 net=3791
rlabel metal2 366 -2290 366 -2290 0 net=3159
rlabel metal2 121 -2292 121 -2292 0 net=7087
rlabel metal2 121 -2294 121 -2294 0 net=3925
rlabel metal2 401 -2296 401 -2296 0 net=4543
rlabel metal2 422 -2298 422 -2298 0 net=4351
rlabel metal2 555 -2298 555 -2298 0 net=4659
rlabel metal2 422 -2300 422 -2300 0 net=4770
rlabel metal2 464 -2302 464 -2302 0 net=2546
rlabel metal2 590 -2302 590 -2302 0 net=5375
rlabel metal2 464 -2304 464 -2304 0 net=4899
rlabel metal2 590 -2306 590 -2306 0 net=4747
rlabel metal2 562 -2308 562 -2308 0 net=2730
rlabel metal2 471 -2310 471 -2310 0 net=4261
rlabel metal2 51 -2321 51 -2321 0 net=1876
rlabel metal2 187 -2321 187 -2321 0 net=864
rlabel metal2 383 -2321 383 -2321 0 net=4262
rlabel metal2 492 -2321 492 -2321 0 net=7516
rlabel metal2 884 -2321 884 -2321 0 net=5581
rlabel metal2 968 -2321 968 -2321 0 net=6868
rlabel metal2 982 -2321 982 -2321 0 net=2315
rlabel metal2 996 -2321 996 -2321 0 net=7086
rlabel metal2 1038 -2321 1038 -2321 0 net=6614
rlabel metal2 65 -2323 65 -2323 0 net=1410
rlabel metal2 89 -2323 89 -2323 0 net=5786
rlabel metal2 772 -2323 772 -2323 0 net=6259
rlabel metal2 898 -2323 898 -2323 0 net=7419
rlabel metal2 989 -2323 989 -2323 0 net=6007
rlabel metal2 44 -2325 44 -2325 0 net=5453
rlabel metal2 135 -2325 135 -2325 0 net=1131
rlabel metal2 306 -2325 306 -2325 0 net=2673
rlabel metal2 492 -2325 492 -2325 0 net=4355
rlabel metal2 632 -2325 632 -2325 0 net=5178
rlabel metal2 698 -2325 698 -2325 0 net=7224
rlabel metal2 891 -2325 891 -2325 0 net=6125
rlabel metal2 138 -2327 138 -2327 0 net=2696
rlabel metal2 310 -2327 310 -2327 0 net=4486
rlabel metal2 457 -2327 457 -2327 0 net=3792
rlabel metal2 152 -2329 152 -2329 0 net=1656
rlabel metal2 275 -2329 275 -2329 0 net=1800
rlabel metal2 520 -2329 520 -2329 0 net=3685
rlabel metal2 520 -2329 520 -2329 0 net=3685
rlabel metal2 558 -2329 558 -2329 0 net=7144
rlabel metal2 114 -2331 114 -2331 0 net=2523
rlabel metal2 292 -2331 292 -2331 0 net=1225
rlabel metal2 338 -2331 338 -2331 0 net=4400
rlabel metal2 352 -2331 352 -2331 0 net=3408
rlabel metal2 446 -2331 446 -2331 0 net=6022
rlabel metal2 716 -2331 716 -2331 0 net=5811
rlabel metal2 751 -2331 751 -2331 0 net=7471
rlabel metal2 114 -2333 114 -2333 0 net=2647
rlabel metal2 205 -2333 205 -2333 0 net=3091
rlabel metal2 338 -2333 338 -2333 0 net=3161
rlabel metal2 387 -2333 387 -2333 0 net=6070
rlabel metal2 548 -2333 548 -2333 0 net=3229
rlabel metal2 716 -2333 716 -2333 0 net=7205
rlabel metal2 93 -2335 93 -2335 0 net=1091
rlabel metal2 233 -2335 233 -2335 0 net=1867
rlabel metal2 359 -2335 359 -2335 0 net=3976
rlabel metal2 387 -2335 387 -2335 0 net=1479
rlabel metal2 429 -2335 429 -2335 0 net=3964
rlabel metal2 562 -2335 562 -2335 0 net=6180
rlabel metal2 772 -2335 772 -2335 0 net=7623
rlabel metal2 93 -2337 93 -2337 0 net=1843
rlabel metal2 163 -2337 163 -2337 0 net=1579
rlabel metal2 359 -2337 359 -2337 0 net=5839
rlabel metal2 534 -2337 534 -2337 0 net=5377
rlabel metal2 632 -2337 632 -2337 0 net=6003
rlabel metal2 702 -2337 702 -2337 0 net=7221
rlabel metal2 121 -2339 121 -2339 0 net=3927
rlabel metal2 394 -2339 394 -2339 0 net=2827
rlabel metal2 394 -2339 394 -2339 0 net=2827
rlabel metal2 401 -2339 401 -2339 0 net=4545
rlabel metal2 453 -2339 453 -2339 0 net=4641
rlabel metal2 555 -2339 555 -2339 0 net=4661
rlabel metal2 569 -2339 569 -2339 0 net=4748
rlabel metal2 604 -2339 604 -2339 0 net=4621
rlabel metal2 614 -2339 614 -2339 0 net=6400
rlabel metal2 779 -2339 779 -2339 0 net=6671
rlabel metal2 121 -2341 121 -2341 0 net=1485
rlabel metal2 226 -2341 226 -2341 0 net=3255
rlabel metal2 415 -2341 415 -2341 0 net=7088
rlabel metal2 569 -2341 569 -2341 0 net=4669
rlabel metal2 618 -2341 618 -2341 0 net=7576
rlabel metal2 149 -2343 149 -2343 0 net=4649
rlabel metal2 324 -2343 324 -2343 0 net=2367
rlabel metal2 429 -2343 429 -2343 0 net=4901
rlabel metal2 485 -2343 485 -2343 0 net=4353
rlabel metal2 555 -2343 555 -2343 0 net=7119
rlabel metal2 667 -2343 667 -2343 0 net=7503
rlabel metal2 72 -2345 72 -2345 0 net=2454
rlabel metal2 572 -2345 572 -2345 0 net=6514
rlabel metal2 730 -2345 730 -2345 0 net=6291
rlabel metal2 793 -2345 793 -2345 0 net=7523
rlabel metal2 72 -2347 72 -2347 0 net=7007
rlabel metal2 436 -2347 436 -2347 0 net=3875
rlabel metal2 436 -2347 436 -2347 0 net=3875
rlabel metal2 457 -2347 457 -2347 0 net=4145
rlabel metal2 576 -2347 576 -2347 0 net=5490
rlabel metal2 730 -2347 730 -2347 0 net=6623
rlabel metal2 758 -2347 758 -2347 0 net=6733
rlabel metal2 107 -2349 107 -2349 0 net=3985
rlabel metal2 464 -2349 464 -2349 0 net=4513
rlabel metal2 576 -2349 576 -2349 0 net=4705
rlabel metal2 590 -2349 590 -2349 0 net=4995
rlabel metal2 604 -2349 604 -2349 0 net=5867
rlabel metal2 660 -2349 660 -2349 0 net=6603
rlabel metal2 765 -2349 765 -2349 0 net=7481
rlabel metal2 107 -2351 107 -2351 0 net=3221
rlabel metal2 478 -2351 478 -2351 0 net=4497
rlabel metal2 583 -2351 583 -2351 0 net=6527
rlabel metal2 719 -2351 719 -2351 0 net=1
rlabel metal2 156 -2353 156 -2353 0 net=1105
rlabel metal2 226 -2353 226 -2353 0 net=2297
rlabel metal2 236 -2353 236 -2353 0 net=764
rlabel metal2 128 -2355 128 -2355 0 net=4583
rlabel metal2 240 -2355 240 -2355 0 net=4101
rlabel metal2 240 -2355 240 -2355 0 net=4101
rlabel metal2 247 -2355 247 -2355 0 net=3248
rlabel metal2 478 -2355 478 -2355 0 net=6839
rlabel metal2 597 -2355 597 -2355 0 net=5437
rlabel metal2 674 -2355 674 -2355 0 net=6891
rlabel metal2 128 -2357 128 -2357 0 net=4071
rlabel metal2 254 -2357 254 -2357 0 net=4611
rlabel metal2 499 -2357 499 -2357 0 net=3754
rlabel metal2 639 -2357 639 -2357 0 net=6469
rlabel metal2 191 -2359 191 -2359 0 net=2373
rlabel metal2 254 -2359 254 -2359 0 net=4487
rlabel metal2 527 -2359 527 -2359 0 net=2513
rlabel metal2 170 -2361 170 -2361 0 net=1645
rlabel metal2 219 -2361 219 -2361 0 net=2205
rlabel metal2 271 -2361 271 -2361 0 net=3441
rlabel metal2 681 -2361 681 -2361 0 net=6881
rlabel metal2 142 -2363 142 -2363 0 net=1330
rlabel metal2 289 -2363 289 -2363 0 net=5907
rlabel metal2 723 -2363 723 -2363 0 net=6345
rlabel metal2 100 -2365 100 -2365 0 net=3485
rlabel metal2 303 -2365 303 -2365 0 net=2111
rlabel metal2 79 -2367 79 -2367 0 net=3822
rlabel metal2 317 -2367 317 -2367 0 net=2677
rlabel metal2 408 -2367 408 -2367 0 net=4171
rlabel metal2 58 -2369 58 -2369 0 net=6937
rlabel metal2 100 -2369 100 -2369 0 net=7233
rlabel metal2 331 -2369 331 -2369 0 net=3083
rlabel metal2 408 -2369 408 -2369 0 net=3361
rlabel metal2 142 -2371 142 -2371 0 net=6929
rlabel metal2 653 -2371 653 -2371 0 net=7031
rlabel metal2 198 -2373 198 -2373 0 net=1781
rlabel metal2 177 -2375 177 -2375 0 net=1067
rlabel metal2 72 -2386 72 -2386 0 net=7008
rlabel metal2 166 -2386 166 -2386 0 net=1068
rlabel metal2 240 -2386 240 -2386 0 net=4103
rlabel metal2 240 -2386 240 -2386 0 net=4103
rlabel metal2 303 -2386 303 -2386 0 net=3084
rlabel metal2 355 -2386 355 -2386 0 net=5908
rlabel metal2 646 -2386 646 -2386 0 net=4622
rlabel metal2 723 -2386 723 -2386 0 net=6625
rlabel metal2 800 -2386 800 -2386 0 net=6261
rlabel metal2 814 -2386 814 -2386 0 net=6673
rlabel metal2 891 -2386 891 -2386 0 net=7421
rlabel metal2 940 -2386 940 -2386 0 net=5582
rlabel metal2 79 -2388 79 -2388 0 net=6938
rlabel metal2 191 -2388 191 -2388 0 net=1646
rlabel metal2 303 -2388 303 -2388 0 net=3257
rlabel metal2 418 -2388 418 -2388 0 net=807
rlabel metal2 730 -2388 730 -2388 0 net=6347
rlabel metal2 779 -2388 779 -2388 0 net=6293
rlabel metal2 898 -2388 898 -2388 0 net=6127
rlabel metal2 898 -2388 898 -2388 0 net=6127
rlabel metal2 975 -2388 975 -2388 0 net=6008
rlabel metal2 86 -2390 86 -2390 0 net=5454
rlabel metal2 156 -2390 156 -2390 0 net=4584
rlabel metal2 177 -2390 177 -2390 0 net=2374
rlabel metal2 282 -2390 282 -2390 0 net=1869
rlabel metal2 422 -2390 422 -2390 0 net=2368
rlabel metal2 688 -2390 688 -2390 0 net=2514
rlabel metal2 978 -2390 978 -2390 0 net=2316
rlabel metal2 93 -2392 93 -2392 0 net=1844
rlabel metal2 219 -2392 219 -2392 0 net=2207
rlabel metal2 429 -2392 429 -2392 0 net=4902
rlabel metal2 499 -2392 499 -2392 0 net=4173
rlabel metal2 530 -2392 530 -2392 0 net=2112
rlabel metal2 691 -2392 691 -2392 0 net=530
rlabel metal2 121 -2394 121 -2394 0 net=1486
rlabel metal2 310 -2394 310 -2394 0 net=4650
rlabel metal2 394 -2394 394 -2394 0 net=2828
rlabel metal2 516 -2394 516 -2394 0 net=7222
rlabel metal2 135 -2396 135 -2396 0 net=1132
rlabel metal2 453 -2396 453 -2396 0 net=7032
rlabel metal2 142 -2398 142 -2398 0 net=6931
rlabel metal2 205 -2398 205 -2398 0 net=1093
rlabel metal2 247 -2398 247 -2398 0 net=2525
rlabel metal2 268 -2398 268 -2398 0 net=3499
rlabel metal2 310 -2398 310 -2398 0 net=3363
rlabel metal2 443 -2398 443 -2398 0 net=4546
rlabel metal2 576 -2398 576 -2398 0 net=4707
rlabel metal2 653 -2398 653 -2398 0 net=6893
rlabel metal2 261 -2400 261 -2400 0 net=3987
rlabel metal2 345 -2400 345 -2400 0 net=6939
rlabel metal2 436 -2400 436 -2400 0 net=3877
rlabel metal2 450 -2400 450 -2400 0 net=4514
rlabel metal2 499 -2400 499 -2400 0 net=4499
rlabel metal2 516 -2400 516 -2400 0 net=6528
rlabel metal2 674 -2400 674 -2400 0 net=7207
rlabel metal2 254 -2402 254 -2402 0 net=4488
rlabel metal2 352 -2402 352 -2402 0 net=1581
rlabel metal2 548 -2402 548 -2402 0 net=4643
rlabel metal2 716 -2402 716 -2402 0 net=7473
rlabel metal2 128 -2404 128 -2404 0 net=4073
rlabel metal2 296 -2404 296 -2404 0 net=1227
rlabel metal2 415 -2404 415 -2404 0 net=3443
rlabel metal2 492 -2404 492 -2404 0 net=4356
rlabel metal2 513 -2404 513 -2404 0 net=5275
rlabel metal2 709 -2404 709 -2404 0 net=3231
rlabel metal2 212 -2406 212 -2406 0 net=1107
rlabel metal2 359 -2406 359 -2406 0 net=5841
rlabel metal2 436 -2406 436 -2406 0 net=4147
rlabel metal2 460 -2406 460 -2406 0 net=4354
rlabel metal2 492 -2406 492 -2406 0 net=5379
rlabel metal2 548 -2406 548 -2406 0 net=2179
rlabel metal2 576 -2406 576 -2406 0 net=5439
rlabel metal2 289 -2408 289 -2408 0 net=3487
rlabel metal2 366 -2408 366 -2408 0 net=3928
rlabel metal2 100 -2410 100 -2410 0 net=7235
rlabel metal2 369 -2410 369 -2410 0 net=1480
rlabel metal2 478 -2410 478 -2410 0 net=6841
rlabel metal2 555 -2410 555 -2410 0 net=2675
rlabel metal2 114 -2412 114 -2412 0 net=2649
rlabel metal2 523 -2412 523 -2412 0 net=4670
rlabel metal2 597 -2412 597 -2412 0 net=5869
rlabel metal2 611 -2412 611 -2412 0 net=6005
rlabel metal2 331 -2414 331 -2414 0 net=1783
rlabel metal2 604 -2414 604 -2414 0 net=7505
rlabel metal2 233 -2416 233 -2416 0 net=5565
rlabel metal2 373 -2416 373 -2416 0 net=4612
rlabel metal2 632 -2416 632 -2416 0 net=6605
rlabel metal2 667 -2416 667 -2416 0 net=6883
rlabel metal2 226 -2418 226 -2418 0 net=2299
rlabel metal2 338 -2418 338 -2418 0 net=3163
rlabel metal2 471 -2418 471 -2418 0 net=2674
rlabel metal2 618 -2418 618 -2418 0 net=7121
rlabel metal2 681 -2418 681 -2418 0 net=7482
rlabel metal2 107 -2420 107 -2420 0 net=3223
rlabel metal2 317 -2420 317 -2420 0 net=2679
rlabel metal2 471 -2420 471 -2420 0 net=4663
rlabel metal2 618 -2420 618 -2420 0 net=6471
rlabel metal2 758 -2420 758 -2420 0 net=6735
rlabel metal2 275 -2422 275 -2422 0 net=3093
rlabel metal2 562 -2422 562 -2422 0 net=4997
rlabel metal2 737 -2422 737 -2422 0 net=5813
rlabel metal2 275 -2424 275 -2424 0 net=3697
rlabel metal2 520 -2424 520 -2424 0 net=3687
rlabel metal2 737 -2424 737 -2424 0 net=7625
rlabel metal2 282 -2426 282 -2426 0 net=2853
rlabel metal2 429 -2426 429 -2426 0 net=2623
rlabel metal2 772 -2426 772 -2426 0 net=7525
rlabel metal2 226 -2437 226 -2437 0 net=3224
rlabel metal2 380 -2437 380 -2437 0 net=4664
rlabel metal2 509 -2437 509 -2437 0 net=5440
rlabel metal2 607 -2437 607 -2437 0 net=6472
rlabel metal2 639 -2437 639 -2437 0 net=5233
rlabel metal2 702 -2437 702 -2437 0 net=7475
rlabel metal2 723 -2437 723 -2437 0 net=6627
rlabel metal2 723 -2437 723 -2437 0 net=6627
rlabel metal2 744 -2437 744 -2437 0 net=5814
rlabel metal2 807 -2437 807 -2437 0 net=6262
rlabel metal2 828 -2437 828 -2437 0 net=6675
rlabel metal2 828 -2437 828 -2437 0 net=6675
rlabel metal2 898 -2437 898 -2437 0 net=6128
rlabel metal2 219 -2439 219 -2439 0 net=1095
rlabel metal2 233 -2439 233 -2439 0 net=2301
rlabel metal2 261 -2439 261 -2439 0 net=3988
rlabel metal2 387 -2439 387 -2439 0 net=2651
rlabel metal2 569 -2439 569 -2439 0 net=6006
rlabel metal2 614 -2439 614 -2439 0 net=837
rlabel metal2 233 -2441 233 -2441 0 net=2526
rlabel metal2 275 -2441 275 -2441 0 net=3698
rlabel metal2 387 -2441 387 -2441 0 net=2625
rlabel metal2 432 -2441 432 -2441 0 net=4998
rlabel metal2 572 -2441 572 -2441 0 net=5870
rlabel metal2 611 -2441 611 -2441 0 net=6894
rlabel metal2 660 -2441 660 -2441 0 net=7123
rlabel metal2 688 -2441 688 -2441 0 net=7626
rlabel metal2 747 -2441 747 -2441 0 net=6736
rlabel metal2 800 -2441 800 -2441 0 net=6295
rlabel metal2 891 -2441 891 -2441 0 net=7423
rlabel metal2 236 -2443 236 -2443 0 net=548
rlabel metal2 331 -2443 331 -2443 0 net=5566
rlabel metal2 460 -2443 460 -2443 0 net=928
rlabel metal2 240 -2445 240 -2445 0 net=4105
rlabel metal2 240 -2445 240 -2445 0 net=4105
rlabel metal2 282 -2445 282 -2445 0 net=2854
rlabel metal2 450 -2445 450 -2445 0 net=809
rlabel metal2 509 -2445 509 -2445 0 net=5276
rlabel metal2 590 -2445 590 -2445 0 net=3689
rlabel metal2 625 -2445 625 -2445 0 net=4709
rlabel metal2 660 -2445 660 -2445 0 net=7209
rlabel metal2 730 -2445 730 -2445 0 net=6349
rlabel metal2 751 -2445 751 -2445 0 net=3232
rlabel metal2 296 -2447 296 -2447 0 net=1109
rlabel metal2 338 -2447 338 -2447 0 net=2681
rlabel metal2 401 -2447 401 -2447 0 net=1870
rlabel metal2 457 -2447 457 -2447 0 net=5491
rlabel metal2 576 -2447 576 -2447 0 net=7507
rlabel metal2 625 -2447 625 -2447 0 net=6009
rlabel metal2 663 -2447 663 -2447 0 net=1
rlabel metal2 751 -2447 751 -2447 0 net=7526
rlabel metal2 254 -2449 254 -2449 0 net=4075
rlabel metal2 310 -2449 310 -2449 0 net=3365
rlabel metal2 373 -2449 373 -2449 0 net=3165
rlabel metal2 408 -2449 408 -2449 0 net=5843
rlabel metal2 408 -2449 408 -2449 0 net=5843
rlabel metal2 453 -2449 453 -2449 0 net=4500
rlabel metal2 597 -2449 597 -2449 0 net=6607
rlabel metal2 646 -2449 646 -2449 0 net=4645
rlabel metal2 198 -2451 198 -2451 0 net=6932
rlabel metal2 268 -2451 268 -2451 0 net=3501
rlabel metal2 317 -2451 317 -2451 0 net=3094
rlabel metal2 464 -2451 464 -2451 0 net=3445
rlabel metal2 499 -2451 499 -2451 0 net=6843
rlabel metal2 541 -2451 541 -2451 0 net=1583
rlabel metal2 646 -2451 646 -2451 0 net=6884
rlabel metal2 341 -2453 341 -2453 0 net=2180
rlabel metal2 345 -2455 345 -2455 0 net=6941
rlabel metal2 443 -2455 443 -2455 0 net=3879
rlabel metal2 478 -2455 478 -2455 0 net=1785
rlabel metal2 303 -2457 303 -2457 0 net=3258
rlabel metal2 348 -2457 348 -2457 0 net=2676
rlabel metal2 394 -2459 394 -2459 0 net=1228
rlabel metal2 478 -2459 478 -2459 0 net=6677
rlabel metal2 527 -2459 527 -2459 0 net=4175
rlabel metal2 359 -2461 359 -2461 0 net=3489
rlabel metal2 422 -2461 422 -2461 0 net=2209
rlabel metal2 492 -2461 492 -2461 0 net=5381
rlabel metal2 289 -2463 289 -2463 0 net=7237
rlabel metal2 415 -2463 415 -2463 0 net=5505
rlabel metal2 422 -2465 422 -2465 0 net=4149
rlabel metal2 436 -2467 436 -2467 0 net=6695
rlabel metal2 226 -2478 226 -2478 0 net=1097
rlabel metal2 226 -2478 226 -2478 0 net=1097
rlabel metal2 240 -2478 240 -2478 0 net=4107
rlabel metal2 240 -2478 240 -2478 0 net=4107
rlabel metal2 247 -2478 247 -2478 0 net=2302
rlabel metal2 296 -2478 296 -2478 0 net=4076
rlabel metal2 359 -2478 359 -2478 0 net=7239
rlabel metal2 390 -2478 390 -2478 0 net=5492
rlabel metal2 492 -2478 492 -2478 0 net=5506
rlabel metal2 513 -2478 513 -2478 0 net=2652
rlabel metal2 649 -2478 649 -2478 0 net=4710
rlabel metal2 674 -2478 674 -2478 0 net=7124
rlabel metal2 723 -2478 723 -2478 0 net=6628
rlabel metal2 723 -2478 723 -2478 0 net=6628
rlabel metal2 726 -2478 726 -2478 0 net=774
rlabel metal2 310 -2480 310 -2480 0 net=3502
rlabel metal2 359 -2480 359 -2480 0 net=2627
rlabel metal2 394 -2480 394 -2480 0 net=3490
rlabel metal2 432 -2480 432 -2480 0 net=6844
rlabel metal2 527 -2480 527 -2480 0 net=5383
rlabel metal2 541 -2480 541 -2480 0 net=4176
rlabel metal2 604 -2480 604 -2480 0 net=5234
rlabel metal2 653 -2480 653 -2480 0 net=7210
rlabel metal2 688 -2480 688 -2480 0 net=4647
rlabel metal2 744 -2480 744 -2480 0 net=6350
rlabel metal2 807 -2480 807 -2480 0 net=6296
rlabel metal2 828 -2480 828 -2480 0 net=6676
rlabel metal2 898 -2480 898 -2480 0 net=7425
rlabel metal2 331 -2482 331 -2482 0 net=1110
rlabel metal2 373 -2482 373 -2482 0 net=6942
rlabel metal2 401 -2482 401 -2482 0 net=5844
rlabel metal2 443 -2482 443 -2482 0 net=3446
rlabel metal2 548 -2482 548 -2482 0 net=1786
rlabel metal2 632 -2482 632 -2482 0 net=1585
rlabel metal2 688 -2482 688 -2482 0 net=7476
rlabel metal2 352 -2484 352 -2484 0 net=3367
rlabel metal2 404 -2484 404 -2484 0 net=4150
rlabel metal2 446 -2484 446 -2484 0 net=3880
rlabel metal2 485 -2484 485 -2484 0 net=2210
rlabel metal2 551 -2484 551 -2484 0 net=7508
rlabel metal2 597 -2484 597 -2484 0 net=6609
rlabel metal2 614 -2484 614 -2484 0 net=6010
rlabel metal2 366 -2486 366 -2486 0 net=2682
rlabel metal2 453 -2486 453 -2486 0 net=6678
rlabel metal2 618 -2486 618 -2486 0 net=3691
rlabel metal2 366 -2488 366 -2488 0 net=6696
rlabel metal2 226 -2499 226 -2499 0 net=1098
rlabel metal2 236 -2499 236 -2499 0 net=4108
rlabel metal2 359 -2499 359 -2499 0 net=2628
rlabel metal2 373 -2499 373 -2499 0 net=3368
rlabel metal2 397 -2499 397 -2499 0 net=3168
rlabel metal2 534 -2499 534 -2499 0 net=5384
rlabel metal2 558 -2499 558 -2499 0 net=478
rlabel metal2 380 -2501 380 -2501 0 net=7240
rlabel metal2 604 -2501 604 -2501 0 net=6610
rlabel metal2 632 -2501 632 -2501 0 net=3692
rlabel metal2 660 -2501 660 -2501 0 net=1586
rlabel metal2 702 -2501 702 -2501 0 net=4648
rlabel metal2 898 -2501 898 -2501 0 net=7426
<< end >>
