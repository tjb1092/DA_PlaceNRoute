magic
tech scmos
timestamp 1555071770 
<< pdiffusion >>
rect 1 -10 7 -4
rect 8 -10 14 -4
rect 15 -10 21 -4
rect 22 -10 28 -4
rect 29 -10 35 -4
rect 134 -10 137 -4
rect 141 -10 147 -4
rect 148 -10 151 -4
rect 155 -10 161 -4
rect 176 -10 182 -4
rect 1 -27 7 -21
rect 8 -27 14 -21
rect 15 -27 21 -21
rect 22 -27 28 -21
rect 99 -27 105 -21
rect 106 -27 109 -21
rect 120 -27 126 -21
rect 127 -27 133 -21
rect 134 -27 137 -21
rect 141 -27 147 -21
rect 148 -27 154 -21
rect 155 -27 158 -21
rect 162 -27 165 -21
rect 169 -27 172 -21
rect 176 -27 182 -21
rect 183 -27 186 -21
rect 190 -27 196 -21
rect 1 -46 7 -40
rect 8 -46 14 -40
rect 15 -46 21 -40
rect 78 -46 81 -40
rect 85 -46 88 -40
rect 92 -46 95 -40
rect 99 -46 105 -40
rect 106 -46 112 -40
rect 113 -46 119 -40
rect 120 -46 123 -40
rect 127 -46 130 -40
rect 134 -46 137 -40
rect 141 -46 147 -40
rect 148 -46 154 -40
rect 155 -46 161 -40
rect 162 -46 165 -40
rect 169 -46 172 -40
rect 176 -46 182 -40
rect 183 -46 186 -40
rect 190 -46 196 -40
rect 197 -46 200 -40
rect 204 -46 207 -40
rect 211 -46 214 -40
rect 218 -46 221 -40
rect 225 -46 228 -40
rect 1 -71 7 -65
rect 8 -71 14 -65
rect 15 -71 21 -65
rect 78 -71 81 -65
rect 85 -71 88 -65
rect 92 -71 95 -65
rect 99 -71 102 -65
rect 106 -71 112 -65
rect 113 -71 116 -65
rect 120 -71 126 -65
rect 127 -71 133 -65
rect 134 -71 140 -65
rect 141 -71 147 -65
rect 148 -71 154 -65
rect 155 -71 161 -65
rect 162 -71 165 -65
rect 169 -71 172 -65
rect 176 -71 179 -65
rect 183 -71 189 -65
rect 190 -71 193 -65
rect 197 -71 203 -65
rect 204 -71 207 -65
rect 211 -71 214 -65
rect 218 -71 224 -65
rect 225 -71 228 -65
rect 232 -71 235 -65
rect 1 -100 7 -94
rect 8 -100 14 -94
rect 64 -100 67 -94
rect 71 -100 74 -94
rect 78 -100 81 -94
rect 85 -100 91 -94
rect 92 -100 98 -94
rect 99 -100 102 -94
rect 106 -100 112 -94
rect 113 -100 116 -94
rect 120 -100 123 -94
rect 127 -100 133 -94
rect 134 -100 140 -94
rect 141 -100 147 -94
rect 148 -100 154 -94
rect 155 -100 158 -94
rect 162 -100 165 -94
rect 169 -100 175 -94
rect 176 -100 179 -94
rect 183 -100 186 -94
rect 190 -100 193 -94
rect 197 -100 200 -94
rect 204 -100 210 -94
rect 211 -100 214 -94
rect 218 -100 224 -94
rect 225 -100 228 -94
rect 232 -100 235 -94
rect 239 -100 245 -94
rect 246 -100 249 -94
rect 253 -100 256 -94
rect 260 -100 266 -94
rect 267 -100 270 -94
rect 281 -100 284 -94
rect 1 -125 7 -119
rect 29 -125 35 -119
rect 43 -125 49 -119
rect 50 -125 53 -119
rect 57 -125 60 -119
rect 64 -125 67 -119
rect 71 -125 77 -119
rect 78 -125 84 -119
rect 85 -125 88 -119
rect 92 -125 95 -119
rect 99 -125 102 -119
rect 106 -125 109 -119
rect 113 -125 119 -119
rect 120 -125 123 -119
rect 127 -125 133 -119
rect 134 -125 140 -119
rect 141 -125 144 -119
rect 148 -125 151 -119
rect 155 -125 161 -119
rect 162 -125 165 -119
rect 169 -125 172 -119
rect 176 -125 179 -119
rect 183 -125 189 -119
rect 190 -125 196 -119
rect 197 -125 203 -119
rect 204 -125 207 -119
rect 211 -125 214 -119
rect 218 -125 224 -119
rect 225 -125 228 -119
rect 232 -125 235 -119
rect 239 -125 242 -119
rect 246 -125 249 -119
rect 253 -125 256 -119
rect 260 -125 263 -119
rect 267 -125 273 -119
rect 274 -125 277 -119
rect 281 -125 284 -119
rect 288 -125 291 -119
rect 295 -125 301 -119
rect 302 -125 305 -119
rect 323 -125 329 -119
rect 15 -154 21 -148
rect 22 -154 25 -148
rect 29 -154 35 -148
rect 36 -154 39 -148
rect 43 -154 49 -148
rect 50 -154 56 -148
rect 57 -154 60 -148
rect 64 -154 70 -148
rect 71 -154 77 -148
rect 78 -154 81 -148
rect 85 -154 88 -148
rect 92 -154 98 -148
rect 99 -154 102 -148
rect 106 -154 109 -148
rect 113 -154 119 -148
rect 120 -154 123 -148
rect 127 -154 133 -148
rect 134 -154 137 -148
rect 141 -154 144 -148
rect 148 -154 154 -148
rect 155 -154 158 -148
rect 162 -154 168 -148
rect 169 -154 175 -148
rect 176 -154 182 -148
rect 183 -154 186 -148
rect 190 -154 193 -148
rect 197 -154 203 -148
rect 204 -154 207 -148
rect 211 -154 217 -148
rect 218 -154 224 -148
rect 225 -154 228 -148
rect 232 -154 238 -148
rect 239 -154 242 -148
rect 246 -154 249 -148
rect 253 -154 256 -148
rect 260 -154 263 -148
rect 267 -154 270 -148
rect 274 -154 277 -148
rect 281 -154 284 -148
rect 288 -154 291 -148
rect 295 -154 298 -148
rect 302 -154 305 -148
rect 309 -154 312 -148
rect 316 -154 319 -148
rect 323 -154 326 -148
rect 330 -154 336 -148
rect 337 -154 343 -148
rect 344 -154 347 -148
rect 15 -193 21 -187
rect 43 -193 46 -187
rect 50 -193 53 -187
rect 57 -193 63 -187
rect 64 -193 70 -187
rect 71 -193 74 -187
rect 78 -193 81 -187
rect 85 -193 88 -187
rect 92 -193 95 -187
rect 99 -193 102 -187
rect 106 -193 109 -187
rect 113 -193 119 -187
rect 120 -193 126 -187
rect 127 -193 130 -187
rect 134 -193 137 -187
rect 141 -193 147 -187
rect 148 -193 151 -187
rect 155 -193 161 -187
rect 162 -193 165 -187
rect 169 -193 175 -187
rect 176 -193 182 -187
rect 183 -193 189 -187
rect 190 -193 193 -187
rect 197 -193 200 -187
rect 204 -193 210 -187
rect 211 -193 217 -187
rect 218 -193 221 -187
rect 225 -193 231 -187
rect 232 -193 235 -187
rect 239 -193 245 -187
rect 246 -193 249 -187
rect 253 -193 256 -187
rect 260 -193 263 -187
rect 267 -193 270 -187
rect 274 -193 277 -187
rect 281 -193 284 -187
rect 288 -193 291 -187
rect 295 -193 301 -187
rect 302 -193 308 -187
rect 309 -193 312 -187
rect 316 -193 322 -187
rect 323 -193 326 -187
rect 351 -193 357 -187
rect 358 -193 364 -187
rect 29 -224 32 -218
rect 36 -224 42 -218
rect 43 -224 46 -218
rect 50 -224 56 -218
rect 57 -224 60 -218
rect 64 -224 67 -218
rect 71 -224 74 -218
rect 78 -224 84 -218
rect 85 -224 91 -218
rect 92 -224 95 -218
rect 99 -224 105 -218
rect 106 -224 112 -218
rect 113 -224 116 -218
rect 120 -224 123 -218
rect 127 -224 130 -218
rect 134 -224 140 -218
rect 141 -224 144 -218
rect 148 -224 154 -218
rect 155 -224 161 -218
rect 162 -224 165 -218
rect 169 -224 172 -218
rect 176 -224 179 -218
rect 183 -224 189 -218
rect 190 -224 193 -218
rect 197 -224 200 -218
rect 204 -224 207 -218
rect 211 -224 217 -218
rect 218 -224 221 -218
rect 225 -224 228 -218
rect 232 -224 238 -218
rect 239 -224 242 -218
rect 246 -224 252 -218
rect 253 -224 256 -218
rect 260 -224 263 -218
rect 267 -224 270 -218
rect 274 -224 277 -218
rect 281 -224 284 -218
rect 288 -224 291 -218
rect 295 -224 298 -218
rect 302 -224 305 -218
rect 309 -224 312 -218
rect 316 -224 322 -218
rect 323 -224 329 -218
rect 330 -224 336 -218
rect 337 -224 343 -218
rect 344 -224 347 -218
rect 351 -224 357 -218
rect 358 -224 361 -218
rect 365 -224 368 -218
rect 372 -224 378 -218
rect 379 -224 382 -218
rect 386 -224 392 -218
rect 8 -253 11 -247
rect 15 -253 18 -247
rect 22 -253 25 -247
rect 29 -253 35 -247
rect 36 -253 42 -247
rect 43 -253 46 -247
rect 50 -253 56 -247
rect 57 -253 60 -247
rect 64 -253 67 -247
rect 71 -253 74 -247
rect 78 -253 84 -247
rect 85 -253 91 -247
rect 92 -253 95 -247
rect 99 -253 102 -247
rect 106 -253 112 -247
rect 113 -253 119 -247
rect 120 -253 123 -247
rect 127 -253 133 -247
rect 134 -253 137 -247
rect 141 -253 147 -247
rect 148 -253 154 -247
rect 155 -253 158 -247
rect 162 -253 165 -247
rect 169 -253 175 -247
rect 176 -253 179 -247
rect 183 -253 186 -247
rect 190 -253 193 -247
rect 197 -253 200 -247
rect 204 -253 210 -247
rect 211 -253 214 -247
rect 218 -253 224 -247
rect 225 -253 228 -247
rect 232 -253 235 -247
rect 239 -253 242 -247
rect 246 -253 249 -247
rect 253 -253 256 -247
rect 260 -253 263 -247
rect 267 -253 273 -247
rect 274 -253 277 -247
rect 281 -253 284 -247
rect 288 -253 291 -247
rect 295 -253 298 -247
rect 302 -253 305 -247
rect 309 -253 312 -247
rect 316 -253 319 -247
rect 323 -253 329 -247
rect 330 -253 333 -247
rect 337 -253 343 -247
rect 344 -253 350 -247
rect 351 -253 354 -247
rect 379 -253 385 -247
rect 386 -253 392 -247
rect 393 -253 396 -247
rect 1 -300 4 -294
rect 8 -300 14 -294
rect 15 -300 18 -294
rect 22 -300 25 -294
rect 29 -300 35 -294
rect 36 -300 39 -294
rect 43 -300 46 -294
rect 50 -300 56 -294
rect 57 -300 60 -294
rect 64 -300 70 -294
rect 71 -300 77 -294
rect 78 -300 84 -294
rect 85 -300 88 -294
rect 92 -300 98 -294
rect 99 -300 102 -294
rect 106 -300 109 -294
rect 113 -300 119 -294
rect 120 -300 123 -294
rect 127 -300 133 -294
rect 134 -300 137 -294
rect 141 -300 144 -294
rect 148 -300 154 -294
rect 155 -300 161 -294
rect 162 -300 165 -294
rect 169 -300 175 -294
rect 176 -300 182 -294
rect 183 -300 189 -294
rect 190 -300 196 -294
rect 197 -300 200 -294
rect 204 -300 210 -294
rect 211 -300 217 -294
rect 218 -300 221 -294
rect 225 -300 228 -294
rect 232 -300 238 -294
rect 239 -300 245 -294
rect 246 -300 249 -294
rect 253 -300 256 -294
rect 260 -300 263 -294
rect 267 -300 270 -294
rect 274 -300 277 -294
rect 281 -300 284 -294
rect 288 -300 291 -294
rect 295 -300 298 -294
rect 302 -300 305 -294
rect 309 -300 312 -294
rect 316 -300 319 -294
rect 323 -300 326 -294
rect 330 -300 333 -294
rect 337 -300 340 -294
rect 344 -300 347 -294
rect 29 -347 32 -341
rect 36 -347 39 -341
rect 43 -347 46 -341
rect 50 -347 56 -341
rect 57 -347 60 -341
rect 64 -347 67 -341
rect 71 -347 77 -341
rect 78 -347 81 -341
rect 85 -347 88 -341
rect 92 -347 95 -341
rect 99 -347 105 -341
rect 106 -347 112 -341
rect 113 -347 119 -341
rect 120 -347 126 -341
rect 127 -347 130 -341
rect 134 -347 140 -341
rect 141 -347 147 -341
rect 148 -347 154 -341
rect 155 -347 161 -341
rect 162 -347 165 -341
rect 169 -347 172 -341
rect 176 -347 179 -341
rect 183 -347 189 -341
rect 190 -347 196 -341
rect 197 -347 203 -341
rect 204 -347 210 -341
rect 211 -347 217 -341
rect 218 -347 221 -341
rect 225 -347 231 -341
rect 232 -347 235 -341
rect 239 -347 245 -341
rect 246 -347 249 -341
rect 253 -347 256 -341
rect 260 -347 263 -341
rect 267 -347 270 -341
rect 274 -347 277 -341
rect 281 -347 284 -341
rect 288 -347 291 -341
rect 295 -347 301 -341
rect 302 -347 305 -341
rect 309 -347 312 -341
rect 316 -347 319 -341
rect 323 -347 326 -341
rect 1 -382 4 -376
rect 8 -382 11 -376
rect 15 -382 18 -376
rect 22 -382 25 -376
rect 29 -382 35 -376
rect 36 -382 39 -376
rect 43 -382 46 -376
rect 50 -382 53 -376
rect 57 -382 63 -376
rect 64 -382 70 -376
rect 71 -382 77 -376
rect 78 -382 81 -376
rect 85 -382 91 -376
rect 92 -382 98 -376
rect 99 -382 102 -376
rect 106 -382 109 -376
rect 113 -382 119 -376
rect 120 -382 123 -376
rect 127 -382 130 -376
rect 134 -382 140 -376
rect 141 -382 147 -376
rect 148 -382 151 -376
rect 155 -382 161 -376
rect 162 -382 168 -376
rect 169 -382 175 -376
rect 176 -382 182 -376
rect 183 -382 189 -376
rect 190 -382 196 -376
rect 197 -382 200 -376
rect 204 -382 207 -376
rect 211 -382 217 -376
rect 218 -382 221 -376
rect 225 -382 228 -376
rect 232 -382 235 -376
rect 239 -382 242 -376
rect 246 -382 249 -376
rect 253 -382 256 -376
rect 260 -382 266 -376
rect 267 -382 270 -376
rect 274 -382 277 -376
rect 281 -382 284 -376
rect 288 -382 291 -376
rect 295 -382 298 -376
rect 302 -382 308 -376
rect 309 -382 312 -376
rect 316 -382 319 -376
rect 323 -382 326 -376
rect 330 -382 333 -376
rect 337 -382 340 -376
rect 344 -382 347 -376
rect 22 -423 25 -417
rect 29 -423 32 -417
rect 36 -423 42 -417
rect 43 -423 46 -417
rect 50 -423 56 -417
rect 57 -423 60 -417
rect 64 -423 67 -417
rect 71 -423 77 -417
rect 78 -423 84 -417
rect 85 -423 88 -417
rect 92 -423 98 -417
rect 99 -423 105 -417
rect 106 -423 112 -417
rect 127 -423 130 -417
rect 134 -423 137 -417
rect 141 -423 144 -417
rect 148 -423 154 -417
rect 155 -423 158 -417
rect 162 -423 165 -417
rect 169 -423 175 -417
rect 176 -423 179 -417
rect 183 -423 186 -417
rect 190 -423 193 -417
rect 197 -423 203 -417
rect 204 -423 207 -417
rect 211 -423 217 -417
rect 218 -423 224 -417
rect 225 -423 231 -417
rect 232 -423 235 -417
rect 239 -423 245 -417
rect 246 -423 249 -417
rect 253 -423 256 -417
rect 260 -423 263 -417
rect 267 -423 273 -417
rect 274 -423 277 -417
rect 281 -423 287 -417
rect 288 -423 294 -417
rect 295 -423 298 -417
rect 302 -423 305 -417
rect 309 -423 312 -417
rect 316 -423 319 -417
rect 1 -454 4 -448
rect 8 -454 11 -448
rect 15 -454 18 -448
rect 22 -454 25 -448
rect 29 -454 32 -448
rect 36 -454 39 -448
rect 43 -454 49 -448
rect 50 -454 53 -448
rect 57 -454 63 -448
rect 64 -454 67 -448
rect 71 -454 77 -448
rect 78 -454 84 -448
rect 85 -454 91 -448
rect 92 -454 95 -448
rect 99 -454 105 -448
rect 106 -454 112 -448
rect 113 -454 116 -448
rect 120 -454 123 -448
rect 127 -454 133 -448
rect 134 -454 140 -448
rect 141 -454 144 -448
rect 148 -454 151 -448
rect 155 -454 161 -448
rect 162 -454 165 -448
rect 169 -454 175 -448
rect 176 -454 179 -448
rect 183 -454 186 -448
rect 190 -454 196 -448
rect 197 -454 203 -448
rect 204 -454 207 -448
rect 211 -454 217 -448
rect 218 -454 224 -448
rect 225 -454 228 -448
rect 232 -454 238 -448
rect 239 -454 242 -448
rect 246 -454 249 -448
rect 253 -454 256 -448
rect 260 -454 263 -448
rect 267 -454 270 -448
rect 274 -454 277 -448
rect 281 -454 284 -448
rect 288 -454 291 -448
rect 295 -454 298 -448
rect 302 -454 305 -448
rect 309 -454 312 -448
rect 316 -454 319 -448
rect 323 -454 329 -448
rect 330 -454 336 -448
rect 337 -454 340 -448
rect 36 -495 42 -489
rect 43 -495 46 -489
rect 50 -495 53 -489
rect 57 -495 60 -489
rect 64 -495 67 -489
rect 71 -495 77 -489
rect 78 -495 84 -489
rect 85 -495 88 -489
rect 92 -495 95 -489
rect 99 -495 102 -489
rect 106 -495 109 -489
rect 113 -495 116 -489
rect 120 -495 126 -489
rect 127 -495 133 -489
rect 134 -495 140 -489
rect 141 -495 147 -489
rect 148 -495 151 -489
rect 155 -495 158 -489
rect 162 -495 165 -489
rect 169 -495 172 -489
rect 176 -495 182 -489
rect 183 -495 186 -489
rect 190 -495 193 -489
rect 197 -495 203 -489
rect 204 -495 207 -489
rect 211 -495 217 -489
rect 218 -495 224 -489
rect 225 -495 228 -489
rect 232 -495 235 -489
rect 239 -495 242 -489
rect 246 -495 249 -489
rect 253 -495 259 -489
rect 260 -495 263 -489
rect 267 -495 270 -489
rect 274 -495 277 -489
rect 281 -495 287 -489
rect 288 -495 291 -489
rect 295 -495 298 -489
rect 302 -495 305 -489
rect 309 -495 312 -489
rect 316 -495 322 -489
rect 323 -495 329 -489
rect 330 -495 333 -489
rect 337 -495 340 -489
rect 344 -495 350 -489
rect 351 -495 354 -489
rect 358 -495 361 -489
rect 365 -495 371 -489
rect 15 -532 18 -526
rect 22 -532 25 -526
rect 29 -532 32 -526
rect 36 -532 42 -526
rect 43 -532 49 -526
rect 50 -532 53 -526
rect 57 -532 63 -526
rect 64 -532 67 -526
rect 71 -532 74 -526
rect 78 -532 84 -526
rect 85 -532 88 -526
rect 92 -532 95 -526
rect 99 -532 105 -526
rect 106 -532 109 -526
rect 113 -532 116 -526
rect 120 -532 126 -526
rect 127 -532 130 -526
rect 134 -532 140 -526
rect 141 -532 144 -526
rect 148 -532 151 -526
rect 155 -532 161 -526
rect 162 -532 168 -526
rect 169 -532 172 -526
rect 176 -532 182 -526
rect 183 -532 186 -526
rect 190 -532 196 -526
rect 197 -532 203 -526
rect 204 -532 210 -526
rect 211 -532 217 -526
rect 218 -532 221 -526
rect 225 -532 231 -526
rect 232 -532 235 -526
rect 239 -532 242 -526
rect 246 -532 249 -526
rect 253 -532 256 -526
rect 260 -532 263 -526
rect 267 -532 273 -526
rect 274 -532 277 -526
rect 281 -532 284 -526
rect 288 -532 291 -526
rect 295 -532 298 -526
rect 302 -532 305 -526
rect 309 -532 312 -526
rect 316 -532 319 -526
rect 323 -532 326 -526
rect 330 -532 336 -526
rect 337 -532 340 -526
rect 344 -532 347 -526
rect 351 -532 354 -526
rect 8 -575 11 -569
rect 15 -575 18 -569
rect 22 -575 25 -569
rect 29 -575 35 -569
rect 36 -575 42 -569
rect 43 -575 49 -569
rect 50 -575 53 -569
rect 57 -575 63 -569
rect 64 -575 70 -569
rect 71 -575 74 -569
rect 78 -575 84 -569
rect 85 -575 88 -569
rect 92 -575 95 -569
rect 99 -575 102 -569
rect 106 -575 112 -569
rect 113 -575 119 -569
rect 120 -575 123 -569
rect 127 -575 130 -569
rect 134 -575 140 -569
rect 141 -575 144 -569
rect 148 -575 154 -569
rect 155 -575 158 -569
rect 162 -575 168 -569
rect 169 -575 172 -569
rect 176 -575 182 -569
rect 183 -575 186 -569
rect 190 -575 193 -569
rect 197 -575 200 -569
rect 204 -575 207 -569
rect 211 -575 214 -569
rect 218 -575 224 -569
rect 225 -575 228 -569
rect 232 -575 238 -569
rect 239 -575 245 -569
rect 246 -575 252 -569
rect 253 -575 256 -569
rect 260 -575 263 -569
rect 267 -575 270 -569
rect 274 -575 277 -569
rect 281 -575 284 -569
rect 288 -575 291 -569
rect 295 -575 298 -569
rect 302 -575 305 -569
rect 309 -575 312 -569
rect 316 -575 319 -569
rect 323 -575 326 -569
rect 330 -575 333 -569
rect 337 -575 340 -569
rect 344 -575 347 -569
rect 351 -575 354 -569
rect 358 -575 364 -569
rect 365 -575 371 -569
rect 43 -612 49 -606
rect 50 -612 53 -606
rect 64 -612 70 -606
rect 71 -612 74 -606
rect 78 -612 84 -606
rect 85 -612 88 -606
rect 92 -612 95 -606
rect 99 -612 105 -606
rect 106 -612 112 -606
rect 113 -612 116 -606
rect 120 -612 126 -606
rect 127 -612 130 -606
rect 134 -612 137 -606
rect 141 -612 147 -606
rect 148 -612 154 -606
rect 155 -612 158 -606
rect 162 -612 168 -606
rect 169 -612 172 -606
rect 176 -612 179 -606
rect 183 -612 189 -606
rect 190 -612 196 -606
rect 197 -612 200 -606
rect 204 -612 207 -606
rect 211 -612 217 -606
rect 218 -612 221 -606
rect 225 -612 231 -606
rect 232 -612 235 -606
rect 239 -612 242 -606
rect 246 -612 252 -606
rect 253 -612 259 -606
rect 260 -612 266 -606
rect 267 -612 270 -606
rect 274 -612 280 -606
rect 281 -612 284 -606
rect 288 -612 294 -606
rect 309 -612 312 -606
rect 43 -643 49 -637
rect 50 -643 53 -637
rect 57 -643 60 -637
rect 64 -643 70 -637
rect 71 -643 74 -637
rect 78 -643 84 -637
rect 85 -643 88 -637
rect 92 -643 98 -637
rect 99 -643 105 -637
rect 106 -643 109 -637
rect 113 -643 116 -637
rect 120 -643 126 -637
rect 127 -643 130 -637
rect 134 -643 140 -637
rect 141 -643 147 -637
rect 148 -643 154 -637
rect 155 -643 158 -637
rect 162 -643 165 -637
rect 169 -643 175 -637
rect 176 -643 182 -637
rect 183 -643 186 -637
rect 190 -643 196 -637
rect 197 -643 200 -637
rect 204 -643 210 -637
rect 211 -643 214 -637
rect 218 -643 221 -637
rect 225 -643 228 -637
rect 232 -643 235 -637
rect 239 -643 242 -637
rect 246 -643 249 -637
rect 253 -643 256 -637
rect 260 -643 263 -637
rect 267 -643 270 -637
rect 274 -643 277 -637
rect 281 -643 284 -637
rect 288 -643 294 -637
rect 295 -643 301 -637
rect 302 -643 305 -637
rect 309 -643 315 -637
rect 43 -670 46 -664
rect 50 -670 56 -664
rect 57 -670 63 -664
rect 64 -670 67 -664
rect 71 -670 74 -664
rect 78 -670 81 -664
rect 85 -670 91 -664
rect 92 -670 98 -664
rect 99 -670 105 -664
rect 106 -670 109 -664
rect 113 -670 116 -664
rect 120 -670 126 -664
rect 134 -670 140 -664
rect 141 -670 147 -664
rect 148 -670 151 -664
rect 169 -670 172 -664
rect 176 -670 182 -664
rect 183 -670 186 -664
rect 190 -670 193 -664
rect 197 -670 203 -664
rect 204 -670 207 -664
rect 211 -670 217 -664
rect 218 -670 224 -664
rect 225 -670 228 -664
rect 232 -670 235 -664
rect 239 -670 245 -664
rect 253 -670 256 -664
rect 260 -670 266 -664
rect 267 -670 270 -664
rect 274 -670 280 -664
rect 281 -670 287 -664
rect 288 -670 294 -664
rect 43 -685 49 -679
rect 50 -685 53 -679
rect 57 -685 60 -679
rect 64 -685 70 -679
rect 71 -685 77 -679
rect 78 -685 81 -679
rect 85 -685 91 -679
rect 92 -685 98 -679
rect 99 -685 105 -679
rect 106 -685 112 -679
rect 113 -685 119 -679
rect 120 -685 123 -679
rect 127 -685 130 -679
rect 134 -685 137 -679
rect 141 -685 147 -679
rect 148 -685 154 -679
rect 190 -685 196 -679
rect 197 -685 203 -679
rect 204 -685 207 -679
rect 211 -685 214 -679
rect 218 -685 224 -679
rect 225 -685 228 -679
rect 232 -685 238 -679
rect 239 -685 245 -679
rect 246 -685 249 -679
rect 253 -685 256 -679
rect 260 -685 266 -679
rect 274 -685 277 -679
rect 281 -685 287 -679
<< polysilicon >>
rect 135 -5 136 -3
rect 135 -11 136 -9
rect 142 -5 143 -3
rect 145 -5 146 -3
rect 149 -5 150 -3
rect 149 -11 150 -9
rect 159 -11 160 -9
rect 177 -11 178 -9
rect 100 -22 101 -20
rect 107 -22 108 -20
rect 107 -28 108 -26
rect 121 -22 122 -20
rect 128 -22 129 -20
rect 135 -22 136 -20
rect 135 -28 136 -26
rect 142 -22 143 -20
rect 145 -22 146 -20
rect 142 -28 143 -26
rect 152 -22 153 -20
rect 152 -28 153 -26
rect 156 -22 157 -20
rect 156 -28 157 -26
rect 163 -22 164 -20
rect 163 -28 164 -26
rect 170 -22 171 -20
rect 170 -28 171 -26
rect 177 -22 178 -20
rect 180 -22 181 -20
rect 184 -22 185 -20
rect 184 -28 185 -26
rect 191 -28 192 -26
rect 79 -41 80 -39
rect 79 -47 80 -45
rect 86 -41 87 -39
rect 86 -47 87 -45
rect 93 -41 94 -39
rect 93 -47 94 -45
rect 100 -41 101 -39
rect 103 -41 104 -39
rect 107 -47 108 -45
rect 110 -47 111 -45
rect 117 -41 118 -39
rect 114 -47 115 -45
rect 121 -41 122 -39
rect 121 -47 122 -45
rect 128 -41 129 -39
rect 128 -47 129 -45
rect 135 -41 136 -39
rect 135 -47 136 -45
rect 142 -41 143 -39
rect 142 -47 143 -45
rect 145 -47 146 -45
rect 149 -41 150 -39
rect 152 -41 153 -39
rect 149 -47 150 -45
rect 159 -41 160 -39
rect 156 -47 157 -45
rect 163 -41 164 -39
rect 163 -47 164 -45
rect 170 -41 171 -39
rect 170 -47 171 -45
rect 180 -41 181 -39
rect 180 -47 181 -45
rect 184 -41 185 -39
rect 184 -47 185 -45
rect 194 -41 195 -39
rect 191 -47 192 -45
rect 198 -41 199 -39
rect 198 -47 199 -45
rect 205 -41 206 -39
rect 205 -47 206 -45
rect 212 -41 213 -39
rect 212 -47 213 -45
rect 219 -41 220 -39
rect 219 -47 220 -45
rect 226 -41 227 -39
rect 226 -47 227 -45
rect 79 -66 80 -64
rect 79 -72 80 -70
rect 86 -66 87 -64
rect 86 -72 87 -70
rect 93 -66 94 -64
rect 93 -72 94 -70
rect 100 -66 101 -64
rect 100 -72 101 -70
rect 110 -66 111 -64
rect 107 -72 108 -70
rect 114 -66 115 -64
rect 114 -72 115 -70
rect 121 -72 122 -70
rect 124 -72 125 -70
rect 131 -66 132 -64
rect 131 -72 132 -70
rect 138 -66 139 -64
rect 135 -72 136 -70
rect 138 -72 139 -70
rect 142 -66 143 -64
rect 145 -66 146 -64
rect 142 -72 143 -70
rect 149 -66 150 -64
rect 152 -66 153 -64
rect 156 -66 157 -64
rect 156 -72 157 -70
rect 159 -72 160 -70
rect 163 -66 164 -64
rect 163 -72 164 -70
rect 170 -66 171 -64
rect 170 -72 171 -70
rect 177 -66 178 -64
rect 177 -72 178 -70
rect 187 -66 188 -64
rect 191 -66 192 -64
rect 191 -72 192 -70
rect 198 -72 199 -70
rect 205 -66 206 -64
rect 205 -72 206 -70
rect 212 -66 213 -64
rect 212 -72 213 -70
rect 222 -66 223 -64
rect 226 -66 227 -64
rect 226 -72 227 -70
rect 233 -66 234 -64
rect 233 -72 234 -70
rect 65 -95 66 -93
rect 65 -101 66 -99
rect 72 -95 73 -93
rect 72 -101 73 -99
rect 79 -95 80 -93
rect 79 -101 80 -99
rect 86 -95 87 -93
rect 93 -95 94 -93
rect 93 -101 94 -99
rect 100 -95 101 -93
rect 100 -101 101 -99
rect 107 -95 108 -93
rect 107 -101 108 -99
rect 114 -95 115 -93
rect 114 -101 115 -99
rect 121 -95 122 -93
rect 121 -101 122 -99
rect 128 -95 129 -93
rect 131 -101 132 -99
rect 138 -95 139 -93
rect 135 -101 136 -99
rect 142 -95 143 -93
rect 142 -101 143 -99
rect 152 -95 153 -93
rect 149 -101 150 -99
rect 152 -101 153 -99
rect 156 -95 157 -93
rect 156 -101 157 -99
rect 163 -95 164 -93
rect 163 -101 164 -99
rect 170 -95 171 -93
rect 173 -101 174 -99
rect 177 -95 178 -93
rect 177 -101 178 -99
rect 184 -95 185 -93
rect 184 -101 185 -99
rect 191 -95 192 -93
rect 191 -101 192 -99
rect 198 -95 199 -93
rect 198 -101 199 -99
rect 205 -95 206 -93
rect 205 -101 206 -99
rect 212 -95 213 -93
rect 212 -101 213 -99
rect 219 -95 220 -93
rect 222 -95 223 -93
rect 219 -101 220 -99
rect 226 -95 227 -93
rect 226 -101 227 -99
rect 233 -95 234 -93
rect 233 -101 234 -99
rect 240 -95 241 -93
rect 243 -95 244 -93
rect 243 -101 244 -99
rect 247 -95 248 -93
rect 247 -101 248 -99
rect 254 -95 255 -93
rect 254 -101 255 -99
rect 261 -95 262 -93
rect 264 -101 265 -99
rect 268 -95 269 -93
rect 268 -101 269 -99
rect 282 -95 283 -93
rect 282 -101 283 -99
rect 33 -126 34 -124
rect 44 -120 45 -118
rect 51 -120 52 -118
rect 51 -126 52 -124
rect 58 -120 59 -118
rect 58 -126 59 -124
rect 65 -120 66 -118
rect 65 -126 66 -124
rect 75 -120 76 -118
rect 79 -126 80 -124
rect 82 -126 83 -124
rect 86 -120 87 -118
rect 86 -126 87 -124
rect 93 -120 94 -118
rect 93 -126 94 -124
rect 100 -120 101 -118
rect 100 -126 101 -124
rect 107 -120 108 -118
rect 107 -126 108 -124
rect 114 -120 115 -118
rect 117 -120 118 -118
rect 114 -126 115 -124
rect 121 -120 122 -118
rect 121 -126 122 -124
rect 128 -120 129 -118
rect 128 -126 129 -124
rect 131 -126 132 -124
rect 138 -120 139 -118
rect 142 -120 143 -118
rect 142 -126 143 -124
rect 149 -120 150 -118
rect 149 -126 150 -124
rect 156 -120 157 -118
rect 159 -120 160 -118
rect 156 -126 157 -124
rect 159 -126 160 -124
rect 163 -120 164 -118
rect 163 -126 164 -124
rect 170 -120 171 -118
rect 170 -126 171 -124
rect 177 -120 178 -118
rect 177 -126 178 -124
rect 184 -120 185 -118
rect 184 -126 185 -124
rect 191 -126 192 -124
rect 194 -126 195 -124
rect 201 -120 202 -118
rect 198 -126 199 -124
rect 205 -120 206 -118
rect 205 -126 206 -124
rect 212 -120 213 -118
rect 212 -126 213 -124
rect 219 -120 220 -118
rect 222 -120 223 -118
rect 226 -120 227 -118
rect 226 -126 227 -124
rect 233 -120 234 -118
rect 233 -126 234 -124
rect 240 -120 241 -118
rect 240 -126 241 -124
rect 247 -120 248 -118
rect 247 -126 248 -124
rect 254 -120 255 -118
rect 254 -126 255 -124
rect 261 -120 262 -118
rect 261 -126 262 -124
rect 271 -126 272 -124
rect 275 -120 276 -118
rect 275 -126 276 -124
rect 282 -120 283 -118
rect 282 -126 283 -124
rect 289 -120 290 -118
rect 289 -126 290 -124
rect 296 -120 297 -118
rect 299 -120 300 -118
rect 299 -126 300 -124
rect 303 -120 304 -118
rect 303 -126 304 -124
rect 324 -126 325 -124
rect 19 -149 20 -147
rect 23 -149 24 -147
rect 23 -155 24 -153
rect 30 -149 31 -147
rect 37 -149 38 -147
rect 37 -155 38 -153
rect 47 -149 48 -147
rect 51 -155 52 -153
rect 58 -149 59 -147
rect 58 -155 59 -153
rect 65 -149 66 -147
rect 68 -149 69 -147
rect 68 -155 69 -153
rect 72 -149 73 -147
rect 79 -149 80 -147
rect 79 -155 80 -153
rect 86 -149 87 -147
rect 86 -155 87 -153
rect 93 -149 94 -147
rect 96 -149 97 -147
rect 93 -155 94 -153
rect 100 -149 101 -147
rect 100 -155 101 -153
rect 107 -149 108 -147
rect 107 -155 108 -153
rect 114 -149 115 -147
rect 114 -155 115 -153
rect 121 -149 122 -147
rect 121 -155 122 -153
rect 128 -155 129 -153
rect 135 -149 136 -147
rect 135 -155 136 -153
rect 142 -149 143 -147
rect 142 -155 143 -153
rect 149 -149 150 -147
rect 152 -149 153 -147
rect 149 -155 150 -153
rect 152 -155 153 -153
rect 156 -149 157 -147
rect 156 -155 157 -153
rect 163 -149 164 -147
rect 166 -149 167 -147
rect 163 -155 164 -153
rect 166 -155 167 -153
rect 170 -149 171 -147
rect 173 -149 174 -147
rect 173 -155 174 -153
rect 177 -149 178 -147
rect 180 -155 181 -153
rect 184 -149 185 -147
rect 184 -155 185 -153
rect 191 -149 192 -147
rect 191 -155 192 -153
rect 201 -149 202 -147
rect 198 -155 199 -153
rect 201 -155 202 -153
rect 205 -149 206 -147
rect 205 -155 206 -153
rect 212 -155 213 -153
rect 215 -155 216 -153
rect 219 -149 220 -147
rect 226 -149 227 -147
rect 226 -155 227 -153
rect 236 -149 237 -147
rect 233 -155 234 -153
rect 240 -149 241 -147
rect 240 -155 241 -153
rect 247 -149 248 -147
rect 247 -155 248 -153
rect 254 -149 255 -147
rect 254 -155 255 -153
rect 261 -149 262 -147
rect 261 -155 262 -153
rect 268 -149 269 -147
rect 268 -155 269 -153
rect 275 -149 276 -147
rect 275 -155 276 -153
rect 282 -149 283 -147
rect 282 -155 283 -153
rect 289 -149 290 -147
rect 289 -155 290 -153
rect 296 -149 297 -147
rect 296 -155 297 -153
rect 303 -149 304 -147
rect 303 -155 304 -153
rect 310 -149 311 -147
rect 310 -155 311 -153
rect 317 -149 318 -147
rect 317 -155 318 -153
rect 324 -149 325 -147
rect 324 -155 325 -153
rect 331 -149 332 -147
rect 334 -155 335 -153
rect 341 -149 342 -147
rect 345 -149 346 -147
rect 345 -155 346 -153
rect 19 -188 20 -186
rect 44 -188 45 -186
rect 44 -194 45 -192
rect 51 -188 52 -186
rect 51 -194 52 -192
rect 58 -188 59 -186
rect 61 -188 62 -186
rect 61 -194 62 -192
rect 68 -194 69 -192
rect 72 -188 73 -186
rect 72 -194 73 -192
rect 79 -188 80 -186
rect 79 -194 80 -192
rect 86 -188 87 -186
rect 86 -194 87 -192
rect 93 -188 94 -186
rect 93 -194 94 -192
rect 100 -188 101 -186
rect 100 -194 101 -192
rect 107 -188 108 -186
rect 107 -194 108 -192
rect 114 -188 115 -186
rect 117 -188 118 -186
rect 114 -194 115 -192
rect 117 -194 118 -192
rect 121 -188 122 -186
rect 124 -188 125 -186
rect 128 -188 129 -186
rect 128 -194 129 -192
rect 135 -188 136 -186
rect 135 -194 136 -192
rect 142 -194 143 -192
rect 145 -194 146 -192
rect 149 -188 150 -186
rect 149 -194 150 -192
rect 159 -188 160 -186
rect 159 -194 160 -192
rect 163 -188 164 -186
rect 163 -194 164 -192
rect 173 -188 174 -186
rect 177 -188 178 -186
rect 180 -188 181 -186
rect 180 -194 181 -192
rect 184 -188 185 -186
rect 191 -188 192 -186
rect 191 -194 192 -192
rect 198 -188 199 -186
rect 198 -194 199 -192
rect 205 -188 206 -186
rect 208 -194 209 -192
rect 212 -188 213 -186
rect 215 -194 216 -192
rect 219 -188 220 -186
rect 219 -194 220 -192
rect 226 -188 227 -186
rect 226 -194 227 -192
rect 229 -194 230 -192
rect 233 -188 234 -186
rect 233 -194 234 -192
rect 240 -194 241 -192
rect 243 -194 244 -192
rect 247 -188 248 -186
rect 247 -194 248 -192
rect 254 -188 255 -186
rect 254 -194 255 -192
rect 261 -188 262 -186
rect 261 -194 262 -192
rect 268 -188 269 -186
rect 268 -194 269 -192
rect 275 -188 276 -186
rect 275 -194 276 -192
rect 282 -188 283 -186
rect 282 -194 283 -192
rect 289 -188 290 -186
rect 289 -194 290 -192
rect 296 -188 297 -186
rect 299 -188 300 -186
rect 296 -194 297 -192
rect 303 -188 304 -186
rect 306 -188 307 -186
rect 303 -194 304 -192
rect 310 -188 311 -186
rect 310 -194 311 -192
rect 317 -188 318 -186
rect 324 -188 325 -186
rect 324 -194 325 -192
rect 352 -194 353 -192
rect 359 -188 360 -186
rect 359 -194 360 -192
rect 30 -219 31 -217
rect 30 -225 31 -223
rect 37 -219 38 -217
rect 40 -219 41 -217
rect 40 -225 41 -223
rect 44 -219 45 -217
rect 44 -225 45 -223
rect 54 -219 55 -217
rect 51 -225 52 -223
rect 58 -219 59 -217
rect 58 -225 59 -223
rect 65 -219 66 -217
rect 65 -225 66 -223
rect 72 -219 73 -217
rect 72 -225 73 -223
rect 79 -219 80 -217
rect 82 -219 83 -217
rect 86 -219 87 -217
rect 89 -225 90 -223
rect 93 -219 94 -217
rect 93 -225 94 -223
rect 100 -219 101 -217
rect 103 -219 104 -217
rect 107 -219 108 -217
rect 110 -225 111 -223
rect 114 -219 115 -217
rect 114 -225 115 -223
rect 121 -219 122 -217
rect 121 -225 122 -223
rect 128 -219 129 -217
rect 128 -225 129 -223
rect 135 -219 136 -217
rect 138 -219 139 -217
rect 135 -225 136 -223
rect 142 -219 143 -217
rect 142 -225 143 -223
rect 149 -219 150 -217
rect 149 -225 150 -223
rect 152 -225 153 -223
rect 159 -219 160 -217
rect 156 -225 157 -223
rect 159 -225 160 -223
rect 163 -219 164 -217
rect 163 -225 164 -223
rect 170 -219 171 -217
rect 170 -225 171 -223
rect 177 -219 178 -217
rect 177 -225 178 -223
rect 184 -219 185 -217
rect 187 -219 188 -217
rect 187 -225 188 -223
rect 191 -219 192 -217
rect 191 -225 192 -223
rect 198 -219 199 -217
rect 198 -225 199 -223
rect 205 -219 206 -217
rect 205 -225 206 -223
rect 212 -219 213 -217
rect 215 -219 216 -217
rect 212 -225 213 -223
rect 215 -225 216 -223
rect 219 -219 220 -217
rect 219 -225 220 -223
rect 226 -219 227 -217
rect 226 -225 227 -223
rect 233 -225 234 -223
rect 240 -219 241 -217
rect 240 -225 241 -223
rect 247 -219 248 -217
rect 250 -225 251 -223
rect 254 -219 255 -217
rect 254 -225 255 -223
rect 261 -219 262 -217
rect 261 -225 262 -223
rect 268 -219 269 -217
rect 268 -225 269 -223
rect 275 -219 276 -217
rect 275 -225 276 -223
rect 282 -219 283 -217
rect 282 -225 283 -223
rect 289 -219 290 -217
rect 289 -225 290 -223
rect 296 -219 297 -217
rect 296 -225 297 -223
rect 303 -219 304 -217
rect 303 -225 304 -223
rect 310 -219 311 -217
rect 310 -225 311 -223
rect 320 -225 321 -223
rect 324 -219 325 -217
rect 327 -219 328 -217
rect 327 -225 328 -223
rect 331 -219 332 -217
rect 334 -225 335 -223
rect 341 -219 342 -217
rect 345 -219 346 -217
rect 345 -225 346 -223
rect 352 -219 353 -217
rect 355 -225 356 -223
rect 359 -219 360 -217
rect 359 -225 360 -223
rect 366 -219 367 -217
rect 366 -225 367 -223
rect 373 -219 374 -217
rect 373 -225 374 -223
rect 380 -219 381 -217
rect 380 -225 381 -223
rect 390 -219 391 -217
rect 387 -225 388 -223
rect 9 -248 10 -246
rect 9 -254 10 -252
rect 16 -248 17 -246
rect 16 -254 17 -252
rect 23 -248 24 -246
rect 23 -254 24 -252
rect 33 -248 34 -246
rect 33 -254 34 -252
rect 37 -248 38 -246
rect 44 -248 45 -246
rect 44 -254 45 -252
rect 54 -248 55 -246
rect 51 -254 52 -252
rect 58 -248 59 -246
rect 58 -254 59 -252
rect 65 -248 66 -246
rect 65 -254 66 -252
rect 72 -248 73 -246
rect 72 -254 73 -252
rect 79 -248 80 -246
rect 79 -254 80 -252
rect 86 -248 87 -246
rect 86 -254 87 -252
rect 89 -254 90 -252
rect 93 -248 94 -246
rect 93 -254 94 -252
rect 100 -248 101 -246
rect 100 -254 101 -252
rect 107 -248 108 -246
rect 110 -248 111 -246
rect 107 -254 108 -252
rect 114 -248 115 -246
rect 114 -254 115 -252
rect 121 -248 122 -246
rect 121 -254 122 -252
rect 131 -254 132 -252
rect 135 -248 136 -246
rect 135 -254 136 -252
rect 142 -254 143 -252
rect 145 -254 146 -252
rect 149 -248 150 -246
rect 152 -248 153 -246
rect 149 -254 150 -252
rect 156 -248 157 -246
rect 156 -254 157 -252
rect 163 -248 164 -246
rect 163 -254 164 -252
rect 170 -248 171 -246
rect 173 -248 174 -246
rect 170 -254 171 -252
rect 173 -254 174 -252
rect 177 -248 178 -246
rect 177 -254 178 -252
rect 184 -248 185 -246
rect 184 -254 185 -252
rect 191 -248 192 -246
rect 191 -254 192 -252
rect 198 -248 199 -246
rect 198 -254 199 -252
rect 208 -248 209 -246
rect 205 -254 206 -252
rect 212 -248 213 -246
rect 212 -254 213 -252
rect 222 -248 223 -246
rect 219 -254 220 -252
rect 222 -254 223 -252
rect 226 -248 227 -246
rect 226 -254 227 -252
rect 233 -248 234 -246
rect 233 -254 234 -252
rect 240 -248 241 -246
rect 240 -254 241 -252
rect 247 -248 248 -246
rect 247 -254 248 -252
rect 254 -248 255 -246
rect 254 -254 255 -252
rect 261 -248 262 -246
rect 261 -254 262 -252
rect 268 -248 269 -246
rect 268 -254 269 -252
rect 275 -248 276 -246
rect 275 -254 276 -252
rect 282 -248 283 -246
rect 282 -254 283 -252
rect 289 -248 290 -246
rect 289 -254 290 -252
rect 296 -248 297 -246
rect 296 -254 297 -252
rect 303 -248 304 -246
rect 303 -254 304 -252
rect 310 -248 311 -246
rect 310 -254 311 -252
rect 317 -248 318 -246
rect 317 -254 318 -252
rect 327 -248 328 -246
rect 331 -248 332 -246
rect 331 -254 332 -252
rect 338 -248 339 -246
rect 345 -254 346 -252
rect 352 -248 353 -246
rect 352 -254 353 -252
rect 380 -248 381 -246
rect 387 -254 388 -252
rect 394 -248 395 -246
rect 394 -254 395 -252
rect 2 -295 3 -293
rect 2 -301 3 -299
rect 9 -295 10 -293
rect 16 -295 17 -293
rect 16 -301 17 -299
rect 23 -295 24 -293
rect 23 -301 24 -299
rect 30 -301 31 -299
rect 37 -295 38 -293
rect 37 -301 38 -299
rect 44 -295 45 -293
rect 44 -301 45 -299
rect 54 -295 55 -293
rect 51 -301 52 -299
rect 58 -295 59 -293
rect 58 -301 59 -299
rect 65 -295 66 -293
rect 68 -295 69 -293
rect 65 -301 66 -299
rect 72 -295 73 -293
rect 75 -295 76 -293
rect 79 -295 80 -293
rect 82 -295 83 -293
rect 79 -301 80 -299
rect 86 -295 87 -293
rect 86 -301 87 -299
rect 96 -295 97 -293
rect 96 -301 97 -299
rect 100 -295 101 -293
rect 100 -301 101 -299
rect 107 -295 108 -293
rect 107 -301 108 -299
rect 114 -295 115 -293
rect 117 -301 118 -299
rect 121 -295 122 -293
rect 121 -301 122 -299
rect 128 -295 129 -293
rect 131 -301 132 -299
rect 135 -295 136 -293
rect 135 -301 136 -299
rect 142 -295 143 -293
rect 142 -301 143 -299
rect 149 -295 150 -293
rect 152 -295 153 -293
rect 149 -301 150 -299
rect 156 -295 157 -293
rect 159 -295 160 -293
rect 156 -301 157 -299
rect 163 -295 164 -293
rect 163 -301 164 -299
rect 170 -295 171 -293
rect 170 -301 171 -299
rect 173 -301 174 -299
rect 177 -295 178 -293
rect 180 -295 181 -293
rect 177 -301 178 -299
rect 187 -295 188 -293
rect 184 -301 185 -299
rect 187 -301 188 -299
rect 191 -295 192 -293
rect 194 -295 195 -293
rect 191 -301 192 -299
rect 194 -301 195 -299
rect 198 -295 199 -293
rect 198 -301 199 -299
rect 208 -295 209 -293
rect 205 -301 206 -299
rect 208 -301 209 -299
rect 212 -295 213 -293
rect 215 -295 216 -293
rect 212 -301 213 -299
rect 215 -301 216 -299
rect 219 -295 220 -293
rect 219 -301 220 -299
rect 226 -295 227 -293
rect 226 -301 227 -299
rect 233 -295 234 -293
rect 243 -295 244 -293
rect 243 -301 244 -299
rect 247 -295 248 -293
rect 247 -301 248 -299
rect 254 -295 255 -293
rect 254 -301 255 -299
rect 261 -295 262 -293
rect 261 -301 262 -299
rect 268 -295 269 -293
rect 268 -301 269 -299
rect 275 -295 276 -293
rect 275 -301 276 -299
rect 282 -295 283 -293
rect 282 -301 283 -299
rect 289 -295 290 -293
rect 289 -301 290 -299
rect 296 -295 297 -293
rect 296 -301 297 -299
rect 303 -295 304 -293
rect 303 -301 304 -299
rect 310 -295 311 -293
rect 310 -301 311 -299
rect 317 -295 318 -293
rect 317 -301 318 -299
rect 324 -295 325 -293
rect 324 -301 325 -299
rect 331 -295 332 -293
rect 331 -301 332 -299
rect 338 -295 339 -293
rect 338 -301 339 -299
rect 345 -295 346 -293
rect 345 -301 346 -299
rect 30 -342 31 -340
rect 30 -348 31 -346
rect 37 -342 38 -340
rect 37 -348 38 -346
rect 44 -342 45 -340
rect 44 -348 45 -346
rect 54 -342 55 -340
rect 58 -342 59 -340
rect 58 -348 59 -346
rect 65 -342 66 -340
rect 65 -348 66 -346
rect 75 -342 76 -340
rect 79 -342 80 -340
rect 79 -348 80 -346
rect 86 -342 87 -340
rect 86 -348 87 -346
rect 93 -342 94 -340
rect 93 -348 94 -346
rect 103 -342 104 -340
rect 103 -348 104 -346
rect 110 -342 111 -340
rect 107 -348 108 -346
rect 114 -342 115 -340
rect 117 -348 118 -346
rect 121 -342 122 -340
rect 128 -342 129 -340
rect 128 -348 129 -346
rect 135 -342 136 -340
rect 138 -342 139 -340
rect 135 -348 136 -346
rect 142 -342 143 -340
rect 145 -342 146 -340
rect 145 -348 146 -346
rect 149 -342 150 -340
rect 152 -342 153 -340
rect 152 -348 153 -346
rect 156 -342 157 -340
rect 163 -342 164 -340
rect 163 -348 164 -346
rect 170 -342 171 -340
rect 170 -348 171 -346
rect 177 -342 178 -340
rect 177 -348 178 -346
rect 184 -342 185 -340
rect 187 -342 188 -340
rect 184 -348 185 -346
rect 191 -348 192 -346
rect 194 -348 195 -346
rect 198 -342 199 -340
rect 201 -342 202 -340
rect 201 -348 202 -346
rect 208 -342 209 -340
rect 205 -348 206 -346
rect 212 -342 213 -340
rect 215 -342 216 -340
rect 212 -348 213 -346
rect 219 -342 220 -340
rect 219 -348 220 -346
rect 229 -342 230 -340
rect 233 -342 234 -340
rect 233 -348 234 -346
rect 240 -342 241 -340
rect 243 -348 244 -346
rect 247 -342 248 -340
rect 247 -348 248 -346
rect 254 -342 255 -340
rect 254 -348 255 -346
rect 261 -342 262 -340
rect 261 -348 262 -346
rect 268 -342 269 -340
rect 268 -348 269 -346
rect 275 -342 276 -340
rect 275 -348 276 -346
rect 282 -342 283 -340
rect 282 -348 283 -346
rect 289 -342 290 -340
rect 289 -348 290 -346
rect 296 -342 297 -340
rect 299 -348 300 -346
rect 303 -342 304 -340
rect 303 -348 304 -346
rect 310 -342 311 -340
rect 310 -348 311 -346
rect 317 -342 318 -340
rect 317 -348 318 -346
rect 324 -342 325 -340
rect 324 -348 325 -346
rect 2 -377 3 -375
rect 2 -383 3 -381
rect 9 -377 10 -375
rect 9 -383 10 -381
rect 16 -377 17 -375
rect 16 -383 17 -381
rect 23 -377 24 -375
rect 23 -383 24 -381
rect 30 -383 31 -381
rect 37 -377 38 -375
rect 37 -383 38 -381
rect 44 -377 45 -375
rect 44 -383 45 -381
rect 51 -377 52 -375
rect 51 -383 52 -381
rect 58 -383 59 -381
rect 61 -383 62 -381
rect 65 -377 66 -375
rect 68 -383 69 -381
rect 72 -377 73 -375
rect 75 -377 76 -375
rect 75 -383 76 -381
rect 79 -377 80 -375
rect 79 -383 80 -381
rect 86 -377 87 -375
rect 89 -377 90 -375
rect 89 -383 90 -381
rect 93 -377 94 -375
rect 96 -377 97 -375
rect 93 -383 94 -381
rect 100 -377 101 -375
rect 100 -383 101 -381
rect 107 -377 108 -375
rect 107 -383 108 -381
rect 114 -377 115 -375
rect 117 -377 118 -375
rect 114 -383 115 -381
rect 117 -383 118 -381
rect 121 -377 122 -375
rect 121 -383 122 -381
rect 128 -377 129 -375
rect 128 -383 129 -381
rect 135 -377 136 -375
rect 138 -383 139 -381
rect 142 -377 143 -375
rect 145 -377 146 -375
rect 142 -383 143 -381
rect 149 -377 150 -375
rect 149 -383 150 -381
rect 156 -383 157 -381
rect 163 -377 164 -375
rect 166 -377 167 -375
rect 166 -383 167 -381
rect 170 -377 171 -375
rect 173 -377 174 -375
rect 170 -383 171 -381
rect 180 -377 181 -375
rect 177 -383 178 -381
rect 180 -383 181 -381
rect 184 -383 185 -381
rect 191 -377 192 -375
rect 191 -383 192 -381
rect 194 -383 195 -381
rect 198 -377 199 -375
rect 198 -383 199 -381
rect 205 -377 206 -375
rect 205 -383 206 -381
rect 212 -377 213 -375
rect 215 -377 216 -375
rect 215 -383 216 -381
rect 219 -377 220 -375
rect 219 -383 220 -381
rect 226 -377 227 -375
rect 226 -383 227 -381
rect 233 -377 234 -375
rect 233 -383 234 -381
rect 240 -377 241 -375
rect 240 -383 241 -381
rect 247 -377 248 -375
rect 247 -383 248 -381
rect 254 -377 255 -375
rect 254 -383 255 -381
rect 264 -377 265 -375
rect 261 -383 262 -381
rect 268 -377 269 -375
rect 268 -383 269 -381
rect 275 -377 276 -375
rect 275 -383 276 -381
rect 282 -377 283 -375
rect 282 -383 283 -381
rect 289 -377 290 -375
rect 289 -383 290 -381
rect 296 -377 297 -375
rect 296 -383 297 -381
rect 306 -383 307 -381
rect 310 -377 311 -375
rect 310 -383 311 -381
rect 317 -377 318 -375
rect 317 -383 318 -381
rect 324 -377 325 -375
rect 324 -383 325 -381
rect 331 -377 332 -375
rect 331 -383 332 -381
rect 338 -377 339 -375
rect 338 -383 339 -381
rect 345 -377 346 -375
rect 345 -383 346 -381
rect 23 -418 24 -416
rect 23 -424 24 -422
rect 30 -418 31 -416
rect 30 -424 31 -422
rect 40 -418 41 -416
rect 37 -424 38 -422
rect 44 -418 45 -416
rect 44 -424 45 -422
rect 51 -418 52 -416
rect 54 -418 55 -416
rect 54 -424 55 -422
rect 58 -418 59 -416
rect 58 -424 59 -422
rect 65 -418 66 -416
rect 65 -424 66 -422
rect 75 -418 76 -416
rect 72 -424 73 -422
rect 79 -418 80 -416
rect 82 -418 83 -416
rect 86 -418 87 -416
rect 86 -424 87 -422
rect 96 -418 97 -416
rect 93 -424 94 -422
rect 96 -424 97 -422
rect 103 -418 104 -416
rect 107 -418 108 -416
rect 107 -424 108 -422
rect 128 -418 129 -416
rect 128 -424 129 -422
rect 135 -418 136 -416
rect 135 -424 136 -422
rect 142 -418 143 -416
rect 142 -424 143 -422
rect 149 -418 150 -416
rect 152 -418 153 -416
rect 156 -418 157 -416
rect 156 -424 157 -422
rect 163 -418 164 -416
rect 163 -424 164 -422
rect 170 -424 171 -422
rect 173 -424 174 -422
rect 177 -418 178 -416
rect 177 -424 178 -422
rect 184 -418 185 -416
rect 184 -424 185 -422
rect 191 -418 192 -416
rect 191 -424 192 -422
rect 198 -418 199 -416
rect 201 -418 202 -416
rect 201 -424 202 -422
rect 205 -418 206 -416
rect 205 -424 206 -422
rect 212 -418 213 -416
rect 215 -418 216 -416
rect 219 -418 220 -416
rect 219 -424 220 -422
rect 222 -424 223 -422
rect 226 -418 227 -416
rect 226 -424 227 -422
rect 229 -424 230 -422
rect 233 -418 234 -416
rect 233 -424 234 -422
rect 243 -418 244 -416
rect 247 -418 248 -416
rect 247 -424 248 -422
rect 254 -418 255 -416
rect 254 -424 255 -422
rect 261 -418 262 -416
rect 261 -424 262 -422
rect 268 -418 269 -416
rect 271 -418 272 -416
rect 268 -424 269 -422
rect 275 -418 276 -416
rect 275 -424 276 -422
rect 282 -418 283 -416
rect 285 -418 286 -416
rect 282 -424 283 -422
rect 289 -418 290 -416
rect 292 -418 293 -416
rect 296 -418 297 -416
rect 296 -424 297 -422
rect 303 -418 304 -416
rect 303 -424 304 -422
rect 310 -418 311 -416
rect 310 -424 311 -422
rect 317 -418 318 -416
rect 317 -424 318 -422
rect 2 -449 3 -447
rect 2 -455 3 -453
rect 9 -449 10 -447
rect 9 -455 10 -453
rect 16 -449 17 -447
rect 16 -455 17 -453
rect 23 -449 24 -447
rect 23 -455 24 -453
rect 30 -449 31 -447
rect 30 -455 31 -453
rect 37 -449 38 -447
rect 37 -455 38 -453
rect 47 -449 48 -447
rect 44 -455 45 -453
rect 51 -449 52 -447
rect 51 -455 52 -453
rect 58 -449 59 -447
rect 58 -455 59 -453
rect 61 -455 62 -453
rect 65 -449 66 -447
rect 65 -455 66 -453
rect 72 -449 73 -447
rect 75 -455 76 -453
rect 79 -449 80 -447
rect 82 -449 83 -447
rect 79 -455 80 -453
rect 89 -449 90 -447
rect 86 -455 87 -453
rect 89 -455 90 -453
rect 93 -449 94 -447
rect 93 -455 94 -453
rect 103 -449 104 -447
rect 100 -455 101 -453
rect 103 -455 104 -453
rect 107 -449 108 -447
rect 110 -449 111 -447
rect 110 -455 111 -453
rect 114 -449 115 -447
rect 114 -455 115 -453
rect 121 -449 122 -447
rect 121 -455 122 -453
rect 128 -449 129 -447
rect 131 -449 132 -447
rect 128 -455 129 -453
rect 135 -449 136 -447
rect 135 -455 136 -453
rect 138 -455 139 -453
rect 142 -449 143 -447
rect 142 -455 143 -453
rect 149 -449 150 -447
rect 149 -455 150 -453
rect 156 -449 157 -447
rect 159 -455 160 -453
rect 163 -449 164 -447
rect 163 -455 164 -453
rect 170 -449 171 -447
rect 173 -455 174 -453
rect 177 -449 178 -447
rect 177 -455 178 -453
rect 184 -449 185 -447
rect 184 -455 185 -453
rect 191 -449 192 -447
rect 194 -449 195 -447
rect 194 -455 195 -453
rect 201 -449 202 -447
rect 205 -449 206 -447
rect 205 -455 206 -453
rect 212 -449 213 -447
rect 212 -455 213 -453
rect 215 -455 216 -453
rect 219 -449 220 -447
rect 219 -455 220 -453
rect 226 -449 227 -447
rect 226 -455 227 -453
rect 233 -449 234 -447
rect 233 -455 234 -453
rect 236 -455 237 -453
rect 240 -449 241 -447
rect 240 -455 241 -453
rect 247 -449 248 -447
rect 247 -455 248 -453
rect 254 -449 255 -447
rect 254 -455 255 -453
rect 261 -449 262 -447
rect 261 -455 262 -453
rect 268 -449 269 -447
rect 268 -455 269 -453
rect 275 -449 276 -447
rect 275 -455 276 -453
rect 282 -449 283 -447
rect 282 -455 283 -453
rect 289 -449 290 -447
rect 289 -455 290 -453
rect 296 -449 297 -447
rect 296 -455 297 -453
rect 303 -449 304 -447
rect 303 -455 304 -453
rect 310 -449 311 -447
rect 310 -455 311 -453
rect 317 -449 318 -447
rect 317 -455 318 -453
rect 324 -449 325 -447
rect 327 -449 328 -447
rect 327 -455 328 -453
rect 334 -455 335 -453
rect 338 -449 339 -447
rect 338 -455 339 -453
rect 40 -490 41 -488
rect 44 -490 45 -488
rect 44 -496 45 -494
rect 51 -490 52 -488
rect 51 -496 52 -494
rect 58 -490 59 -488
rect 58 -496 59 -494
rect 65 -490 66 -488
rect 65 -496 66 -494
rect 75 -490 76 -488
rect 72 -496 73 -494
rect 82 -496 83 -494
rect 86 -490 87 -488
rect 86 -496 87 -494
rect 93 -490 94 -488
rect 93 -496 94 -494
rect 100 -490 101 -488
rect 100 -496 101 -494
rect 107 -490 108 -488
rect 107 -496 108 -494
rect 114 -490 115 -488
rect 114 -496 115 -494
rect 121 -490 122 -488
rect 124 -496 125 -494
rect 128 -490 129 -488
rect 131 -490 132 -488
rect 128 -496 129 -494
rect 138 -490 139 -488
rect 138 -496 139 -494
rect 142 -490 143 -488
rect 145 -490 146 -488
rect 145 -496 146 -494
rect 149 -490 150 -488
rect 149 -496 150 -494
rect 156 -490 157 -488
rect 156 -496 157 -494
rect 163 -490 164 -488
rect 163 -496 164 -494
rect 170 -490 171 -488
rect 170 -496 171 -494
rect 177 -490 178 -488
rect 180 -490 181 -488
rect 180 -496 181 -494
rect 184 -490 185 -488
rect 184 -496 185 -494
rect 191 -490 192 -488
rect 191 -496 192 -494
rect 198 -490 199 -488
rect 198 -496 199 -494
rect 201 -496 202 -494
rect 205 -490 206 -488
rect 205 -496 206 -494
rect 215 -490 216 -488
rect 219 -490 220 -488
rect 222 -490 223 -488
rect 222 -496 223 -494
rect 226 -490 227 -488
rect 226 -496 227 -494
rect 233 -490 234 -488
rect 233 -496 234 -494
rect 240 -490 241 -488
rect 240 -496 241 -494
rect 247 -490 248 -488
rect 247 -496 248 -494
rect 254 -496 255 -494
rect 257 -496 258 -494
rect 261 -490 262 -488
rect 261 -496 262 -494
rect 268 -490 269 -488
rect 268 -496 269 -494
rect 275 -490 276 -488
rect 275 -496 276 -494
rect 282 -496 283 -494
rect 289 -490 290 -488
rect 289 -496 290 -494
rect 296 -490 297 -488
rect 296 -496 297 -494
rect 303 -490 304 -488
rect 303 -496 304 -494
rect 310 -490 311 -488
rect 310 -496 311 -494
rect 317 -490 318 -488
rect 320 -490 321 -488
rect 320 -496 321 -494
rect 327 -496 328 -494
rect 331 -490 332 -488
rect 331 -496 332 -494
rect 338 -490 339 -488
rect 338 -496 339 -494
rect 348 -496 349 -494
rect 352 -490 353 -488
rect 352 -496 353 -494
rect 359 -490 360 -488
rect 359 -496 360 -494
rect 366 -490 367 -488
rect 16 -527 17 -525
rect 16 -533 17 -531
rect 23 -527 24 -525
rect 23 -533 24 -531
rect 30 -527 31 -525
rect 30 -533 31 -531
rect 37 -533 38 -531
rect 44 -527 45 -525
rect 44 -533 45 -531
rect 51 -527 52 -525
rect 51 -533 52 -531
rect 61 -527 62 -525
rect 58 -533 59 -531
rect 61 -533 62 -531
rect 65 -527 66 -525
rect 65 -533 66 -531
rect 72 -527 73 -525
rect 72 -533 73 -531
rect 79 -527 80 -525
rect 82 -527 83 -525
rect 82 -533 83 -531
rect 86 -527 87 -525
rect 86 -533 87 -531
rect 93 -527 94 -525
rect 93 -533 94 -531
rect 100 -527 101 -525
rect 103 -527 104 -525
rect 103 -533 104 -531
rect 107 -527 108 -525
rect 107 -533 108 -531
rect 114 -527 115 -525
rect 114 -533 115 -531
rect 121 -527 122 -525
rect 124 -533 125 -531
rect 128 -527 129 -525
rect 128 -533 129 -531
rect 135 -527 136 -525
rect 135 -533 136 -531
rect 138 -533 139 -531
rect 142 -527 143 -525
rect 142 -533 143 -531
rect 149 -527 150 -525
rect 149 -533 150 -531
rect 156 -527 157 -525
rect 159 -527 160 -525
rect 156 -533 157 -531
rect 159 -533 160 -531
rect 163 -527 164 -525
rect 166 -527 167 -525
rect 163 -533 164 -531
rect 166 -533 167 -531
rect 170 -527 171 -525
rect 170 -533 171 -531
rect 177 -527 178 -525
rect 180 -527 181 -525
rect 180 -533 181 -531
rect 184 -527 185 -525
rect 184 -533 185 -531
rect 194 -527 195 -525
rect 191 -533 192 -531
rect 194 -533 195 -531
rect 198 -527 199 -525
rect 201 -527 202 -525
rect 201 -533 202 -531
rect 205 -527 206 -525
rect 208 -533 209 -531
rect 212 -527 213 -525
rect 212 -533 213 -531
rect 215 -533 216 -531
rect 219 -527 220 -525
rect 219 -533 220 -531
rect 226 -527 227 -525
rect 229 -527 230 -525
rect 233 -527 234 -525
rect 233 -533 234 -531
rect 240 -527 241 -525
rect 240 -533 241 -531
rect 247 -527 248 -525
rect 247 -533 248 -531
rect 254 -527 255 -525
rect 254 -533 255 -531
rect 261 -527 262 -525
rect 261 -533 262 -531
rect 271 -527 272 -525
rect 268 -533 269 -531
rect 271 -533 272 -531
rect 275 -527 276 -525
rect 275 -533 276 -531
rect 282 -527 283 -525
rect 282 -533 283 -531
rect 289 -527 290 -525
rect 289 -533 290 -531
rect 296 -527 297 -525
rect 296 -533 297 -531
rect 303 -527 304 -525
rect 303 -533 304 -531
rect 310 -527 311 -525
rect 310 -533 311 -531
rect 317 -527 318 -525
rect 317 -533 318 -531
rect 324 -527 325 -525
rect 324 -533 325 -531
rect 331 -527 332 -525
rect 331 -533 332 -531
rect 338 -527 339 -525
rect 338 -533 339 -531
rect 345 -527 346 -525
rect 345 -533 346 -531
rect 352 -527 353 -525
rect 352 -533 353 -531
rect 9 -570 10 -568
rect 9 -576 10 -574
rect 16 -570 17 -568
rect 16 -576 17 -574
rect 23 -570 24 -568
rect 23 -576 24 -574
rect 33 -570 34 -568
rect 40 -570 41 -568
rect 44 -576 45 -574
rect 51 -570 52 -568
rect 51 -576 52 -574
rect 58 -570 59 -568
rect 61 -570 62 -568
rect 61 -576 62 -574
rect 65 -570 66 -568
rect 68 -570 69 -568
rect 72 -570 73 -568
rect 72 -576 73 -574
rect 82 -570 83 -568
rect 79 -576 80 -574
rect 86 -570 87 -568
rect 86 -576 87 -574
rect 93 -570 94 -568
rect 93 -576 94 -574
rect 100 -570 101 -568
rect 100 -576 101 -574
rect 107 -570 108 -568
rect 117 -570 118 -568
rect 114 -576 115 -574
rect 121 -570 122 -568
rect 121 -576 122 -574
rect 128 -570 129 -568
rect 128 -576 129 -574
rect 135 -570 136 -568
rect 135 -576 136 -574
rect 142 -570 143 -568
rect 142 -576 143 -574
rect 149 -576 150 -574
rect 156 -570 157 -568
rect 156 -576 157 -574
rect 163 -570 164 -568
rect 166 -570 167 -568
rect 163 -576 164 -574
rect 170 -570 171 -568
rect 170 -576 171 -574
rect 177 -570 178 -568
rect 177 -576 178 -574
rect 180 -576 181 -574
rect 184 -570 185 -568
rect 184 -576 185 -574
rect 191 -570 192 -568
rect 191 -576 192 -574
rect 198 -570 199 -568
rect 198 -576 199 -574
rect 205 -570 206 -568
rect 205 -576 206 -574
rect 212 -570 213 -568
rect 212 -576 213 -574
rect 219 -570 220 -568
rect 222 -570 223 -568
rect 219 -576 220 -574
rect 222 -576 223 -574
rect 226 -570 227 -568
rect 226 -576 227 -574
rect 233 -570 234 -568
rect 233 -576 234 -574
rect 236 -576 237 -574
rect 243 -570 244 -568
rect 240 -576 241 -574
rect 243 -576 244 -574
rect 247 -570 248 -568
rect 250 -570 251 -568
rect 250 -576 251 -574
rect 254 -570 255 -568
rect 254 -576 255 -574
rect 261 -570 262 -568
rect 261 -576 262 -574
rect 268 -570 269 -568
rect 268 -576 269 -574
rect 275 -570 276 -568
rect 275 -576 276 -574
rect 282 -570 283 -568
rect 282 -576 283 -574
rect 289 -570 290 -568
rect 289 -576 290 -574
rect 296 -570 297 -568
rect 296 -576 297 -574
rect 303 -570 304 -568
rect 303 -576 304 -574
rect 310 -570 311 -568
rect 310 -576 311 -574
rect 317 -570 318 -568
rect 317 -576 318 -574
rect 324 -570 325 -568
rect 324 -576 325 -574
rect 331 -570 332 -568
rect 331 -576 332 -574
rect 338 -570 339 -568
rect 338 -576 339 -574
rect 345 -570 346 -568
rect 345 -576 346 -574
rect 352 -570 353 -568
rect 352 -576 353 -574
rect 362 -570 363 -568
rect 359 -576 360 -574
rect 369 -570 370 -568
rect 369 -576 370 -574
rect 44 -607 45 -605
rect 47 -607 48 -605
rect 51 -607 52 -605
rect 51 -613 52 -611
rect 68 -607 69 -605
rect 68 -613 69 -611
rect 72 -607 73 -605
rect 72 -613 73 -611
rect 79 -607 80 -605
rect 86 -607 87 -605
rect 86 -613 87 -611
rect 93 -607 94 -605
rect 93 -613 94 -611
rect 100 -607 101 -605
rect 103 -607 104 -605
rect 110 -607 111 -605
rect 110 -613 111 -611
rect 114 -607 115 -605
rect 114 -613 115 -611
rect 121 -607 122 -605
rect 121 -613 122 -611
rect 124 -613 125 -611
rect 128 -607 129 -605
rect 128 -613 129 -611
rect 135 -607 136 -605
rect 135 -613 136 -611
rect 145 -607 146 -605
rect 142 -613 143 -611
rect 149 -607 150 -605
rect 152 -607 153 -605
rect 156 -607 157 -605
rect 156 -613 157 -611
rect 163 -607 164 -605
rect 163 -613 164 -611
rect 166 -613 167 -611
rect 170 -607 171 -605
rect 170 -613 171 -611
rect 177 -607 178 -605
rect 177 -613 178 -611
rect 187 -607 188 -605
rect 184 -613 185 -611
rect 187 -613 188 -611
rect 191 -607 192 -605
rect 191 -613 192 -611
rect 194 -613 195 -611
rect 198 -607 199 -605
rect 198 -613 199 -611
rect 205 -607 206 -605
rect 205 -613 206 -611
rect 212 -607 213 -605
rect 212 -613 213 -611
rect 219 -607 220 -605
rect 219 -613 220 -611
rect 229 -607 230 -605
rect 233 -607 234 -605
rect 233 -613 234 -611
rect 240 -607 241 -605
rect 240 -613 241 -611
rect 247 -607 248 -605
rect 250 -607 251 -605
rect 250 -613 251 -611
rect 254 -607 255 -605
rect 257 -607 258 -605
rect 257 -613 258 -611
rect 261 -607 262 -605
rect 264 -607 265 -605
rect 268 -607 269 -605
rect 268 -613 269 -611
rect 275 -607 276 -605
rect 275 -613 276 -611
rect 282 -607 283 -605
rect 282 -613 283 -611
rect 292 -607 293 -605
rect 289 -613 290 -611
rect 310 -607 311 -605
rect 310 -613 311 -611
rect 44 -644 45 -642
rect 51 -638 52 -636
rect 51 -644 52 -642
rect 58 -638 59 -636
rect 58 -644 59 -642
rect 65 -638 66 -636
rect 68 -638 69 -636
rect 65 -644 66 -642
rect 72 -638 73 -636
rect 72 -644 73 -642
rect 79 -638 80 -636
rect 79 -644 80 -642
rect 82 -644 83 -642
rect 86 -638 87 -636
rect 86 -644 87 -642
rect 96 -638 97 -636
rect 93 -644 94 -642
rect 96 -644 97 -642
rect 100 -638 101 -636
rect 103 -638 104 -636
rect 107 -638 108 -636
rect 107 -644 108 -642
rect 114 -638 115 -636
rect 114 -644 115 -642
rect 124 -644 125 -642
rect 128 -638 129 -636
rect 128 -644 129 -642
rect 138 -638 139 -636
rect 142 -638 143 -636
rect 142 -644 143 -642
rect 149 -644 150 -642
rect 152 -644 153 -642
rect 156 -638 157 -636
rect 156 -644 157 -642
rect 163 -638 164 -636
rect 163 -644 164 -642
rect 170 -638 171 -636
rect 173 -644 174 -642
rect 177 -638 178 -636
rect 180 -644 181 -642
rect 184 -638 185 -636
rect 184 -644 185 -642
rect 191 -644 192 -642
rect 194 -644 195 -642
rect 198 -638 199 -636
rect 198 -644 199 -642
rect 208 -638 209 -636
rect 208 -644 209 -642
rect 212 -638 213 -636
rect 212 -644 213 -642
rect 219 -638 220 -636
rect 219 -644 220 -642
rect 226 -638 227 -636
rect 226 -644 227 -642
rect 233 -638 234 -636
rect 233 -644 234 -642
rect 240 -638 241 -636
rect 240 -644 241 -642
rect 247 -638 248 -636
rect 247 -644 248 -642
rect 254 -638 255 -636
rect 254 -644 255 -642
rect 261 -638 262 -636
rect 261 -644 262 -642
rect 268 -638 269 -636
rect 268 -644 269 -642
rect 275 -638 276 -636
rect 275 -644 276 -642
rect 282 -638 283 -636
rect 282 -644 283 -642
rect 289 -638 290 -636
rect 292 -638 293 -636
rect 299 -638 300 -636
rect 303 -638 304 -636
rect 303 -644 304 -642
rect 313 -638 314 -636
rect 310 -644 311 -642
rect 44 -665 45 -663
rect 44 -671 45 -669
rect 54 -665 55 -663
rect 58 -671 59 -669
rect 65 -665 66 -663
rect 65 -671 66 -669
rect 72 -665 73 -663
rect 72 -671 73 -669
rect 79 -665 80 -663
rect 79 -671 80 -669
rect 89 -665 90 -663
rect 86 -671 87 -669
rect 93 -671 94 -669
rect 96 -671 97 -669
rect 100 -665 101 -663
rect 100 -671 101 -669
rect 107 -665 108 -663
rect 107 -671 108 -669
rect 114 -665 115 -663
rect 114 -671 115 -669
rect 121 -665 122 -663
rect 124 -671 125 -669
rect 135 -665 136 -663
rect 138 -671 139 -669
rect 142 -665 143 -663
rect 149 -665 150 -663
rect 149 -671 150 -669
rect 170 -665 171 -663
rect 170 -671 171 -669
rect 180 -671 181 -669
rect 184 -665 185 -663
rect 184 -671 185 -669
rect 191 -665 192 -663
rect 191 -671 192 -669
rect 201 -665 202 -663
rect 201 -671 202 -669
rect 205 -665 206 -663
rect 205 -671 206 -669
rect 212 -665 213 -663
rect 222 -665 223 -663
rect 219 -671 220 -669
rect 226 -665 227 -663
rect 226 -671 227 -669
rect 233 -665 234 -663
rect 233 -671 234 -669
rect 240 -665 241 -663
rect 243 -665 244 -663
rect 240 -671 241 -669
rect 243 -671 244 -669
rect 254 -665 255 -663
rect 254 -671 255 -669
rect 261 -665 262 -663
rect 264 -665 265 -663
rect 268 -665 269 -663
rect 268 -671 269 -669
rect 278 -665 279 -663
rect 282 -665 283 -663
rect 285 -671 286 -669
rect 292 -665 293 -663
rect 292 -671 293 -669
rect 44 -686 45 -684
rect 51 -680 52 -678
rect 51 -686 52 -684
rect 58 -680 59 -678
rect 58 -686 59 -684
rect 65 -680 66 -678
rect 72 -680 73 -678
rect 72 -686 73 -684
rect 79 -680 80 -678
rect 79 -686 80 -684
rect 86 -686 87 -684
rect 93 -686 94 -684
rect 103 -680 104 -678
rect 107 -686 108 -684
rect 114 -686 115 -684
rect 117 -686 118 -684
rect 121 -680 122 -678
rect 121 -686 122 -684
rect 128 -680 129 -678
rect 128 -686 129 -684
rect 135 -680 136 -678
rect 135 -686 136 -684
rect 145 -680 146 -678
rect 142 -686 143 -684
rect 145 -686 146 -684
rect 152 -686 153 -684
rect 191 -680 192 -678
rect 201 -680 202 -678
rect 198 -686 199 -684
rect 205 -680 206 -678
rect 205 -686 206 -684
rect 212 -680 213 -678
rect 212 -686 213 -684
rect 222 -686 223 -684
rect 226 -680 227 -678
rect 226 -686 227 -684
rect 233 -686 234 -684
rect 240 -680 241 -678
rect 243 -686 244 -684
rect 247 -680 248 -678
rect 247 -686 248 -684
rect 254 -680 255 -678
rect 254 -686 255 -684
rect 264 -686 265 -684
rect 275 -680 276 -678
rect 275 -686 276 -684
rect 285 -686 286 -684
<< metal1 >>
rect 135 0 146 1
rect 142 -2 150 -1
rect 100 -13 108 -12
rect 121 -13 164 -12
rect 177 -13 181 -12
rect 128 -15 171 -14
rect 177 -15 185 -14
rect 135 -17 143 -16
rect 149 -17 160 -16
rect 135 -19 146 -18
rect 152 -19 157 -18
rect 79 -30 118 -29
rect 128 -30 136 -29
rect 142 -30 153 -29
rect 159 -30 220 -29
rect 86 -32 150 -31
rect 170 -32 227 -31
rect 93 -34 104 -33
rect 121 -34 143 -33
rect 170 -34 185 -33
rect 191 -34 213 -33
rect 100 -36 108 -35
rect 135 -36 153 -35
rect 163 -36 185 -35
rect 194 -36 199 -35
rect 156 -38 164 -37
rect 180 -38 206 -37
rect 79 -49 108 -48
rect 114 -49 122 -48
rect 128 -49 178 -48
rect 180 -49 220 -48
rect 222 -49 234 -48
rect 79 -51 139 -50
rect 145 -51 206 -50
rect 86 -53 111 -52
rect 114 -53 136 -52
rect 145 -53 227 -52
rect 86 -55 94 -54
rect 100 -55 153 -54
rect 156 -55 185 -54
rect 191 -55 206 -54
rect 93 -57 157 -56
rect 170 -57 227 -56
rect 131 -59 143 -58
rect 149 -59 213 -58
rect 110 -61 143 -60
rect 163 -61 171 -60
rect 187 -61 192 -60
rect 198 -61 213 -60
rect 149 -63 164 -62
rect 72 -74 125 -73
rect 135 -74 157 -73
rect 159 -74 227 -73
rect 243 -74 269 -73
rect 79 -76 129 -75
rect 138 -76 178 -75
rect 184 -76 199 -75
rect 205 -76 220 -75
rect 222 -76 255 -75
rect 261 -76 283 -75
rect 79 -78 94 -77
rect 121 -78 132 -77
rect 138 -78 213 -77
rect 86 -80 108 -79
rect 142 -80 213 -79
rect 65 -82 87 -81
rect 93 -82 108 -81
rect 152 -82 199 -81
rect 205 -82 248 -81
rect 100 -84 122 -83
rect 156 -84 241 -83
rect 100 -86 143 -85
rect 163 -86 178 -85
rect 191 -86 227 -85
rect 114 -88 164 -87
rect 114 -90 171 -89
rect 170 -92 192 -91
rect 44 -103 52 -102
rect 65 -103 129 -102
rect 142 -103 178 -102
rect 198 -103 223 -102
rect 254 -103 265 -102
rect 268 -103 297 -102
rect 299 -103 304 -102
rect 65 -105 76 -104
rect 79 -105 108 -104
rect 131 -105 143 -104
rect 149 -105 157 -104
rect 159 -105 244 -104
rect 247 -105 255 -104
rect 282 -105 290 -104
rect 72 -107 174 -106
rect 205 -107 283 -106
rect 86 -109 94 -108
rect 100 -109 108 -108
rect 117 -109 150 -108
rect 152 -109 164 -108
rect 170 -109 185 -108
rect 212 -109 241 -108
rect 93 -111 136 -110
rect 138 -111 206 -110
rect 212 -111 220 -110
rect 226 -111 248 -110
rect 100 -113 122 -112
rect 156 -113 262 -112
rect 114 -115 122 -114
rect 163 -115 202 -114
rect 219 -115 276 -114
rect 58 -117 115 -116
rect 177 -117 185 -116
rect 191 -117 227 -116
rect 19 -128 24 -127
rect 30 -128 34 -127
rect 47 -128 52 -127
rect 58 -128 97 -127
rect 100 -128 129 -127
rect 135 -128 178 -127
rect 184 -128 213 -127
rect 240 -128 269 -127
rect 289 -128 300 -127
rect 310 -128 325 -127
rect 331 -128 346 -127
rect 58 -130 73 -129
rect 79 -130 87 -129
rect 107 -130 115 -129
rect 149 -130 157 -129
rect 159 -130 171 -129
rect 177 -130 255 -129
rect 271 -130 290 -129
rect 296 -130 304 -129
rect 324 -130 342 -129
rect 65 -132 83 -131
rect 93 -132 115 -131
rect 121 -132 150 -131
rect 156 -132 220 -131
rect 254 -132 262 -131
rect 275 -132 304 -131
rect 37 -134 66 -133
rect 68 -134 87 -133
rect 93 -134 101 -133
rect 107 -134 167 -133
rect 191 -134 234 -133
rect 236 -134 262 -133
rect 79 -136 174 -135
rect 198 -136 283 -135
rect 121 -138 153 -137
rect 163 -138 241 -137
rect 247 -138 283 -137
rect 163 -140 185 -139
rect 201 -140 276 -139
rect 170 -142 192 -141
rect 205 -142 318 -141
rect 194 -144 206 -143
rect 226 -144 248 -143
rect 131 -146 227 -145
rect 19 -157 24 -156
rect 37 -157 69 -156
rect 72 -157 108 -156
rect 114 -157 125 -156
rect 152 -157 206 -156
rect 212 -157 276 -156
rect 296 -157 307 -156
rect 310 -157 335 -156
rect 345 -157 360 -156
rect 44 -159 101 -158
rect 107 -159 129 -158
rect 163 -159 269 -158
rect 296 -159 311 -158
rect 51 -161 62 -160
rect 79 -161 118 -160
rect 128 -161 160 -160
rect 163 -161 192 -160
rect 201 -161 248 -160
rect 303 -161 314 -160
rect 51 -163 59 -162
rect 86 -163 94 -162
rect 114 -163 181 -162
rect 184 -163 216 -162
rect 219 -163 227 -162
rect 303 -163 325 -162
rect 58 -165 80 -164
rect 86 -165 234 -164
rect 313 -165 325 -164
rect 93 -167 136 -166
rect 149 -167 192 -166
rect 198 -167 248 -166
rect 135 -169 178 -168
rect 180 -169 318 -168
rect 142 -171 150 -170
rect 156 -171 185 -170
rect 198 -171 241 -170
rect 268 -171 318 -170
rect 166 -173 227 -172
rect 233 -173 300 -172
rect 173 -175 290 -174
rect 121 -177 174 -176
rect 205 -177 276 -176
rect 100 -179 122 -178
rect 254 -179 290 -178
rect 254 -181 283 -180
rect 261 -183 283 -182
rect 212 -185 262 -184
rect 30 -196 73 -195
rect 79 -196 83 -195
rect 86 -196 146 -195
rect 159 -196 220 -195
rect 229 -196 283 -195
rect 296 -196 325 -195
rect 331 -196 346 -195
rect 359 -196 391 -195
rect 37 -198 62 -197
rect 72 -198 115 -197
rect 121 -198 139 -197
rect 159 -198 262 -197
rect 296 -198 311 -197
rect 352 -198 360 -197
rect 373 -198 381 -197
rect 40 -200 55 -199
rect 58 -200 87 -199
rect 100 -200 206 -199
rect 212 -200 255 -199
rect 303 -200 311 -199
rect 352 -200 367 -199
rect 44 -202 115 -201
rect 135 -202 171 -201
rect 180 -202 328 -201
rect 44 -204 80 -203
rect 103 -204 118 -203
rect 135 -204 283 -203
rect 303 -204 342 -203
rect 51 -206 69 -205
rect 107 -206 143 -205
rect 163 -206 178 -205
rect 187 -206 199 -205
rect 215 -206 220 -205
rect 240 -206 276 -205
rect 65 -208 101 -207
rect 128 -208 143 -207
rect 149 -208 164 -207
rect 184 -208 199 -207
rect 233 -208 276 -207
rect 107 -210 129 -209
rect 149 -210 209 -209
rect 243 -210 269 -209
rect 215 -212 269 -211
rect 247 -214 262 -213
rect 240 -216 248 -215
rect 254 -216 325 -215
rect 9 -227 41 -226
rect 54 -227 101 -226
rect 107 -227 122 -226
rect 128 -227 157 -226
rect 177 -227 216 -226
rect 222 -227 290 -226
rect 310 -227 332 -226
rect 334 -227 374 -226
rect 387 -227 395 -226
rect 16 -229 45 -228
rect 79 -229 157 -228
rect 159 -229 178 -228
rect 212 -229 339 -228
rect 345 -229 353 -228
rect 355 -229 360 -228
rect 23 -231 59 -230
rect 93 -231 213 -230
rect 233 -231 276 -230
rect 282 -231 318 -230
rect 327 -231 367 -230
rect 30 -233 90 -232
rect 93 -233 188 -232
rect 226 -233 276 -232
rect 289 -233 321 -232
rect 33 -235 311 -234
rect 37 -237 111 -236
rect 114 -237 136 -236
rect 149 -237 174 -236
rect 198 -237 227 -236
rect 233 -237 255 -236
rect 268 -237 283 -236
rect 303 -237 328 -236
rect 51 -239 111 -238
rect 114 -239 122 -238
rect 135 -239 143 -238
rect 149 -239 164 -238
rect 191 -239 199 -238
rect 205 -239 304 -238
rect 58 -241 73 -240
rect 152 -241 164 -240
rect 170 -241 192 -240
rect 208 -241 255 -240
rect 44 -243 153 -242
rect 170 -243 185 -242
rect 240 -243 248 -242
rect 250 -243 262 -242
rect 72 -245 87 -244
rect 219 -245 241 -244
rect 261 -245 269 -244
rect 9 -256 34 -255
rect 37 -256 199 -255
rect 205 -256 234 -255
rect 268 -256 297 -255
rect 345 -256 353 -255
rect 387 -256 395 -255
rect 9 -258 69 -257
rect 72 -258 83 -257
rect 89 -258 115 -257
rect 128 -258 227 -257
rect 16 -260 143 -259
rect 145 -260 339 -259
rect 16 -262 115 -261
rect 135 -262 143 -261
rect 149 -262 346 -261
rect 23 -264 76 -263
rect 79 -264 192 -263
rect 208 -264 248 -263
rect 23 -266 80 -265
rect 93 -266 132 -265
rect 149 -266 304 -265
rect 51 -268 164 -267
rect 173 -268 213 -267
rect 215 -268 318 -267
rect 54 -270 244 -269
rect 289 -270 304 -269
rect 310 -270 318 -269
rect 58 -272 87 -271
rect 100 -272 136 -271
rect 156 -272 220 -271
rect 226 -272 241 -271
rect 254 -272 311 -271
rect 58 -274 66 -273
rect 72 -274 87 -273
rect 100 -274 153 -273
rect 159 -274 248 -273
rect 254 -274 276 -273
rect 2 -276 66 -275
rect 107 -276 164 -275
rect 170 -276 220 -275
rect 233 -276 290 -275
rect 107 -278 122 -277
rect 170 -278 199 -277
rect 212 -278 325 -277
rect 121 -280 188 -279
rect 191 -280 332 -279
rect 156 -282 332 -281
rect 177 -284 269 -283
rect 44 -286 178 -285
rect 180 -286 262 -285
rect 44 -288 97 -287
rect 184 -288 297 -287
rect 194 -290 276 -289
rect 222 -292 262 -291
rect 2 -303 31 -302
rect 44 -303 192 -302
rect 205 -303 290 -302
rect 16 -305 76 -304
rect 79 -305 150 -304
rect 170 -305 269 -304
rect 23 -307 55 -306
rect 65 -307 164 -306
rect 187 -307 255 -306
rect 261 -307 290 -306
rect 30 -309 59 -308
rect 65 -309 132 -308
rect 135 -309 174 -308
rect 212 -309 304 -308
rect 37 -311 188 -310
rect 212 -311 262 -310
rect 282 -311 304 -310
rect 37 -313 209 -312
rect 215 -313 234 -312
rect 240 -313 283 -312
rect 44 -315 104 -314
rect 107 -315 146 -314
rect 163 -315 185 -314
rect 208 -315 269 -314
rect 51 -317 139 -316
rect 142 -317 150 -316
rect 184 -317 255 -316
rect 58 -319 115 -318
rect 117 -319 325 -318
rect 79 -321 153 -320
rect 215 -321 332 -320
rect 86 -323 94 -322
rect 96 -323 297 -322
rect 324 -323 339 -322
rect 86 -325 122 -324
rect 128 -325 195 -324
rect 229 -325 318 -324
rect 100 -327 171 -326
rect 226 -327 318 -326
rect 110 -329 346 -328
rect 135 -331 248 -330
rect 142 -333 178 -332
rect 219 -333 248 -332
rect 121 -335 178 -334
rect 198 -335 220 -334
rect 243 -335 311 -334
rect 198 -337 276 -336
rect 296 -337 311 -336
rect 201 -339 276 -338
rect 2 -350 115 -349
rect 121 -350 136 -349
rect 145 -350 199 -349
rect 205 -350 318 -349
rect 16 -352 66 -351
rect 79 -352 90 -351
rect 93 -352 101 -351
rect 103 -352 164 -351
rect 173 -352 339 -351
rect 23 -354 108 -353
rect 145 -354 192 -353
rect 215 -354 241 -353
rect 243 -354 276 -353
rect 289 -354 318 -353
rect 30 -356 73 -355
rect 75 -356 80 -355
rect 86 -356 118 -355
rect 149 -356 167 -355
rect 177 -356 202 -355
rect 219 -356 332 -355
rect 9 -358 87 -357
rect 93 -358 192 -357
rect 226 -358 234 -357
rect 268 -358 297 -357
rect 299 -358 325 -357
rect 37 -360 136 -359
rect 152 -360 276 -359
rect 303 -360 346 -359
rect 37 -362 97 -361
rect 117 -362 283 -361
rect 44 -364 143 -363
rect 163 -364 290 -363
rect 44 -366 181 -365
rect 184 -366 325 -365
rect 51 -368 66 -367
rect 128 -368 220 -367
rect 233 -368 248 -367
rect 254 -368 269 -367
rect 58 -370 108 -369
rect 128 -370 213 -369
rect 247 -370 265 -369
rect 194 -372 255 -371
rect 261 -372 283 -371
rect 205 -374 213 -373
rect 9 -385 55 -384
rect 68 -385 297 -384
rect 306 -385 311 -384
rect 16 -387 62 -386
rect 75 -387 104 -386
rect 107 -387 118 -386
rect 128 -387 213 -386
rect 215 -387 332 -386
rect 23 -389 83 -388
rect 86 -389 115 -388
rect 128 -389 150 -388
rect 152 -389 199 -388
rect 205 -389 216 -388
rect 261 -389 318 -388
rect 2 -391 24 -390
rect 37 -391 76 -390
rect 93 -391 101 -390
rect 135 -391 143 -390
rect 156 -391 192 -390
rect 194 -391 283 -390
rect 285 -391 297 -390
rect 44 -393 90 -392
rect 96 -393 122 -392
rect 138 -393 192 -392
rect 201 -393 262 -392
rect 271 -393 318 -392
rect 44 -395 59 -394
rect 142 -395 150 -394
rect 163 -395 199 -394
rect 205 -395 244 -394
rect 282 -395 346 -394
rect 51 -397 66 -396
rect 166 -397 220 -396
rect 289 -397 304 -396
rect 40 -399 52 -398
rect 58 -399 80 -398
rect 170 -399 255 -398
rect 292 -399 311 -398
rect 79 -401 108 -400
rect 177 -401 325 -400
rect 177 -403 185 -402
rect 219 -403 227 -402
rect 240 -403 255 -402
rect 156 -405 227 -404
rect 180 -407 290 -406
rect 184 -409 248 -408
rect 247 -411 276 -410
rect 268 -413 276 -412
rect 268 -415 339 -414
rect 2 -426 132 -425
rect 135 -426 227 -425
rect 229 -426 241 -425
rect 254 -426 290 -425
rect 317 -426 328 -425
rect 9 -428 45 -427
rect 47 -428 52 -427
rect 54 -428 66 -427
rect 72 -428 97 -427
rect 114 -428 143 -427
rect 149 -428 164 -427
rect 170 -428 178 -427
rect 201 -428 234 -427
rect 268 -428 304 -427
rect 324 -428 339 -427
rect 16 -430 59 -429
rect 65 -430 94 -429
rect 107 -430 164 -429
rect 170 -430 185 -429
rect 205 -430 213 -429
rect 222 -430 318 -429
rect 23 -432 59 -431
rect 79 -432 94 -431
rect 107 -432 122 -431
rect 142 -432 157 -431
rect 184 -432 195 -431
rect 201 -432 206 -431
rect 226 -432 283 -431
rect 23 -434 136 -433
rect 233 -434 255 -433
rect 261 -434 304 -433
rect 30 -436 38 -435
rect 72 -436 283 -435
rect 30 -438 87 -437
rect 110 -438 178 -437
rect 219 -438 262 -437
rect 268 -438 297 -437
rect 37 -440 90 -439
rect 173 -440 220 -439
rect 82 -442 104 -441
rect 191 -442 297 -441
rect 191 -444 248 -443
rect 156 -446 248 -445
rect 2 -457 90 -456
rect 107 -457 139 -456
rect 170 -457 174 -456
rect 177 -457 192 -456
rect 198 -457 318 -456
rect 320 -457 353 -456
rect 359 -457 367 -456
rect 9 -459 45 -458
rect 75 -459 164 -458
rect 194 -459 318 -458
rect 331 -459 339 -458
rect 16 -461 80 -460
rect 93 -461 164 -460
rect 205 -461 213 -460
rect 215 -461 283 -460
rect 310 -461 335 -460
rect 23 -463 41 -462
rect 44 -463 132 -462
rect 135 -463 304 -462
rect 327 -463 339 -462
rect 30 -465 104 -464
rect 110 -465 297 -464
rect 37 -467 59 -466
rect 93 -467 143 -466
rect 184 -467 206 -466
rect 219 -467 304 -466
rect 51 -469 59 -468
rect 100 -469 178 -468
rect 180 -469 185 -468
rect 219 -469 297 -468
rect 51 -471 76 -470
rect 100 -471 146 -470
rect 233 -471 290 -470
rect 114 -473 160 -472
rect 233 -473 269 -472
rect 275 -473 290 -472
rect 114 -475 122 -474
rect 128 -475 223 -474
rect 247 -475 276 -474
rect 121 -477 150 -476
rect 215 -477 248 -476
rect 254 -477 311 -476
rect 86 -479 150 -478
rect 65 -481 87 -480
rect 128 -481 262 -480
rect 61 -483 66 -482
rect 138 -483 157 -482
rect 240 -483 262 -482
rect 142 -485 269 -484
rect 236 -487 241 -486
rect 16 -498 52 -497
rect 65 -498 83 -497
rect 103 -498 181 -497
rect 184 -498 258 -497
rect 282 -498 304 -497
rect 310 -498 325 -497
rect 331 -498 349 -497
rect 23 -500 80 -499
rect 114 -500 146 -499
rect 149 -500 185 -499
rect 198 -500 272 -499
rect 275 -500 311 -499
rect 320 -500 339 -499
rect 345 -500 360 -499
rect 30 -502 62 -501
rect 72 -502 87 -501
rect 93 -502 115 -501
rect 121 -502 150 -501
rect 177 -502 339 -501
rect 58 -504 66 -503
rect 72 -504 101 -503
rect 135 -504 195 -503
rect 201 -504 269 -503
rect 296 -504 332 -503
rect 44 -506 101 -505
rect 138 -506 164 -505
rect 180 -506 220 -505
rect 222 -506 318 -505
rect 44 -508 52 -507
rect 86 -508 157 -507
rect 163 -508 171 -507
rect 201 -508 227 -507
rect 229 -508 283 -507
rect 93 -510 129 -509
rect 142 -510 199 -509
rect 226 -510 276 -509
rect 82 -512 129 -511
rect 156 -512 206 -511
rect 233 -512 328 -511
rect 107 -514 171 -513
rect 247 -514 304 -513
rect 107 -516 167 -515
rect 191 -516 248 -515
rect 254 -516 290 -515
rect 124 -518 290 -517
rect 159 -520 234 -519
rect 261 -520 297 -519
rect 205 -522 262 -521
rect 212 -524 255 -523
rect 9 -535 34 -534
rect 37 -535 41 -534
rect 61 -535 94 -534
rect 100 -535 167 -534
rect 201 -535 206 -534
rect 208 -535 318 -534
rect 331 -535 346 -534
rect 352 -535 363 -534
rect 16 -537 83 -536
rect 86 -537 195 -536
rect 212 -537 311 -536
rect 331 -537 370 -536
rect 16 -539 83 -538
rect 93 -539 216 -538
rect 222 -539 304 -538
rect 23 -541 118 -540
rect 121 -541 136 -540
rect 138 -541 241 -540
rect 250 -541 304 -540
rect 23 -543 59 -542
rect 68 -543 87 -542
rect 114 -543 181 -542
rect 191 -543 318 -542
rect 30 -545 45 -544
rect 58 -545 104 -544
rect 124 -545 248 -544
rect 268 -545 311 -544
rect 135 -547 213 -546
rect 226 -547 244 -546
rect 247 -547 346 -546
rect 156 -549 255 -548
rect 261 -549 269 -548
rect 271 -549 325 -548
rect 107 -551 157 -550
rect 159 -551 171 -550
rect 177 -551 192 -550
rect 233 -551 262 -550
rect 324 -551 339 -550
rect 72 -553 108 -552
rect 163 -553 276 -552
rect 61 -555 73 -554
rect 163 -555 276 -554
rect 166 -557 199 -556
rect 233 -557 353 -556
rect 170 -559 185 -558
rect 254 -559 297 -558
rect 149 -561 185 -560
rect 289 -561 297 -560
rect 282 -563 290 -562
rect 219 -565 283 -564
rect 219 -567 339 -566
rect 9 -578 62 -577
rect 68 -578 80 -577
rect 93 -578 104 -577
rect 114 -578 213 -577
rect 219 -578 325 -577
rect 345 -578 370 -577
rect 23 -580 48 -579
rect 79 -580 111 -579
rect 114 -580 136 -579
rect 149 -580 185 -579
rect 212 -580 276 -579
rect 289 -580 360 -579
rect 44 -582 52 -581
rect 93 -582 122 -581
rect 128 -582 164 -581
rect 177 -582 332 -581
rect 44 -584 52 -583
rect 100 -584 129 -583
rect 135 -584 171 -583
rect 180 -584 283 -583
rect 16 -586 101 -585
rect 121 -586 146 -585
rect 149 -586 171 -585
rect 219 -586 227 -585
rect 229 -586 258 -585
rect 261 -586 276 -585
rect 152 -588 192 -587
rect 233 -588 311 -587
rect 156 -590 223 -589
rect 233 -590 262 -589
rect 264 -590 353 -589
rect 142 -592 157 -591
rect 163 -592 178 -591
rect 191 -592 199 -591
rect 236 -592 241 -591
rect 243 -592 304 -591
rect 310 -592 339 -591
rect 187 -594 199 -593
rect 240 -594 293 -593
rect 247 -596 297 -595
rect 250 -598 318 -597
rect 254 -600 283 -599
rect 254 -602 269 -601
rect 250 -604 269 -603
rect 65 -615 69 -614
rect 79 -615 108 -614
rect 110 -615 115 -614
rect 128 -615 164 -614
rect 187 -615 241 -614
rect 261 -615 269 -614
rect 289 -615 314 -614
rect 58 -617 69 -616
rect 86 -617 97 -616
rect 100 -617 122 -616
rect 128 -617 139 -616
rect 142 -617 171 -616
rect 194 -617 220 -616
rect 226 -617 251 -616
rect 268 -617 293 -616
rect 303 -617 311 -616
rect 86 -619 104 -618
rect 114 -619 136 -618
rect 142 -619 192 -618
rect 198 -619 255 -618
rect 275 -619 290 -618
rect 93 -621 125 -620
rect 156 -621 185 -620
rect 233 -621 241 -620
rect 257 -621 276 -620
rect 156 -623 209 -622
rect 233 -623 283 -622
rect 163 -625 213 -624
rect 282 -625 300 -624
rect 166 -627 220 -626
rect 170 -629 199 -628
rect 177 -631 213 -630
rect 177 -633 248 -632
rect 184 -635 206 -634
rect 44 -646 52 -645
rect 65 -646 83 -645
rect 96 -646 101 -645
rect 114 -646 153 -645
rect 156 -646 171 -645
rect 173 -646 241 -645
rect 243 -646 262 -645
rect 292 -646 304 -645
rect 44 -648 55 -647
rect 58 -648 66 -647
rect 72 -648 80 -647
rect 107 -648 115 -647
rect 121 -648 136 -647
rect 149 -648 220 -647
rect 247 -648 311 -647
rect 72 -650 87 -649
rect 93 -650 108 -649
rect 124 -650 164 -649
rect 180 -650 213 -649
rect 261 -650 283 -649
rect 79 -652 90 -651
rect 128 -652 143 -651
rect 184 -652 206 -651
rect 208 -652 276 -651
rect 142 -654 150 -653
rect 184 -654 223 -653
rect 268 -654 283 -653
rect 191 -656 199 -655
rect 201 -656 255 -655
rect 268 -656 279 -655
rect 191 -658 213 -657
rect 254 -658 265 -657
rect 194 -660 227 -659
rect 226 -662 241 -661
rect 44 -673 52 -672
rect 58 -673 66 -672
rect 72 -673 87 -672
rect 93 -673 101 -672
rect 103 -673 108 -672
rect 114 -673 129 -672
rect 135 -673 139 -672
rect 145 -673 150 -672
rect 170 -673 181 -672
rect 184 -673 202 -672
rect 212 -673 227 -672
rect 240 -673 248 -672
rect 268 -673 276 -672
rect 285 -673 293 -672
rect 58 -675 66 -674
rect 72 -675 97 -674
rect 121 -675 125 -674
rect 191 -675 220 -674
rect 226 -675 234 -674
rect 240 -675 244 -674
rect 191 -677 202 -676
rect 44 -688 52 -687
rect 58 -688 73 -687
rect 79 -688 87 -687
rect 93 -688 115 -687
rect 117 -688 122 -687
rect 135 -688 146 -687
rect 198 -688 206 -687
rect 212 -688 223 -687
rect 226 -688 244 -687
rect 254 -688 265 -687
rect 275 -688 286 -687
rect 107 -690 129 -689
rect 142 -690 153 -689
rect 233 -690 248 -689
<< m2contact >>
rect 135 0 136 1
rect 145 0 146 1
rect 142 -2 143 -1
rect 149 -2 150 -1
rect 100 -13 101 -12
rect 107 -13 108 -12
rect 121 -13 122 -12
rect 163 -13 164 -12
rect 177 -13 178 -12
rect 180 -13 181 -12
rect 128 -15 129 -14
rect 170 -15 171 -14
rect 177 -15 178 -14
rect 184 -15 185 -14
rect 135 -17 136 -16
rect 142 -17 143 -16
rect 149 -17 150 -16
rect 159 -17 160 -16
rect 135 -19 136 -18
rect 145 -19 146 -18
rect 152 -19 153 -18
rect 156 -19 157 -18
rect 79 -30 80 -29
rect 117 -30 118 -29
rect 128 -30 129 -29
rect 135 -30 136 -29
rect 142 -30 143 -29
rect 152 -30 153 -29
rect 159 -30 160 -29
rect 219 -30 220 -29
rect 86 -32 87 -31
rect 149 -32 150 -31
rect 170 -32 171 -31
rect 226 -32 227 -31
rect 93 -34 94 -33
rect 103 -34 104 -33
rect 121 -34 122 -33
rect 142 -34 143 -33
rect 170 -34 171 -33
rect 184 -34 185 -33
rect 191 -34 192 -33
rect 212 -34 213 -33
rect 100 -36 101 -35
rect 107 -36 108 -35
rect 135 -36 136 -35
rect 152 -36 153 -35
rect 163 -36 164 -35
rect 184 -36 185 -35
rect 194 -36 195 -35
rect 198 -36 199 -35
rect 156 -38 157 -37
rect 163 -38 164 -37
rect 180 -38 181 -37
rect 205 -38 206 -37
rect 79 -49 80 -48
rect 107 -49 108 -48
rect 114 -49 115 -48
rect 121 -49 122 -48
rect 128 -49 129 -48
rect 177 -49 178 -48
rect 180 -49 181 -48
rect 219 -49 220 -48
rect 222 -49 223 -48
rect 233 -49 234 -48
rect 79 -51 80 -50
rect 138 -51 139 -50
rect 145 -51 146 -50
rect 205 -51 206 -50
rect 86 -53 87 -52
rect 110 -53 111 -52
rect 114 -53 115 -52
rect 135 -53 136 -52
rect 145 -53 146 -52
rect 226 -53 227 -52
rect 86 -55 87 -54
rect 93 -55 94 -54
rect 100 -55 101 -54
rect 152 -55 153 -54
rect 156 -55 157 -54
rect 184 -55 185 -54
rect 191 -55 192 -54
rect 205 -55 206 -54
rect 93 -57 94 -56
rect 156 -57 157 -56
rect 170 -57 171 -56
rect 226 -57 227 -56
rect 131 -59 132 -58
rect 142 -59 143 -58
rect 149 -59 150 -58
rect 212 -59 213 -58
rect 110 -61 111 -60
rect 142 -61 143 -60
rect 163 -61 164 -60
rect 170 -61 171 -60
rect 187 -61 188 -60
rect 191 -61 192 -60
rect 198 -61 199 -60
rect 212 -61 213 -60
rect 149 -63 150 -62
rect 163 -63 164 -62
rect 72 -74 73 -73
rect 124 -74 125 -73
rect 135 -74 136 -73
rect 156 -74 157 -73
rect 159 -74 160 -73
rect 226 -74 227 -73
rect 243 -74 244 -73
rect 268 -74 269 -73
rect 79 -76 80 -75
rect 128 -76 129 -75
rect 138 -76 139 -75
rect 177 -76 178 -75
rect 184 -76 185 -75
rect 198 -76 199 -75
rect 205 -76 206 -75
rect 219 -76 220 -75
rect 222 -76 223 -75
rect 254 -76 255 -75
rect 261 -76 262 -75
rect 282 -76 283 -75
rect 79 -78 80 -77
rect 93 -78 94 -77
rect 121 -78 122 -77
rect 131 -78 132 -77
rect 138 -78 139 -77
rect 212 -78 213 -77
rect 86 -80 87 -79
rect 107 -80 108 -79
rect 142 -80 143 -79
rect 212 -80 213 -79
rect 65 -82 66 -81
rect 86 -82 87 -81
rect 93 -82 94 -81
rect 107 -82 108 -81
rect 152 -82 153 -81
rect 198 -82 199 -81
rect 205 -82 206 -81
rect 247 -82 248 -81
rect 100 -84 101 -83
rect 121 -84 122 -83
rect 156 -84 157 -83
rect 240 -84 241 -83
rect 100 -86 101 -85
rect 142 -86 143 -85
rect 163 -86 164 -85
rect 177 -86 178 -85
rect 191 -86 192 -85
rect 226 -86 227 -85
rect 114 -88 115 -87
rect 163 -88 164 -87
rect 114 -90 115 -89
rect 170 -90 171 -89
rect 170 -92 171 -91
rect 191 -92 192 -91
rect 44 -103 45 -102
rect 51 -103 52 -102
rect 65 -103 66 -102
rect 128 -103 129 -102
rect 142 -103 143 -102
rect 177 -103 178 -102
rect 198 -103 199 -102
rect 222 -103 223 -102
rect 254 -103 255 -102
rect 264 -103 265 -102
rect 268 -103 269 -102
rect 296 -103 297 -102
rect 299 -103 300 -102
rect 303 -103 304 -102
rect 65 -105 66 -104
rect 75 -105 76 -104
rect 79 -105 80 -104
rect 107 -105 108 -104
rect 131 -105 132 -104
rect 142 -105 143 -104
rect 149 -105 150 -104
rect 156 -105 157 -104
rect 159 -105 160 -104
rect 243 -105 244 -104
rect 247 -105 248 -104
rect 254 -105 255 -104
rect 282 -105 283 -104
rect 289 -105 290 -104
rect 72 -107 73 -106
rect 173 -107 174 -106
rect 205 -107 206 -106
rect 282 -107 283 -106
rect 86 -109 87 -108
rect 93 -109 94 -108
rect 100 -109 101 -108
rect 107 -109 108 -108
rect 117 -109 118 -108
rect 149 -109 150 -108
rect 152 -109 153 -108
rect 163 -109 164 -108
rect 170 -109 171 -108
rect 184 -109 185 -108
rect 212 -109 213 -108
rect 240 -109 241 -108
rect 93 -111 94 -110
rect 135 -111 136 -110
rect 138 -111 139 -110
rect 205 -111 206 -110
rect 212 -111 213 -110
rect 219 -111 220 -110
rect 226 -111 227 -110
rect 247 -111 248 -110
rect 100 -113 101 -112
rect 121 -113 122 -112
rect 156 -113 157 -112
rect 261 -113 262 -112
rect 114 -115 115 -114
rect 121 -115 122 -114
rect 163 -115 164 -114
rect 201 -115 202 -114
rect 219 -115 220 -114
rect 275 -115 276 -114
rect 58 -117 59 -116
rect 114 -117 115 -116
rect 177 -117 178 -116
rect 184 -117 185 -116
rect 191 -117 192 -116
rect 226 -117 227 -116
rect 19 -128 20 -127
rect 23 -128 24 -127
rect 30 -128 31 -127
rect 33 -128 34 -127
rect 47 -128 48 -127
rect 51 -128 52 -127
rect 58 -128 59 -127
rect 96 -128 97 -127
rect 100 -128 101 -127
rect 128 -128 129 -127
rect 135 -128 136 -127
rect 177 -128 178 -127
rect 184 -128 185 -127
rect 212 -128 213 -127
rect 240 -128 241 -127
rect 268 -128 269 -127
rect 289 -128 290 -127
rect 299 -128 300 -127
rect 310 -128 311 -127
rect 324 -128 325 -127
rect 331 -128 332 -127
rect 345 -128 346 -127
rect 58 -130 59 -129
rect 72 -130 73 -129
rect 79 -130 80 -129
rect 86 -130 87 -129
rect 107 -130 108 -129
rect 114 -130 115 -129
rect 149 -130 150 -129
rect 156 -130 157 -129
rect 159 -130 160 -129
rect 170 -130 171 -129
rect 177 -130 178 -129
rect 254 -130 255 -129
rect 271 -130 272 -129
rect 289 -130 290 -129
rect 296 -130 297 -129
rect 303 -130 304 -129
rect 324 -130 325 -129
rect 341 -130 342 -129
rect 65 -132 66 -131
rect 82 -132 83 -131
rect 93 -132 94 -131
rect 114 -132 115 -131
rect 121 -132 122 -131
rect 149 -132 150 -131
rect 156 -132 157 -131
rect 219 -132 220 -131
rect 254 -132 255 -131
rect 261 -132 262 -131
rect 275 -132 276 -131
rect 303 -132 304 -131
rect 37 -134 38 -133
rect 65 -134 66 -133
rect 68 -134 69 -133
rect 86 -134 87 -133
rect 93 -134 94 -133
rect 100 -134 101 -133
rect 107 -134 108 -133
rect 166 -134 167 -133
rect 191 -134 192 -133
rect 233 -134 234 -133
rect 236 -134 237 -133
rect 261 -134 262 -133
rect 79 -136 80 -135
rect 173 -136 174 -135
rect 198 -136 199 -135
rect 282 -136 283 -135
rect 121 -138 122 -137
rect 152 -138 153 -137
rect 163 -138 164 -137
rect 240 -138 241 -137
rect 247 -138 248 -137
rect 282 -138 283 -137
rect 163 -140 164 -139
rect 184 -140 185 -139
rect 201 -140 202 -139
rect 275 -140 276 -139
rect 170 -142 171 -141
rect 191 -142 192 -141
rect 205 -142 206 -141
rect 317 -142 318 -141
rect 194 -144 195 -143
rect 205 -144 206 -143
rect 226 -144 227 -143
rect 247 -144 248 -143
rect 131 -146 132 -145
rect 226 -146 227 -145
rect 19 -157 20 -156
rect 23 -157 24 -156
rect 37 -157 38 -156
rect 68 -157 69 -156
rect 72 -157 73 -156
rect 107 -157 108 -156
rect 114 -157 115 -156
rect 124 -157 125 -156
rect 152 -157 153 -156
rect 205 -157 206 -156
rect 212 -157 213 -156
rect 275 -157 276 -156
rect 296 -157 297 -156
rect 306 -157 307 -156
rect 310 -157 311 -156
rect 334 -157 335 -156
rect 345 -157 346 -156
rect 359 -157 360 -156
rect 44 -159 45 -158
rect 100 -159 101 -158
rect 107 -159 108 -158
rect 128 -159 129 -158
rect 163 -159 164 -158
rect 268 -159 269 -158
rect 296 -159 297 -158
rect 310 -159 311 -158
rect 51 -161 52 -160
rect 61 -161 62 -160
rect 79 -161 80 -160
rect 117 -161 118 -160
rect 128 -161 129 -160
rect 159 -161 160 -160
rect 163 -161 164 -160
rect 191 -161 192 -160
rect 201 -161 202 -160
rect 247 -161 248 -160
rect 303 -161 304 -160
rect 313 -161 314 -160
rect 51 -163 52 -162
rect 58 -163 59 -162
rect 86 -163 87 -162
rect 93 -163 94 -162
rect 114 -163 115 -162
rect 180 -163 181 -162
rect 184 -163 185 -162
rect 215 -163 216 -162
rect 219 -163 220 -162
rect 226 -163 227 -162
rect 303 -163 304 -162
rect 324 -163 325 -162
rect 58 -165 59 -164
rect 79 -165 80 -164
rect 86 -165 87 -164
rect 233 -165 234 -164
rect 313 -165 314 -164
rect 324 -165 325 -164
rect 93 -167 94 -166
rect 135 -167 136 -166
rect 149 -167 150 -166
rect 191 -167 192 -166
rect 198 -167 199 -166
rect 247 -167 248 -166
rect 135 -169 136 -168
rect 177 -169 178 -168
rect 180 -169 181 -168
rect 317 -169 318 -168
rect 142 -171 143 -170
rect 149 -171 150 -170
rect 156 -171 157 -170
rect 184 -171 185 -170
rect 198 -171 199 -170
rect 240 -171 241 -170
rect 268 -171 269 -170
rect 317 -171 318 -170
rect 166 -173 167 -172
rect 226 -173 227 -172
rect 233 -173 234 -172
rect 299 -173 300 -172
rect 173 -175 174 -174
rect 289 -175 290 -174
rect 121 -177 122 -176
rect 173 -177 174 -176
rect 205 -177 206 -176
rect 275 -177 276 -176
rect 100 -179 101 -178
rect 121 -179 122 -178
rect 254 -179 255 -178
rect 289 -179 290 -178
rect 254 -181 255 -180
rect 282 -181 283 -180
rect 261 -183 262 -182
rect 282 -183 283 -182
rect 212 -185 213 -184
rect 261 -185 262 -184
rect 30 -196 31 -195
rect 72 -196 73 -195
rect 79 -196 80 -195
rect 82 -196 83 -195
rect 86 -196 87 -195
rect 145 -196 146 -195
rect 159 -196 160 -195
rect 219 -196 220 -195
rect 229 -196 230 -195
rect 282 -196 283 -195
rect 296 -196 297 -195
rect 324 -196 325 -195
rect 331 -196 332 -195
rect 345 -196 346 -195
rect 359 -196 360 -195
rect 390 -196 391 -195
rect 37 -198 38 -197
rect 61 -198 62 -197
rect 72 -198 73 -197
rect 114 -198 115 -197
rect 121 -198 122 -197
rect 138 -198 139 -197
rect 159 -198 160 -197
rect 261 -198 262 -197
rect 296 -198 297 -197
rect 310 -198 311 -197
rect 352 -198 353 -197
rect 359 -198 360 -197
rect 373 -198 374 -197
rect 380 -198 381 -197
rect 40 -200 41 -199
rect 54 -200 55 -199
rect 58 -200 59 -199
rect 86 -200 87 -199
rect 100 -200 101 -199
rect 205 -200 206 -199
rect 212 -200 213 -199
rect 254 -200 255 -199
rect 303 -200 304 -199
rect 310 -200 311 -199
rect 352 -200 353 -199
rect 366 -200 367 -199
rect 44 -202 45 -201
rect 114 -202 115 -201
rect 135 -202 136 -201
rect 170 -202 171 -201
rect 180 -202 181 -201
rect 327 -202 328 -201
rect 44 -204 45 -203
rect 79 -204 80 -203
rect 103 -204 104 -203
rect 117 -204 118 -203
rect 135 -204 136 -203
rect 282 -204 283 -203
rect 303 -204 304 -203
rect 341 -204 342 -203
rect 51 -206 52 -205
rect 68 -206 69 -205
rect 107 -206 108 -205
rect 142 -206 143 -205
rect 163 -206 164 -205
rect 177 -206 178 -205
rect 187 -206 188 -205
rect 198 -206 199 -205
rect 215 -206 216 -205
rect 219 -206 220 -205
rect 240 -206 241 -205
rect 275 -206 276 -205
rect 65 -208 66 -207
rect 100 -208 101 -207
rect 128 -208 129 -207
rect 142 -208 143 -207
rect 149 -208 150 -207
rect 163 -208 164 -207
rect 184 -208 185 -207
rect 198 -208 199 -207
rect 233 -208 234 -207
rect 275 -208 276 -207
rect 107 -210 108 -209
rect 128 -210 129 -209
rect 149 -210 150 -209
rect 208 -210 209 -209
rect 243 -210 244 -209
rect 268 -210 269 -209
rect 215 -212 216 -211
rect 268 -212 269 -211
rect 247 -214 248 -213
rect 261 -214 262 -213
rect 240 -216 241 -215
rect 247 -216 248 -215
rect 254 -216 255 -215
rect 324 -216 325 -215
rect 9 -227 10 -226
rect 40 -227 41 -226
rect 54 -227 55 -226
rect 100 -227 101 -226
rect 107 -227 108 -226
rect 121 -227 122 -226
rect 128 -227 129 -226
rect 156 -227 157 -226
rect 177 -227 178 -226
rect 215 -227 216 -226
rect 222 -227 223 -226
rect 289 -227 290 -226
rect 310 -227 311 -226
rect 331 -227 332 -226
rect 334 -227 335 -226
rect 373 -227 374 -226
rect 387 -227 388 -226
rect 394 -227 395 -226
rect 16 -229 17 -228
rect 44 -229 45 -228
rect 79 -229 80 -228
rect 156 -229 157 -228
rect 159 -229 160 -228
rect 177 -229 178 -228
rect 212 -229 213 -228
rect 338 -229 339 -228
rect 345 -229 346 -228
rect 352 -229 353 -228
rect 355 -229 356 -228
rect 359 -229 360 -228
rect 23 -231 24 -230
rect 58 -231 59 -230
rect 93 -231 94 -230
rect 212 -231 213 -230
rect 233 -231 234 -230
rect 275 -231 276 -230
rect 282 -231 283 -230
rect 317 -231 318 -230
rect 327 -231 328 -230
rect 366 -231 367 -230
rect 30 -233 31 -232
rect 89 -233 90 -232
rect 93 -233 94 -232
rect 187 -233 188 -232
rect 226 -233 227 -232
rect 275 -233 276 -232
rect 289 -233 290 -232
rect 320 -233 321 -232
rect 33 -235 34 -234
rect 310 -235 311 -234
rect 37 -237 38 -236
rect 110 -237 111 -236
rect 114 -237 115 -236
rect 135 -237 136 -236
rect 149 -237 150 -236
rect 173 -237 174 -236
rect 198 -237 199 -236
rect 226 -237 227 -236
rect 233 -237 234 -236
rect 254 -237 255 -236
rect 268 -237 269 -236
rect 282 -237 283 -236
rect 303 -237 304 -236
rect 327 -237 328 -236
rect 51 -239 52 -238
rect 110 -239 111 -238
rect 114 -239 115 -238
rect 121 -239 122 -238
rect 135 -239 136 -238
rect 142 -239 143 -238
rect 149 -239 150 -238
rect 163 -239 164 -238
rect 191 -239 192 -238
rect 198 -239 199 -238
rect 205 -239 206 -238
rect 303 -239 304 -238
rect 58 -241 59 -240
rect 72 -241 73 -240
rect 152 -241 153 -240
rect 163 -241 164 -240
rect 170 -241 171 -240
rect 191 -241 192 -240
rect 208 -241 209 -240
rect 254 -241 255 -240
rect 44 -243 45 -242
rect 152 -243 153 -242
rect 170 -243 171 -242
rect 184 -243 185 -242
rect 240 -243 241 -242
rect 247 -243 248 -242
rect 250 -243 251 -242
rect 261 -243 262 -242
rect 72 -245 73 -244
rect 86 -245 87 -244
rect 219 -245 220 -244
rect 240 -245 241 -244
rect 261 -245 262 -244
rect 268 -245 269 -244
rect 9 -256 10 -255
rect 33 -256 34 -255
rect 37 -256 38 -255
rect 198 -256 199 -255
rect 205 -256 206 -255
rect 233 -256 234 -255
rect 268 -256 269 -255
rect 296 -256 297 -255
rect 345 -256 346 -255
rect 352 -256 353 -255
rect 387 -256 388 -255
rect 394 -256 395 -255
rect 9 -258 10 -257
rect 68 -258 69 -257
rect 72 -258 73 -257
rect 82 -258 83 -257
rect 89 -258 90 -257
rect 114 -258 115 -257
rect 128 -258 129 -257
rect 226 -258 227 -257
rect 16 -260 17 -259
rect 142 -260 143 -259
rect 145 -260 146 -259
rect 338 -260 339 -259
rect 16 -262 17 -261
rect 114 -262 115 -261
rect 135 -262 136 -261
rect 142 -262 143 -261
rect 149 -262 150 -261
rect 345 -262 346 -261
rect 23 -264 24 -263
rect 75 -264 76 -263
rect 79 -264 80 -263
rect 191 -264 192 -263
rect 208 -264 209 -263
rect 247 -264 248 -263
rect 23 -266 24 -265
rect 79 -266 80 -265
rect 93 -266 94 -265
rect 131 -266 132 -265
rect 149 -266 150 -265
rect 303 -266 304 -265
rect 51 -268 52 -267
rect 163 -268 164 -267
rect 173 -268 174 -267
rect 212 -268 213 -267
rect 215 -268 216 -267
rect 317 -268 318 -267
rect 54 -270 55 -269
rect 243 -270 244 -269
rect 289 -270 290 -269
rect 303 -270 304 -269
rect 310 -270 311 -269
rect 317 -270 318 -269
rect 58 -272 59 -271
rect 86 -272 87 -271
rect 100 -272 101 -271
rect 135 -272 136 -271
rect 156 -272 157 -271
rect 219 -272 220 -271
rect 226 -272 227 -271
rect 240 -272 241 -271
rect 254 -272 255 -271
rect 310 -272 311 -271
rect 58 -274 59 -273
rect 65 -274 66 -273
rect 72 -274 73 -273
rect 86 -274 87 -273
rect 100 -274 101 -273
rect 152 -274 153 -273
rect 159 -274 160 -273
rect 247 -274 248 -273
rect 254 -274 255 -273
rect 275 -274 276 -273
rect 2 -276 3 -275
rect 65 -276 66 -275
rect 107 -276 108 -275
rect 163 -276 164 -275
rect 170 -276 171 -275
rect 219 -276 220 -275
rect 233 -276 234 -275
rect 289 -276 290 -275
rect 107 -278 108 -277
rect 121 -278 122 -277
rect 170 -278 171 -277
rect 198 -278 199 -277
rect 212 -278 213 -277
rect 324 -278 325 -277
rect 121 -280 122 -279
rect 187 -280 188 -279
rect 191 -280 192 -279
rect 331 -280 332 -279
rect 156 -282 157 -281
rect 331 -282 332 -281
rect 177 -284 178 -283
rect 268 -284 269 -283
rect 44 -286 45 -285
rect 177 -286 178 -285
rect 180 -286 181 -285
rect 261 -286 262 -285
rect 44 -288 45 -287
rect 96 -288 97 -287
rect 184 -288 185 -287
rect 296 -288 297 -287
rect 194 -290 195 -289
rect 275 -290 276 -289
rect 222 -292 223 -291
rect 261 -292 262 -291
rect 2 -303 3 -302
rect 30 -303 31 -302
rect 44 -303 45 -302
rect 191 -303 192 -302
rect 205 -303 206 -302
rect 289 -303 290 -302
rect 16 -305 17 -304
rect 75 -305 76 -304
rect 79 -305 80 -304
rect 149 -305 150 -304
rect 170 -305 171 -304
rect 268 -305 269 -304
rect 23 -307 24 -306
rect 54 -307 55 -306
rect 65 -307 66 -306
rect 163 -307 164 -306
rect 187 -307 188 -306
rect 254 -307 255 -306
rect 261 -307 262 -306
rect 289 -307 290 -306
rect 30 -309 31 -308
rect 58 -309 59 -308
rect 65 -309 66 -308
rect 131 -309 132 -308
rect 135 -309 136 -308
rect 173 -309 174 -308
rect 212 -309 213 -308
rect 303 -309 304 -308
rect 37 -311 38 -310
rect 187 -311 188 -310
rect 212 -311 213 -310
rect 261 -311 262 -310
rect 282 -311 283 -310
rect 303 -311 304 -310
rect 37 -313 38 -312
rect 208 -313 209 -312
rect 215 -313 216 -312
rect 233 -313 234 -312
rect 240 -313 241 -312
rect 282 -313 283 -312
rect 44 -315 45 -314
rect 103 -315 104 -314
rect 107 -315 108 -314
rect 145 -315 146 -314
rect 163 -315 164 -314
rect 184 -315 185 -314
rect 208 -315 209 -314
rect 268 -315 269 -314
rect 51 -317 52 -316
rect 138 -317 139 -316
rect 142 -317 143 -316
rect 149 -317 150 -316
rect 184 -317 185 -316
rect 254 -317 255 -316
rect 58 -319 59 -318
rect 114 -319 115 -318
rect 117 -319 118 -318
rect 324 -319 325 -318
rect 79 -321 80 -320
rect 152 -321 153 -320
rect 215 -321 216 -320
rect 331 -321 332 -320
rect 86 -323 87 -322
rect 93 -323 94 -322
rect 96 -323 97 -322
rect 296 -323 297 -322
rect 324 -323 325 -322
rect 338 -323 339 -322
rect 86 -325 87 -324
rect 121 -325 122 -324
rect 128 -325 129 -324
rect 194 -325 195 -324
rect 229 -325 230 -324
rect 317 -325 318 -324
rect 100 -327 101 -326
rect 170 -327 171 -326
rect 226 -327 227 -326
rect 317 -327 318 -326
rect 110 -329 111 -328
rect 345 -329 346 -328
rect 135 -331 136 -330
rect 247 -331 248 -330
rect 142 -333 143 -332
rect 177 -333 178 -332
rect 219 -333 220 -332
rect 247 -333 248 -332
rect 121 -335 122 -334
rect 177 -335 178 -334
rect 198 -335 199 -334
rect 219 -335 220 -334
rect 243 -335 244 -334
rect 310 -335 311 -334
rect 198 -337 199 -336
rect 275 -337 276 -336
rect 296 -337 297 -336
rect 310 -337 311 -336
rect 201 -339 202 -338
rect 275 -339 276 -338
rect 2 -350 3 -349
rect 114 -350 115 -349
rect 121 -350 122 -349
rect 135 -350 136 -349
rect 145 -350 146 -349
rect 198 -350 199 -349
rect 205 -350 206 -349
rect 317 -350 318 -349
rect 16 -352 17 -351
rect 65 -352 66 -351
rect 79 -352 80 -351
rect 89 -352 90 -351
rect 93 -352 94 -351
rect 100 -352 101 -351
rect 103 -352 104 -351
rect 163 -352 164 -351
rect 173 -352 174 -351
rect 338 -352 339 -351
rect 23 -354 24 -353
rect 107 -354 108 -353
rect 145 -354 146 -353
rect 191 -354 192 -353
rect 215 -354 216 -353
rect 240 -354 241 -353
rect 243 -354 244 -353
rect 275 -354 276 -353
rect 289 -354 290 -353
rect 317 -354 318 -353
rect 30 -356 31 -355
rect 72 -356 73 -355
rect 75 -356 76 -355
rect 79 -356 80 -355
rect 86 -356 87 -355
rect 117 -356 118 -355
rect 149 -356 150 -355
rect 166 -356 167 -355
rect 177 -356 178 -355
rect 201 -356 202 -355
rect 219 -356 220 -355
rect 331 -356 332 -355
rect 9 -358 10 -357
rect 86 -358 87 -357
rect 93 -358 94 -357
rect 191 -358 192 -357
rect 226 -358 227 -357
rect 233 -358 234 -357
rect 268 -358 269 -357
rect 296 -358 297 -357
rect 299 -358 300 -357
rect 324 -358 325 -357
rect 37 -360 38 -359
rect 135 -360 136 -359
rect 152 -360 153 -359
rect 275 -360 276 -359
rect 303 -360 304 -359
rect 345 -360 346 -359
rect 37 -362 38 -361
rect 96 -362 97 -361
rect 117 -362 118 -361
rect 282 -362 283 -361
rect 44 -364 45 -363
rect 142 -364 143 -363
rect 163 -364 164 -363
rect 289 -364 290 -363
rect 44 -366 45 -365
rect 180 -366 181 -365
rect 184 -366 185 -365
rect 324 -366 325 -365
rect 51 -368 52 -367
rect 65 -368 66 -367
rect 128 -368 129 -367
rect 219 -368 220 -367
rect 233 -368 234 -367
rect 247 -368 248 -367
rect 254 -368 255 -367
rect 268 -368 269 -367
rect 58 -370 59 -369
rect 107 -370 108 -369
rect 128 -370 129 -369
rect 212 -370 213 -369
rect 247 -370 248 -369
rect 264 -370 265 -369
rect 194 -372 195 -371
rect 254 -372 255 -371
rect 261 -372 262 -371
rect 282 -372 283 -371
rect 205 -374 206 -373
rect 212 -374 213 -373
rect 9 -385 10 -384
rect 54 -385 55 -384
rect 68 -385 69 -384
rect 296 -385 297 -384
rect 306 -385 307 -384
rect 310 -385 311 -384
rect 16 -387 17 -386
rect 61 -387 62 -386
rect 75 -387 76 -386
rect 103 -387 104 -386
rect 107 -387 108 -386
rect 117 -387 118 -386
rect 128 -387 129 -386
rect 212 -387 213 -386
rect 215 -387 216 -386
rect 331 -387 332 -386
rect 23 -389 24 -388
rect 82 -389 83 -388
rect 86 -389 87 -388
rect 114 -389 115 -388
rect 128 -389 129 -388
rect 149 -389 150 -388
rect 152 -389 153 -388
rect 198 -389 199 -388
rect 205 -389 206 -388
rect 215 -389 216 -388
rect 261 -389 262 -388
rect 317 -389 318 -388
rect 2 -391 3 -390
rect 23 -391 24 -390
rect 37 -391 38 -390
rect 75 -391 76 -390
rect 93 -391 94 -390
rect 100 -391 101 -390
rect 135 -391 136 -390
rect 142 -391 143 -390
rect 156 -391 157 -390
rect 191 -391 192 -390
rect 194 -391 195 -390
rect 282 -391 283 -390
rect 285 -391 286 -390
rect 296 -391 297 -390
rect 44 -393 45 -392
rect 89 -393 90 -392
rect 96 -393 97 -392
rect 121 -393 122 -392
rect 138 -393 139 -392
rect 191 -393 192 -392
rect 201 -393 202 -392
rect 261 -393 262 -392
rect 271 -393 272 -392
rect 317 -393 318 -392
rect 44 -395 45 -394
rect 58 -395 59 -394
rect 142 -395 143 -394
rect 149 -395 150 -394
rect 163 -395 164 -394
rect 198 -395 199 -394
rect 205 -395 206 -394
rect 243 -395 244 -394
rect 282 -395 283 -394
rect 345 -395 346 -394
rect 51 -397 52 -396
rect 65 -397 66 -396
rect 166 -397 167 -396
rect 219 -397 220 -396
rect 289 -397 290 -396
rect 303 -397 304 -396
rect 40 -399 41 -398
rect 51 -399 52 -398
rect 58 -399 59 -398
rect 79 -399 80 -398
rect 170 -399 171 -398
rect 254 -399 255 -398
rect 292 -399 293 -398
rect 310 -399 311 -398
rect 79 -401 80 -400
rect 107 -401 108 -400
rect 177 -401 178 -400
rect 324 -401 325 -400
rect 177 -403 178 -402
rect 184 -403 185 -402
rect 219 -403 220 -402
rect 226 -403 227 -402
rect 240 -403 241 -402
rect 254 -403 255 -402
rect 156 -405 157 -404
rect 226 -405 227 -404
rect 180 -407 181 -406
rect 289 -407 290 -406
rect 184 -409 185 -408
rect 247 -409 248 -408
rect 247 -411 248 -410
rect 275 -411 276 -410
rect 268 -413 269 -412
rect 275 -413 276 -412
rect 268 -415 269 -414
rect 338 -415 339 -414
rect 2 -426 3 -425
rect 131 -426 132 -425
rect 135 -426 136 -425
rect 226 -426 227 -425
rect 229 -426 230 -425
rect 240 -426 241 -425
rect 254 -426 255 -425
rect 289 -426 290 -425
rect 317 -426 318 -425
rect 327 -426 328 -425
rect 9 -428 10 -427
rect 44 -428 45 -427
rect 47 -428 48 -427
rect 51 -428 52 -427
rect 54 -428 55 -427
rect 65 -428 66 -427
rect 72 -428 73 -427
rect 96 -428 97 -427
rect 114 -428 115 -427
rect 142 -428 143 -427
rect 149 -428 150 -427
rect 163 -428 164 -427
rect 170 -428 171 -427
rect 177 -428 178 -427
rect 201 -428 202 -427
rect 233 -428 234 -427
rect 268 -428 269 -427
rect 303 -428 304 -427
rect 324 -428 325 -427
rect 338 -428 339 -427
rect 16 -430 17 -429
rect 58 -430 59 -429
rect 65 -430 66 -429
rect 93 -430 94 -429
rect 107 -430 108 -429
rect 163 -430 164 -429
rect 170 -430 171 -429
rect 184 -430 185 -429
rect 205 -430 206 -429
rect 212 -430 213 -429
rect 222 -430 223 -429
rect 317 -430 318 -429
rect 23 -432 24 -431
rect 58 -432 59 -431
rect 79 -432 80 -431
rect 93 -432 94 -431
rect 107 -432 108 -431
rect 121 -432 122 -431
rect 142 -432 143 -431
rect 156 -432 157 -431
rect 184 -432 185 -431
rect 194 -432 195 -431
rect 201 -432 202 -431
rect 205 -432 206 -431
rect 226 -432 227 -431
rect 282 -432 283 -431
rect 23 -434 24 -433
rect 135 -434 136 -433
rect 233 -434 234 -433
rect 254 -434 255 -433
rect 261 -434 262 -433
rect 303 -434 304 -433
rect 30 -436 31 -435
rect 37 -436 38 -435
rect 72 -436 73 -435
rect 282 -436 283 -435
rect 30 -438 31 -437
rect 86 -438 87 -437
rect 110 -438 111 -437
rect 177 -438 178 -437
rect 219 -438 220 -437
rect 261 -438 262 -437
rect 268 -438 269 -437
rect 296 -438 297 -437
rect 37 -440 38 -439
rect 89 -440 90 -439
rect 173 -440 174 -439
rect 219 -440 220 -439
rect 82 -442 83 -441
rect 103 -442 104 -441
rect 191 -442 192 -441
rect 296 -442 297 -441
rect 191 -444 192 -443
rect 247 -444 248 -443
rect 156 -446 157 -445
rect 247 -446 248 -445
rect 2 -457 3 -456
rect 89 -457 90 -456
rect 107 -457 108 -456
rect 138 -457 139 -456
rect 170 -457 171 -456
rect 173 -457 174 -456
rect 177 -457 178 -456
rect 191 -457 192 -456
rect 198 -457 199 -456
rect 317 -457 318 -456
rect 320 -457 321 -456
rect 352 -457 353 -456
rect 359 -457 360 -456
rect 366 -457 367 -456
rect 9 -459 10 -458
rect 44 -459 45 -458
rect 75 -459 76 -458
rect 163 -459 164 -458
rect 194 -459 195 -458
rect 317 -459 318 -458
rect 331 -459 332 -458
rect 338 -459 339 -458
rect 16 -461 17 -460
rect 79 -461 80 -460
rect 93 -461 94 -460
rect 163 -461 164 -460
rect 205 -461 206 -460
rect 212 -461 213 -460
rect 215 -461 216 -460
rect 282 -461 283 -460
rect 310 -461 311 -460
rect 334 -461 335 -460
rect 23 -463 24 -462
rect 40 -463 41 -462
rect 44 -463 45 -462
rect 131 -463 132 -462
rect 135 -463 136 -462
rect 303 -463 304 -462
rect 327 -463 328 -462
rect 338 -463 339 -462
rect 30 -465 31 -464
rect 103 -465 104 -464
rect 110 -465 111 -464
rect 296 -465 297 -464
rect 37 -467 38 -466
rect 58 -467 59 -466
rect 93 -467 94 -466
rect 142 -467 143 -466
rect 184 -467 185 -466
rect 205 -467 206 -466
rect 219 -467 220 -466
rect 303 -467 304 -466
rect 51 -469 52 -468
rect 58 -469 59 -468
rect 100 -469 101 -468
rect 177 -469 178 -468
rect 180 -469 181 -468
rect 184 -469 185 -468
rect 219 -469 220 -468
rect 296 -469 297 -468
rect 51 -471 52 -470
rect 75 -471 76 -470
rect 100 -471 101 -470
rect 145 -471 146 -470
rect 233 -471 234 -470
rect 289 -471 290 -470
rect 114 -473 115 -472
rect 159 -473 160 -472
rect 233 -473 234 -472
rect 268 -473 269 -472
rect 275 -473 276 -472
rect 289 -473 290 -472
rect 114 -475 115 -474
rect 121 -475 122 -474
rect 128 -475 129 -474
rect 222 -475 223 -474
rect 247 -475 248 -474
rect 275 -475 276 -474
rect 121 -477 122 -476
rect 149 -477 150 -476
rect 215 -477 216 -476
rect 247 -477 248 -476
rect 254 -477 255 -476
rect 310 -477 311 -476
rect 86 -479 87 -478
rect 149 -479 150 -478
rect 65 -481 66 -480
rect 86 -481 87 -480
rect 128 -481 129 -480
rect 261 -481 262 -480
rect 61 -483 62 -482
rect 65 -483 66 -482
rect 138 -483 139 -482
rect 156 -483 157 -482
rect 240 -483 241 -482
rect 261 -483 262 -482
rect 142 -485 143 -484
rect 268 -485 269 -484
rect 236 -487 237 -486
rect 240 -487 241 -486
rect 16 -498 17 -497
rect 51 -498 52 -497
rect 65 -498 66 -497
rect 82 -498 83 -497
rect 103 -498 104 -497
rect 180 -498 181 -497
rect 184 -498 185 -497
rect 257 -498 258 -497
rect 282 -498 283 -497
rect 303 -498 304 -497
rect 310 -498 311 -497
rect 324 -498 325 -497
rect 331 -498 332 -497
rect 348 -498 349 -497
rect 23 -500 24 -499
rect 79 -500 80 -499
rect 114 -500 115 -499
rect 145 -500 146 -499
rect 149 -500 150 -499
rect 184 -500 185 -499
rect 198 -500 199 -499
rect 271 -500 272 -499
rect 275 -500 276 -499
rect 310 -500 311 -499
rect 320 -500 321 -499
rect 338 -500 339 -499
rect 345 -500 346 -499
rect 359 -500 360 -499
rect 30 -502 31 -501
rect 61 -502 62 -501
rect 72 -502 73 -501
rect 86 -502 87 -501
rect 93 -502 94 -501
rect 114 -502 115 -501
rect 121 -502 122 -501
rect 149 -502 150 -501
rect 177 -502 178 -501
rect 338 -502 339 -501
rect 58 -504 59 -503
rect 65 -504 66 -503
rect 72 -504 73 -503
rect 100 -504 101 -503
rect 135 -504 136 -503
rect 194 -504 195 -503
rect 201 -504 202 -503
rect 268 -504 269 -503
rect 296 -504 297 -503
rect 331 -504 332 -503
rect 44 -506 45 -505
rect 100 -506 101 -505
rect 138 -506 139 -505
rect 163 -506 164 -505
rect 180 -506 181 -505
rect 219 -506 220 -505
rect 222 -506 223 -505
rect 317 -506 318 -505
rect 44 -508 45 -507
rect 51 -508 52 -507
rect 86 -508 87 -507
rect 156 -508 157 -507
rect 163 -508 164 -507
rect 170 -508 171 -507
rect 201 -508 202 -507
rect 226 -508 227 -507
rect 229 -508 230 -507
rect 282 -508 283 -507
rect 93 -510 94 -509
rect 128 -510 129 -509
rect 142 -510 143 -509
rect 198 -510 199 -509
rect 226 -510 227 -509
rect 275 -510 276 -509
rect 82 -512 83 -511
rect 128 -512 129 -511
rect 156 -512 157 -511
rect 205 -512 206 -511
rect 233 -512 234 -511
rect 327 -512 328 -511
rect 107 -514 108 -513
rect 170 -514 171 -513
rect 247 -514 248 -513
rect 303 -514 304 -513
rect 107 -516 108 -515
rect 166 -516 167 -515
rect 191 -516 192 -515
rect 247 -516 248 -515
rect 254 -516 255 -515
rect 289 -516 290 -515
rect 124 -518 125 -517
rect 289 -518 290 -517
rect 159 -520 160 -519
rect 233 -520 234 -519
rect 261 -520 262 -519
rect 296 -520 297 -519
rect 205 -522 206 -521
rect 261 -522 262 -521
rect 212 -524 213 -523
rect 254 -524 255 -523
rect 9 -535 10 -534
rect 33 -535 34 -534
rect 37 -535 38 -534
rect 40 -535 41 -534
rect 61 -535 62 -534
rect 93 -535 94 -534
rect 100 -535 101 -534
rect 166 -535 167 -534
rect 201 -535 202 -534
rect 205 -535 206 -534
rect 208 -535 209 -534
rect 317 -535 318 -534
rect 331 -535 332 -534
rect 345 -535 346 -534
rect 352 -535 353 -534
rect 362 -535 363 -534
rect 16 -537 17 -536
rect 82 -537 83 -536
rect 86 -537 87 -536
rect 194 -537 195 -536
rect 212 -537 213 -536
rect 310 -537 311 -536
rect 331 -537 332 -536
rect 369 -537 370 -536
rect 16 -539 17 -538
rect 82 -539 83 -538
rect 93 -539 94 -538
rect 215 -539 216 -538
rect 222 -539 223 -538
rect 303 -539 304 -538
rect 23 -541 24 -540
rect 117 -541 118 -540
rect 121 -541 122 -540
rect 135 -541 136 -540
rect 138 -541 139 -540
rect 240 -541 241 -540
rect 250 -541 251 -540
rect 303 -541 304 -540
rect 23 -543 24 -542
rect 58 -543 59 -542
rect 68 -543 69 -542
rect 86 -543 87 -542
rect 114 -543 115 -542
rect 180 -543 181 -542
rect 191 -543 192 -542
rect 317 -543 318 -542
rect 30 -545 31 -544
rect 44 -545 45 -544
rect 58 -545 59 -544
rect 103 -545 104 -544
rect 124 -545 125 -544
rect 247 -545 248 -544
rect 268 -545 269 -544
rect 310 -545 311 -544
rect 135 -547 136 -546
rect 212 -547 213 -546
rect 226 -547 227 -546
rect 243 -547 244 -546
rect 247 -547 248 -546
rect 345 -547 346 -546
rect 156 -549 157 -548
rect 254 -549 255 -548
rect 261 -549 262 -548
rect 268 -549 269 -548
rect 271 -549 272 -548
rect 324 -549 325 -548
rect 107 -551 108 -550
rect 156 -551 157 -550
rect 159 -551 160 -550
rect 170 -551 171 -550
rect 177 -551 178 -550
rect 191 -551 192 -550
rect 233 -551 234 -550
rect 261 -551 262 -550
rect 324 -551 325 -550
rect 338 -551 339 -550
rect 72 -553 73 -552
rect 107 -553 108 -552
rect 163 -553 164 -552
rect 275 -553 276 -552
rect 61 -555 62 -554
rect 72 -555 73 -554
rect 163 -555 164 -554
rect 275 -555 276 -554
rect 166 -557 167 -556
rect 198 -557 199 -556
rect 233 -557 234 -556
rect 352 -557 353 -556
rect 170 -559 171 -558
rect 184 -559 185 -558
rect 254 -559 255 -558
rect 296 -559 297 -558
rect 149 -561 150 -560
rect 184 -561 185 -560
rect 289 -561 290 -560
rect 296 -561 297 -560
rect 282 -563 283 -562
rect 289 -563 290 -562
rect 219 -565 220 -564
rect 282 -565 283 -564
rect 219 -567 220 -566
rect 338 -567 339 -566
rect 9 -578 10 -577
rect 61 -578 62 -577
rect 68 -578 69 -577
rect 79 -578 80 -577
rect 93 -578 94 -577
rect 103 -578 104 -577
rect 114 -578 115 -577
rect 212 -578 213 -577
rect 219 -578 220 -577
rect 324 -578 325 -577
rect 345 -578 346 -577
rect 369 -578 370 -577
rect 23 -580 24 -579
rect 47 -580 48 -579
rect 79 -580 80 -579
rect 110 -580 111 -579
rect 114 -580 115 -579
rect 135 -580 136 -579
rect 149 -580 150 -579
rect 184 -580 185 -579
rect 212 -580 213 -579
rect 275 -580 276 -579
rect 289 -580 290 -579
rect 359 -580 360 -579
rect 44 -582 45 -581
rect 51 -582 52 -581
rect 93 -582 94 -581
rect 121 -582 122 -581
rect 128 -582 129 -581
rect 163 -582 164 -581
rect 177 -582 178 -581
rect 331 -582 332 -581
rect 44 -584 45 -583
rect 51 -584 52 -583
rect 100 -584 101 -583
rect 128 -584 129 -583
rect 135 -584 136 -583
rect 170 -584 171 -583
rect 180 -584 181 -583
rect 282 -584 283 -583
rect 16 -586 17 -585
rect 100 -586 101 -585
rect 121 -586 122 -585
rect 145 -586 146 -585
rect 149 -586 150 -585
rect 170 -586 171 -585
rect 219 -586 220 -585
rect 226 -586 227 -585
rect 229 -586 230 -585
rect 257 -586 258 -585
rect 261 -586 262 -585
rect 275 -586 276 -585
rect 152 -588 153 -587
rect 191 -588 192 -587
rect 233 -588 234 -587
rect 310 -588 311 -587
rect 156 -590 157 -589
rect 222 -590 223 -589
rect 233 -590 234 -589
rect 261 -590 262 -589
rect 264 -590 265 -589
rect 352 -590 353 -589
rect 142 -592 143 -591
rect 156 -592 157 -591
rect 163 -592 164 -591
rect 177 -592 178 -591
rect 191 -592 192 -591
rect 198 -592 199 -591
rect 236 -592 237 -591
rect 240 -592 241 -591
rect 243 -592 244 -591
rect 303 -592 304 -591
rect 310 -592 311 -591
rect 338 -592 339 -591
rect 187 -594 188 -593
rect 198 -594 199 -593
rect 240 -594 241 -593
rect 292 -594 293 -593
rect 247 -596 248 -595
rect 296 -596 297 -595
rect 250 -598 251 -597
rect 317 -598 318 -597
rect 254 -600 255 -599
rect 282 -600 283 -599
rect 254 -602 255 -601
rect 268 -602 269 -601
rect 250 -604 251 -603
rect 268 -604 269 -603
rect 65 -615 66 -614
rect 68 -615 69 -614
rect 79 -615 80 -614
rect 107 -615 108 -614
rect 110 -615 111 -614
rect 114 -615 115 -614
rect 128 -615 129 -614
rect 163 -615 164 -614
rect 187 -615 188 -614
rect 240 -615 241 -614
rect 261 -615 262 -614
rect 268 -615 269 -614
rect 289 -615 290 -614
rect 313 -615 314 -614
rect 58 -617 59 -616
rect 68 -617 69 -616
rect 86 -617 87 -616
rect 96 -617 97 -616
rect 100 -617 101 -616
rect 121 -617 122 -616
rect 128 -617 129 -616
rect 138 -617 139 -616
rect 142 -617 143 -616
rect 170 -617 171 -616
rect 194 -617 195 -616
rect 219 -617 220 -616
rect 226 -617 227 -616
rect 250 -617 251 -616
rect 268 -617 269 -616
rect 292 -617 293 -616
rect 303 -617 304 -616
rect 310 -617 311 -616
rect 86 -619 87 -618
rect 103 -619 104 -618
rect 114 -619 115 -618
rect 135 -619 136 -618
rect 142 -619 143 -618
rect 191 -619 192 -618
rect 198 -619 199 -618
rect 254 -619 255 -618
rect 275 -619 276 -618
rect 289 -619 290 -618
rect 93 -621 94 -620
rect 124 -621 125 -620
rect 156 -621 157 -620
rect 184 -621 185 -620
rect 233 -621 234 -620
rect 240 -621 241 -620
rect 257 -621 258 -620
rect 275 -621 276 -620
rect 156 -623 157 -622
rect 208 -623 209 -622
rect 233 -623 234 -622
rect 282 -623 283 -622
rect 163 -625 164 -624
rect 212 -625 213 -624
rect 282 -625 283 -624
rect 299 -625 300 -624
rect 166 -627 167 -626
rect 219 -627 220 -626
rect 170 -629 171 -628
rect 198 -629 199 -628
rect 177 -631 178 -630
rect 212 -631 213 -630
rect 177 -633 178 -632
rect 247 -633 248 -632
rect 184 -635 185 -634
rect 205 -635 206 -634
rect 44 -646 45 -645
rect 51 -646 52 -645
rect 65 -646 66 -645
rect 82 -646 83 -645
rect 96 -646 97 -645
rect 100 -646 101 -645
rect 114 -646 115 -645
rect 152 -646 153 -645
rect 156 -646 157 -645
rect 170 -646 171 -645
rect 173 -646 174 -645
rect 240 -646 241 -645
rect 243 -646 244 -645
rect 261 -646 262 -645
rect 292 -646 293 -645
rect 303 -646 304 -645
rect 44 -648 45 -647
rect 54 -648 55 -647
rect 58 -648 59 -647
rect 65 -648 66 -647
rect 72 -648 73 -647
rect 79 -648 80 -647
rect 107 -648 108 -647
rect 114 -648 115 -647
rect 121 -648 122 -647
rect 135 -648 136 -647
rect 149 -648 150 -647
rect 219 -648 220 -647
rect 247 -648 248 -647
rect 310 -648 311 -647
rect 72 -650 73 -649
rect 86 -650 87 -649
rect 93 -650 94 -649
rect 107 -650 108 -649
rect 124 -650 125 -649
rect 163 -650 164 -649
rect 180 -650 181 -649
rect 212 -650 213 -649
rect 261 -650 262 -649
rect 282 -650 283 -649
rect 79 -652 80 -651
rect 89 -652 90 -651
rect 128 -652 129 -651
rect 142 -652 143 -651
rect 184 -652 185 -651
rect 205 -652 206 -651
rect 208 -652 209 -651
rect 275 -652 276 -651
rect 142 -654 143 -653
rect 149 -654 150 -653
rect 184 -654 185 -653
rect 222 -654 223 -653
rect 268 -654 269 -653
rect 282 -654 283 -653
rect 191 -656 192 -655
rect 198 -656 199 -655
rect 201 -656 202 -655
rect 254 -656 255 -655
rect 268 -656 269 -655
rect 278 -656 279 -655
rect 191 -658 192 -657
rect 212 -658 213 -657
rect 254 -658 255 -657
rect 264 -658 265 -657
rect 194 -660 195 -659
rect 226 -660 227 -659
rect 226 -662 227 -661
rect 240 -662 241 -661
rect 44 -673 45 -672
rect 51 -673 52 -672
rect 58 -673 59 -672
rect 65 -673 66 -672
rect 72 -673 73 -672
rect 86 -673 87 -672
rect 93 -673 94 -672
rect 100 -673 101 -672
rect 103 -673 104 -672
rect 107 -673 108 -672
rect 114 -673 115 -672
rect 128 -673 129 -672
rect 135 -673 136 -672
rect 138 -673 139 -672
rect 145 -673 146 -672
rect 149 -673 150 -672
rect 170 -673 171 -672
rect 180 -673 181 -672
rect 184 -673 185 -672
rect 201 -673 202 -672
rect 212 -673 213 -672
rect 226 -673 227 -672
rect 240 -673 241 -672
rect 247 -673 248 -672
rect 268 -673 269 -672
rect 275 -673 276 -672
rect 285 -673 286 -672
rect 292 -673 293 -672
rect 58 -675 59 -674
rect 65 -675 66 -674
rect 72 -675 73 -674
rect 96 -675 97 -674
rect 121 -675 122 -674
rect 124 -675 125 -674
rect 191 -675 192 -674
rect 219 -675 220 -674
rect 226 -675 227 -674
rect 233 -675 234 -674
rect 240 -675 241 -674
rect 243 -675 244 -674
rect 191 -677 192 -676
rect 201 -677 202 -676
rect 44 -688 45 -687
rect 51 -688 52 -687
rect 58 -688 59 -687
rect 72 -688 73 -687
rect 79 -688 80 -687
rect 86 -688 87 -687
rect 93 -688 94 -687
rect 114 -688 115 -687
rect 117 -688 118 -687
rect 121 -688 122 -687
rect 135 -688 136 -687
rect 145 -688 146 -687
rect 198 -688 199 -687
rect 205 -688 206 -687
rect 212 -688 213 -687
rect 222 -688 223 -687
rect 226 -688 227 -687
rect 243 -688 244 -687
rect 254 -688 255 -687
rect 264 -688 265 -687
rect 275 -688 276 -687
rect 285 -688 286 -687
rect 107 -690 108 -689
rect 128 -690 129 -689
rect 142 -690 143 -689
rect 152 -690 153 -689
rect 233 -690 234 -689
rect 247 -690 248 -689
<< metal2 >>
rect 135 -3 136 1
rect 145 -3 146 1
rect 142 -3 143 -1
rect 149 -3 150 -1
rect 100 -20 101 -12
rect 107 -20 108 -12
rect 121 -20 122 -12
rect 163 -20 164 -12
rect 177 -13 178 -11
rect 180 -20 181 -12
rect 128 -20 129 -14
rect 170 -20 171 -14
rect 177 -20 178 -14
rect 184 -20 185 -14
rect 135 -17 136 -11
rect 142 -20 143 -16
rect 149 -17 150 -11
rect 159 -17 160 -11
rect 135 -20 136 -18
rect 145 -20 146 -18
rect 152 -20 153 -18
rect 156 -20 157 -18
rect 79 -39 80 -29
rect 117 -39 118 -29
rect 128 -39 129 -29
rect 135 -30 136 -28
rect 142 -30 143 -28
rect 152 -30 153 -28
rect 159 -39 160 -29
rect 219 -39 220 -29
rect 86 -39 87 -31
rect 149 -39 150 -31
rect 170 -32 171 -28
rect 226 -39 227 -31
rect 93 -39 94 -33
rect 103 -39 104 -33
rect 121 -39 122 -33
rect 142 -39 143 -33
rect 170 -39 171 -33
rect 184 -34 185 -28
rect 191 -34 192 -28
rect 212 -39 213 -33
rect 100 -39 101 -35
rect 107 -36 108 -28
rect 135 -39 136 -35
rect 152 -39 153 -35
rect 163 -36 164 -28
rect 184 -39 185 -35
rect 194 -39 195 -35
rect 198 -39 199 -35
rect 156 -38 157 -28
rect 163 -39 164 -37
rect 180 -39 181 -37
rect 205 -39 206 -37
rect 79 -49 80 -47
rect 107 -49 108 -47
rect 114 -49 115 -47
rect 121 -49 122 -47
rect 128 -49 129 -47
rect 177 -64 178 -48
rect 180 -49 181 -47
rect 219 -49 220 -47
rect 222 -64 223 -48
rect 233 -64 234 -48
rect 79 -64 80 -50
rect 138 -64 139 -50
rect 145 -51 146 -47
rect 205 -51 206 -47
rect 86 -53 87 -47
rect 110 -53 111 -47
rect 114 -64 115 -52
rect 135 -53 136 -47
rect 145 -64 146 -52
rect 226 -53 227 -47
rect 86 -64 87 -54
rect 93 -55 94 -47
rect 100 -64 101 -54
rect 152 -64 153 -54
rect 156 -55 157 -47
rect 184 -55 185 -47
rect 191 -55 192 -47
rect 205 -64 206 -54
rect 93 -64 94 -56
rect 156 -64 157 -56
rect 170 -57 171 -47
rect 226 -64 227 -56
rect 131 -64 132 -58
rect 142 -59 143 -47
rect 149 -59 150 -47
rect 212 -59 213 -47
rect 110 -64 111 -60
rect 142 -64 143 -60
rect 163 -61 164 -47
rect 170 -64 171 -60
rect 187 -64 188 -60
rect 191 -64 192 -60
rect 198 -61 199 -47
rect 212 -64 213 -60
rect 149 -64 150 -62
rect 163 -64 164 -62
rect 72 -93 73 -73
rect 124 -74 125 -72
rect 135 -74 136 -72
rect 156 -74 157 -72
rect 159 -74 160 -72
rect 226 -74 227 -72
rect 233 -74 234 -72
rect 233 -93 234 -73
rect 233 -74 234 -72
rect 233 -93 234 -73
rect 243 -93 244 -73
rect 268 -93 269 -73
rect 79 -76 80 -72
rect 128 -93 129 -75
rect 138 -76 139 -72
rect 177 -76 178 -72
rect 184 -93 185 -75
rect 198 -76 199 -72
rect 205 -76 206 -72
rect 219 -93 220 -75
rect 222 -93 223 -75
rect 254 -93 255 -75
rect 261 -93 262 -75
rect 282 -93 283 -75
rect 79 -93 80 -77
rect 93 -78 94 -72
rect 121 -78 122 -72
rect 131 -78 132 -72
rect 138 -93 139 -77
rect 212 -78 213 -72
rect 86 -80 87 -72
rect 107 -80 108 -72
rect 142 -80 143 -72
rect 212 -93 213 -79
rect 65 -93 66 -81
rect 86 -93 87 -81
rect 93 -93 94 -81
rect 107 -93 108 -81
rect 152 -93 153 -81
rect 198 -93 199 -81
rect 205 -93 206 -81
rect 247 -93 248 -81
rect 100 -84 101 -72
rect 121 -93 122 -83
rect 156 -93 157 -83
rect 240 -93 241 -83
rect 100 -93 101 -85
rect 142 -93 143 -85
rect 163 -86 164 -72
rect 177 -93 178 -85
rect 191 -86 192 -72
rect 226 -93 227 -85
rect 114 -88 115 -72
rect 163 -93 164 -87
rect 114 -93 115 -89
rect 170 -90 171 -72
rect 170 -93 171 -91
rect 191 -93 192 -91
rect 44 -118 45 -102
rect 51 -118 52 -102
rect 65 -103 66 -101
rect 128 -118 129 -102
rect 142 -103 143 -101
rect 177 -103 178 -101
rect 198 -103 199 -101
rect 222 -118 223 -102
rect 233 -103 234 -101
rect 233 -118 234 -102
rect 233 -103 234 -101
rect 233 -118 234 -102
rect 254 -103 255 -101
rect 264 -103 265 -101
rect 268 -103 269 -101
rect 296 -118 297 -102
rect 299 -118 300 -102
rect 303 -118 304 -102
rect 65 -118 66 -104
rect 75 -118 76 -104
rect 79 -105 80 -101
rect 107 -105 108 -101
rect 131 -105 132 -101
rect 142 -118 143 -104
rect 149 -105 150 -101
rect 156 -105 157 -101
rect 159 -118 160 -104
rect 243 -105 244 -101
rect 247 -105 248 -101
rect 254 -118 255 -104
rect 282 -105 283 -101
rect 289 -118 290 -104
rect 72 -107 73 -101
rect 173 -107 174 -101
rect 205 -107 206 -101
rect 282 -118 283 -106
rect 86 -118 87 -108
rect 93 -109 94 -101
rect 100 -109 101 -101
rect 107 -118 108 -108
rect 117 -118 118 -108
rect 149 -118 150 -108
rect 152 -109 153 -101
rect 163 -109 164 -101
rect 170 -118 171 -108
rect 184 -109 185 -101
rect 212 -109 213 -101
rect 240 -118 241 -108
rect 93 -118 94 -110
rect 135 -111 136 -101
rect 138 -118 139 -110
rect 205 -118 206 -110
rect 212 -118 213 -110
rect 219 -111 220 -101
rect 226 -111 227 -101
rect 247 -118 248 -110
rect 100 -118 101 -112
rect 121 -113 122 -101
rect 156 -118 157 -112
rect 261 -118 262 -112
rect 114 -115 115 -101
rect 121 -118 122 -114
rect 163 -118 164 -114
rect 201 -118 202 -114
rect 219 -118 220 -114
rect 275 -118 276 -114
rect 58 -118 59 -116
rect 114 -118 115 -116
rect 177 -118 178 -116
rect 184 -118 185 -116
rect 191 -117 192 -101
rect 226 -118 227 -116
rect 19 -147 20 -127
rect 23 -147 24 -127
rect 30 -147 31 -127
rect 33 -128 34 -126
rect 47 -147 48 -127
rect 51 -128 52 -126
rect 58 -128 59 -126
rect 96 -147 97 -127
rect 100 -128 101 -126
rect 128 -128 129 -126
rect 135 -147 136 -127
rect 177 -128 178 -126
rect 184 -128 185 -126
rect 212 -128 213 -126
rect 240 -128 241 -126
rect 268 -147 269 -127
rect 289 -128 290 -126
rect 299 -128 300 -126
rect 310 -147 311 -127
rect 324 -128 325 -126
rect 331 -147 332 -127
rect 345 -147 346 -127
rect 58 -147 59 -129
rect 72 -147 73 -129
rect 79 -130 80 -126
rect 86 -130 87 -126
rect 107 -130 108 -126
rect 114 -130 115 -126
rect 142 -130 143 -126
rect 142 -147 143 -129
rect 142 -130 143 -126
rect 142 -147 143 -129
rect 149 -130 150 -126
rect 156 -130 157 -126
rect 159 -130 160 -126
rect 170 -130 171 -126
rect 177 -147 178 -129
rect 254 -130 255 -126
rect 271 -130 272 -126
rect 289 -147 290 -129
rect 296 -147 297 -129
rect 303 -130 304 -126
rect 324 -147 325 -129
rect 341 -147 342 -129
rect 65 -132 66 -126
rect 82 -132 83 -126
rect 93 -132 94 -126
rect 114 -147 115 -131
rect 121 -132 122 -126
rect 149 -147 150 -131
rect 156 -147 157 -131
rect 219 -147 220 -131
rect 254 -147 255 -131
rect 261 -132 262 -126
rect 275 -132 276 -126
rect 303 -147 304 -131
rect 37 -147 38 -133
rect 65 -147 66 -133
rect 68 -147 69 -133
rect 86 -147 87 -133
rect 93 -147 94 -133
rect 100 -147 101 -133
rect 107 -147 108 -133
rect 166 -147 167 -133
rect 191 -134 192 -126
rect 233 -134 234 -126
rect 236 -147 237 -133
rect 261 -147 262 -133
rect 79 -147 80 -135
rect 173 -147 174 -135
rect 198 -136 199 -126
rect 282 -136 283 -126
rect 121 -147 122 -137
rect 152 -147 153 -137
rect 163 -138 164 -126
rect 240 -147 241 -137
rect 247 -138 248 -126
rect 282 -147 283 -137
rect 163 -147 164 -139
rect 184 -147 185 -139
rect 201 -147 202 -139
rect 275 -147 276 -139
rect 170 -147 171 -141
rect 191 -147 192 -141
rect 205 -142 206 -126
rect 317 -147 318 -141
rect 194 -144 195 -126
rect 205 -147 206 -143
rect 226 -144 227 -126
rect 247 -147 248 -143
rect 131 -146 132 -126
rect 226 -147 227 -145
rect 19 -186 20 -156
rect 23 -157 24 -155
rect 37 -157 38 -155
rect 68 -157 69 -155
rect 72 -186 73 -156
rect 107 -157 108 -155
rect 114 -157 115 -155
rect 124 -186 125 -156
rect 152 -157 153 -155
rect 205 -157 206 -155
rect 212 -157 213 -155
rect 275 -157 276 -155
rect 296 -157 297 -155
rect 306 -186 307 -156
rect 310 -157 311 -155
rect 334 -157 335 -155
rect 345 -157 346 -155
rect 359 -186 360 -156
rect 44 -186 45 -158
rect 100 -159 101 -155
rect 107 -186 108 -158
rect 128 -159 129 -155
rect 163 -159 164 -155
rect 268 -159 269 -155
rect 296 -186 297 -158
rect 310 -186 311 -158
rect 51 -161 52 -155
rect 61 -186 62 -160
rect 79 -161 80 -155
rect 117 -186 118 -160
rect 128 -186 129 -160
rect 159 -186 160 -160
rect 163 -186 164 -160
rect 191 -161 192 -155
rect 201 -161 202 -155
rect 247 -161 248 -155
rect 303 -161 304 -155
rect 313 -165 314 -160
rect 51 -186 52 -162
rect 58 -163 59 -155
rect 86 -163 87 -155
rect 93 -163 94 -155
rect 114 -186 115 -162
rect 180 -163 181 -155
rect 184 -163 185 -155
rect 215 -163 216 -155
rect 219 -186 220 -162
rect 226 -163 227 -155
rect 303 -186 304 -162
rect 324 -163 325 -155
rect 58 -186 59 -164
rect 79 -186 80 -164
rect 86 -186 87 -164
rect 233 -165 234 -155
rect 324 -186 325 -164
rect 93 -186 94 -166
rect 135 -167 136 -155
rect 149 -167 150 -155
rect 191 -186 192 -166
rect 198 -167 199 -155
rect 247 -186 248 -166
rect 135 -186 136 -168
rect 177 -186 178 -168
rect 180 -186 181 -168
rect 317 -169 318 -155
rect 142 -171 143 -155
rect 149 -186 150 -170
rect 156 -171 157 -155
rect 184 -186 185 -170
rect 198 -186 199 -170
rect 240 -171 241 -155
rect 268 -186 269 -170
rect 317 -186 318 -170
rect 166 -173 167 -155
rect 226 -186 227 -172
rect 233 -186 234 -172
rect 299 -186 300 -172
rect 173 -175 174 -155
rect 289 -175 290 -155
rect 121 -177 122 -155
rect 173 -186 174 -176
rect 205 -186 206 -176
rect 275 -186 276 -176
rect 100 -186 101 -178
rect 121 -186 122 -178
rect 254 -179 255 -155
rect 289 -186 290 -178
rect 254 -186 255 -180
rect 282 -181 283 -155
rect 261 -183 262 -155
rect 282 -186 283 -182
rect 212 -186 213 -184
rect 261 -186 262 -184
rect 30 -217 31 -195
rect 72 -196 73 -194
rect 79 -196 80 -194
rect 82 -217 83 -195
rect 86 -196 87 -194
rect 145 -196 146 -194
rect 159 -196 160 -194
rect 219 -196 220 -194
rect 226 -196 227 -194
rect 226 -217 227 -195
rect 226 -196 227 -194
rect 226 -217 227 -195
rect 229 -196 230 -194
rect 282 -196 283 -194
rect 289 -196 290 -194
rect 289 -217 290 -195
rect 289 -196 290 -194
rect 289 -217 290 -195
rect 296 -196 297 -194
rect 324 -196 325 -194
rect 331 -217 332 -195
rect 345 -217 346 -195
rect 359 -196 360 -194
rect 390 -217 391 -195
rect 37 -217 38 -197
rect 61 -198 62 -194
rect 72 -217 73 -197
rect 114 -198 115 -194
rect 121 -217 122 -197
rect 138 -217 139 -197
rect 159 -217 160 -197
rect 261 -198 262 -194
rect 296 -217 297 -197
rect 310 -198 311 -194
rect 352 -198 353 -194
rect 359 -217 360 -197
rect 373 -217 374 -197
rect 380 -217 381 -197
rect 40 -217 41 -199
rect 54 -217 55 -199
rect 58 -217 59 -199
rect 86 -217 87 -199
rect 93 -200 94 -194
rect 93 -217 94 -199
rect 93 -200 94 -194
rect 93 -217 94 -199
rect 100 -200 101 -194
rect 205 -217 206 -199
rect 212 -217 213 -199
rect 254 -200 255 -194
rect 303 -200 304 -194
rect 310 -217 311 -199
rect 352 -217 353 -199
rect 366 -217 367 -199
rect 44 -202 45 -194
rect 114 -217 115 -201
rect 135 -202 136 -194
rect 170 -217 171 -201
rect 180 -202 181 -194
rect 327 -217 328 -201
rect 44 -217 45 -203
rect 79 -217 80 -203
rect 103 -217 104 -203
rect 117 -204 118 -194
rect 135 -217 136 -203
rect 282 -217 283 -203
rect 303 -217 304 -203
rect 341 -217 342 -203
rect 51 -206 52 -194
rect 68 -206 69 -194
rect 107 -206 108 -194
rect 142 -206 143 -194
rect 163 -206 164 -194
rect 177 -217 178 -205
rect 187 -217 188 -205
rect 198 -206 199 -194
rect 215 -206 216 -194
rect 219 -217 220 -205
rect 240 -206 241 -194
rect 275 -206 276 -194
rect 65 -217 66 -207
rect 100 -217 101 -207
rect 128 -208 129 -194
rect 142 -217 143 -207
rect 149 -208 150 -194
rect 163 -217 164 -207
rect 184 -217 185 -207
rect 198 -217 199 -207
rect 233 -208 234 -194
rect 275 -217 276 -207
rect 107 -217 108 -209
rect 128 -217 129 -209
rect 149 -217 150 -209
rect 208 -210 209 -194
rect 243 -210 244 -194
rect 268 -210 269 -194
rect 191 -212 192 -194
rect 191 -217 192 -211
rect 191 -212 192 -194
rect 191 -217 192 -211
rect 215 -217 216 -211
rect 268 -217 269 -211
rect 247 -214 248 -194
rect 261 -217 262 -213
rect 240 -217 241 -215
rect 247 -217 248 -215
rect 254 -217 255 -215
rect 324 -217 325 -215
rect 9 -246 10 -226
rect 40 -227 41 -225
rect 54 -246 55 -226
rect 100 -246 101 -226
rect 107 -246 108 -226
rect 121 -227 122 -225
rect 128 -227 129 -225
rect 156 -227 157 -225
rect 177 -227 178 -225
rect 215 -227 216 -225
rect 222 -246 223 -226
rect 289 -227 290 -225
rect 296 -227 297 -225
rect 296 -246 297 -226
rect 296 -227 297 -225
rect 296 -246 297 -226
rect 310 -227 311 -225
rect 331 -246 332 -226
rect 334 -227 335 -225
rect 373 -227 374 -225
rect 380 -227 381 -225
rect 380 -246 381 -226
rect 380 -227 381 -225
rect 380 -246 381 -226
rect 387 -227 388 -225
rect 394 -246 395 -226
rect 16 -246 17 -228
rect 44 -229 45 -225
rect 65 -229 66 -225
rect 65 -246 66 -228
rect 65 -229 66 -225
rect 65 -246 66 -228
rect 79 -246 80 -228
rect 156 -246 157 -228
rect 159 -229 160 -225
rect 177 -246 178 -228
rect 212 -229 213 -225
rect 338 -246 339 -228
rect 345 -229 346 -225
rect 352 -246 353 -228
rect 355 -229 356 -225
rect 359 -229 360 -225
rect 23 -246 24 -230
rect 58 -231 59 -225
rect 93 -231 94 -225
rect 212 -246 213 -230
rect 233 -231 234 -225
rect 275 -231 276 -225
rect 282 -231 283 -225
rect 317 -246 318 -230
rect 327 -231 328 -225
rect 366 -231 367 -225
rect 30 -233 31 -225
rect 89 -233 90 -225
rect 93 -246 94 -232
rect 187 -233 188 -225
rect 226 -233 227 -225
rect 275 -246 276 -232
rect 289 -246 290 -232
rect 320 -233 321 -225
rect 33 -246 34 -234
rect 310 -246 311 -234
rect 37 -246 38 -236
rect 110 -237 111 -225
rect 114 -237 115 -225
rect 135 -237 136 -225
rect 149 -237 150 -225
rect 173 -246 174 -236
rect 198 -237 199 -225
rect 226 -246 227 -236
rect 233 -246 234 -236
rect 254 -237 255 -225
rect 268 -237 269 -225
rect 282 -246 283 -236
rect 303 -237 304 -225
rect 327 -246 328 -236
rect 51 -239 52 -225
rect 110 -246 111 -238
rect 114 -246 115 -238
rect 121 -246 122 -238
rect 135 -246 136 -238
rect 142 -239 143 -225
rect 149 -246 150 -238
rect 163 -239 164 -225
rect 191 -239 192 -225
rect 198 -246 199 -238
rect 205 -239 206 -225
rect 303 -246 304 -238
rect 58 -246 59 -240
rect 72 -241 73 -225
rect 152 -241 153 -225
rect 163 -246 164 -240
rect 170 -241 171 -225
rect 191 -246 192 -240
rect 208 -246 209 -240
rect 254 -246 255 -240
rect 44 -246 45 -242
rect 152 -246 153 -242
rect 170 -246 171 -242
rect 184 -246 185 -242
rect 240 -243 241 -225
rect 247 -246 248 -242
rect 250 -243 251 -225
rect 261 -243 262 -225
rect 72 -246 73 -244
rect 86 -246 87 -244
rect 219 -245 220 -225
rect 240 -246 241 -244
rect 261 -246 262 -244
rect 268 -246 269 -244
rect 9 -256 10 -254
rect 33 -256 34 -254
rect 37 -293 38 -255
rect 198 -256 199 -254
rect 205 -256 206 -254
rect 233 -256 234 -254
rect 268 -256 269 -254
rect 296 -256 297 -254
rect 345 -256 346 -254
rect 352 -256 353 -254
rect 387 -256 388 -254
rect 394 -256 395 -254
rect 9 -293 10 -257
rect 68 -293 69 -257
rect 72 -258 73 -254
rect 82 -293 83 -257
rect 89 -258 90 -254
rect 114 -258 115 -254
rect 128 -293 129 -257
rect 226 -258 227 -254
rect 282 -258 283 -254
rect 282 -293 283 -257
rect 282 -258 283 -254
rect 282 -293 283 -257
rect 16 -260 17 -254
rect 142 -260 143 -254
rect 145 -260 146 -254
rect 338 -293 339 -259
rect 16 -293 17 -261
rect 114 -293 115 -261
rect 135 -262 136 -254
rect 142 -293 143 -261
rect 149 -262 150 -254
rect 345 -293 346 -261
rect 23 -264 24 -254
rect 75 -293 76 -263
rect 79 -264 80 -254
rect 191 -264 192 -254
rect 208 -293 209 -263
rect 247 -264 248 -254
rect 23 -293 24 -265
rect 79 -293 80 -265
rect 93 -266 94 -254
rect 131 -266 132 -254
rect 149 -293 150 -265
rect 303 -266 304 -254
rect 51 -268 52 -254
rect 163 -268 164 -254
rect 173 -268 174 -254
rect 212 -268 213 -254
rect 215 -293 216 -267
rect 317 -268 318 -254
rect 54 -293 55 -269
rect 243 -293 244 -269
rect 289 -270 290 -254
rect 303 -293 304 -269
rect 310 -270 311 -254
rect 317 -293 318 -269
rect 58 -272 59 -254
rect 86 -272 87 -254
rect 100 -272 101 -254
rect 135 -293 136 -271
rect 156 -272 157 -254
rect 219 -272 220 -254
rect 226 -293 227 -271
rect 240 -272 241 -254
rect 254 -272 255 -254
rect 310 -293 311 -271
rect 58 -293 59 -273
rect 65 -274 66 -254
rect 72 -293 73 -273
rect 86 -293 87 -273
rect 100 -293 101 -273
rect 152 -293 153 -273
rect 159 -293 160 -273
rect 247 -293 248 -273
rect 254 -293 255 -273
rect 275 -274 276 -254
rect 2 -293 3 -275
rect 65 -293 66 -275
rect 107 -276 108 -254
rect 163 -293 164 -275
rect 170 -276 171 -254
rect 219 -293 220 -275
rect 233 -293 234 -275
rect 289 -293 290 -275
rect 107 -293 108 -277
rect 121 -278 122 -254
rect 170 -293 171 -277
rect 198 -293 199 -277
rect 212 -293 213 -277
rect 324 -293 325 -277
rect 121 -293 122 -279
rect 187 -293 188 -279
rect 191 -293 192 -279
rect 331 -280 332 -254
rect 156 -293 157 -281
rect 331 -293 332 -281
rect 177 -284 178 -254
rect 268 -293 269 -283
rect 44 -286 45 -254
rect 177 -293 178 -285
rect 180 -293 181 -285
rect 261 -286 262 -254
rect 44 -293 45 -287
rect 96 -293 97 -287
rect 184 -288 185 -254
rect 296 -293 297 -287
rect 194 -293 195 -289
rect 275 -293 276 -289
rect 222 -292 223 -254
rect 261 -293 262 -291
rect 2 -303 3 -301
rect 30 -303 31 -301
rect 44 -303 45 -301
rect 191 -303 192 -301
rect 205 -303 206 -301
rect 289 -303 290 -301
rect 16 -305 17 -301
rect 75 -340 76 -304
rect 79 -305 80 -301
rect 149 -305 150 -301
rect 156 -305 157 -301
rect 156 -340 157 -304
rect 156 -305 157 -301
rect 156 -340 157 -304
rect 170 -305 171 -301
rect 268 -305 269 -301
rect 23 -307 24 -301
rect 54 -340 55 -306
rect 65 -307 66 -301
rect 163 -307 164 -301
rect 187 -307 188 -301
rect 254 -307 255 -301
rect 261 -307 262 -301
rect 289 -340 290 -306
rect 30 -340 31 -308
rect 58 -309 59 -301
rect 65 -340 66 -308
rect 131 -309 132 -301
rect 135 -309 136 -301
rect 173 -309 174 -301
rect 212 -309 213 -301
rect 303 -309 304 -301
rect 37 -311 38 -301
rect 187 -340 188 -310
rect 212 -340 213 -310
rect 261 -340 262 -310
rect 282 -311 283 -301
rect 303 -340 304 -310
rect 37 -340 38 -312
rect 208 -313 209 -301
rect 215 -313 216 -301
rect 233 -340 234 -312
rect 240 -340 241 -312
rect 282 -340 283 -312
rect 44 -340 45 -314
rect 103 -340 104 -314
rect 107 -315 108 -301
rect 145 -340 146 -314
rect 163 -340 164 -314
rect 184 -315 185 -301
rect 208 -340 209 -314
rect 268 -340 269 -314
rect 51 -317 52 -301
rect 138 -340 139 -316
rect 142 -317 143 -301
rect 149 -340 150 -316
rect 184 -340 185 -316
rect 254 -340 255 -316
rect 58 -340 59 -318
rect 114 -340 115 -318
rect 117 -319 118 -301
rect 324 -319 325 -301
rect 79 -340 80 -320
rect 152 -340 153 -320
rect 215 -340 216 -320
rect 331 -321 332 -301
rect 86 -323 87 -301
rect 93 -340 94 -322
rect 96 -323 97 -301
rect 296 -323 297 -301
rect 324 -340 325 -322
rect 338 -323 339 -301
rect 86 -340 87 -324
rect 121 -325 122 -301
rect 128 -340 129 -324
rect 194 -325 195 -301
rect 229 -340 230 -324
rect 317 -325 318 -301
rect 100 -327 101 -301
rect 170 -340 171 -326
rect 226 -327 227 -301
rect 317 -340 318 -326
rect 110 -340 111 -328
rect 345 -329 346 -301
rect 135 -340 136 -330
rect 247 -331 248 -301
rect 142 -340 143 -332
rect 177 -333 178 -301
rect 219 -333 220 -301
rect 247 -340 248 -332
rect 121 -340 122 -334
rect 177 -340 178 -334
rect 198 -335 199 -301
rect 219 -340 220 -334
rect 243 -335 244 -301
rect 310 -335 311 -301
rect 198 -340 199 -336
rect 275 -337 276 -301
rect 296 -340 297 -336
rect 310 -340 311 -336
rect 201 -340 202 -338
rect 275 -340 276 -338
rect 2 -375 3 -349
rect 114 -375 115 -349
rect 121 -375 122 -349
rect 135 -350 136 -348
rect 145 -350 146 -348
rect 198 -375 199 -349
rect 205 -350 206 -348
rect 317 -350 318 -348
rect 16 -375 17 -351
rect 65 -352 66 -348
rect 79 -352 80 -348
rect 89 -375 90 -351
rect 93 -352 94 -348
rect 100 -375 101 -351
rect 103 -352 104 -348
rect 163 -352 164 -348
rect 170 -352 171 -348
rect 170 -375 171 -351
rect 170 -352 171 -348
rect 170 -375 171 -351
rect 173 -375 174 -351
rect 338 -375 339 -351
rect 23 -375 24 -353
rect 107 -354 108 -348
rect 145 -375 146 -353
rect 191 -354 192 -348
rect 215 -375 216 -353
rect 240 -375 241 -353
rect 243 -354 244 -348
rect 275 -354 276 -348
rect 289 -354 290 -348
rect 317 -375 318 -353
rect 30 -356 31 -348
rect 72 -375 73 -355
rect 75 -375 76 -355
rect 79 -375 80 -355
rect 86 -356 87 -348
rect 117 -356 118 -348
rect 149 -375 150 -355
rect 166 -375 167 -355
rect 177 -356 178 -348
rect 201 -356 202 -348
rect 219 -356 220 -348
rect 331 -375 332 -355
rect 9 -375 10 -357
rect 86 -375 87 -357
rect 93 -375 94 -357
rect 191 -375 192 -357
rect 226 -375 227 -357
rect 233 -358 234 -348
rect 268 -358 269 -348
rect 296 -375 297 -357
rect 299 -358 300 -348
rect 324 -358 325 -348
rect 37 -360 38 -348
rect 135 -375 136 -359
rect 152 -360 153 -348
rect 275 -375 276 -359
rect 303 -360 304 -348
rect 345 -375 346 -359
rect 37 -375 38 -361
rect 96 -375 97 -361
rect 117 -375 118 -361
rect 282 -362 283 -348
rect 310 -362 311 -348
rect 310 -375 311 -361
rect 310 -362 311 -348
rect 310 -375 311 -361
rect 44 -364 45 -348
rect 142 -375 143 -363
rect 163 -375 164 -363
rect 289 -375 290 -363
rect 44 -375 45 -365
rect 180 -375 181 -365
rect 184 -366 185 -348
rect 324 -375 325 -365
rect 51 -375 52 -367
rect 65 -375 66 -367
rect 128 -368 129 -348
rect 219 -375 220 -367
rect 233 -375 234 -367
rect 247 -368 248 -348
rect 254 -368 255 -348
rect 268 -375 269 -367
rect 58 -370 59 -348
rect 107 -375 108 -369
rect 128 -375 129 -369
rect 212 -370 213 -348
rect 247 -375 248 -369
rect 264 -375 265 -369
rect 194 -372 195 -348
rect 254 -375 255 -371
rect 261 -372 262 -348
rect 282 -375 283 -371
rect 205 -375 206 -373
rect 212 -375 213 -373
rect 9 -385 10 -383
rect 54 -416 55 -384
rect 68 -385 69 -383
rect 296 -385 297 -383
rect 306 -385 307 -383
rect 310 -385 311 -383
rect 16 -387 17 -383
rect 61 -387 62 -383
rect 75 -387 76 -383
rect 103 -416 104 -386
rect 107 -387 108 -383
rect 117 -387 118 -383
rect 128 -387 129 -383
rect 212 -416 213 -386
rect 215 -387 216 -383
rect 331 -387 332 -383
rect 23 -389 24 -383
rect 82 -416 83 -388
rect 86 -416 87 -388
rect 114 -389 115 -383
rect 128 -416 129 -388
rect 149 -389 150 -383
rect 152 -416 153 -388
rect 198 -389 199 -383
rect 205 -389 206 -383
rect 215 -416 216 -388
rect 233 -389 234 -383
rect 233 -416 234 -388
rect 233 -389 234 -383
rect 233 -416 234 -388
rect 261 -389 262 -383
rect 317 -389 318 -383
rect 2 -391 3 -383
rect 23 -416 24 -390
rect 30 -391 31 -383
rect 30 -416 31 -390
rect 30 -391 31 -383
rect 30 -416 31 -390
rect 37 -391 38 -383
rect 75 -416 76 -390
rect 93 -391 94 -383
rect 100 -391 101 -383
rect 135 -416 136 -390
rect 142 -391 143 -383
rect 156 -391 157 -383
rect 191 -391 192 -383
rect 194 -391 195 -383
rect 282 -391 283 -383
rect 285 -416 286 -390
rect 296 -416 297 -390
rect 44 -393 45 -383
rect 89 -393 90 -383
rect 96 -416 97 -392
rect 121 -393 122 -383
rect 138 -393 139 -383
rect 191 -416 192 -392
rect 201 -416 202 -392
rect 261 -416 262 -392
rect 271 -416 272 -392
rect 317 -416 318 -392
rect 44 -416 45 -394
rect 58 -395 59 -383
rect 142 -416 143 -394
rect 149 -416 150 -394
rect 163 -416 164 -394
rect 198 -416 199 -394
rect 205 -416 206 -394
rect 243 -416 244 -394
rect 282 -416 283 -394
rect 345 -395 346 -383
rect 51 -397 52 -383
rect 65 -416 66 -396
rect 166 -397 167 -383
rect 219 -397 220 -383
rect 289 -397 290 -383
rect 303 -416 304 -396
rect 40 -416 41 -398
rect 51 -416 52 -398
rect 58 -416 59 -398
rect 79 -399 80 -383
rect 170 -399 171 -383
rect 254 -399 255 -383
rect 292 -416 293 -398
rect 310 -416 311 -398
rect 79 -416 80 -400
rect 107 -416 108 -400
rect 177 -401 178 -383
rect 324 -401 325 -383
rect 177 -416 178 -402
rect 184 -403 185 -383
rect 219 -416 220 -402
rect 226 -403 227 -383
rect 240 -403 241 -383
rect 254 -416 255 -402
rect 156 -416 157 -404
rect 226 -416 227 -404
rect 180 -407 181 -383
rect 289 -416 290 -406
rect 184 -416 185 -408
rect 247 -409 248 -383
rect 247 -416 248 -410
rect 275 -411 276 -383
rect 268 -413 269 -383
rect 275 -416 276 -412
rect 268 -416 269 -414
rect 338 -415 339 -383
rect 2 -447 3 -425
rect 131 -447 132 -425
rect 135 -426 136 -424
rect 226 -426 227 -424
rect 229 -426 230 -424
rect 240 -447 241 -425
rect 254 -426 255 -424
rect 289 -447 290 -425
rect 310 -426 311 -424
rect 310 -447 311 -425
rect 310 -426 311 -424
rect 310 -447 311 -425
rect 317 -426 318 -424
rect 327 -447 328 -425
rect 9 -447 10 -427
rect 44 -428 45 -424
rect 47 -447 48 -427
rect 51 -447 52 -427
rect 54 -428 55 -424
rect 65 -428 66 -424
rect 72 -428 73 -424
rect 96 -428 97 -424
rect 114 -447 115 -427
rect 142 -428 143 -424
rect 149 -447 150 -427
rect 163 -428 164 -424
rect 170 -428 171 -424
rect 177 -428 178 -424
rect 201 -428 202 -424
rect 233 -428 234 -424
rect 268 -428 269 -424
rect 303 -428 304 -424
rect 324 -447 325 -427
rect 338 -447 339 -427
rect 16 -447 17 -429
rect 58 -430 59 -424
rect 65 -447 66 -429
rect 93 -430 94 -424
rect 107 -430 108 -424
rect 163 -447 164 -429
rect 170 -447 171 -429
rect 184 -430 185 -424
rect 205 -430 206 -424
rect 212 -447 213 -429
rect 222 -430 223 -424
rect 317 -447 318 -429
rect 23 -432 24 -424
rect 58 -447 59 -431
rect 79 -447 80 -431
rect 93 -447 94 -431
rect 107 -447 108 -431
rect 121 -447 122 -431
rect 128 -432 129 -424
rect 128 -447 129 -431
rect 128 -432 129 -424
rect 128 -447 129 -431
rect 142 -447 143 -431
rect 156 -432 157 -424
rect 184 -447 185 -431
rect 194 -447 195 -431
rect 201 -447 202 -431
rect 205 -447 206 -431
rect 226 -447 227 -431
rect 282 -432 283 -424
rect 23 -447 24 -433
rect 135 -447 136 -433
rect 233 -447 234 -433
rect 254 -447 255 -433
rect 261 -434 262 -424
rect 303 -447 304 -433
rect 30 -436 31 -424
rect 37 -436 38 -424
rect 72 -447 73 -435
rect 282 -447 283 -435
rect 30 -447 31 -437
rect 86 -438 87 -424
rect 110 -447 111 -437
rect 177 -447 178 -437
rect 219 -438 220 -424
rect 261 -447 262 -437
rect 268 -447 269 -437
rect 296 -438 297 -424
rect 37 -447 38 -439
rect 89 -447 90 -439
rect 173 -440 174 -424
rect 219 -447 220 -439
rect 275 -440 276 -424
rect 275 -447 276 -439
rect 275 -440 276 -424
rect 275 -447 276 -439
rect 82 -447 83 -441
rect 103 -447 104 -441
rect 191 -442 192 -424
rect 296 -447 297 -441
rect 191 -447 192 -443
rect 247 -444 248 -424
rect 156 -447 157 -445
rect 247 -447 248 -445
rect 2 -457 3 -455
rect 89 -457 90 -455
rect 107 -488 108 -456
rect 138 -457 139 -455
rect 170 -488 171 -456
rect 173 -457 174 -455
rect 177 -457 178 -455
rect 191 -488 192 -456
rect 198 -488 199 -456
rect 317 -457 318 -455
rect 320 -488 321 -456
rect 352 -488 353 -456
rect 359 -488 360 -456
rect 366 -488 367 -456
rect 9 -459 10 -455
rect 44 -459 45 -455
rect 75 -459 76 -455
rect 163 -459 164 -455
rect 194 -459 195 -455
rect 317 -488 318 -458
rect 331 -488 332 -458
rect 338 -459 339 -455
rect 16 -461 17 -455
rect 79 -461 80 -455
rect 93 -461 94 -455
rect 163 -488 164 -460
rect 205 -461 206 -455
rect 212 -461 213 -455
rect 215 -461 216 -455
rect 282 -461 283 -455
rect 310 -461 311 -455
rect 334 -461 335 -455
rect 23 -463 24 -455
rect 40 -488 41 -462
rect 44 -488 45 -462
rect 131 -488 132 -462
rect 135 -463 136 -455
rect 303 -463 304 -455
rect 327 -463 328 -455
rect 338 -488 339 -462
rect 30 -465 31 -455
rect 103 -465 104 -455
rect 110 -465 111 -455
rect 296 -465 297 -455
rect 37 -467 38 -455
rect 58 -467 59 -455
rect 93 -488 94 -466
rect 142 -467 143 -455
rect 184 -467 185 -455
rect 205 -488 206 -466
rect 219 -467 220 -455
rect 303 -488 304 -466
rect 51 -469 52 -455
rect 58 -488 59 -468
rect 100 -469 101 -455
rect 177 -488 178 -468
rect 180 -488 181 -468
rect 184 -488 185 -468
rect 219 -488 220 -468
rect 296 -488 297 -468
rect 51 -488 52 -470
rect 75 -488 76 -470
rect 100 -488 101 -470
rect 145 -488 146 -470
rect 226 -471 227 -455
rect 226 -488 227 -470
rect 226 -471 227 -455
rect 226 -488 227 -470
rect 233 -471 234 -455
rect 289 -471 290 -455
rect 114 -473 115 -455
rect 159 -473 160 -455
rect 233 -488 234 -472
rect 268 -473 269 -455
rect 275 -473 276 -455
rect 289 -488 290 -472
rect 114 -488 115 -474
rect 121 -475 122 -455
rect 128 -475 129 -455
rect 222 -488 223 -474
rect 247 -475 248 -455
rect 275 -488 276 -474
rect 121 -488 122 -476
rect 149 -477 150 -455
rect 215 -488 216 -476
rect 247 -488 248 -476
rect 254 -477 255 -455
rect 310 -488 311 -476
rect 86 -479 87 -455
rect 149 -488 150 -478
rect 65 -481 66 -455
rect 86 -488 87 -480
rect 128 -488 129 -480
rect 261 -481 262 -455
rect 61 -483 62 -455
rect 65 -488 66 -482
rect 138 -488 139 -482
rect 156 -488 157 -482
rect 240 -483 241 -455
rect 261 -488 262 -482
rect 142 -488 143 -484
rect 268 -488 269 -484
rect 236 -487 237 -455
rect 240 -488 241 -486
rect 16 -525 17 -497
rect 51 -498 52 -496
rect 65 -498 66 -496
rect 82 -498 83 -496
rect 103 -525 104 -497
rect 180 -498 181 -496
rect 184 -498 185 -496
rect 257 -498 258 -496
rect 282 -498 283 -496
rect 303 -498 304 -496
rect 310 -498 311 -496
rect 324 -525 325 -497
rect 331 -498 332 -496
rect 348 -498 349 -496
rect 352 -498 353 -496
rect 352 -525 353 -497
rect 352 -498 353 -496
rect 352 -525 353 -497
rect 23 -525 24 -499
rect 79 -525 80 -499
rect 114 -500 115 -496
rect 145 -500 146 -496
rect 149 -500 150 -496
rect 184 -525 185 -499
rect 198 -500 199 -496
rect 271 -525 272 -499
rect 275 -500 276 -496
rect 310 -525 311 -499
rect 320 -500 321 -496
rect 338 -500 339 -496
rect 345 -525 346 -499
rect 359 -500 360 -496
rect 30 -525 31 -501
rect 61 -525 62 -501
rect 72 -502 73 -496
rect 86 -502 87 -496
rect 93 -502 94 -496
rect 114 -525 115 -501
rect 121 -525 122 -501
rect 149 -525 150 -501
rect 177 -525 178 -501
rect 338 -525 339 -501
rect 58 -504 59 -496
rect 65 -525 66 -503
rect 72 -525 73 -503
rect 100 -504 101 -496
rect 135 -525 136 -503
rect 194 -525 195 -503
rect 201 -504 202 -496
rect 268 -504 269 -496
rect 296 -504 297 -496
rect 331 -525 332 -503
rect 44 -506 45 -496
rect 100 -525 101 -505
rect 138 -506 139 -496
rect 163 -506 164 -496
rect 180 -525 181 -505
rect 219 -525 220 -505
rect 222 -506 223 -496
rect 317 -525 318 -505
rect 44 -525 45 -507
rect 51 -525 52 -507
rect 86 -525 87 -507
rect 156 -508 157 -496
rect 163 -525 164 -507
rect 170 -508 171 -496
rect 201 -525 202 -507
rect 226 -508 227 -496
rect 229 -525 230 -507
rect 282 -525 283 -507
rect 93 -525 94 -509
rect 128 -510 129 -496
rect 142 -525 143 -509
rect 198 -525 199 -509
rect 226 -525 227 -509
rect 275 -525 276 -509
rect 82 -525 83 -511
rect 128 -525 129 -511
rect 156 -525 157 -511
rect 205 -512 206 -496
rect 233 -512 234 -496
rect 327 -512 328 -496
rect 107 -514 108 -496
rect 170 -525 171 -513
rect 240 -514 241 -496
rect 240 -525 241 -513
rect 240 -514 241 -496
rect 240 -525 241 -513
rect 247 -514 248 -496
rect 303 -525 304 -513
rect 107 -525 108 -515
rect 166 -525 167 -515
rect 191 -516 192 -496
rect 247 -525 248 -515
rect 254 -516 255 -496
rect 289 -516 290 -496
rect 124 -518 125 -496
rect 289 -525 290 -517
rect 159 -525 160 -519
rect 233 -525 234 -519
rect 261 -520 262 -496
rect 296 -525 297 -519
rect 205 -525 206 -521
rect 261 -525 262 -521
rect 212 -525 213 -523
rect 254 -525 255 -523
rect 9 -568 10 -534
rect 33 -568 34 -534
rect 37 -535 38 -533
rect 40 -568 41 -534
rect 51 -535 52 -533
rect 51 -568 52 -534
rect 51 -535 52 -533
rect 51 -568 52 -534
rect 61 -535 62 -533
rect 93 -535 94 -533
rect 100 -568 101 -534
rect 166 -535 167 -533
rect 201 -535 202 -533
rect 205 -568 206 -534
rect 208 -535 209 -533
rect 317 -535 318 -533
rect 331 -535 332 -533
rect 345 -535 346 -533
rect 352 -535 353 -533
rect 362 -568 363 -534
rect 16 -537 17 -533
rect 82 -537 83 -533
rect 86 -537 87 -533
rect 194 -537 195 -533
rect 212 -537 213 -533
rect 310 -537 311 -533
rect 331 -568 332 -536
rect 369 -568 370 -536
rect 16 -568 17 -538
rect 82 -568 83 -538
rect 93 -568 94 -538
rect 215 -539 216 -533
rect 222 -568 223 -538
rect 303 -539 304 -533
rect 23 -541 24 -533
rect 117 -568 118 -540
rect 121 -568 122 -540
rect 135 -541 136 -533
rect 138 -541 139 -533
rect 240 -541 241 -533
rect 250 -568 251 -540
rect 303 -568 304 -540
rect 23 -568 24 -542
rect 58 -543 59 -533
rect 65 -543 66 -533
rect 65 -568 66 -542
rect 65 -543 66 -533
rect 65 -568 66 -542
rect 68 -568 69 -542
rect 86 -568 87 -542
rect 114 -543 115 -533
rect 180 -543 181 -533
rect 191 -543 192 -533
rect 317 -568 318 -542
rect 30 -545 31 -533
rect 44 -545 45 -533
rect 58 -568 59 -544
rect 103 -545 104 -533
rect 124 -545 125 -533
rect 247 -545 248 -533
rect 268 -545 269 -533
rect 310 -568 311 -544
rect 128 -547 129 -533
rect 128 -568 129 -546
rect 128 -547 129 -533
rect 128 -568 129 -546
rect 135 -568 136 -546
rect 212 -568 213 -546
rect 226 -568 227 -546
rect 243 -568 244 -546
rect 247 -568 248 -546
rect 345 -568 346 -546
rect 142 -549 143 -533
rect 142 -568 143 -548
rect 142 -549 143 -533
rect 142 -568 143 -548
rect 156 -549 157 -533
rect 254 -549 255 -533
rect 261 -549 262 -533
rect 268 -568 269 -548
rect 271 -549 272 -533
rect 324 -549 325 -533
rect 107 -551 108 -533
rect 156 -568 157 -550
rect 159 -551 160 -533
rect 170 -551 171 -533
rect 177 -568 178 -550
rect 191 -568 192 -550
rect 233 -551 234 -533
rect 261 -568 262 -550
rect 324 -568 325 -550
rect 338 -551 339 -533
rect 72 -553 73 -533
rect 107 -568 108 -552
rect 163 -553 164 -533
rect 275 -553 276 -533
rect 61 -568 62 -554
rect 72 -568 73 -554
rect 163 -568 164 -554
rect 275 -568 276 -554
rect 166 -568 167 -556
rect 198 -568 199 -556
rect 233 -568 234 -556
rect 352 -568 353 -556
rect 170 -568 171 -558
rect 184 -559 185 -533
rect 254 -568 255 -558
rect 296 -559 297 -533
rect 149 -561 150 -533
rect 184 -568 185 -560
rect 289 -561 290 -533
rect 296 -568 297 -560
rect 282 -563 283 -533
rect 289 -568 290 -562
rect 219 -565 220 -533
rect 282 -568 283 -564
rect 219 -568 220 -566
rect 338 -568 339 -566
rect 9 -578 10 -576
rect 61 -578 62 -576
rect 68 -605 69 -577
rect 79 -578 80 -576
rect 86 -578 87 -576
rect 86 -605 87 -577
rect 86 -578 87 -576
rect 86 -605 87 -577
rect 93 -578 94 -576
rect 103 -605 104 -577
rect 114 -578 115 -576
rect 212 -578 213 -576
rect 219 -578 220 -576
rect 324 -578 325 -576
rect 345 -578 346 -576
rect 369 -578 370 -576
rect 23 -580 24 -576
rect 47 -605 48 -579
rect 72 -580 73 -576
rect 72 -605 73 -579
rect 72 -580 73 -576
rect 72 -605 73 -579
rect 79 -605 80 -579
rect 110 -605 111 -579
rect 114 -605 115 -579
rect 135 -580 136 -576
rect 149 -580 150 -576
rect 184 -580 185 -576
rect 205 -580 206 -576
rect 205 -605 206 -579
rect 205 -580 206 -576
rect 205 -605 206 -579
rect 212 -605 213 -579
rect 275 -580 276 -576
rect 289 -580 290 -576
rect 359 -580 360 -576
rect 44 -582 45 -576
rect 51 -582 52 -576
rect 93 -605 94 -581
rect 121 -582 122 -576
rect 128 -582 129 -576
rect 163 -582 164 -576
rect 177 -582 178 -576
rect 331 -582 332 -576
rect 44 -605 45 -583
rect 51 -605 52 -583
rect 100 -584 101 -576
rect 128 -605 129 -583
rect 135 -605 136 -583
rect 170 -584 171 -576
rect 180 -584 181 -576
rect 282 -584 283 -576
rect 16 -586 17 -576
rect 100 -605 101 -585
rect 121 -605 122 -585
rect 145 -605 146 -585
rect 149 -605 150 -585
rect 170 -605 171 -585
rect 219 -605 220 -585
rect 226 -586 227 -576
rect 229 -605 230 -585
rect 257 -605 258 -585
rect 261 -586 262 -576
rect 275 -605 276 -585
rect 152 -605 153 -587
rect 191 -588 192 -576
rect 233 -588 234 -576
rect 310 -588 311 -576
rect 156 -590 157 -576
rect 222 -590 223 -576
rect 233 -605 234 -589
rect 261 -605 262 -589
rect 264 -605 265 -589
rect 352 -590 353 -576
rect 142 -592 143 -576
rect 156 -605 157 -591
rect 163 -605 164 -591
rect 177 -605 178 -591
rect 191 -605 192 -591
rect 198 -592 199 -576
rect 236 -592 237 -576
rect 240 -592 241 -576
rect 243 -592 244 -576
rect 303 -592 304 -576
rect 310 -605 311 -591
rect 338 -592 339 -576
rect 187 -605 188 -593
rect 198 -605 199 -593
rect 240 -605 241 -593
rect 292 -605 293 -593
rect 247 -605 248 -595
rect 296 -596 297 -576
rect 250 -598 251 -576
rect 317 -598 318 -576
rect 254 -600 255 -576
rect 282 -605 283 -599
rect 254 -605 255 -601
rect 268 -602 269 -576
rect 250 -605 251 -603
rect 268 -605 269 -603
rect 51 -615 52 -613
rect 51 -636 52 -614
rect 51 -615 52 -613
rect 51 -636 52 -614
rect 65 -636 66 -614
rect 68 -615 69 -613
rect 72 -615 73 -613
rect 72 -636 73 -614
rect 72 -615 73 -613
rect 72 -636 73 -614
rect 79 -636 80 -614
rect 107 -636 108 -614
rect 110 -615 111 -613
rect 114 -615 115 -613
rect 128 -615 129 -613
rect 163 -615 164 -613
rect 187 -615 188 -613
rect 240 -615 241 -613
rect 261 -636 262 -614
rect 268 -615 269 -613
rect 289 -615 290 -613
rect 313 -636 314 -614
rect 58 -636 59 -616
rect 68 -636 69 -616
rect 86 -617 87 -613
rect 96 -636 97 -616
rect 100 -636 101 -616
rect 121 -617 122 -613
rect 128 -636 129 -616
rect 138 -636 139 -616
rect 142 -617 143 -613
rect 170 -617 171 -613
rect 194 -617 195 -613
rect 219 -617 220 -613
rect 226 -636 227 -616
rect 250 -617 251 -613
rect 268 -636 269 -616
rect 292 -636 293 -616
rect 303 -636 304 -616
rect 310 -617 311 -613
rect 86 -636 87 -618
rect 103 -636 104 -618
rect 114 -636 115 -618
rect 135 -619 136 -613
rect 142 -636 143 -618
rect 191 -619 192 -613
rect 198 -619 199 -613
rect 254 -636 255 -618
rect 275 -619 276 -613
rect 289 -636 290 -618
rect 93 -621 94 -613
rect 124 -621 125 -613
rect 156 -621 157 -613
rect 184 -621 185 -613
rect 233 -621 234 -613
rect 240 -636 241 -620
rect 257 -621 258 -613
rect 275 -636 276 -620
rect 156 -636 157 -622
rect 208 -636 209 -622
rect 233 -636 234 -622
rect 282 -623 283 -613
rect 163 -636 164 -624
rect 212 -625 213 -613
rect 282 -636 283 -624
rect 299 -636 300 -624
rect 166 -627 167 -613
rect 219 -636 220 -626
rect 170 -636 171 -628
rect 198 -636 199 -628
rect 177 -631 178 -613
rect 212 -636 213 -630
rect 177 -636 178 -632
rect 247 -636 248 -632
rect 184 -636 185 -634
rect 205 -635 206 -613
rect 44 -646 45 -644
rect 51 -646 52 -644
rect 65 -646 66 -644
rect 82 -646 83 -644
rect 96 -646 97 -644
rect 100 -663 101 -645
rect 114 -646 115 -644
rect 152 -646 153 -644
rect 156 -646 157 -644
rect 170 -663 171 -645
rect 173 -646 174 -644
rect 240 -646 241 -644
rect 243 -663 244 -645
rect 261 -646 262 -644
rect 292 -663 293 -645
rect 303 -646 304 -644
rect 44 -663 45 -647
rect 54 -663 55 -647
rect 58 -648 59 -644
rect 65 -663 66 -647
rect 72 -648 73 -644
rect 79 -648 80 -644
rect 107 -648 108 -644
rect 114 -663 115 -647
rect 121 -663 122 -647
rect 135 -663 136 -647
rect 149 -648 150 -644
rect 219 -648 220 -644
rect 233 -648 234 -644
rect 233 -663 234 -647
rect 233 -648 234 -644
rect 233 -663 234 -647
rect 247 -648 248 -644
rect 310 -648 311 -644
rect 72 -663 73 -649
rect 86 -650 87 -644
rect 93 -650 94 -644
rect 107 -663 108 -649
rect 124 -650 125 -644
rect 163 -650 164 -644
rect 180 -650 181 -644
rect 212 -650 213 -644
rect 261 -663 262 -649
rect 282 -650 283 -644
rect 79 -663 80 -651
rect 89 -663 90 -651
rect 128 -652 129 -644
rect 142 -652 143 -644
rect 184 -652 185 -644
rect 205 -663 206 -651
rect 208 -652 209 -644
rect 275 -652 276 -644
rect 142 -663 143 -653
rect 149 -663 150 -653
rect 184 -663 185 -653
rect 222 -663 223 -653
rect 268 -654 269 -644
rect 282 -663 283 -653
rect 191 -656 192 -644
rect 198 -656 199 -644
rect 201 -663 202 -655
rect 254 -656 255 -644
rect 268 -663 269 -655
rect 278 -663 279 -655
rect 191 -663 192 -657
rect 212 -663 213 -657
rect 254 -663 255 -657
rect 264 -663 265 -657
rect 194 -660 195 -644
rect 226 -660 227 -644
rect 226 -663 227 -661
rect 240 -663 241 -661
rect 44 -673 45 -671
rect 51 -678 52 -672
rect 58 -673 59 -671
rect 65 -673 66 -671
rect 72 -673 73 -671
rect 86 -673 87 -671
rect 93 -673 94 -671
rect 100 -673 101 -671
rect 103 -678 104 -672
rect 107 -673 108 -671
rect 114 -673 115 -671
rect 128 -678 129 -672
rect 135 -678 136 -672
rect 138 -673 139 -671
rect 145 -678 146 -672
rect 149 -673 150 -671
rect 170 -673 171 -671
rect 180 -673 181 -671
rect 184 -673 185 -671
rect 201 -673 202 -671
rect 205 -673 206 -671
rect 205 -678 206 -672
rect 205 -673 206 -671
rect 205 -678 206 -672
rect 212 -678 213 -672
rect 226 -673 227 -671
rect 240 -673 241 -671
rect 247 -678 248 -672
rect 254 -673 255 -671
rect 254 -678 255 -672
rect 254 -673 255 -671
rect 254 -678 255 -672
rect 268 -673 269 -671
rect 275 -678 276 -672
rect 285 -673 286 -671
rect 292 -673 293 -671
rect 58 -678 59 -674
rect 65 -678 66 -674
rect 72 -678 73 -674
rect 96 -675 97 -671
rect 121 -678 122 -674
rect 124 -675 125 -671
rect 191 -675 192 -671
rect 219 -675 220 -671
rect 226 -678 227 -674
rect 233 -675 234 -671
rect 240 -678 241 -674
rect 243 -675 244 -671
rect 79 -677 80 -671
rect 79 -678 80 -676
rect 79 -677 80 -671
rect 79 -678 80 -676
rect 191 -678 192 -676
rect 201 -678 202 -676
rect 44 -688 45 -686
rect 51 -688 52 -686
rect 58 -688 59 -686
rect 72 -688 73 -686
rect 79 -688 80 -686
rect 86 -688 87 -686
rect 93 -688 94 -686
rect 114 -688 115 -686
rect 117 -688 118 -686
rect 121 -688 122 -686
rect 135 -688 136 -686
rect 145 -688 146 -686
rect 198 -688 199 -686
rect 205 -688 206 -686
rect 212 -688 213 -686
rect 222 -688 223 -686
rect 226 -688 227 -686
rect 243 -688 244 -686
rect 254 -688 255 -686
rect 264 -688 265 -686
rect 275 -688 276 -686
rect 285 -688 286 -686
rect 107 -690 108 -686
rect 128 -690 129 -686
rect 142 -690 143 -686
rect 152 -690 153 -686
rect 233 -690 234 -686
rect 247 -690 248 -686
<< labels >>
rlabel pdiffusion 3 -8 3 -8 0 cellNo=17
rlabel pdiffusion 10 -8 10 -8 0 cellNo=21
rlabel pdiffusion 17 -8 17 -8 0 cellNo=42
rlabel pdiffusion 24 -8 24 -8 0 cellNo=81
rlabel pdiffusion 31 -8 31 -8 0 cellNo=276
rlabel pdiffusion 136 -8 136 -8 0 feedthrough
rlabel pdiffusion 143 -8 143 -8 0 cellNo=283
rlabel pdiffusion 150 -8 150 -8 0 feedthrough
rlabel pdiffusion 157 -8 157 -8 0 cellNo=106
rlabel pdiffusion 178 -8 178 -8 0 cellNo=137
rlabel pdiffusion 3 -25 3 -25 0 cellNo=25
rlabel pdiffusion 10 -25 10 -25 0 cellNo=355
rlabel pdiffusion 17 -25 17 -25 0 cellNo=69
rlabel pdiffusion 24 -25 24 -25 0 cellNo=152
rlabel pdiffusion 101 -25 101 -25 0 cellNo=338
rlabel pdiffusion 108 -25 108 -25 0 feedthrough
rlabel pdiffusion 122 -25 122 -25 0 cellNo=177
rlabel pdiffusion 129 -25 129 -25 0 cellNo=74
rlabel pdiffusion 136 -25 136 -25 0 feedthrough
rlabel pdiffusion 143 -25 143 -25 0 cellNo=36
rlabel pdiffusion 150 -25 150 -25 0 cellNo=56
rlabel pdiffusion 157 -25 157 -25 0 feedthrough
rlabel pdiffusion 164 -25 164 -25 0 feedthrough
rlabel pdiffusion 171 -25 171 -25 0 feedthrough
rlabel pdiffusion 178 -25 178 -25 0 cellNo=309
rlabel pdiffusion 185 -25 185 -25 0 feedthrough
rlabel pdiffusion 192 -25 192 -25 0 cellNo=24
rlabel pdiffusion 3 -44 3 -44 0 cellNo=45
rlabel pdiffusion 10 -44 10 -44 0 cellNo=64
rlabel pdiffusion 17 -44 17 -44 0 cellNo=114
rlabel pdiffusion 80 -44 80 -44 0 feedthrough
rlabel pdiffusion 87 -44 87 -44 0 feedthrough
rlabel pdiffusion 94 -44 94 -44 0 feedthrough
rlabel pdiffusion 101 -44 101 -44 0 cellNo=103
rlabel pdiffusion 108 -44 108 -44 0 cellNo=318
rlabel pdiffusion 115 -44 115 -44 0 cellNo=37
rlabel pdiffusion 122 -44 122 -44 0 feedthrough
rlabel pdiffusion 129 -44 129 -44 0 feedthrough
rlabel pdiffusion 136 -44 136 -44 0 feedthrough
rlabel pdiffusion 143 -44 143 -44 0 cellNo=101
rlabel pdiffusion 150 -44 150 -44 0 cellNo=232
rlabel pdiffusion 157 -44 157 -44 0 cellNo=29
rlabel pdiffusion 164 -44 164 -44 0 feedthrough
rlabel pdiffusion 171 -44 171 -44 0 feedthrough
rlabel pdiffusion 178 -44 178 -44 0 cellNo=181
rlabel pdiffusion 185 -44 185 -44 0 feedthrough
rlabel pdiffusion 192 -44 192 -44 0 cellNo=122
rlabel pdiffusion 199 -44 199 -44 0 feedthrough
rlabel pdiffusion 206 -44 206 -44 0 feedthrough
rlabel pdiffusion 213 -44 213 -44 0 feedthrough
rlabel pdiffusion 220 -44 220 -44 0 feedthrough
rlabel pdiffusion 227 -44 227 -44 0 feedthrough
rlabel pdiffusion 3 -69 3 -69 0 cellNo=63
rlabel pdiffusion 10 -69 10 -69 0 cellNo=100
rlabel pdiffusion 17 -69 17 -69 0 cellNo=221
rlabel pdiffusion 80 -69 80 -69 0 feedthrough
rlabel pdiffusion 87 -69 87 -69 0 feedthrough
rlabel pdiffusion 94 -69 94 -69 0 feedthrough
rlabel pdiffusion 101 -69 101 -69 0 feedthrough
rlabel pdiffusion 108 -69 108 -69 0 cellNo=173
rlabel pdiffusion 115 -69 115 -69 0 feedthrough
rlabel pdiffusion 122 -69 122 -69 0 cellNo=104
rlabel pdiffusion 129 -69 129 -69 0 cellNo=203
rlabel pdiffusion 136 -69 136 -69 0 cellNo=160
rlabel pdiffusion 143 -69 143 -69 0 cellNo=337
rlabel pdiffusion 150 -69 150 -69 0 cellNo=164
rlabel pdiffusion 157 -69 157 -69 0 cellNo=108
rlabel pdiffusion 164 -69 164 -69 0 feedthrough
rlabel pdiffusion 171 -69 171 -69 0 feedthrough
rlabel pdiffusion 178 -69 178 -69 0 feedthrough
rlabel pdiffusion 185 -69 185 -69 0 cellNo=256
rlabel pdiffusion 192 -69 192 -69 0 feedthrough
rlabel pdiffusion 199 -69 199 -69 0 cellNo=296
rlabel pdiffusion 206 -69 206 -69 0 feedthrough
rlabel pdiffusion 213 -69 213 -69 0 feedthrough
rlabel pdiffusion 220 -69 220 -69 0 cellNo=252
rlabel pdiffusion 227 -69 227 -69 0 feedthrough
rlabel pdiffusion 234 -69 234 -69 0 feedthrough
rlabel pdiffusion 3 -98 3 -98 0 cellNo=82
rlabel pdiffusion 10 -98 10 -98 0 cellNo=335
rlabel pdiffusion 66 -98 66 -98 0 feedthrough
rlabel pdiffusion 73 -98 73 -98 0 feedthrough
rlabel pdiffusion 80 -98 80 -98 0 feedthrough
rlabel pdiffusion 87 -98 87 -98 0 cellNo=46
rlabel pdiffusion 94 -98 94 -98 0 cellNo=7
rlabel pdiffusion 101 -98 101 -98 0 feedthrough
rlabel pdiffusion 108 -98 108 -98 0 cellNo=218
rlabel pdiffusion 115 -98 115 -98 0 feedthrough
rlabel pdiffusion 122 -98 122 -98 0 feedthrough
rlabel pdiffusion 129 -98 129 -98 0 cellNo=275
rlabel pdiffusion 136 -98 136 -98 0 cellNo=27
rlabel pdiffusion 143 -98 143 -98 0 cellNo=130
rlabel pdiffusion 150 -98 150 -98 0 cellNo=272
rlabel pdiffusion 157 -98 157 -98 0 feedthrough
rlabel pdiffusion 164 -98 164 -98 0 feedthrough
rlabel pdiffusion 171 -98 171 -98 0 cellNo=350
rlabel pdiffusion 178 -98 178 -98 0 feedthrough
rlabel pdiffusion 185 -98 185 -98 0 feedthrough
rlabel pdiffusion 192 -98 192 -98 0 feedthrough
rlabel pdiffusion 199 -98 199 -98 0 feedthrough
rlabel pdiffusion 206 -98 206 -98 0 cellNo=31
rlabel pdiffusion 213 -98 213 -98 0 feedthrough
rlabel pdiffusion 220 -98 220 -98 0 cellNo=298
rlabel pdiffusion 227 -98 227 -98 0 feedthrough
rlabel pdiffusion 234 -98 234 -98 0 feedthrough
rlabel pdiffusion 241 -98 241 -98 0 cellNo=68
rlabel pdiffusion 248 -98 248 -98 0 feedthrough
rlabel pdiffusion 255 -98 255 -98 0 feedthrough
rlabel pdiffusion 262 -98 262 -98 0 cellNo=211
rlabel pdiffusion 269 -98 269 -98 0 feedthrough
rlabel pdiffusion 283 -98 283 -98 0 feedthrough
rlabel pdiffusion 3 -123 3 -123 0 cellNo=190
rlabel pdiffusion 31 -123 31 -123 0 cellNo=58
rlabel pdiffusion 45 -123 45 -123 0 cellNo=226
rlabel pdiffusion 52 -123 52 -123 0 feedthrough
rlabel pdiffusion 59 -123 59 -123 0 feedthrough
rlabel pdiffusion 66 -123 66 -123 0 feedthrough
rlabel pdiffusion 73 -123 73 -123 0 cellNo=136
rlabel pdiffusion 80 -123 80 -123 0 cellNo=132
rlabel pdiffusion 87 -123 87 -123 0 feedthrough
rlabel pdiffusion 94 -123 94 -123 0 feedthrough
rlabel pdiffusion 101 -123 101 -123 0 feedthrough
rlabel pdiffusion 108 -123 108 -123 0 feedthrough
rlabel pdiffusion 115 -123 115 -123 0 cellNo=111
rlabel pdiffusion 122 -123 122 -123 0 feedthrough
rlabel pdiffusion 129 -123 129 -123 0 cellNo=38
rlabel pdiffusion 136 -123 136 -123 0 cellNo=61
rlabel pdiffusion 143 -123 143 -123 0 feedthrough
rlabel pdiffusion 150 -123 150 -123 0 feedthrough
rlabel pdiffusion 157 -123 157 -123 0 cellNo=133
rlabel pdiffusion 164 -123 164 -123 0 feedthrough
rlabel pdiffusion 171 -123 171 -123 0 feedthrough
rlabel pdiffusion 178 -123 178 -123 0 feedthrough
rlabel pdiffusion 185 -123 185 -123 0 cellNo=34
rlabel pdiffusion 192 -123 192 -123 0 cellNo=163
rlabel pdiffusion 199 -123 199 -123 0 cellNo=43
rlabel pdiffusion 206 -123 206 -123 0 feedthrough
rlabel pdiffusion 213 -123 213 -123 0 feedthrough
rlabel pdiffusion 220 -123 220 -123 0 cellNo=288
rlabel pdiffusion 227 -123 227 -123 0 feedthrough
rlabel pdiffusion 234 -123 234 -123 0 feedthrough
rlabel pdiffusion 241 -123 241 -123 0 feedthrough
rlabel pdiffusion 248 -123 248 -123 0 feedthrough
rlabel pdiffusion 255 -123 255 -123 0 feedthrough
rlabel pdiffusion 262 -123 262 -123 0 feedthrough
rlabel pdiffusion 269 -123 269 -123 0 cellNo=14
rlabel pdiffusion 276 -123 276 -123 0 feedthrough
rlabel pdiffusion 283 -123 283 -123 0 feedthrough
rlabel pdiffusion 290 -123 290 -123 0 feedthrough
rlabel pdiffusion 297 -123 297 -123 0 cellNo=135
rlabel pdiffusion 304 -123 304 -123 0 feedthrough
rlabel pdiffusion 325 -123 325 -123 0 cellNo=50
rlabel pdiffusion 17 -152 17 -152 0 cellNo=156
rlabel pdiffusion 24 -152 24 -152 0 feedthrough
rlabel pdiffusion 31 -152 31 -152 0 cellNo=305
rlabel pdiffusion 38 -152 38 -152 0 feedthrough
rlabel pdiffusion 45 -152 45 -152 0 cellNo=102
rlabel pdiffusion 52 -152 52 -152 0 cellNo=174
rlabel pdiffusion 59 -152 59 -152 0 feedthrough
rlabel pdiffusion 66 -152 66 -152 0 cellNo=48
rlabel pdiffusion 73 -152 73 -152 0 cellNo=53
rlabel pdiffusion 80 -152 80 -152 0 feedthrough
rlabel pdiffusion 87 -152 87 -152 0 feedthrough
rlabel pdiffusion 94 -152 94 -152 0 cellNo=265
rlabel pdiffusion 101 -152 101 -152 0 feedthrough
rlabel pdiffusion 108 -152 108 -152 0 feedthrough
rlabel pdiffusion 115 -152 115 -152 0 cellNo=112
rlabel pdiffusion 122 -152 122 -152 0 feedthrough
rlabel pdiffusion 129 -152 129 -152 0 cellNo=51
rlabel pdiffusion 136 -152 136 -152 0 feedthrough
rlabel pdiffusion 143 -152 143 -152 0 feedthrough
rlabel pdiffusion 150 -152 150 -152 0 cellNo=332
rlabel pdiffusion 157 -152 157 -152 0 feedthrough
rlabel pdiffusion 164 -152 164 -152 0 cellNo=346
rlabel pdiffusion 171 -152 171 -152 0 cellNo=223
rlabel pdiffusion 178 -152 178 -152 0 cellNo=127
rlabel pdiffusion 185 -152 185 -152 0 feedthrough
rlabel pdiffusion 192 -152 192 -152 0 feedthrough
rlabel pdiffusion 199 -152 199 -152 0 cellNo=60
rlabel pdiffusion 206 -152 206 -152 0 feedthrough
rlabel pdiffusion 213 -152 213 -152 0 cellNo=179
rlabel pdiffusion 220 -152 220 -152 0 cellNo=105
rlabel pdiffusion 227 -152 227 -152 0 feedthrough
rlabel pdiffusion 234 -152 234 -152 0 cellNo=67
rlabel pdiffusion 241 -152 241 -152 0 feedthrough
rlabel pdiffusion 248 -152 248 -152 0 feedthrough
rlabel pdiffusion 255 -152 255 -152 0 feedthrough
rlabel pdiffusion 262 -152 262 -152 0 feedthrough
rlabel pdiffusion 269 -152 269 -152 0 feedthrough
rlabel pdiffusion 276 -152 276 -152 0 feedthrough
rlabel pdiffusion 283 -152 283 -152 0 feedthrough
rlabel pdiffusion 290 -152 290 -152 0 feedthrough
rlabel pdiffusion 297 -152 297 -152 0 feedthrough
rlabel pdiffusion 304 -152 304 -152 0 feedthrough
rlabel pdiffusion 311 -152 311 -152 0 feedthrough
rlabel pdiffusion 318 -152 318 -152 0 feedthrough
rlabel pdiffusion 325 -152 325 -152 0 feedthrough
rlabel pdiffusion 332 -152 332 -152 0 cellNo=92
rlabel pdiffusion 339 -152 339 -152 0 cellNo=66
rlabel pdiffusion 346 -152 346 -152 0 feedthrough
rlabel pdiffusion 17 -191 17 -191 0 cellNo=8
rlabel pdiffusion 45 -191 45 -191 0 feedthrough
rlabel pdiffusion 52 -191 52 -191 0 feedthrough
rlabel pdiffusion 59 -191 59 -191 0 cellNo=15
rlabel pdiffusion 66 -191 66 -191 0 cellNo=214
rlabel pdiffusion 73 -191 73 -191 0 feedthrough
rlabel pdiffusion 80 -191 80 -191 0 feedthrough
rlabel pdiffusion 87 -191 87 -191 0 feedthrough
rlabel pdiffusion 94 -191 94 -191 0 feedthrough
rlabel pdiffusion 101 -191 101 -191 0 feedthrough
rlabel pdiffusion 108 -191 108 -191 0 feedthrough
rlabel pdiffusion 115 -191 115 -191 0 cellNo=250
rlabel pdiffusion 122 -191 122 -191 0 cellNo=22
rlabel pdiffusion 129 -191 129 -191 0 feedthrough
rlabel pdiffusion 136 -191 136 -191 0 feedthrough
rlabel pdiffusion 143 -191 143 -191 0 cellNo=6
rlabel pdiffusion 150 -191 150 -191 0 feedthrough
rlabel pdiffusion 157 -191 157 -191 0 cellNo=324
rlabel pdiffusion 164 -191 164 -191 0 feedthrough
rlabel pdiffusion 171 -191 171 -191 0 cellNo=95
rlabel pdiffusion 178 -191 178 -191 0 cellNo=216
rlabel pdiffusion 185 -191 185 -191 0 cellNo=10
rlabel pdiffusion 192 -191 192 -191 0 feedthrough
rlabel pdiffusion 199 -191 199 -191 0 feedthrough
rlabel pdiffusion 206 -191 206 -191 0 cellNo=193
rlabel pdiffusion 213 -191 213 -191 0 cellNo=210
rlabel pdiffusion 220 -191 220 -191 0 feedthrough
rlabel pdiffusion 227 -191 227 -191 0 cellNo=282
rlabel pdiffusion 234 -191 234 -191 0 feedthrough
rlabel pdiffusion 241 -191 241 -191 0 cellNo=326
rlabel pdiffusion 248 -191 248 -191 0 feedthrough
rlabel pdiffusion 255 -191 255 -191 0 feedthrough
rlabel pdiffusion 262 -191 262 -191 0 feedthrough
rlabel pdiffusion 269 -191 269 -191 0 feedthrough
rlabel pdiffusion 276 -191 276 -191 0 feedthrough
rlabel pdiffusion 283 -191 283 -191 0 feedthrough
rlabel pdiffusion 290 -191 290 -191 0 feedthrough
rlabel pdiffusion 297 -191 297 -191 0 cellNo=12
rlabel pdiffusion 304 -191 304 -191 0 cellNo=229
rlabel pdiffusion 311 -191 311 -191 0 feedthrough
rlabel pdiffusion 318 -191 318 -191 0 cellNo=254
rlabel pdiffusion 325 -191 325 -191 0 feedthrough
rlabel pdiffusion 353 -191 353 -191 0 cellNo=157
rlabel pdiffusion 360 -191 360 -191 0 cellNo=247
rlabel pdiffusion 31 -222 31 -222 0 feedthrough
rlabel pdiffusion 38 -222 38 -222 0 cellNo=98
rlabel pdiffusion 45 -222 45 -222 0 feedthrough
rlabel pdiffusion 52 -222 52 -222 0 cellNo=62
rlabel pdiffusion 59 -222 59 -222 0 feedthrough
rlabel pdiffusion 66 -222 66 -222 0 feedthrough
rlabel pdiffusion 73 -222 73 -222 0 feedthrough
rlabel pdiffusion 80 -222 80 -222 0 cellNo=76
rlabel pdiffusion 87 -222 87 -222 0 cellNo=73
rlabel pdiffusion 94 -222 94 -222 0 feedthrough
rlabel pdiffusion 101 -222 101 -222 0 cellNo=70
rlabel pdiffusion 108 -222 108 -222 0 cellNo=97
rlabel pdiffusion 115 -222 115 -222 0 feedthrough
rlabel pdiffusion 122 -222 122 -222 0 feedthrough
rlabel pdiffusion 129 -222 129 -222 0 feedthrough
rlabel pdiffusion 136 -222 136 -222 0 cellNo=88
rlabel pdiffusion 143 -222 143 -222 0 feedthrough
rlabel pdiffusion 150 -222 150 -222 0 cellNo=5
rlabel pdiffusion 157 -222 157 -222 0 cellNo=233
rlabel pdiffusion 164 -222 164 -222 0 feedthrough
rlabel pdiffusion 171 -222 171 -222 0 feedthrough
rlabel pdiffusion 178 -222 178 -222 0 feedthrough
rlabel pdiffusion 185 -222 185 -222 0 cellNo=93
rlabel pdiffusion 192 -222 192 -222 0 feedthrough
rlabel pdiffusion 199 -222 199 -222 0 feedthrough
rlabel pdiffusion 206 -222 206 -222 0 feedthrough
rlabel pdiffusion 213 -222 213 -222 0 cellNo=9
rlabel pdiffusion 220 -222 220 -222 0 feedthrough
rlabel pdiffusion 227 -222 227 -222 0 feedthrough
rlabel pdiffusion 234 -222 234 -222 0 cellNo=300
rlabel pdiffusion 241 -222 241 -222 0 feedthrough
rlabel pdiffusion 248 -222 248 -222 0 cellNo=225
rlabel pdiffusion 255 -222 255 -222 0 feedthrough
rlabel pdiffusion 262 -222 262 -222 0 feedthrough
rlabel pdiffusion 269 -222 269 -222 0 feedthrough
rlabel pdiffusion 276 -222 276 -222 0 feedthrough
rlabel pdiffusion 283 -222 283 -222 0 feedthrough
rlabel pdiffusion 290 -222 290 -222 0 feedthrough
rlabel pdiffusion 297 -222 297 -222 0 feedthrough
rlabel pdiffusion 304 -222 304 -222 0 feedthrough
rlabel pdiffusion 311 -222 311 -222 0 feedthrough
rlabel pdiffusion 318 -222 318 -222 0 cellNo=201
rlabel pdiffusion 325 -222 325 -222 0 cellNo=317
rlabel pdiffusion 332 -222 332 -222 0 cellNo=99
rlabel pdiffusion 339 -222 339 -222 0 cellNo=244
rlabel pdiffusion 346 -222 346 -222 0 feedthrough
rlabel pdiffusion 353 -222 353 -222 0 cellNo=189
rlabel pdiffusion 360 -222 360 -222 0 feedthrough
rlabel pdiffusion 367 -222 367 -222 0 feedthrough
rlabel pdiffusion 374 -222 374 -222 0 cellNo=199
rlabel pdiffusion 381 -222 381 -222 0 feedthrough
rlabel pdiffusion 388 -222 388 -222 0 cellNo=342
rlabel pdiffusion 10 -251 10 -251 0 feedthrough
rlabel pdiffusion 17 -251 17 -251 0 feedthrough
rlabel pdiffusion 24 -251 24 -251 0 feedthrough
rlabel pdiffusion 31 -251 31 -251 0 cellNo=246
rlabel pdiffusion 38 -251 38 -251 0 cellNo=328
rlabel pdiffusion 45 -251 45 -251 0 feedthrough
rlabel pdiffusion 52 -251 52 -251 0 cellNo=80
rlabel pdiffusion 59 -251 59 -251 0 feedthrough
rlabel pdiffusion 66 -251 66 -251 0 feedthrough
rlabel pdiffusion 73 -251 73 -251 0 feedthrough
rlabel pdiffusion 80 -251 80 -251 0 cellNo=314
rlabel pdiffusion 87 -251 87 -251 0 cellNo=33
rlabel pdiffusion 94 -251 94 -251 0 feedthrough
rlabel pdiffusion 101 -251 101 -251 0 feedthrough
rlabel pdiffusion 108 -251 108 -251 0 cellNo=302
rlabel pdiffusion 115 -251 115 -251 0 cellNo=87
rlabel pdiffusion 122 -251 122 -251 0 feedthrough
rlabel pdiffusion 129 -251 129 -251 0 cellNo=28
rlabel pdiffusion 136 -251 136 -251 0 feedthrough
rlabel pdiffusion 143 -251 143 -251 0 cellNo=212
rlabel pdiffusion 150 -251 150 -251 0 cellNo=269
rlabel pdiffusion 157 -251 157 -251 0 feedthrough
rlabel pdiffusion 164 -251 164 -251 0 feedthrough
rlabel pdiffusion 171 -251 171 -251 0 cellNo=359
rlabel pdiffusion 178 -251 178 -251 0 feedthrough
rlabel pdiffusion 185 -251 185 -251 0 feedthrough
rlabel pdiffusion 192 -251 192 -251 0 feedthrough
rlabel pdiffusion 199 -251 199 -251 0 feedthrough
rlabel pdiffusion 206 -251 206 -251 0 cellNo=339
rlabel pdiffusion 213 -251 213 -251 0 feedthrough
rlabel pdiffusion 220 -251 220 -251 0 cellNo=125
rlabel pdiffusion 227 -251 227 -251 0 feedthrough
rlabel pdiffusion 234 -251 234 -251 0 feedthrough
rlabel pdiffusion 241 -251 241 -251 0 feedthrough
rlabel pdiffusion 248 -251 248 -251 0 feedthrough
rlabel pdiffusion 255 -251 255 -251 0 feedthrough
rlabel pdiffusion 262 -251 262 -251 0 feedthrough
rlabel pdiffusion 269 -251 269 -251 0 cellNo=228
rlabel pdiffusion 276 -251 276 -251 0 feedthrough
rlabel pdiffusion 283 -251 283 -251 0 feedthrough
rlabel pdiffusion 290 -251 290 -251 0 feedthrough
rlabel pdiffusion 297 -251 297 -251 0 feedthrough
rlabel pdiffusion 304 -251 304 -251 0 feedthrough
rlabel pdiffusion 311 -251 311 -251 0 feedthrough
rlabel pdiffusion 318 -251 318 -251 0 feedthrough
rlabel pdiffusion 325 -251 325 -251 0 cellNo=251
rlabel pdiffusion 332 -251 332 -251 0 feedthrough
rlabel pdiffusion 339 -251 339 -251 0 cellNo=240
rlabel pdiffusion 346 -251 346 -251 0 cellNo=154
rlabel pdiffusion 353 -251 353 -251 0 feedthrough
rlabel pdiffusion 381 -251 381 -251 0 cellNo=208
rlabel pdiffusion 388 -251 388 -251 0 cellNo=59
rlabel pdiffusion 395 -251 395 -251 0 feedthrough
rlabel pdiffusion 3 -298 3 -298 0 feedthrough
rlabel pdiffusion 10 -298 10 -298 0 cellNo=344
rlabel pdiffusion 17 -298 17 -298 0 feedthrough
rlabel pdiffusion 24 -298 24 -298 0 feedthrough
rlabel pdiffusion 31 -298 31 -298 0 cellNo=273
rlabel pdiffusion 38 -298 38 -298 0 feedthrough
rlabel pdiffusion 45 -298 45 -298 0 feedthrough
rlabel pdiffusion 52 -298 52 -298 0 cellNo=20
rlabel pdiffusion 59 -298 59 -298 0 feedthrough
rlabel pdiffusion 66 -298 66 -298 0 cellNo=224
rlabel pdiffusion 73 -298 73 -298 0 cellNo=26
rlabel pdiffusion 80 -298 80 -298 0 cellNo=316
rlabel pdiffusion 87 -298 87 -298 0 feedthrough
rlabel pdiffusion 94 -298 94 -298 0 cellNo=90
rlabel pdiffusion 101 -298 101 -298 0 feedthrough
rlabel pdiffusion 108 -298 108 -298 0 feedthrough
rlabel pdiffusion 115 -298 115 -298 0 cellNo=94
rlabel pdiffusion 122 -298 122 -298 0 feedthrough
rlabel pdiffusion 129 -298 129 -298 0 cellNo=148
rlabel pdiffusion 136 -298 136 -298 0 feedthrough
rlabel pdiffusion 143 -298 143 -298 0 feedthrough
rlabel pdiffusion 150 -298 150 -298 0 cellNo=284
rlabel pdiffusion 157 -298 157 -298 0 cellNo=260
rlabel pdiffusion 164 -298 164 -298 0 feedthrough
rlabel pdiffusion 171 -298 171 -298 0 cellNo=30
rlabel pdiffusion 178 -298 178 -298 0 cellNo=1
rlabel pdiffusion 185 -298 185 -298 0 cellNo=162
rlabel pdiffusion 192 -298 192 -298 0 cellNo=129
rlabel pdiffusion 199 -298 199 -298 0 feedthrough
rlabel pdiffusion 206 -298 206 -298 0 cellNo=131
rlabel pdiffusion 213 -298 213 -298 0 cellNo=71
rlabel pdiffusion 220 -298 220 -298 0 feedthrough
rlabel pdiffusion 227 -298 227 -298 0 feedthrough
rlabel pdiffusion 234 -298 234 -298 0 cellNo=290
rlabel pdiffusion 241 -298 241 -298 0 cellNo=235
rlabel pdiffusion 248 -298 248 -298 0 feedthrough
rlabel pdiffusion 255 -298 255 -298 0 feedthrough
rlabel pdiffusion 262 -298 262 -298 0 feedthrough
rlabel pdiffusion 269 -298 269 -298 0 feedthrough
rlabel pdiffusion 276 -298 276 -298 0 feedthrough
rlabel pdiffusion 283 -298 283 -298 0 feedthrough
rlabel pdiffusion 290 -298 290 -298 0 feedthrough
rlabel pdiffusion 297 -298 297 -298 0 feedthrough
rlabel pdiffusion 304 -298 304 -298 0 feedthrough
rlabel pdiffusion 311 -298 311 -298 0 feedthrough
rlabel pdiffusion 318 -298 318 -298 0 feedthrough
rlabel pdiffusion 325 -298 325 -298 0 feedthrough
rlabel pdiffusion 332 -298 332 -298 0 feedthrough
rlabel pdiffusion 339 -298 339 -298 0 feedthrough
rlabel pdiffusion 346 -298 346 -298 0 feedthrough
rlabel pdiffusion 31 -345 31 -345 0 feedthrough
rlabel pdiffusion 38 -345 38 -345 0 feedthrough
rlabel pdiffusion 45 -345 45 -345 0 feedthrough
rlabel pdiffusion 52 -345 52 -345 0 cellNo=3
rlabel pdiffusion 59 -345 59 -345 0 feedthrough
rlabel pdiffusion 66 -345 66 -345 0 feedthrough
rlabel pdiffusion 73 -345 73 -345 0 cellNo=277
rlabel pdiffusion 80 -345 80 -345 0 feedthrough
rlabel pdiffusion 87 -345 87 -345 0 feedthrough
rlabel pdiffusion 94 -345 94 -345 0 feedthrough
rlabel pdiffusion 101 -345 101 -345 0 cellNo=44
rlabel pdiffusion 108 -345 108 -345 0 cellNo=85
rlabel pdiffusion 115 -345 115 -345 0 cellNo=185
rlabel pdiffusion 122 -345 122 -345 0 cellNo=167
rlabel pdiffusion 129 -345 129 -345 0 feedthrough
rlabel pdiffusion 136 -345 136 -345 0 cellNo=77
rlabel pdiffusion 143 -345 143 -345 0 cellNo=249
rlabel pdiffusion 150 -345 150 -345 0 cellNo=222
rlabel pdiffusion 157 -345 157 -345 0 cellNo=304
rlabel pdiffusion 164 -345 164 -345 0 feedthrough
rlabel pdiffusion 171 -345 171 -345 0 feedthrough
rlabel pdiffusion 178 -345 178 -345 0 feedthrough
rlabel pdiffusion 185 -345 185 -345 0 cellNo=75
rlabel pdiffusion 192 -345 192 -345 0 cellNo=204
rlabel pdiffusion 199 -345 199 -345 0 cellNo=171
rlabel pdiffusion 206 -345 206 -345 0 cellNo=49
rlabel pdiffusion 213 -345 213 -345 0 cellNo=334
rlabel pdiffusion 220 -345 220 -345 0 feedthrough
rlabel pdiffusion 227 -345 227 -345 0 cellNo=289
rlabel pdiffusion 234 -345 234 -345 0 feedthrough
rlabel pdiffusion 241 -345 241 -345 0 cellNo=237
rlabel pdiffusion 248 -345 248 -345 0 feedthrough
rlabel pdiffusion 255 -345 255 -345 0 feedthrough
rlabel pdiffusion 262 -345 262 -345 0 feedthrough
rlabel pdiffusion 269 -345 269 -345 0 feedthrough
rlabel pdiffusion 276 -345 276 -345 0 feedthrough
rlabel pdiffusion 283 -345 283 -345 0 feedthrough
rlabel pdiffusion 290 -345 290 -345 0 feedthrough
rlabel pdiffusion 297 -345 297 -345 0 cellNo=336
rlabel pdiffusion 304 -345 304 -345 0 feedthrough
rlabel pdiffusion 311 -345 311 -345 0 feedthrough
rlabel pdiffusion 318 -345 318 -345 0 feedthrough
rlabel pdiffusion 325 -345 325 -345 0 feedthrough
rlabel pdiffusion 3 -380 3 -380 0 feedthrough
rlabel pdiffusion 10 -380 10 -380 0 feedthrough
rlabel pdiffusion 17 -380 17 -380 0 feedthrough
rlabel pdiffusion 24 -380 24 -380 0 feedthrough
rlabel pdiffusion 31 -380 31 -380 0 cellNo=310
rlabel pdiffusion 38 -380 38 -380 0 feedthrough
rlabel pdiffusion 45 -380 45 -380 0 feedthrough
rlabel pdiffusion 52 -380 52 -380 0 feedthrough
rlabel pdiffusion 59 -380 59 -380 0 cellNo=255
rlabel pdiffusion 66 -380 66 -380 0 cellNo=313
rlabel pdiffusion 73 -380 73 -380 0 cellNo=241
rlabel pdiffusion 80 -380 80 -380 0 feedthrough
rlabel pdiffusion 87 -380 87 -380 0 cellNo=267
rlabel pdiffusion 94 -380 94 -380 0 cellNo=65
rlabel pdiffusion 101 -380 101 -380 0 feedthrough
rlabel pdiffusion 108 -380 108 -380 0 feedthrough
rlabel pdiffusion 115 -380 115 -380 0 cellNo=86
rlabel pdiffusion 122 -380 122 -380 0 feedthrough
rlabel pdiffusion 129 -380 129 -380 0 feedthrough
rlabel pdiffusion 136 -380 136 -380 0 cellNo=227
rlabel pdiffusion 143 -380 143 -380 0 cellNo=281
rlabel pdiffusion 150 -380 150 -380 0 feedthrough
rlabel pdiffusion 157 -380 157 -380 0 cellNo=215
rlabel pdiffusion 164 -380 164 -380 0 cellNo=121
rlabel pdiffusion 171 -380 171 -380 0 cellNo=47
rlabel pdiffusion 178 -380 178 -380 0 cellNo=119
rlabel pdiffusion 185 -380 185 -380 0 cellNo=183
rlabel pdiffusion 192 -380 192 -380 0 cellNo=72
rlabel pdiffusion 199 -380 199 -380 0 feedthrough
rlabel pdiffusion 206 -380 206 -380 0 feedthrough
rlabel pdiffusion 213 -380 213 -380 0 cellNo=188
rlabel pdiffusion 220 -380 220 -380 0 feedthrough
rlabel pdiffusion 227 -380 227 -380 0 feedthrough
rlabel pdiffusion 234 -380 234 -380 0 feedthrough
rlabel pdiffusion 241 -380 241 -380 0 feedthrough
rlabel pdiffusion 248 -380 248 -380 0 feedthrough
rlabel pdiffusion 255 -380 255 -380 0 feedthrough
rlabel pdiffusion 262 -380 262 -380 0 cellNo=243
rlabel pdiffusion 269 -380 269 -380 0 feedthrough
rlabel pdiffusion 276 -380 276 -380 0 feedthrough
rlabel pdiffusion 283 -380 283 -380 0 feedthrough
rlabel pdiffusion 290 -380 290 -380 0 feedthrough
rlabel pdiffusion 297 -380 297 -380 0 feedthrough
rlabel pdiffusion 304 -380 304 -380 0 cellNo=182
rlabel pdiffusion 311 -380 311 -380 0 feedthrough
rlabel pdiffusion 318 -380 318 -380 0 feedthrough
rlabel pdiffusion 325 -380 325 -380 0 feedthrough
rlabel pdiffusion 332 -380 332 -380 0 feedthrough
rlabel pdiffusion 339 -380 339 -380 0 feedthrough
rlabel pdiffusion 346 -380 346 -380 0 feedthrough
rlabel pdiffusion 24 -421 24 -421 0 feedthrough
rlabel pdiffusion 31 -421 31 -421 0 feedthrough
rlabel pdiffusion 38 -421 38 -421 0 cellNo=139
rlabel pdiffusion 45 -421 45 -421 0 feedthrough
rlabel pdiffusion 52 -421 52 -421 0 cellNo=41
rlabel pdiffusion 59 -421 59 -421 0 feedthrough
rlabel pdiffusion 66 -421 66 -421 0 feedthrough
rlabel pdiffusion 73 -421 73 -421 0 cellNo=262
rlabel pdiffusion 80 -421 80 -421 0 cellNo=323
rlabel pdiffusion 87 -421 87 -421 0 feedthrough
rlabel pdiffusion 94 -421 94 -421 0 cellNo=124
rlabel pdiffusion 101 -421 101 -421 0 cellNo=308
rlabel pdiffusion 108 -421 108 -421 0 cellNo=322
rlabel pdiffusion 129 -421 129 -421 0 feedthrough
rlabel pdiffusion 136 -421 136 -421 0 feedthrough
rlabel pdiffusion 143 -421 143 -421 0 feedthrough
rlabel pdiffusion 150 -421 150 -421 0 cellNo=138
rlabel pdiffusion 157 -421 157 -421 0 feedthrough
rlabel pdiffusion 164 -421 164 -421 0 feedthrough
rlabel pdiffusion 171 -421 171 -421 0 cellNo=261
rlabel pdiffusion 178 -421 178 -421 0 feedthrough
rlabel pdiffusion 185 -421 185 -421 0 feedthrough
rlabel pdiffusion 192 -421 192 -421 0 feedthrough
rlabel pdiffusion 199 -421 199 -421 0 cellNo=187
rlabel pdiffusion 206 -421 206 -421 0 feedthrough
rlabel pdiffusion 213 -421 213 -421 0 cellNo=245
rlabel pdiffusion 220 -421 220 -421 0 cellNo=57
rlabel pdiffusion 227 -421 227 -421 0 cellNo=312
rlabel pdiffusion 234 -421 234 -421 0 feedthrough
rlabel pdiffusion 241 -421 241 -421 0 cellNo=206
rlabel pdiffusion 248 -421 248 -421 0 feedthrough
rlabel pdiffusion 255 -421 255 -421 0 feedthrough
rlabel pdiffusion 262 -421 262 -421 0 feedthrough
rlabel pdiffusion 269 -421 269 -421 0 cellNo=343
rlabel pdiffusion 276 -421 276 -421 0 feedthrough
rlabel pdiffusion 283 -421 283 -421 0 cellNo=146
rlabel pdiffusion 290 -421 290 -421 0 cellNo=120
rlabel pdiffusion 297 -421 297 -421 0 feedthrough
rlabel pdiffusion 304 -421 304 -421 0 feedthrough
rlabel pdiffusion 311 -421 311 -421 0 feedthrough
rlabel pdiffusion 318 -421 318 -421 0 feedthrough
rlabel pdiffusion 3 -452 3 -452 0 feedthrough
rlabel pdiffusion 10 -452 10 -452 0 feedthrough
rlabel pdiffusion 17 -452 17 -452 0 feedthrough
rlabel pdiffusion 24 -452 24 -452 0 feedthrough
rlabel pdiffusion 31 -452 31 -452 0 feedthrough
rlabel pdiffusion 38 -452 38 -452 0 feedthrough
rlabel pdiffusion 45 -452 45 -452 0 cellNo=161
rlabel pdiffusion 52 -452 52 -452 0 feedthrough
rlabel pdiffusion 59 -452 59 -452 0 cellNo=293
rlabel pdiffusion 66 -452 66 -452 0 feedthrough
rlabel pdiffusion 73 -452 73 -452 0 cellNo=153
rlabel pdiffusion 80 -452 80 -452 0 cellNo=319
rlabel pdiffusion 87 -452 87 -452 0 cellNo=196
rlabel pdiffusion 94 -452 94 -452 0 feedthrough
rlabel pdiffusion 101 -452 101 -452 0 cellNo=333
rlabel pdiffusion 108 -452 108 -452 0 cellNo=107
rlabel pdiffusion 115 -452 115 -452 0 feedthrough
rlabel pdiffusion 122 -452 122 -452 0 feedthrough
rlabel pdiffusion 129 -452 129 -452 0 cellNo=175
rlabel pdiffusion 136 -452 136 -452 0 cellNo=169
rlabel pdiffusion 143 -452 143 -452 0 feedthrough
rlabel pdiffusion 150 -452 150 -452 0 feedthrough
rlabel pdiffusion 157 -452 157 -452 0 cellNo=79
rlabel pdiffusion 164 -452 164 -452 0 feedthrough
rlabel pdiffusion 171 -452 171 -452 0 cellNo=4
rlabel pdiffusion 178 -452 178 -452 0 feedthrough
rlabel pdiffusion 185 -452 185 -452 0 feedthrough
rlabel pdiffusion 192 -452 192 -452 0 cellNo=217
rlabel pdiffusion 199 -452 199 -452 0 cellNo=195
rlabel pdiffusion 206 -452 206 -452 0 feedthrough
rlabel pdiffusion 213 -452 213 -452 0 cellNo=230
rlabel pdiffusion 220 -452 220 -452 0 cellNo=194
rlabel pdiffusion 227 -452 227 -452 0 feedthrough
rlabel pdiffusion 234 -452 234 -452 0 cellNo=266
rlabel pdiffusion 241 -452 241 -452 0 feedthrough
rlabel pdiffusion 248 -452 248 -452 0 feedthrough
rlabel pdiffusion 255 -452 255 -452 0 feedthrough
rlabel pdiffusion 262 -452 262 -452 0 feedthrough
rlabel pdiffusion 269 -452 269 -452 0 feedthrough
rlabel pdiffusion 276 -452 276 -452 0 feedthrough
rlabel pdiffusion 283 -452 283 -452 0 feedthrough
rlabel pdiffusion 290 -452 290 -452 0 feedthrough
rlabel pdiffusion 297 -452 297 -452 0 feedthrough
rlabel pdiffusion 304 -452 304 -452 0 feedthrough
rlabel pdiffusion 311 -452 311 -452 0 feedthrough
rlabel pdiffusion 318 -452 318 -452 0 feedthrough
rlabel pdiffusion 325 -452 325 -452 0 cellNo=271
rlabel pdiffusion 332 -452 332 -452 0 cellNo=52
rlabel pdiffusion 339 -452 339 -452 0 feedthrough
rlabel pdiffusion 38 -493 38 -493 0 cellNo=295
rlabel pdiffusion 45 -493 45 -493 0 feedthrough
rlabel pdiffusion 52 -493 52 -493 0 feedthrough
rlabel pdiffusion 59 -493 59 -493 0 feedthrough
rlabel pdiffusion 66 -493 66 -493 0 feedthrough
rlabel pdiffusion 73 -493 73 -493 0 cellNo=123
rlabel pdiffusion 80 -493 80 -493 0 cellNo=140
rlabel pdiffusion 87 -493 87 -493 0 feedthrough
rlabel pdiffusion 94 -493 94 -493 0 feedthrough
rlabel pdiffusion 101 -493 101 -493 0 feedthrough
rlabel pdiffusion 108 -493 108 -493 0 feedthrough
rlabel pdiffusion 115 -493 115 -493 0 feedthrough
rlabel pdiffusion 122 -493 122 -493 0 cellNo=354
rlabel pdiffusion 129 -493 129 -493 0 cellNo=197
rlabel pdiffusion 136 -493 136 -493 0 cellNo=2
rlabel pdiffusion 143 -493 143 -493 0 cellNo=231
rlabel pdiffusion 150 -493 150 -493 0 feedthrough
rlabel pdiffusion 157 -493 157 -493 0 feedthrough
rlabel pdiffusion 164 -493 164 -493 0 feedthrough
rlabel pdiffusion 171 -493 171 -493 0 feedthrough
rlabel pdiffusion 178 -493 178 -493 0 cellNo=78
rlabel pdiffusion 185 -493 185 -493 0 feedthrough
rlabel pdiffusion 192 -493 192 -493 0 feedthrough
rlabel pdiffusion 199 -493 199 -493 0 cellNo=145
rlabel pdiffusion 206 -493 206 -493 0 feedthrough
rlabel pdiffusion 213 -493 213 -493 0 cellNo=109
rlabel pdiffusion 220 -493 220 -493 0 cellNo=147
rlabel pdiffusion 227 -493 227 -493 0 feedthrough
rlabel pdiffusion 234 -493 234 -493 0 feedthrough
rlabel pdiffusion 241 -493 241 -493 0 feedthrough
rlabel pdiffusion 248 -493 248 -493 0 feedthrough
rlabel pdiffusion 255 -493 255 -493 0 cellNo=259
rlabel pdiffusion 262 -493 262 -493 0 feedthrough
rlabel pdiffusion 269 -493 269 -493 0 feedthrough
rlabel pdiffusion 276 -493 276 -493 0 feedthrough
rlabel pdiffusion 283 -493 283 -493 0 cellNo=32
rlabel pdiffusion 290 -493 290 -493 0 feedthrough
rlabel pdiffusion 297 -493 297 -493 0 feedthrough
rlabel pdiffusion 304 -493 304 -493 0 feedthrough
rlabel pdiffusion 311 -493 311 -493 0 feedthrough
rlabel pdiffusion 318 -493 318 -493 0 cellNo=242
rlabel pdiffusion 325 -493 325 -493 0 cellNo=287
rlabel pdiffusion 332 -493 332 -493 0 feedthrough
rlabel pdiffusion 339 -493 339 -493 0 feedthrough
rlabel pdiffusion 346 -493 346 -493 0 cellNo=307
rlabel pdiffusion 353 -493 353 -493 0 feedthrough
rlabel pdiffusion 360 -493 360 -493 0 feedthrough
rlabel pdiffusion 367 -493 367 -493 0 cellNo=303
rlabel pdiffusion 17 -530 17 -530 0 feedthrough
rlabel pdiffusion 24 -530 24 -530 0 feedthrough
rlabel pdiffusion 31 -530 31 -530 0 feedthrough
rlabel pdiffusion 38 -530 38 -530 0 cellNo=170
rlabel pdiffusion 45 -530 45 -530 0 cellNo=294
rlabel pdiffusion 52 -530 52 -530 0 feedthrough
rlabel pdiffusion 59 -530 59 -530 0 cellNo=151
rlabel pdiffusion 66 -530 66 -530 0 feedthrough
rlabel pdiffusion 73 -530 73 -530 0 feedthrough
rlabel pdiffusion 80 -530 80 -530 0 cellNo=116
rlabel pdiffusion 87 -530 87 -530 0 feedthrough
rlabel pdiffusion 94 -530 94 -530 0 feedthrough
rlabel pdiffusion 101 -530 101 -530 0 cellNo=200
rlabel pdiffusion 108 -530 108 -530 0 feedthrough
rlabel pdiffusion 115 -530 115 -530 0 feedthrough
rlabel pdiffusion 122 -530 122 -530 0 cellNo=239
rlabel pdiffusion 129 -530 129 -530 0 feedthrough
rlabel pdiffusion 136 -530 136 -530 0 cellNo=39
rlabel pdiffusion 143 -530 143 -530 0 feedthrough
rlabel pdiffusion 150 -530 150 -530 0 feedthrough
rlabel pdiffusion 157 -530 157 -530 0 cellNo=16
rlabel pdiffusion 164 -530 164 -530 0 cellNo=166
rlabel pdiffusion 171 -530 171 -530 0 feedthrough
rlabel pdiffusion 178 -530 178 -530 0 cellNo=270
rlabel pdiffusion 185 -530 185 -530 0 feedthrough
rlabel pdiffusion 192 -530 192 -530 0 cellNo=54
rlabel pdiffusion 199 -530 199 -530 0 cellNo=159
rlabel pdiffusion 206 -530 206 -530 0 cellNo=144
rlabel pdiffusion 213 -530 213 -530 0 cellNo=345
rlabel pdiffusion 220 -530 220 -530 0 feedthrough
rlabel pdiffusion 227 -530 227 -530 0 cellNo=142
rlabel pdiffusion 234 -530 234 -530 0 feedthrough
rlabel pdiffusion 241 -530 241 -530 0 feedthrough
rlabel pdiffusion 248 -530 248 -530 0 feedthrough
rlabel pdiffusion 255 -530 255 -530 0 feedthrough
rlabel pdiffusion 262 -530 262 -530 0 feedthrough
rlabel pdiffusion 269 -530 269 -530 0 cellNo=172
rlabel pdiffusion 276 -530 276 -530 0 feedthrough
rlabel pdiffusion 283 -530 283 -530 0 feedthrough
rlabel pdiffusion 290 -530 290 -530 0 feedthrough
rlabel pdiffusion 297 -530 297 -530 0 feedthrough
rlabel pdiffusion 304 -530 304 -530 0 feedthrough
rlabel pdiffusion 311 -530 311 -530 0 feedthrough
rlabel pdiffusion 318 -530 318 -530 0 feedthrough
rlabel pdiffusion 325 -530 325 -530 0 feedthrough
rlabel pdiffusion 332 -530 332 -530 0 cellNo=213
rlabel pdiffusion 339 -530 339 -530 0 feedthrough
rlabel pdiffusion 346 -530 346 -530 0 feedthrough
rlabel pdiffusion 353 -530 353 -530 0 feedthrough
rlabel pdiffusion 10 -573 10 -573 0 feedthrough
rlabel pdiffusion 17 -573 17 -573 0 feedthrough
rlabel pdiffusion 24 -573 24 -573 0 feedthrough
rlabel pdiffusion 31 -573 31 -573 0 cellNo=202
rlabel pdiffusion 38 -573 38 -573 0 cellNo=128
rlabel pdiffusion 45 -573 45 -573 0 cellNo=96
rlabel pdiffusion 52 -573 52 -573 0 feedthrough
rlabel pdiffusion 59 -573 59 -573 0 cellNo=150
rlabel pdiffusion 66 -573 66 -573 0 cellNo=253
rlabel pdiffusion 73 -573 73 -573 0 feedthrough
rlabel pdiffusion 80 -573 80 -573 0 cellNo=329
rlabel pdiffusion 87 -573 87 -573 0 feedthrough
rlabel pdiffusion 94 -573 94 -573 0 feedthrough
rlabel pdiffusion 101 -573 101 -573 0 feedthrough
rlabel pdiffusion 108 -573 108 -573 0 cellNo=89
rlabel pdiffusion 115 -573 115 -573 0 cellNo=352
rlabel pdiffusion 122 -573 122 -573 0 feedthrough
rlabel pdiffusion 129 -573 129 -573 0 feedthrough
rlabel pdiffusion 136 -573 136 -573 0 cellNo=168
rlabel pdiffusion 143 -573 143 -573 0 feedthrough
rlabel pdiffusion 150 -573 150 -573 0 cellNo=357
rlabel pdiffusion 157 -573 157 -573 0 feedthrough
rlabel pdiffusion 164 -573 164 -573 0 cellNo=84
rlabel pdiffusion 171 -573 171 -573 0 feedthrough
rlabel pdiffusion 178 -573 178 -573 0 cellNo=40
rlabel pdiffusion 185 -573 185 -573 0 feedthrough
rlabel pdiffusion 192 -573 192 -573 0 feedthrough
rlabel pdiffusion 199 -573 199 -573 0 feedthrough
rlabel pdiffusion 206 -573 206 -573 0 feedthrough
rlabel pdiffusion 213 -573 213 -573 0 feedthrough
rlabel pdiffusion 220 -573 220 -573 0 cellNo=353
rlabel pdiffusion 227 -573 227 -573 0 feedthrough
rlabel pdiffusion 234 -573 234 -573 0 cellNo=192
rlabel pdiffusion 241 -573 241 -573 0 cellNo=347
rlabel pdiffusion 248 -573 248 -573 0 cellNo=219
rlabel pdiffusion 255 -573 255 -573 0 feedthrough
rlabel pdiffusion 262 -573 262 -573 0 feedthrough
rlabel pdiffusion 269 -573 269 -573 0 feedthrough
rlabel pdiffusion 276 -573 276 -573 0 feedthrough
rlabel pdiffusion 283 -573 283 -573 0 feedthrough
rlabel pdiffusion 290 -573 290 -573 0 feedthrough
rlabel pdiffusion 297 -573 297 -573 0 feedthrough
rlabel pdiffusion 304 -573 304 -573 0 feedthrough
rlabel pdiffusion 311 -573 311 -573 0 feedthrough
rlabel pdiffusion 318 -573 318 -573 0 feedthrough
rlabel pdiffusion 325 -573 325 -573 0 feedthrough
rlabel pdiffusion 332 -573 332 -573 0 feedthrough
rlabel pdiffusion 339 -573 339 -573 0 feedthrough
rlabel pdiffusion 346 -573 346 -573 0 feedthrough
rlabel pdiffusion 353 -573 353 -573 0 feedthrough
rlabel pdiffusion 360 -573 360 -573 0 cellNo=180
rlabel pdiffusion 367 -573 367 -573 0 cellNo=176
rlabel pdiffusion 45 -610 45 -610 0 cellNo=348
rlabel pdiffusion 52 -610 52 -610 0 feedthrough
rlabel pdiffusion 66 -610 66 -610 0 cellNo=264
rlabel pdiffusion 73 -610 73 -610 0 feedthrough
rlabel pdiffusion 80 -610 80 -610 0 cellNo=321
rlabel pdiffusion 87 -610 87 -610 0 feedthrough
rlabel pdiffusion 94 -610 94 -610 0 feedthrough
rlabel pdiffusion 101 -610 101 -610 0 cellNo=178
rlabel pdiffusion 108 -610 108 -610 0 cellNo=19
rlabel pdiffusion 115 -610 115 -610 0 feedthrough
rlabel pdiffusion 122 -610 122 -610 0 cellNo=55
rlabel pdiffusion 129 -610 129 -610 0 feedthrough
rlabel pdiffusion 136 -610 136 -610 0 feedthrough
rlabel pdiffusion 143 -610 143 -610 0 cellNo=340
rlabel pdiffusion 150 -610 150 -610 0 cellNo=113
rlabel pdiffusion 157 -610 157 -610 0 feedthrough
rlabel pdiffusion 164 -610 164 -610 0 cellNo=278
rlabel pdiffusion 171 -610 171 -610 0 feedthrough
rlabel pdiffusion 178 -610 178 -610 0 feedthrough
rlabel pdiffusion 185 -610 185 -610 0 cellNo=83
rlabel pdiffusion 192 -610 192 -610 0 cellNo=220
rlabel pdiffusion 199 -610 199 -610 0 feedthrough
rlabel pdiffusion 206 -610 206 -610 0 feedthrough
rlabel pdiffusion 213 -610 213 -610 0 cellNo=351
rlabel pdiffusion 220 -610 220 -610 0 feedthrough
rlabel pdiffusion 227 -610 227 -610 0 cellNo=191
rlabel pdiffusion 234 -610 234 -610 0 feedthrough
rlabel pdiffusion 241 -610 241 -610 0 feedthrough
rlabel pdiffusion 248 -610 248 -610 0 cellNo=248
rlabel pdiffusion 255 -610 255 -610 0 cellNo=349
rlabel pdiffusion 262 -610 262 -610 0 cellNo=356
rlabel pdiffusion 269 -610 269 -610 0 feedthrough
rlabel pdiffusion 276 -610 276 -610 0 cellNo=115
rlabel pdiffusion 283 -610 283 -610 0 feedthrough
rlabel pdiffusion 290 -610 290 -610 0 cellNo=165
rlabel pdiffusion 311 -610 311 -610 0 feedthrough
rlabel pdiffusion 45 -641 45 -641 0 cellNo=91
rlabel pdiffusion 52 -641 52 -641 0 feedthrough
rlabel pdiffusion 59 -641 59 -641 0 feedthrough
rlabel pdiffusion 66 -641 66 -641 0 cellNo=134
rlabel pdiffusion 73 -641 73 -641 0 feedthrough
rlabel pdiffusion 80 -641 80 -641 0 cellNo=263
rlabel pdiffusion 87 -641 87 -641 0 feedthrough
rlabel pdiffusion 94 -641 94 -641 0 cellNo=315
rlabel pdiffusion 101 -641 101 -641 0 cellNo=126
rlabel pdiffusion 108 -641 108 -641 0 feedthrough
rlabel pdiffusion 115 -641 115 -641 0 feedthrough
rlabel pdiffusion 122 -641 122 -641 0 cellNo=18
rlabel pdiffusion 129 -641 129 -641 0 feedthrough
rlabel pdiffusion 136 -641 136 -641 0 cellNo=285
rlabel pdiffusion 143 -641 143 -641 0 cellNo=155
rlabel pdiffusion 150 -641 150 -641 0 cellNo=257
rlabel pdiffusion 157 -641 157 -641 0 feedthrough
rlabel pdiffusion 164 -641 164 -641 0 feedthrough
rlabel pdiffusion 171 -641 171 -641 0 cellNo=360
rlabel pdiffusion 178 -641 178 -641 0 cellNo=331
rlabel pdiffusion 185 -641 185 -641 0 feedthrough
rlabel pdiffusion 192 -641 192 -641 0 cellNo=258
rlabel pdiffusion 199 -641 199 -641 0 feedthrough
rlabel pdiffusion 206 -641 206 -641 0 cellNo=320
rlabel pdiffusion 213 -641 213 -641 0 feedthrough
rlabel pdiffusion 220 -641 220 -641 0 feedthrough
rlabel pdiffusion 227 -641 227 -641 0 feedthrough
rlabel pdiffusion 234 -641 234 -641 0 feedthrough
rlabel pdiffusion 241 -641 241 -641 0 feedthrough
rlabel pdiffusion 248 -641 248 -641 0 feedthrough
rlabel pdiffusion 255 -641 255 -641 0 feedthrough
rlabel pdiffusion 262 -641 262 -641 0 feedthrough
rlabel pdiffusion 269 -641 269 -641 0 feedthrough
rlabel pdiffusion 276 -641 276 -641 0 feedthrough
rlabel pdiffusion 283 -641 283 -641 0 feedthrough
rlabel pdiffusion 290 -641 290 -641 0 cellNo=186
rlabel pdiffusion 297 -641 297 -641 0 cellNo=297
rlabel pdiffusion 304 -641 304 -641 0 feedthrough
rlabel pdiffusion 311 -641 311 -641 0 cellNo=280
rlabel pdiffusion 45 -668 45 -668 0 feedthrough
rlabel pdiffusion 52 -668 52 -668 0 cellNo=291
rlabel pdiffusion 59 -668 59 -668 0 cellNo=13
rlabel pdiffusion 66 -668 66 -668 0 feedthrough
rlabel pdiffusion 73 -668 73 -668 0 feedthrough
rlabel pdiffusion 80 -668 80 -668 0 feedthrough
rlabel pdiffusion 87 -668 87 -668 0 cellNo=158
rlabel pdiffusion 94 -668 94 -668 0 cellNo=143
rlabel pdiffusion 101 -668 101 -668 0 cellNo=184
rlabel pdiffusion 108 -668 108 -668 0 feedthrough
rlabel pdiffusion 115 -668 115 -668 0 feedthrough
rlabel pdiffusion 122 -668 122 -668 0 cellNo=207
rlabel pdiffusion 136 -668 136 -668 0 cellNo=330
rlabel pdiffusion 143 -668 143 -668 0 cellNo=118
rlabel pdiffusion 150 -668 150 -668 0 feedthrough
rlabel pdiffusion 171 -668 171 -668 0 feedthrough
rlabel pdiffusion 178 -668 178 -668 0 cellNo=117
rlabel pdiffusion 185 -668 185 -668 0 feedthrough
rlabel pdiffusion 192 -668 192 -668 0 feedthrough
rlabel pdiffusion 199 -668 199 -668 0 cellNo=327
rlabel pdiffusion 206 -668 206 -668 0 feedthrough
rlabel pdiffusion 213 -668 213 -668 0 cellNo=292
rlabel pdiffusion 220 -668 220 -668 0 cellNo=301
rlabel pdiffusion 227 -668 227 -668 0 feedthrough
rlabel pdiffusion 234 -668 234 -668 0 feedthrough
rlabel pdiffusion 241 -668 241 -668 0 cellNo=299
rlabel pdiffusion 255 -668 255 -668 0 feedthrough
rlabel pdiffusion 262 -668 262 -668 0 cellNo=274
rlabel pdiffusion 269 -668 269 -668 0 feedthrough
rlabel pdiffusion 276 -668 276 -668 0 cellNo=198
rlabel pdiffusion 283 -668 283 -668 0 cellNo=141
rlabel pdiffusion 290 -668 290 -668 0 cellNo=110
rlabel pdiffusion 45 -683 45 -683 0 cellNo=279
rlabel pdiffusion 52 -683 52 -683 0 feedthrough
rlabel pdiffusion 59 -683 59 -683 0 feedthrough
rlabel pdiffusion 66 -683 66 -683 0 cellNo=311
rlabel pdiffusion 73 -683 73 -683 0 cellNo=234
rlabel pdiffusion 80 -683 80 -683 0 feedthrough
rlabel pdiffusion 87 -683 87 -683 0 cellNo=11
rlabel pdiffusion 94 -683 94 -683 0 cellNo=268
rlabel pdiffusion 101 -683 101 -683 0 cellNo=358
rlabel pdiffusion 108 -683 108 -683 0 cellNo=23
rlabel pdiffusion 115 -683 115 -683 0 cellNo=236
rlabel pdiffusion 122 -683 122 -683 0 feedthrough
rlabel pdiffusion 129 -683 129 -683 0 feedthrough
rlabel pdiffusion 136 -683 136 -683 0 feedthrough
rlabel pdiffusion 143 -683 143 -683 0 cellNo=149
rlabel pdiffusion 150 -683 150 -683 0 cellNo=238
rlabel pdiffusion 192 -683 192 -683 0 cellNo=286
rlabel pdiffusion 199 -683 199 -683 0 cellNo=341
rlabel pdiffusion 206 -683 206 -683 0 feedthrough
rlabel pdiffusion 213 -683 213 -683 0 feedthrough
rlabel pdiffusion 220 -683 220 -683 0 cellNo=205
rlabel pdiffusion 227 -683 227 -683 0 feedthrough
rlabel pdiffusion 234 -683 234 -683 0 cellNo=209
rlabel pdiffusion 241 -683 241 -683 0 cellNo=306
rlabel pdiffusion 248 -683 248 -683 0 feedthrough
rlabel pdiffusion 255 -683 255 -683 0 feedthrough
rlabel pdiffusion 262 -683 262 -683 0 cellNo=325
rlabel pdiffusion 276 -683 276 -683 0 feedthrough
rlabel pdiffusion 283 -683 283 -683 0 cellNo=35
rlabel polysilicon 135 -4 135 -4 0 1
rlabel polysilicon 135 -10 135 -10 0 3
rlabel polysilicon 142 -4 142 -4 0 1
rlabel polysilicon 145 -4 145 -4 0 2
rlabel polysilicon 149 -4 149 -4 0 1
rlabel polysilicon 149 -10 149 -10 0 3
rlabel polysilicon 159 -10 159 -10 0 4
rlabel polysilicon 177 -10 177 -10 0 3
rlabel polysilicon 100 -21 100 -21 0 1
rlabel polysilicon 107 -21 107 -21 0 1
rlabel polysilicon 107 -27 107 -27 0 3
rlabel polysilicon 121 -21 121 -21 0 1
rlabel polysilicon 128 -21 128 -21 0 1
rlabel polysilicon 135 -21 135 -21 0 1
rlabel polysilicon 135 -27 135 -27 0 3
rlabel polysilicon 142 -21 142 -21 0 1
rlabel polysilicon 145 -21 145 -21 0 2
rlabel polysilicon 142 -27 142 -27 0 3
rlabel polysilicon 152 -21 152 -21 0 2
rlabel polysilicon 152 -27 152 -27 0 4
rlabel polysilicon 156 -21 156 -21 0 1
rlabel polysilicon 156 -27 156 -27 0 3
rlabel polysilicon 163 -21 163 -21 0 1
rlabel polysilicon 163 -27 163 -27 0 3
rlabel polysilicon 170 -21 170 -21 0 1
rlabel polysilicon 170 -27 170 -27 0 3
rlabel polysilicon 177 -21 177 -21 0 1
rlabel polysilicon 180 -21 180 -21 0 2
rlabel polysilicon 184 -21 184 -21 0 1
rlabel polysilicon 184 -27 184 -27 0 3
rlabel polysilicon 191 -27 191 -27 0 3
rlabel polysilicon 79 -40 79 -40 0 1
rlabel polysilicon 79 -46 79 -46 0 3
rlabel polysilicon 86 -40 86 -40 0 1
rlabel polysilicon 86 -46 86 -46 0 3
rlabel polysilicon 93 -40 93 -40 0 1
rlabel polysilicon 93 -46 93 -46 0 3
rlabel polysilicon 100 -40 100 -40 0 1
rlabel polysilicon 103 -40 103 -40 0 2
rlabel polysilicon 107 -46 107 -46 0 3
rlabel polysilicon 110 -46 110 -46 0 4
rlabel polysilicon 117 -40 117 -40 0 2
rlabel polysilicon 114 -46 114 -46 0 3
rlabel polysilicon 121 -40 121 -40 0 1
rlabel polysilicon 121 -46 121 -46 0 3
rlabel polysilicon 128 -40 128 -40 0 1
rlabel polysilicon 128 -46 128 -46 0 3
rlabel polysilicon 135 -40 135 -40 0 1
rlabel polysilicon 135 -46 135 -46 0 3
rlabel polysilicon 142 -40 142 -40 0 1
rlabel polysilicon 142 -46 142 -46 0 3
rlabel polysilicon 145 -46 145 -46 0 4
rlabel polysilicon 149 -40 149 -40 0 1
rlabel polysilicon 152 -40 152 -40 0 2
rlabel polysilicon 149 -46 149 -46 0 3
rlabel polysilicon 159 -40 159 -40 0 2
rlabel polysilicon 156 -46 156 -46 0 3
rlabel polysilicon 163 -40 163 -40 0 1
rlabel polysilicon 163 -46 163 -46 0 3
rlabel polysilicon 170 -40 170 -40 0 1
rlabel polysilicon 170 -46 170 -46 0 3
rlabel polysilicon 180 -40 180 -40 0 2
rlabel polysilicon 180 -46 180 -46 0 4
rlabel polysilicon 184 -40 184 -40 0 1
rlabel polysilicon 184 -46 184 -46 0 3
rlabel polysilicon 194 -40 194 -40 0 2
rlabel polysilicon 191 -46 191 -46 0 3
rlabel polysilicon 198 -40 198 -40 0 1
rlabel polysilicon 198 -46 198 -46 0 3
rlabel polysilicon 205 -40 205 -40 0 1
rlabel polysilicon 205 -46 205 -46 0 3
rlabel polysilicon 212 -40 212 -40 0 1
rlabel polysilicon 212 -46 212 -46 0 3
rlabel polysilicon 219 -40 219 -40 0 1
rlabel polysilicon 219 -46 219 -46 0 3
rlabel polysilicon 226 -40 226 -40 0 1
rlabel polysilicon 226 -46 226 -46 0 3
rlabel polysilicon 79 -65 79 -65 0 1
rlabel polysilicon 79 -71 79 -71 0 3
rlabel polysilicon 86 -65 86 -65 0 1
rlabel polysilicon 86 -71 86 -71 0 3
rlabel polysilicon 93 -65 93 -65 0 1
rlabel polysilicon 93 -71 93 -71 0 3
rlabel polysilicon 100 -65 100 -65 0 1
rlabel polysilicon 100 -71 100 -71 0 3
rlabel polysilicon 110 -65 110 -65 0 2
rlabel polysilicon 107 -71 107 -71 0 3
rlabel polysilicon 114 -65 114 -65 0 1
rlabel polysilicon 114 -71 114 -71 0 3
rlabel polysilicon 121 -71 121 -71 0 3
rlabel polysilicon 124 -71 124 -71 0 4
rlabel polysilicon 131 -65 131 -65 0 2
rlabel polysilicon 131 -71 131 -71 0 4
rlabel polysilicon 138 -65 138 -65 0 2
rlabel polysilicon 135 -71 135 -71 0 3
rlabel polysilicon 138 -71 138 -71 0 4
rlabel polysilicon 142 -65 142 -65 0 1
rlabel polysilicon 145 -65 145 -65 0 2
rlabel polysilicon 142 -71 142 -71 0 3
rlabel polysilicon 149 -65 149 -65 0 1
rlabel polysilicon 152 -65 152 -65 0 2
rlabel polysilicon 156 -65 156 -65 0 1
rlabel polysilicon 156 -71 156 -71 0 3
rlabel polysilicon 159 -71 159 -71 0 4
rlabel polysilicon 163 -65 163 -65 0 1
rlabel polysilicon 163 -71 163 -71 0 3
rlabel polysilicon 170 -65 170 -65 0 1
rlabel polysilicon 170 -71 170 -71 0 3
rlabel polysilicon 177 -65 177 -65 0 1
rlabel polysilicon 177 -71 177 -71 0 3
rlabel polysilicon 187 -65 187 -65 0 2
rlabel polysilicon 191 -65 191 -65 0 1
rlabel polysilicon 191 -71 191 -71 0 3
rlabel polysilicon 198 -71 198 -71 0 3
rlabel polysilicon 205 -65 205 -65 0 1
rlabel polysilicon 205 -71 205 -71 0 3
rlabel polysilicon 212 -65 212 -65 0 1
rlabel polysilicon 212 -71 212 -71 0 3
rlabel polysilicon 222 -65 222 -65 0 2
rlabel polysilicon 226 -65 226 -65 0 1
rlabel polysilicon 226 -71 226 -71 0 3
rlabel polysilicon 233 -65 233 -65 0 1
rlabel polysilicon 233 -71 233 -71 0 3
rlabel polysilicon 65 -94 65 -94 0 1
rlabel polysilicon 65 -100 65 -100 0 3
rlabel polysilicon 72 -94 72 -94 0 1
rlabel polysilicon 72 -100 72 -100 0 3
rlabel polysilicon 79 -94 79 -94 0 1
rlabel polysilicon 79 -100 79 -100 0 3
rlabel polysilicon 86 -94 86 -94 0 1
rlabel polysilicon 93 -94 93 -94 0 1
rlabel polysilicon 93 -100 93 -100 0 3
rlabel polysilicon 100 -94 100 -94 0 1
rlabel polysilicon 100 -100 100 -100 0 3
rlabel polysilicon 107 -94 107 -94 0 1
rlabel polysilicon 107 -100 107 -100 0 3
rlabel polysilicon 114 -94 114 -94 0 1
rlabel polysilicon 114 -100 114 -100 0 3
rlabel polysilicon 121 -94 121 -94 0 1
rlabel polysilicon 121 -100 121 -100 0 3
rlabel polysilicon 128 -94 128 -94 0 1
rlabel polysilicon 131 -100 131 -100 0 4
rlabel polysilicon 138 -94 138 -94 0 2
rlabel polysilicon 135 -100 135 -100 0 3
rlabel polysilicon 142 -94 142 -94 0 1
rlabel polysilicon 142 -100 142 -100 0 3
rlabel polysilicon 152 -94 152 -94 0 2
rlabel polysilicon 149 -100 149 -100 0 3
rlabel polysilicon 152 -100 152 -100 0 4
rlabel polysilicon 156 -94 156 -94 0 1
rlabel polysilicon 156 -100 156 -100 0 3
rlabel polysilicon 163 -94 163 -94 0 1
rlabel polysilicon 163 -100 163 -100 0 3
rlabel polysilicon 170 -94 170 -94 0 1
rlabel polysilicon 173 -100 173 -100 0 4
rlabel polysilicon 177 -94 177 -94 0 1
rlabel polysilicon 177 -100 177 -100 0 3
rlabel polysilicon 184 -94 184 -94 0 1
rlabel polysilicon 184 -100 184 -100 0 3
rlabel polysilicon 191 -94 191 -94 0 1
rlabel polysilicon 191 -100 191 -100 0 3
rlabel polysilicon 198 -94 198 -94 0 1
rlabel polysilicon 198 -100 198 -100 0 3
rlabel polysilicon 205 -94 205 -94 0 1
rlabel polysilicon 205 -100 205 -100 0 3
rlabel polysilicon 212 -94 212 -94 0 1
rlabel polysilicon 212 -100 212 -100 0 3
rlabel polysilicon 219 -94 219 -94 0 1
rlabel polysilicon 222 -94 222 -94 0 2
rlabel polysilicon 219 -100 219 -100 0 3
rlabel polysilicon 226 -94 226 -94 0 1
rlabel polysilicon 226 -100 226 -100 0 3
rlabel polysilicon 233 -94 233 -94 0 1
rlabel polysilicon 233 -100 233 -100 0 3
rlabel polysilicon 240 -94 240 -94 0 1
rlabel polysilicon 243 -94 243 -94 0 2
rlabel polysilicon 243 -100 243 -100 0 4
rlabel polysilicon 247 -94 247 -94 0 1
rlabel polysilicon 247 -100 247 -100 0 3
rlabel polysilicon 254 -94 254 -94 0 1
rlabel polysilicon 254 -100 254 -100 0 3
rlabel polysilicon 261 -94 261 -94 0 1
rlabel polysilicon 264 -100 264 -100 0 4
rlabel polysilicon 268 -94 268 -94 0 1
rlabel polysilicon 268 -100 268 -100 0 3
rlabel polysilicon 282 -94 282 -94 0 1
rlabel polysilicon 282 -100 282 -100 0 3
rlabel polysilicon 33 -125 33 -125 0 4
rlabel polysilicon 44 -119 44 -119 0 1
rlabel polysilicon 51 -119 51 -119 0 1
rlabel polysilicon 51 -125 51 -125 0 3
rlabel polysilicon 58 -119 58 -119 0 1
rlabel polysilicon 58 -125 58 -125 0 3
rlabel polysilicon 65 -119 65 -119 0 1
rlabel polysilicon 65 -125 65 -125 0 3
rlabel polysilicon 75 -119 75 -119 0 2
rlabel polysilicon 79 -125 79 -125 0 3
rlabel polysilicon 82 -125 82 -125 0 4
rlabel polysilicon 86 -119 86 -119 0 1
rlabel polysilicon 86 -125 86 -125 0 3
rlabel polysilicon 93 -119 93 -119 0 1
rlabel polysilicon 93 -125 93 -125 0 3
rlabel polysilicon 100 -119 100 -119 0 1
rlabel polysilicon 100 -125 100 -125 0 3
rlabel polysilicon 107 -119 107 -119 0 1
rlabel polysilicon 107 -125 107 -125 0 3
rlabel polysilicon 114 -119 114 -119 0 1
rlabel polysilicon 117 -119 117 -119 0 2
rlabel polysilicon 114 -125 114 -125 0 3
rlabel polysilicon 121 -119 121 -119 0 1
rlabel polysilicon 121 -125 121 -125 0 3
rlabel polysilicon 128 -119 128 -119 0 1
rlabel polysilicon 128 -125 128 -125 0 3
rlabel polysilicon 131 -125 131 -125 0 4
rlabel polysilicon 138 -119 138 -119 0 2
rlabel polysilicon 142 -119 142 -119 0 1
rlabel polysilicon 142 -125 142 -125 0 3
rlabel polysilicon 149 -119 149 -119 0 1
rlabel polysilicon 149 -125 149 -125 0 3
rlabel polysilicon 156 -119 156 -119 0 1
rlabel polysilicon 159 -119 159 -119 0 2
rlabel polysilicon 156 -125 156 -125 0 3
rlabel polysilicon 159 -125 159 -125 0 4
rlabel polysilicon 163 -119 163 -119 0 1
rlabel polysilicon 163 -125 163 -125 0 3
rlabel polysilicon 170 -119 170 -119 0 1
rlabel polysilicon 170 -125 170 -125 0 3
rlabel polysilicon 177 -119 177 -119 0 1
rlabel polysilicon 177 -125 177 -125 0 3
rlabel polysilicon 184 -119 184 -119 0 1
rlabel polysilicon 184 -125 184 -125 0 3
rlabel polysilicon 191 -125 191 -125 0 3
rlabel polysilicon 194 -125 194 -125 0 4
rlabel polysilicon 201 -119 201 -119 0 2
rlabel polysilicon 198 -125 198 -125 0 3
rlabel polysilicon 205 -119 205 -119 0 1
rlabel polysilicon 205 -125 205 -125 0 3
rlabel polysilicon 212 -119 212 -119 0 1
rlabel polysilicon 212 -125 212 -125 0 3
rlabel polysilicon 219 -119 219 -119 0 1
rlabel polysilicon 222 -119 222 -119 0 2
rlabel polysilicon 226 -119 226 -119 0 1
rlabel polysilicon 226 -125 226 -125 0 3
rlabel polysilicon 233 -119 233 -119 0 1
rlabel polysilicon 233 -125 233 -125 0 3
rlabel polysilicon 240 -119 240 -119 0 1
rlabel polysilicon 240 -125 240 -125 0 3
rlabel polysilicon 247 -119 247 -119 0 1
rlabel polysilicon 247 -125 247 -125 0 3
rlabel polysilicon 254 -119 254 -119 0 1
rlabel polysilicon 254 -125 254 -125 0 3
rlabel polysilicon 261 -119 261 -119 0 1
rlabel polysilicon 261 -125 261 -125 0 3
rlabel polysilicon 271 -125 271 -125 0 4
rlabel polysilicon 275 -119 275 -119 0 1
rlabel polysilicon 275 -125 275 -125 0 3
rlabel polysilicon 282 -119 282 -119 0 1
rlabel polysilicon 282 -125 282 -125 0 3
rlabel polysilicon 289 -119 289 -119 0 1
rlabel polysilicon 289 -125 289 -125 0 3
rlabel polysilicon 296 -119 296 -119 0 1
rlabel polysilicon 299 -119 299 -119 0 2
rlabel polysilicon 299 -125 299 -125 0 4
rlabel polysilicon 303 -119 303 -119 0 1
rlabel polysilicon 303 -125 303 -125 0 3
rlabel polysilicon 324 -125 324 -125 0 3
rlabel polysilicon 19 -148 19 -148 0 2
rlabel polysilicon 23 -148 23 -148 0 1
rlabel polysilicon 23 -154 23 -154 0 3
rlabel polysilicon 30 -148 30 -148 0 1
rlabel polysilicon 37 -148 37 -148 0 1
rlabel polysilicon 37 -154 37 -154 0 3
rlabel polysilicon 47 -148 47 -148 0 2
rlabel polysilicon 51 -154 51 -154 0 3
rlabel polysilicon 58 -148 58 -148 0 1
rlabel polysilicon 58 -154 58 -154 0 3
rlabel polysilicon 65 -148 65 -148 0 1
rlabel polysilicon 68 -148 68 -148 0 2
rlabel polysilicon 68 -154 68 -154 0 4
rlabel polysilicon 72 -148 72 -148 0 1
rlabel polysilicon 79 -148 79 -148 0 1
rlabel polysilicon 79 -154 79 -154 0 3
rlabel polysilicon 86 -148 86 -148 0 1
rlabel polysilicon 86 -154 86 -154 0 3
rlabel polysilicon 93 -148 93 -148 0 1
rlabel polysilicon 96 -148 96 -148 0 2
rlabel polysilicon 93 -154 93 -154 0 3
rlabel polysilicon 100 -148 100 -148 0 1
rlabel polysilicon 100 -154 100 -154 0 3
rlabel polysilicon 107 -148 107 -148 0 1
rlabel polysilicon 107 -154 107 -154 0 3
rlabel polysilicon 114 -148 114 -148 0 1
rlabel polysilicon 114 -154 114 -154 0 3
rlabel polysilicon 121 -148 121 -148 0 1
rlabel polysilicon 121 -154 121 -154 0 3
rlabel polysilicon 128 -154 128 -154 0 3
rlabel polysilicon 135 -148 135 -148 0 1
rlabel polysilicon 135 -154 135 -154 0 3
rlabel polysilicon 142 -148 142 -148 0 1
rlabel polysilicon 142 -154 142 -154 0 3
rlabel polysilicon 149 -148 149 -148 0 1
rlabel polysilicon 152 -148 152 -148 0 2
rlabel polysilicon 149 -154 149 -154 0 3
rlabel polysilicon 152 -154 152 -154 0 4
rlabel polysilicon 156 -148 156 -148 0 1
rlabel polysilicon 156 -154 156 -154 0 3
rlabel polysilicon 163 -148 163 -148 0 1
rlabel polysilicon 166 -148 166 -148 0 2
rlabel polysilicon 163 -154 163 -154 0 3
rlabel polysilicon 166 -154 166 -154 0 4
rlabel polysilicon 170 -148 170 -148 0 1
rlabel polysilicon 173 -148 173 -148 0 2
rlabel polysilicon 173 -154 173 -154 0 4
rlabel polysilicon 177 -148 177 -148 0 1
rlabel polysilicon 180 -154 180 -154 0 4
rlabel polysilicon 184 -148 184 -148 0 1
rlabel polysilicon 184 -154 184 -154 0 3
rlabel polysilicon 191 -148 191 -148 0 1
rlabel polysilicon 191 -154 191 -154 0 3
rlabel polysilicon 201 -148 201 -148 0 2
rlabel polysilicon 198 -154 198 -154 0 3
rlabel polysilicon 201 -154 201 -154 0 4
rlabel polysilicon 205 -148 205 -148 0 1
rlabel polysilicon 205 -154 205 -154 0 3
rlabel polysilicon 212 -154 212 -154 0 3
rlabel polysilicon 215 -154 215 -154 0 4
rlabel polysilicon 219 -148 219 -148 0 1
rlabel polysilicon 226 -148 226 -148 0 1
rlabel polysilicon 226 -154 226 -154 0 3
rlabel polysilicon 236 -148 236 -148 0 2
rlabel polysilicon 233 -154 233 -154 0 3
rlabel polysilicon 240 -148 240 -148 0 1
rlabel polysilicon 240 -154 240 -154 0 3
rlabel polysilicon 247 -148 247 -148 0 1
rlabel polysilicon 247 -154 247 -154 0 3
rlabel polysilicon 254 -148 254 -148 0 1
rlabel polysilicon 254 -154 254 -154 0 3
rlabel polysilicon 261 -148 261 -148 0 1
rlabel polysilicon 261 -154 261 -154 0 3
rlabel polysilicon 268 -148 268 -148 0 1
rlabel polysilicon 268 -154 268 -154 0 3
rlabel polysilicon 275 -148 275 -148 0 1
rlabel polysilicon 275 -154 275 -154 0 3
rlabel polysilicon 282 -148 282 -148 0 1
rlabel polysilicon 282 -154 282 -154 0 3
rlabel polysilicon 289 -148 289 -148 0 1
rlabel polysilicon 289 -154 289 -154 0 3
rlabel polysilicon 296 -148 296 -148 0 1
rlabel polysilicon 296 -154 296 -154 0 3
rlabel polysilicon 303 -148 303 -148 0 1
rlabel polysilicon 303 -154 303 -154 0 3
rlabel polysilicon 310 -148 310 -148 0 1
rlabel polysilicon 310 -154 310 -154 0 3
rlabel polysilicon 317 -148 317 -148 0 1
rlabel polysilicon 317 -154 317 -154 0 3
rlabel polysilicon 324 -148 324 -148 0 1
rlabel polysilicon 324 -154 324 -154 0 3
rlabel polysilicon 331 -148 331 -148 0 1
rlabel polysilicon 334 -154 334 -154 0 4
rlabel polysilicon 341 -148 341 -148 0 2
rlabel polysilicon 345 -148 345 -148 0 1
rlabel polysilicon 345 -154 345 -154 0 3
rlabel polysilicon 19 -187 19 -187 0 2
rlabel polysilicon 44 -187 44 -187 0 1
rlabel polysilicon 44 -193 44 -193 0 3
rlabel polysilicon 51 -187 51 -187 0 1
rlabel polysilicon 51 -193 51 -193 0 3
rlabel polysilicon 58 -187 58 -187 0 1
rlabel polysilicon 61 -187 61 -187 0 2
rlabel polysilicon 61 -193 61 -193 0 4
rlabel polysilicon 68 -193 68 -193 0 4
rlabel polysilicon 72 -187 72 -187 0 1
rlabel polysilicon 72 -193 72 -193 0 3
rlabel polysilicon 79 -187 79 -187 0 1
rlabel polysilicon 79 -193 79 -193 0 3
rlabel polysilicon 86 -187 86 -187 0 1
rlabel polysilicon 86 -193 86 -193 0 3
rlabel polysilicon 93 -187 93 -187 0 1
rlabel polysilicon 93 -193 93 -193 0 3
rlabel polysilicon 100 -187 100 -187 0 1
rlabel polysilicon 100 -193 100 -193 0 3
rlabel polysilicon 107 -187 107 -187 0 1
rlabel polysilicon 107 -193 107 -193 0 3
rlabel polysilicon 114 -187 114 -187 0 1
rlabel polysilicon 117 -187 117 -187 0 2
rlabel polysilicon 114 -193 114 -193 0 3
rlabel polysilicon 117 -193 117 -193 0 4
rlabel polysilicon 121 -187 121 -187 0 1
rlabel polysilicon 124 -187 124 -187 0 2
rlabel polysilicon 128 -187 128 -187 0 1
rlabel polysilicon 128 -193 128 -193 0 3
rlabel polysilicon 135 -187 135 -187 0 1
rlabel polysilicon 135 -193 135 -193 0 3
rlabel polysilicon 142 -193 142 -193 0 3
rlabel polysilicon 145 -193 145 -193 0 4
rlabel polysilicon 149 -187 149 -187 0 1
rlabel polysilicon 149 -193 149 -193 0 3
rlabel polysilicon 159 -187 159 -187 0 2
rlabel polysilicon 159 -193 159 -193 0 4
rlabel polysilicon 163 -187 163 -187 0 1
rlabel polysilicon 163 -193 163 -193 0 3
rlabel polysilicon 173 -187 173 -187 0 2
rlabel polysilicon 177 -187 177 -187 0 1
rlabel polysilicon 180 -187 180 -187 0 2
rlabel polysilicon 180 -193 180 -193 0 4
rlabel polysilicon 184 -187 184 -187 0 1
rlabel polysilicon 191 -187 191 -187 0 1
rlabel polysilicon 191 -193 191 -193 0 3
rlabel polysilicon 198 -187 198 -187 0 1
rlabel polysilicon 198 -193 198 -193 0 3
rlabel polysilicon 205 -187 205 -187 0 1
rlabel polysilicon 208 -193 208 -193 0 4
rlabel polysilicon 212 -187 212 -187 0 1
rlabel polysilicon 215 -193 215 -193 0 4
rlabel polysilicon 219 -187 219 -187 0 1
rlabel polysilicon 219 -193 219 -193 0 3
rlabel polysilicon 226 -187 226 -187 0 1
rlabel polysilicon 226 -193 226 -193 0 3
rlabel polysilicon 229 -193 229 -193 0 4
rlabel polysilicon 233 -187 233 -187 0 1
rlabel polysilicon 233 -193 233 -193 0 3
rlabel polysilicon 240 -193 240 -193 0 3
rlabel polysilicon 243 -193 243 -193 0 4
rlabel polysilicon 247 -187 247 -187 0 1
rlabel polysilicon 247 -193 247 -193 0 3
rlabel polysilicon 254 -187 254 -187 0 1
rlabel polysilicon 254 -193 254 -193 0 3
rlabel polysilicon 261 -187 261 -187 0 1
rlabel polysilicon 261 -193 261 -193 0 3
rlabel polysilicon 268 -187 268 -187 0 1
rlabel polysilicon 268 -193 268 -193 0 3
rlabel polysilicon 275 -187 275 -187 0 1
rlabel polysilicon 275 -193 275 -193 0 3
rlabel polysilicon 282 -187 282 -187 0 1
rlabel polysilicon 282 -193 282 -193 0 3
rlabel polysilicon 289 -187 289 -187 0 1
rlabel polysilicon 289 -193 289 -193 0 3
rlabel polysilicon 296 -187 296 -187 0 1
rlabel polysilicon 299 -187 299 -187 0 2
rlabel polysilicon 296 -193 296 -193 0 3
rlabel polysilicon 303 -187 303 -187 0 1
rlabel polysilicon 306 -187 306 -187 0 2
rlabel polysilicon 303 -193 303 -193 0 3
rlabel polysilicon 310 -187 310 -187 0 1
rlabel polysilicon 310 -193 310 -193 0 3
rlabel polysilicon 317 -187 317 -187 0 1
rlabel polysilicon 324 -187 324 -187 0 1
rlabel polysilicon 324 -193 324 -193 0 3
rlabel polysilicon 352 -193 352 -193 0 3
rlabel polysilicon 359 -187 359 -187 0 1
rlabel polysilicon 359 -193 359 -193 0 3
rlabel polysilicon 30 -218 30 -218 0 1
rlabel polysilicon 30 -224 30 -224 0 3
rlabel polysilicon 37 -218 37 -218 0 1
rlabel polysilicon 40 -218 40 -218 0 2
rlabel polysilicon 40 -224 40 -224 0 4
rlabel polysilicon 44 -218 44 -218 0 1
rlabel polysilicon 44 -224 44 -224 0 3
rlabel polysilicon 54 -218 54 -218 0 2
rlabel polysilicon 51 -224 51 -224 0 3
rlabel polysilicon 58 -218 58 -218 0 1
rlabel polysilicon 58 -224 58 -224 0 3
rlabel polysilicon 65 -218 65 -218 0 1
rlabel polysilicon 65 -224 65 -224 0 3
rlabel polysilicon 72 -218 72 -218 0 1
rlabel polysilicon 72 -224 72 -224 0 3
rlabel polysilicon 79 -218 79 -218 0 1
rlabel polysilicon 82 -218 82 -218 0 2
rlabel polysilicon 86 -218 86 -218 0 1
rlabel polysilicon 89 -224 89 -224 0 4
rlabel polysilicon 93 -218 93 -218 0 1
rlabel polysilicon 93 -224 93 -224 0 3
rlabel polysilicon 100 -218 100 -218 0 1
rlabel polysilicon 103 -218 103 -218 0 2
rlabel polysilicon 107 -218 107 -218 0 1
rlabel polysilicon 110 -224 110 -224 0 4
rlabel polysilicon 114 -218 114 -218 0 1
rlabel polysilicon 114 -224 114 -224 0 3
rlabel polysilicon 121 -218 121 -218 0 1
rlabel polysilicon 121 -224 121 -224 0 3
rlabel polysilicon 128 -218 128 -218 0 1
rlabel polysilicon 128 -224 128 -224 0 3
rlabel polysilicon 135 -218 135 -218 0 1
rlabel polysilicon 138 -218 138 -218 0 2
rlabel polysilicon 135 -224 135 -224 0 3
rlabel polysilicon 142 -218 142 -218 0 1
rlabel polysilicon 142 -224 142 -224 0 3
rlabel polysilicon 149 -218 149 -218 0 1
rlabel polysilicon 149 -224 149 -224 0 3
rlabel polysilicon 152 -224 152 -224 0 4
rlabel polysilicon 159 -218 159 -218 0 2
rlabel polysilicon 156 -224 156 -224 0 3
rlabel polysilicon 159 -224 159 -224 0 4
rlabel polysilicon 163 -218 163 -218 0 1
rlabel polysilicon 163 -224 163 -224 0 3
rlabel polysilicon 170 -218 170 -218 0 1
rlabel polysilicon 170 -224 170 -224 0 3
rlabel polysilicon 177 -218 177 -218 0 1
rlabel polysilicon 177 -224 177 -224 0 3
rlabel polysilicon 184 -218 184 -218 0 1
rlabel polysilicon 187 -218 187 -218 0 2
rlabel polysilicon 187 -224 187 -224 0 4
rlabel polysilicon 191 -218 191 -218 0 1
rlabel polysilicon 191 -224 191 -224 0 3
rlabel polysilicon 198 -218 198 -218 0 1
rlabel polysilicon 198 -224 198 -224 0 3
rlabel polysilicon 205 -218 205 -218 0 1
rlabel polysilicon 205 -224 205 -224 0 3
rlabel polysilicon 212 -218 212 -218 0 1
rlabel polysilicon 215 -218 215 -218 0 2
rlabel polysilicon 212 -224 212 -224 0 3
rlabel polysilicon 215 -224 215 -224 0 4
rlabel polysilicon 219 -218 219 -218 0 1
rlabel polysilicon 219 -224 219 -224 0 3
rlabel polysilicon 226 -218 226 -218 0 1
rlabel polysilicon 226 -224 226 -224 0 3
rlabel polysilicon 233 -224 233 -224 0 3
rlabel polysilicon 240 -218 240 -218 0 1
rlabel polysilicon 240 -224 240 -224 0 3
rlabel polysilicon 247 -218 247 -218 0 1
rlabel polysilicon 250 -224 250 -224 0 4
rlabel polysilicon 254 -218 254 -218 0 1
rlabel polysilicon 254 -224 254 -224 0 3
rlabel polysilicon 261 -218 261 -218 0 1
rlabel polysilicon 261 -224 261 -224 0 3
rlabel polysilicon 268 -218 268 -218 0 1
rlabel polysilicon 268 -224 268 -224 0 3
rlabel polysilicon 275 -218 275 -218 0 1
rlabel polysilicon 275 -224 275 -224 0 3
rlabel polysilicon 282 -218 282 -218 0 1
rlabel polysilicon 282 -224 282 -224 0 3
rlabel polysilicon 289 -218 289 -218 0 1
rlabel polysilicon 289 -224 289 -224 0 3
rlabel polysilicon 296 -218 296 -218 0 1
rlabel polysilicon 296 -224 296 -224 0 3
rlabel polysilicon 303 -218 303 -218 0 1
rlabel polysilicon 303 -224 303 -224 0 3
rlabel polysilicon 310 -218 310 -218 0 1
rlabel polysilicon 310 -224 310 -224 0 3
rlabel polysilicon 320 -224 320 -224 0 4
rlabel polysilicon 324 -218 324 -218 0 1
rlabel polysilicon 327 -218 327 -218 0 2
rlabel polysilicon 327 -224 327 -224 0 4
rlabel polysilicon 331 -218 331 -218 0 1
rlabel polysilicon 334 -224 334 -224 0 4
rlabel polysilicon 341 -218 341 -218 0 2
rlabel polysilicon 345 -218 345 -218 0 1
rlabel polysilicon 345 -224 345 -224 0 3
rlabel polysilicon 352 -218 352 -218 0 1
rlabel polysilicon 355 -224 355 -224 0 4
rlabel polysilicon 359 -218 359 -218 0 1
rlabel polysilicon 359 -224 359 -224 0 3
rlabel polysilicon 366 -218 366 -218 0 1
rlabel polysilicon 366 -224 366 -224 0 3
rlabel polysilicon 373 -218 373 -218 0 1
rlabel polysilicon 373 -224 373 -224 0 3
rlabel polysilicon 380 -218 380 -218 0 1
rlabel polysilicon 380 -224 380 -224 0 3
rlabel polysilicon 390 -218 390 -218 0 2
rlabel polysilicon 387 -224 387 -224 0 3
rlabel polysilicon 9 -247 9 -247 0 1
rlabel polysilicon 9 -253 9 -253 0 3
rlabel polysilicon 16 -247 16 -247 0 1
rlabel polysilicon 16 -253 16 -253 0 3
rlabel polysilicon 23 -247 23 -247 0 1
rlabel polysilicon 23 -253 23 -253 0 3
rlabel polysilicon 33 -247 33 -247 0 2
rlabel polysilicon 33 -253 33 -253 0 4
rlabel polysilicon 37 -247 37 -247 0 1
rlabel polysilicon 44 -247 44 -247 0 1
rlabel polysilicon 44 -253 44 -253 0 3
rlabel polysilicon 54 -247 54 -247 0 2
rlabel polysilicon 51 -253 51 -253 0 3
rlabel polysilicon 58 -247 58 -247 0 1
rlabel polysilicon 58 -253 58 -253 0 3
rlabel polysilicon 65 -247 65 -247 0 1
rlabel polysilicon 65 -253 65 -253 0 3
rlabel polysilicon 72 -247 72 -247 0 1
rlabel polysilicon 72 -253 72 -253 0 3
rlabel polysilicon 79 -247 79 -247 0 1
rlabel polysilicon 79 -253 79 -253 0 3
rlabel polysilicon 86 -247 86 -247 0 1
rlabel polysilicon 86 -253 86 -253 0 3
rlabel polysilicon 89 -253 89 -253 0 4
rlabel polysilicon 93 -247 93 -247 0 1
rlabel polysilicon 93 -253 93 -253 0 3
rlabel polysilicon 100 -247 100 -247 0 1
rlabel polysilicon 100 -253 100 -253 0 3
rlabel polysilicon 107 -247 107 -247 0 1
rlabel polysilicon 110 -247 110 -247 0 2
rlabel polysilicon 107 -253 107 -253 0 3
rlabel polysilicon 114 -247 114 -247 0 1
rlabel polysilicon 114 -253 114 -253 0 3
rlabel polysilicon 121 -247 121 -247 0 1
rlabel polysilicon 121 -253 121 -253 0 3
rlabel polysilicon 131 -253 131 -253 0 4
rlabel polysilicon 135 -247 135 -247 0 1
rlabel polysilicon 135 -253 135 -253 0 3
rlabel polysilicon 142 -253 142 -253 0 3
rlabel polysilicon 145 -253 145 -253 0 4
rlabel polysilicon 149 -247 149 -247 0 1
rlabel polysilicon 152 -247 152 -247 0 2
rlabel polysilicon 149 -253 149 -253 0 3
rlabel polysilicon 156 -247 156 -247 0 1
rlabel polysilicon 156 -253 156 -253 0 3
rlabel polysilicon 163 -247 163 -247 0 1
rlabel polysilicon 163 -253 163 -253 0 3
rlabel polysilicon 170 -247 170 -247 0 1
rlabel polysilicon 173 -247 173 -247 0 2
rlabel polysilicon 170 -253 170 -253 0 3
rlabel polysilicon 173 -253 173 -253 0 4
rlabel polysilicon 177 -247 177 -247 0 1
rlabel polysilicon 177 -253 177 -253 0 3
rlabel polysilicon 184 -247 184 -247 0 1
rlabel polysilicon 184 -253 184 -253 0 3
rlabel polysilicon 191 -247 191 -247 0 1
rlabel polysilicon 191 -253 191 -253 0 3
rlabel polysilicon 198 -247 198 -247 0 1
rlabel polysilicon 198 -253 198 -253 0 3
rlabel polysilicon 208 -247 208 -247 0 2
rlabel polysilicon 205 -253 205 -253 0 3
rlabel polysilicon 212 -247 212 -247 0 1
rlabel polysilicon 212 -253 212 -253 0 3
rlabel polysilicon 222 -247 222 -247 0 2
rlabel polysilicon 219 -253 219 -253 0 3
rlabel polysilicon 222 -253 222 -253 0 4
rlabel polysilicon 226 -247 226 -247 0 1
rlabel polysilicon 226 -253 226 -253 0 3
rlabel polysilicon 233 -247 233 -247 0 1
rlabel polysilicon 233 -253 233 -253 0 3
rlabel polysilicon 240 -247 240 -247 0 1
rlabel polysilicon 240 -253 240 -253 0 3
rlabel polysilicon 247 -247 247 -247 0 1
rlabel polysilicon 247 -253 247 -253 0 3
rlabel polysilicon 254 -247 254 -247 0 1
rlabel polysilicon 254 -253 254 -253 0 3
rlabel polysilicon 261 -247 261 -247 0 1
rlabel polysilicon 261 -253 261 -253 0 3
rlabel polysilicon 268 -247 268 -247 0 1
rlabel polysilicon 268 -253 268 -253 0 3
rlabel polysilicon 275 -247 275 -247 0 1
rlabel polysilicon 275 -253 275 -253 0 3
rlabel polysilicon 282 -247 282 -247 0 1
rlabel polysilicon 282 -253 282 -253 0 3
rlabel polysilicon 289 -247 289 -247 0 1
rlabel polysilicon 289 -253 289 -253 0 3
rlabel polysilicon 296 -247 296 -247 0 1
rlabel polysilicon 296 -253 296 -253 0 3
rlabel polysilicon 303 -247 303 -247 0 1
rlabel polysilicon 303 -253 303 -253 0 3
rlabel polysilicon 310 -247 310 -247 0 1
rlabel polysilicon 310 -253 310 -253 0 3
rlabel polysilicon 317 -247 317 -247 0 1
rlabel polysilicon 317 -253 317 -253 0 3
rlabel polysilicon 327 -247 327 -247 0 2
rlabel polysilicon 331 -247 331 -247 0 1
rlabel polysilicon 331 -253 331 -253 0 3
rlabel polysilicon 338 -247 338 -247 0 1
rlabel polysilicon 345 -253 345 -253 0 3
rlabel polysilicon 352 -247 352 -247 0 1
rlabel polysilicon 352 -253 352 -253 0 3
rlabel polysilicon 380 -247 380 -247 0 1
rlabel polysilicon 387 -253 387 -253 0 3
rlabel polysilicon 394 -247 394 -247 0 1
rlabel polysilicon 394 -253 394 -253 0 3
rlabel polysilicon 2 -294 2 -294 0 1
rlabel polysilicon 2 -300 2 -300 0 3
rlabel polysilicon 9 -294 9 -294 0 1
rlabel polysilicon 16 -294 16 -294 0 1
rlabel polysilicon 16 -300 16 -300 0 3
rlabel polysilicon 23 -294 23 -294 0 1
rlabel polysilicon 23 -300 23 -300 0 3
rlabel polysilicon 30 -300 30 -300 0 3
rlabel polysilicon 37 -294 37 -294 0 1
rlabel polysilicon 37 -300 37 -300 0 3
rlabel polysilicon 44 -294 44 -294 0 1
rlabel polysilicon 44 -300 44 -300 0 3
rlabel polysilicon 54 -294 54 -294 0 2
rlabel polysilicon 51 -300 51 -300 0 3
rlabel polysilicon 58 -294 58 -294 0 1
rlabel polysilicon 58 -300 58 -300 0 3
rlabel polysilicon 65 -294 65 -294 0 1
rlabel polysilicon 68 -294 68 -294 0 2
rlabel polysilicon 65 -300 65 -300 0 3
rlabel polysilicon 72 -294 72 -294 0 1
rlabel polysilicon 75 -294 75 -294 0 2
rlabel polysilicon 79 -294 79 -294 0 1
rlabel polysilicon 82 -294 82 -294 0 2
rlabel polysilicon 79 -300 79 -300 0 3
rlabel polysilicon 86 -294 86 -294 0 1
rlabel polysilicon 86 -300 86 -300 0 3
rlabel polysilicon 96 -294 96 -294 0 2
rlabel polysilicon 96 -300 96 -300 0 4
rlabel polysilicon 100 -294 100 -294 0 1
rlabel polysilicon 100 -300 100 -300 0 3
rlabel polysilicon 107 -294 107 -294 0 1
rlabel polysilicon 107 -300 107 -300 0 3
rlabel polysilicon 114 -294 114 -294 0 1
rlabel polysilicon 117 -300 117 -300 0 4
rlabel polysilicon 121 -294 121 -294 0 1
rlabel polysilicon 121 -300 121 -300 0 3
rlabel polysilicon 128 -294 128 -294 0 1
rlabel polysilicon 131 -300 131 -300 0 4
rlabel polysilicon 135 -294 135 -294 0 1
rlabel polysilicon 135 -300 135 -300 0 3
rlabel polysilicon 142 -294 142 -294 0 1
rlabel polysilicon 142 -300 142 -300 0 3
rlabel polysilicon 149 -294 149 -294 0 1
rlabel polysilicon 152 -294 152 -294 0 2
rlabel polysilicon 149 -300 149 -300 0 3
rlabel polysilicon 156 -294 156 -294 0 1
rlabel polysilicon 159 -294 159 -294 0 2
rlabel polysilicon 156 -300 156 -300 0 3
rlabel polysilicon 163 -294 163 -294 0 1
rlabel polysilicon 163 -300 163 -300 0 3
rlabel polysilicon 170 -294 170 -294 0 1
rlabel polysilicon 170 -300 170 -300 0 3
rlabel polysilicon 173 -300 173 -300 0 4
rlabel polysilicon 177 -294 177 -294 0 1
rlabel polysilicon 180 -294 180 -294 0 2
rlabel polysilicon 177 -300 177 -300 0 3
rlabel polysilicon 187 -294 187 -294 0 2
rlabel polysilicon 184 -300 184 -300 0 3
rlabel polysilicon 187 -300 187 -300 0 4
rlabel polysilicon 191 -294 191 -294 0 1
rlabel polysilicon 194 -294 194 -294 0 2
rlabel polysilicon 191 -300 191 -300 0 3
rlabel polysilicon 194 -300 194 -300 0 4
rlabel polysilicon 198 -294 198 -294 0 1
rlabel polysilicon 198 -300 198 -300 0 3
rlabel polysilicon 208 -294 208 -294 0 2
rlabel polysilicon 205 -300 205 -300 0 3
rlabel polysilicon 208 -300 208 -300 0 4
rlabel polysilicon 212 -294 212 -294 0 1
rlabel polysilicon 215 -294 215 -294 0 2
rlabel polysilicon 212 -300 212 -300 0 3
rlabel polysilicon 215 -300 215 -300 0 4
rlabel polysilicon 219 -294 219 -294 0 1
rlabel polysilicon 219 -300 219 -300 0 3
rlabel polysilicon 226 -294 226 -294 0 1
rlabel polysilicon 226 -300 226 -300 0 3
rlabel polysilicon 233 -294 233 -294 0 1
rlabel polysilicon 243 -294 243 -294 0 2
rlabel polysilicon 243 -300 243 -300 0 4
rlabel polysilicon 247 -294 247 -294 0 1
rlabel polysilicon 247 -300 247 -300 0 3
rlabel polysilicon 254 -294 254 -294 0 1
rlabel polysilicon 254 -300 254 -300 0 3
rlabel polysilicon 261 -294 261 -294 0 1
rlabel polysilicon 261 -300 261 -300 0 3
rlabel polysilicon 268 -294 268 -294 0 1
rlabel polysilicon 268 -300 268 -300 0 3
rlabel polysilicon 275 -294 275 -294 0 1
rlabel polysilicon 275 -300 275 -300 0 3
rlabel polysilicon 282 -294 282 -294 0 1
rlabel polysilicon 282 -300 282 -300 0 3
rlabel polysilicon 289 -294 289 -294 0 1
rlabel polysilicon 289 -300 289 -300 0 3
rlabel polysilicon 296 -294 296 -294 0 1
rlabel polysilicon 296 -300 296 -300 0 3
rlabel polysilicon 303 -294 303 -294 0 1
rlabel polysilicon 303 -300 303 -300 0 3
rlabel polysilicon 310 -294 310 -294 0 1
rlabel polysilicon 310 -300 310 -300 0 3
rlabel polysilicon 317 -294 317 -294 0 1
rlabel polysilicon 317 -300 317 -300 0 3
rlabel polysilicon 324 -294 324 -294 0 1
rlabel polysilicon 324 -300 324 -300 0 3
rlabel polysilicon 331 -294 331 -294 0 1
rlabel polysilicon 331 -300 331 -300 0 3
rlabel polysilicon 338 -294 338 -294 0 1
rlabel polysilicon 338 -300 338 -300 0 3
rlabel polysilicon 345 -294 345 -294 0 1
rlabel polysilicon 345 -300 345 -300 0 3
rlabel polysilicon 30 -341 30 -341 0 1
rlabel polysilicon 30 -347 30 -347 0 3
rlabel polysilicon 37 -341 37 -341 0 1
rlabel polysilicon 37 -347 37 -347 0 3
rlabel polysilicon 44 -341 44 -341 0 1
rlabel polysilicon 44 -347 44 -347 0 3
rlabel polysilicon 54 -341 54 -341 0 2
rlabel polysilicon 58 -341 58 -341 0 1
rlabel polysilicon 58 -347 58 -347 0 3
rlabel polysilicon 65 -341 65 -341 0 1
rlabel polysilicon 65 -347 65 -347 0 3
rlabel polysilicon 75 -341 75 -341 0 2
rlabel polysilicon 79 -341 79 -341 0 1
rlabel polysilicon 79 -347 79 -347 0 3
rlabel polysilicon 86 -341 86 -341 0 1
rlabel polysilicon 86 -347 86 -347 0 3
rlabel polysilicon 93 -341 93 -341 0 1
rlabel polysilicon 93 -347 93 -347 0 3
rlabel polysilicon 103 -341 103 -341 0 2
rlabel polysilicon 103 -347 103 -347 0 4
rlabel polysilicon 110 -341 110 -341 0 2
rlabel polysilicon 107 -347 107 -347 0 3
rlabel polysilicon 114 -341 114 -341 0 1
rlabel polysilicon 117 -347 117 -347 0 4
rlabel polysilicon 121 -341 121 -341 0 1
rlabel polysilicon 128 -341 128 -341 0 1
rlabel polysilicon 128 -347 128 -347 0 3
rlabel polysilicon 135 -341 135 -341 0 1
rlabel polysilicon 138 -341 138 -341 0 2
rlabel polysilicon 135 -347 135 -347 0 3
rlabel polysilicon 142 -341 142 -341 0 1
rlabel polysilicon 145 -341 145 -341 0 2
rlabel polysilicon 145 -347 145 -347 0 4
rlabel polysilicon 149 -341 149 -341 0 1
rlabel polysilicon 152 -341 152 -341 0 2
rlabel polysilicon 152 -347 152 -347 0 4
rlabel polysilicon 156 -341 156 -341 0 1
rlabel polysilicon 163 -341 163 -341 0 1
rlabel polysilicon 163 -347 163 -347 0 3
rlabel polysilicon 170 -341 170 -341 0 1
rlabel polysilicon 170 -347 170 -347 0 3
rlabel polysilicon 177 -341 177 -341 0 1
rlabel polysilicon 177 -347 177 -347 0 3
rlabel polysilicon 184 -341 184 -341 0 1
rlabel polysilicon 187 -341 187 -341 0 2
rlabel polysilicon 184 -347 184 -347 0 3
rlabel polysilicon 191 -347 191 -347 0 3
rlabel polysilicon 194 -347 194 -347 0 4
rlabel polysilicon 198 -341 198 -341 0 1
rlabel polysilicon 201 -341 201 -341 0 2
rlabel polysilicon 201 -347 201 -347 0 4
rlabel polysilicon 208 -341 208 -341 0 2
rlabel polysilicon 205 -347 205 -347 0 3
rlabel polysilicon 212 -341 212 -341 0 1
rlabel polysilicon 215 -341 215 -341 0 2
rlabel polysilicon 212 -347 212 -347 0 3
rlabel polysilicon 219 -341 219 -341 0 1
rlabel polysilicon 219 -347 219 -347 0 3
rlabel polysilicon 229 -341 229 -341 0 2
rlabel polysilicon 233 -341 233 -341 0 1
rlabel polysilicon 233 -347 233 -347 0 3
rlabel polysilicon 240 -341 240 -341 0 1
rlabel polysilicon 243 -347 243 -347 0 4
rlabel polysilicon 247 -341 247 -341 0 1
rlabel polysilicon 247 -347 247 -347 0 3
rlabel polysilicon 254 -341 254 -341 0 1
rlabel polysilicon 254 -347 254 -347 0 3
rlabel polysilicon 261 -341 261 -341 0 1
rlabel polysilicon 261 -347 261 -347 0 3
rlabel polysilicon 268 -341 268 -341 0 1
rlabel polysilicon 268 -347 268 -347 0 3
rlabel polysilicon 275 -341 275 -341 0 1
rlabel polysilicon 275 -347 275 -347 0 3
rlabel polysilicon 282 -341 282 -341 0 1
rlabel polysilicon 282 -347 282 -347 0 3
rlabel polysilicon 289 -341 289 -341 0 1
rlabel polysilicon 289 -347 289 -347 0 3
rlabel polysilicon 296 -341 296 -341 0 1
rlabel polysilicon 299 -347 299 -347 0 4
rlabel polysilicon 303 -341 303 -341 0 1
rlabel polysilicon 303 -347 303 -347 0 3
rlabel polysilicon 310 -341 310 -341 0 1
rlabel polysilicon 310 -347 310 -347 0 3
rlabel polysilicon 317 -341 317 -341 0 1
rlabel polysilicon 317 -347 317 -347 0 3
rlabel polysilicon 324 -341 324 -341 0 1
rlabel polysilicon 324 -347 324 -347 0 3
rlabel polysilicon 2 -376 2 -376 0 1
rlabel polysilicon 2 -382 2 -382 0 3
rlabel polysilicon 9 -376 9 -376 0 1
rlabel polysilicon 9 -382 9 -382 0 3
rlabel polysilicon 16 -376 16 -376 0 1
rlabel polysilicon 16 -382 16 -382 0 3
rlabel polysilicon 23 -376 23 -376 0 1
rlabel polysilicon 23 -382 23 -382 0 3
rlabel polysilicon 30 -382 30 -382 0 3
rlabel polysilicon 37 -376 37 -376 0 1
rlabel polysilicon 37 -382 37 -382 0 3
rlabel polysilicon 44 -376 44 -376 0 1
rlabel polysilicon 44 -382 44 -382 0 3
rlabel polysilicon 51 -376 51 -376 0 1
rlabel polysilicon 51 -382 51 -382 0 3
rlabel polysilicon 58 -382 58 -382 0 3
rlabel polysilicon 61 -382 61 -382 0 4
rlabel polysilicon 65 -376 65 -376 0 1
rlabel polysilicon 68 -382 68 -382 0 4
rlabel polysilicon 72 -376 72 -376 0 1
rlabel polysilicon 75 -376 75 -376 0 2
rlabel polysilicon 75 -382 75 -382 0 4
rlabel polysilicon 79 -376 79 -376 0 1
rlabel polysilicon 79 -382 79 -382 0 3
rlabel polysilicon 86 -376 86 -376 0 1
rlabel polysilicon 89 -376 89 -376 0 2
rlabel polysilicon 89 -382 89 -382 0 4
rlabel polysilicon 93 -376 93 -376 0 1
rlabel polysilicon 96 -376 96 -376 0 2
rlabel polysilicon 93 -382 93 -382 0 3
rlabel polysilicon 100 -376 100 -376 0 1
rlabel polysilicon 100 -382 100 -382 0 3
rlabel polysilicon 107 -376 107 -376 0 1
rlabel polysilicon 107 -382 107 -382 0 3
rlabel polysilicon 114 -376 114 -376 0 1
rlabel polysilicon 117 -376 117 -376 0 2
rlabel polysilicon 114 -382 114 -382 0 3
rlabel polysilicon 117 -382 117 -382 0 4
rlabel polysilicon 121 -376 121 -376 0 1
rlabel polysilicon 121 -382 121 -382 0 3
rlabel polysilicon 128 -376 128 -376 0 1
rlabel polysilicon 128 -382 128 -382 0 3
rlabel polysilicon 135 -376 135 -376 0 1
rlabel polysilicon 138 -382 138 -382 0 4
rlabel polysilicon 142 -376 142 -376 0 1
rlabel polysilicon 145 -376 145 -376 0 2
rlabel polysilicon 142 -382 142 -382 0 3
rlabel polysilicon 149 -376 149 -376 0 1
rlabel polysilicon 149 -382 149 -382 0 3
rlabel polysilicon 156 -382 156 -382 0 3
rlabel polysilicon 163 -376 163 -376 0 1
rlabel polysilicon 166 -376 166 -376 0 2
rlabel polysilicon 166 -382 166 -382 0 4
rlabel polysilicon 170 -376 170 -376 0 1
rlabel polysilicon 173 -376 173 -376 0 2
rlabel polysilicon 170 -382 170 -382 0 3
rlabel polysilicon 180 -376 180 -376 0 2
rlabel polysilicon 177 -382 177 -382 0 3
rlabel polysilicon 180 -382 180 -382 0 4
rlabel polysilicon 184 -382 184 -382 0 3
rlabel polysilicon 191 -376 191 -376 0 1
rlabel polysilicon 191 -382 191 -382 0 3
rlabel polysilicon 194 -382 194 -382 0 4
rlabel polysilicon 198 -376 198 -376 0 1
rlabel polysilicon 198 -382 198 -382 0 3
rlabel polysilicon 205 -376 205 -376 0 1
rlabel polysilicon 205 -382 205 -382 0 3
rlabel polysilicon 212 -376 212 -376 0 1
rlabel polysilicon 215 -376 215 -376 0 2
rlabel polysilicon 215 -382 215 -382 0 4
rlabel polysilicon 219 -376 219 -376 0 1
rlabel polysilicon 219 -382 219 -382 0 3
rlabel polysilicon 226 -376 226 -376 0 1
rlabel polysilicon 226 -382 226 -382 0 3
rlabel polysilicon 233 -376 233 -376 0 1
rlabel polysilicon 233 -382 233 -382 0 3
rlabel polysilicon 240 -376 240 -376 0 1
rlabel polysilicon 240 -382 240 -382 0 3
rlabel polysilicon 247 -376 247 -376 0 1
rlabel polysilicon 247 -382 247 -382 0 3
rlabel polysilicon 254 -376 254 -376 0 1
rlabel polysilicon 254 -382 254 -382 0 3
rlabel polysilicon 264 -376 264 -376 0 2
rlabel polysilicon 261 -382 261 -382 0 3
rlabel polysilicon 268 -376 268 -376 0 1
rlabel polysilicon 268 -382 268 -382 0 3
rlabel polysilicon 275 -376 275 -376 0 1
rlabel polysilicon 275 -382 275 -382 0 3
rlabel polysilicon 282 -376 282 -376 0 1
rlabel polysilicon 282 -382 282 -382 0 3
rlabel polysilicon 289 -376 289 -376 0 1
rlabel polysilicon 289 -382 289 -382 0 3
rlabel polysilicon 296 -376 296 -376 0 1
rlabel polysilicon 296 -382 296 -382 0 3
rlabel polysilicon 306 -382 306 -382 0 4
rlabel polysilicon 310 -376 310 -376 0 1
rlabel polysilicon 310 -382 310 -382 0 3
rlabel polysilicon 317 -376 317 -376 0 1
rlabel polysilicon 317 -382 317 -382 0 3
rlabel polysilicon 324 -376 324 -376 0 1
rlabel polysilicon 324 -382 324 -382 0 3
rlabel polysilicon 331 -376 331 -376 0 1
rlabel polysilicon 331 -382 331 -382 0 3
rlabel polysilicon 338 -376 338 -376 0 1
rlabel polysilicon 338 -382 338 -382 0 3
rlabel polysilicon 345 -376 345 -376 0 1
rlabel polysilicon 345 -382 345 -382 0 3
rlabel polysilicon 23 -417 23 -417 0 1
rlabel polysilicon 23 -423 23 -423 0 3
rlabel polysilicon 30 -417 30 -417 0 1
rlabel polysilicon 30 -423 30 -423 0 3
rlabel polysilicon 40 -417 40 -417 0 2
rlabel polysilicon 37 -423 37 -423 0 3
rlabel polysilicon 44 -417 44 -417 0 1
rlabel polysilicon 44 -423 44 -423 0 3
rlabel polysilicon 51 -417 51 -417 0 1
rlabel polysilicon 54 -417 54 -417 0 2
rlabel polysilicon 54 -423 54 -423 0 4
rlabel polysilicon 58 -417 58 -417 0 1
rlabel polysilicon 58 -423 58 -423 0 3
rlabel polysilicon 65 -417 65 -417 0 1
rlabel polysilicon 65 -423 65 -423 0 3
rlabel polysilicon 75 -417 75 -417 0 2
rlabel polysilicon 72 -423 72 -423 0 3
rlabel polysilicon 79 -417 79 -417 0 1
rlabel polysilicon 82 -417 82 -417 0 2
rlabel polysilicon 86 -417 86 -417 0 1
rlabel polysilicon 86 -423 86 -423 0 3
rlabel polysilicon 96 -417 96 -417 0 2
rlabel polysilicon 93 -423 93 -423 0 3
rlabel polysilicon 96 -423 96 -423 0 4
rlabel polysilicon 103 -417 103 -417 0 2
rlabel polysilicon 107 -417 107 -417 0 1
rlabel polysilicon 107 -423 107 -423 0 3
rlabel polysilicon 128 -417 128 -417 0 1
rlabel polysilicon 128 -423 128 -423 0 3
rlabel polysilicon 135 -417 135 -417 0 1
rlabel polysilicon 135 -423 135 -423 0 3
rlabel polysilicon 142 -417 142 -417 0 1
rlabel polysilicon 142 -423 142 -423 0 3
rlabel polysilicon 149 -417 149 -417 0 1
rlabel polysilicon 152 -417 152 -417 0 2
rlabel polysilicon 156 -417 156 -417 0 1
rlabel polysilicon 156 -423 156 -423 0 3
rlabel polysilicon 163 -417 163 -417 0 1
rlabel polysilicon 163 -423 163 -423 0 3
rlabel polysilicon 170 -423 170 -423 0 3
rlabel polysilicon 173 -423 173 -423 0 4
rlabel polysilicon 177 -417 177 -417 0 1
rlabel polysilicon 177 -423 177 -423 0 3
rlabel polysilicon 184 -417 184 -417 0 1
rlabel polysilicon 184 -423 184 -423 0 3
rlabel polysilicon 191 -417 191 -417 0 1
rlabel polysilicon 191 -423 191 -423 0 3
rlabel polysilicon 198 -417 198 -417 0 1
rlabel polysilicon 201 -417 201 -417 0 2
rlabel polysilicon 201 -423 201 -423 0 4
rlabel polysilicon 205 -417 205 -417 0 1
rlabel polysilicon 205 -423 205 -423 0 3
rlabel polysilicon 212 -417 212 -417 0 1
rlabel polysilicon 215 -417 215 -417 0 2
rlabel polysilicon 219 -417 219 -417 0 1
rlabel polysilicon 219 -423 219 -423 0 3
rlabel polysilicon 222 -423 222 -423 0 4
rlabel polysilicon 226 -417 226 -417 0 1
rlabel polysilicon 226 -423 226 -423 0 3
rlabel polysilicon 229 -423 229 -423 0 4
rlabel polysilicon 233 -417 233 -417 0 1
rlabel polysilicon 233 -423 233 -423 0 3
rlabel polysilicon 243 -417 243 -417 0 2
rlabel polysilicon 247 -417 247 -417 0 1
rlabel polysilicon 247 -423 247 -423 0 3
rlabel polysilicon 254 -417 254 -417 0 1
rlabel polysilicon 254 -423 254 -423 0 3
rlabel polysilicon 261 -417 261 -417 0 1
rlabel polysilicon 261 -423 261 -423 0 3
rlabel polysilicon 268 -417 268 -417 0 1
rlabel polysilicon 271 -417 271 -417 0 2
rlabel polysilicon 268 -423 268 -423 0 3
rlabel polysilicon 275 -417 275 -417 0 1
rlabel polysilicon 275 -423 275 -423 0 3
rlabel polysilicon 282 -417 282 -417 0 1
rlabel polysilicon 285 -417 285 -417 0 2
rlabel polysilicon 282 -423 282 -423 0 3
rlabel polysilicon 289 -417 289 -417 0 1
rlabel polysilicon 292 -417 292 -417 0 2
rlabel polysilicon 296 -417 296 -417 0 1
rlabel polysilicon 296 -423 296 -423 0 3
rlabel polysilicon 303 -417 303 -417 0 1
rlabel polysilicon 303 -423 303 -423 0 3
rlabel polysilicon 310 -417 310 -417 0 1
rlabel polysilicon 310 -423 310 -423 0 3
rlabel polysilicon 317 -417 317 -417 0 1
rlabel polysilicon 317 -423 317 -423 0 3
rlabel polysilicon 2 -448 2 -448 0 1
rlabel polysilicon 2 -454 2 -454 0 3
rlabel polysilicon 9 -448 9 -448 0 1
rlabel polysilicon 9 -454 9 -454 0 3
rlabel polysilicon 16 -448 16 -448 0 1
rlabel polysilicon 16 -454 16 -454 0 3
rlabel polysilicon 23 -448 23 -448 0 1
rlabel polysilicon 23 -454 23 -454 0 3
rlabel polysilicon 30 -448 30 -448 0 1
rlabel polysilicon 30 -454 30 -454 0 3
rlabel polysilicon 37 -448 37 -448 0 1
rlabel polysilicon 37 -454 37 -454 0 3
rlabel polysilicon 47 -448 47 -448 0 2
rlabel polysilicon 44 -454 44 -454 0 3
rlabel polysilicon 51 -448 51 -448 0 1
rlabel polysilicon 51 -454 51 -454 0 3
rlabel polysilicon 58 -448 58 -448 0 1
rlabel polysilicon 58 -454 58 -454 0 3
rlabel polysilicon 61 -454 61 -454 0 4
rlabel polysilicon 65 -448 65 -448 0 1
rlabel polysilicon 65 -454 65 -454 0 3
rlabel polysilicon 72 -448 72 -448 0 1
rlabel polysilicon 75 -454 75 -454 0 4
rlabel polysilicon 79 -448 79 -448 0 1
rlabel polysilicon 82 -448 82 -448 0 2
rlabel polysilicon 79 -454 79 -454 0 3
rlabel polysilicon 89 -448 89 -448 0 2
rlabel polysilicon 86 -454 86 -454 0 3
rlabel polysilicon 89 -454 89 -454 0 4
rlabel polysilicon 93 -448 93 -448 0 1
rlabel polysilicon 93 -454 93 -454 0 3
rlabel polysilicon 103 -448 103 -448 0 2
rlabel polysilicon 100 -454 100 -454 0 3
rlabel polysilicon 103 -454 103 -454 0 4
rlabel polysilicon 107 -448 107 -448 0 1
rlabel polysilicon 110 -448 110 -448 0 2
rlabel polysilicon 110 -454 110 -454 0 4
rlabel polysilicon 114 -448 114 -448 0 1
rlabel polysilicon 114 -454 114 -454 0 3
rlabel polysilicon 121 -448 121 -448 0 1
rlabel polysilicon 121 -454 121 -454 0 3
rlabel polysilicon 128 -448 128 -448 0 1
rlabel polysilicon 131 -448 131 -448 0 2
rlabel polysilicon 128 -454 128 -454 0 3
rlabel polysilicon 135 -448 135 -448 0 1
rlabel polysilicon 135 -454 135 -454 0 3
rlabel polysilicon 138 -454 138 -454 0 4
rlabel polysilicon 142 -448 142 -448 0 1
rlabel polysilicon 142 -454 142 -454 0 3
rlabel polysilicon 149 -448 149 -448 0 1
rlabel polysilicon 149 -454 149 -454 0 3
rlabel polysilicon 156 -448 156 -448 0 1
rlabel polysilicon 159 -454 159 -454 0 4
rlabel polysilicon 163 -448 163 -448 0 1
rlabel polysilicon 163 -454 163 -454 0 3
rlabel polysilicon 170 -448 170 -448 0 1
rlabel polysilicon 173 -454 173 -454 0 4
rlabel polysilicon 177 -448 177 -448 0 1
rlabel polysilicon 177 -454 177 -454 0 3
rlabel polysilicon 184 -448 184 -448 0 1
rlabel polysilicon 184 -454 184 -454 0 3
rlabel polysilicon 191 -448 191 -448 0 1
rlabel polysilicon 194 -448 194 -448 0 2
rlabel polysilicon 194 -454 194 -454 0 4
rlabel polysilicon 201 -448 201 -448 0 2
rlabel polysilicon 205 -448 205 -448 0 1
rlabel polysilicon 205 -454 205 -454 0 3
rlabel polysilicon 212 -448 212 -448 0 1
rlabel polysilicon 212 -454 212 -454 0 3
rlabel polysilicon 215 -454 215 -454 0 4
rlabel polysilicon 219 -448 219 -448 0 1
rlabel polysilicon 219 -454 219 -454 0 3
rlabel polysilicon 226 -448 226 -448 0 1
rlabel polysilicon 226 -454 226 -454 0 3
rlabel polysilicon 233 -448 233 -448 0 1
rlabel polysilicon 233 -454 233 -454 0 3
rlabel polysilicon 236 -454 236 -454 0 4
rlabel polysilicon 240 -448 240 -448 0 1
rlabel polysilicon 240 -454 240 -454 0 3
rlabel polysilicon 247 -448 247 -448 0 1
rlabel polysilicon 247 -454 247 -454 0 3
rlabel polysilicon 254 -448 254 -448 0 1
rlabel polysilicon 254 -454 254 -454 0 3
rlabel polysilicon 261 -448 261 -448 0 1
rlabel polysilicon 261 -454 261 -454 0 3
rlabel polysilicon 268 -448 268 -448 0 1
rlabel polysilicon 268 -454 268 -454 0 3
rlabel polysilicon 275 -448 275 -448 0 1
rlabel polysilicon 275 -454 275 -454 0 3
rlabel polysilicon 282 -448 282 -448 0 1
rlabel polysilicon 282 -454 282 -454 0 3
rlabel polysilicon 289 -448 289 -448 0 1
rlabel polysilicon 289 -454 289 -454 0 3
rlabel polysilicon 296 -448 296 -448 0 1
rlabel polysilicon 296 -454 296 -454 0 3
rlabel polysilicon 303 -448 303 -448 0 1
rlabel polysilicon 303 -454 303 -454 0 3
rlabel polysilicon 310 -448 310 -448 0 1
rlabel polysilicon 310 -454 310 -454 0 3
rlabel polysilicon 317 -448 317 -448 0 1
rlabel polysilicon 317 -454 317 -454 0 3
rlabel polysilicon 324 -448 324 -448 0 1
rlabel polysilicon 327 -448 327 -448 0 2
rlabel polysilicon 327 -454 327 -454 0 4
rlabel polysilicon 334 -454 334 -454 0 4
rlabel polysilicon 338 -448 338 -448 0 1
rlabel polysilicon 338 -454 338 -454 0 3
rlabel polysilicon 40 -489 40 -489 0 2
rlabel polysilicon 44 -489 44 -489 0 1
rlabel polysilicon 44 -495 44 -495 0 3
rlabel polysilicon 51 -489 51 -489 0 1
rlabel polysilicon 51 -495 51 -495 0 3
rlabel polysilicon 58 -489 58 -489 0 1
rlabel polysilicon 58 -495 58 -495 0 3
rlabel polysilicon 65 -489 65 -489 0 1
rlabel polysilicon 65 -495 65 -495 0 3
rlabel polysilicon 75 -489 75 -489 0 2
rlabel polysilicon 72 -495 72 -495 0 3
rlabel polysilicon 82 -495 82 -495 0 4
rlabel polysilicon 86 -489 86 -489 0 1
rlabel polysilicon 86 -495 86 -495 0 3
rlabel polysilicon 93 -489 93 -489 0 1
rlabel polysilicon 93 -495 93 -495 0 3
rlabel polysilicon 100 -489 100 -489 0 1
rlabel polysilicon 100 -495 100 -495 0 3
rlabel polysilicon 107 -489 107 -489 0 1
rlabel polysilicon 107 -495 107 -495 0 3
rlabel polysilicon 114 -489 114 -489 0 1
rlabel polysilicon 114 -495 114 -495 0 3
rlabel polysilicon 121 -489 121 -489 0 1
rlabel polysilicon 124 -495 124 -495 0 4
rlabel polysilicon 128 -489 128 -489 0 1
rlabel polysilicon 131 -489 131 -489 0 2
rlabel polysilicon 128 -495 128 -495 0 3
rlabel polysilicon 138 -489 138 -489 0 2
rlabel polysilicon 138 -495 138 -495 0 4
rlabel polysilicon 142 -489 142 -489 0 1
rlabel polysilicon 145 -489 145 -489 0 2
rlabel polysilicon 145 -495 145 -495 0 4
rlabel polysilicon 149 -489 149 -489 0 1
rlabel polysilicon 149 -495 149 -495 0 3
rlabel polysilicon 156 -489 156 -489 0 1
rlabel polysilicon 156 -495 156 -495 0 3
rlabel polysilicon 163 -489 163 -489 0 1
rlabel polysilicon 163 -495 163 -495 0 3
rlabel polysilicon 170 -489 170 -489 0 1
rlabel polysilicon 170 -495 170 -495 0 3
rlabel polysilicon 177 -489 177 -489 0 1
rlabel polysilicon 180 -489 180 -489 0 2
rlabel polysilicon 180 -495 180 -495 0 4
rlabel polysilicon 184 -489 184 -489 0 1
rlabel polysilicon 184 -495 184 -495 0 3
rlabel polysilicon 191 -489 191 -489 0 1
rlabel polysilicon 191 -495 191 -495 0 3
rlabel polysilicon 198 -489 198 -489 0 1
rlabel polysilicon 198 -495 198 -495 0 3
rlabel polysilicon 201 -495 201 -495 0 4
rlabel polysilicon 205 -489 205 -489 0 1
rlabel polysilicon 205 -495 205 -495 0 3
rlabel polysilicon 215 -489 215 -489 0 2
rlabel polysilicon 219 -489 219 -489 0 1
rlabel polysilicon 222 -489 222 -489 0 2
rlabel polysilicon 222 -495 222 -495 0 4
rlabel polysilicon 226 -489 226 -489 0 1
rlabel polysilicon 226 -495 226 -495 0 3
rlabel polysilicon 233 -489 233 -489 0 1
rlabel polysilicon 233 -495 233 -495 0 3
rlabel polysilicon 240 -489 240 -489 0 1
rlabel polysilicon 240 -495 240 -495 0 3
rlabel polysilicon 247 -489 247 -489 0 1
rlabel polysilicon 247 -495 247 -495 0 3
rlabel polysilicon 254 -495 254 -495 0 3
rlabel polysilicon 257 -495 257 -495 0 4
rlabel polysilicon 261 -489 261 -489 0 1
rlabel polysilicon 261 -495 261 -495 0 3
rlabel polysilicon 268 -489 268 -489 0 1
rlabel polysilicon 268 -495 268 -495 0 3
rlabel polysilicon 275 -489 275 -489 0 1
rlabel polysilicon 275 -495 275 -495 0 3
rlabel polysilicon 282 -495 282 -495 0 3
rlabel polysilicon 289 -489 289 -489 0 1
rlabel polysilicon 289 -495 289 -495 0 3
rlabel polysilicon 296 -489 296 -489 0 1
rlabel polysilicon 296 -495 296 -495 0 3
rlabel polysilicon 303 -489 303 -489 0 1
rlabel polysilicon 303 -495 303 -495 0 3
rlabel polysilicon 310 -489 310 -489 0 1
rlabel polysilicon 310 -495 310 -495 0 3
rlabel polysilicon 317 -489 317 -489 0 1
rlabel polysilicon 320 -489 320 -489 0 2
rlabel polysilicon 320 -495 320 -495 0 4
rlabel polysilicon 327 -495 327 -495 0 4
rlabel polysilicon 331 -489 331 -489 0 1
rlabel polysilicon 331 -495 331 -495 0 3
rlabel polysilicon 338 -489 338 -489 0 1
rlabel polysilicon 338 -495 338 -495 0 3
rlabel polysilicon 348 -495 348 -495 0 4
rlabel polysilicon 352 -489 352 -489 0 1
rlabel polysilicon 352 -495 352 -495 0 3
rlabel polysilicon 359 -489 359 -489 0 1
rlabel polysilicon 359 -495 359 -495 0 3
rlabel polysilicon 366 -489 366 -489 0 1
rlabel polysilicon 16 -526 16 -526 0 1
rlabel polysilicon 16 -532 16 -532 0 3
rlabel polysilicon 23 -526 23 -526 0 1
rlabel polysilicon 23 -532 23 -532 0 3
rlabel polysilicon 30 -526 30 -526 0 1
rlabel polysilicon 30 -532 30 -532 0 3
rlabel polysilicon 37 -532 37 -532 0 3
rlabel polysilicon 44 -526 44 -526 0 1
rlabel polysilicon 44 -532 44 -532 0 3
rlabel polysilicon 51 -526 51 -526 0 1
rlabel polysilicon 51 -532 51 -532 0 3
rlabel polysilicon 61 -526 61 -526 0 2
rlabel polysilicon 58 -532 58 -532 0 3
rlabel polysilicon 61 -532 61 -532 0 4
rlabel polysilicon 65 -526 65 -526 0 1
rlabel polysilicon 65 -532 65 -532 0 3
rlabel polysilicon 72 -526 72 -526 0 1
rlabel polysilicon 72 -532 72 -532 0 3
rlabel polysilicon 79 -526 79 -526 0 1
rlabel polysilicon 82 -526 82 -526 0 2
rlabel polysilicon 82 -532 82 -532 0 4
rlabel polysilicon 86 -526 86 -526 0 1
rlabel polysilicon 86 -532 86 -532 0 3
rlabel polysilicon 93 -526 93 -526 0 1
rlabel polysilicon 93 -532 93 -532 0 3
rlabel polysilicon 100 -526 100 -526 0 1
rlabel polysilicon 103 -526 103 -526 0 2
rlabel polysilicon 103 -532 103 -532 0 4
rlabel polysilicon 107 -526 107 -526 0 1
rlabel polysilicon 107 -532 107 -532 0 3
rlabel polysilicon 114 -526 114 -526 0 1
rlabel polysilicon 114 -532 114 -532 0 3
rlabel polysilicon 121 -526 121 -526 0 1
rlabel polysilicon 124 -532 124 -532 0 4
rlabel polysilicon 128 -526 128 -526 0 1
rlabel polysilicon 128 -532 128 -532 0 3
rlabel polysilicon 135 -526 135 -526 0 1
rlabel polysilicon 135 -532 135 -532 0 3
rlabel polysilicon 138 -532 138 -532 0 4
rlabel polysilicon 142 -526 142 -526 0 1
rlabel polysilicon 142 -532 142 -532 0 3
rlabel polysilicon 149 -526 149 -526 0 1
rlabel polysilicon 149 -532 149 -532 0 3
rlabel polysilicon 156 -526 156 -526 0 1
rlabel polysilicon 159 -526 159 -526 0 2
rlabel polysilicon 156 -532 156 -532 0 3
rlabel polysilicon 159 -532 159 -532 0 4
rlabel polysilicon 163 -526 163 -526 0 1
rlabel polysilicon 166 -526 166 -526 0 2
rlabel polysilicon 163 -532 163 -532 0 3
rlabel polysilicon 166 -532 166 -532 0 4
rlabel polysilicon 170 -526 170 -526 0 1
rlabel polysilicon 170 -532 170 -532 0 3
rlabel polysilicon 177 -526 177 -526 0 1
rlabel polysilicon 180 -526 180 -526 0 2
rlabel polysilicon 180 -532 180 -532 0 4
rlabel polysilicon 184 -526 184 -526 0 1
rlabel polysilicon 184 -532 184 -532 0 3
rlabel polysilicon 194 -526 194 -526 0 2
rlabel polysilicon 191 -532 191 -532 0 3
rlabel polysilicon 194 -532 194 -532 0 4
rlabel polysilicon 198 -526 198 -526 0 1
rlabel polysilicon 201 -526 201 -526 0 2
rlabel polysilicon 201 -532 201 -532 0 4
rlabel polysilicon 205 -526 205 -526 0 1
rlabel polysilicon 208 -532 208 -532 0 4
rlabel polysilicon 212 -526 212 -526 0 1
rlabel polysilicon 212 -532 212 -532 0 3
rlabel polysilicon 215 -532 215 -532 0 4
rlabel polysilicon 219 -526 219 -526 0 1
rlabel polysilicon 219 -532 219 -532 0 3
rlabel polysilicon 226 -526 226 -526 0 1
rlabel polysilicon 229 -526 229 -526 0 2
rlabel polysilicon 233 -526 233 -526 0 1
rlabel polysilicon 233 -532 233 -532 0 3
rlabel polysilicon 240 -526 240 -526 0 1
rlabel polysilicon 240 -532 240 -532 0 3
rlabel polysilicon 247 -526 247 -526 0 1
rlabel polysilicon 247 -532 247 -532 0 3
rlabel polysilicon 254 -526 254 -526 0 1
rlabel polysilicon 254 -532 254 -532 0 3
rlabel polysilicon 261 -526 261 -526 0 1
rlabel polysilicon 261 -532 261 -532 0 3
rlabel polysilicon 271 -526 271 -526 0 2
rlabel polysilicon 268 -532 268 -532 0 3
rlabel polysilicon 271 -532 271 -532 0 4
rlabel polysilicon 275 -526 275 -526 0 1
rlabel polysilicon 275 -532 275 -532 0 3
rlabel polysilicon 282 -526 282 -526 0 1
rlabel polysilicon 282 -532 282 -532 0 3
rlabel polysilicon 289 -526 289 -526 0 1
rlabel polysilicon 289 -532 289 -532 0 3
rlabel polysilicon 296 -526 296 -526 0 1
rlabel polysilicon 296 -532 296 -532 0 3
rlabel polysilicon 303 -526 303 -526 0 1
rlabel polysilicon 303 -532 303 -532 0 3
rlabel polysilicon 310 -526 310 -526 0 1
rlabel polysilicon 310 -532 310 -532 0 3
rlabel polysilicon 317 -526 317 -526 0 1
rlabel polysilicon 317 -532 317 -532 0 3
rlabel polysilicon 324 -526 324 -526 0 1
rlabel polysilicon 324 -532 324 -532 0 3
rlabel polysilicon 331 -526 331 -526 0 1
rlabel polysilicon 331 -532 331 -532 0 3
rlabel polysilicon 338 -526 338 -526 0 1
rlabel polysilicon 338 -532 338 -532 0 3
rlabel polysilicon 345 -526 345 -526 0 1
rlabel polysilicon 345 -532 345 -532 0 3
rlabel polysilicon 352 -526 352 -526 0 1
rlabel polysilicon 352 -532 352 -532 0 3
rlabel polysilicon 9 -569 9 -569 0 1
rlabel polysilicon 9 -575 9 -575 0 3
rlabel polysilicon 16 -569 16 -569 0 1
rlabel polysilicon 16 -575 16 -575 0 3
rlabel polysilicon 23 -569 23 -569 0 1
rlabel polysilicon 23 -575 23 -575 0 3
rlabel polysilicon 33 -569 33 -569 0 2
rlabel polysilicon 40 -569 40 -569 0 2
rlabel polysilicon 44 -575 44 -575 0 3
rlabel polysilicon 51 -569 51 -569 0 1
rlabel polysilicon 51 -575 51 -575 0 3
rlabel polysilicon 58 -569 58 -569 0 1
rlabel polysilicon 61 -569 61 -569 0 2
rlabel polysilicon 61 -575 61 -575 0 4
rlabel polysilicon 65 -569 65 -569 0 1
rlabel polysilicon 68 -569 68 -569 0 2
rlabel polysilicon 72 -569 72 -569 0 1
rlabel polysilicon 72 -575 72 -575 0 3
rlabel polysilicon 82 -569 82 -569 0 2
rlabel polysilicon 79 -575 79 -575 0 3
rlabel polysilicon 86 -569 86 -569 0 1
rlabel polysilicon 86 -575 86 -575 0 3
rlabel polysilicon 93 -569 93 -569 0 1
rlabel polysilicon 93 -575 93 -575 0 3
rlabel polysilicon 100 -569 100 -569 0 1
rlabel polysilicon 100 -575 100 -575 0 3
rlabel polysilicon 107 -569 107 -569 0 1
rlabel polysilicon 117 -569 117 -569 0 2
rlabel polysilicon 114 -575 114 -575 0 3
rlabel polysilicon 121 -569 121 -569 0 1
rlabel polysilicon 121 -575 121 -575 0 3
rlabel polysilicon 128 -569 128 -569 0 1
rlabel polysilicon 128 -575 128 -575 0 3
rlabel polysilicon 135 -569 135 -569 0 1
rlabel polysilicon 135 -575 135 -575 0 3
rlabel polysilicon 142 -569 142 -569 0 1
rlabel polysilicon 142 -575 142 -575 0 3
rlabel polysilicon 149 -575 149 -575 0 3
rlabel polysilicon 156 -569 156 -569 0 1
rlabel polysilicon 156 -575 156 -575 0 3
rlabel polysilicon 163 -569 163 -569 0 1
rlabel polysilicon 166 -569 166 -569 0 2
rlabel polysilicon 163 -575 163 -575 0 3
rlabel polysilicon 170 -569 170 -569 0 1
rlabel polysilicon 170 -575 170 -575 0 3
rlabel polysilicon 177 -569 177 -569 0 1
rlabel polysilicon 177 -575 177 -575 0 3
rlabel polysilicon 180 -575 180 -575 0 4
rlabel polysilicon 184 -569 184 -569 0 1
rlabel polysilicon 184 -575 184 -575 0 3
rlabel polysilicon 191 -569 191 -569 0 1
rlabel polysilicon 191 -575 191 -575 0 3
rlabel polysilicon 198 -569 198 -569 0 1
rlabel polysilicon 198 -575 198 -575 0 3
rlabel polysilicon 205 -569 205 -569 0 1
rlabel polysilicon 205 -575 205 -575 0 3
rlabel polysilicon 212 -569 212 -569 0 1
rlabel polysilicon 212 -575 212 -575 0 3
rlabel polysilicon 219 -569 219 -569 0 1
rlabel polysilicon 222 -569 222 -569 0 2
rlabel polysilicon 219 -575 219 -575 0 3
rlabel polysilicon 222 -575 222 -575 0 4
rlabel polysilicon 226 -569 226 -569 0 1
rlabel polysilicon 226 -575 226 -575 0 3
rlabel polysilicon 233 -569 233 -569 0 1
rlabel polysilicon 233 -575 233 -575 0 3
rlabel polysilicon 236 -575 236 -575 0 4
rlabel polysilicon 243 -569 243 -569 0 2
rlabel polysilicon 240 -575 240 -575 0 3
rlabel polysilicon 243 -575 243 -575 0 4
rlabel polysilicon 247 -569 247 -569 0 1
rlabel polysilicon 250 -569 250 -569 0 2
rlabel polysilicon 250 -575 250 -575 0 4
rlabel polysilicon 254 -569 254 -569 0 1
rlabel polysilicon 254 -575 254 -575 0 3
rlabel polysilicon 261 -569 261 -569 0 1
rlabel polysilicon 261 -575 261 -575 0 3
rlabel polysilicon 268 -569 268 -569 0 1
rlabel polysilicon 268 -575 268 -575 0 3
rlabel polysilicon 275 -569 275 -569 0 1
rlabel polysilicon 275 -575 275 -575 0 3
rlabel polysilicon 282 -569 282 -569 0 1
rlabel polysilicon 282 -575 282 -575 0 3
rlabel polysilicon 289 -569 289 -569 0 1
rlabel polysilicon 289 -575 289 -575 0 3
rlabel polysilicon 296 -569 296 -569 0 1
rlabel polysilicon 296 -575 296 -575 0 3
rlabel polysilicon 303 -569 303 -569 0 1
rlabel polysilicon 303 -575 303 -575 0 3
rlabel polysilicon 310 -569 310 -569 0 1
rlabel polysilicon 310 -575 310 -575 0 3
rlabel polysilicon 317 -569 317 -569 0 1
rlabel polysilicon 317 -575 317 -575 0 3
rlabel polysilicon 324 -569 324 -569 0 1
rlabel polysilicon 324 -575 324 -575 0 3
rlabel polysilicon 331 -569 331 -569 0 1
rlabel polysilicon 331 -575 331 -575 0 3
rlabel polysilicon 338 -569 338 -569 0 1
rlabel polysilicon 338 -575 338 -575 0 3
rlabel polysilicon 345 -569 345 -569 0 1
rlabel polysilicon 345 -575 345 -575 0 3
rlabel polysilicon 352 -569 352 -569 0 1
rlabel polysilicon 352 -575 352 -575 0 3
rlabel polysilicon 362 -569 362 -569 0 2
rlabel polysilicon 359 -575 359 -575 0 3
rlabel polysilicon 369 -569 369 -569 0 2
rlabel polysilicon 369 -575 369 -575 0 4
rlabel polysilicon 44 -606 44 -606 0 1
rlabel polysilicon 47 -606 47 -606 0 2
rlabel polysilicon 51 -606 51 -606 0 1
rlabel polysilicon 51 -612 51 -612 0 3
rlabel polysilicon 68 -606 68 -606 0 2
rlabel polysilicon 68 -612 68 -612 0 4
rlabel polysilicon 72 -606 72 -606 0 1
rlabel polysilicon 72 -612 72 -612 0 3
rlabel polysilicon 79 -606 79 -606 0 1
rlabel polysilicon 86 -606 86 -606 0 1
rlabel polysilicon 86 -612 86 -612 0 3
rlabel polysilicon 93 -606 93 -606 0 1
rlabel polysilicon 93 -612 93 -612 0 3
rlabel polysilicon 100 -606 100 -606 0 1
rlabel polysilicon 103 -606 103 -606 0 2
rlabel polysilicon 110 -606 110 -606 0 2
rlabel polysilicon 110 -612 110 -612 0 4
rlabel polysilicon 114 -606 114 -606 0 1
rlabel polysilicon 114 -612 114 -612 0 3
rlabel polysilicon 121 -606 121 -606 0 1
rlabel polysilicon 121 -612 121 -612 0 3
rlabel polysilicon 124 -612 124 -612 0 4
rlabel polysilicon 128 -606 128 -606 0 1
rlabel polysilicon 128 -612 128 -612 0 3
rlabel polysilicon 135 -606 135 -606 0 1
rlabel polysilicon 135 -612 135 -612 0 3
rlabel polysilicon 145 -606 145 -606 0 2
rlabel polysilicon 142 -612 142 -612 0 3
rlabel polysilicon 149 -606 149 -606 0 1
rlabel polysilicon 152 -606 152 -606 0 2
rlabel polysilicon 156 -606 156 -606 0 1
rlabel polysilicon 156 -612 156 -612 0 3
rlabel polysilicon 163 -606 163 -606 0 1
rlabel polysilicon 163 -612 163 -612 0 3
rlabel polysilicon 166 -612 166 -612 0 4
rlabel polysilicon 170 -606 170 -606 0 1
rlabel polysilicon 170 -612 170 -612 0 3
rlabel polysilicon 177 -606 177 -606 0 1
rlabel polysilicon 177 -612 177 -612 0 3
rlabel polysilicon 187 -606 187 -606 0 2
rlabel polysilicon 184 -612 184 -612 0 3
rlabel polysilicon 187 -612 187 -612 0 4
rlabel polysilicon 191 -606 191 -606 0 1
rlabel polysilicon 191 -612 191 -612 0 3
rlabel polysilicon 194 -612 194 -612 0 4
rlabel polysilicon 198 -606 198 -606 0 1
rlabel polysilicon 198 -612 198 -612 0 3
rlabel polysilicon 205 -606 205 -606 0 1
rlabel polysilicon 205 -612 205 -612 0 3
rlabel polysilicon 212 -606 212 -606 0 1
rlabel polysilicon 212 -612 212 -612 0 3
rlabel polysilicon 219 -606 219 -606 0 1
rlabel polysilicon 219 -612 219 -612 0 3
rlabel polysilicon 229 -606 229 -606 0 2
rlabel polysilicon 233 -606 233 -606 0 1
rlabel polysilicon 233 -612 233 -612 0 3
rlabel polysilicon 240 -606 240 -606 0 1
rlabel polysilicon 240 -612 240 -612 0 3
rlabel polysilicon 247 -606 247 -606 0 1
rlabel polysilicon 250 -606 250 -606 0 2
rlabel polysilicon 250 -612 250 -612 0 4
rlabel polysilicon 254 -606 254 -606 0 1
rlabel polysilicon 257 -606 257 -606 0 2
rlabel polysilicon 257 -612 257 -612 0 4
rlabel polysilicon 261 -606 261 -606 0 1
rlabel polysilicon 264 -606 264 -606 0 2
rlabel polysilicon 268 -606 268 -606 0 1
rlabel polysilicon 268 -612 268 -612 0 3
rlabel polysilicon 275 -606 275 -606 0 1
rlabel polysilicon 275 -612 275 -612 0 3
rlabel polysilicon 282 -606 282 -606 0 1
rlabel polysilicon 282 -612 282 -612 0 3
rlabel polysilicon 292 -606 292 -606 0 2
rlabel polysilicon 289 -612 289 -612 0 3
rlabel polysilicon 310 -606 310 -606 0 1
rlabel polysilicon 310 -612 310 -612 0 3
rlabel polysilicon 44 -643 44 -643 0 3
rlabel polysilicon 51 -637 51 -637 0 1
rlabel polysilicon 51 -643 51 -643 0 3
rlabel polysilicon 58 -637 58 -637 0 1
rlabel polysilicon 58 -643 58 -643 0 3
rlabel polysilicon 65 -637 65 -637 0 1
rlabel polysilicon 68 -637 68 -637 0 2
rlabel polysilicon 65 -643 65 -643 0 3
rlabel polysilicon 72 -637 72 -637 0 1
rlabel polysilicon 72 -643 72 -643 0 3
rlabel polysilicon 79 -637 79 -637 0 1
rlabel polysilicon 79 -643 79 -643 0 3
rlabel polysilicon 82 -643 82 -643 0 4
rlabel polysilicon 86 -637 86 -637 0 1
rlabel polysilicon 86 -643 86 -643 0 3
rlabel polysilicon 96 -637 96 -637 0 2
rlabel polysilicon 93 -643 93 -643 0 3
rlabel polysilicon 96 -643 96 -643 0 4
rlabel polysilicon 100 -637 100 -637 0 1
rlabel polysilicon 103 -637 103 -637 0 2
rlabel polysilicon 107 -637 107 -637 0 1
rlabel polysilicon 107 -643 107 -643 0 3
rlabel polysilicon 114 -637 114 -637 0 1
rlabel polysilicon 114 -643 114 -643 0 3
rlabel polysilicon 124 -643 124 -643 0 4
rlabel polysilicon 128 -637 128 -637 0 1
rlabel polysilicon 128 -643 128 -643 0 3
rlabel polysilicon 138 -637 138 -637 0 2
rlabel polysilicon 142 -637 142 -637 0 1
rlabel polysilicon 142 -643 142 -643 0 3
rlabel polysilicon 149 -643 149 -643 0 3
rlabel polysilicon 152 -643 152 -643 0 4
rlabel polysilicon 156 -637 156 -637 0 1
rlabel polysilicon 156 -643 156 -643 0 3
rlabel polysilicon 163 -637 163 -637 0 1
rlabel polysilicon 163 -643 163 -643 0 3
rlabel polysilicon 170 -637 170 -637 0 1
rlabel polysilicon 173 -643 173 -643 0 4
rlabel polysilicon 177 -637 177 -637 0 1
rlabel polysilicon 180 -643 180 -643 0 4
rlabel polysilicon 184 -637 184 -637 0 1
rlabel polysilicon 184 -643 184 -643 0 3
rlabel polysilicon 191 -643 191 -643 0 3
rlabel polysilicon 194 -643 194 -643 0 4
rlabel polysilicon 198 -637 198 -637 0 1
rlabel polysilicon 198 -643 198 -643 0 3
rlabel polysilicon 208 -637 208 -637 0 2
rlabel polysilicon 208 -643 208 -643 0 4
rlabel polysilicon 212 -637 212 -637 0 1
rlabel polysilicon 212 -643 212 -643 0 3
rlabel polysilicon 219 -637 219 -637 0 1
rlabel polysilicon 219 -643 219 -643 0 3
rlabel polysilicon 226 -637 226 -637 0 1
rlabel polysilicon 226 -643 226 -643 0 3
rlabel polysilicon 233 -637 233 -637 0 1
rlabel polysilicon 233 -643 233 -643 0 3
rlabel polysilicon 240 -637 240 -637 0 1
rlabel polysilicon 240 -643 240 -643 0 3
rlabel polysilicon 247 -637 247 -637 0 1
rlabel polysilicon 247 -643 247 -643 0 3
rlabel polysilicon 254 -637 254 -637 0 1
rlabel polysilicon 254 -643 254 -643 0 3
rlabel polysilicon 261 -637 261 -637 0 1
rlabel polysilicon 261 -643 261 -643 0 3
rlabel polysilicon 268 -637 268 -637 0 1
rlabel polysilicon 268 -643 268 -643 0 3
rlabel polysilicon 275 -637 275 -637 0 1
rlabel polysilicon 275 -643 275 -643 0 3
rlabel polysilicon 282 -637 282 -637 0 1
rlabel polysilicon 282 -643 282 -643 0 3
rlabel polysilicon 289 -637 289 -637 0 1
rlabel polysilicon 292 -637 292 -637 0 2
rlabel polysilicon 299 -637 299 -637 0 2
rlabel polysilicon 303 -637 303 -637 0 1
rlabel polysilicon 303 -643 303 -643 0 3
rlabel polysilicon 313 -637 313 -637 0 2
rlabel polysilicon 310 -643 310 -643 0 3
rlabel polysilicon 44 -664 44 -664 0 1
rlabel polysilicon 44 -670 44 -670 0 3
rlabel polysilicon 54 -664 54 -664 0 2
rlabel polysilicon 58 -670 58 -670 0 3
rlabel polysilicon 65 -664 65 -664 0 1
rlabel polysilicon 65 -670 65 -670 0 3
rlabel polysilicon 72 -664 72 -664 0 1
rlabel polysilicon 72 -670 72 -670 0 3
rlabel polysilicon 79 -664 79 -664 0 1
rlabel polysilicon 79 -670 79 -670 0 3
rlabel polysilicon 89 -664 89 -664 0 2
rlabel polysilicon 86 -670 86 -670 0 3
rlabel polysilicon 93 -670 93 -670 0 3
rlabel polysilicon 96 -670 96 -670 0 4
rlabel polysilicon 100 -664 100 -664 0 1
rlabel polysilicon 100 -670 100 -670 0 3
rlabel polysilicon 107 -664 107 -664 0 1
rlabel polysilicon 107 -670 107 -670 0 3
rlabel polysilicon 114 -664 114 -664 0 1
rlabel polysilicon 114 -670 114 -670 0 3
rlabel polysilicon 121 -664 121 -664 0 1
rlabel polysilicon 124 -670 124 -670 0 4
rlabel polysilicon 135 -664 135 -664 0 1
rlabel polysilicon 138 -670 138 -670 0 4
rlabel polysilicon 142 -664 142 -664 0 1
rlabel polysilicon 149 -664 149 -664 0 1
rlabel polysilicon 149 -670 149 -670 0 3
rlabel polysilicon 170 -664 170 -664 0 1
rlabel polysilicon 170 -670 170 -670 0 3
rlabel polysilicon 180 -670 180 -670 0 4
rlabel polysilicon 184 -664 184 -664 0 1
rlabel polysilicon 184 -670 184 -670 0 3
rlabel polysilicon 191 -664 191 -664 0 1
rlabel polysilicon 191 -670 191 -670 0 3
rlabel polysilicon 201 -664 201 -664 0 2
rlabel polysilicon 201 -670 201 -670 0 4
rlabel polysilicon 205 -664 205 -664 0 1
rlabel polysilicon 205 -670 205 -670 0 3
rlabel polysilicon 212 -664 212 -664 0 1
rlabel polysilicon 222 -664 222 -664 0 2
rlabel polysilicon 219 -670 219 -670 0 3
rlabel polysilicon 226 -664 226 -664 0 1
rlabel polysilicon 226 -670 226 -670 0 3
rlabel polysilicon 233 -664 233 -664 0 1
rlabel polysilicon 233 -670 233 -670 0 3
rlabel polysilicon 240 -664 240 -664 0 1
rlabel polysilicon 243 -664 243 -664 0 2
rlabel polysilicon 240 -670 240 -670 0 3
rlabel polysilicon 243 -670 243 -670 0 4
rlabel polysilicon 254 -664 254 -664 0 1
rlabel polysilicon 254 -670 254 -670 0 3
rlabel polysilicon 261 -664 261 -664 0 1
rlabel polysilicon 264 -664 264 -664 0 2
rlabel polysilicon 268 -664 268 -664 0 1
rlabel polysilicon 268 -670 268 -670 0 3
rlabel polysilicon 278 -664 278 -664 0 2
rlabel polysilicon 282 -664 282 -664 0 1
rlabel polysilicon 285 -670 285 -670 0 4
rlabel polysilicon 292 -664 292 -664 0 2
rlabel polysilicon 292 -670 292 -670 0 4
rlabel polysilicon 44 -685 44 -685 0 3
rlabel polysilicon 51 -679 51 -679 0 1
rlabel polysilicon 51 -685 51 -685 0 3
rlabel polysilicon 58 -679 58 -679 0 1
rlabel polysilicon 58 -685 58 -685 0 3
rlabel polysilicon 65 -679 65 -679 0 1
rlabel polysilicon 72 -679 72 -679 0 1
rlabel polysilicon 72 -685 72 -685 0 3
rlabel polysilicon 79 -679 79 -679 0 1
rlabel polysilicon 79 -685 79 -685 0 3
rlabel polysilicon 86 -685 86 -685 0 3
rlabel polysilicon 93 -685 93 -685 0 3
rlabel polysilicon 103 -679 103 -679 0 2
rlabel polysilicon 107 -685 107 -685 0 3
rlabel polysilicon 114 -685 114 -685 0 3
rlabel polysilicon 117 -685 117 -685 0 4
rlabel polysilicon 121 -679 121 -679 0 1
rlabel polysilicon 121 -685 121 -685 0 3
rlabel polysilicon 128 -679 128 -679 0 1
rlabel polysilicon 128 -685 128 -685 0 3
rlabel polysilicon 135 -679 135 -679 0 1
rlabel polysilicon 135 -685 135 -685 0 3
rlabel polysilicon 145 -679 145 -679 0 2
rlabel polysilicon 142 -685 142 -685 0 3
rlabel polysilicon 145 -685 145 -685 0 4
rlabel polysilicon 152 -685 152 -685 0 4
rlabel polysilicon 191 -679 191 -679 0 1
rlabel polysilicon 201 -679 201 -679 0 2
rlabel polysilicon 198 -685 198 -685 0 3
rlabel polysilicon 205 -679 205 -679 0 1
rlabel polysilicon 205 -685 205 -685 0 3
rlabel polysilicon 212 -679 212 -679 0 1
rlabel polysilicon 212 -685 212 -685 0 3
rlabel polysilicon 222 -685 222 -685 0 4
rlabel polysilicon 226 -679 226 -679 0 1
rlabel polysilicon 226 -685 226 -685 0 3
rlabel polysilicon 233 -685 233 -685 0 3
rlabel polysilicon 240 -679 240 -679 0 1
rlabel polysilicon 243 -685 243 -685 0 4
rlabel polysilicon 247 -679 247 -679 0 1
rlabel polysilicon 247 -685 247 -685 0 3
rlabel polysilicon 254 -679 254 -679 0 1
rlabel polysilicon 254 -685 254 -685 0 3
rlabel polysilicon 264 -685 264 -685 0 4
rlabel polysilicon 275 -679 275 -679 0 1
rlabel polysilicon 275 -685 275 -685 0 3
rlabel polysilicon 285 -685 285 -685 0 4
rlabel metal2 135 1 135 1 0 net=689
rlabel metal2 142 -1 142 -1 0 net=881
rlabel metal2 100 -12 100 -12 0 net=777
rlabel metal2 121 -12 121 -12 0 net=753
rlabel metal2 177 -12 177 -12 0 net=136
rlabel metal2 128 -14 128 -14 0 net=1207
rlabel metal2 177 -14 177 -14 0 net=1213
rlabel metal2 135 -16 135 -16 0 net=690
rlabel metal2 149 -16 149 -16 0 net=882
rlabel metal2 135 -18 135 -18 0 net=623
rlabel metal2 152 -18 152 -18 0 net=727
rlabel metal2 79 -29 79 -29 0 net=373
rlabel metal2 128 -29 128 -29 0 net=625
rlabel metal2 142 -29 142 -29 0 net=41
rlabel metal2 159 -29 159 -29 0 net=1131
rlabel metal2 86 -31 86 -31 0 net=1073
rlabel metal2 170 -31 170 -31 0 net=1209
rlabel metal2 93 -33 93 -33 0 net=693
rlabel metal2 121 -33 121 -33 0 net=563
rlabel metal2 170 -33 170 -33 0 net=1215
rlabel metal2 191 -33 191 -33 0 net=1107
rlabel metal2 100 -35 100 -35 0 net=778
rlabel metal2 135 -35 135 -35 0 net=509
rlabel metal2 163 -35 163 -35 0 net=755
rlabel metal2 194 -35 194 -35 0 net=1141
rlabel metal2 156 -37 156 -37 0 net=729
rlabel metal2 180 -37 180 -37 0 net=965
rlabel metal2 79 -48 79 -48 0 net=374
rlabel metal2 114 -48 114 -48 0 net=564
rlabel metal2 128 -48 128 -48 0 net=627
rlabel metal2 180 -48 180 -48 0 net=1132
rlabel metal2 222 -48 222 -48 0 net=983
rlabel metal2 79 -50 79 -50 0 net=893
rlabel metal2 145 -50 145 -50 0 net=966
rlabel metal2 86 -52 86 -52 0 net=1074
rlabel metal2 114 -52 114 -52 0 net=511
rlabel metal2 145 -52 145 -52 0 net=1210
rlabel metal2 86 -54 86 -54 0 net=695
rlabel metal2 100 -54 100 -54 0 net=479
rlabel metal2 156 -54 156 -54 0 net=756
rlabel metal2 191 -54 191 -54 0 net=907
rlabel metal2 93 -56 93 -56 0 net=603
rlabel metal2 170 -56 170 -56 0 net=1217
rlabel metal2 131 -58 131 -58 0 net=117
rlabel metal2 149 -58 149 -58 0 net=1108
rlabel metal2 110 -60 110 -60 0 net=337
rlabel metal2 163 -60 163 -60 0 net=731
rlabel metal2 187 -60 187 -60 0 net=947
rlabel metal2 198 -60 198 -60 0 net=1143
rlabel metal2 149 -62 149 -62 0 net=791
rlabel metal2 72 -73 72 -73 0 net=829
rlabel metal2 135 -73 135 -73 0 net=326
rlabel metal2 159 -73 159 -73 0 net=1218
rlabel metal2 233 -73 233 -73 0 net=985
rlabel metal2 233 -73 233 -73 0 net=985
rlabel metal2 243 -73 243 -73 0 net=651
rlabel metal2 79 -75 79 -75 0 net=894
rlabel metal2 138 -75 138 -75 0 net=628
rlabel metal2 184 -75 184 -75 0 net=819
rlabel metal2 205 -75 205 -75 0 net=908
rlabel metal2 222 -75 222 -75 0 net=451
rlabel metal2 261 -75 261 -75 0 net=1325
rlabel metal2 79 -77 79 -77 0 net=605
rlabel metal2 121 -77 121 -77 0 net=101
rlabel metal2 138 -77 138 -77 0 net=1144
rlabel metal2 86 -79 86 -79 0 net=696
rlabel metal2 142 -79 142 -79 0 net=873
rlabel metal2 65 -81 65 -81 0 net=379
rlabel metal2 93 -81 93 -81 0 net=186
rlabel metal2 152 -81 152 -81 0 net=1127
rlabel metal2 205 -81 205 -81 0 net=1249
rlabel metal2 100 -83 100 -83 0 net=481
rlabel metal2 156 -83 156 -83 0 net=499
rlabel metal2 100 -85 100 -85 0 net=795
rlabel metal2 163 -85 163 -85 0 net=793
rlabel metal2 191 -85 191 -85 0 net=949
rlabel metal2 114 -87 114 -87 0 net=513
rlabel metal2 114 -89 114 -89 0 net=733
rlabel metal2 170 -91 170 -91 0 net=785
rlabel metal2 44 -102 44 -102 0 net=613
rlabel metal2 65 -102 65 -102 0 net=380
rlabel metal2 142 -102 142 -102 0 net=794
rlabel metal2 198 -102 198 -102 0 net=1128
rlabel metal2 233 -102 233 -102 0 net=987
rlabel metal2 233 -102 233 -102 0 net=987
rlabel metal2 254 -102 254 -102 0 net=452
rlabel metal2 268 -102 268 -102 0 net=652
rlabel metal2 299 -102 299 -102 0 net=1111
rlabel metal2 65 -104 65 -104 0 net=1313
rlabel metal2 79 -104 79 -104 0 net=606
rlabel metal2 131 -104 131 -104 0 net=501
rlabel metal2 149 -104 149 -104 0 net=500
rlabel metal2 159 -104 159 -104 0 net=48
rlabel metal2 247 -104 247 -104 0 net=1251
rlabel metal2 282 -104 282 -104 0 net=1327
rlabel metal2 72 -106 72 -106 0 net=830
rlabel metal2 205 -106 205 -106 0 net=1289
rlabel metal2 86 -108 86 -108 0 net=725
rlabel metal2 100 -108 100 -108 0 net=797
rlabel metal2 117 -108 117 -108 0 net=635
rlabel metal2 152 -108 152 -108 0 net=514
rlabel metal2 170 -108 170 -108 0 net=821
rlabel metal2 212 -108 212 -108 0 net=875
rlabel metal2 93 -110 93 -110 0 net=1175
rlabel metal2 138 -110 138 -110 0 net=1339
rlabel metal2 212 -110 212 -110 0 net=823
rlabel metal2 226 -110 226 -110 0 net=951
rlabel metal2 100 -112 100 -112 0 net=483
rlabel metal2 156 -112 156 -112 0 net=1097
rlabel metal2 114 -114 114 -114 0 net=735
rlabel metal2 163 -114 163 -114 0 net=683
rlabel metal2 219 -114 219 -114 0 net=1135
rlabel metal2 58 -116 58 -116 0 net=1319
rlabel metal2 177 -116 177 -116 0 net=579
rlabel metal2 191 -116 191 -116 0 net=787
rlabel metal2 19 -127 19 -127 0 net=485
rlabel metal2 30 -127 30 -127 0 net=21
rlabel metal2 47 -127 47 -127 0 net=614
rlabel metal2 58 -127 58 -127 0 net=1320
rlabel metal2 100 -127 100 -127 0 net=484
rlabel metal2 135 -127 135 -127 0 net=581
rlabel metal2 184 -127 184 -127 0 net=824
rlabel metal2 240 -127 240 -127 0 net=877
rlabel metal2 289 -127 289 -127 0 net=1328
rlabel metal2 310 -127 310 -127 0 net=1295
rlabel metal2 331 -127 331 -127 0 net=1231
rlabel metal2 58 -129 58 -129 0 net=531
rlabel metal2 79 -129 79 -129 0 net=726
rlabel metal2 107 -129 107 -129 0 net=798
rlabel metal2 142 -129 142 -129 0 net=503
rlabel metal2 142 -129 142 -129 0 net=503
rlabel metal2 149 -129 149 -129 0 net=636
rlabel metal2 159 -129 159 -129 0 net=822
rlabel metal2 177 -129 177 -129 0 net=1252
rlabel metal2 271 -129 271 -129 0 net=1105
rlabel metal2 296 -129 296 -129 0 net=1113
rlabel metal2 324 -129 324 -129 0 net=937
rlabel metal2 65 -131 65 -131 0 net=1314
rlabel metal2 93 -131 93 -131 0 net=1176
rlabel metal2 121 -131 121 -131 0 net=736
rlabel metal2 156 -131 156 -131 0 net=637
rlabel metal2 254 -131 254 -131 0 net=1099
rlabel metal2 275 -131 275 -131 0 net=1137
rlabel metal2 37 -133 37 -133 0 net=443
rlabel metal2 68 -133 68 -133 0 net=963
rlabel metal2 93 -133 93 -133 0 net=437
rlabel metal2 107 -133 107 -133 0 net=617
rlabel metal2 191 -133 191 -133 0 net=988
rlabel metal2 236 -133 236 -133 0 net=1259
rlabel metal2 79 -135 79 -135 0 net=769
rlabel metal2 198 -135 198 -135 0 net=1290
rlabel metal2 121 -137 121 -137 0 net=701
rlabel metal2 163 -137 163 -137 0 net=685
rlabel metal2 247 -137 247 -137 0 net=953
rlabel metal2 163 -139 163 -139 0 net=493
rlabel metal2 201 -139 201 -139 0 net=1083
rlabel metal2 170 -141 170 -141 0 net=469
rlabel metal2 205 -141 205 -141 0 net=1341
rlabel metal2 194 -143 194 -143 0 net=565
rlabel metal2 226 -143 226 -143 0 net=789
rlabel metal2 131 -145 131 -145 0 net=629
rlabel metal2 19 -156 19 -156 0 net=486
rlabel metal2 37 -156 37 -156 0 net=444
rlabel metal2 72 -156 72 -156 0 net=619
rlabel metal2 114 -156 114 -156 0 net=50
rlabel metal2 152 -156 152 -156 0 net=566
rlabel metal2 212 -156 212 -156 0 net=1084
rlabel metal2 296 -156 296 -156 0 net=1114
rlabel metal2 310 -156 310 -156 0 net=1296
rlabel metal2 345 -156 345 -156 0 net=1232
rlabel metal2 44 -158 44 -158 0 net=439
rlabel metal2 107 -158 107 -158 0 net=745
rlabel metal2 163 -158 163 -158 0 net=878
rlabel metal2 296 -158 296 -158 0 net=1163
rlabel metal2 51 -160 51 -160 0 net=335
rlabel metal2 79 -160 79 -160 0 net=770
rlabel metal2 128 -160 128 -160 0 net=555
rlabel metal2 163 -160 163 -160 0 net=471
rlabel metal2 201 -160 201 -160 0 net=790
rlabel metal2 303 -160 303 -160 0 net=1139
rlabel metal2 51 -162 51 -162 0 net=533
rlabel metal2 86 -162 86 -162 0 net=964
rlabel metal2 114 -162 114 -162 0 net=47
rlabel metal2 184 -162 184 -162 0 net=494
rlabel metal2 219 -162 219 -162 0 net=631
rlabel metal2 303 -162 303 -162 0 net=938
rlabel metal2 58 -164 58 -164 0 net=901
rlabel metal2 86 -164 86 -164 0 net=1071
rlabel metal2 93 -166 93 -166 0 net=583
rlabel metal2 149 -166 149 -166 0 net=595
rlabel metal2 198 -166 198 -166 0 net=973
rlabel metal2 135 -168 135 -168 0 net=453
rlabel metal2 180 -168 180 -168 0 net=1342
rlabel metal2 142 -170 142 -170 0 net=505
rlabel metal2 156 -170 156 -170 0 net=638
rlabel metal2 198 -170 198 -170 0 net=687
rlabel metal2 268 -170 268 -170 0 net=813
rlabel metal2 166 -172 166 -172 0 net=77
rlabel metal2 233 -172 233 -172 0 net=721
rlabel metal2 173 -174 173 -174 0 net=1106
rlabel metal2 121 -176 121 -176 0 net=702
rlabel metal2 205 -176 205 -176 0 net=1157
rlabel metal2 100 -178 100 -178 0 net=1237
rlabel metal2 254 -178 254 -178 0 net=1101
rlabel metal2 254 -180 254 -180 0 net=955
rlabel metal2 261 -182 261 -182 0 net=1261
rlabel metal2 212 -184 212 -184 0 net=1095
rlabel metal2 30 -195 30 -195 0 net=621
rlabel metal2 79 -195 79 -195 0 net=902
rlabel metal2 86 -195 86 -195 0 net=1072
rlabel metal2 159 -195 159 -195 0 net=632
rlabel metal2 226 -195 226 -195 0 net=913
rlabel metal2 226 -195 226 -195 0 net=913
rlabel metal2 229 -195 229 -195 0 net=1262
rlabel metal2 289 -195 289 -195 0 net=1103
rlabel metal2 289 -195 289 -195 0 net=1103
rlabel metal2 296 -195 296 -195 0 net=1140
rlabel metal2 331 -195 331 -195 0 net=1369
rlabel metal2 359 -195 359 -195 0 net=213
rlabel metal2 37 -197 37 -197 0 net=344
rlabel metal2 72 -197 72 -197 0 net=575
rlabel metal2 121 -197 121 -197 0 net=737
rlabel metal2 159 -197 159 -197 0 net=1096
rlabel metal2 296 -197 296 -197 0 net=1165
rlabel metal2 352 -197 352 -197 0 net=1025
rlabel metal2 373 -197 373 -197 0 net=1253
rlabel metal2 40 -199 40 -199 0 net=243
rlabel metal2 58 -199 58 -199 0 net=739
rlabel metal2 93 -199 93 -199 0 net=585
rlabel metal2 93 -199 93 -199 0 net=585
rlabel metal2 100 -199 100 -199 0 net=1239
rlabel metal2 212 -199 212 -199 0 net=956
rlabel metal2 303 -199 303 -199 0 net=1349
rlabel metal2 352 -199 352 -199 0 net=743
rlabel metal2 44 -201 44 -201 0 net=441
rlabel metal2 135 -201 135 -201 0 net=455
rlabel metal2 180 -201 180 -201 0 net=187
rlabel metal2 44 -203 44 -203 0 net=991
rlabel metal2 103 -203 103 -203 0 net=137
rlabel metal2 135 -203 135 -203 0 net=1303
rlabel metal2 303 -203 303 -203 0 net=1063
rlabel metal2 51 -205 51 -205 0 net=534
rlabel metal2 107 -205 107 -205 0 net=746
rlabel metal2 163 -205 163 -205 0 net=473
rlabel metal2 187 -205 187 -205 0 net=688
rlabel metal2 215 -205 215 -205 0 net=841
rlabel metal2 240 -205 240 -205 0 net=1158
rlabel metal2 65 -207 65 -207 0 net=655
rlabel metal2 128 -207 128 -207 0 net=557
rlabel metal2 149 -207 149 -207 0 net=507
rlabel metal2 184 -207 184 -207 0 net=771
rlabel metal2 233 -207 233 -207 0 net=723
rlabel metal2 107 -209 107 -209 0 net=775
rlabel metal2 149 -209 149 -209 0 net=251
rlabel metal2 243 -209 243 -209 0 net=814
rlabel metal2 191 -211 191 -211 0 net=597
rlabel metal2 191 -211 191 -211 0 net=597
rlabel metal2 215 -211 215 -211 0 net=927
rlabel metal2 247 -213 247 -213 0 net=975
rlabel metal2 240 -215 240 -215 0 net=805
rlabel metal2 254 -215 254 -215 0 net=779
rlabel metal2 9 -226 9 -226 0 net=1211
rlabel metal2 54 -226 54 -226 0 net=459
rlabel metal2 107 -226 107 -226 0 net=738
rlabel metal2 128 -226 128 -226 0 net=776
rlabel metal2 177 -226 177 -226 0 net=474
rlabel metal2 222 -226 222 -226 0 net=1104
rlabel metal2 296 -226 296 -226 0 net=1167
rlabel metal2 296 -226 296 -226 0 net=1167
rlabel metal2 310 -226 310 -226 0 net=1351
rlabel metal2 334 -226 334 -226 0 net=132
rlabel metal2 380 -226 380 -226 0 net=1254
rlabel metal2 380 -226 380 -226 0 net=1254
rlabel metal2 387 -226 387 -226 0 net=1145
rlabel metal2 16 -228 16 -228 0 net=993
rlabel metal2 65 -228 65 -228 0 net=657
rlabel metal2 65 -228 65 -228 0 net=657
rlabel metal2 79 -228 79 -228 0 net=467
rlabel metal2 159 -228 159 -228 0 net=921
rlabel metal2 212 -228 212 -228 0 net=57
rlabel metal2 345 -228 345 -228 0 net=1371
rlabel metal2 355 -228 355 -228 0 net=1026
rlabel metal2 23 -230 23 -230 0 net=741
rlabel metal2 93 -230 93 -230 0 net=587
rlabel metal2 233 -230 233 -230 0 net=724
rlabel metal2 282 -230 282 -230 0 net=1305
rlabel metal2 327 -230 327 -230 0 net=744
rlabel metal2 30 -232 30 -232 0 net=622
rlabel metal2 93 -232 93 -232 0 net=537
rlabel metal2 226 -232 226 -232 0 net=915
rlabel metal2 289 -232 289 -232 0 net=1035
rlabel metal2 33 -234 33 -234 0 net=1079
rlabel metal2 37 -236 37 -236 0 net=26
rlabel metal2 114 -236 114 -236 0 net=442
rlabel metal2 149 -236 149 -236 0 net=73
rlabel metal2 198 -236 198 -236 0 net=773
rlabel metal2 233 -236 233 -236 0 net=781
rlabel metal2 268 -236 268 -236 0 net=929
rlabel metal2 303 -236 303 -236 0 net=1064
rlabel metal2 51 -238 51 -238 0 net=342
rlabel metal2 114 -238 114 -238 0 net=409
rlabel metal2 135 -238 135 -238 0 net=559
rlabel metal2 149 -238 149 -238 0 net=508
rlabel metal2 191 -238 191 -238 0 net=599
rlabel metal2 205 -238 205 -238 0 net=1241
rlabel metal2 58 -240 58 -240 0 net=577
rlabel metal2 152 -240 152 -240 0 net=1133
rlabel metal2 170 -240 170 -240 0 net=457
rlabel metal2 208 -240 208 -240 0 net=1059
rlabel metal2 44 -242 44 -242 0 net=751
rlabel metal2 170 -242 170 -242 0 net=1007
rlabel metal2 240 -242 240 -242 0 net=807
rlabel metal2 250 -242 250 -242 0 net=976
rlabel metal2 72 -244 72 -244 0 net=491
rlabel metal2 219 -244 219 -244 0 net=843
rlabel metal2 261 -244 261 -244 0 net=1171
rlabel metal2 9 -255 9 -255 0 net=1212
rlabel metal2 37 -255 37 -255 0 net=601
rlabel metal2 205 -255 205 -255 0 net=782
rlabel metal2 268 -255 268 -255 0 net=1168
rlabel metal2 345 -255 345 -255 0 net=1372
rlabel metal2 387 -255 387 -255 0 net=1146
rlabel metal2 9 -257 9 -257 0 net=302
rlabel metal2 72 -257 72 -257 0 net=492
rlabel metal2 89 -257 89 -257 0 net=89
rlabel metal2 128 -257 128 -257 0 net=774
rlabel metal2 282 -257 282 -257 0 net=931
rlabel metal2 282 -257 282 -257 0 net=931
rlabel metal2 16 -259 16 -259 0 net=994
rlabel metal2 145 -259 145 -259 0 net=1321
rlabel metal2 16 -261 16 -261 0 net=447
rlabel metal2 135 -261 135 -261 0 net=561
rlabel metal2 149 -261 149 -261 0 net=1317
rlabel metal2 23 -263 23 -263 0 net=742
rlabel metal2 79 -263 79 -263 0 net=458
rlabel metal2 208 -263 208 -263 0 net=808
rlabel metal2 23 -265 23 -265 0 net=897
rlabel metal2 93 -265 93 -265 0 net=538
rlabel metal2 149 -265 149 -265 0 net=1242
rlabel metal2 51 -267 51 -267 0 net=1134
rlabel metal2 173 -267 173 -267 0 net=588
rlabel metal2 215 -267 215 -267 0 net=1306
rlabel metal2 54 -269 54 -269 0 net=158
rlabel metal2 289 -269 289 -269 0 net=1037
rlabel metal2 310 -269 310 -269 0 net=1081
rlabel metal2 58 -271 58 -271 0 net=578
rlabel metal2 100 -271 100 -271 0 net=461
rlabel metal2 156 -271 156 -271 0 net=468
rlabel metal2 226 -271 226 -271 0 net=845
rlabel metal2 254 -271 254 -271 0 net=1061
rlabel metal2 58 -273 58 -273 0 net=659
rlabel metal2 72 -273 72 -273 0 net=387
rlabel metal2 100 -273 100 -273 0 net=433
rlabel metal2 159 -273 159 -273 0 net=871
rlabel metal2 254 -273 254 -273 0 net=917
rlabel metal2 2 -275 2 -275 0 net=989
rlabel metal2 107 -275 107 -275 0 net=717
rlabel metal2 170 -275 170 -275 0 net=939
rlabel metal2 233 -275 233 -275 0 net=903
rlabel metal2 107 -277 107 -277 0 net=411
rlabel metal2 170 -277 170 -277 0 net=835
rlabel metal2 212 -277 212 -277 0 net=1205
rlabel metal2 121 -279 121 -279 0 net=639
rlabel metal2 191 -279 191 -279 0 net=1352
rlabel metal2 156 -281 156 -281 0 net=1223
rlabel metal2 177 -283 177 -283 0 net=923
rlabel metal2 44 -285 44 -285 0 net=752
rlabel metal2 180 -285 180 -285 0 net=1172
rlabel metal2 44 -287 44 -287 0 net=643
rlabel metal2 184 -287 184 -287 0 net=1009
rlabel metal2 194 -289 194 -289 0 net=957
rlabel metal2 222 -291 222 -291 0 net=1199
rlabel metal2 2 -302 2 -302 0 net=990
rlabel metal2 44 -302 44 -302 0 net=644
rlabel metal2 205 -302 205 -302 0 net=904
rlabel metal2 16 -304 16 -304 0 net=448
rlabel metal2 79 -304 79 -304 0 net=83
rlabel metal2 156 -304 156 -304 0 net=150
rlabel metal2 156 -304 156 -304 0 net=150
rlabel metal2 170 -304 170 -304 0 net=924
rlabel metal2 23 -306 23 -306 0 net=898
rlabel metal2 65 -306 65 -306 0 net=718
rlabel metal2 187 -306 187 -306 0 net=918
rlabel metal2 261 -306 261 -306 0 net=1201
rlabel metal2 30 -308 30 -308 0 net=661
rlabel metal2 65 -308 65 -308 0 net=697
rlabel metal2 135 -308 135 -308 0 net=462
rlabel metal2 212 -308 212 -308 0 net=1038
rlabel metal2 37 -310 37 -310 0 net=602
rlabel metal2 212 -310 212 -310 0 net=1153
rlabel metal2 282 -310 282 -310 0 net=933
rlabel metal2 37 -312 37 -312 0 net=1265
rlabel metal2 215 -312 215 -312 0 net=979
rlabel metal2 240 -312 240 -312 0 net=1247
rlabel metal2 44 -314 44 -314 0 net=863
rlabel metal2 107 -314 107 -314 0 net=412
rlabel metal2 163 -314 163 -314 0 net=691
rlabel metal2 208 -314 208 -314 0 net=1183
rlabel metal2 51 -316 51 -316 0 net=167
rlabel metal2 142 -316 142 -316 0 net=562
rlabel metal2 184 -316 184 -316 0 net=1085
rlabel metal2 58 -318 58 -318 0 net=369
rlabel metal2 117 -318 117 -318 0 net=1206
rlabel metal2 79 -320 79 -320 0 net=681
rlabel metal2 215 -320 215 -320 0 net=1224
rlabel metal2 86 -322 86 -322 0 net=389
rlabel metal2 96 -322 96 -322 0 net=1010
rlabel metal2 324 -322 324 -322 0 net=1323
rlabel metal2 86 -324 86 -324 0 net=641
rlabel metal2 128 -324 128 -324 0 net=1067
rlabel metal2 229 -324 229 -324 0 net=1082
rlabel metal2 100 -326 100 -326 0 net=435
rlabel metal2 226 -326 226 -326 0 net=847
rlabel metal2 110 -328 110 -328 0 net=1318
rlabel metal2 135 -330 135 -330 0 net=872
rlabel metal2 142 -332 142 -332 0 net=358
rlabel metal2 219 -332 219 -332 0 net=941
rlabel metal2 121 -334 121 -334 0 net=535
rlabel metal2 198 -334 198 -334 0 net=837
rlabel metal2 243 -334 243 -334 0 net=1062
rlabel metal2 198 -336 198 -336 0 net=958
rlabel metal2 296 -336 296 -336 0 net=1123
rlabel metal2 201 -338 201 -338 0 net=1193
rlabel metal2 2 -349 2 -349 0 net=1195
rlabel metal2 121 -349 121 -349 0 net=401
rlabel metal2 145 -349 145 -349 0 net=569
rlabel metal2 205 -349 205 -349 0 net=848
rlabel metal2 16 -351 16 -351 0 net=699
rlabel metal2 79 -351 79 -351 0 net=682
rlabel metal2 93 -351 93 -351 0 net=391
rlabel metal2 103 -351 103 -351 0 net=692
rlabel metal2 170 -351 170 -351 0 net=436
rlabel metal2 170 -351 170 -351 0 net=436
rlabel metal2 173 -351 173 -351 0 net=1291
rlabel metal2 23 -353 23 -353 0 net=589
rlabel metal2 145 -353 145 -353 0 net=43
rlabel metal2 215 -353 215 -353 0 net=1177
rlabel metal2 243 -353 243 -353 0 net=1194
rlabel metal2 289 -353 289 -353 0 net=1203
rlabel metal2 30 -355 30 -355 0 net=662
rlabel metal2 75 -355 75 -355 0 net=607
rlabel metal2 86 -355 86 -355 0 net=642
rlabel metal2 149 -355 149 -355 0 net=417
rlabel metal2 177 -355 177 -355 0 net=536
rlabel metal2 219 -355 219 -355 0 net=839
rlabel metal2 9 -357 9 -357 0 net=1343
rlabel metal2 93 -357 93 -357 0 net=172
rlabel metal2 226 -357 226 -357 0 net=981
rlabel metal2 268 -357 268 -357 0 net=1185
rlabel metal2 299 -357 299 -357 0 net=1324
rlabel metal2 37 -359 37 -359 0 net=1266
rlabel metal2 152 -359 152 -359 0 net=959
rlabel metal2 303 -359 303 -359 0 net=935
rlabel metal2 37 -361 37 -361 0 net=407
rlabel metal2 117 -361 117 -361 0 net=1248
rlabel metal2 310 -361 310 -361 0 net=1125
rlabel metal2 310 -361 310 -361 0 net=1125
rlabel metal2 44 -363 44 -363 0 net=864
rlabel metal2 163 -363 163 -363 0 net=1021
rlabel metal2 44 -365 44 -365 0 net=709
rlabel metal2 184 -365 184 -365 0 net=1257
rlabel metal2 51 -367 51 -367 0 net=487
rlabel metal2 128 -367 128 -367 0 net=1069
rlabel metal2 233 -367 233 -367 0 net=943
rlabel metal2 254 -367 254 -367 0 net=1087
rlabel metal2 58 -369 58 -369 0 net=371
rlabel metal2 128 -369 128 -369 0 net=707
rlabel metal2 247 -369 247 -369 0 net=849
rlabel metal2 194 -371 194 -371 0 net=1129
rlabel metal2 261 -371 261 -371 0 net=1155
rlabel metal2 205 -373 205 -373 0 net=895
rlabel metal2 9 -384 9 -384 0 net=1344
rlabel metal2 68 -384 68 -384 0 net=1186
rlabel metal2 306 -384 306 -384 0 net=1126
rlabel metal2 16 -386 16 -386 0 net=700
rlabel metal2 75 -386 75 -386 0 net=102
rlabel metal2 107 -386 107 -386 0 net=372
rlabel metal2 128 -386 128 -386 0 net=708
rlabel metal2 215 -386 215 -386 0 net=840
rlabel metal2 23 -388 23 -388 0 net=590
rlabel metal2 86 -388 86 -388 0 net=747
rlabel metal2 128 -388 128 -388 0 net=419
rlabel metal2 152 -388 152 -388 0 net=570
rlabel metal2 205 -388 205 -388 0 net=896
rlabel metal2 233 -388 233 -388 0 net=945
rlabel metal2 233 -388 233 -388 0 net=945
rlabel metal2 261 -388 261 -388 0 net=1204
rlabel metal2 2 -390 2 -390 0 net=1197
rlabel metal2 30 -390 30 -390 0 net=571
rlabel metal2 30 -390 30 -390 0 net=571
rlabel metal2 37 -390 37 -390 0 net=408
rlabel metal2 93 -390 93 -390 0 net=392
rlabel metal2 135 -390 135 -390 0 net=825
rlabel metal2 156 -390 156 -390 0 net=254
rlabel metal2 194 -390 194 -390 0 net=1156
rlabel metal2 285 -390 285 -390 0 net=865
rlabel metal2 44 -392 44 -392 0 net=710
rlabel metal2 96 -392 96 -392 0 net=402
rlabel metal2 138 -392 138 -392 0 net=1233
rlabel metal2 201 -392 201 -392 0 net=1243
rlabel metal2 271 -392 271 -392 0 net=1293
rlabel metal2 44 -394 44 -394 0 net=711
rlabel metal2 142 -394 142 -394 0 net=757
rlabel metal2 163 -394 163 -394 0 net=703
rlabel metal2 205 -394 205 -394 0 net=995
rlabel metal2 282 -394 282 -394 0 net=936
rlabel metal2 51 -396 51 -396 0 net=489
rlabel metal2 166 -396 166 -396 0 net=1070
rlabel metal2 289 -396 289 -396 0 net=1023
rlabel metal2 40 -398 40 -398 0 net=79
rlabel metal2 58 -398 58 -398 0 net=609
rlabel metal2 170 -398 170 -398 0 net=1130
rlabel metal2 292 -398 292 -398 0 net=1285
rlabel metal2 79 -400 79 -400 0 net=128
rlabel metal2 177 -400 177 -400 0 net=1258
rlabel metal2 177 -402 177 -402 0 net=861
rlabel metal2 219 -402 219 -402 0 net=982
rlabel metal2 240 -402 240 -402 0 net=1179
rlabel metal2 156 -404 156 -404 0 net=361
rlabel metal2 180 -406 180 -406 0 net=195
rlabel metal2 184 -408 184 -408 0 net=851
rlabel metal2 247 -410 247 -410 0 net=961
rlabel metal2 268 -412 268 -412 0 net=1089
rlabel metal2 268 -414 268 -414 0 net=1292
rlabel metal2 2 -425 2 -425 0 net=1263
rlabel metal2 135 -425 135 -425 0 net=826
rlabel metal2 229 -425 229 -425 0 net=1039
rlabel metal2 254 -425 254 -425 0 net=1181
rlabel metal2 310 -425 310 -425 0 net=1287
rlabel metal2 310 -425 310 -425 0 net=1287
rlabel metal2 317 -425 317 -425 0 net=1294
rlabel metal2 9 -427 9 -427 0 net=713
rlabel metal2 47 -427 47 -427 0 net=763
rlabel metal2 54 -427 54 -427 0 net=490
rlabel metal2 72 -427 72 -427 0 net=221
rlabel metal2 114 -427 114 -427 0 net=759
rlabel metal2 149 -427 149 -427 0 net=705
rlabel metal2 170 -427 170 -427 0 net=862
rlabel metal2 201 -427 201 -427 0 net=946
rlabel metal2 268 -427 268 -427 0 net=1024
rlabel metal2 324 -427 324 -427 0 net=883
rlabel metal2 16 -429 16 -429 0 net=611
rlabel metal2 65 -429 65 -429 0 net=427
rlabel metal2 107 -429 107 -429 0 net=799
rlabel metal2 170 -429 170 -429 0 net=852
rlabel metal2 205 -429 205 -429 0 net=996
rlabel metal2 222 -429 222 -429 0 net=1345
rlabel metal2 23 -431 23 -431 0 net=1198
rlabel metal2 79 -431 79 -431 0 net=1075
rlabel metal2 107 -431 107 -431 0 net=677
rlabel metal2 128 -431 128 -431 0 net=420
rlabel metal2 128 -431 128 -431 0 net=420
rlabel metal2 142 -431 142 -431 0 net=363
rlabel metal2 184 -431 184 -431 0 net=801
rlabel metal2 201 -431 201 -431 0 net=977
rlabel metal2 226 -431 226 -431 0 net=815
rlabel metal2 23 -433 23 -433 0 net=653
rlabel metal2 233 -433 233 -433 0 net=1361
rlabel metal2 261 -433 261 -433 0 net=1245
rlabel metal2 30 -435 30 -435 0 net=572
rlabel metal2 72 -435 72 -435 0 net=1003
rlabel metal2 30 -437 30 -437 0 net=749
rlabel metal2 110 -437 110 -437 0 net=1147
rlabel metal2 219 -437 219 -437 0 net=879
rlabel metal2 268 -437 268 -437 0 net=867
rlabel metal2 37 -439 37 -439 0 net=385
rlabel metal2 173 -439 173 -439 0 net=63
rlabel metal2 275 -439 275 -439 0 net=1091
rlabel metal2 275 -439 275 -439 0 net=1091
rlabel metal2 82 -441 82 -441 0 net=42
rlabel metal2 191 -441 191 -441 0 net=1235
rlabel metal2 191 -443 191 -443 0 net=962
rlabel metal2 156 -445 156 -445 0 net=1267
rlabel metal2 2 -456 2 -456 0 net=1264
rlabel metal2 107 -456 107 -456 0 net=591
rlabel metal2 170 -456 170 -456 0 net=919
rlabel metal2 177 -456 177 -456 0 net=1149
rlabel metal2 198 -456 198 -456 0 net=1346
rlabel metal2 320 -456 320 -456 0 net=1335
rlabel metal2 359 -456 359 -456 0 net=1297
rlabel metal2 9 -458 9 -458 0 net=714
rlabel metal2 75 -458 75 -458 0 net=800
rlabel metal2 194 -458 194 -458 0 net=294
rlabel metal2 331 -458 331 -458 0 net=885
rlabel metal2 16 -460 16 -460 0 net=612
rlabel metal2 93 -460 93 -460 0 net=1077
rlabel metal2 205 -460 205 -460 0 net=978
rlabel metal2 215 -460 215 -460 0 net=1004
rlabel metal2 310 -460 310 -460 0 net=1288
rlabel metal2 23 -462 23 -462 0 net=654
rlabel metal2 44 -462 44 -462 0 net=719
rlabel metal2 135 -462 135 -462 0 net=1246
rlabel metal2 327 -462 327 -462 0 net=1109
rlabel metal2 30 -464 30 -464 0 net=750
rlabel metal2 110 -464 110 -464 0 net=1236
rlabel metal2 37 -466 37 -466 0 net=386
rlabel metal2 93 -466 93 -466 0 net=365
rlabel metal2 184 -466 184 -466 0 net=803
rlabel metal2 219 -466 219 -466 0 net=1359
rlabel metal2 51 -468 51 -468 0 net=765
rlabel metal2 100 -468 100 -468 0 net=169
rlabel metal2 180 -468 180 -468 0 net=1311
rlabel metal2 219 -468 219 -468 0 net=1225
rlabel metal2 51 -470 51 -470 0 net=909
rlabel metal2 100 -470 100 -470 0 net=647
rlabel metal2 226 -470 226 -470 0 net=817
rlabel metal2 226 -470 226 -470 0 net=817
rlabel metal2 233 -470 233 -470 0 net=1182
rlabel metal2 114 -472 114 -472 0 net=760
rlabel metal2 233 -472 233 -472 0 net=869
rlabel metal2 275 -472 275 -472 0 net=1093
rlabel metal2 114 -474 114 -474 0 net=679
rlabel metal2 128 -474 128 -474 0 net=269
rlabel metal2 247 -474 247 -474 0 net=1269
rlabel metal2 121 -476 121 -476 0 net=706
rlabel metal2 215 -476 215 -476 0 net=1159
rlabel metal2 254 -476 254 -476 0 net=1363
rlabel metal2 86 -478 86 -478 0 net=521
rlabel metal2 65 -480 65 -480 0 net=429
rlabel metal2 128 -480 128 -480 0 net=880
rlabel metal2 61 -482 61 -482 0 net=1001
rlabel metal2 138 -482 138 -482 0 net=1055
rlabel metal2 240 -482 240 -482 0 net=1041
rlabel metal2 142 -484 142 -484 0 net=1005
rlabel metal2 236 -486 236 -486 0 net=831
rlabel metal2 16 -497 16 -497 0 net=911
rlabel metal2 65 -497 65 -497 0 net=1002
rlabel metal2 103 -497 103 -497 0 net=290
rlabel metal2 184 -497 184 -497 0 net=1312
rlabel metal2 282 -497 282 -497 0 net=1360
rlabel metal2 310 -497 310 -497 0 net=1365
rlabel metal2 331 -497 331 -497 0 net=886
rlabel metal2 352 -497 352 -497 0 net=1337
rlabel metal2 352 -497 352 -497 0 net=1337
rlabel metal2 23 -499 23 -499 0 net=1315
rlabel metal2 114 -499 114 -499 0 net=680
rlabel metal2 149 -499 149 -499 0 net=523
rlabel metal2 198 -499 198 -499 0 net=161
rlabel metal2 275 -499 275 -499 0 net=1271
rlabel metal2 320 -499 320 -499 0 net=1110
rlabel metal2 345 -499 345 -499 0 net=1299
rlabel metal2 30 -501 30 -501 0 net=1169
rlabel metal2 72 -501 72 -501 0 net=430
rlabel metal2 93 -501 93 -501 0 net=367
rlabel metal2 121 -501 121 -501 0 net=475
rlabel metal2 177 -501 177 -501 0 net=1307
rlabel metal2 58 -503 58 -503 0 net=767
rlabel metal2 72 -503 72 -503 0 net=649
rlabel metal2 135 -503 135 -503 0 net=348
rlabel metal2 201 -503 201 -503 0 net=1006
rlabel metal2 296 -503 296 -503 0 net=1226
rlabel metal2 44 -505 44 -505 0 net=720
rlabel metal2 138 -505 138 -505 0 net=1078
rlabel metal2 180 -505 180 -505 0 net=967
rlabel metal2 222 -505 222 -505 0 net=1273
rlabel metal2 44 -507 44 -507 0 net=539
rlabel metal2 86 -507 86 -507 0 net=1057
rlabel metal2 163 -507 163 -507 0 net=920
rlabel metal2 201 -507 201 -507 0 net=818
rlabel metal2 229 -507 229 -507 0 net=1011
rlabel metal2 93 -509 93 -509 0 net=567
rlabel metal2 142 -509 142 -509 0 net=515
rlabel metal2 226 -509 226 -509 0 net=615
rlabel metal2 82 -511 82 -511 0 net=397
rlabel metal2 156 -511 156 -511 0 net=804
rlabel metal2 233 -511 233 -511 0 net=870
rlabel metal2 107 -513 107 -513 0 net=593
rlabel metal2 240 -513 240 -513 0 net=833
rlabel metal2 240 -513 240 -513 0 net=833
rlabel metal2 247 -513 247 -513 0 net=1161
rlabel metal2 107 -515 107 -515 0 net=375
rlabel metal2 191 -515 191 -515 0 net=1151
rlabel metal2 254 -515 254 -515 0 net=1094
rlabel metal2 124 -517 124 -517 0 net=1027
rlabel metal2 159 -519 159 -519 0 net=855
rlabel metal2 261 -519 261 -519 0 net=1043
rlabel metal2 205 -521 205 -521 0 net=887
rlabel metal2 212 -523 212 -523 0 net=665
rlabel metal2 9 -534 9 -534 0 net=1229
rlabel metal2 37 -534 37 -534 0 net=108
rlabel metal2 51 -534 51 -534 0 net=541
rlabel metal2 51 -534 51 -534 0 net=541
rlabel metal2 61 -534 61 -534 0 net=568
rlabel metal2 100 -534 100 -534 0 net=393
rlabel metal2 201 -534 201 -534 0 net=667
rlabel metal2 208 -534 208 -534 0 net=1274
rlabel metal2 331 -534 331 -534 0 net=1300
rlabel metal2 352 -534 352 -534 0 net=1338
rlabel metal2 16 -536 16 -536 0 net=912
rlabel metal2 86 -536 86 -536 0 net=1058
rlabel metal2 212 -536 212 -536 0 net=1272
rlabel metal2 331 -536 331 -536 0 net=549
rlabel metal2 16 -538 16 -538 0 net=925
rlabel metal2 93 -538 93 -538 0 net=663
rlabel metal2 222 -538 222 -538 0 net=1162
rlabel metal2 23 -540 23 -540 0 net=1316
rlabel metal2 121 -540 121 -540 0 net=1115
rlabel metal2 138 -540 138 -540 0 net=834
rlabel metal2 250 -540 250 -540 0 net=1173
rlabel metal2 23 -542 23 -542 0 net=899
rlabel metal2 65 -542 65 -542 0 net=768
rlabel metal2 65 -542 65 -542 0 net=768
rlabel metal2 68 -542 68 -542 0 net=551
rlabel metal2 114 -542 114 -542 0 net=368
rlabel metal2 191 -542 191 -542 0 net=633
rlabel metal2 30 -544 30 -544 0 net=1170
rlabel metal2 58 -544 58 -544 0 net=259
rlabel metal2 124 -544 124 -544 0 net=1152
rlabel metal2 268 -544 268 -544 0 net=1255
rlabel metal2 128 -546 128 -546 0 net=399
rlabel metal2 128 -546 128 -546 0 net=399
rlabel metal2 135 -546 135 -546 0 net=405
rlabel metal2 226 -546 226 -546 0 net=1119
rlabel metal2 247 -546 247 -546 0 net=827
rlabel metal2 142 -548 142 -548 0 net=517
rlabel metal2 142 -548 142 -548 0 net=517
rlabel metal2 156 -548 156 -548 0 net=666
rlabel metal2 261 -548 261 -548 0 net=889
rlabel metal2 271 -548 271 -548 0 net=1366
rlabel metal2 107 -550 107 -550 0 net=377
rlabel metal2 159 -550 159 -550 0 net=594
rlabel metal2 177 -550 177 -550 0 net=445
rlabel metal2 233 -550 233 -550 0 net=857
rlabel metal2 324 -550 324 -550 0 net=1309
rlabel metal2 72 -552 72 -552 0 net=650
rlabel metal2 163 -552 163 -552 0 net=616
rlabel metal2 61 -554 61 -554 0 net=1015
rlabel metal2 163 -554 163 -554 0 net=905
rlabel metal2 166 -556 166 -556 0 net=421
rlabel metal2 233 -556 233 -556 0 net=1333
rlabel metal2 170 -558 170 -558 0 net=525
rlabel metal2 254 -558 254 -558 0 net=1045
rlabel metal2 149 -560 149 -560 0 net=477
rlabel metal2 289 -560 289 -560 0 net=1029
rlabel metal2 282 -562 282 -562 0 net=1013
rlabel metal2 219 -564 219 -564 0 net=969
rlabel metal2 219 -566 219 -566 0 net=1187
rlabel metal2 9 -577 9 -577 0 net=1230
rlabel metal2 68 -577 68 -577 0 net=31
rlabel metal2 86 -577 86 -577 0 net=553
rlabel metal2 86 -577 86 -577 0 net=553
rlabel metal2 93 -577 93 -577 0 net=664
rlabel metal2 114 -577 114 -577 0 net=406
rlabel metal2 219 -577 219 -577 0 net=1310
rlabel metal2 345 -577 345 -577 0 net=828
rlabel metal2 23 -579 23 -579 0 net=900
rlabel metal2 72 -579 72 -579 0 net=1017
rlabel metal2 72 -579 72 -579 0 net=1017
rlabel metal2 79 -579 79 -579 0 net=182
rlabel metal2 114 -579 114 -579 0 net=1367
rlabel metal2 149 -579 149 -579 0 net=478
rlabel metal2 205 -579 205 -579 0 net=669
rlabel metal2 205 -579 205 -579 0 net=669
rlabel metal2 212 -579 212 -579 0 net=906
rlabel metal2 289 -579 289 -579 0 net=1014
rlabel metal2 44 -581 44 -581 0 net=542
rlabel metal2 93 -581 93 -581 0 net=1117
rlabel metal2 128 -581 128 -581 0 net=400
rlabel metal2 177 -581 177 -581 0 net=550
rlabel metal2 44 -583 44 -583 0 net=413
rlabel metal2 100 -583 100 -583 0 net=395
rlabel metal2 135 -583 135 -583 0 net=527
rlabel metal2 180 -583 180 -583 0 net=970
rlabel metal2 16 -585 16 -585 0 net=926
rlabel metal2 121 -585 121 -585 0 net=139
rlabel metal2 149 -585 149 -585 0 net=1065
rlabel metal2 219 -585 219 -585 0 net=1121
rlabel metal2 229 -585 229 -585 0 net=181
rlabel metal2 261 -585 261 -585 0 net=858
rlabel metal2 152 -587 152 -587 0 net=446
rlabel metal2 233 -587 233 -587 0 net=1256
rlabel metal2 156 -589 156 -589 0 net=378
rlabel metal2 233 -589 233 -589 0 net=1281
rlabel metal2 264 -589 264 -589 0 net=1334
rlabel metal2 142 -591 142 -591 0 net=519
rlabel metal2 163 -591 163 -591 0 net=809
rlabel metal2 191 -591 191 -591 0 net=422
rlabel metal2 236 -591 236 -591 0 net=270
rlabel metal2 243 -591 243 -591 0 net=1174
rlabel metal2 310 -591 310 -591 0 net=1189
rlabel metal2 187 -593 187 -593 0 net=1353
rlabel metal2 240 -593 240 -593 0 net=403
rlabel metal2 247 -595 247 -595 0 net=1030
rlabel metal2 250 -597 250 -597 0 net=634
rlabel metal2 254 -599 254 -599 0 net=1047
rlabel metal2 254 -601 254 -601 0 net=890
rlabel metal2 250 -603 250 -603 0 net=1329
rlabel metal2 51 -614 51 -614 0 net=415
rlabel metal2 51 -614 51 -614 0 net=415
rlabel metal2 65 -614 65 -614 0 net=11
rlabel metal2 72 -614 72 -614 0 net=1019
rlabel metal2 72 -614 72 -614 0 net=1019
rlabel metal2 79 -614 79 -614 0 net=1275
rlabel metal2 110 -614 110 -614 0 net=1368
rlabel metal2 128 -614 128 -614 0 net=396
rlabel metal2 187 -614 187 -614 0 net=404
rlabel metal2 261 -614 261 -614 0 net=1331
rlabel metal2 289 -614 289 -614 0 net=239
rlabel metal2 58 -616 58 -616 0 net=545
rlabel metal2 86 -616 86 -616 0 net=554
rlabel metal2 100 -616 100 -616 0 net=309
rlabel metal2 128 -616 128 -616 0 net=783
rlabel metal2 142 -616 142 -616 0 net=1066
rlabel metal2 194 -616 194 -616 0 net=1122
rlabel metal2 226 -616 226 -616 0 net=1227
rlabel metal2 268 -616 268 -616 0 net=1347
rlabel metal2 303 -616 303 -616 0 net=1191
rlabel metal2 86 -618 86 -618 0 net=463
rlabel metal2 114 -618 114 -618 0 net=529
rlabel metal2 142 -618 142 -618 0 net=354
rlabel metal2 198 -618 198 -618 0 net=1355
rlabel metal2 275 -618 275 -618 0 net=287
rlabel metal2 93 -620 93 -620 0 net=1118
rlabel metal2 156 -620 156 -620 0 net=520
rlabel metal2 233 -620 233 -620 0 net=1283
rlabel metal2 257 -620 257 -620 0 net=1357
rlabel metal2 156 -622 156 -622 0 net=381
rlabel metal2 233 -622 233 -622 0 net=1049
rlabel metal2 163 -624 163 -624 0 net=761
rlabel metal2 282 -624 282 -624 0 net=1373
rlabel metal2 166 -626 166 -626 0 net=971
rlabel metal2 170 -628 170 -628 0 net=715
rlabel metal2 177 -630 177 -630 0 net=811
rlabel metal2 177 -632 177 -632 0 net=1301
rlabel metal2 184 -634 184 -634 0 net=671
rlabel metal2 44 -645 44 -645 0 net=416
rlabel metal2 65 -645 65 -645 0 net=317
rlabel metal2 96 -645 96 -645 0 net=291
rlabel metal2 114 -645 114 -645 0 net=530
rlabel metal2 156 -645 156 -645 0 net=383
rlabel metal2 173 -645 173 -645 0 net=1284
rlabel metal2 243 -645 243 -645 0 net=1332
rlabel metal2 292 -645 292 -645 0 net=1192
rlabel metal2 44 -647 44 -647 0 net=997
rlabel metal2 58 -647 58 -647 0 net=547
rlabel metal2 72 -647 72 -647 0 net=1020
rlabel metal2 107 -647 107 -647 0 net=1277
rlabel metal2 121 -647 121 -647 0 net=22
rlabel metal2 149 -647 149 -647 0 net=972
rlabel metal2 233 -647 233 -647 0 net=1051
rlabel metal2 233 -647 233 -647 0 net=1051
rlabel metal2 247 -647 247 -647 0 net=1302
rlabel metal2 72 -649 72 -649 0 net=465
rlabel metal2 93 -649 93 -649 0 net=645
rlabel metal2 124 -649 124 -649 0 net=762
rlabel metal2 180 -649 180 -649 0 net=812
rlabel metal2 261 -649 261 -649 0 net=1374
rlabel metal2 79 -651 79 -651 0 net=423
rlabel metal2 128 -651 128 -651 0 net=784
rlabel metal2 184 -651 184 -651 0 net=673
rlabel metal2 208 -651 208 -651 0 net=1358
rlabel metal2 142 -653 142 -653 0 net=543
rlabel metal2 184 -653 184 -653 0 net=859
rlabel metal2 268 -653 268 -653 0 net=1348
rlabel metal2 191 -655 191 -655 0 net=716
rlabel metal2 201 -655 201 -655 0 net=1356
rlabel metal2 268 -655 268 -655 0 net=1219
rlabel metal2 191 -657 191 -657 0 net=573
rlabel metal2 254 -657 254 -657 0 net=1031
rlabel metal2 194 -659 194 -659 0 net=1228
rlabel metal2 226 -661 226 -661 0 net=495
rlabel metal2 44 -672 44 -672 0 net=999
rlabel metal2 58 -672 58 -672 0 net=548
rlabel metal2 72 -672 72 -672 0 net=466
rlabel metal2 93 -672 93 -672 0 net=32
rlabel metal2 103 -672 103 -672 0 net=646
rlabel metal2 114 -672 114 -672 0 net=1279
rlabel metal2 135 -672 135 -672 0 net=449
rlabel metal2 145 -672 145 -672 0 net=544
rlabel metal2 170 -672 170 -672 0 net=384
rlabel metal2 184 -672 184 -672 0 net=860
rlabel metal2 205 -672 205 -672 0 net=675
rlabel metal2 205 -672 205 -672 0 net=675
rlabel metal2 212 -672 212 -672 0 net=497
rlabel metal2 240 -672 240 -672 0 net=853
rlabel metal2 254 -672 254 -672 0 net=1033
rlabel metal2 254 -672 254 -672 0 net=1033
rlabel metal2 268 -672 268 -672 0 net=1221
rlabel metal2 285 -672 285 -672 0 net=339
rlabel metal2 58 -674 58 -674 0 net=891
rlabel metal2 72 -674 72 -674 0 net=100
rlabel metal2 121 -674 121 -674 0 net=431
rlabel metal2 191 -674 191 -674 0 net=574
rlabel metal2 226 -674 226 -674 0 net=1053
rlabel metal2 240 -674 240 -674 0 net=55
rlabel metal2 79 -676 79 -676 0 net=425
rlabel metal2 79 -676 79 -676 0 net=425
rlabel metal2 191 -676 191 -676 0 net=260
rlabel metal2 44 -687 44 -687 0 net=1000
rlabel metal2 58 -687 58 -687 0 net=892
rlabel metal2 79 -687 79 -687 0 net=426
rlabel metal2 93 -687 93 -687 0 net=353
rlabel metal2 117 -687 117 -687 0 net=432
rlabel metal2 135 -687 135 -687 0 net=450
rlabel metal2 198 -687 198 -687 0 net=676
rlabel metal2 212 -687 212 -687 0 net=498
rlabel metal2 226 -687 226 -687 0 net=1054
rlabel metal2 254 -687 254 -687 0 net=1034
rlabel metal2 275 -687 275 -687 0 net=1222
rlabel metal2 107 -689 107 -689 0 net=1280
rlabel metal2 142 -689 142 -689 0 net=320
rlabel metal2 233 -689 233 -689 0 net=854
<< end >>
