magic
tech scmos
timestamp 1555016756 
<< pdiffusion >>
rect 1 -14 7 -8
rect 8 -14 14 -8
rect 15 -14 21 -8
rect 22 -14 28 -8
rect 29 -14 35 -8
rect 36 -14 42 -8
rect 43 -14 49 -8
rect 50 -14 56 -8
rect 57 -14 63 -8
rect 92 -14 95 -8
rect 113 -14 116 -8
rect 120 -14 126 -8
rect 127 -14 130 -8
rect 134 -14 140 -8
rect 141 -14 147 -8
rect 148 -14 154 -8
rect 155 -14 161 -8
rect 162 -14 165 -8
rect 169 -14 172 -8
rect 176 -14 182 -8
rect 183 -14 186 -8
rect 190 -14 196 -8
rect 197 -14 200 -8
rect 204 -14 207 -8
rect 211 -14 214 -8
rect 218 -14 224 -8
rect 225 -14 231 -8
rect 232 -14 238 -8
rect 239 -14 242 -8
rect 253 -14 259 -8
rect 260 -14 263 -8
rect 288 -14 294 -8
rect 337 -14 343 -8
rect 1 -41 7 -35
rect 8 -41 14 -35
rect 15 -41 21 -35
rect 29 -41 35 -35
rect 36 -41 42 -35
rect 43 -41 49 -35
rect 50 -41 56 -35
rect 64 -41 70 -35
rect 71 -41 74 -35
rect 78 -41 84 -35
rect 92 -41 95 -35
rect 99 -41 105 -35
rect 106 -41 112 -35
rect 113 -41 119 -35
rect 120 -41 126 -35
rect 127 -41 133 -35
rect 134 -41 137 -35
rect 141 -41 147 -35
rect 148 -41 154 -35
rect 155 -41 161 -35
rect 162 -41 168 -35
rect 169 -41 172 -35
rect 176 -41 179 -35
rect 183 -41 186 -35
rect 190 -41 193 -35
rect 197 -41 200 -35
rect 204 -41 210 -35
rect 211 -41 214 -35
rect 218 -41 221 -35
rect 225 -41 228 -35
rect 232 -41 235 -35
rect 239 -41 242 -35
rect 246 -41 249 -35
rect 253 -41 256 -35
rect 267 -41 273 -35
rect 274 -41 277 -35
rect 281 -41 287 -35
rect 288 -41 294 -35
rect 295 -41 298 -35
rect 309 -41 315 -35
rect 316 -41 319 -35
rect 323 -41 326 -35
rect 330 -41 336 -35
rect 337 -41 340 -35
rect 344 -41 347 -35
rect 351 -41 354 -35
rect 386 -41 389 -35
rect 400 -41 406 -35
rect 1 -76 7 -70
rect 15 -76 18 -70
rect 22 -76 25 -70
rect 29 -76 35 -70
rect 36 -76 42 -70
rect 43 -76 46 -70
rect 50 -76 56 -70
rect 57 -76 63 -70
rect 64 -76 67 -70
rect 71 -76 77 -70
rect 78 -76 84 -70
rect 85 -76 91 -70
rect 92 -76 95 -70
rect 99 -76 102 -70
rect 106 -76 112 -70
rect 113 -76 119 -70
rect 120 -76 123 -70
rect 127 -76 130 -70
rect 134 -76 137 -70
rect 141 -76 144 -70
rect 148 -76 154 -70
rect 155 -76 158 -70
rect 162 -76 165 -70
rect 169 -76 172 -70
rect 176 -76 182 -70
rect 183 -76 189 -70
rect 190 -76 196 -70
rect 197 -76 203 -70
rect 204 -76 210 -70
rect 211 -76 214 -70
rect 218 -76 224 -70
rect 225 -76 228 -70
rect 232 -76 235 -70
rect 239 -76 242 -70
rect 246 -76 252 -70
rect 253 -76 256 -70
rect 260 -76 266 -70
rect 267 -76 273 -70
rect 274 -76 277 -70
rect 281 -76 287 -70
rect 288 -76 291 -70
rect 295 -76 301 -70
rect 302 -76 308 -70
rect 309 -76 312 -70
rect 316 -76 319 -70
rect 323 -76 326 -70
rect 330 -76 333 -70
rect 337 -76 343 -70
rect 344 -76 347 -70
rect 351 -76 357 -70
rect 358 -76 361 -70
rect 365 -76 368 -70
rect 372 -76 375 -70
rect 379 -76 382 -70
rect 386 -76 389 -70
rect 393 -76 399 -70
rect 400 -76 403 -70
rect 407 -76 410 -70
rect 414 -76 417 -70
rect 421 -76 424 -70
rect 428 -76 434 -70
rect 435 -76 438 -70
rect 1 -129 7 -123
rect 8 -129 14 -123
rect 15 -129 21 -123
rect 22 -129 28 -123
rect 29 -129 35 -123
rect 36 -129 42 -123
rect 43 -129 49 -123
rect 50 -129 56 -123
rect 57 -129 60 -123
rect 64 -129 70 -123
rect 71 -129 77 -123
rect 78 -129 81 -123
rect 85 -129 88 -123
rect 92 -129 95 -123
rect 99 -129 105 -123
rect 106 -129 109 -123
rect 113 -129 119 -123
rect 120 -129 123 -123
rect 127 -129 130 -123
rect 134 -129 140 -123
rect 141 -129 144 -123
rect 148 -129 151 -123
rect 155 -129 161 -123
rect 162 -129 165 -123
rect 169 -129 175 -123
rect 176 -129 182 -123
rect 183 -129 189 -123
rect 190 -129 193 -123
rect 197 -129 200 -123
rect 204 -129 207 -123
rect 211 -129 214 -123
rect 218 -129 221 -123
rect 225 -129 228 -123
rect 232 -129 235 -123
rect 239 -129 245 -123
rect 246 -129 249 -123
rect 253 -129 259 -123
rect 260 -129 263 -123
rect 267 -129 270 -123
rect 274 -129 277 -123
rect 281 -129 287 -123
rect 288 -129 294 -123
rect 295 -129 298 -123
rect 302 -129 305 -123
rect 309 -129 312 -123
rect 316 -129 319 -123
rect 323 -129 329 -123
rect 330 -129 336 -123
rect 337 -129 343 -123
rect 344 -129 347 -123
rect 351 -129 357 -123
rect 358 -129 361 -123
rect 365 -129 368 -123
rect 372 -129 378 -123
rect 379 -129 385 -123
rect 386 -129 389 -123
rect 393 -129 396 -123
rect 400 -129 403 -123
rect 407 -129 410 -123
rect 414 -129 417 -123
rect 421 -129 424 -123
rect 428 -129 431 -123
rect 435 -129 438 -123
rect 442 -129 445 -123
rect 449 -129 452 -123
rect 456 -129 459 -123
rect 463 -129 466 -123
rect 470 -129 473 -123
rect 477 -129 480 -123
rect 484 -129 487 -123
rect 491 -129 494 -123
rect 498 -129 501 -123
rect 505 -129 508 -123
rect 512 -129 515 -123
rect 519 -129 522 -123
rect 1 -204 7 -198
rect 8 -204 14 -198
rect 15 -204 21 -198
rect 22 -204 28 -198
rect 29 -204 35 -198
rect 36 -204 42 -198
rect 43 -204 46 -198
rect 50 -204 56 -198
rect 57 -204 60 -198
rect 64 -204 67 -198
rect 71 -204 74 -198
rect 78 -204 81 -198
rect 85 -204 91 -198
rect 92 -204 95 -198
rect 99 -204 102 -198
rect 106 -204 109 -198
rect 113 -204 119 -198
rect 120 -204 123 -198
rect 127 -204 130 -198
rect 134 -204 140 -198
rect 141 -204 147 -198
rect 148 -204 154 -198
rect 155 -204 158 -198
rect 162 -204 165 -198
rect 169 -204 172 -198
rect 176 -204 182 -198
rect 183 -204 189 -198
rect 190 -204 193 -198
rect 197 -204 203 -198
rect 204 -204 210 -198
rect 211 -204 217 -198
rect 218 -204 221 -198
rect 225 -204 228 -198
rect 232 -204 235 -198
rect 239 -204 242 -198
rect 246 -204 252 -198
rect 253 -204 259 -198
rect 260 -204 263 -198
rect 267 -204 273 -198
rect 274 -204 277 -198
rect 281 -204 287 -198
rect 288 -204 294 -198
rect 295 -204 298 -198
rect 302 -204 305 -198
rect 309 -204 315 -198
rect 316 -204 319 -198
rect 323 -204 326 -198
rect 330 -204 333 -198
rect 337 -204 343 -198
rect 344 -204 347 -198
rect 351 -204 354 -198
rect 358 -204 361 -198
rect 365 -204 368 -198
rect 372 -204 375 -198
rect 379 -204 382 -198
rect 386 -204 392 -198
rect 393 -204 396 -198
rect 400 -204 403 -198
rect 407 -204 413 -198
rect 414 -204 417 -198
rect 421 -204 427 -198
rect 428 -204 431 -198
rect 435 -204 438 -198
rect 442 -204 445 -198
rect 449 -204 452 -198
rect 456 -204 459 -198
rect 463 -204 466 -198
rect 470 -204 473 -198
rect 477 -204 480 -198
rect 484 -204 487 -198
rect 491 -204 494 -198
rect 498 -204 501 -198
rect 505 -204 508 -198
rect 512 -204 515 -198
rect 519 -204 522 -198
rect 526 -204 529 -198
rect 533 -204 536 -198
rect 540 -204 543 -198
rect 547 -204 550 -198
rect 554 -204 557 -198
rect 561 -204 564 -198
rect 568 -204 571 -198
rect 575 -204 578 -198
rect 582 -204 585 -198
rect 589 -204 592 -198
rect 596 -204 599 -198
rect 603 -204 606 -198
rect 610 -204 613 -198
rect 617 -204 620 -198
rect 624 -204 627 -198
rect 631 -204 634 -198
rect 638 -204 641 -198
rect 645 -204 648 -198
rect 652 -204 655 -198
rect 659 -204 662 -198
rect 1 -277 7 -271
rect 8 -277 14 -271
rect 15 -277 21 -271
rect 22 -277 28 -271
rect 29 -277 32 -271
rect 36 -277 42 -271
rect 43 -277 49 -271
rect 50 -277 53 -271
rect 57 -277 63 -271
rect 64 -277 67 -271
rect 71 -277 74 -271
rect 78 -277 84 -271
rect 85 -277 91 -271
rect 92 -277 95 -271
rect 99 -277 105 -271
rect 106 -277 109 -271
rect 113 -277 116 -271
rect 120 -277 126 -271
rect 127 -277 130 -271
rect 134 -277 137 -271
rect 141 -277 144 -271
rect 148 -277 151 -271
rect 155 -277 161 -271
rect 162 -277 165 -271
rect 169 -277 172 -271
rect 176 -277 182 -271
rect 183 -277 186 -271
rect 190 -277 193 -271
rect 197 -277 200 -271
rect 204 -277 207 -271
rect 211 -277 214 -271
rect 218 -277 221 -271
rect 225 -277 228 -271
rect 232 -277 235 -271
rect 239 -277 245 -271
rect 246 -277 252 -271
rect 253 -277 259 -271
rect 260 -277 263 -271
rect 267 -277 273 -271
rect 274 -277 280 -271
rect 281 -277 287 -271
rect 288 -277 291 -271
rect 295 -277 301 -271
rect 302 -277 308 -271
rect 309 -277 312 -271
rect 316 -277 322 -271
rect 323 -277 326 -271
rect 330 -277 336 -271
rect 337 -277 340 -271
rect 344 -277 347 -271
rect 351 -277 357 -271
rect 358 -277 361 -271
rect 365 -277 371 -271
rect 372 -277 375 -271
rect 379 -277 382 -271
rect 386 -277 389 -271
rect 393 -277 396 -271
rect 400 -277 403 -271
rect 407 -277 410 -271
rect 414 -277 417 -271
rect 421 -277 424 -271
rect 428 -277 431 -271
rect 435 -277 438 -271
rect 442 -277 445 -271
rect 449 -277 452 -271
rect 456 -277 459 -271
rect 463 -277 466 -271
rect 470 -277 473 -271
rect 477 -277 480 -271
rect 484 -277 487 -271
rect 491 -277 494 -271
rect 498 -277 501 -271
rect 505 -277 508 -271
rect 512 -277 515 -271
rect 519 -277 522 -271
rect 526 -277 529 -271
rect 533 -277 536 -271
rect 540 -277 543 -271
rect 547 -277 550 -271
rect 561 -277 564 -271
rect 568 -277 571 -271
rect 575 -277 578 -271
rect 582 -277 585 -271
rect 589 -277 592 -271
rect 596 -277 599 -271
rect 603 -277 606 -271
rect 610 -277 613 -271
rect 617 -277 623 -271
rect 624 -277 627 -271
rect 631 -277 634 -271
rect 638 -277 644 -271
rect 666 -277 669 -271
rect 1 -342 7 -336
rect 8 -342 14 -336
rect 15 -342 21 -336
rect 22 -342 28 -336
rect 29 -342 35 -336
rect 36 -342 39 -336
rect 43 -342 49 -336
rect 50 -342 56 -336
rect 57 -342 60 -336
rect 64 -342 70 -336
rect 71 -342 77 -336
rect 78 -342 84 -336
rect 85 -342 91 -336
rect 92 -342 95 -336
rect 99 -342 105 -336
rect 106 -342 109 -336
rect 113 -342 116 -336
rect 120 -342 123 -336
rect 127 -342 130 -336
rect 134 -342 140 -336
rect 141 -342 147 -336
rect 148 -342 151 -336
rect 155 -342 161 -336
rect 162 -342 168 -336
rect 169 -342 172 -336
rect 176 -342 179 -336
rect 183 -342 189 -336
rect 190 -342 193 -336
rect 197 -342 203 -336
rect 204 -342 207 -336
rect 211 -342 214 -336
rect 218 -342 221 -336
rect 225 -342 228 -336
rect 232 -342 235 -336
rect 239 -342 245 -336
rect 246 -342 249 -336
rect 253 -342 256 -336
rect 260 -342 263 -336
rect 267 -342 270 -336
rect 274 -342 277 -336
rect 281 -342 284 -336
rect 288 -342 291 -336
rect 295 -342 298 -336
rect 302 -342 305 -336
rect 309 -342 315 -336
rect 316 -342 322 -336
rect 323 -342 329 -336
rect 330 -342 333 -336
rect 337 -342 343 -336
rect 344 -342 347 -336
rect 351 -342 357 -336
rect 358 -342 364 -336
rect 365 -342 368 -336
rect 372 -342 375 -336
rect 379 -342 382 -336
rect 386 -342 392 -336
rect 393 -342 396 -336
rect 400 -342 403 -336
rect 407 -342 410 -336
rect 414 -342 417 -336
rect 421 -342 424 -336
rect 428 -342 431 -336
rect 435 -342 438 -336
rect 442 -342 445 -336
rect 449 -342 452 -336
rect 456 -342 459 -336
rect 463 -342 466 -336
rect 470 -342 473 -336
rect 477 -342 480 -336
rect 484 -342 487 -336
rect 491 -342 497 -336
rect 498 -342 501 -336
rect 505 -342 508 -336
rect 512 -342 515 -336
rect 519 -342 522 -336
rect 526 -342 529 -336
rect 533 -342 536 -336
rect 540 -342 543 -336
rect 547 -342 550 -336
rect 554 -342 557 -336
rect 561 -342 564 -336
rect 568 -342 571 -336
rect 575 -342 578 -336
rect 582 -342 585 -336
rect 589 -342 592 -336
rect 603 -342 606 -336
rect 610 -342 613 -336
rect 617 -342 620 -336
rect 624 -342 627 -336
rect 631 -342 634 -336
rect 638 -342 641 -336
rect 645 -342 648 -336
rect 652 -342 655 -336
rect 659 -342 662 -336
rect 666 -342 669 -336
rect 673 -342 676 -336
rect 708 -342 711 -336
rect 1 -409 7 -403
rect 8 -409 14 -403
rect 22 -409 25 -403
rect 29 -409 35 -403
rect 36 -409 39 -403
rect 43 -409 46 -403
rect 50 -409 53 -403
rect 57 -409 60 -403
rect 64 -409 70 -403
rect 71 -409 74 -403
rect 78 -409 81 -403
rect 85 -409 88 -403
rect 92 -409 98 -403
rect 99 -409 102 -403
rect 106 -409 112 -403
rect 113 -409 119 -403
rect 120 -409 126 -403
rect 127 -409 130 -403
rect 134 -409 137 -403
rect 141 -409 144 -403
rect 148 -409 151 -403
rect 155 -409 161 -403
rect 162 -409 165 -403
rect 169 -409 172 -403
rect 176 -409 179 -403
rect 183 -409 189 -403
rect 190 -409 193 -403
rect 197 -409 200 -403
rect 204 -409 207 -403
rect 211 -409 214 -403
rect 218 -409 221 -403
rect 225 -409 231 -403
rect 232 -409 235 -403
rect 239 -409 245 -403
rect 246 -409 249 -403
rect 253 -409 256 -403
rect 260 -409 263 -403
rect 267 -409 270 -403
rect 274 -409 277 -403
rect 281 -409 287 -403
rect 288 -409 291 -403
rect 295 -409 298 -403
rect 302 -409 305 -403
rect 309 -409 312 -403
rect 316 -409 319 -403
rect 323 -409 329 -403
rect 330 -409 336 -403
rect 337 -409 343 -403
rect 344 -409 347 -403
rect 351 -409 357 -403
rect 358 -409 361 -403
rect 365 -409 368 -403
rect 372 -409 378 -403
rect 379 -409 385 -403
rect 386 -409 392 -403
rect 393 -409 396 -403
rect 400 -409 403 -403
rect 407 -409 413 -403
rect 414 -409 417 -403
rect 421 -409 424 -403
rect 428 -409 434 -403
rect 435 -409 438 -403
rect 442 -409 445 -403
rect 449 -409 452 -403
rect 456 -409 459 -403
rect 463 -409 469 -403
rect 470 -409 473 -403
rect 477 -409 483 -403
rect 484 -409 487 -403
rect 491 -409 494 -403
rect 498 -409 504 -403
rect 505 -409 508 -403
rect 512 -409 515 -403
rect 519 -409 522 -403
rect 526 -409 529 -403
rect 533 -409 536 -403
rect 540 -409 543 -403
rect 547 -409 550 -403
rect 554 -409 557 -403
rect 561 -409 564 -403
rect 568 -409 571 -403
rect 575 -409 578 -403
rect 582 -409 585 -403
rect 589 -409 592 -403
rect 596 -409 599 -403
rect 603 -409 606 -403
rect 610 -409 613 -403
rect 617 -409 620 -403
rect 624 -409 627 -403
rect 631 -409 637 -403
rect 638 -409 641 -403
rect 645 -409 648 -403
rect 652 -409 658 -403
rect 659 -409 662 -403
rect 666 -409 669 -403
rect 715 -409 718 -403
rect 1 -474 7 -468
rect 8 -474 11 -468
rect 15 -474 18 -468
rect 22 -474 28 -468
rect 29 -474 32 -468
rect 36 -474 39 -468
rect 43 -474 46 -468
rect 50 -474 53 -468
rect 57 -474 60 -468
rect 64 -474 70 -468
rect 71 -474 77 -468
rect 78 -474 84 -468
rect 85 -474 88 -468
rect 92 -474 95 -468
rect 99 -474 105 -468
rect 106 -474 109 -468
rect 113 -474 116 -468
rect 120 -474 123 -468
rect 127 -474 130 -468
rect 134 -474 137 -468
rect 141 -474 147 -468
rect 148 -474 151 -468
rect 155 -474 158 -468
rect 162 -474 168 -468
rect 169 -474 175 -468
rect 176 -474 182 -468
rect 183 -474 189 -468
rect 190 -474 196 -468
rect 197 -474 200 -468
rect 204 -474 207 -468
rect 211 -474 214 -468
rect 218 -474 221 -468
rect 225 -474 228 -468
rect 232 -474 235 -468
rect 239 -474 242 -468
rect 246 -474 249 -468
rect 253 -474 256 -468
rect 260 -474 263 -468
rect 267 -474 270 -468
rect 274 -474 277 -468
rect 281 -474 284 -468
rect 288 -474 291 -468
rect 295 -474 298 -468
rect 302 -474 305 -468
rect 309 -474 315 -468
rect 316 -474 319 -468
rect 323 -474 326 -468
rect 330 -474 333 -468
rect 337 -474 340 -468
rect 344 -474 347 -468
rect 351 -474 354 -468
rect 358 -474 364 -468
rect 365 -474 371 -468
rect 372 -474 375 -468
rect 379 -474 385 -468
rect 386 -474 392 -468
rect 393 -474 399 -468
rect 400 -474 403 -468
rect 407 -474 413 -468
rect 414 -474 420 -468
rect 421 -474 427 -468
rect 428 -474 434 -468
rect 435 -474 441 -468
rect 442 -474 448 -468
rect 449 -474 455 -468
rect 456 -474 459 -468
rect 463 -474 466 -468
rect 470 -474 473 -468
rect 477 -474 480 -468
rect 484 -474 487 -468
rect 491 -474 494 -468
rect 498 -474 501 -468
rect 505 -474 508 -468
rect 512 -474 515 -468
rect 519 -474 522 -468
rect 526 -474 529 -468
rect 533 -474 536 -468
rect 540 -474 543 -468
rect 547 -474 550 -468
rect 554 -474 557 -468
rect 561 -474 564 -468
rect 568 -474 571 -468
rect 575 -474 578 -468
rect 582 -474 585 -468
rect 589 -474 592 -468
rect 596 -474 599 -468
rect 603 -474 606 -468
rect 610 -474 613 -468
rect 624 -474 627 -468
rect 631 -474 634 -468
rect 638 -474 641 -468
rect 645 -474 648 -468
rect 652 -474 655 -468
rect 666 -474 669 -468
rect 673 -474 676 -468
rect 680 -474 683 -468
rect 687 -474 690 -468
rect 694 -474 697 -468
rect 701 -474 704 -468
rect 708 -474 714 -468
rect 715 -474 721 -468
rect 722 -474 725 -468
rect 729 -474 732 -468
rect 1 -559 7 -553
rect 8 -559 14 -553
rect 15 -559 21 -553
rect 22 -559 25 -553
rect 29 -559 35 -553
rect 36 -559 42 -553
rect 43 -559 46 -553
rect 50 -559 56 -553
rect 57 -559 63 -553
rect 64 -559 70 -553
rect 71 -559 77 -553
rect 78 -559 81 -553
rect 85 -559 88 -553
rect 92 -559 95 -553
rect 99 -559 105 -553
rect 106 -559 109 -553
rect 113 -559 116 -553
rect 120 -559 126 -553
rect 127 -559 130 -553
rect 134 -559 137 -553
rect 141 -559 147 -553
rect 148 -559 154 -553
rect 155 -559 158 -553
rect 162 -559 168 -553
rect 169 -559 172 -553
rect 176 -559 182 -553
rect 183 -559 189 -553
rect 190 -559 193 -553
rect 197 -559 200 -553
rect 204 -559 207 -553
rect 211 -559 217 -553
rect 218 -559 221 -553
rect 225 -559 228 -553
rect 232 -559 238 -553
rect 239 -559 245 -553
rect 246 -559 249 -553
rect 253 -559 256 -553
rect 260 -559 263 -553
rect 267 -559 270 -553
rect 274 -559 277 -553
rect 281 -559 284 -553
rect 288 -559 291 -553
rect 295 -559 298 -553
rect 302 -559 308 -553
rect 309 -559 312 -553
rect 316 -559 322 -553
rect 323 -559 326 -553
rect 330 -559 333 -553
rect 337 -559 340 -553
rect 344 -559 347 -553
rect 351 -559 354 -553
rect 358 -559 361 -553
rect 365 -559 371 -553
rect 372 -559 375 -553
rect 379 -559 385 -553
rect 386 -559 389 -553
rect 393 -559 399 -553
rect 400 -559 403 -553
rect 407 -559 410 -553
rect 414 -559 417 -553
rect 421 -559 427 -553
rect 428 -559 434 -553
rect 435 -559 438 -553
rect 442 -559 448 -553
rect 449 -559 452 -553
rect 456 -559 459 -553
rect 463 -559 466 -553
rect 470 -559 473 -553
rect 477 -559 480 -553
rect 484 -559 487 -553
rect 491 -559 494 -553
rect 498 -559 501 -553
rect 505 -559 508 -553
rect 512 -559 515 -553
rect 519 -559 522 -553
rect 526 -559 529 -553
rect 533 -559 536 -553
rect 540 -559 543 -553
rect 547 -559 550 -553
rect 554 -559 557 -553
rect 561 -559 564 -553
rect 568 -559 571 -553
rect 575 -559 578 -553
rect 582 -559 585 -553
rect 589 -559 592 -553
rect 596 -559 599 -553
rect 603 -559 606 -553
rect 610 -559 613 -553
rect 617 -559 620 -553
rect 624 -559 627 -553
rect 631 -559 634 -553
rect 638 -559 641 -553
rect 645 -559 648 -553
rect 652 -559 655 -553
rect 659 -559 662 -553
rect 666 -559 669 -553
rect 673 -559 676 -553
rect 680 -559 683 -553
rect 687 -559 690 -553
rect 694 -559 697 -553
rect 701 -559 704 -553
rect 708 -559 711 -553
rect 715 -559 718 -553
rect 722 -559 725 -553
rect 729 -559 732 -553
rect 736 -559 739 -553
rect 743 -559 746 -553
rect 750 -559 753 -553
rect 778 -559 781 -553
rect 1 -652 7 -646
rect 8 -652 14 -646
rect 15 -652 18 -646
rect 22 -652 25 -646
rect 29 -652 35 -646
rect 36 -652 42 -646
rect 43 -652 49 -646
rect 50 -652 53 -646
rect 57 -652 60 -646
rect 64 -652 67 -646
rect 71 -652 74 -646
rect 78 -652 81 -646
rect 85 -652 88 -646
rect 92 -652 98 -646
rect 99 -652 102 -646
rect 106 -652 112 -646
rect 113 -652 119 -646
rect 120 -652 126 -646
rect 127 -652 133 -646
rect 134 -652 137 -646
rect 141 -652 147 -646
rect 148 -652 154 -646
rect 155 -652 158 -646
rect 162 -652 168 -646
rect 169 -652 172 -646
rect 176 -652 179 -646
rect 183 -652 189 -646
rect 190 -652 193 -646
rect 197 -652 200 -646
rect 204 -652 207 -646
rect 211 -652 214 -646
rect 218 -652 221 -646
rect 225 -652 228 -646
rect 232 -652 235 -646
rect 239 -652 242 -646
rect 246 -652 249 -646
rect 253 -652 256 -646
rect 260 -652 263 -646
rect 267 -652 270 -646
rect 274 -652 280 -646
rect 281 -652 284 -646
rect 288 -652 294 -646
rect 295 -652 298 -646
rect 302 -652 305 -646
rect 309 -652 312 -646
rect 316 -652 319 -646
rect 323 -652 326 -646
rect 330 -652 333 -646
rect 337 -652 340 -646
rect 344 -652 350 -646
rect 351 -652 357 -646
rect 358 -652 361 -646
rect 365 -652 371 -646
rect 372 -652 375 -646
rect 379 -652 382 -646
rect 386 -652 392 -646
rect 393 -652 399 -646
rect 400 -652 403 -646
rect 407 -652 413 -646
rect 414 -652 420 -646
rect 421 -652 427 -646
rect 428 -652 431 -646
rect 435 -652 438 -646
rect 442 -652 448 -646
rect 449 -652 452 -646
rect 456 -652 459 -646
rect 463 -652 466 -646
rect 470 -652 473 -646
rect 477 -652 480 -646
rect 484 -652 487 -646
rect 498 -652 501 -646
rect 505 -652 508 -646
rect 512 -652 518 -646
rect 519 -652 522 -646
rect 526 -652 529 -646
rect 533 -652 536 -646
rect 540 -652 543 -646
rect 547 -652 550 -646
rect 554 -652 557 -646
rect 561 -652 564 -646
rect 568 -652 571 -646
rect 575 -652 578 -646
rect 582 -652 585 -646
rect 589 -652 592 -646
rect 596 -652 599 -646
rect 603 -652 606 -646
rect 610 -652 613 -646
rect 617 -652 620 -646
rect 624 -652 627 -646
rect 631 -652 634 -646
rect 638 -652 641 -646
rect 645 -652 648 -646
rect 652 -652 655 -646
rect 659 -652 665 -646
rect 666 -652 669 -646
rect 673 -652 676 -646
rect 680 -652 683 -646
rect 687 -652 690 -646
rect 694 -652 697 -646
rect 701 -652 704 -646
rect 708 -652 711 -646
rect 715 -652 718 -646
rect 722 -652 725 -646
rect 729 -652 732 -646
rect 736 -652 739 -646
rect 806 -652 809 -646
rect 1 -733 7 -727
rect 8 -733 11 -727
rect 15 -733 18 -727
rect 22 -733 25 -727
rect 29 -733 32 -727
rect 36 -733 39 -727
rect 43 -733 46 -727
rect 50 -733 56 -727
rect 57 -733 63 -727
rect 64 -733 70 -727
rect 71 -733 77 -727
rect 78 -733 81 -727
rect 85 -733 88 -727
rect 92 -733 98 -727
rect 99 -733 102 -727
rect 106 -733 109 -727
rect 113 -733 119 -727
rect 120 -733 126 -727
rect 127 -733 130 -727
rect 134 -733 137 -727
rect 141 -733 144 -727
rect 148 -733 151 -727
rect 155 -733 161 -727
rect 162 -733 168 -727
rect 169 -733 175 -727
rect 176 -733 179 -727
rect 183 -733 186 -727
rect 190 -733 193 -727
rect 197 -733 200 -727
rect 204 -733 207 -727
rect 211 -733 214 -727
rect 218 -733 221 -727
rect 225 -733 228 -727
rect 232 -733 238 -727
rect 239 -733 245 -727
rect 246 -733 249 -727
rect 253 -733 259 -727
rect 260 -733 263 -727
rect 267 -733 270 -727
rect 274 -733 277 -727
rect 281 -733 284 -727
rect 288 -733 294 -727
rect 295 -733 298 -727
rect 302 -733 305 -727
rect 309 -733 312 -727
rect 316 -733 319 -727
rect 323 -733 326 -727
rect 330 -733 336 -727
rect 337 -733 340 -727
rect 344 -733 347 -727
rect 351 -733 354 -727
rect 358 -733 361 -727
rect 365 -733 371 -727
rect 372 -733 375 -727
rect 379 -733 382 -727
rect 386 -733 389 -727
rect 393 -733 399 -727
rect 400 -733 403 -727
rect 407 -733 413 -727
rect 414 -733 417 -727
rect 421 -733 424 -727
rect 428 -733 434 -727
rect 435 -733 441 -727
rect 442 -733 445 -727
rect 449 -733 455 -727
rect 456 -733 459 -727
rect 463 -733 469 -727
rect 470 -733 476 -727
rect 477 -733 480 -727
rect 484 -733 487 -727
rect 491 -733 494 -727
rect 498 -733 501 -727
rect 505 -733 508 -727
rect 512 -733 515 -727
rect 519 -733 522 -727
rect 526 -733 529 -727
rect 533 -733 536 -727
rect 540 -733 543 -727
rect 547 -733 550 -727
rect 554 -733 557 -727
rect 561 -733 564 -727
rect 568 -733 571 -727
rect 575 -733 578 -727
rect 582 -733 585 -727
rect 589 -733 592 -727
rect 596 -733 602 -727
rect 603 -733 606 -727
rect 610 -733 613 -727
rect 617 -733 620 -727
rect 624 -733 627 -727
rect 631 -733 634 -727
rect 638 -733 641 -727
rect 645 -733 648 -727
rect 652 -733 655 -727
rect 659 -733 662 -727
rect 666 -733 669 -727
rect 673 -733 676 -727
rect 680 -733 683 -727
rect 687 -733 690 -727
rect 694 -733 697 -727
rect 701 -733 704 -727
rect 708 -733 711 -727
rect 715 -733 718 -727
rect 722 -733 725 -727
rect 729 -733 732 -727
rect 736 -733 739 -727
rect 743 -733 746 -727
rect 750 -733 753 -727
rect 757 -733 760 -727
rect 764 -733 767 -727
rect 771 -733 774 -727
rect 778 -733 781 -727
rect 785 -733 788 -727
rect 792 -733 795 -727
rect 799 -733 802 -727
rect 806 -733 809 -727
rect 813 -733 819 -727
rect 820 -733 826 -727
rect 827 -733 830 -727
rect 1 -822 7 -816
rect 8 -822 11 -816
rect 15 -822 21 -816
rect 22 -822 25 -816
rect 29 -822 32 -816
rect 36 -822 42 -816
rect 43 -822 49 -816
rect 50 -822 56 -816
rect 57 -822 60 -816
rect 64 -822 70 -816
rect 71 -822 77 -816
rect 78 -822 84 -816
rect 85 -822 88 -816
rect 92 -822 98 -816
rect 99 -822 102 -816
rect 106 -822 109 -816
rect 113 -822 116 -816
rect 120 -822 123 -816
rect 127 -822 130 -816
rect 134 -822 137 -816
rect 141 -822 144 -816
rect 148 -822 154 -816
rect 155 -822 158 -816
rect 162 -822 165 -816
rect 169 -822 172 -816
rect 176 -822 179 -816
rect 183 -822 189 -816
rect 190 -822 193 -816
rect 197 -822 200 -816
rect 204 -822 207 -816
rect 211 -822 214 -816
rect 218 -822 221 -816
rect 225 -822 228 -816
rect 232 -822 235 -816
rect 239 -822 242 -816
rect 246 -822 249 -816
rect 253 -822 256 -816
rect 260 -822 263 -816
rect 267 -822 273 -816
rect 274 -822 277 -816
rect 281 -822 284 -816
rect 288 -822 291 -816
rect 295 -822 298 -816
rect 302 -822 308 -816
rect 309 -822 312 -816
rect 316 -822 319 -816
rect 323 -822 326 -816
rect 330 -822 336 -816
rect 337 -822 343 -816
rect 344 -822 350 -816
rect 351 -822 357 -816
rect 358 -822 361 -816
rect 365 -822 371 -816
rect 372 -822 375 -816
rect 379 -822 385 -816
rect 386 -822 392 -816
rect 393 -822 396 -816
rect 400 -822 406 -816
rect 407 -822 410 -816
rect 414 -822 417 -816
rect 421 -822 424 -816
rect 428 -822 434 -816
rect 435 -822 441 -816
rect 442 -822 448 -816
rect 449 -822 455 -816
rect 456 -822 459 -816
rect 463 -822 466 -816
rect 470 -822 473 -816
rect 477 -822 480 -816
rect 484 -822 487 -816
rect 491 -822 494 -816
rect 498 -822 501 -816
rect 505 -822 508 -816
rect 512 -822 515 -816
rect 519 -822 522 -816
rect 526 -822 529 -816
rect 533 -822 536 -816
rect 540 -822 543 -816
rect 547 -822 550 -816
rect 554 -822 560 -816
rect 561 -822 564 -816
rect 568 -822 571 -816
rect 575 -822 578 -816
rect 582 -822 585 -816
rect 589 -822 595 -816
rect 596 -822 599 -816
rect 603 -822 606 -816
rect 610 -822 613 -816
rect 617 -822 620 -816
rect 624 -822 627 -816
rect 631 -822 634 -816
rect 638 -822 641 -816
rect 645 -822 648 -816
rect 652 -822 655 -816
rect 659 -822 662 -816
rect 666 -822 669 -816
rect 673 -822 676 -816
rect 680 -822 683 -816
rect 687 -822 690 -816
rect 694 -822 697 -816
rect 701 -822 704 -816
rect 708 -822 711 -816
rect 715 -822 718 -816
rect 722 -822 725 -816
rect 729 -822 732 -816
rect 736 -822 739 -816
rect 743 -822 746 -816
rect 750 -822 753 -816
rect 757 -822 760 -816
rect 764 -822 767 -816
rect 771 -822 774 -816
rect 778 -822 781 -816
rect 785 -822 788 -816
rect 792 -822 795 -816
rect 1 -907 7 -901
rect 8 -907 14 -901
rect 15 -907 18 -901
rect 22 -907 28 -901
rect 29 -907 32 -901
rect 36 -907 42 -901
rect 43 -907 46 -901
rect 50 -907 56 -901
rect 57 -907 60 -901
rect 64 -907 67 -901
rect 71 -907 74 -901
rect 78 -907 81 -901
rect 85 -907 88 -901
rect 92 -907 95 -901
rect 99 -907 105 -901
rect 106 -907 109 -901
rect 113 -907 119 -901
rect 120 -907 123 -901
rect 127 -907 130 -901
rect 134 -907 140 -901
rect 141 -907 147 -901
rect 148 -907 151 -901
rect 155 -907 158 -901
rect 162 -907 165 -901
rect 169 -907 175 -901
rect 176 -907 182 -901
rect 183 -907 186 -901
rect 190 -907 193 -901
rect 197 -907 200 -901
rect 204 -907 207 -901
rect 211 -907 214 -901
rect 218 -907 221 -901
rect 225 -907 228 -901
rect 232 -907 235 -901
rect 239 -907 242 -901
rect 246 -907 249 -901
rect 253 -907 259 -901
rect 260 -907 263 -901
rect 267 -907 270 -901
rect 274 -907 280 -901
rect 281 -907 287 -901
rect 288 -907 294 -901
rect 295 -907 301 -901
rect 302 -907 308 -901
rect 309 -907 312 -901
rect 316 -907 319 -901
rect 323 -907 326 -901
rect 330 -907 333 -901
rect 337 -907 343 -901
rect 344 -907 347 -901
rect 351 -907 354 -901
rect 358 -907 364 -901
rect 365 -907 368 -901
rect 372 -907 375 -901
rect 379 -907 382 -901
rect 386 -907 389 -901
rect 393 -907 396 -901
rect 400 -907 406 -901
rect 407 -907 413 -901
rect 414 -907 417 -901
rect 421 -907 424 -901
rect 428 -907 431 -901
rect 435 -907 438 -901
rect 442 -907 445 -901
rect 449 -907 455 -901
rect 456 -907 459 -901
rect 463 -907 466 -901
rect 470 -907 473 -901
rect 477 -907 480 -901
rect 484 -907 487 -901
rect 491 -907 494 -901
rect 498 -907 501 -901
rect 505 -907 511 -901
rect 512 -907 515 -901
rect 519 -907 522 -901
rect 526 -907 532 -901
rect 533 -907 539 -901
rect 540 -907 543 -901
rect 554 -907 557 -901
rect 561 -907 564 -901
rect 568 -907 571 -901
rect 575 -907 578 -901
rect 582 -907 585 -901
rect 589 -907 595 -901
rect 596 -907 599 -901
rect 603 -907 606 -901
rect 617 -907 620 -901
rect 624 -907 627 -901
rect 631 -907 634 -901
rect 638 -907 641 -901
rect 645 -907 648 -901
rect 652 -907 655 -901
rect 659 -907 662 -901
rect 666 -907 669 -901
rect 673 -907 676 -901
rect 680 -907 683 -901
rect 687 -907 690 -901
rect 694 -907 700 -901
rect 701 -907 704 -901
rect 708 -907 711 -901
rect 736 -907 739 -901
rect 757 -907 760 -901
rect 1 -990 4 -984
rect 8 -990 14 -984
rect 15 -990 18 -984
rect 22 -990 28 -984
rect 29 -990 32 -984
rect 36 -990 39 -984
rect 43 -990 49 -984
rect 50 -990 56 -984
rect 57 -990 63 -984
rect 64 -990 70 -984
rect 71 -990 74 -984
rect 78 -990 81 -984
rect 85 -990 91 -984
rect 92 -990 95 -984
rect 99 -990 102 -984
rect 106 -990 112 -984
rect 113 -990 116 -984
rect 120 -990 123 -984
rect 127 -990 130 -984
rect 134 -990 140 -984
rect 141 -990 147 -984
rect 148 -990 154 -984
rect 155 -990 158 -984
rect 162 -990 165 -984
rect 169 -990 172 -984
rect 176 -990 182 -984
rect 183 -990 189 -984
rect 190 -990 193 -984
rect 197 -990 200 -984
rect 204 -990 207 -984
rect 211 -990 214 -984
rect 218 -990 221 -984
rect 225 -990 231 -984
rect 232 -990 235 -984
rect 239 -990 242 -984
rect 246 -990 252 -984
rect 253 -990 256 -984
rect 260 -990 263 -984
rect 267 -990 270 -984
rect 274 -990 277 -984
rect 281 -990 284 -984
rect 288 -990 294 -984
rect 295 -990 298 -984
rect 302 -990 305 -984
rect 309 -990 315 -984
rect 316 -990 319 -984
rect 323 -990 326 -984
rect 330 -990 333 -984
rect 337 -990 340 -984
rect 344 -990 347 -984
rect 351 -990 354 -984
rect 358 -990 364 -984
rect 365 -990 368 -984
rect 372 -990 375 -984
rect 379 -990 385 -984
rect 386 -990 389 -984
rect 393 -990 399 -984
rect 400 -990 403 -984
rect 407 -990 413 -984
rect 414 -990 417 -984
rect 421 -990 424 -984
rect 428 -990 431 -984
rect 435 -990 438 -984
rect 442 -990 448 -984
rect 449 -990 452 -984
rect 456 -990 459 -984
rect 463 -990 466 -984
rect 470 -990 473 -984
rect 477 -990 480 -984
rect 484 -990 490 -984
rect 491 -990 494 -984
rect 498 -990 504 -984
rect 505 -990 508 -984
rect 512 -990 515 -984
rect 519 -990 522 -984
rect 526 -990 529 -984
rect 533 -990 536 -984
rect 540 -990 543 -984
rect 547 -990 550 -984
rect 554 -990 557 -984
rect 561 -990 564 -984
rect 568 -990 571 -984
rect 575 -990 578 -984
rect 582 -990 585 -984
rect 589 -990 592 -984
rect 603 -990 609 -984
rect 610 -990 613 -984
rect 617 -990 623 -984
rect 624 -990 627 -984
rect 631 -990 634 -984
rect 638 -990 641 -984
rect 645 -990 648 -984
rect 652 -990 655 -984
rect 659 -990 662 -984
rect 666 -990 669 -984
rect 673 -990 676 -984
rect 680 -990 683 -984
rect 687 -990 690 -984
rect 694 -990 697 -984
rect 701 -990 704 -984
rect 708 -990 711 -984
rect 715 -990 718 -984
rect 722 -990 728 -984
rect 750 -990 753 -984
rect 8 -1065 14 -1059
rect 15 -1065 18 -1059
rect 22 -1065 28 -1059
rect 29 -1065 35 -1059
rect 36 -1065 39 -1059
rect 43 -1065 49 -1059
rect 50 -1065 56 -1059
rect 57 -1065 60 -1059
rect 64 -1065 67 -1059
rect 71 -1065 77 -1059
rect 78 -1065 81 -1059
rect 85 -1065 88 -1059
rect 92 -1065 95 -1059
rect 99 -1065 105 -1059
rect 106 -1065 109 -1059
rect 113 -1065 119 -1059
rect 120 -1065 123 -1059
rect 127 -1065 130 -1059
rect 134 -1065 140 -1059
rect 141 -1065 144 -1059
rect 148 -1065 151 -1059
rect 155 -1065 158 -1059
rect 162 -1065 165 -1059
rect 169 -1065 175 -1059
rect 176 -1065 179 -1059
rect 183 -1065 189 -1059
rect 190 -1065 193 -1059
rect 197 -1065 200 -1059
rect 204 -1065 207 -1059
rect 211 -1065 214 -1059
rect 218 -1065 221 -1059
rect 225 -1065 228 -1059
rect 232 -1065 235 -1059
rect 239 -1065 242 -1059
rect 246 -1065 249 -1059
rect 253 -1065 256 -1059
rect 260 -1065 263 -1059
rect 267 -1065 273 -1059
rect 274 -1065 277 -1059
rect 281 -1065 287 -1059
rect 288 -1065 291 -1059
rect 295 -1065 298 -1059
rect 302 -1065 308 -1059
rect 309 -1065 315 -1059
rect 316 -1065 322 -1059
rect 323 -1065 326 -1059
rect 330 -1065 333 -1059
rect 337 -1065 340 -1059
rect 344 -1065 347 -1059
rect 351 -1065 357 -1059
rect 358 -1065 364 -1059
rect 365 -1065 371 -1059
rect 372 -1065 378 -1059
rect 379 -1065 382 -1059
rect 386 -1065 389 -1059
rect 393 -1065 399 -1059
rect 400 -1065 406 -1059
rect 407 -1065 410 -1059
rect 414 -1065 420 -1059
rect 421 -1065 427 -1059
rect 428 -1065 431 -1059
rect 435 -1065 438 -1059
rect 442 -1065 445 -1059
rect 449 -1065 455 -1059
rect 456 -1065 459 -1059
rect 463 -1065 466 -1059
rect 470 -1065 473 -1059
rect 477 -1065 480 -1059
rect 484 -1065 487 -1059
rect 491 -1065 494 -1059
rect 498 -1065 501 -1059
rect 505 -1065 508 -1059
rect 512 -1065 515 -1059
rect 519 -1065 522 -1059
rect 526 -1065 529 -1059
rect 533 -1065 536 -1059
rect 540 -1065 543 -1059
rect 547 -1065 550 -1059
rect 554 -1065 557 -1059
rect 561 -1065 564 -1059
rect 568 -1065 571 -1059
rect 575 -1065 578 -1059
rect 582 -1065 585 -1059
rect 589 -1065 592 -1059
rect 596 -1065 599 -1059
rect 603 -1065 609 -1059
rect 610 -1065 613 -1059
rect 617 -1065 620 -1059
rect 624 -1065 627 -1059
rect 631 -1065 634 -1059
rect 638 -1065 641 -1059
rect 645 -1065 648 -1059
rect 652 -1065 655 -1059
rect 659 -1065 662 -1059
rect 666 -1065 669 -1059
rect 673 -1065 676 -1059
rect 680 -1065 683 -1059
rect 687 -1065 690 -1059
rect 694 -1065 697 -1059
rect 701 -1065 704 -1059
rect 708 -1065 711 -1059
rect 715 -1065 718 -1059
rect 722 -1065 725 -1059
rect 729 -1065 732 -1059
rect 750 -1065 756 -1059
rect 757 -1065 760 -1059
rect 8 -1132 11 -1126
rect 15 -1132 18 -1126
rect 22 -1132 28 -1126
rect 36 -1132 39 -1126
rect 43 -1132 46 -1126
rect 50 -1132 53 -1126
rect 57 -1132 60 -1126
rect 64 -1132 67 -1126
rect 71 -1132 74 -1126
rect 78 -1132 81 -1126
rect 85 -1132 91 -1126
rect 92 -1132 95 -1126
rect 99 -1132 102 -1126
rect 106 -1132 109 -1126
rect 113 -1132 119 -1126
rect 120 -1132 123 -1126
rect 127 -1132 130 -1126
rect 134 -1132 140 -1126
rect 141 -1132 144 -1126
rect 148 -1132 154 -1126
rect 155 -1132 158 -1126
rect 162 -1132 168 -1126
rect 169 -1132 172 -1126
rect 176 -1132 182 -1126
rect 183 -1132 189 -1126
rect 190 -1132 196 -1126
rect 197 -1132 200 -1126
rect 204 -1132 210 -1126
rect 211 -1132 214 -1126
rect 218 -1132 221 -1126
rect 225 -1132 228 -1126
rect 232 -1132 238 -1126
rect 239 -1132 242 -1126
rect 246 -1132 252 -1126
rect 253 -1132 256 -1126
rect 260 -1132 263 -1126
rect 267 -1132 270 -1126
rect 274 -1132 277 -1126
rect 281 -1132 287 -1126
rect 288 -1132 294 -1126
rect 295 -1132 298 -1126
rect 302 -1132 305 -1126
rect 309 -1132 312 -1126
rect 316 -1132 322 -1126
rect 323 -1132 329 -1126
rect 330 -1132 333 -1126
rect 337 -1132 340 -1126
rect 344 -1132 347 -1126
rect 351 -1132 357 -1126
rect 358 -1132 361 -1126
rect 365 -1132 371 -1126
rect 372 -1132 375 -1126
rect 379 -1132 385 -1126
rect 386 -1132 389 -1126
rect 393 -1132 396 -1126
rect 400 -1132 403 -1126
rect 407 -1132 410 -1126
rect 414 -1132 417 -1126
rect 421 -1132 427 -1126
rect 428 -1132 434 -1126
rect 435 -1132 441 -1126
rect 442 -1132 445 -1126
rect 449 -1132 452 -1126
rect 456 -1132 459 -1126
rect 463 -1132 466 -1126
rect 470 -1132 476 -1126
rect 477 -1132 480 -1126
rect 484 -1132 487 -1126
rect 491 -1132 494 -1126
rect 498 -1132 501 -1126
rect 505 -1132 511 -1126
rect 512 -1132 515 -1126
rect 519 -1132 522 -1126
rect 526 -1132 529 -1126
rect 533 -1132 536 -1126
rect 540 -1132 543 -1126
rect 547 -1132 550 -1126
rect 554 -1132 557 -1126
rect 561 -1132 564 -1126
rect 568 -1132 571 -1126
rect 575 -1132 578 -1126
rect 582 -1132 585 -1126
rect 589 -1132 592 -1126
rect 596 -1132 599 -1126
rect 603 -1132 606 -1126
rect 624 -1132 627 -1126
rect 631 -1132 634 -1126
rect 638 -1132 641 -1126
rect 645 -1132 648 -1126
rect 652 -1132 655 -1126
rect 659 -1132 662 -1126
rect 666 -1132 669 -1126
rect 673 -1132 676 -1126
rect 680 -1132 683 -1126
rect 694 -1132 697 -1126
rect 701 -1132 704 -1126
rect 708 -1132 711 -1126
rect 715 -1132 718 -1126
rect 722 -1132 725 -1126
rect 729 -1132 732 -1126
rect 736 -1132 742 -1126
rect 743 -1132 749 -1126
rect 750 -1132 756 -1126
rect 757 -1132 760 -1126
rect 778 -1132 781 -1126
rect 785 -1132 788 -1126
rect 792 -1132 795 -1126
rect 813 -1132 816 -1126
rect 8 -1213 11 -1207
rect 15 -1213 18 -1207
rect 22 -1213 25 -1207
rect 29 -1213 35 -1207
rect 36 -1213 42 -1207
rect 43 -1213 46 -1207
rect 50 -1213 56 -1207
rect 57 -1213 60 -1207
rect 64 -1213 70 -1207
rect 71 -1213 74 -1207
rect 78 -1213 81 -1207
rect 85 -1213 91 -1207
rect 92 -1213 95 -1207
rect 99 -1213 102 -1207
rect 106 -1213 109 -1207
rect 113 -1213 119 -1207
rect 120 -1213 123 -1207
rect 127 -1213 130 -1207
rect 134 -1213 137 -1207
rect 141 -1213 147 -1207
rect 148 -1213 151 -1207
rect 155 -1213 158 -1207
rect 162 -1213 168 -1207
rect 169 -1213 172 -1207
rect 176 -1213 179 -1207
rect 183 -1213 189 -1207
rect 190 -1213 193 -1207
rect 197 -1213 200 -1207
rect 204 -1213 207 -1207
rect 211 -1213 214 -1207
rect 218 -1213 221 -1207
rect 225 -1213 228 -1207
rect 232 -1213 238 -1207
rect 239 -1213 242 -1207
rect 246 -1213 249 -1207
rect 253 -1213 259 -1207
rect 260 -1213 263 -1207
rect 267 -1213 270 -1207
rect 274 -1213 280 -1207
rect 281 -1213 284 -1207
rect 288 -1213 291 -1207
rect 295 -1213 298 -1207
rect 302 -1213 305 -1207
rect 309 -1213 312 -1207
rect 316 -1213 322 -1207
rect 323 -1213 329 -1207
rect 330 -1213 333 -1207
rect 337 -1213 343 -1207
rect 344 -1213 350 -1207
rect 351 -1213 354 -1207
rect 358 -1213 361 -1207
rect 365 -1213 371 -1207
rect 372 -1213 375 -1207
rect 379 -1213 382 -1207
rect 386 -1213 392 -1207
rect 393 -1213 399 -1207
rect 400 -1213 406 -1207
rect 407 -1213 413 -1207
rect 414 -1213 417 -1207
rect 421 -1213 424 -1207
rect 428 -1213 431 -1207
rect 435 -1213 438 -1207
rect 442 -1213 445 -1207
rect 449 -1213 452 -1207
rect 456 -1213 459 -1207
rect 463 -1213 469 -1207
rect 470 -1213 476 -1207
rect 477 -1213 483 -1207
rect 484 -1213 487 -1207
rect 491 -1213 494 -1207
rect 498 -1213 501 -1207
rect 505 -1213 508 -1207
rect 512 -1213 515 -1207
rect 519 -1213 522 -1207
rect 526 -1213 529 -1207
rect 533 -1213 536 -1207
rect 540 -1213 546 -1207
rect 547 -1213 550 -1207
rect 554 -1213 557 -1207
rect 561 -1213 564 -1207
rect 568 -1213 571 -1207
rect 575 -1213 578 -1207
rect 582 -1213 585 -1207
rect 589 -1213 595 -1207
rect 596 -1213 599 -1207
rect 603 -1213 606 -1207
rect 610 -1213 613 -1207
rect 617 -1213 620 -1207
rect 624 -1213 627 -1207
rect 631 -1213 634 -1207
rect 638 -1213 641 -1207
rect 645 -1213 648 -1207
rect 652 -1213 655 -1207
rect 659 -1213 665 -1207
rect 666 -1213 669 -1207
rect 673 -1213 676 -1207
rect 680 -1213 683 -1207
rect 687 -1213 690 -1207
rect 694 -1213 697 -1207
rect 701 -1213 704 -1207
rect 708 -1213 711 -1207
rect 715 -1213 718 -1207
rect 722 -1213 725 -1207
rect 729 -1213 732 -1207
rect 743 -1213 746 -1207
rect 750 -1213 753 -1207
rect 757 -1213 760 -1207
rect 764 -1213 767 -1207
rect 771 -1213 774 -1207
rect 778 -1213 781 -1207
rect 785 -1213 788 -1207
rect 792 -1213 795 -1207
rect 799 -1213 802 -1207
rect 1 -1306 4 -1300
rect 8 -1306 11 -1300
rect 15 -1306 18 -1300
rect 22 -1306 25 -1300
rect 29 -1306 32 -1300
rect 36 -1306 39 -1300
rect 43 -1306 46 -1300
rect 50 -1306 53 -1300
rect 57 -1306 60 -1300
rect 64 -1306 70 -1300
rect 71 -1306 77 -1300
rect 78 -1306 81 -1300
rect 85 -1306 88 -1300
rect 92 -1306 95 -1300
rect 99 -1306 102 -1300
rect 106 -1306 109 -1300
rect 113 -1306 119 -1300
rect 120 -1306 123 -1300
rect 127 -1306 130 -1300
rect 134 -1306 137 -1300
rect 141 -1306 147 -1300
rect 148 -1306 151 -1300
rect 155 -1306 158 -1300
rect 162 -1306 168 -1300
rect 169 -1306 172 -1300
rect 176 -1306 179 -1300
rect 183 -1306 189 -1300
rect 190 -1306 193 -1300
rect 197 -1306 203 -1300
rect 204 -1306 207 -1300
rect 211 -1306 214 -1300
rect 218 -1306 221 -1300
rect 225 -1306 231 -1300
rect 232 -1306 235 -1300
rect 239 -1306 242 -1300
rect 246 -1306 249 -1300
rect 253 -1306 256 -1300
rect 260 -1306 263 -1300
rect 267 -1306 270 -1300
rect 274 -1306 277 -1300
rect 281 -1306 284 -1300
rect 288 -1306 291 -1300
rect 295 -1306 298 -1300
rect 302 -1306 308 -1300
rect 309 -1306 315 -1300
rect 316 -1306 319 -1300
rect 323 -1306 326 -1300
rect 330 -1306 336 -1300
rect 337 -1306 343 -1300
rect 344 -1306 347 -1300
rect 351 -1306 357 -1300
rect 358 -1306 364 -1300
rect 365 -1306 371 -1300
rect 372 -1306 375 -1300
rect 379 -1306 382 -1300
rect 386 -1306 389 -1300
rect 393 -1306 396 -1300
rect 400 -1306 406 -1300
rect 407 -1306 413 -1300
rect 414 -1306 417 -1300
rect 421 -1306 427 -1300
rect 428 -1306 431 -1300
rect 435 -1306 438 -1300
rect 442 -1306 445 -1300
rect 449 -1306 455 -1300
rect 456 -1306 462 -1300
rect 463 -1306 466 -1300
rect 470 -1306 473 -1300
rect 477 -1306 480 -1300
rect 484 -1306 487 -1300
rect 491 -1306 494 -1300
rect 498 -1306 501 -1300
rect 505 -1306 508 -1300
rect 512 -1306 515 -1300
rect 519 -1306 522 -1300
rect 526 -1306 529 -1300
rect 533 -1306 539 -1300
rect 540 -1306 543 -1300
rect 547 -1306 550 -1300
rect 554 -1306 557 -1300
rect 561 -1306 564 -1300
rect 568 -1306 574 -1300
rect 575 -1306 578 -1300
rect 582 -1306 585 -1300
rect 589 -1306 592 -1300
rect 596 -1306 599 -1300
rect 603 -1306 606 -1300
rect 610 -1306 613 -1300
rect 617 -1306 620 -1300
rect 624 -1306 627 -1300
rect 631 -1306 634 -1300
rect 638 -1306 641 -1300
rect 645 -1306 651 -1300
rect 652 -1306 655 -1300
rect 659 -1306 662 -1300
rect 666 -1306 669 -1300
rect 673 -1306 676 -1300
rect 680 -1306 683 -1300
rect 687 -1306 690 -1300
rect 694 -1306 697 -1300
rect 701 -1306 704 -1300
rect 708 -1306 711 -1300
rect 715 -1306 718 -1300
rect 722 -1306 725 -1300
rect 729 -1306 732 -1300
rect 736 -1306 739 -1300
rect 743 -1306 746 -1300
rect 750 -1306 753 -1300
rect 757 -1306 760 -1300
rect 764 -1306 770 -1300
rect 771 -1306 777 -1300
rect 778 -1306 784 -1300
rect 785 -1306 791 -1300
rect 8 -1383 14 -1377
rect 22 -1383 25 -1377
rect 29 -1383 32 -1377
rect 36 -1383 42 -1377
rect 43 -1383 46 -1377
rect 50 -1383 53 -1377
rect 57 -1383 60 -1377
rect 64 -1383 67 -1377
rect 71 -1383 77 -1377
rect 78 -1383 84 -1377
rect 85 -1383 91 -1377
rect 92 -1383 98 -1377
rect 99 -1383 102 -1377
rect 106 -1383 109 -1377
rect 113 -1383 119 -1377
rect 120 -1383 123 -1377
rect 127 -1383 130 -1377
rect 134 -1383 137 -1377
rect 141 -1383 147 -1377
rect 148 -1383 151 -1377
rect 155 -1383 158 -1377
rect 162 -1383 168 -1377
rect 169 -1383 172 -1377
rect 176 -1383 182 -1377
rect 183 -1383 189 -1377
rect 190 -1383 193 -1377
rect 197 -1383 200 -1377
rect 204 -1383 207 -1377
rect 211 -1383 217 -1377
rect 218 -1383 221 -1377
rect 225 -1383 228 -1377
rect 232 -1383 235 -1377
rect 239 -1383 242 -1377
rect 246 -1383 249 -1377
rect 253 -1383 256 -1377
rect 260 -1383 263 -1377
rect 267 -1383 270 -1377
rect 274 -1383 280 -1377
rect 281 -1383 284 -1377
rect 288 -1383 291 -1377
rect 295 -1383 301 -1377
rect 302 -1383 305 -1377
rect 309 -1383 312 -1377
rect 316 -1383 322 -1377
rect 323 -1383 326 -1377
rect 330 -1383 336 -1377
rect 337 -1383 340 -1377
rect 344 -1383 350 -1377
rect 351 -1383 354 -1377
rect 358 -1383 361 -1377
rect 365 -1383 368 -1377
rect 372 -1383 375 -1377
rect 379 -1383 382 -1377
rect 386 -1383 389 -1377
rect 393 -1383 396 -1377
rect 400 -1383 406 -1377
rect 407 -1383 413 -1377
rect 414 -1383 417 -1377
rect 421 -1383 424 -1377
rect 428 -1383 431 -1377
rect 435 -1383 438 -1377
rect 442 -1383 448 -1377
rect 449 -1383 452 -1377
rect 456 -1383 459 -1377
rect 463 -1383 466 -1377
rect 470 -1383 473 -1377
rect 477 -1383 483 -1377
rect 484 -1383 487 -1377
rect 491 -1383 494 -1377
rect 498 -1383 501 -1377
rect 505 -1383 508 -1377
rect 512 -1383 518 -1377
rect 519 -1383 522 -1377
rect 526 -1383 529 -1377
rect 533 -1383 536 -1377
rect 540 -1383 543 -1377
rect 547 -1383 550 -1377
rect 554 -1383 557 -1377
rect 561 -1383 567 -1377
rect 568 -1383 574 -1377
rect 575 -1383 578 -1377
rect 582 -1383 585 -1377
rect 589 -1383 592 -1377
rect 596 -1383 599 -1377
rect 603 -1383 606 -1377
rect 610 -1383 613 -1377
rect 617 -1383 620 -1377
rect 631 -1383 634 -1377
rect 638 -1383 641 -1377
rect 645 -1383 648 -1377
rect 652 -1383 655 -1377
rect 659 -1383 662 -1377
rect 666 -1383 669 -1377
rect 673 -1383 676 -1377
rect 680 -1383 683 -1377
rect 687 -1383 693 -1377
rect 694 -1383 697 -1377
rect 701 -1383 707 -1377
rect 708 -1383 711 -1377
rect 715 -1383 721 -1377
rect 757 -1383 760 -1377
rect 778 -1383 781 -1377
rect 799 -1383 802 -1377
rect 8 -1452 11 -1446
rect 15 -1452 18 -1446
rect 22 -1452 25 -1446
rect 29 -1452 32 -1446
rect 36 -1452 39 -1446
rect 43 -1452 46 -1446
rect 50 -1452 56 -1446
rect 57 -1452 60 -1446
rect 64 -1452 67 -1446
rect 71 -1452 77 -1446
rect 78 -1452 81 -1446
rect 85 -1452 88 -1446
rect 92 -1452 95 -1446
rect 99 -1452 105 -1446
rect 106 -1452 109 -1446
rect 113 -1452 119 -1446
rect 120 -1452 126 -1446
rect 127 -1452 130 -1446
rect 134 -1452 140 -1446
rect 141 -1452 144 -1446
rect 148 -1452 151 -1446
rect 155 -1452 161 -1446
rect 162 -1452 165 -1446
rect 169 -1452 172 -1446
rect 176 -1452 179 -1446
rect 183 -1452 189 -1446
rect 190 -1452 193 -1446
rect 197 -1452 200 -1446
rect 204 -1452 207 -1446
rect 211 -1452 214 -1446
rect 218 -1452 221 -1446
rect 225 -1452 228 -1446
rect 232 -1452 235 -1446
rect 239 -1452 242 -1446
rect 246 -1452 249 -1446
rect 253 -1452 259 -1446
rect 260 -1452 263 -1446
rect 267 -1452 273 -1446
rect 274 -1452 277 -1446
rect 281 -1452 284 -1446
rect 288 -1452 291 -1446
rect 295 -1452 298 -1446
rect 302 -1452 305 -1446
rect 309 -1452 312 -1446
rect 316 -1452 319 -1446
rect 323 -1452 326 -1446
rect 330 -1452 336 -1446
rect 337 -1452 340 -1446
rect 344 -1452 347 -1446
rect 351 -1452 354 -1446
rect 358 -1452 361 -1446
rect 365 -1452 368 -1446
rect 372 -1452 375 -1446
rect 379 -1452 385 -1446
rect 386 -1452 389 -1446
rect 393 -1452 399 -1446
rect 400 -1452 406 -1446
rect 407 -1452 413 -1446
rect 414 -1452 417 -1446
rect 421 -1452 424 -1446
rect 428 -1452 434 -1446
rect 435 -1452 441 -1446
rect 442 -1452 445 -1446
rect 449 -1452 452 -1446
rect 456 -1452 459 -1446
rect 463 -1452 466 -1446
rect 470 -1452 476 -1446
rect 477 -1452 480 -1446
rect 484 -1452 490 -1446
rect 491 -1452 494 -1446
rect 498 -1452 501 -1446
rect 505 -1452 511 -1446
rect 512 -1452 515 -1446
rect 519 -1452 522 -1446
rect 526 -1452 529 -1446
rect 533 -1452 536 -1446
rect 540 -1452 543 -1446
rect 547 -1452 553 -1446
rect 554 -1452 557 -1446
rect 561 -1452 564 -1446
rect 568 -1452 571 -1446
rect 575 -1452 578 -1446
rect 582 -1452 585 -1446
rect 589 -1452 592 -1446
rect 596 -1452 599 -1446
rect 603 -1452 606 -1446
rect 610 -1452 613 -1446
rect 617 -1452 620 -1446
rect 624 -1452 627 -1446
rect 631 -1452 634 -1446
rect 638 -1452 641 -1446
rect 645 -1452 648 -1446
rect 652 -1452 655 -1446
rect 659 -1452 662 -1446
rect 666 -1452 669 -1446
rect 673 -1452 676 -1446
rect 680 -1452 683 -1446
rect 687 -1452 690 -1446
rect 694 -1452 697 -1446
rect 701 -1452 704 -1446
rect 708 -1452 711 -1446
rect 715 -1452 718 -1446
rect 722 -1452 725 -1446
rect 729 -1452 732 -1446
rect 736 -1452 739 -1446
rect 743 -1452 746 -1446
rect 750 -1452 753 -1446
rect 764 -1452 770 -1446
rect 771 -1452 774 -1446
rect 778 -1452 784 -1446
rect 785 -1452 791 -1446
rect 792 -1452 798 -1446
rect 799 -1452 805 -1446
rect 806 -1452 809 -1446
rect 813 -1452 819 -1446
rect 827 -1452 830 -1446
rect 834 -1452 837 -1446
rect 1 -1531 7 -1525
rect 8 -1531 11 -1525
rect 15 -1531 18 -1525
rect 22 -1531 25 -1525
rect 29 -1531 32 -1525
rect 36 -1531 39 -1525
rect 43 -1531 46 -1525
rect 50 -1531 56 -1525
rect 57 -1531 60 -1525
rect 64 -1531 67 -1525
rect 71 -1531 77 -1525
rect 78 -1531 81 -1525
rect 85 -1531 88 -1525
rect 92 -1531 98 -1525
rect 99 -1531 102 -1525
rect 106 -1531 109 -1525
rect 113 -1531 116 -1525
rect 120 -1531 123 -1525
rect 127 -1531 130 -1525
rect 134 -1531 140 -1525
rect 141 -1531 144 -1525
rect 148 -1531 151 -1525
rect 155 -1531 158 -1525
rect 162 -1531 168 -1525
rect 169 -1531 175 -1525
rect 176 -1531 182 -1525
rect 183 -1531 189 -1525
rect 190 -1531 193 -1525
rect 197 -1531 200 -1525
rect 204 -1531 210 -1525
rect 211 -1531 214 -1525
rect 218 -1531 221 -1525
rect 225 -1531 228 -1525
rect 232 -1531 238 -1525
rect 239 -1531 245 -1525
rect 246 -1531 252 -1525
rect 253 -1531 259 -1525
rect 260 -1531 263 -1525
rect 267 -1531 273 -1525
rect 274 -1531 277 -1525
rect 281 -1531 284 -1525
rect 288 -1531 291 -1525
rect 295 -1531 298 -1525
rect 302 -1531 308 -1525
rect 309 -1531 312 -1525
rect 316 -1531 319 -1525
rect 323 -1531 326 -1525
rect 330 -1531 336 -1525
rect 337 -1531 343 -1525
rect 344 -1531 347 -1525
rect 351 -1531 354 -1525
rect 358 -1531 364 -1525
rect 365 -1531 371 -1525
rect 372 -1531 375 -1525
rect 379 -1531 385 -1525
rect 386 -1531 392 -1525
rect 393 -1531 396 -1525
rect 400 -1531 403 -1525
rect 407 -1531 410 -1525
rect 414 -1531 420 -1525
rect 421 -1531 424 -1525
rect 428 -1531 431 -1525
rect 435 -1531 441 -1525
rect 442 -1531 445 -1525
rect 449 -1531 452 -1525
rect 456 -1531 459 -1525
rect 463 -1531 466 -1525
rect 470 -1531 473 -1525
rect 477 -1531 480 -1525
rect 484 -1531 487 -1525
rect 491 -1531 494 -1525
rect 498 -1531 501 -1525
rect 505 -1531 508 -1525
rect 512 -1531 515 -1525
rect 519 -1531 525 -1525
rect 526 -1531 529 -1525
rect 533 -1531 536 -1525
rect 540 -1531 543 -1525
rect 547 -1531 550 -1525
rect 554 -1531 557 -1525
rect 561 -1531 564 -1525
rect 568 -1531 571 -1525
rect 575 -1531 578 -1525
rect 582 -1531 585 -1525
rect 589 -1531 592 -1525
rect 596 -1531 602 -1525
rect 603 -1531 606 -1525
rect 610 -1531 613 -1525
rect 617 -1531 623 -1525
rect 624 -1531 627 -1525
rect 631 -1531 634 -1525
rect 638 -1531 641 -1525
rect 645 -1531 648 -1525
rect 652 -1531 655 -1525
rect 659 -1531 662 -1525
rect 666 -1531 669 -1525
rect 673 -1531 676 -1525
rect 680 -1531 683 -1525
rect 687 -1531 690 -1525
rect 694 -1531 697 -1525
rect 701 -1531 704 -1525
rect 708 -1531 711 -1525
rect 715 -1531 718 -1525
rect 722 -1531 725 -1525
rect 729 -1531 732 -1525
rect 736 -1531 739 -1525
rect 743 -1531 746 -1525
rect 750 -1531 753 -1525
rect 1 -1610 7 -1604
rect 8 -1610 14 -1604
rect 15 -1610 18 -1604
rect 22 -1610 25 -1604
rect 29 -1610 35 -1604
rect 36 -1610 39 -1604
rect 43 -1610 49 -1604
rect 50 -1610 53 -1604
rect 57 -1610 60 -1604
rect 64 -1610 67 -1604
rect 71 -1610 74 -1604
rect 78 -1610 84 -1604
rect 85 -1610 91 -1604
rect 92 -1610 95 -1604
rect 99 -1610 105 -1604
rect 106 -1610 109 -1604
rect 113 -1610 119 -1604
rect 120 -1610 123 -1604
rect 127 -1610 130 -1604
rect 134 -1610 140 -1604
rect 141 -1610 147 -1604
rect 148 -1610 154 -1604
rect 155 -1610 158 -1604
rect 162 -1610 165 -1604
rect 169 -1610 172 -1604
rect 176 -1610 179 -1604
rect 183 -1610 186 -1604
rect 190 -1610 196 -1604
rect 197 -1610 200 -1604
rect 204 -1610 207 -1604
rect 211 -1610 214 -1604
rect 218 -1610 224 -1604
rect 225 -1610 228 -1604
rect 232 -1610 238 -1604
rect 239 -1610 242 -1604
rect 246 -1610 249 -1604
rect 253 -1610 256 -1604
rect 260 -1610 263 -1604
rect 267 -1610 270 -1604
rect 274 -1610 280 -1604
rect 281 -1610 284 -1604
rect 288 -1610 291 -1604
rect 295 -1610 298 -1604
rect 302 -1610 308 -1604
rect 309 -1610 315 -1604
rect 316 -1610 322 -1604
rect 323 -1610 326 -1604
rect 330 -1610 333 -1604
rect 337 -1610 343 -1604
rect 344 -1610 347 -1604
rect 351 -1610 354 -1604
rect 358 -1610 364 -1604
rect 365 -1610 371 -1604
rect 372 -1610 375 -1604
rect 379 -1610 382 -1604
rect 386 -1610 389 -1604
rect 393 -1610 396 -1604
rect 400 -1610 403 -1604
rect 407 -1610 413 -1604
rect 414 -1610 417 -1604
rect 421 -1610 424 -1604
rect 428 -1610 431 -1604
rect 435 -1610 441 -1604
rect 442 -1610 448 -1604
rect 449 -1610 452 -1604
rect 456 -1610 459 -1604
rect 463 -1610 466 -1604
rect 470 -1610 476 -1604
rect 477 -1610 480 -1604
rect 484 -1610 490 -1604
rect 491 -1610 494 -1604
rect 498 -1610 501 -1604
rect 505 -1610 508 -1604
rect 512 -1610 515 -1604
rect 519 -1610 522 -1604
rect 526 -1610 529 -1604
rect 533 -1610 536 -1604
rect 540 -1610 543 -1604
rect 547 -1610 550 -1604
rect 554 -1610 560 -1604
rect 561 -1610 564 -1604
rect 568 -1610 571 -1604
rect 575 -1610 578 -1604
rect 582 -1610 585 -1604
rect 589 -1610 592 -1604
rect 596 -1610 599 -1604
rect 603 -1610 606 -1604
rect 610 -1610 613 -1604
rect 617 -1610 620 -1604
rect 624 -1610 627 -1604
rect 631 -1610 634 -1604
rect 638 -1610 641 -1604
rect 645 -1610 648 -1604
rect 652 -1610 655 -1604
rect 659 -1610 662 -1604
rect 666 -1610 669 -1604
rect 673 -1610 676 -1604
rect 680 -1610 683 -1604
rect 8 -1679 11 -1673
rect 15 -1679 18 -1673
rect 22 -1679 25 -1673
rect 29 -1679 35 -1673
rect 36 -1679 39 -1673
rect 43 -1679 49 -1673
rect 50 -1679 56 -1673
rect 57 -1679 60 -1673
rect 64 -1679 67 -1673
rect 71 -1679 74 -1673
rect 78 -1679 81 -1673
rect 85 -1679 91 -1673
rect 92 -1679 95 -1673
rect 99 -1679 105 -1673
rect 106 -1679 112 -1673
rect 113 -1679 119 -1673
rect 120 -1679 123 -1673
rect 127 -1679 130 -1673
rect 134 -1679 137 -1673
rect 141 -1679 147 -1673
rect 148 -1679 151 -1673
rect 155 -1679 158 -1673
rect 162 -1679 165 -1673
rect 169 -1679 175 -1673
rect 176 -1679 179 -1673
rect 183 -1679 189 -1673
rect 190 -1679 196 -1673
rect 197 -1679 200 -1673
rect 204 -1679 207 -1673
rect 211 -1679 214 -1673
rect 218 -1679 221 -1673
rect 225 -1679 228 -1673
rect 232 -1679 238 -1673
rect 239 -1679 245 -1673
rect 246 -1679 249 -1673
rect 253 -1679 256 -1673
rect 260 -1679 266 -1673
rect 267 -1679 270 -1673
rect 274 -1679 277 -1673
rect 281 -1679 284 -1673
rect 288 -1679 294 -1673
rect 295 -1679 301 -1673
rect 302 -1679 308 -1673
rect 309 -1679 312 -1673
rect 316 -1679 319 -1673
rect 323 -1679 326 -1673
rect 330 -1679 336 -1673
rect 337 -1679 343 -1673
rect 344 -1679 347 -1673
rect 351 -1679 357 -1673
rect 358 -1679 364 -1673
rect 365 -1679 371 -1673
rect 372 -1679 378 -1673
rect 379 -1679 382 -1673
rect 386 -1679 392 -1673
rect 393 -1679 396 -1673
rect 400 -1679 403 -1673
rect 407 -1679 410 -1673
rect 414 -1679 417 -1673
rect 421 -1679 424 -1673
rect 428 -1679 431 -1673
rect 435 -1679 438 -1673
rect 442 -1679 445 -1673
rect 449 -1679 452 -1673
rect 456 -1679 459 -1673
rect 463 -1679 466 -1673
rect 470 -1679 473 -1673
rect 477 -1679 480 -1673
rect 484 -1679 487 -1673
rect 491 -1679 494 -1673
rect 498 -1679 501 -1673
rect 505 -1679 508 -1673
rect 512 -1679 515 -1673
rect 519 -1679 522 -1673
rect 526 -1679 529 -1673
rect 533 -1679 536 -1673
rect 540 -1679 543 -1673
rect 547 -1679 550 -1673
rect 554 -1679 557 -1673
rect 561 -1679 564 -1673
rect 568 -1679 571 -1673
rect 575 -1679 578 -1673
rect 582 -1679 585 -1673
rect 589 -1679 592 -1673
rect 596 -1679 599 -1673
rect 610 -1679 613 -1673
rect 617 -1679 623 -1673
rect 645 -1679 651 -1673
rect 659 -1679 662 -1673
rect 673 -1679 679 -1673
rect 680 -1679 683 -1673
rect 8 -1736 11 -1730
rect 15 -1736 18 -1730
rect 22 -1736 25 -1730
rect 29 -1736 35 -1730
rect 36 -1736 42 -1730
rect 43 -1736 46 -1730
rect 50 -1736 53 -1730
rect 57 -1736 60 -1730
rect 64 -1736 67 -1730
rect 71 -1736 74 -1730
rect 78 -1736 81 -1730
rect 85 -1736 88 -1730
rect 92 -1736 98 -1730
rect 99 -1736 105 -1730
rect 106 -1736 109 -1730
rect 113 -1736 116 -1730
rect 120 -1736 126 -1730
rect 127 -1736 133 -1730
rect 134 -1736 137 -1730
rect 141 -1736 147 -1730
rect 148 -1736 154 -1730
rect 155 -1736 161 -1730
rect 162 -1736 165 -1730
rect 169 -1736 172 -1730
rect 176 -1736 182 -1730
rect 183 -1736 189 -1730
rect 190 -1736 193 -1730
rect 197 -1736 200 -1730
rect 204 -1736 210 -1730
rect 211 -1736 214 -1730
rect 218 -1736 221 -1730
rect 225 -1736 228 -1730
rect 232 -1736 235 -1730
rect 239 -1736 245 -1730
rect 246 -1736 252 -1730
rect 253 -1736 259 -1730
rect 260 -1736 263 -1730
rect 267 -1736 273 -1730
rect 274 -1736 277 -1730
rect 281 -1736 284 -1730
rect 288 -1736 294 -1730
rect 295 -1736 298 -1730
rect 302 -1736 305 -1730
rect 309 -1736 315 -1730
rect 316 -1736 322 -1730
rect 323 -1736 326 -1730
rect 330 -1736 333 -1730
rect 337 -1736 343 -1730
rect 344 -1736 347 -1730
rect 351 -1736 357 -1730
rect 358 -1736 364 -1730
rect 365 -1736 368 -1730
rect 372 -1736 378 -1730
rect 379 -1736 382 -1730
rect 393 -1736 396 -1730
rect 400 -1736 403 -1730
rect 407 -1736 410 -1730
rect 414 -1736 417 -1730
rect 421 -1736 424 -1730
rect 428 -1736 431 -1730
rect 435 -1736 438 -1730
rect 442 -1736 448 -1730
rect 456 -1736 462 -1730
rect 463 -1736 466 -1730
rect 470 -1736 473 -1730
rect 477 -1736 480 -1730
rect 484 -1736 487 -1730
rect 491 -1736 494 -1730
rect 498 -1736 501 -1730
rect 519 -1736 522 -1730
rect 526 -1736 529 -1730
rect 554 -1736 557 -1730
rect 575 -1736 581 -1730
rect 617 -1736 620 -1730
rect 652 -1736 655 -1730
rect 666 -1736 672 -1730
rect 673 -1736 676 -1730
rect 36 -1777 39 -1771
rect 50 -1777 53 -1771
rect 57 -1777 63 -1771
rect 64 -1777 67 -1771
rect 71 -1777 74 -1771
rect 85 -1777 88 -1771
rect 92 -1777 95 -1771
rect 99 -1777 105 -1771
rect 106 -1777 112 -1771
rect 113 -1777 119 -1771
rect 120 -1777 126 -1771
rect 127 -1777 130 -1771
rect 134 -1777 137 -1771
rect 141 -1777 144 -1771
rect 148 -1777 154 -1771
rect 155 -1777 161 -1771
rect 162 -1777 168 -1771
rect 169 -1777 175 -1771
rect 176 -1777 182 -1771
rect 183 -1777 189 -1771
rect 190 -1777 193 -1771
rect 197 -1777 200 -1771
rect 204 -1777 210 -1771
rect 211 -1777 217 -1771
rect 218 -1777 221 -1771
rect 225 -1777 228 -1771
rect 232 -1777 235 -1771
rect 239 -1777 242 -1771
rect 253 -1777 259 -1771
rect 260 -1777 263 -1771
rect 267 -1777 270 -1771
rect 274 -1777 280 -1771
rect 288 -1777 291 -1771
rect 295 -1777 298 -1771
rect 309 -1777 312 -1771
rect 316 -1777 319 -1771
rect 323 -1777 326 -1771
rect 330 -1777 336 -1771
rect 337 -1777 340 -1771
rect 344 -1777 347 -1771
rect 351 -1777 354 -1771
rect 365 -1777 368 -1771
rect 379 -1777 385 -1771
rect 400 -1777 406 -1771
rect 414 -1777 420 -1771
rect 421 -1777 424 -1771
rect 428 -1777 431 -1771
rect 449 -1777 455 -1771
rect 456 -1777 462 -1771
rect 463 -1777 466 -1771
rect 470 -1777 473 -1771
rect 477 -1777 480 -1771
rect 484 -1777 490 -1771
rect 498 -1777 504 -1771
rect 512 -1777 515 -1771
rect 519 -1777 522 -1771
rect 526 -1777 529 -1771
rect 533 -1777 536 -1771
rect 540 -1777 546 -1771
rect 547 -1777 550 -1771
rect 561 -1777 567 -1771
rect 610 -1777 616 -1771
rect 617 -1777 620 -1771
rect 631 -1777 634 -1771
rect 50 -1806 53 -1800
rect 57 -1806 63 -1800
rect 85 -1806 91 -1800
rect 99 -1806 105 -1800
rect 106 -1806 112 -1800
rect 113 -1806 119 -1800
rect 120 -1806 126 -1800
rect 127 -1806 133 -1800
rect 134 -1806 140 -1800
rect 141 -1806 147 -1800
rect 148 -1806 151 -1800
rect 155 -1806 158 -1800
rect 169 -1806 175 -1800
rect 176 -1806 182 -1800
rect 183 -1806 189 -1800
rect 204 -1806 207 -1800
rect 232 -1806 235 -1800
rect 246 -1806 252 -1800
rect 253 -1806 259 -1800
rect 260 -1806 266 -1800
rect 267 -1806 273 -1800
rect 309 -1806 315 -1800
rect 351 -1806 354 -1800
rect 372 -1806 378 -1800
rect 386 -1806 392 -1800
rect 407 -1806 413 -1800
rect 414 -1806 420 -1800
rect 463 -1806 469 -1800
rect 470 -1806 473 -1800
rect 477 -1806 483 -1800
rect 498 -1806 504 -1800
rect 519 -1806 522 -1800
rect 526 -1806 532 -1800
rect 638 -1806 644 -1800
<< polysilicon >>
rect 47 -15 48 -13
rect 58 -9 59 -7
rect 93 -9 94 -7
rect 93 -15 94 -13
rect 114 -9 115 -7
rect 114 -15 115 -13
rect 124 -9 125 -7
rect 128 -9 129 -7
rect 128 -15 129 -13
rect 135 -9 136 -7
rect 142 -9 143 -7
rect 152 -9 153 -7
rect 156 -9 157 -7
rect 163 -9 164 -7
rect 163 -15 164 -13
rect 170 -9 171 -7
rect 170 -15 171 -13
rect 177 -9 178 -7
rect 177 -15 178 -13
rect 184 -9 185 -7
rect 184 -15 185 -13
rect 191 -9 192 -7
rect 198 -9 199 -7
rect 198 -15 199 -13
rect 205 -9 206 -7
rect 205 -15 206 -13
rect 212 -9 213 -7
rect 212 -15 213 -13
rect 222 -15 223 -13
rect 226 -15 227 -13
rect 236 -9 237 -7
rect 233 -15 234 -13
rect 240 -9 241 -7
rect 240 -15 241 -13
rect 257 -9 258 -7
rect 261 -9 262 -7
rect 261 -15 262 -13
rect 289 -15 290 -13
rect 338 -9 339 -7
rect 338 -15 339 -13
rect 44 -36 45 -34
rect 51 -42 52 -40
rect 72 -36 73 -34
rect 72 -42 73 -40
rect 79 -36 80 -34
rect 93 -36 94 -34
rect 93 -42 94 -40
rect 103 -36 104 -34
rect 107 -42 108 -40
rect 117 -42 118 -40
rect 124 -36 125 -34
rect 128 -36 129 -34
rect 131 -36 132 -34
rect 135 -36 136 -34
rect 135 -42 136 -40
rect 142 -36 143 -34
rect 149 -36 150 -34
rect 156 -42 157 -40
rect 163 -36 164 -34
rect 170 -36 171 -34
rect 170 -42 171 -40
rect 177 -36 178 -34
rect 177 -42 178 -40
rect 184 -36 185 -34
rect 184 -42 185 -40
rect 191 -36 192 -34
rect 191 -42 192 -40
rect 198 -36 199 -34
rect 198 -42 199 -40
rect 205 -36 206 -34
rect 205 -42 206 -40
rect 208 -42 209 -40
rect 212 -36 213 -34
rect 212 -42 213 -40
rect 219 -36 220 -34
rect 219 -42 220 -40
rect 226 -36 227 -34
rect 226 -42 227 -40
rect 233 -36 234 -34
rect 233 -42 234 -40
rect 240 -36 241 -34
rect 240 -42 241 -40
rect 247 -36 248 -34
rect 247 -42 248 -40
rect 254 -36 255 -34
rect 254 -42 255 -40
rect 271 -36 272 -34
rect 271 -42 272 -40
rect 275 -36 276 -34
rect 275 -42 276 -40
rect 282 -36 283 -34
rect 285 -36 286 -34
rect 292 -42 293 -40
rect 296 -36 297 -34
rect 296 -42 297 -40
rect 313 -36 314 -34
rect 317 -36 318 -34
rect 317 -42 318 -40
rect 324 -36 325 -34
rect 324 -42 325 -40
rect 334 -36 335 -34
rect 338 -36 339 -34
rect 338 -42 339 -40
rect 345 -36 346 -34
rect 345 -42 346 -40
rect 352 -36 353 -34
rect 352 -42 353 -40
rect 387 -36 388 -34
rect 387 -42 388 -40
rect 404 -42 405 -40
rect 16 -71 17 -69
rect 16 -77 17 -75
rect 23 -71 24 -69
rect 23 -77 24 -75
rect 37 -77 38 -75
rect 44 -71 45 -69
rect 44 -77 45 -75
rect 58 -71 59 -69
rect 61 -71 62 -69
rect 65 -71 66 -69
rect 65 -77 66 -75
rect 72 -77 73 -75
rect 82 -71 83 -69
rect 86 -71 87 -69
rect 93 -71 94 -69
rect 93 -77 94 -75
rect 100 -71 101 -69
rect 100 -77 101 -75
rect 110 -71 111 -69
rect 114 -71 115 -69
rect 121 -71 122 -69
rect 121 -77 122 -75
rect 128 -71 129 -69
rect 128 -77 129 -75
rect 135 -71 136 -69
rect 135 -77 136 -75
rect 142 -71 143 -69
rect 142 -77 143 -75
rect 152 -71 153 -69
rect 149 -77 150 -75
rect 152 -77 153 -75
rect 156 -71 157 -69
rect 156 -77 157 -75
rect 163 -71 164 -69
rect 163 -77 164 -75
rect 170 -71 171 -69
rect 170 -77 171 -75
rect 177 -71 178 -69
rect 180 -71 181 -69
rect 184 -71 185 -69
rect 184 -77 185 -75
rect 187 -77 188 -75
rect 194 -71 195 -69
rect 194 -77 195 -75
rect 198 -71 199 -69
rect 198 -77 199 -75
rect 205 -71 206 -69
rect 205 -77 206 -75
rect 208 -77 209 -75
rect 212 -71 213 -69
rect 212 -77 213 -75
rect 222 -71 223 -69
rect 222 -77 223 -75
rect 226 -71 227 -69
rect 226 -77 227 -75
rect 233 -71 234 -69
rect 233 -77 234 -75
rect 240 -71 241 -69
rect 240 -77 241 -75
rect 247 -77 248 -75
rect 250 -77 251 -75
rect 254 -71 255 -69
rect 254 -77 255 -75
rect 261 -71 262 -69
rect 261 -77 262 -75
rect 268 -71 269 -69
rect 271 -71 272 -69
rect 275 -71 276 -69
rect 275 -77 276 -75
rect 282 -71 283 -69
rect 289 -71 290 -69
rect 289 -77 290 -75
rect 299 -71 300 -69
rect 299 -77 300 -75
rect 303 -77 304 -75
rect 306 -77 307 -75
rect 310 -71 311 -69
rect 310 -77 311 -75
rect 317 -71 318 -69
rect 317 -77 318 -75
rect 324 -71 325 -69
rect 324 -77 325 -75
rect 331 -71 332 -69
rect 331 -77 332 -75
rect 341 -71 342 -69
rect 345 -71 346 -69
rect 345 -77 346 -75
rect 359 -71 360 -69
rect 359 -77 360 -75
rect 366 -71 367 -69
rect 366 -77 367 -75
rect 373 -71 374 -69
rect 373 -77 374 -75
rect 380 -71 381 -69
rect 380 -77 381 -75
rect 387 -71 388 -69
rect 387 -77 388 -75
rect 394 -71 395 -69
rect 397 -77 398 -75
rect 401 -71 402 -69
rect 401 -77 402 -75
rect 408 -71 409 -69
rect 408 -77 409 -75
rect 415 -71 416 -69
rect 415 -77 416 -75
rect 422 -71 423 -69
rect 422 -77 423 -75
rect 436 -71 437 -69
rect 436 -77 437 -75
rect 44 -130 45 -128
rect 51 -130 52 -128
rect 58 -124 59 -122
rect 58 -130 59 -128
rect 65 -130 66 -128
rect 75 -130 76 -128
rect 79 -124 80 -122
rect 79 -130 80 -128
rect 86 -124 87 -122
rect 86 -130 87 -128
rect 93 -124 94 -122
rect 93 -130 94 -128
rect 100 -130 101 -128
rect 103 -130 104 -128
rect 107 -124 108 -122
rect 107 -130 108 -128
rect 114 -124 115 -122
rect 121 -124 122 -122
rect 121 -130 122 -128
rect 128 -124 129 -122
rect 128 -130 129 -128
rect 135 -130 136 -128
rect 138 -130 139 -128
rect 142 -124 143 -122
rect 142 -130 143 -128
rect 149 -124 150 -122
rect 149 -130 150 -128
rect 156 -124 157 -122
rect 159 -130 160 -128
rect 163 -124 164 -122
rect 163 -130 164 -128
rect 173 -124 174 -122
rect 170 -130 171 -128
rect 177 -124 178 -122
rect 177 -130 178 -128
rect 180 -130 181 -128
rect 187 -124 188 -122
rect 187 -130 188 -128
rect 191 -124 192 -122
rect 191 -130 192 -128
rect 198 -124 199 -122
rect 198 -130 199 -128
rect 205 -124 206 -122
rect 205 -130 206 -128
rect 212 -124 213 -122
rect 212 -130 213 -128
rect 219 -124 220 -122
rect 219 -130 220 -128
rect 226 -124 227 -122
rect 226 -130 227 -128
rect 233 -124 234 -122
rect 233 -130 234 -128
rect 240 -130 241 -128
rect 243 -130 244 -128
rect 247 -124 248 -122
rect 247 -130 248 -128
rect 254 -124 255 -122
rect 261 -124 262 -122
rect 261 -130 262 -128
rect 268 -124 269 -122
rect 268 -130 269 -128
rect 275 -124 276 -122
rect 275 -130 276 -128
rect 282 -124 283 -122
rect 285 -124 286 -122
rect 282 -130 283 -128
rect 289 -124 290 -122
rect 292 -124 293 -122
rect 289 -130 290 -128
rect 296 -124 297 -122
rect 296 -130 297 -128
rect 303 -124 304 -122
rect 303 -130 304 -128
rect 310 -124 311 -122
rect 310 -130 311 -128
rect 317 -124 318 -122
rect 317 -130 318 -128
rect 324 -130 325 -128
rect 327 -130 328 -128
rect 331 -124 332 -122
rect 334 -124 335 -122
rect 334 -130 335 -128
rect 338 -124 339 -122
rect 345 -124 346 -122
rect 345 -130 346 -128
rect 352 -130 353 -128
rect 359 -124 360 -122
rect 359 -130 360 -128
rect 366 -124 367 -122
rect 366 -130 367 -128
rect 373 -124 374 -122
rect 373 -130 374 -128
rect 380 -124 381 -122
rect 383 -130 384 -128
rect 387 -124 388 -122
rect 387 -130 388 -128
rect 394 -124 395 -122
rect 394 -130 395 -128
rect 401 -124 402 -122
rect 401 -130 402 -128
rect 408 -124 409 -122
rect 408 -130 409 -128
rect 415 -124 416 -122
rect 415 -130 416 -128
rect 422 -124 423 -122
rect 422 -130 423 -128
rect 429 -124 430 -122
rect 429 -130 430 -128
rect 436 -124 437 -122
rect 436 -130 437 -128
rect 443 -124 444 -122
rect 443 -130 444 -128
rect 450 -124 451 -122
rect 450 -130 451 -128
rect 457 -124 458 -122
rect 457 -130 458 -128
rect 464 -124 465 -122
rect 464 -130 465 -128
rect 471 -124 472 -122
rect 471 -130 472 -128
rect 478 -124 479 -122
rect 478 -130 479 -128
rect 485 -124 486 -122
rect 485 -130 486 -128
rect 492 -124 493 -122
rect 492 -130 493 -128
rect 499 -124 500 -122
rect 499 -130 500 -128
rect 506 -124 507 -122
rect 506 -130 507 -128
rect 513 -124 514 -122
rect 513 -130 514 -128
rect 520 -124 521 -122
rect 520 -130 521 -128
rect 12 -199 13 -197
rect 16 -205 17 -203
rect 23 -205 24 -203
rect 30 -205 31 -203
rect 33 -205 34 -203
rect 44 -199 45 -197
rect 44 -205 45 -203
rect 58 -199 59 -197
rect 58 -205 59 -203
rect 65 -199 66 -197
rect 65 -205 66 -203
rect 72 -199 73 -197
rect 72 -205 73 -203
rect 79 -199 80 -197
rect 79 -205 80 -203
rect 89 -199 90 -197
rect 89 -205 90 -203
rect 93 -199 94 -197
rect 93 -205 94 -203
rect 100 -199 101 -197
rect 100 -205 101 -203
rect 107 -199 108 -197
rect 107 -205 108 -203
rect 117 -199 118 -197
rect 114 -205 115 -203
rect 121 -199 122 -197
rect 121 -205 122 -203
rect 128 -199 129 -197
rect 128 -205 129 -203
rect 135 -199 136 -197
rect 135 -205 136 -203
rect 142 -199 143 -197
rect 142 -205 143 -203
rect 149 -199 150 -197
rect 152 -199 153 -197
rect 152 -205 153 -203
rect 156 -199 157 -197
rect 156 -205 157 -203
rect 163 -199 164 -197
rect 163 -205 164 -203
rect 170 -199 171 -197
rect 170 -205 171 -203
rect 177 -199 178 -197
rect 180 -199 181 -197
rect 180 -205 181 -203
rect 187 -199 188 -197
rect 187 -205 188 -203
rect 191 -199 192 -197
rect 191 -205 192 -203
rect 198 -199 199 -197
rect 198 -205 199 -203
rect 201 -205 202 -203
rect 208 -205 209 -203
rect 212 -205 213 -203
rect 215 -205 216 -203
rect 219 -199 220 -197
rect 219 -205 220 -203
rect 226 -199 227 -197
rect 226 -205 227 -203
rect 233 -199 234 -197
rect 233 -205 234 -203
rect 240 -199 241 -197
rect 240 -205 241 -203
rect 250 -199 251 -197
rect 247 -205 248 -203
rect 250 -205 251 -203
rect 254 -199 255 -197
rect 254 -205 255 -203
rect 257 -205 258 -203
rect 261 -199 262 -197
rect 261 -205 262 -203
rect 271 -199 272 -197
rect 268 -205 269 -203
rect 275 -199 276 -197
rect 275 -205 276 -203
rect 282 -199 283 -197
rect 285 -199 286 -197
rect 282 -205 283 -203
rect 285 -205 286 -203
rect 289 -199 290 -197
rect 292 -199 293 -197
rect 292 -205 293 -203
rect 296 -199 297 -197
rect 296 -205 297 -203
rect 303 -199 304 -197
rect 303 -205 304 -203
rect 313 -205 314 -203
rect 317 -199 318 -197
rect 317 -205 318 -203
rect 324 -199 325 -197
rect 324 -205 325 -203
rect 331 -199 332 -197
rect 331 -205 332 -203
rect 341 -199 342 -197
rect 338 -205 339 -203
rect 345 -199 346 -197
rect 345 -205 346 -203
rect 352 -199 353 -197
rect 352 -205 353 -203
rect 359 -199 360 -197
rect 359 -205 360 -203
rect 366 -199 367 -197
rect 366 -205 367 -203
rect 373 -199 374 -197
rect 373 -205 374 -203
rect 380 -199 381 -197
rect 380 -205 381 -203
rect 387 -199 388 -197
rect 390 -199 391 -197
rect 387 -205 388 -203
rect 394 -199 395 -197
rect 394 -205 395 -203
rect 401 -199 402 -197
rect 401 -205 402 -203
rect 408 -199 409 -197
rect 411 -205 412 -203
rect 415 -199 416 -197
rect 415 -205 416 -203
rect 422 -199 423 -197
rect 425 -205 426 -203
rect 429 -199 430 -197
rect 429 -205 430 -203
rect 436 -199 437 -197
rect 436 -205 437 -203
rect 443 -199 444 -197
rect 443 -205 444 -203
rect 450 -199 451 -197
rect 450 -205 451 -203
rect 457 -199 458 -197
rect 457 -205 458 -203
rect 464 -199 465 -197
rect 464 -205 465 -203
rect 471 -199 472 -197
rect 471 -205 472 -203
rect 478 -199 479 -197
rect 478 -205 479 -203
rect 485 -199 486 -197
rect 485 -205 486 -203
rect 492 -199 493 -197
rect 492 -205 493 -203
rect 499 -199 500 -197
rect 499 -205 500 -203
rect 506 -199 507 -197
rect 506 -205 507 -203
rect 513 -199 514 -197
rect 513 -205 514 -203
rect 520 -199 521 -197
rect 520 -205 521 -203
rect 527 -199 528 -197
rect 527 -205 528 -203
rect 534 -199 535 -197
rect 534 -205 535 -203
rect 541 -199 542 -197
rect 541 -205 542 -203
rect 548 -199 549 -197
rect 548 -205 549 -203
rect 555 -199 556 -197
rect 555 -205 556 -203
rect 562 -199 563 -197
rect 562 -205 563 -203
rect 569 -199 570 -197
rect 569 -205 570 -203
rect 576 -199 577 -197
rect 576 -205 577 -203
rect 583 -199 584 -197
rect 583 -205 584 -203
rect 590 -199 591 -197
rect 590 -205 591 -203
rect 597 -199 598 -197
rect 597 -205 598 -203
rect 604 -199 605 -197
rect 604 -205 605 -203
rect 611 -199 612 -197
rect 611 -205 612 -203
rect 618 -199 619 -197
rect 618 -205 619 -203
rect 625 -199 626 -197
rect 625 -205 626 -203
rect 632 -199 633 -197
rect 632 -205 633 -203
rect 639 -199 640 -197
rect 639 -205 640 -203
rect 646 -199 647 -197
rect 646 -205 647 -203
rect 653 -199 654 -197
rect 653 -205 654 -203
rect 660 -199 661 -197
rect 660 -205 661 -203
rect 16 -272 17 -270
rect 30 -272 31 -270
rect 30 -278 31 -276
rect 44 -278 45 -276
rect 51 -272 52 -270
rect 51 -278 52 -276
rect 58 -272 59 -270
rect 58 -278 59 -276
rect 65 -272 66 -270
rect 65 -278 66 -276
rect 72 -272 73 -270
rect 72 -278 73 -276
rect 82 -272 83 -270
rect 79 -278 80 -276
rect 89 -272 90 -270
rect 89 -278 90 -276
rect 93 -272 94 -270
rect 93 -278 94 -276
rect 100 -272 101 -270
rect 103 -272 104 -270
rect 100 -278 101 -276
rect 107 -272 108 -270
rect 107 -278 108 -276
rect 114 -272 115 -270
rect 114 -278 115 -276
rect 121 -272 122 -270
rect 124 -272 125 -270
rect 121 -278 122 -276
rect 128 -272 129 -270
rect 128 -278 129 -276
rect 135 -272 136 -270
rect 135 -278 136 -276
rect 142 -272 143 -270
rect 142 -278 143 -276
rect 149 -272 150 -270
rect 149 -278 150 -276
rect 156 -272 157 -270
rect 159 -278 160 -276
rect 163 -272 164 -270
rect 163 -278 164 -276
rect 170 -272 171 -270
rect 170 -278 171 -276
rect 177 -272 178 -270
rect 180 -272 181 -270
rect 177 -278 178 -276
rect 184 -272 185 -270
rect 184 -278 185 -276
rect 191 -272 192 -270
rect 191 -278 192 -276
rect 198 -272 199 -270
rect 198 -278 199 -276
rect 205 -272 206 -270
rect 205 -278 206 -276
rect 212 -272 213 -270
rect 212 -278 213 -276
rect 219 -272 220 -270
rect 219 -278 220 -276
rect 226 -272 227 -270
rect 226 -278 227 -276
rect 233 -272 234 -270
rect 233 -278 234 -276
rect 240 -272 241 -270
rect 243 -272 244 -270
rect 250 -278 251 -276
rect 257 -272 258 -270
rect 254 -278 255 -276
rect 261 -272 262 -270
rect 261 -278 262 -276
rect 268 -272 269 -270
rect 268 -278 269 -276
rect 278 -272 279 -270
rect 282 -272 283 -270
rect 285 -272 286 -270
rect 282 -278 283 -276
rect 285 -278 286 -276
rect 289 -272 290 -270
rect 289 -278 290 -276
rect 299 -272 300 -270
rect 296 -278 297 -276
rect 299 -278 300 -276
rect 303 -272 304 -270
rect 306 -272 307 -270
rect 303 -278 304 -276
rect 306 -278 307 -276
rect 310 -272 311 -270
rect 310 -278 311 -276
rect 320 -272 321 -270
rect 317 -278 318 -276
rect 320 -278 321 -276
rect 324 -272 325 -270
rect 324 -278 325 -276
rect 331 -272 332 -270
rect 334 -272 335 -270
rect 334 -278 335 -276
rect 338 -272 339 -270
rect 338 -278 339 -276
rect 345 -272 346 -270
rect 345 -278 346 -276
rect 352 -278 353 -276
rect 355 -278 356 -276
rect 359 -272 360 -270
rect 359 -278 360 -276
rect 366 -272 367 -270
rect 369 -278 370 -276
rect 373 -272 374 -270
rect 373 -278 374 -276
rect 380 -272 381 -270
rect 380 -278 381 -276
rect 387 -272 388 -270
rect 387 -278 388 -276
rect 394 -272 395 -270
rect 394 -278 395 -276
rect 401 -272 402 -270
rect 401 -278 402 -276
rect 408 -272 409 -270
rect 408 -278 409 -276
rect 415 -272 416 -270
rect 415 -278 416 -276
rect 422 -272 423 -270
rect 422 -278 423 -276
rect 429 -272 430 -270
rect 429 -278 430 -276
rect 436 -272 437 -270
rect 436 -278 437 -276
rect 443 -272 444 -270
rect 443 -278 444 -276
rect 450 -272 451 -270
rect 450 -278 451 -276
rect 457 -272 458 -270
rect 457 -278 458 -276
rect 464 -272 465 -270
rect 464 -278 465 -276
rect 471 -272 472 -270
rect 471 -278 472 -276
rect 478 -272 479 -270
rect 478 -278 479 -276
rect 485 -272 486 -270
rect 485 -278 486 -276
rect 492 -272 493 -270
rect 492 -278 493 -276
rect 499 -272 500 -270
rect 499 -278 500 -276
rect 506 -272 507 -270
rect 506 -278 507 -276
rect 513 -272 514 -270
rect 513 -278 514 -276
rect 520 -272 521 -270
rect 520 -278 521 -276
rect 527 -272 528 -270
rect 527 -278 528 -276
rect 534 -272 535 -270
rect 534 -278 535 -276
rect 541 -272 542 -270
rect 541 -278 542 -276
rect 548 -272 549 -270
rect 548 -278 549 -276
rect 562 -272 563 -270
rect 562 -278 563 -276
rect 569 -272 570 -270
rect 569 -278 570 -276
rect 576 -272 577 -270
rect 576 -278 577 -276
rect 583 -272 584 -270
rect 583 -278 584 -276
rect 590 -272 591 -270
rect 590 -278 591 -276
rect 597 -272 598 -270
rect 597 -278 598 -276
rect 604 -272 605 -270
rect 604 -278 605 -276
rect 611 -272 612 -270
rect 611 -278 612 -276
rect 618 -272 619 -270
rect 625 -272 626 -270
rect 625 -278 626 -276
rect 632 -272 633 -270
rect 632 -278 633 -276
rect 639 -278 640 -276
rect 667 -272 668 -270
rect 667 -278 668 -276
rect 9 -343 10 -341
rect 12 -343 13 -341
rect 16 -337 17 -335
rect 23 -337 24 -335
rect 30 -337 31 -335
rect 37 -337 38 -335
rect 37 -343 38 -341
rect 47 -337 48 -335
rect 44 -343 45 -341
rect 51 -337 52 -335
rect 54 -337 55 -335
rect 58 -337 59 -335
rect 58 -343 59 -341
rect 65 -337 66 -335
rect 68 -343 69 -341
rect 72 -337 73 -335
rect 75 -343 76 -341
rect 79 -337 80 -335
rect 82 -337 83 -335
rect 79 -343 80 -341
rect 89 -337 90 -335
rect 86 -343 87 -341
rect 89 -343 90 -341
rect 93 -337 94 -335
rect 93 -343 94 -341
rect 100 -343 101 -341
rect 107 -337 108 -335
rect 107 -343 108 -341
rect 114 -337 115 -335
rect 114 -343 115 -341
rect 121 -337 122 -335
rect 121 -343 122 -341
rect 128 -337 129 -335
rect 128 -343 129 -341
rect 135 -337 136 -335
rect 135 -343 136 -341
rect 142 -337 143 -335
rect 145 -337 146 -335
rect 142 -343 143 -341
rect 149 -337 150 -335
rect 149 -343 150 -341
rect 159 -337 160 -335
rect 156 -343 157 -341
rect 163 -343 164 -341
rect 170 -337 171 -335
rect 170 -343 171 -341
rect 177 -337 178 -335
rect 177 -343 178 -341
rect 184 -337 185 -335
rect 187 -337 188 -335
rect 191 -337 192 -335
rect 191 -343 192 -341
rect 201 -337 202 -335
rect 201 -343 202 -341
rect 205 -337 206 -335
rect 205 -343 206 -341
rect 212 -337 213 -335
rect 212 -343 213 -341
rect 219 -337 220 -335
rect 219 -343 220 -341
rect 226 -337 227 -335
rect 226 -343 227 -341
rect 233 -337 234 -335
rect 233 -343 234 -341
rect 240 -337 241 -335
rect 247 -337 248 -335
rect 247 -343 248 -341
rect 254 -337 255 -335
rect 254 -343 255 -341
rect 261 -337 262 -335
rect 261 -343 262 -341
rect 268 -337 269 -335
rect 268 -343 269 -341
rect 275 -337 276 -335
rect 275 -343 276 -341
rect 282 -337 283 -335
rect 282 -343 283 -341
rect 289 -337 290 -335
rect 289 -343 290 -341
rect 296 -337 297 -335
rect 296 -343 297 -341
rect 303 -337 304 -335
rect 303 -343 304 -341
rect 313 -337 314 -335
rect 310 -343 311 -341
rect 313 -343 314 -341
rect 317 -337 318 -335
rect 320 -337 321 -335
rect 324 -337 325 -335
rect 324 -343 325 -341
rect 327 -343 328 -341
rect 331 -337 332 -335
rect 331 -343 332 -341
rect 341 -337 342 -335
rect 341 -343 342 -341
rect 345 -337 346 -335
rect 345 -343 346 -341
rect 352 -343 353 -341
rect 355 -343 356 -341
rect 362 -337 363 -335
rect 359 -343 360 -341
rect 362 -343 363 -341
rect 366 -337 367 -335
rect 366 -343 367 -341
rect 373 -337 374 -335
rect 373 -343 374 -341
rect 380 -337 381 -335
rect 380 -343 381 -341
rect 387 -337 388 -335
rect 390 -337 391 -335
rect 390 -343 391 -341
rect 394 -337 395 -335
rect 394 -343 395 -341
rect 401 -337 402 -335
rect 401 -343 402 -341
rect 408 -337 409 -335
rect 408 -343 409 -341
rect 415 -337 416 -335
rect 415 -343 416 -341
rect 422 -337 423 -335
rect 422 -343 423 -341
rect 429 -337 430 -335
rect 429 -343 430 -341
rect 436 -337 437 -335
rect 436 -343 437 -341
rect 443 -337 444 -335
rect 443 -343 444 -341
rect 450 -337 451 -335
rect 450 -343 451 -341
rect 457 -337 458 -335
rect 457 -343 458 -341
rect 464 -337 465 -335
rect 464 -343 465 -341
rect 471 -337 472 -335
rect 471 -343 472 -341
rect 478 -337 479 -335
rect 478 -343 479 -341
rect 485 -337 486 -335
rect 485 -343 486 -341
rect 492 -343 493 -341
rect 495 -343 496 -341
rect 499 -337 500 -335
rect 499 -343 500 -341
rect 506 -337 507 -335
rect 506 -343 507 -341
rect 513 -337 514 -335
rect 513 -343 514 -341
rect 520 -337 521 -335
rect 520 -343 521 -341
rect 527 -337 528 -335
rect 527 -343 528 -341
rect 534 -337 535 -335
rect 534 -343 535 -341
rect 541 -337 542 -335
rect 541 -343 542 -341
rect 548 -337 549 -335
rect 548 -343 549 -341
rect 555 -337 556 -335
rect 555 -343 556 -341
rect 562 -337 563 -335
rect 562 -343 563 -341
rect 569 -337 570 -335
rect 569 -343 570 -341
rect 576 -337 577 -335
rect 576 -343 577 -341
rect 583 -337 584 -335
rect 583 -343 584 -341
rect 590 -337 591 -335
rect 590 -343 591 -341
rect 604 -337 605 -335
rect 604 -343 605 -341
rect 611 -337 612 -335
rect 611 -343 612 -341
rect 618 -337 619 -335
rect 618 -343 619 -341
rect 625 -337 626 -335
rect 625 -343 626 -341
rect 632 -337 633 -335
rect 632 -343 633 -341
rect 639 -337 640 -335
rect 639 -343 640 -341
rect 646 -337 647 -335
rect 646 -343 647 -341
rect 653 -337 654 -335
rect 653 -343 654 -341
rect 660 -337 661 -335
rect 660 -343 661 -341
rect 667 -337 668 -335
rect 667 -343 668 -341
rect 674 -337 675 -335
rect 674 -343 675 -341
rect 709 -337 710 -335
rect 709 -343 710 -341
rect 23 -404 24 -402
rect 23 -410 24 -408
rect 30 -404 31 -402
rect 37 -404 38 -402
rect 37 -410 38 -408
rect 44 -404 45 -402
rect 44 -410 45 -408
rect 51 -404 52 -402
rect 51 -410 52 -408
rect 58 -404 59 -402
rect 58 -410 59 -408
rect 65 -404 66 -402
rect 68 -410 69 -408
rect 72 -404 73 -402
rect 72 -410 73 -408
rect 79 -404 80 -402
rect 79 -410 80 -408
rect 86 -404 87 -402
rect 86 -410 87 -408
rect 93 -404 94 -402
rect 93 -410 94 -408
rect 96 -410 97 -408
rect 100 -404 101 -402
rect 100 -410 101 -408
rect 110 -404 111 -402
rect 110 -410 111 -408
rect 117 -404 118 -402
rect 121 -404 122 -402
rect 121 -410 122 -408
rect 124 -410 125 -408
rect 128 -404 129 -402
rect 128 -410 129 -408
rect 135 -404 136 -402
rect 135 -410 136 -408
rect 142 -404 143 -402
rect 142 -410 143 -408
rect 149 -404 150 -402
rect 149 -410 150 -408
rect 156 -404 157 -402
rect 163 -404 164 -402
rect 163 -410 164 -408
rect 170 -404 171 -402
rect 170 -410 171 -408
rect 177 -404 178 -402
rect 177 -410 178 -408
rect 187 -404 188 -402
rect 184 -410 185 -408
rect 191 -404 192 -402
rect 191 -410 192 -408
rect 198 -404 199 -402
rect 198 -410 199 -408
rect 205 -404 206 -402
rect 205 -410 206 -408
rect 212 -404 213 -402
rect 212 -410 213 -408
rect 219 -404 220 -402
rect 219 -410 220 -408
rect 226 -404 227 -402
rect 229 -410 230 -408
rect 233 -404 234 -402
rect 233 -410 234 -408
rect 243 -404 244 -402
rect 240 -410 241 -408
rect 243 -410 244 -408
rect 247 -404 248 -402
rect 247 -410 248 -408
rect 254 -404 255 -402
rect 254 -410 255 -408
rect 261 -404 262 -402
rect 261 -410 262 -408
rect 268 -404 269 -402
rect 268 -410 269 -408
rect 275 -404 276 -402
rect 275 -410 276 -408
rect 282 -404 283 -402
rect 282 -410 283 -408
rect 285 -410 286 -408
rect 289 -404 290 -402
rect 289 -410 290 -408
rect 296 -404 297 -402
rect 296 -410 297 -408
rect 303 -404 304 -402
rect 303 -410 304 -408
rect 310 -404 311 -402
rect 310 -410 311 -408
rect 317 -404 318 -402
rect 317 -410 318 -408
rect 324 -404 325 -402
rect 327 -410 328 -408
rect 334 -404 335 -402
rect 338 -404 339 -402
rect 341 -410 342 -408
rect 345 -404 346 -402
rect 345 -410 346 -408
rect 355 -404 356 -402
rect 352 -410 353 -408
rect 359 -404 360 -402
rect 359 -410 360 -408
rect 366 -404 367 -402
rect 366 -410 367 -408
rect 373 -404 374 -402
rect 373 -410 374 -408
rect 380 -404 381 -402
rect 383 -404 384 -402
rect 380 -410 381 -408
rect 383 -410 384 -408
rect 387 -404 388 -402
rect 390 -404 391 -402
rect 387 -410 388 -408
rect 390 -410 391 -408
rect 394 -404 395 -402
rect 394 -410 395 -408
rect 401 -404 402 -402
rect 401 -410 402 -408
rect 411 -404 412 -402
rect 415 -404 416 -402
rect 415 -410 416 -408
rect 422 -404 423 -402
rect 422 -410 423 -408
rect 432 -410 433 -408
rect 436 -404 437 -402
rect 436 -410 437 -408
rect 443 -404 444 -402
rect 443 -410 444 -408
rect 450 -404 451 -402
rect 450 -410 451 -408
rect 457 -404 458 -402
rect 457 -410 458 -408
rect 467 -404 468 -402
rect 464 -410 465 -408
rect 471 -404 472 -402
rect 471 -410 472 -408
rect 481 -404 482 -402
rect 478 -410 479 -408
rect 481 -410 482 -408
rect 485 -404 486 -402
rect 485 -410 486 -408
rect 492 -404 493 -402
rect 492 -410 493 -408
rect 502 -410 503 -408
rect 506 -404 507 -402
rect 506 -410 507 -408
rect 513 -404 514 -402
rect 513 -410 514 -408
rect 520 -404 521 -402
rect 520 -410 521 -408
rect 527 -404 528 -402
rect 527 -410 528 -408
rect 534 -404 535 -402
rect 534 -410 535 -408
rect 541 -404 542 -402
rect 541 -410 542 -408
rect 548 -404 549 -402
rect 548 -410 549 -408
rect 555 -404 556 -402
rect 555 -410 556 -408
rect 562 -404 563 -402
rect 562 -410 563 -408
rect 569 -404 570 -402
rect 569 -410 570 -408
rect 576 -404 577 -402
rect 576 -410 577 -408
rect 583 -404 584 -402
rect 583 -410 584 -408
rect 590 -404 591 -402
rect 590 -410 591 -408
rect 597 -404 598 -402
rect 597 -410 598 -408
rect 604 -404 605 -402
rect 604 -410 605 -408
rect 611 -404 612 -402
rect 611 -410 612 -408
rect 618 -404 619 -402
rect 618 -410 619 -408
rect 625 -404 626 -402
rect 625 -410 626 -408
rect 635 -404 636 -402
rect 639 -404 640 -402
rect 639 -410 640 -408
rect 646 -404 647 -402
rect 646 -410 647 -408
rect 653 -404 654 -402
rect 656 -410 657 -408
rect 660 -404 661 -402
rect 660 -410 661 -408
rect 667 -404 668 -402
rect 667 -410 668 -408
rect 716 -404 717 -402
rect 716 -410 717 -408
rect 9 -469 10 -467
rect 9 -475 10 -473
rect 16 -469 17 -467
rect 16 -475 17 -473
rect 26 -475 27 -473
rect 30 -469 31 -467
rect 30 -475 31 -473
rect 37 -469 38 -467
rect 37 -475 38 -473
rect 44 -469 45 -467
rect 44 -475 45 -473
rect 51 -469 52 -467
rect 51 -475 52 -473
rect 58 -469 59 -467
rect 58 -475 59 -473
rect 65 -469 66 -467
rect 68 -475 69 -473
rect 72 -469 73 -467
rect 75 -475 76 -473
rect 82 -469 83 -467
rect 79 -475 80 -473
rect 86 -469 87 -467
rect 86 -475 87 -473
rect 93 -469 94 -467
rect 93 -475 94 -473
rect 100 -469 101 -467
rect 103 -469 104 -467
rect 107 -469 108 -467
rect 107 -475 108 -473
rect 114 -469 115 -467
rect 114 -475 115 -473
rect 121 -469 122 -467
rect 121 -475 122 -473
rect 128 -469 129 -467
rect 128 -475 129 -473
rect 135 -469 136 -467
rect 135 -475 136 -473
rect 142 -475 143 -473
rect 145 -475 146 -473
rect 149 -469 150 -467
rect 149 -475 150 -473
rect 156 -469 157 -467
rect 156 -475 157 -473
rect 166 -469 167 -467
rect 163 -475 164 -473
rect 170 -469 171 -467
rect 170 -475 171 -473
rect 177 -469 178 -467
rect 180 -469 181 -467
rect 177 -475 178 -473
rect 180 -475 181 -473
rect 184 -469 185 -467
rect 187 -475 188 -473
rect 191 -469 192 -467
rect 194 -469 195 -467
rect 191 -475 192 -473
rect 198 -469 199 -467
rect 198 -475 199 -473
rect 205 -469 206 -467
rect 205 -475 206 -473
rect 212 -469 213 -467
rect 212 -475 213 -473
rect 219 -469 220 -467
rect 219 -475 220 -473
rect 226 -469 227 -467
rect 226 -475 227 -473
rect 233 -469 234 -467
rect 233 -475 234 -473
rect 240 -469 241 -467
rect 240 -475 241 -473
rect 247 -469 248 -467
rect 247 -475 248 -473
rect 254 -469 255 -467
rect 254 -475 255 -473
rect 261 -469 262 -467
rect 261 -475 262 -473
rect 268 -469 269 -467
rect 268 -475 269 -473
rect 275 -469 276 -467
rect 275 -475 276 -473
rect 282 -469 283 -467
rect 282 -475 283 -473
rect 289 -469 290 -467
rect 289 -475 290 -473
rect 296 -469 297 -467
rect 296 -475 297 -473
rect 303 -469 304 -467
rect 303 -475 304 -473
rect 313 -469 314 -467
rect 310 -475 311 -473
rect 317 -469 318 -467
rect 317 -475 318 -473
rect 324 -469 325 -467
rect 324 -475 325 -473
rect 331 -469 332 -467
rect 331 -475 332 -473
rect 338 -469 339 -467
rect 338 -475 339 -473
rect 345 -469 346 -467
rect 345 -475 346 -473
rect 352 -469 353 -467
rect 352 -475 353 -473
rect 359 -469 360 -467
rect 359 -475 360 -473
rect 366 -469 367 -467
rect 366 -475 367 -473
rect 373 -469 374 -467
rect 373 -475 374 -473
rect 380 -469 381 -467
rect 383 -475 384 -473
rect 387 -469 388 -467
rect 390 -469 391 -467
rect 387 -475 388 -473
rect 390 -475 391 -473
rect 394 -469 395 -467
rect 394 -475 395 -473
rect 401 -469 402 -467
rect 401 -475 402 -473
rect 408 -469 409 -467
rect 411 -469 412 -467
rect 408 -475 409 -473
rect 411 -475 412 -473
rect 418 -469 419 -467
rect 422 -469 423 -467
rect 425 -469 426 -467
rect 429 -475 430 -473
rect 432 -475 433 -473
rect 436 -469 437 -467
rect 439 -469 440 -467
rect 439 -475 440 -473
rect 446 -469 447 -467
rect 443 -475 444 -473
rect 446 -475 447 -473
rect 453 -469 454 -467
rect 453 -475 454 -473
rect 457 -469 458 -467
rect 457 -475 458 -473
rect 464 -469 465 -467
rect 464 -475 465 -473
rect 471 -469 472 -467
rect 471 -475 472 -473
rect 478 -469 479 -467
rect 478 -475 479 -473
rect 485 -469 486 -467
rect 485 -475 486 -473
rect 492 -469 493 -467
rect 492 -475 493 -473
rect 499 -469 500 -467
rect 499 -475 500 -473
rect 506 -469 507 -467
rect 506 -475 507 -473
rect 513 -469 514 -467
rect 513 -475 514 -473
rect 520 -469 521 -467
rect 520 -475 521 -473
rect 527 -469 528 -467
rect 527 -475 528 -473
rect 534 -469 535 -467
rect 534 -475 535 -473
rect 541 -469 542 -467
rect 541 -475 542 -473
rect 548 -469 549 -467
rect 548 -475 549 -473
rect 555 -469 556 -467
rect 555 -475 556 -473
rect 562 -469 563 -467
rect 562 -475 563 -473
rect 569 -469 570 -467
rect 569 -475 570 -473
rect 576 -469 577 -467
rect 576 -475 577 -473
rect 583 -469 584 -467
rect 583 -475 584 -473
rect 590 -469 591 -467
rect 590 -475 591 -473
rect 597 -469 598 -467
rect 597 -475 598 -473
rect 604 -469 605 -467
rect 604 -475 605 -473
rect 611 -469 612 -467
rect 611 -475 612 -473
rect 625 -469 626 -467
rect 625 -475 626 -473
rect 632 -469 633 -467
rect 632 -475 633 -473
rect 639 -469 640 -467
rect 639 -475 640 -473
rect 646 -469 647 -467
rect 646 -475 647 -473
rect 653 -469 654 -467
rect 653 -475 654 -473
rect 667 -469 668 -467
rect 667 -475 668 -473
rect 674 -469 675 -467
rect 674 -475 675 -473
rect 681 -469 682 -467
rect 681 -475 682 -473
rect 688 -469 689 -467
rect 688 -475 689 -473
rect 695 -469 696 -467
rect 695 -475 696 -473
rect 702 -469 703 -467
rect 702 -475 703 -473
rect 709 -469 710 -467
rect 716 -475 717 -473
rect 719 -475 720 -473
rect 723 -469 724 -467
rect 723 -475 724 -473
rect 730 -469 731 -467
rect 730 -475 731 -473
rect 23 -554 24 -552
rect 23 -560 24 -558
rect 40 -560 41 -558
rect 44 -554 45 -552
rect 44 -560 45 -558
rect 51 -554 52 -552
rect 51 -560 52 -558
rect 54 -560 55 -558
rect 61 -554 62 -552
rect 61 -560 62 -558
rect 65 -554 66 -552
rect 68 -554 69 -552
rect 65 -560 66 -558
rect 75 -554 76 -552
rect 72 -560 73 -558
rect 75 -560 76 -558
rect 79 -554 80 -552
rect 79 -560 80 -558
rect 86 -554 87 -552
rect 86 -560 87 -558
rect 93 -554 94 -552
rect 93 -560 94 -558
rect 103 -560 104 -558
rect 107 -554 108 -552
rect 107 -560 108 -558
rect 114 -554 115 -552
rect 114 -560 115 -558
rect 121 -554 122 -552
rect 124 -554 125 -552
rect 128 -554 129 -552
rect 128 -560 129 -558
rect 135 -554 136 -552
rect 135 -560 136 -558
rect 145 -554 146 -552
rect 142 -560 143 -558
rect 152 -554 153 -552
rect 156 -554 157 -552
rect 156 -560 157 -558
rect 163 -554 164 -552
rect 163 -560 164 -558
rect 166 -560 167 -558
rect 170 -554 171 -552
rect 170 -560 171 -558
rect 177 -560 178 -558
rect 184 -560 185 -558
rect 187 -560 188 -558
rect 191 -554 192 -552
rect 191 -560 192 -558
rect 198 -554 199 -552
rect 198 -560 199 -558
rect 205 -554 206 -552
rect 205 -560 206 -558
rect 212 -554 213 -552
rect 212 -560 213 -558
rect 215 -560 216 -558
rect 219 -554 220 -552
rect 219 -560 220 -558
rect 226 -554 227 -552
rect 226 -560 227 -558
rect 233 -554 234 -552
rect 233 -560 234 -558
rect 236 -560 237 -558
rect 240 -554 241 -552
rect 243 -554 244 -552
rect 240 -560 241 -558
rect 247 -554 248 -552
rect 247 -560 248 -558
rect 254 -554 255 -552
rect 254 -560 255 -558
rect 261 -554 262 -552
rect 261 -560 262 -558
rect 268 -554 269 -552
rect 268 -560 269 -558
rect 275 -554 276 -552
rect 275 -560 276 -558
rect 282 -554 283 -552
rect 282 -560 283 -558
rect 289 -554 290 -552
rect 289 -560 290 -558
rect 296 -554 297 -552
rect 296 -560 297 -558
rect 303 -554 304 -552
rect 303 -560 304 -558
rect 306 -560 307 -558
rect 310 -554 311 -552
rect 310 -560 311 -558
rect 317 -554 318 -552
rect 320 -554 321 -552
rect 317 -560 318 -558
rect 320 -560 321 -558
rect 324 -554 325 -552
rect 324 -560 325 -558
rect 331 -554 332 -552
rect 331 -560 332 -558
rect 338 -554 339 -552
rect 338 -560 339 -558
rect 345 -554 346 -552
rect 345 -560 346 -558
rect 352 -554 353 -552
rect 352 -560 353 -558
rect 359 -554 360 -552
rect 359 -560 360 -558
rect 369 -554 370 -552
rect 366 -560 367 -558
rect 369 -560 370 -558
rect 373 -554 374 -552
rect 373 -560 374 -558
rect 380 -560 381 -558
rect 383 -560 384 -558
rect 387 -554 388 -552
rect 387 -560 388 -558
rect 397 -554 398 -552
rect 394 -560 395 -558
rect 397 -560 398 -558
rect 401 -554 402 -552
rect 401 -560 402 -558
rect 408 -554 409 -552
rect 408 -560 409 -558
rect 415 -554 416 -552
rect 415 -560 416 -558
rect 422 -554 423 -552
rect 425 -560 426 -558
rect 432 -554 433 -552
rect 429 -560 430 -558
rect 432 -560 433 -558
rect 436 -554 437 -552
rect 436 -560 437 -558
rect 443 -554 444 -552
rect 446 -554 447 -552
rect 446 -560 447 -558
rect 450 -554 451 -552
rect 450 -560 451 -558
rect 457 -554 458 -552
rect 457 -560 458 -558
rect 464 -554 465 -552
rect 464 -560 465 -558
rect 471 -554 472 -552
rect 471 -560 472 -558
rect 478 -554 479 -552
rect 478 -560 479 -558
rect 485 -554 486 -552
rect 485 -560 486 -558
rect 492 -554 493 -552
rect 492 -560 493 -558
rect 499 -554 500 -552
rect 499 -560 500 -558
rect 506 -554 507 -552
rect 506 -560 507 -558
rect 513 -554 514 -552
rect 513 -560 514 -558
rect 520 -554 521 -552
rect 520 -560 521 -558
rect 527 -554 528 -552
rect 527 -560 528 -558
rect 534 -554 535 -552
rect 534 -560 535 -558
rect 541 -554 542 -552
rect 541 -560 542 -558
rect 548 -554 549 -552
rect 548 -560 549 -558
rect 555 -554 556 -552
rect 555 -560 556 -558
rect 562 -554 563 -552
rect 562 -560 563 -558
rect 569 -554 570 -552
rect 569 -560 570 -558
rect 576 -554 577 -552
rect 576 -560 577 -558
rect 583 -554 584 -552
rect 583 -560 584 -558
rect 590 -554 591 -552
rect 590 -560 591 -558
rect 597 -554 598 -552
rect 597 -560 598 -558
rect 604 -554 605 -552
rect 604 -560 605 -558
rect 611 -554 612 -552
rect 611 -560 612 -558
rect 618 -554 619 -552
rect 618 -560 619 -558
rect 625 -554 626 -552
rect 625 -560 626 -558
rect 632 -554 633 -552
rect 632 -560 633 -558
rect 639 -554 640 -552
rect 639 -560 640 -558
rect 646 -554 647 -552
rect 646 -560 647 -558
rect 653 -554 654 -552
rect 653 -560 654 -558
rect 660 -554 661 -552
rect 660 -560 661 -558
rect 667 -554 668 -552
rect 667 -560 668 -558
rect 674 -554 675 -552
rect 674 -560 675 -558
rect 681 -554 682 -552
rect 681 -560 682 -558
rect 688 -554 689 -552
rect 688 -560 689 -558
rect 695 -554 696 -552
rect 695 -560 696 -558
rect 702 -554 703 -552
rect 702 -560 703 -558
rect 709 -554 710 -552
rect 709 -560 710 -558
rect 716 -554 717 -552
rect 716 -560 717 -558
rect 723 -554 724 -552
rect 723 -560 724 -558
rect 730 -554 731 -552
rect 730 -560 731 -558
rect 737 -554 738 -552
rect 737 -560 738 -558
rect 744 -554 745 -552
rect 744 -560 745 -558
rect 751 -554 752 -552
rect 751 -560 752 -558
rect 779 -554 780 -552
rect 779 -560 780 -558
rect 16 -647 17 -645
rect 16 -653 17 -651
rect 23 -647 24 -645
rect 23 -653 24 -651
rect 30 -647 31 -645
rect 33 -647 34 -645
rect 40 -647 41 -645
rect 47 -647 48 -645
rect 44 -653 45 -651
rect 47 -653 48 -651
rect 51 -647 52 -645
rect 51 -653 52 -651
rect 58 -647 59 -645
rect 58 -653 59 -651
rect 65 -647 66 -645
rect 65 -653 66 -651
rect 72 -647 73 -645
rect 72 -653 73 -651
rect 79 -647 80 -645
rect 79 -653 80 -651
rect 86 -647 87 -645
rect 86 -653 87 -651
rect 93 -647 94 -645
rect 96 -647 97 -645
rect 100 -647 101 -645
rect 100 -653 101 -651
rect 107 -653 108 -651
rect 110 -653 111 -651
rect 114 -653 115 -651
rect 117 -653 118 -651
rect 124 -647 125 -645
rect 121 -653 122 -651
rect 124 -653 125 -651
rect 128 -647 129 -645
rect 131 -653 132 -651
rect 135 -647 136 -645
rect 135 -653 136 -651
rect 142 -647 143 -645
rect 142 -653 143 -651
rect 145 -653 146 -651
rect 149 -647 150 -645
rect 152 -653 153 -651
rect 156 -647 157 -645
rect 156 -653 157 -651
rect 163 -653 164 -651
rect 166 -653 167 -651
rect 170 -647 171 -645
rect 170 -653 171 -651
rect 177 -647 178 -645
rect 177 -653 178 -651
rect 184 -647 185 -645
rect 187 -647 188 -645
rect 184 -653 185 -651
rect 191 -647 192 -645
rect 191 -653 192 -651
rect 198 -647 199 -645
rect 198 -653 199 -651
rect 205 -647 206 -645
rect 205 -653 206 -651
rect 212 -647 213 -645
rect 212 -653 213 -651
rect 219 -647 220 -645
rect 219 -653 220 -651
rect 226 -647 227 -645
rect 226 -653 227 -651
rect 233 -647 234 -645
rect 233 -653 234 -651
rect 240 -647 241 -645
rect 240 -653 241 -651
rect 247 -647 248 -645
rect 247 -653 248 -651
rect 254 -647 255 -645
rect 254 -653 255 -651
rect 261 -647 262 -645
rect 261 -653 262 -651
rect 268 -647 269 -645
rect 268 -653 269 -651
rect 275 -647 276 -645
rect 278 -647 279 -645
rect 275 -653 276 -651
rect 278 -653 279 -651
rect 282 -647 283 -645
rect 282 -653 283 -651
rect 289 -647 290 -645
rect 292 -647 293 -645
rect 289 -653 290 -651
rect 292 -653 293 -651
rect 296 -647 297 -645
rect 296 -653 297 -651
rect 303 -647 304 -645
rect 303 -653 304 -651
rect 310 -647 311 -645
rect 310 -653 311 -651
rect 317 -647 318 -645
rect 317 -653 318 -651
rect 324 -647 325 -645
rect 324 -653 325 -651
rect 331 -647 332 -645
rect 331 -653 332 -651
rect 338 -647 339 -645
rect 338 -653 339 -651
rect 345 -647 346 -645
rect 348 -647 349 -645
rect 348 -653 349 -651
rect 352 -647 353 -645
rect 355 -647 356 -645
rect 352 -653 353 -651
rect 359 -647 360 -645
rect 359 -653 360 -651
rect 366 -647 367 -645
rect 369 -647 370 -645
rect 366 -653 367 -651
rect 369 -653 370 -651
rect 373 -647 374 -645
rect 373 -653 374 -651
rect 380 -647 381 -645
rect 380 -653 381 -651
rect 387 -647 388 -645
rect 390 -647 391 -645
rect 390 -653 391 -651
rect 394 -647 395 -645
rect 394 -653 395 -651
rect 401 -647 402 -645
rect 401 -653 402 -651
rect 411 -647 412 -645
rect 408 -653 409 -651
rect 411 -653 412 -651
rect 415 -647 416 -645
rect 418 -647 419 -645
rect 418 -653 419 -651
rect 425 -647 426 -645
rect 422 -653 423 -651
rect 429 -647 430 -645
rect 429 -653 430 -651
rect 436 -647 437 -645
rect 436 -653 437 -651
rect 443 -647 444 -645
rect 446 -647 447 -645
rect 443 -653 444 -651
rect 446 -653 447 -651
rect 450 -647 451 -645
rect 450 -653 451 -651
rect 457 -647 458 -645
rect 457 -653 458 -651
rect 464 -647 465 -645
rect 464 -653 465 -651
rect 471 -647 472 -645
rect 471 -653 472 -651
rect 478 -647 479 -645
rect 478 -653 479 -651
rect 485 -647 486 -645
rect 485 -653 486 -651
rect 499 -647 500 -645
rect 499 -653 500 -651
rect 506 -647 507 -645
rect 506 -653 507 -651
rect 513 -647 514 -645
rect 516 -647 517 -645
rect 520 -647 521 -645
rect 520 -653 521 -651
rect 527 -647 528 -645
rect 527 -653 528 -651
rect 534 -647 535 -645
rect 534 -653 535 -651
rect 541 -647 542 -645
rect 541 -653 542 -651
rect 548 -647 549 -645
rect 548 -653 549 -651
rect 555 -647 556 -645
rect 555 -653 556 -651
rect 562 -647 563 -645
rect 562 -653 563 -651
rect 569 -647 570 -645
rect 569 -653 570 -651
rect 576 -647 577 -645
rect 576 -653 577 -651
rect 583 -647 584 -645
rect 583 -653 584 -651
rect 590 -647 591 -645
rect 590 -653 591 -651
rect 597 -647 598 -645
rect 597 -653 598 -651
rect 604 -647 605 -645
rect 604 -653 605 -651
rect 611 -647 612 -645
rect 611 -653 612 -651
rect 618 -647 619 -645
rect 618 -653 619 -651
rect 625 -647 626 -645
rect 625 -653 626 -651
rect 632 -647 633 -645
rect 632 -653 633 -651
rect 639 -647 640 -645
rect 639 -653 640 -651
rect 646 -647 647 -645
rect 646 -653 647 -651
rect 653 -647 654 -645
rect 653 -653 654 -651
rect 660 -647 661 -645
rect 667 -647 668 -645
rect 667 -653 668 -651
rect 674 -647 675 -645
rect 674 -653 675 -651
rect 681 -647 682 -645
rect 681 -653 682 -651
rect 688 -647 689 -645
rect 688 -653 689 -651
rect 695 -647 696 -645
rect 695 -653 696 -651
rect 702 -647 703 -645
rect 702 -653 703 -651
rect 709 -647 710 -645
rect 709 -653 710 -651
rect 716 -647 717 -645
rect 716 -653 717 -651
rect 723 -647 724 -645
rect 723 -653 724 -651
rect 730 -647 731 -645
rect 730 -653 731 -651
rect 737 -647 738 -645
rect 737 -653 738 -651
rect 807 -647 808 -645
rect 807 -653 808 -651
rect 9 -728 10 -726
rect 9 -734 10 -732
rect 16 -728 17 -726
rect 16 -734 17 -732
rect 23 -728 24 -726
rect 23 -734 24 -732
rect 30 -728 31 -726
rect 30 -734 31 -732
rect 37 -728 38 -726
rect 37 -734 38 -732
rect 44 -728 45 -726
rect 44 -734 45 -732
rect 51 -734 52 -732
rect 58 -728 59 -726
rect 58 -734 59 -732
rect 65 -728 66 -726
rect 65 -734 66 -732
rect 68 -734 69 -732
rect 72 -734 73 -732
rect 75 -734 76 -732
rect 79 -728 80 -726
rect 79 -734 80 -732
rect 86 -728 87 -726
rect 86 -734 87 -732
rect 93 -728 94 -726
rect 96 -728 97 -726
rect 93 -734 94 -732
rect 100 -728 101 -726
rect 100 -734 101 -732
rect 107 -728 108 -726
rect 107 -734 108 -732
rect 114 -728 115 -726
rect 117 -728 118 -726
rect 117 -734 118 -732
rect 121 -728 122 -726
rect 124 -728 125 -726
rect 124 -734 125 -732
rect 128 -728 129 -726
rect 128 -734 129 -732
rect 135 -728 136 -726
rect 135 -734 136 -732
rect 142 -728 143 -726
rect 142 -734 143 -732
rect 149 -728 150 -726
rect 149 -734 150 -732
rect 156 -728 157 -726
rect 156 -734 157 -732
rect 159 -734 160 -732
rect 163 -728 164 -726
rect 166 -728 167 -726
rect 173 -728 174 -726
rect 177 -728 178 -726
rect 177 -734 178 -732
rect 184 -728 185 -726
rect 184 -734 185 -732
rect 191 -728 192 -726
rect 191 -734 192 -732
rect 198 -728 199 -726
rect 198 -734 199 -732
rect 205 -728 206 -726
rect 205 -734 206 -732
rect 212 -728 213 -726
rect 212 -734 213 -732
rect 219 -728 220 -726
rect 219 -734 220 -732
rect 226 -728 227 -726
rect 226 -734 227 -732
rect 233 -728 234 -726
rect 236 -728 237 -726
rect 233 -734 234 -732
rect 236 -734 237 -732
rect 240 -728 241 -726
rect 243 -728 244 -726
rect 240 -734 241 -732
rect 247 -728 248 -726
rect 247 -734 248 -732
rect 254 -728 255 -726
rect 257 -728 258 -726
rect 261 -728 262 -726
rect 261 -734 262 -732
rect 268 -728 269 -726
rect 268 -734 269 -732
rect 275 -728 276 -726
rect 275 -734 276 -732
rect 282 -728 283 -726
rect 282 -734 283 -732
rect 289 -728 290 -726
rect 289 -734 290 -732
rect 292 -734 293 -732
rect 296 -728 297 -726
rect 296 -734 297 -732
rect 303 -728 304 -726
rect 303 -734 304 -732
rect 310 -728 311 -726
rect 310 -734 311 -732
rect 317 -728 318 -726
rect 317 -734 318 -732
rect 324 -728 325 -726
rect 324 -734 325 -732
rect 331 -728 332 -726
rect 334 -728 335 -726
rect 331 -734 332 -732
rect 338 -728 339 -726
rect 338 -734 339 -732
rect 345 -728 346 -726
rect 345 -734 346 -732
rect 352 -728 353 -726
rect 352 -734 353 -732
rect 359 -728 360 -726
rect 359 -734 360 -732
rect 369 -728 370 -726
rect 366 -734 367 -732
rect 373 -728 374 -726
rect 373 -734 374 -732
rect 380 -728 381 -726
rect 380 -734 381 -732
rect 387 -728 388 -726
rect 387 -734 388 -732
rect 394 -728 395 -726
rect 397 -728 398 -726
rect 394 -734 395 -732
rect 401 -728 402 -726
rect 401 -734 402 -732
rect 408 -728 409 -726
rect 411 -728 412 -726
rect 408 -734 409 -732
rect 411 -734 412 -732
rect 415 -728 416 -726
rect 415 -734 416 -732
rect 422 -728 423 -726
rect 422 -734 423 -732
rect 429 -728 430 -726
rect 432 -728 433 -726
rect 429 -734 430 -732
rect 436 -728 437 -726
rect 439 -728 440 -726
rect 436 -734 437 -732
rect 443 -728 444 -726
rect 443 -734 444 -732
rect 450 -734 451 -732
rect 457 -728 458 -726
rect 457 -734 458 -732
rect 467 -728 468 -726
rect 464 -734 465 -732
rect 467 -734 468 -732
rect 474 -728 475 -726
rect 471 -734 472 -732
rect 474 -734 475 -732
rect 478 -728 479 -726
rect 478 -734 479 -732
rect 485 -728 486 -726
rect 485 -734 486 -732
rect 492 -728 493 -726
rect 492 -734 493 -732
rect 499 -728 500 -726
rect 499 -734 500 -732
rect 506 -728 507 -726
rect 506 -734 507 -732
rect 513 -728 514 -726
rect 513 -734 514 -732
rect 520 -728 521 -726
rect 520 -734 521 -732
rect 527 -728 528 -726
rect 527 -734 528 -732
rect 534 -728 535 -726
rect 534 -734 535 -732
rect 541 -728 542 -726
rect 541 -734 542 -732
rect 548 -728 549 -726
rect 548 -734 549 -732
rect 555 -728 556 -726
rect 555 -734 556 -732
rect 562 -728 563 -726
rect 562 -734 563 -732
rect 569 -728 570 -726
rect 569 -734 570 -732
rect 576 -728 577 -726
rect 576 -734 577 -732
rect 583 -728 584 -726
rect 583 -734 584 -732
rect 590 -728 591 -726
rect 590 -734 591 -732
rect 600 -734 601 -732
rect 604 -728 605 -726
rect 604 -734 605 -732
rect 611 -728 612 -726
rect 611 -734 612 -732
rect 618 -728 619 -726
rect 618 -734 619 -732
rect 625 -728 626 -726
rect 625 -734 626 -732
rect 632 -728 633 -726
rect 632 -734 633 -732
rect 639 -728 640 -726
rect 639 -734 640 -732
rect 646 -728 647 -726
rect 646 -734 647 -732
rect 653 -728 654 -726
rect 653 -734 654 -732
rect 660 -728 661 -726
rect 660 -734 661 -732
rect 667 -728 668 -726
rect 667 -734 668 -732
rect 674 -728 675 -726
rect 674 -734 675 -732
rect 681 -728 682 -726
rect 681 -734 682 -732
rect 688 -728 689 -726
rect 688 -734 689 -732
rect 695 -728 696 -726
rect 695 -734 696 -732
rect 702 -728 703 -726
rect 702 -734 703 -732
rect 709 -728 710 -726
rect 709 -734 710 -732
rect 716 -728 717 -726
rect 716 -734 717 -732
rect 723 -728 724 -726
rect 723 -734 724 -732
rect 730 -728 731 -726
rect 730 -734 731 -732
rect 737 -728 738 -726
rect 737 -734 738 -732
rect 744 -728 745 -726
rect 744 -734 745 -732
rect 751 -728 752 -726
rect 751 -734 752 -732
rect 758 -728 759 -726
rect 758 -734 759 -732
rect 765 -728 766 -726
rect 765 -734 766 -732
rect 772 -728 773 -726
rect 772 -734 773 -732
rect 779 -728 780 -726
rect 779 -734 780 -732
rect 786 -728 787 -726
rect 786 -734 787 -732
rect 793 -728 794 -726
rect 793 -734 794 -732
rect 800 -728 801 -726
rect 800 -734 801 -732
rect 807 -728 808 -726
rect 807 -734 808 -732
rect 814 -728 815 -726
rect 814 -734 815 -732
rect 817 -734 818 -732
rect 824 -728 825 -726
rect 821 -734 822 -732
rect 824 -734 825 -732
rect 828 -728 829 -726
rect 828 -734 829 -732
rect 9 -817 10 -815
rect 9 -823 10 -821
rect 16 -817 17 -815
rect 23 -817 24 -815
rect 23 -823 24 -821
rect 30 -817 31 -815
rect 30 -823 31 -821
rect 37 -817 38 -815
rect 40 -817 41 -815
rect 37 -823 38 -821
rect 47 -817 48 -815
rect 44 -823 45 -821
rect 51 -823 52 -821
rect 58 -817 59 -815
rect 58 -823 59 -821
rect 65 -823 66 -821
rect 68 -823 69 -821
rect 72 -817 73 -815
rect 72 -823 73 -821
rect 82 -817 83 -815
rect 82 -823 83 -821
rect 86 -817 87 -815
rect 86 -823 87 -821
rect 93 -817 94 -815
rect 96 -817 97 -815
rect 93 -823 94 -821
rect 96 -823 97 -821
rect 100 -817 101 -815
rect 100 -823 101 -821
rect 107 -817 108 -815
rect 107 -823 108 -821
rect 114 -817 115 -815
rect 114 -823 115 -821
rect 121 -817 122 -815
rect 121 -823 122 -821
rect 128 -817 129 -815
rect 128 -823 129 -821
rect 135 -817 136 -815
rect 135 -823 136 -821
rect 142 -817 143 -815
rect 142 -823 143 -821
rect 149 -817 150 -815
rect 149 -823 150 -821
rect 152 -823 153 -821
rect 156 -817 157 -815
rect 156 -823 157 -821
rect 163 -817 164 -815
rect 163 -823 164 -821
rect 170 -817 171 -815
rect 170 -823 171 -821
rect 177 -817 178 -815
rect 177 -823 178 -821
rect 187 -817 188 -815
rect 187 -823 188 -821
rect 191 -817 192 -815
rect 191 -823 192 -821
rect 198 -817 199 -815
rect 198 -823 199 -821
rect 205 -817 206 -815
rect 212 -817 213 -815
rect 212 -823 213 -821
rect 219 -817 220 -815
rect 219 -823 220 -821
rect 226 -817 227 -815
rect 226 -823 227 -821
rect 233 -817 234 -815
rect 233 -823 234 -821
rect 240 -817 241 -815
rect 240 -823 241 -821
rect 247 -817 248 -815
rect 247 -823 248 -821
rect 254 -817 255 -815
rect 254 -823 255 -821
rect 261 -817 262 -815
rect 261 -823 262 -821
rect 268 -817 269 -815
rect 271 -817 272 -815
rect 268 -823 269 -821
rect 275 -817 276 -815
rect 275 -823 276 -821
rect 282 -817 283 -815
rect 282 -823 283 -821
rect 289 -817 290 -815
rect 289 -823 290 -821
rect 296 -817 297 -815
rect 296 -823 297 -821
rect 306 -817 307 -815
rect 303 -823 304 -821
rect 306 -823 307 -821
rect 310 -817 311 -815
rect 310 -823 311 -821
rect 317 -817 318 -815
rect 317 -823 318 -821
rect 324 -817 325 -815
rect 324 -823 325 -821
rect 331 -817 332 -815
rect 331 -823 332 -821
rect 338 -817 339 -815
rect 341 -817 342 -815
rect 338 -823 339 -821
rect 345 -817 346 -815
rect 348 -817 349 -815
rect 345 -823 346 -821
rect 348 -823 349 -821
rect 352 -817 353 -815
rect 352 -823 353 -821
rect 359 -817 360 -815
rect 359 -823 360 -821
rect 366 -817 367 -815
rect 369 -817 370 -815
rect 366 -823 367 -821
rect 369 -823 370 -821
rect 373 -817 374 -815
rect 373 -823 374 -821
rect 380 -817 381 -815
rect 383 -823 384 -821
rect 387 -817 388 -815
rect 390 -817 391 -815
rect 387 -823 388 -821
rect 390 -823 391 -821
rect 394 -817 395 -815
rect 394 -823 395 -821
rect 404 -817 405 -815
rect 404 -823 405 -821
rect 408 -817 409 -815
rect 408 -823 409 -821
rect 415 -817 416 -815
rect 415 -823 416 -821
rect 422 -817 423 -815
rect 422 -823 423 -821
rect 429 -823 430 -821
rect 436 -817 437 -815
rect 439 -817 440 -815
rect 436 -823 437 -821
rect 446 -817 447 -815
rect 443 -823 444 -821
rect 453 -817 454 -815
rect 453 -823 454 -821
rect 457 -817 458 -815
rect 457 -823 458 -821
rect 464 -817 465 -815
rect 464 -823 465 -821
rect 471 -817 472 -815
rect 471 -823 472 -821
rect 478 -817 479 -815
rect 478 -823 479 -821
rect 485 -817 486 -815
rect 485 -823 486 -821
rect 492 -817 493 -815
rect 492 -823 493 -821
rect 499 -817 500 -815
rect 499 -823 500 -821
rect 506 -817 507 -815
rect 506 -823 507 -821
rect 513 -817 514 -815
rect 513 -823 514 -821
rect 520 -817 521 -815
rect 520 -823 521 -821
rect 527 -817 528 -815
rect 527 -823 528 -821
rect 534 -817 535 -815
rect 534 -823 535 -821
rect 541 -817 542 -815
rect 541 -823 542 -821
rect 548 -817 549 -815
rect 548 -823 549 -821
rect 555 -817 556 -815
rect 555 -823 556 -821
rect 562 -817 563 -815
rect 562 -823 563 -821
rect 569 -817 570 -815
rect 569 -823 570 -821
rect 576 -817 577 -815
rect 576 -823 577 -821
rect 583 -817 584 -815
rect 583 -823 584 -821
rect 590 -823 591 -821
rect 597 -817 598 -815
rect 597 -823 598 -821
rect 604 -817 605 -815
rect 604 -823 605 -821
rect 611 -817 612 -815
rect 611 -823 612 -821
rect 618 -817 619 -815
rect 618 -823 619 -821
rect 625 -817 626 -815
rect 625 -823 626 -821
rect 632 -817 633 -815
rect 632 -823 633 -821
rect 635 -823 636 -821
rect 639 -817 640 -815
rect 639 -823 640 -821
rect 646 -817 647 -815
rect 646 -823 647 -821
rect 653 -817 654 -815
rect 653 -823 654 -821
rect 660 -817 661 -815
rect 660 -823 661 -821
rect 667 -817 668 -815
rect 667 -823 668 -821
rect 674 -817 675 -815
rect 674 -823 675 -821
rect 681 -817 682 -815
rect 681 -823 682 -821
rect 688 -817 689 -815
rect 688 -823 689 -821
rect 695 -817 696 -815
rect 695 -823 696 -821
rect 702 -817 703 -815
rect 702 -823 703 -821
rect 709 -817 710 -815
rect 709 -823 710 -821
rect 716 -817 717 -815
rect 716 -823 717 -821
rect 723 -817 724 -815
rect 723 -823 724 -821
rect 730 -817 731 -815
rect 730 -823 731 -821
rect 737 -817 738 -815
rect 737 -823 738 -821
rect 744 -817 745 -815
rect 744 -823 745 -821
rect 751 -817 752 -815
rect 751 -823 752 -821
rect 758 -817 759 -815
rect 758 -823 759 -821
rect 765 -817 766 -815
rect 765 -823 766 -821
rect 772 -817 773 -815
rect 772 -823 773 -821
rect 779 -817 780 -815
rect 779 -823 780 -821
rect 786 -817 787 -815
rect 786 -823 787 -821
rect 793 -817 794 -815
rect 793 -823 794 -821
rect 9 -908 10 -906
rect 16 -902 17 -900
rect 16 -908 17 -906
rect 26 -902 27 -900
rect 23 -908 24 -906
rect 30 -902 31 -900
rect 30 -908 31 -906
rect 37 -902 38 -900
rect 40 -908 41 -906
rect 44 -902 45 -900
rect 44 -908 45 -906
rect 51 -902 52 -900
rect 54 -902 55 -900
rect 58 -902 59 -900
rect 58 -908 59 -906
rect 65 -902 66 -900
rect 65 -908 66 -906
rect 72 -902 73 -900
rect 72 -908 73 -906
rect 79 -902 80 -900
rect 79 -908 80 -906
rect 86 -902 87 -900
rect 86 -908 87 -906
rect 93 -902 94 -900
rect 93 -908 94 -906
rect 100 -908 101 -906
rect 103 -908 104 -906
rect 107 -902 108 -900
rect 107 -908 108 -906
rect 114 -902 115 -900
rect 117 -902 118 -900
rect 117 -908 118 -906
rect 121 -902 122 -900
rect 121 -908 122 -906
rect 128 -902 129 -900
rect 128 -908 129 -906
rect 135 -902 136 -900
rect 135 -908 136 -906
rect 142 -902 143 -900
rect 145 -902 146 -900
rect 145 -908 146 -906
rect 149 -902 150 -900
rect 149 -908 150 -906
rect 156 -902 157 -900
rect 156 -908 157 -906
rect 163 -902 164 -900
rect 163 -908 164 -906
rect 170 -902 171 -900
rect 173 -902 174 -900
rect 173 -908 174 -906
rect 177 -902 178 -900
rect 180 -902 181 -900
rect 180 -908 181 -906
rect 184 -902 185 -900
rect 184 -908 185 -906
rect 191 -902 192 -900
rect 191 -908 192 -906
rect 198 -902 199 -900
rect 198 -908 199 -906
rect 205 -908 206 -906
rect 212 -902 213 -900
rect 212 -908 213 -906
rect 219 -902 220 -900
rect 219 -908 220 -906
rect 226 -902 227 -900
rect 226 -908 227 -906
rect 233 -902 234 -900
rect 233 -908 234 -906
rect 240 -902 241 -900
rect 240 -908 241 -906
rect 247 -902 248 -900
rect 247 -908 248 -906
rect 257 -902 258 -900
rect 254 -908 255 -906
rect 257 -908 258 -906
rect 261 -902 262 -900
rect 261 -908 262 -906
rect 268 -902 269 -900
rect 268 -908 269 -906
rect 275 -902 276 -900
rect 275 -908 276 -906
rect 278 -908 279 -906
rect 285 -902 286 -900
rect 285 -908 286 -906
rect 289 -902 290 -900
rect 299 -902 300 -900
rect 299 -908 300 -906
rect 306 -902 307 -900
rect 306 -908 307 -906
rect 310 -902 311 -900
rect 310 -908 311 -906
rect 317 -902 318 -900
rect 317 -908 318 -906
rect 324 -902 325 -900
rect 324 -908 325 -906
rect 331 -902 332 -900
rect 331 -908 332 -906
rect 341 -902 342 -900
rect 345 -902 346 -900
rect 345 -908 346 -906
rect 352 -902 353 -900
rect 352 -908 353 -906
rect 359 -902 360 -900
rect 362 -902 363 -900
rect 362 -908 363 -906
rect 366 -902 367 -900
rect 366 -908 367 -906
rect 373 -902 374 -900
rect 373 -908 374 -906
rect 380 -902 381 -900
rect 380 -908 381 -906
rect 387 -902 388 -900
rect 387 -908 388 -906
rect 394 -902 395 -900
rect 394 -908 395 -906
rect 404 -902 405 -900
rect 401 -908 402 -906
rect 404 -908 405 -906
rect 411 -902 412 -900
rect 411 -908 412 -906
rect 415 -902 416 -900
rect 415 -908 416 -906
rect 422 -902 423 -900
rect 422 -908 423 -906
rect 429 -902 430 -900
rect 429 -908 430 -906
rect 436 -902 437 -900
rect 436 -908 437 -906
rect 443 -902 444 -900
rect 443 -908 444 -906
rect 450 -902 451 -900
rect 453 -902 454 -900
rect 450 -908 451 -906
rect 457 -902 458 -900
rect 457 -908 458 -906
rect 464 -902 465 -900
rect 464 -908 465 -906
rect 471 -902 472 -900
rect 471 -908 472 -906
rect 478 -902 479 -900
rect 478 -908 479 -906
rect 485 -902 486 -900
rect 485 -908 486 -906
rect 492 -902 493 -900
rect 492 -908 493 -906
rect 499 -902 500 -900
rect 499 -908 500 -906
rect 506 -908 507 -906
rect 509 -908 510 -906
rect 513 -902 514 -900
rect 513 -908 514 -906
rect 520 -902 521 -900
rect 520 -908 521 -906
rect 530 -902 531 -900
rect 527 -908 528 -906
rect 534 -902 535 -900
rect 537 -902 538 -900
rect 537 -908 538 -906
rect 541 -902 542 -900
rect 541 -908 542 -906
rect 555 -902 556 -900
rect 555 -908 556 -906
rect 562 -902 563 -900
rect 562 -908 563 -906
rect 569 -902 570 -900
rect 569 -908 570 -906
rect 576 -902 577 -900
rect 576 -908 577 -906
rect 583 -902 584 -900
rect 583 -908 584 -906
rect 590 -908 591 -906
rect 597 -902 598 -900
rect 597 -908 598 -906
rect 604 -902 605 -900
rect 604 -908 605 -906
rect 618 -902 619 -900
rect 618 -908 619 -906
rect 625 -902 626 -900
rect 625 -908 626 -906
rect 632 -902 633 -900
rect 635 -902 636 -900
rect 632 -908 633 -906
rect 639 -902 640 -900
rect 639 -908 640 -906
rect 646 -902 647 -900
rect 646 -908 647 -906
rect 653 -902 654 -900
rect 653 -908 654 -906
rect 660 -902 661 -900
rect 660 -908 661 -906
rect 667 -902 668 -900
rect 667 -908 668 -906
rect 674 -902 675 -900
rect 674 -908 675 -906
rect 681 -902 682 -900
rect 681 -908 682 -906
rect 688 -902 689 -900
rect 688 -908 689 -906
rect 695 -902 696 -900
rect 695 -908 696 -906
rect 702 -902 703 -900
rect 702 -908 703 -906
rect 709 -902 710 -900
rect 709 -908 710 -906
rect 737 -902 738 -900
rect 737 -908 738 -906
rect 758 -902 759 -900
rect 758 -908 759 -906
rect 2 -985 3 -983
rect 2 -991 3 -989
rect 9 -991 10 -989
rect 16 -985 17 -983
rect 16 -991 17 -989
rect 26 -985 27 -983
rect 26 -991 27 -989
rect 30 -985 31 -983
rect 30 -991 31 -989
rect 37 -985 38 -983
rect 37 -991 38 -989
rect 44 -985 45 -983
rect 47 -985 48 -983
rect 44 -991 45 -989
rect 47 -991 48 -989
rect 51 -985 52 -983
rect 54 -985 55 -983
rect 58 -985 59 -983
rect 61 -985 62 -983
rect 65 -985 66 -983
rect 68 -991 69 -989
rect 72 -985 73 -983
rect 72 -991 73 -989
rect 79 -985 80 -983
rect 79 -991 80 -989
rect 86 -991 87 -989
rect 89 -991 90 -989
rect 93 -985 94 -983
rect 93 -991 94 -989
rect 100 -985 101 -983
rect 100 -991 101 -989
rect 107 -985 108 -983
rect 107 -991 108 -989
rect 114 -985 115 -983
rect 114 -991 115 -989
rect 121 -985 122 -983
rect 121 -991 122 -989
rect 128 -985 129 -983
rect 128 -991 129 -989
rect 135 -985 136 -983
rect 135 -991 136 -989
rect 142 -985 143 -983
rect 145 -985 146 -983
rect 142 -991 143 -989
rect 149 -985 150 -983
rect 152 -985 153 -983
rect 149 -991 150 -989
rect 156 -985 157 -983
rect 156 -991 157 -989
rect 163 -985 164 -983
rect 163 -991 164 -989
rect 170 -985 171 -983
rect 170 -991 171 -989
rect 180 -985 181 -983
rect 177 -991 178 -989
rect 180 -991 181 -989
rect 184 -985 185 -983
rect 187 -985 188 -983
rect 184 -991 185 -989
rect 187 -991 188 -989
rect 191 -985 192 -983
rect 191 -991 192 -989
rect 198 -985 199 -983
rect 198 -991 199 -989
rect 205 -985 206 -983
rect 205 -991 206 -989
rect 212 -985 213 -983
rect 212 -991 213 -989
rect 219 -985 220 -983
rect 219 -991 220 -989
rect 229 -985 230 -983
rect 226 -991 227 -989
rect 233 -985 234 -983
rect 233 -991 234 -989
rect 240 -985 241 -983
rect 240 -991 241 -989
rect 250 -985 251 -983
rect 250 -991 251 -989
rect 254 -985 255 -983
rect 254 -991 255 -989
rect 261 -985 262 -983
rect 261 -991 262 -989
rect 268 -985 269 -983
rect 268 -991 269 -989
rect 275 -985 276 -983
rect 275 -991 276 -989
rect 282 -985 283 -983
rect 282 -991 283 -989
rect 289 -985 290 -983
rect 292 -991 293 -989
rect 296 -985 297 -983
rect 296 -991 297 -989
rect 303 -985 304 -983
rect 303 -991 304 -989
rect 310 -985 311 -983
rect 313 -985 314 -983
rect 310 -991 311 -989
rect 313 -991 314 -989
rect 317 -985 318 -983
rect 317 -991 318 -989
rect 324 -985 325 -983
rect 324 -991 325 -989
rect 331 -985 332 -983
rect 331 -991 332 -989
rect 338 -985 339 -983
rect 338 -991 339 -989
rect 345 -985 346 -983
rect 345 -991 346 -989
rect 352 -985 353 -983
rect 352 -991 353 -989
rect 359 -985 360 -983
rect 362 -985 363 -983
rect 366 -985 367 -983
rect 366 -991 367 -989
rect 373 -985 374 -983
rect 373 -991 374 -989
rect 383 -985 384 -983
rect 383 -991 384 -989
rect 387 -985 388 -983
rect 387 -991 388 -989
rect 394 -985 395 -983
rect 397 -985 398 -983
rect 394 -991 395 -989
rect 397 -991 398 -989
rect 401 -985 402 -983
rect 401 -991 402 -989
rect 408 -985 409 -983
rect 411 -985 412 -983
rect 411 -991 412 -989
rect 415 -985 416 -983
rect 415 -991 416 -989
rect 422 -985 423 -983
rect 422 -991 423 -989
rect 429 -985 430 -983
rect 429 -991 430 -989
rect 436 -985 437 -983
rect 436 -991 437 -989
rect 443 -985 444 -983
rect 446 -991 447 -989
rect 450 -985 451 -983
rect 450 -991 451 -989
rect 457 -985 458 -983
rect 457 -991 458 -989
rect 464 -985 465 -983
rect 464 -991 465 -989
rect 471 -985 472 -983
rect 471 -991 472 -989
rect 478 -985 479 -983
rect 478 -991 479 -989
rect 485 -991 486 -989
rect 488 -991 489 -989
rect 492 -985 493 -983
rect 492 -991 493 -989
rect 499 -985 500 -983
rect 502 -985 503 -983
rect 502 -991 503 -989
rect 506 -985 507 -983
rect 506 -991 507 -989
rect 513 -985 514 -983
rect 513 -991 514 -989
rect 520 -985 521 -983
rect 520 -991 521 -989
rect 527 -985 528 -983
rect 527 -991 528 -989
rect 534 -985 535 -983
rect 534 -991 535 -989
rect 541 -985 542 -983
rect 541 -991 542 -989
rect 548 -985 549 -983
rect 548 -991 549 -989
rect 555 -985 556 -983
rect 555 -991 556 -989
rect 562 -985 563 -983
rect 562 -991 563 -989
rect 569 -985 570 -983
rect 569 -991 570 -989
rect 576 -985 577 -983
rect 576 -991 577 -989
rect 583 -985 584 -983
rect 583 -991 584 -989
rect 590 -985 591 -983
rect 590 -991 591 -989
rect 604 -985 605 -983
rect 607 -985 608 -983
rect 604 -991 605 -989
rect 607 -991 608 -989
rect 611 -985 612 -983
rect 611 -991 612 -989
rect 621 -985 622 -983
rect 621 -991 622 -989
rect 625 -985 626 -983
rect 625 -991 626 -989
rect 632 -985 633 -983
rect 632 -991 633 -989
rect 639 -985 640 -983
rect 639 -991 640 -989
rect 646 -985 647 -983
rect 646 -991 647 -989
rect 653 -985 654 -983
rect 653 -991 654 -989
rect 660 -985 661 -983
rect 660 -991 661 -989
rect 667 -985 668 -983
rect 667 -991 668 -989
rect 674 -985 675 -983
rect 674 -991 675 -989
rect 681 -985 682 -983
rect 681 -991 682 -989
rect 688 -985 689 -983
rect 688 -991 689 -989
rect 695 -985 696 -983
rect 695 -991 696 -989
rect 702 -985 703 -983
rect 702 -991 703 -989
rect 709 -985 710 -983
rect 709 -991 710 -989
rect 716 -985 717 -983
rect 716 -991 717 -989
rect 726 -985 727 -983
rect 751 -985 752 -983
rect 751 -991 752 -989
rect 9 -1066 10 -1064
rect 16 -1060 17 -1058
rect 16 -1066 17 -1064
rect 23 -1060 24 -1058
rect 26 -1066 27 -1064
rect 30 -1060 31 -1058
rect 30 -1066 31 -1064
rect 37 -1060 38 -1058
rect 37 -1066 38 -1064
rect 47 -1066 48 -1064
rect 54 -1060 55 -1058
rect 51 -1066 52 -1064
rect 58 -1060 59 -1058
rect 58 -1066 59 -1064
rect 65 -1060 66 -1058
rect 65 -1066 66 -1064
rect 75 -1060 76 -1058
rect 79 -1060 80 -1058
rect 79 -1066 80 -1064
rect 86 -1060 87 -1058
rect 86 -1066 87 -1064
rect 93 -1060 94 -1058
rect 93 -1066 94 -1064
rect 100 -1060 101 -1058
rect 103 -1060 104 -1058
rect 103 -1066 104 -1064
rect 107 -1060 108 -1058
rect 107 -1066 108 -1064
rect 117 -1060 118 -1058
rect 114 -1066 115 -1064
rect 121 -1060 122 -1058
rect 121 -1066 122 -1064
rect 128 -1060 129 -1058
rect 128 -1066 129 -1064
rect 135 -1060 136 -1058
rect 135 -1066 136 -1064
rect 138 -1066 139 -1064
rect 142 -1060 143 -1058
rect 142 -1066 143 -1064
rect 149 -1060 150 -1058
rect 149 -1066 150 -1064
rect 156 -1060 157 -1058
rect 156 -1066 157 -1064
rect 163 -1060 164 -1058
rect 163 -1066 164 -1064
rect 170 -1060 171 -1058
rect 173 -1066 174 -1064
rect 177 -1060 178 -1058
rect 177 -1066 178 -1064
rect 184 -1060 185 -1058
rect 184 -1066 185 -1064
rect 187 -1066 188 -1064
rect 191 -1060 192 -1058
rect 191 -1066 192 -1064
rect 198 -1060 199 -1058
rect 198 -1066 199 -1064
rect 205 -1060 206 -1058
rect 205 -1066 206 -1064
rect 212 -1060 213 -1058
rect 212 -1066 213 -1064
rect 219 -1060 220 -1058
rect 219 -1066 220 -1064
rect 226 -1060 227 -1058
rect 226 -1066 227 -1064
rect 233 -1060 234 -1058
rect 233 -1066 234 -1064
rect 240 -1060 241 -1058
rect 240 -1066 241 -1064
rect 247 -1060 248 -1058
rect 247 -1066 248 -1064
rect 254 -1060 255 -1058
rect 254 -1066 255 -1064
rect 261 -1060 262 -1058
rect 261 -1066 262 -1064
rect 268 -1060 269 -1058
rect 271 -1066 272 -1064
rect 275 -1060 276 -1058
rect 275 -1066 276 -1064
rect 282 -1066 283 -1064
rect 289 -1060 290 -1058
rect 289 -1066 290 -1064
rect 296 -1060 297 -1058
rect 296 -1066 297 -1064
rect 303 -1060 304 -1058
rect 306 -1060 307 -1058
rect 303 -1066 304 -1064
rect 306 -1066 307 -1064
rect 310 -1060 311 -1058
rect 310 -1066 311 -1064
rect 317 -1060 318 -1058
rect 320 -1060 321 -1058
rect 317 -1066 318 -1064
rect 324 -1060 325 -1058
rect 324 -1066 325 -1064
rect 331 -1060 332 -1058
rect 331 -1066 332 -1064
rect 338 -1060 339 -1058
rect 338 -1066 339 -1064
rect 345 -1060 346 -1058
rect 345 -1066 346 -1064
rect 352 -1060 353 -1058
rect 355 -1060 356 -1058
rect 359 -1060 360 -1058
rect 362 -1060 363 -1058
rect 362 -1066 363 -1064
rect 366 -1060 367 -1058
rect 369 -1060 370 -1058
rect 366 -1066 367 -1064
rect 373 -1060 374 -1058
rect 376 -1066 377 -1064
rect 380 -1060 381 -1058
rect 380 -1066 381 -1064
rect 387 -1060 388 -1058
rect 387 -1066 388 -1064
rect 394 -1060 395 -1058
rect 397 -1066 398 -1064
rect 401 -1060 402 -1058
rect 404 -1060 405 -1058
rect 408 -1060 409 -1058
rect 408 -1066 409 -1064
rect 415 -1066 416 -1064
rect 418 -1066 419 -1064
rect 422 -1060 423 -1058
rect 425 -1060 426 -1058
rect 425 -1066 426 -1064
rect 429 -1060 430 -1058
rect 429 -1066 430 -1064
rect 436 -1060 437 -1058
rect 436 -1066 437 -1064
rect 443 -1060 444 -1058
rect 443 -1066 444 -1064
rect 450 -1060 451 -1058
rect 450 -1066 451 -1064
rect 457 -1060 458 -1058
rect 457 -1066 458 -1064
rect 464 -1060 465 -1058
rect 464 -1066 465 -1064
rect 471 -1060 472 -1058
rect 471 -1066 472 -1064
rect 478 -1060 479 -1058
rect 478 -1066 479 -1064
rect 485 -1060 486 -1058
rect 485 -1066 486 -1064
rect 492 -1060 493 -1058
rect 492 -1066 493 -1064
rect 499 -1060 500 -1058
rect 499 -1066 500 -1064
rect 506 -1060 507 -1058
rect 506 -1066 507 -1064
rect 513 -1060 514 -1058
rect 513 -1066 514 -1064
rect 520 -1060 521 -1058
rect 520 -1066 521 -1064
rect 527 -1060 528 -1058
rect 527 -1066 528 -1064
rect 534 -1060 535 -1058
rect 534 -1066 535 -1064
rect 541 -1060 542 -1058
rect 541 -1066 542 -1064
rect 548 -1060 549 -1058
rect 548 -1066 549 -1064
rect 555 -1060 556 -1058
rect 555 -1066 556 -1064
rect 562 -1060 563 -1058
rect 562 -1066 563 -1064
rect 569 -1060 570 -1058
rect 569 -1066 570 -1064
rect 576 -1060 577 -1058
rect 576 -1066 577 -1064
rect 583 -1060 584 -1058
rect 583 -1066 584 -1064
rect 590 -1060 591 -1058
rect 590 -1066 591 -1064
rect 597 -1060 598 -1058
rect 597 -1066 598 -1064
rect 604 -1066 605 -1064
rect 611 -1060 612 -1058
rect 611 -1066 612 -1064
rect 618 -1060 619 -1058
rect 618 -1066 619 -1064
rect 625 -1060 626 -1058
rect 625 -1066 626 -1064
rect 632 -1060 633 -1058
rect 632 -1066 633 -1064
rect 639 -1060 640 -1058
rect 639 -1066 640 -1064
rect 646 -1060 647 -1058
rect 646 -1066 647 -1064
rect 653 -1060 654 -1058
rect 653 -1066 654 -1064
rect 660 -1060 661 -1058
rect 660 -1066 661 -1064
rect 667 -1060 668 -1058
rect 667 -1066 668 -1064
rect 674 -1060 675 -1058
rect 674 -1066 675 -1064
rect 681 -1060 682 -1058
rect 681 -1066 682 -1064
rect 688 -1060 689 -1058
rect 688 -1066 689 -1064
rect 695 -1060 696 -1058
rect 695 -1066 696 -1064
rect 702 -1060 703 -1058
rect 702 -1066 703 -1064
rect 709 -1060 710 -1058
rect 709 -1066 710 -1064
rect 716 -1060 717 -1058
rect 716 -1066 717 -1064
rect 723 -1060 724 -1058
rect 723 -1066 724 -1064
rect 730 -1060 731 -1058
rect 730 -1066 731 -1064
rect 754 -1066 755 -1064
rect 758 -1060 759 -1058
rect 758 -1066 759 -1064
rect 9 -1127 10 -1125
rect 9 -1133 10 -1131
rect 16 -1127 17 -1125
rect 16 -1133 17 -1131
rect 23 -1127 24 -1125
rect 26 -1133 27 -1131
rect 37 -1127 38 -1125
rect 37 -1133 38 -1131
rect 44 -1127 45 -1125
rect 44 -1133 45 -1131
rect 51 -1127 52 -1125
rect 51 -1133 52 -1131
rect 58 -1127 59 -1125
rect 58 -1133 59 -1131
rect 65 -1127 66 -1125
rect 65 -1133 66 -1131
rect 72 -1127 73 -1125
rect 72 -1133 73 -1131
rect 79 -1127 80 -1125
rect 79 -1133 80 -1131
rect 86 -1127 87 -1125
rect 89 -1127 90 -1125
rect 93 -1127 94 -1125
rect 93 -1133 94 -1131
rect 100 -1127 101 -1125
rect 100 -1133 101 -1131
rect 107 -1127 108 -1125
rect 107 -1133 108 -1131
rect 114 -1127 115 -1125
rect 117 -1127 118 -1125
rect 114 -1133 115 -1131
rect 117 -1133 118 -1131
rect 121 -1127 122 -1125
rect 121 -1133 122 -1131
rect 128 -1127 129 -1125
rect 128 -1133 129 -1131
rect 138 -1127 139 -1125
rect 135 -1133 136 -1131
rect 138 -1133 139 -1131
rect 142 -1127 143 -1125
rect 142 -1133 143 -1131
rect 149 -1127 150 -1125
rect 152 -1133 153 -1131
rect 156 -1127 157 -1125
rect 156 -1133 157 -1131
rect 163 -1127 164 -1125
rect 166 -1127 167 -1125
rect 163 -1133 164 -1131
rect 170 -1127 171 -1125
rect 170 -1133 171 -1131
rect 177 -1127 178 -1125
rect 180 -1127 181 -1125
rect 180 -1133 181 -1131
rect 184 -1127 185 -1125
rect 187 -1127 188 -1125
rect 187 -1133 188 -1131
rect 191 -1127 192 -1125
rect 194 -1127 195 -1125
rect 194 -1133 195 -1131
rect 198 -1127 199 -1125
rect 198 -1133 199 -1131
rect 205 -1127 206 -1125
rect 208 -1127 209 -1125
rect 208 -1133 209 -1131
rect 212 -1127 213 -1125
rect 212 -1133 213 -1131
rect 219 -1127 220 -1125
rect 219 -1133 220 -1131
rect 226 -1127 227 -1125
rect 226 -1133 227 -1131
rect 233 -1127 234 -1125
rect 233 -1133 234 -1131
rect 240 -1127 241 -1125
rect 240 -1133 241 -1131
rect 247 -1127 248 -1125
rect 250 -1127 251 -1125
rect 247 -1133 248 -1131
rect 250 -1133 251 -1131
rect 254 -1127 255 -1125
rect 254 -1133 255 -1131
rect 261 -1127 262 -1125
rect 261 -1133 262 -1131
rect 268 -1127 269 -1125
rect 268 -1133 269 -1131
rect 275 -1127 276 -1125
rect 275 -1133 276 -1131
rect 282 -1127 283 -1125
rect 282 -1133 283 -1131
rect 289 -1127 290 -1125
rect 292 -1133 293 -1131
rect 296 -1127 297 -1125
rect 296 -1133 297 -1131
rect 303 -1127 304 -1125
rect 303 -1133 304 -1131
rect 310 -1127 311 -1125
rect 310 -1133 311 -1131
rect 317 -1127 318 -1125
rect 320 -1127 321 -1125
rect 317 -1133 318 -1131
rect 324 -1127 325 -1125
rect 327 -1127 328 -1125
rect 324 -1133 325 -1131
rect 327 -1133 328 -1131
rect 331 -1127 332 -1125
rect 331 -1133 332 -1131
rect 338 -1127 339 -1125
rect 338 -1133 339 -1131
rect 345 -1127 346 -1125
rect 345 -1133 346 -1131
rect 352 -1133 353 -1131
rect 355 -1133 356 -1131
rect 359 -1127 360 -1125
rect 359 -1133 360 -1131
rect 366 -1127 367 -1125
rect 369 -1127 370 -1125
rect 366 -1133 367 -1131
rect 369 -1133 370 -1131
rect 373 -1127 374 -1125
rect 373 -1133 374 -1131
rect 380 -1127 381 -1125
rect 383 -1127 384 -1125
rect 380 -1133 381 -1131
rect 387 -1127 388 -1125
rect 387 -1133 388 -1131
rect 394 -1127 395 -1125
rect 394 -1133 395 -1131
rect 401 -1127 402 -1125
rect 401 -1133 402 -1131
rect 408 -1127 409 -1125
rect 408 -1133 409 -1131
rect 415 -1127 416 -1125
rect 415 -1133 416 -1131
rect 422 -1127 423 -1125
rect 425 -1127 426 -1125
rect 425 -1133 426 -1131
rect 429 -1127 430 -1125
rect 429 -1133 430 -1131
rect 432 -1133 433 -1131
rect 436 -1127 437 -1125
rect 439 -1127 440 -1125
rect 443 -1127 444 -1125
rect 443 -1133 444 -1131
rect 450 -1127 451 -1125
rect 450 -1133 451 -1131
rect 457 -1127 458 -1125
rect 457 -1133 458 -1131
rect 464 -1127 465 -1125
rect 464 -1133 465 -1131
rect 471 -1127 472 -1125
rect 474 -1127 475 -1125
rect 471 -1133 472 -1131
rect 474 -1133 475 -1131
rect 478 -1127 479 -1125
rect 478 -1133 479 -1131
rect 485 -1127 486 -1125
rect 485 -1133 486 -1131
rect 492 -1127 493 -1125
rect 492 -1133 493 -1131
rect 499 -1127 500 -1125
rect 499 -1133 500 -1131
rect 509 -1127 510 -1125
rect 509 -1133 510 -1131
rect 513 -1127 514 -1125
rect 513 -1133 514 -1131
rect 520 -1127 521 -1125
rect 520 -1133 521 -1131
rect 527 -1127 528 -1125
rect 527 -1133 528 -1131
rect 534 -1127 535 -1125
rect 534 -1133 535 -1131
rect 541 -1127 542 -1125
rect 541 -1133 542 -1131
rect 548 -1127 549 -1125
rect 548 -1133 549 -1131
rect 555 -1127 556 -1125
rect 555 -1133 556 -1131
rect 562 -1127 563 -1125
rect 562 -1133 563 -1131
rect 569 -1127 570 -1125
rect 569 -1133 570 -1131
rect 576 -1127 577 -1125
rect 576 -1133 577 -1131
rect 583 -1127 584 -1125
rect 583 -1133 584 -1131
rect 590 -1127 591 -1125
rect 590 -1133 591 -1131
rect 597 -1127 598 -1125
rect 597 -1133 598 -1131
rect 604 -1127 605 -1125
rect 604 -1133 605 -1131
rect 625 -1127 626 -1125
rect 625 -1133 626 -1131
rect 632 -1127 633 -1125
rect 632 -1133 633 -1131
rect 639 -1127 640 -1125
rect 639 -1133 640 -1131
rect 646 -1127 647 -1125
rect 646 -1133 647 -1131
rect 653 -1127 654 -1125
rect 653 -1133 654 -1131
rect 660 -1127 661 -1125
rect 660 -1133 661 -1131
rect 667 -1127 668 -1125
rect 667 -1133 668 -1131
rect 674 -1127 675 -1125
rect 674 -1133 675 -1131
rect 681 -1127 682 -1125
rect 681 -1133 682 -1131
rect 695 -1127 696 -1125
rect 695 -1133 696 -1131
rect 702 -1127 703 -1125
rect 702 -1133 703 -1131
rect 709 -1127 710 -1125
rect 709 -1133 710 -1131
rect 716 -1127 717 -1125
rect 716 -1133 717 -1131
rect 723 -1127 724 -1125
rect 723 -1133 724 -1131
rect 730 -1127 731 -1125
rect 730 -1133 731 -1131
rect 737 -1127 738 -1125
rect 740 -1127 741 -1125
rect 737 -1133 738 -1131
rect 740 -1133 741 -1131
rect 747 -1133 748 -1131
rect 751 -1127 752 -1125
rect 754 -1127 755 -1125
rect 751 -1133 752 -1131
rect 758 -1127 759 -1125
rect 758 -1133 759 -1131
rect 779 -1127 780 -1125
rect 779 -1133 780 -1131
rect 786 -1127 787 -1125
rect 786 -1133 787 -1131
rect 793 -1127 794 -1125
rect 793 -1133 794 -1131
rect 814 -1127 815 -1125
rect 814 -1133 815 -1131
rect 9 -1208 10 -1206
rect 9 -1214 10 -1212
rect 16 -1208 17 -1206
rect 16 -1214 17 -1212
rect 23 -1208 24 -1206
rect 23 -1214 24 -1212
rect 30 -1208 31 -1206
rect 33 -1208 34 -1206
rect 30 -1214 31 -1212
rect 33 -1214 34 -1212
rect 40 -1208 41 -1206
rect 44 -1208 45 -1206
rect 44 -1214 45 -1212
rect 51 -1208 52 -1206
rect 54 -1208 55 -1206
rect 51 -1214 52 -1212
rect 54 -1214 55 -1212
rect 58 -1208 59 -1206
rect 58 -1214 59 -1212
rect 65 -1208 66 -1206
rect 68 -1208 69 -1206
rect 68 -1214 69 -1212
rect 72 -1208 73 -1206
rect 72 -1214 73 -1212
rect 79 -1208 80 -1206
rect 79 -1214 80 -1212
rect 89 -1214 90 -1212
rect 93 -1208 94 -1206
rect 93 -1214 94 -1212
rect 100 -1208 101 -1206
rect 100 -1214 101 -1212
rect 107 -1208 108 -1206
rect 107 -1214 108 -1212
rect 117 -1208 118 -1206
rect 114 -1214 115 -1212
rect 121 -1208 122 -1206
rect 121 -1214 122 -1212
rect 128 -1208 129 -1206
rect 128 -1214 129 -1212
rect 135 -1208 136 -1206
rect 135 -1214 136 -1212
rect 145 -1208 146 -1206
rect 142 -1214 143 -1212
rect 145 -1214 146 -1212
rect 149 -1208 150 -1206
rect 149 -1214 150 -1212
rect 156 -1208 157 -1206
rect 156 -1214 157 -1212
rect 166 -1208 167 -1206
rect 170 -1208 171 -1206
rect 170 -1214 171 -1212
rect 177 -1208 178 -1206
rect 177 -1214 178 -1212
rect 187 -1208 188 -1206
rect 184 -1214 185 -1212
rect 191 -1208 192 -1206
rect 191 -1214 192 -1212
rect 198 -1208 199 -1206
rect 198 -1214 199 -1212
rect 205 -1208 206 -1206
rect 205 -1214 206 -1212
rect 212 -1208 213 -1206
rect 212 -1214 213 -1212
rect 219 -1208 220 -1206
rect 219 -1214 220 -1212
rect 226 -1208 227 -1206
rect 226 -1214 227 -1212
rect 236 -1208 237 -1206
rect 233 -1214 234 -1212
rect 240 -1208 241 -1206
rect 240 -1214 241 -1212
rect 247 -1208 248 -1206
rect 247 -1214 248 -1212
rect 257 -1208 258 -1206
rect 254 -1214 255 -1212
rect 261 -1208 262 -1206
rect 261 -1214 262 -1212
rect 268 -1208 269 -1206
rect 268 -1214 269 -1212
rect 275 -1208 276 -1206
rect 275 -1214 276 -1212
rect 278 -1214 279 -1212
rect 282 -1208 283 -1206
rect 282 -1214 283 -1212
rect 289 -1208 290 -1206
rect 289 -1214 290 -1212
rect 296 -1208 297 -1206
rect 296 -1214 297 -1212
rect 303 -1208 304 -1206
rect 303 -1214 304 -1212
rect 310 -1208 311 -1206
rect 310 -1214 311 -1212
rect 320 -1208 321 -1206
rect 317 -1214 318 -1212
rect 324 -1208 325 -1206
rect 324 -1214 325 -1212
rect 327 -1214 328 -1212
rect 331 -1208 332 -1206
rect 331 -1214 332 -1212
rect 338 -1208 339 -1206
rect 341 -1208 342 -1206
rect 341 -1214 342 -1212
rect 345 -1208 346 -1206
rect 348 -1208 349 -1206
rect 345 -1214 346 -1212
rect 348 -1214 349 -1212
rect 352 -1208 353 -1206
rect 352 -1214 353 -1212
rect 359 -1208 360 -1206
rect 359 -1214 360 -1212
rect 366 -1208 367 -1206
rect 369 -1208 370 -1206
rect 366 -1214 367 -1212
rect 373 -1208 374 -1206
rect 373 -1214 374 -1212
rect 380 -1208 381 -1206
rect 380 -1214 381 -1212
rect 390 -1208 391 -1206
rect 390 -1214 391 -1212
rect 394 -1208 395 -1206
rect 397 -1208 398 -1206
rect 397 -1214 398 -1212
rect 404 -1208 405 -1206
rect 401 -1214 402 -1212
rect 404 -1214 405 -1212
rect 411 -1208 412 -1206
rect 408 -1214 409 -1212
rect 411 -1214 412 -1212
rect 415 -1208 416 -1206
rect 415 -1214 416 -1212
rect 422 -1208 423 -1206
rect 422 -1214 423 -1212
rect 429 -1208 430 -1206
rect 429 -1214 430 -1212
rect 436 -1208 437 -1206
rect 436 -1214 437 -1212
rect 443 -1208 444 -1206
rect 443 -1214 444 -1212
rect 450 -1208 451 -1206
rect 450 -1214 451 -1212
rect 457 -1208 458 -1206
rect 457 -1214 458 -1212
rect 467 -1208 468 -1206
rect 464 -1214 465 -1212
rect 471 -1208 472 -1206
rect 474 -1214 475 -1212
rect 478 -1208 479 -1206
rect 478 -1214 479 -1212
rect 481 -1214 482 -1212
rect 485 -1208 486 -1206
rect 485 -1214 486 -1212
rect 492 -1208 493 -1206
rect 492 -1214 493 -1212
rect 499 -1208 500 -1206
rect 499 -1214 500 -1212
rect 506 -1208 507 -1206
rect 506 -1214 507 -1212
rect 513 -1208 514 -1206
rect 513 -1214 514 -1212
rect 520 -1208 521 -1206
rect 520 -1214 521 -1212
rect 527 -1208 528 -1206
rect 527 -1214 528 -1212
rect 534 -1208 535 -1206
rect 534 -1214 535 -1212
rect 541 -1214 542 -1212
rect 548 -1208 549 -1206
rect 548 -1214 549 -1212
rect 555 -1208 556 -1206
rect 555 -1214 556 -1212
rect 562 -1208 563 -1206
rect 562 -1214 563 -1212
rect 569 -1208 570 -1206
rect 569 -1214 570 -1212
rect 576 -1208 577 -1206
rect 576 -1214 577 -1212
rect 583 -1208 584 -1206
rect 583 -1214 584 -1212
rect 593 -1208 594 -1206
rect 593 -1214 594 -1212
rect 597 -1208 598 -1206
rect 597 -1214 598 -1212
rect 604 -1208 605 -1206
rect 604 -1214 605 -1212
rect 611 -1208 612 -1206
rect 611 -1214 612 -1212
rect 618 -1208 619 -1206
rect 618 -1214 619 -1212
rect 625 -1208 626 -1206
rect 625 -1214 626 -1212
rect 632 -1208 633 -1206
rect 632 -1214 633 -1212
rect 639 -1208 640 -1206
rect 639 -1214 640 -1212
rect 646 -1208 647 -1206
rect 646 -1214 647 -1212
rect 653 -1208 654 -1206
rect 653 -1214 654 -1212
rect 663 -1214 664 -1212
rect 667 -1208 668 -1206
rect 667 -1214 668 -1212
rect 674 -1208 675 -1206
rect 674 -1214 675 -1212
rect 681 -1208 682 -1206
rect 681 -1214 682 -1212
rect 688 -1208 689 -1206
rect 688 -1214 689 -1212
rect 695 -1208 696 -1206
rect 695 -1214 696 -1212
rect 702 -1208 703 -1206
rect 702 -1214 703 -1212
rect 709 -1208 710 -1206
rect 709 -1214 710 -1212
rect 716 -1208 717 -1206
rect 716 -1214 717 -1212
rect 723 -1208 724 -1206
rect 723 -1214 724 -1212
rect 730 -1208 731 -1206
rect 730 -1214 731 -1212
rect 744 -1208 745 -1206
rect 744 -1214 745 -1212
rect 751 -1208 752 -1206
rect 751 -1214 752 -1212
rect 758 -1208 759 -1206
rect 758 -1214 759 -1212
rect 765 -1208 766 -1206
rect 765 -1214 766 -1212
rect 772 -1208 773 -1206
rect 772 -1214 773 -1212
rect 779 -1208 780 -1206
rect 779 -1214 780 -1212
rect 786 -1208 787 -1206
rect 786 -1214 787 -1212
rect 793 -1208 794 -1206
rect 793 -1214 794 -1212
rect 800 -1208 801 -1206
rect 800 -1214 801 -1212
rect 2 -1301 3 -1299
rect 2 -1307 3 -1305
rect 9 -1301 10 -1299
rect 9 -1307 10 -1305
rect 16 -1301 17 -1299
rect 16 -1307 17 -1305
rect 23 -1301 24 -1299
rect 23 -1307 24 -1305
rect 30 -1301 31 -1299
rect 30 -1307 31 -1305
rect 37 -1301 38 -1299
rect 37 -1307 38 -1305
rect 44 -1301 45 -1299
rect 44 -1307 45 -1305
rect 51 -1301 52 -1299
rect 51 -1307 52 -1305
rect 58 -1301 59 -1299
rect 58 -1307 59 -1305
rect 65 -1301 66 -1299
rect 65 -1307 66 -1305
rect 68 -1307 69 -1305
rect 72 -1301 73 -1299
rect 75 -1301 76 -1299
rect 75 -1307 76 -1305
rect 79 -1301 80 -1299
rect 79 -1307 80 -1305
rect 86 -1301 87 -1299
rect 86 -1307 87 -1305
rect 93 -1301 94 -1299
rect 93 -1307 94 -1305
rect 100 -1301 101 -1299
rect 100 -1307 101 -1305
rect 107 -1301 108 -1299
rect 107 -1307 108 -1305
rect 114 -1307 115 -1305
rect 117 -1307 118 -1305
rect 121 -1301 122 -1299
rect 121 -1307 122 -1305
rect 128 -1301 129 -1299
rect 128 -1307 129 -1305
rect 135 -1301 136 -1299
rect 135 -1307 136 -1305
rect 145 -1301 146 -1299
rect 142 -1307 143 -1305
rect 149 -1301 150 -1299
rect 149 -1307 150 -1305
rect 156 -1301 157 -1299
rect 156 -1307 157 -1305
rect 166 -1301 167 -1299
rect 163 -1307 164 -1305
rect 166 -1307 167 -1305
rect 170 -1301 171 -1299
rect 170 -1307 171 -1305
rect 177 -1301 178 -1299
rect 177 -1307 178 -1305
rect 184 -1301 185 -1299
rect 187 -1301 188 -1299
rect 184 -1307 185 -1305
rect 187 -1307 188 -1305
rect 191 -1301 192 -1299
rect 191 -1307 192 -1305
rect 198 -1301 199 -1299
rect 198 -1307 199 -1305
rect 201 -1307 202 -1305
rect 205 -1301 206 -1299
rect 205 -1307 206 -1305
rect 212 -1301 213 -1299
rect 212 -1307 213 -1305
rect 219 -1301 220 -1299
rect 219 -1307 220 -1305
rect 229 -1307 230 -1305
rect 233 -1301 234 -1299
rect 233 -1307 234 -1305
rect 240 -1301 241 -1299
rect 240 -1307 241 -1305
rect 247 -1301 248 -1299
rect 247 -1307 248 -1305
rect 254 -1301 255 -1299
rect 254 -1307 255 -1305
rect 261 -1301 262 -1299
rect 261 -1307 262 -1305
rect 268 -1301 269 -1299
rect 268 -1307 269 -1305
rect 275 -1301 276 -1299
rect 275 -1307 276 -1305
rect 282 -1301 283 -1299
rect 282 -1307 283 -1305
rect 289 -1301 290 -1299
rect 289 -1307 290 -1305
rect 296 -1301 297 -1299
rect 296 -1307 297 -1305
rect 303 -1301 304 -1299
rect 303 -1307 304 -1305
rect 310 -1301 311 -1299
rect 313 -1307 314 -1305
rect 317 -1301 318 -1299
rect 317 -1307 318 -1305
rect 324 -1301 325 -1299
rect 324 -1307 325 -1305
rect 334 -1301 335 -1299
rect 334 -1307 335 -1305
rect 338 -1301 339 -1299
rect 341 -1301 342 -1299
rect 345 -1301 346 -1299
rect 345 -1307 346 -1305
rect 352 -1307 353 -1305
rect 355 -1307 356 -1305
rect 362 -1301 363 -1299
rect 359 -1307 360 -1305
rect 362 -1307 363 -1305
rect 366 -1307 367 -1305
rect 373 -1301 374 -1299
rect 373 -1307 374 -1305
rect 380 -1301 381 -1299
rect 380 -1307 381 -1305
rect 387 -1301 388 -1299
rect 387 -1307 388 -1305
rect 394 -1301 395 -1299
rect 394 -1307 395 -1305
rect 401 -1301 402 -1299
rect 404 -1301 405 -1299
rect 401 -1307 402 -1305
rect 408 -1301 409 -1299
rect 411 -1301 412 -1299
rect 408 -1307 409 -1305
rect 411 -1307 412 -1305
rect 415 -1301 416 -1299
rect 415 -1307 416 -1305
rect 422 -1301 423 -1299
rect 422 -1307 423 -1305
rect 425 -1307 426 -1305
rect 429 -1301 430 -1299
rect 429 -1307 430 -1305
rect 436 -1301 437 -1299
rect 436 -1307 437 -1305
rect 443 -1301 444 -1299
rect 443 -1307 444 -1305
rect 450 -1301 451 -1299
rect 450 -1307 451 -1305
rect 457 -1301 458 -1299
rect 457 -1307 458 -1305
rect 464 -1301 465 -1299
rect 464 -1307 465 -1305
rect 471 -1301 472 -1299
rect 471 -1307 472 -1305
rect 478 -1301 479 -1299
rect 478 -1307 479 -1305
rect 485 -1301 486 -1299
rect 485 -1307 486 -1305
rect 492 -1301 493 -1299
rect 492 -1307 493 -1305
rect 499 -1301 500 -1299
rect 499 -1307 500 -1305
rect 506 -1301 507 -1299
rect 506 -1307 507 -1305
rect 513 -1301 514 -1299
rect 513 -1307 514 -1305
rect 520 -1301 521 -1299
rect 520 -1307 521 -1305
rect 527 -1301 528 -1299
rect 527 -1307 528 -1305
rect 534 -1301 535 -1299
rect 534 -1307 535 -1305
rect 537 -1307 538 -1305
rect 541 -1301 542 -1299
rect 541 -1307 542 -1305
rect 548 -1301 549 -1299
rect 548 -1307 549 -1305
rect 555 -1301 556 -1299
rect 555 -1307 556 -1305
rect 562 -1301 563 -1299
rect 562 -1307 563 -1305
rect 572 -1301 573 -1299
rect 572 -1307 573 -1305
rect 576 -1301 577 -1299
rect 576 -1307 577 -1305
rect 583 -1301 584 -1299
rect 583 -1307 584 -1305
rect 590 -1301 591 -1299
rect 590 -1307 591 -1305
rect 597 -1301 598 -1299
rect 597 -1307 598 -1305
rect 604 -1301 605 -1299
rect 604 -1307 605 -1305
rect 611 -1301 612 -1299
rect 611 -1307 612 -1305
rect 618 -1301 619 -1299
rect 618 -1307 619 -1305
rect 625 -1301 626 -1299
rect 625 -1307 626 -1305
rect 632 -1301 633 -1299
rect 632 -1307 633 -1305
rect 639 -1301 640 -1299
rect 639 -1307 640 -1305
rect 646 -1301 647 -1299
rect 649 -1301 650 -1299
rect 653 -1301 654 -1299
rect 653 -1307 654 -1305
rect 660 -1301 661 -1299
rect 660 -1307 661 -1305
rect 667 -1301 668 -1299
rect 667 -1307 668 -1305
rect 674 -1301 675 -1299
rect 674 -1307 675 -1305
rect 681 -1301 682 -1299
rect 681 -1307 682 -1305
rect 688 -1301 689 -1299
rect 688 -1307 689 -1305
rect 695 -1301 696 -1299
rect 695 -1307 696 -1305
rect 702 -1301 703 -1299
rect 702 -1307 703 -1305
rect 709 -1301 710 -1299
rect 709 -1307 710 -1305
rect 716 -1301 717 -1299
rect 716 -1307 717 -1305
rect 723 -1301 724 -1299
rect 723 -1307 724 -1305
rect 730 -1301 731 -1299
rect 730 -1307 731 -1305
rect 737 -1301 738 -1299
rect 737 -1307 738 -1305
rect 744 -1301 745 -1299
rect 744 -1307 745 -1305
rect 751 -1301 752 -1299
rect 751 -1307 752 -1305
rect 758 -1301 759 -1299
rect 758 -1307 759 -1305
rect 768 -1307 769 -1305
rect 772 -1301 773 -1299
rect 779 -1301 780 -1299
rect 782 -1301 783 -1299
rect 782 -1307 783 -1305
rect 786 -1301 787 -1299
rect 789 -1301 790 -1299
rect 9 -1378 10 -1376
rect 23 -1378 24 -1376
rect 23 -1384 24 -1382
rect 30 -1378 31 -1376
rect 30 -1384 31 -1382
rect 40 -1378 41 -1376
rect 44 -1378 45 -1376
rect 44 -1384 45 -1382
rect 51 -1378 52 -1376
rect 51 -1384 52 -1382
rect 58 -1378 59 -1376
rect 58 -1384 59 -1382
rect 65 -1378 66 -1376
rect 65 -1384 66 -1382
rect 72 -1378 73 -1376
rect 75 -1384 76 -1382
rect 79 -1378 80 -1376
rect 82 -1378 83 -1376
rect 79 -1384 80 -1382
rect 89 -1384 90 -1382
rect 93 -1378 94 -1376
rect 93 -1384 94 -1382
rect 100 -1378 101 -1376
rect 100 -1384 101 -1382
rect 107 -1378 108 -1376
rect 107 -1384 108 -1382
rect 114 -1378 115 -1376
rect 117 -1378 118 -1376
rect 117 -1384 118 -1382
rect 121 -1378 122 -1376
rect 121 -1384 122 -1382
rect 128 -1378 129 -1376
rect 128 -1384 129 -1382
rect 135 -1378 136 -1376
rect 135 -1384 136 -1382
rect 142 -1378 143 -1376
rect 145 -1378 146 -1376
rect 142 -1384 143 -1382
rect 149 -1378 150 -1376
rect 149 -1384 150 -1382
rect 156 -1378 157 -1376
rect 156 -1384 157 -1382
rect 163 -1378 164 -1376
rect 163 -1384 164 -1382
rect 166 -1384 167 -1382
rect 170 -1378 171 -1376
rect 170 -1384 171 -1382
rect 177 -1378 178 -1376
rect 180 -1378 181 -1376
rect 177 -1384 178 -1382
rect 180 -1384 181 -1382
rect 184 -1378 185 -1376
rect 187 -1378 188 -1376
rect 184 -1384 185 -1382
rect 191 -1378 192 -1376
rect 191 -1384 192 -1382
rect 198 -1378 199 -1376
rect 198 -1384 199 -1382
rect 205 -1378 206 -1376
rect 205 -1384 206 -1382
rect 212 -1378 213 -1376
rect 215 -1378 216 -1376
rect 215 -1384 216 -1382
rect 219 -1378 220 -1376
rect 219 -1384 220 -1382
rect 226 -1378 227 -1376
rect 226 -1384 227 -1382
rect 233 -1378 234 -1376
rect 233 -1384 234 -1382
rect 240 -1378 241 -1376
rect 240 -1384 241 -1382
rect 247 -1378 248 -1376
rect 247 -1384 248 -1382
rect 254 -1378 255 -1376
rect 254 -1384 255 -1382
rect 261 -1378 262 -1376
rect 261 -1384 262 -1382
rect 268 -1378 269 -1376
rect 268 -1384 269 -1382
rect 275 -1378 276 -1376
rect 275 -1384 276 -1382
rect 278 -1384 279 -1382
rect 282 -1378 283 -1376
rect 282 -1384 283 -1382
rect 289 -1378 290 -1376
rect 289 -1384 290 -1382
rect 296 -1378 297 -1376
rect 296 -1384 297 -1382
rect 299 -1384 300 -1382
rect 303 -1378 304 -1376
rect 303 -1384 304 -1382
rect 310 -1378 311 -1376
rect 310 -1384 311 -1382
rect 317 -1378 318 -1376
rect 320 -1378 321 -1376
rect 317 -1384 318 -1382
rect 324 -1378 325 -1376
rect 324 -1384 325 -1382
rect 331 -1378 332 -1376
rect 334 -1378 335 -1376
rect 331 -1384 332 -1382
rect 338 -1378 339 -1376
rect 338 -1384 339 -1382
rect 348 -1378 349 -1376
rect 348 -1384 349 -1382
rect 352 -1378 353 -1376
rect 352 -1384 353 -1382
rect 359 -1378 360 -1376
rect 359 -1384 360 -1382
rect 366 -1378 367 -1376
rect 366 -1384 367 -1382
rect 373 -1378 374 -1376
rect 373 -1384 374 -1382
rect 380 -1378 381 -1376
rect 380 -1384 381 -1382
rect 387 -1378 388 -1376
rect 387 -1384 388 -1382
rect 394 -1378 395 -1376
rect 394 -1384 395 -1382
rect 401 -1378 402 -1376
rect 404 -1378 405 -1376
rect 404 -1384 405 -1382
rect 408 -1378 409 -1376
rect 408 -1384 409 -1382
rect 411 -1384 412 -1382
rect 415 -1378 416 -1376
rect 415 -1384 416 -1382
rect 422 -1378 423 -1376
rect 422 -1384 423 -1382
rect 429 -1378 430 -1376
rect 429 -1384 430 -1382
rect 436 -1378 437 -1376
rect 436 -1384 437 -1382
rect 443 -1378 444 -1376
rect 446 -1378 447 -1376
rect 443 -1384 444 -1382
rect 450 -1378 451 -1376
rect 450 -1384 451 -1382
rect 457 -1378 458 -1376
rect 457 -1384 458 -1382
rect 464 -1378 465 -1376
rect 464 -1384 465 -1382
rect 471 -1378 472 -1376
rect 471 -1384 472 -1382
rect 478 -1378 479 -1376
rect 481 -1378 482 -1376
rect 478 -1384 479 -1382
rect 485 -1378 486 -1376
rect 485 -1384 486 -1382
rect 492 -1378 493 -1376
rect 492 -1384 493 -1382
rect 499 -1378 500 -1376
rect 499 -1384 500 -1382
rect 506 -1378 507 -1376
rect 506 -1384 507 -1382
rect 513 -1378 514 -1376
rect 516 -1378 517 -1376
rect 513 -1384 514 -1382
rect 516 -1384 517 -1382
rect 520 -1378 521 -1376
rect 520 -1384 521 -1382
rect 527 -1378 528 -1376
rect 527 -1384 528 -1382
rect 534 -1378 535 -1376
rect 534 -1384 535 -1382
rect 541 -1378 542 -1376
rect 541 -1384 542 -1382
rect 548 -1378 549 -1376
rect 548 -1384 549 -1382
rect 555 -1378 556 -1376
rect 555 -1384 556 -1382
rect 562 -1378 563 -1376
rect 565 -1378 566 -1376
rect 565 -1384 566 -1382
rect 572 -1384 573 -1382
rect 576 -1378 577 -1376
rect 576 -1384 577 -1382
rect 583 -1378 584 -1376
rect 583 -1384 584 -1382
rect 590 -1378 591 -1376
rect 590 -1384 591 -1382
rect 597 -1378 598 -1376
rect 597 -1384 598 -1382
rect 604 -1378 605 -1376
rect 604 -1384 605 -1382
rect 611 -1378 612 -1376
rect 611 -1384 612 -1382
rect 618 -1378 619 -1376
rect 618 -1384 619 -1382
rect 632 -1378 633 -1376
rect 632 -1384 633 -1382
rect 639 -1378 640 -1376
rect 639 -1384 640 -1382
rect 646 -1378 647 -1376
rect 646 -1384 647 -1382
rect 653 -1378 654 -1376
rect 653 -1384 654 -1382
rect 660 -1378 661 -1376
rect 660 -1384 661 -1382
rect 667 -1378 668 -1376
rect 667 -1384 668 -1382
rect 674 -1378 675 -1376
rect 674 -1384 675 -1382
rect 681 -1378 682 -1376
rect 681 -1384 682 -1382
rect 688 -1378 689 -1376
rect 691 -1378 692 -1376
rect 688 -1384 689 -1382
rect 691 -1384 692 -1382
rect 695 -1378 696 -1376
rect 695 -1384 696 -1382
rect 702 -1378 703 -1376
rect 705 -1378 706 -1376
rect 705 -1384 706 -1382
rect 709 -1378 710 -1376
rect 709 -1384 710 -1382
rect 716 -1384 717 -1382
rect 758 -1378 759 -1376
rect 758 -1384 759 -1382
rect 779 -1378 780 -1376
rect 779 -1384 780 -1382
rect 800 -1378 801 -1376
rect 800 -1384 801 -1382
rect 9 -1447 10 -1445
rect 9 -1453 10 -1451
rect 16 -1447 17 -1445
rect 16 -1453 17 -1451
rect 23 -1447 24 -1445
rect 23 -1453 24 -1451
rect 30 -1447 31 -1445
rect 30 -1453 31 -1451
rect 37 -1447 38 -1445
rect 37 -1453 38 -1451
rect 44 -1447 45 -1445
rect 44 -1453 45 -1451
rect 51 -1447 52 -1445
rect 58 -1447 59 -1445
rect 58 -1453 59 -1451
rect 65 -1447 66 -1445
rect 65 -1453 66 -1451
rect 75 -1447 76 -1445
rect 79 -1447 80 -1445
rect 79 -1453 80 -1451
rect 86 -1447 87 -1445
rect 86 -1453 87 -1451
rect 93 -1447 94 -1445
rect 93 -1453 94 -1451
rect 100 -1447 101 -1445
rect 107 -1447 108 -1445
rect 107 -1453 108 -1451
rect 117 -1447 118 -1445
rect 117 -1453 118 -1451
rect 121 -1453 122 -1451
rect 124 -1453 125 -1451
rect 128 -1447 129 -1445
rect 128 -1453 129 -1451
rect 138 -1447 139 -1445
rect 135 -1453 136 -1451
rect 138 -1453 139 -1451
rect 142 -1447 143 -1445
rect 142 -1453 143 -1451
rect 149 -1447 150 -1445
rect 149 -1453 150 -1451
rect 156 -1453 157 -1451
rect 159 -1453 160 -1451
rect 163 -1447 164 -1445
rect 163 -1453 164 -1451
rect 170 -1447 171 -1445
rect 170 -1453 171 -1451
rect 177 -1447 178 -1445
rect 177 -1453 178 -1451
rect 184 -1453 185 -1451
rect 187 -1453 188 -1451
rect 191 -1447 192 -1445
rect 191 -1453 192 -1451
rect 198 -1447 199 -1445
rect 198 -1453 199 -1451
rect 205 -1447 206 -1445
rect 205 -1453 206 -1451
rect 212 -1447 213 -1445
rect 212 -1453 213 -1451
rect 219 -1447 220 -1445
rect 219 -1453 220 -1451
rect 226 -1447 227 -1445
rect 226 -1453 227 -1451
rect 233 -1447 234 -1445
rect 233 -1453 234 -1451
rect 240 -1447 241 -1445
rect 240 -1453 241 -1451
rect 247 -1447 248 -1445
rect 247 -1453 248 -1451
rect 254 -1447 255 -1445
rect 254 -1453 255 -1451
rect 261 -1447 262 -1445
rect 261 -1453 262 -1451
rect 268 -1447 269 -1445
rect 271 -1447 272 -1445
rect 271 -1453 272 -1451
rect 275 -1447 276 -1445
rect 275 -1453 276 -1451
rect 282 -1447 283 -1445
rect 282 -1453 283 -1451
rect 289 -1447 290 -1445
rect 289 -1453 290 -1451
rect 296 -1447 297 -1445
rect 296 -1453 297 -1451
rect 303 -1447 304 -1445
rect 303 -1453 304 -1451
rect 310 -1447 311 -1445
rect 310 -1453 311 -1451
rect 317 -1447 318 -1445
rect 317 -1453 318 -1451
rect 324 -1447 325 -1445
rect 324 -1453 325 -1451
rect 334 -1447 335 -1445
rect 331 -1453 332 -1451
rect 334 -1453 335 -1451
rect 338 -1447 339 -1445
rect 338 -1453 339 -1451
rect 345 -1447 346 -1445
rect 345 -1453 346 -1451
rect 352 -1447 353 -1445
rect 352 -1453 353 -1451
rect 359 -1447 360 -1445
rect 359 -1453 360 -1451
rect 366 -1447 367 -1445
rect 366 -1453 367 -1451
rect 373 -1447 374 -1445
rect 373 -1453 374 -1451
rect 380 -1447 381 -1445
rect 383 -1447 384 -1445
rect 380 -1453 381 -1451
rect 383 -1453 384 -1451
rect 387 -1447 388 -1445
rect 387 -1453 388 -1451
rect 394 -1447 395 -1445
rect 397 -1453 398 -1451
rect 404 -1447 405 -1445
rect 401 -1453 402 -1451
rect 404 -1453 405 -1451
rect 411 -1447 412 -1445
rect 415 -1447 416 -1445
rect 415 -1453 416 -1451
rect 422 -1447 423 -1445
rect 422 -1453 423 -1451
rect 429 -1447 430 -1445
rect 432 -1447 433 -1445
rect 429 -1453 430 -1451
rect 432 -1453 433 -1451
rect 439 -1447 440 -1445
rect 439 -1453 440 -1451
rect 443 -1447 444 -1445
rect 443 -1453 444 -1451
rect 450 -1447 451 -1445
rect 450 -1453 451 -1451
rect 457 -1447 458 -1445
rect 457 -1453 458 -1451
rect 464 -1447 465 -1445
rect 464 -1453 465 -1451
rect 471 -1453 472 -1451
rect 474 -1453 475 -1451
rect 478 -1447 479 -1445
rect 478 -1453 479 -1451
rect 485 -1447 486 -1445
rect 488 -1447 489 -1445
rect 492 -1447 493 -1445
rect 492 -1453 493 -1451
rect 499 -1447 500 -1445
rect 499 -1453 500 -1451
rect 506 -1447 507 -1445
rect 509 -1447 510 -1445
rect 509 -1453 510 -1451
rect 513 -1447 514 -1445
rect 513 -1453 514 -1451
rect 520 -1447 521 -1445
rect 520 -1453 521 -1451
rect 527 -1447 528 -1445
rect 527 -1453 528 -1451
rect 534 -1447 535 -1445
rect 534 -1453 535 -1451
rect 537 -1453 538 -1451
rect 541 -1447 542 -1445
rect 541 -1453 542 -1451
rect 548 -1447 549 -1445
rect 551 -1447 552 -1445
rect 555 -1447 556 -1445
rect 555 -1453 556 -1451
rect 562 -1447 563 -1445
rect 562 -1453 563 -1451
rect 569 -1447 570 -1445
rect 569 -1453 570 -1451
rect 576 -1447 577 -1445
rect 576 -1453 577 -1451
rect 583 -1447 584 -1445
rect 583 -1453 584 -1451
rect 590 -1447 591 -1445
rect 590 -1453 591 -1451
rect 597 -1447 598 -1445
rect 597 -1453 598 -1451
rect 604 -1447 605 -1445
rect 604 -1453 605 -1451
rect 611 -1447 612 -1445
rect 611 -1453 612 -1451
rect 618 -1447 619 -1445
rect 618 -1453 619 -1451
rect 625 -1447 626 -1445
rect 625 -1453 626 -1451
rect 632 -1447 633 -1445
rect 632 -1453 633 -1451
rect 639 -1447 640 -1445
rect 639 -1453 640 -1451
rect 646 -1447 647 -1445
rect 646 -1453 647 -1451
rect 653 -1447 654 -1445
rect 653 -1453 654 -1451
rect 660 -1447 661 -1445
rect 660 -1453 661 -1451
rect 667 -1447 668 -1445
rect 667 -1453 668 -1451
rect 674 -1447 675 -1445
rect 674 -1453 675 -1451
rect 681 -1447 682 -1445
rect 681 -1453 682 -1451
rect 688 -1447 689 -1445
rect 688 -1453 689 -1451
rect 695 -1447 696 -1445
rect 695 -1453 696 -1451
rect 702 -1447 703 -1445
rect 702 -1453 703 -1451
rect 709 -1447 710 -1445
rect 709 -1453 710 -1451
rect 716 -1447 717 -1445
rect 716 -1453 717 -1451
rect 723 -1447 724 -1445
rect 723 -1453 724 -1451
rect 730 -1447 731 -1445
rect 730 -1453 731 -1451
rect 737 -1447 738 -1445
rect 737 -1453 738 -1451
rect 744 -1447 745 -1445
rect 744 -1453 745 -1451
rect 751 -1447 752 -1445
rect 751 -1453 752 -1451
rect 765 -1447 766 -1445
rect 768 -1447 769 -1445
rect 768 -1453 769 -1451
rect 772 -1447 773 -1445
rect 772 -1453 773 -1451
rect 782 -1447 783 -1445
rect 779 -1453 780 -1451
rect 786 -1447 787 -1445
rect 789 -1447 790 -1445
rect 789 -1453 790 -1451
rect 796 -1447 797 -1445
rect 803 -1447 804 -1445
rect 800 -1453 801 -1451
rect 807 -1447 808 -1445
rect 807 -1453 808 -1451
rect 814 -1453 815 -1451
rect 817 -1453 818 -1451
rect 828 -1447 829 -1445
rect 828 -1453 829 -1451
rect 835 -1447 836 -1445
rect 835 -1453 836 -1451
rect 2 -1532 3 -1530
rect 9 -1526 10 -1524
rect 9 -1532 10 -1530
rect 16 -1526 17 -1524
rect 16 -1532 17 -1530
rect 23 -1526 24 -1524
rect 23 -1532 24 -1530
rect 30 -1526 31 -1524
rect 30 -1532 31 -1530
rect 37 -1526 38 -1524
rect 37 -1532 38 -1530
rect 44 -1526 45 -1524
rect 44 -1532 45 -1530
rect 54 -1526 55 -1524
rect 51 -1532 52 -1530
rect 58 -1526 59 -1524
rect 58 -1532 59 -1530
rect 65 -1526 66 -1524
rect 65 -1532 66 -1530
rect 72 -1526 73 -1524
rect 79 -1526 80 -1524
rect 79 -1532 80 -1530
rect 86 -1526 87 -1524
rect 86 -1532 87 -1530
rect 96 -1526 97 -1524
rect 96 -1532 97 -1530
rect 100 -1532 101 -1530
rect 107 -1526 108 -1524
rect 107 -1532 108 -1530
rect 114 -1526 115 -1524
rect 114 -1532 115 -1530
rect 121 -1526 122 -1524
rect 121 -1532 122 -1530
rect 128 -1526 129 -1524
rect 128 -1532 129 -1530
rect 138 -1526 139 -1524
rect 138 -1532 139 -1530
rect 142 -1526 143 -1524
rect 142 -1532 143 -1530
rect 149 -1526 150 -1524
rect 149 -1532 150 -1530
rect 156 -1526 157 -1524
rect 156 -1532 157 -1530
rect 166 -1526 167 -1524
rect 170 -1526 171 -1524
rect 170 -1532 171 -1530
rect 177 -1526 178 -1524
rect 180 -1526 181 -1524
rect 177 -1532 178 -1530
rect 184 -1532 185 -1530
rect 187 -1532 188 -1530
rect 191 -1526 192 -1524
rect 191 -1532 192 -1530
rect 198 -1526 199 -1524
rect 198 -1532 199 -1530
rect 205 -1532 206 -1530
rect 208 -1532 209 -1530
rect 212 -1526 213 -1524
rect 212 -1532 213 -1530
rect 219 -1526 220 -1524
rect 219 -1532 220 -1530
rect 226 -1526 227 -1524
rect 226 -1532 227 -1530
rect 233 -1526 234 -1524
rect 240 -1526 241 -1524
rect 247 -1526 248 -1524
rect 250 -1526 251 -1524
rect 247 -1532 248 -1530
rect 250 -1532 251 -1530
rect 257 -1526 258 -1524
rect 257 -1532 258 -1530
rect 261 -1526 262 -1524
rect 261 -1532 262 -1530
rect 268 -1526 269 -1524
rect 275 -1526 276 -1524
rect 275 -1532 276 -1530
rect 282 -1526 283 -1524
rect 282 -1532 283 -1530
rect 289 -1526 290 -1524
rect 289 -1532 290 -1530
rect 296 -1526 297 -1524
rect 296 -1532 297 -1530
rect 306 -1526 307 -1524
rect 303 -1532 304 -1530
rect 306 -1532 307 -1530
rect 310 -1526 311 -1524
rect 310 -1532 311 -1530
rect 317 -1526 318 -1524
rect 317 -1532 318 -1530
rect 324 -1526 325 -1524
rect 324 -1532 325 -1530
rect 331 -1526 332 -1524
rect 331 -1532 332 -1530
rect 334 -1532 335 -1530
rect 338 -1526 339 -1524
rect 341 -1526 342 -1524
rect 338 -1532 339 -1530
rect 341 -1532 342 -1530
rect 345 -1526 346 -1524
rect 345 -1532 346 -1530
rect 352 -1526 353 -1524
rect 352 -1532 353 -1530
rect 359 -1526 360 -1524
rect 362 -1526 363 -1524
rect 362 -1532 363 -1530
rect 366 -1526 367 -1524
rect 369 -1526 370 -1524
rect 373 -1526 374 -1524
rect 373 -1532 374 -1530
rect 380 -1526 381 -1524
rect 383 -1526 384 -1524
rect 380 -1532 381 -1530
rect 387 -1526 388 -1524
rect 390 -1526 391 -1524
rect 387 -1532 388 -1530
rect 394 -1526 395 -1524
rect 394 -1532 395 -1530
rect 401 -1526 402 -1524
rect 401 -1532 402 -1530
rect 408 -1526 409 -1524
rect 408 -1532 409 -1530
rect 415 -1526 416 -1524
rect 418 -1526 419 -1524
rect 415 -1532 416 -1530
rect 418 -1532 419 -1530
rect 422 -1526 423 -1524
rect 422 -1532 423 -1530
rect 429 -1526 430 -1524
rect 429 -1532 430 -1530
rect 436 -1526 437 -1524
rect 439 -1526 440 -1524
rect 439 -1532 440 -1530
rect 443 -1526 444 -1524
rect 443 -1532 444 -1530
rect 450 -1526 451 -1524
rect 450 -1532 451 -1530
rect 457 -1526 458 -1524
rect 457 -1532 458 -1530
rect 464 -1526 465 -1524
rect 464 -1532 465 -1530
rect 471 -1526 472 -1524
rect 471 -1532 472 -1530
rect 478 -1526 479 -1524
rect 478 -1532 479 -1530
rect 485 -1526 486 -1524
rect 485 -1532 486 -1530
rect 492 -1526 493 -1524
rect 492 -1532 493 -1530
rect 499 -1526 500 -1524
rect 499 -1532 500 -1530
rect 506 -1526 507 -1524
rect 506 -1532 507 -1530
rect 513 -1526 514 -1524
rect 513 -1532 514 -1530
rect 520 -1526 521 -1524
rect 523 -1526 524 -1524
rect 527 -1526 528 -1524
rect 527 -1532 528 -1530
rect 534 -1526 535 -1524
rect 537 -1526 538 -1524
rect 534 -1532 535 -1530
rect 541 -1526 542 -1524
rect 541 -1532 542 -1530
rect 548 -1526 549 -1524
rect 548 -1532 549 -1530
rect 555 -1526 556 -1524
rect 555 -1532 556 -1530
rect 562 -1526 563 -1524
rect 562 -1532 563 -1530
rect 569 -1526 570 -1524
rect 569 -1532 570 -1530
rect 576 -1526 577 -1524
rect 576 -1532 577 -1530
rect 583 -1526 584 -1524
rect 583 -1532 584 -1530
rect 590 -1526 591 -1524
rect 590 -1532 591 -1530
rect 597 -1526 598 -1524
rect 597 -1532 598 -1530
rect 600 -1532 601 -1530
rect 604 -1526 605 -1524
rect 604 -1532 605 -1530
rect 611 -1526 612 -1524
rect 611 -1532 612 -1530
rect 618 -1526 619 -1524
rect 625 -1526 626 -1524
rect 625 -1532 626 -1530
rect 632 -1526 633 -1524
rect 632 -1532 633 -1530
rect 639 -1526 640 -1524
rect 639 -1532 640 -1530
rect 646 -1526 647 -1524
rect 646 -1532 647 -1530
rect 653 -1526 654 -1524
rect 653 -1532 654 -1530
rect 660 -1526 661 -1524
rect 660 -1532 661 -1530
rect 667 -1526 668 -1524
rect 667 -1532 668 -1530
rect 674 -1526 675 -1524
rect 674 -1532 675 -1530
rect 681 -1526 682 -1524
rect 681 -1532 682 -1530
rect 688 -1526 689 -1524
rect 688 -1532 689 -1530
rect 695 -1526 696 -1524
rect 695 -1532 696 -1530
rect 702 -1526 703 -1524
rect 702 -1532 703 -1530
rect 709 -1526 710 -1524
rect 709 -1532 710 -1530
rect 716 -1526 717 -1524
rect 716 -1532 717 -1530
rect 723 -1526 724 -1524
rect 723 -1532 724 -1530
rect 730 -1526 731 -1524
rect 730 -1532 731 -1530
rect 737 -1526 738 -1524
rect 737 -1532 738 -1530
rect 744 -1526 745 -1524
rect 744 -1532 745 -1530
rect 751 -1526 752 -1524
rect 751 -1532 752 -1530
rect 5 -1611 6 -1609
rect 12 -1605 13 -1603
rect 16 -1605 17 -1603
rect 16 -1611 17 -1609
rect 23 -1605 24 -1603
rect 23 -1611 24 -1609
rect 30 -1605 31 -1603
rect 30 -1611 31 -1609
rect 37 -1605 38 -1603
rect 37 -1611 38 -1609
rect 44 -1605 45 -1603
rect 47 -1611 48 -1609
rect 51 -1605 52 -1603
rect 51 -1611 52 -1609
rect 58 -1605 59 -1603
rect 58 -1611 59 -1609
rect 65 -1605 66 -1603
rect 65 -1611 66 -1609
rect 72 -1605 73 -1603
rect 72 -1611 73 -1609
rect 82 -1605 83 -1603
rect 82 -1611 83 -1609
rect 89 -1605 90 -1603
rect 86 -1611 87 -1609
rect 89 -1611 90 -1609
rect 93 -1605 94 -1603
rect 93 -1611 94 -1609
rect 103 -1605 104 -1603
rect 107 -1605 108 -1603
rect 107 -1611 108 -1609
rect 114 -1605 115 -1603
rect 117 -1605 118 -1603
rect 114 -1611 115 -1609
rect 121 -1605 122 -1603
rect 121 -1611 122 -1609
rect 128 -1605 129 -1603
rect 128 -1611 129 -1609
rect 138 -1605 139 -1603
rect 135 -1611 136 -1609
rect 138 -1611 139 -1609
rect 142 -1611 143 -1609
rect 152 -1605 153 -1603
rect 152 -1611 153 -1609
rect 156 -1605 157 -1603
rect 156 -1611 157 -1609
rect 163 -1605 164 -1603
rect 163 -1611 164 -1609
rect 170 -1605 171 -1603
rect 170 -1611 171 -1609
rect 177 -1605 178 -1603
rect 177 -1611 178 -1609
rect 184 -1605 185 -1603
rect 184 -1611 185 -1609
rect 191 -1605 192 -1603
rect 191 -1611 192 -1609
rect 194 -1611 195 -1609
rect 198 -1605 199 -1603
rect 198 -1611 199 -1609
rect 205 -1605 206 -1603
rect 205 -1611 206 -1609
rect 212 -1605 213 -1603
rect 212 -1611 213 -1609
rect 219 -1605 220 -1603
rect 219 -1611 220 -1609
rect 226 -1605 227 -1603
rect 226 -1611 227 -1609
rect 233 -1605 234 -1603
rect 236 -1605 237 -1603
rect 233 -1611 234 -1609
rect 240 -1605 241 -1603
rect 240 -1611 241 -1609
rect 247 -1605 248 -1603
rect 247 -1611 248 -1609
rect 254 -1605 255 -1603
rect 254 -1611 255 -1609
rect 261 -1605 262 -1603
rect 261 -1611 262 -1609
rect 268 -1605 269 -1603
rect 268 -1611 269 -1609
rect 275 -1605 276 -1603
rect 278 -1605 279 -1603
rect 275 -1611 276 -1609
rect 278 -1611 279 -1609
rect 282 -1605 283 -1603
rect 282 -1611 283 -1609
rect 289 -1605 290 -1603
rect 289 -1611 290 -1609
rect 296 -1605 297 -1603
rect 296 -1611 297 -1609
rect 303 -1605 304 -1603
rect 306 -1605 307 -1603
rect 306 -1611 307 -1609
rect 310 -1605 311 -1603
rect 313 -1605 314 -1603
rect 320 -1605 321 -1603
rect 317 -1611 318 -1609
rect 320 -1611 321 -1609
rect 324 -1605 325 -1603
rect 324 -1611 325 -1609
rect 331 -1605 332 -1603
rect 331 -1611 332 -1609
rect 341 -1605 342 -1603
rect 338 -1611 339 -1609
rect 345 -1605 346 -1603
rect 345 -1611 346 -1609
rect 352 -1605 353 -1603
rect 352 -1611 353 -1609
rect 362 -1605 363 -1603
rect 359 -1611 360 -1609
rect 362 -1611 363 -1609
rect 366 -1605 367 -1603
rect 373 -1605 374 -1603
rect 373 -1611 374 -1609
rect 380 -1605 381 -1603
rect 380 -1611 381 -1609
rect 387 -1605 388 -1603
rect 387 -1611 388 -1609
rect 394 -1605 395 -1603
rect 394 -1611 395 -1609
rect 401 -1605 402 -1603
rect 401 -1611 402 -1609
rect 408 -1605 409 -1603
rect 411 -1605 412 -1603
rect 408 -1611 409 -1609
rect 411 -1611 412 -1609
rect 415 -1605 416 -1603
rect 415 -1611 416 -1609
rect 422 -1605 423 -1603
rect 422 -1611 423 -1609
rect 429 -1605 430 -1603
rect 429 -1611 430 -1609
rect 436 -1605 437 -1603
rect 439 -1611 440 -1609
rect 443 -1605 444 -1603
rect 443 -1611 444 -1609
rect 446 -1611 447 -1609
rect 450 -1605 451 -1603
rect 450 -1611 451 -1609
rect 457 -1605 458 -1603
rect 457 -1611 458 -1609
rect 464 -1605 465 -1603
rect 464 -1611 465 -1609
rect 471 -1605 472 -1603
rect 471 -1611 472 -1609
rect 478 -1605 479 -1603
rect 478 -1611 479 -1609
rect 485 -1605 486 -1603
rect 488 -1605 489 -1603
rect 492 -1605 493 -1603
rect 492 -1611 493 -1609
rect 499 -1605 500 -1603
rect 499 -1611 500 -1609
rect 506 -1605 507 -1603
rect 506 -1611 507 -1609
rect 513 -1605 514 -1603
rect 513 -1611 514 -1609
rect 520 -1605 521 -1603
rect 520 -1611 521 -1609
rect 527 -1605 528 -1603
rect 527 -1611 528 -1609
rect 534 -1605 535 -1603
rect 534 -1611 535 -1609
rect 541 -1605 542 -1603
rect 541 -1611 542 -1609
rect 548 -1605 549 -1603
rect 548 -1611 549 -1609
rect 555 -1611 556 -1609
rect 558 -1611 559 -1609
rect 562 -1605 563 -1603
rect 562 -1611 563 -1609
rect 569 -1605 570 -1603
rect 569 -1611 570 -1609
rect 576 -1605 577 -1603
rect 576 -1611 577 -1609
rect 583 -1605 584 -1603
rect 583 -1611 584 -1609
rect 590 -1605 591 -1603
rect 590 -1611 591 -1609
rect 597 -1605 598 -1603
rect 597 -1611 598 -1609
rect 604 -1605 605 -1603
rect 604 -1611 605 -1609
rect 611 -1605 612 -1603
rect 611 -1611 612 -1609
rect 618 -1605 619 -1603
rect 618 -1611 619 -1609
rect 625 -1605 626 -1603
rect 625 -1611 626 -1609
rect 632 -1605 633 -1603
rect 632 -1611 633 -1609
rect 639 -1605 640 -1603
rect 639 -1611 640 -1609
rect 646 -1605 647 -1603
rect 646 -1611 647 -1609
rect 653 -1605 654 -1603
rect 653 -1611 654 -1609
rect 660 -1605 661 -1603
rect 660 -1611 661 -1609
rect 667 -1605 668 -1603
rect 667 -1611 668 -1609
rect 674 -1605 675 -1603
rect 674 -1611 675 -1609
rect 681 -1605 682 -1603
rect 681 -1611 682 -1609
rect 9 -1674 10 -1672
rect 9 -1680 10 -1678
rect 16 -1674 17 -1672
rect 16 -1680 17 -1678
rect 23 -1674 24 -1672
rect 23 -1680 24 -1678
rect 30 -1674 31 -1672
rect 37 -1674 38 -1672
rect 37 -1680 38 -1678
rect 47 -1680 48 -1678
rect 51 -1674 52 -1672
rect 58 -1674 59 -1672
rect 58 -1680 59 -1678
rect 65 -1674 66 -1672
rect 65 -1680 66 -1678
rect 72 -1674 73 -1672
rect 72 -1680 73 -1678
rect 79 -1674 80 -1672
rect 79 -1680 80 -1678
rect 86 -1674 87 -1672
rect 86 -1680 87 -1678
rect 93 -1674 94 -1672
rect 93 -1680 94 -1678
rect 100 -1674 101 -1672
rect 110 -1674 111 -1672
rect 107 -1680 108 -1678
rect 114 -1674 115 -1672
rect 117 -1674 118 -1672
rect 114 -1680 115 -1678
rect 121 -1674 122 -1672
rect 121 -1680 122 -1678
rect 128 -1674 129 -1672
rect 128 -1680 129 -1678
rect 135 -1674 136 -1672
rect 135 -1680 136 -1678
rect 142 -1680 143 -1678
rect 145 -1680 146 -1678
rect 149 -1674 150 -1672
rect 149 -1680 150 -1678
rect 156 -1674 157 -1672
rect 156 -1680 157 -1678
rect 163 -1674 164 -1672
rect 163 -1680 164 -1678
rect 170 -1674 171 -1672
rect 173 -1674 174 -1672
rect 173 -1680 174 -1678
rect 177 -1674 178 -1672
rect 177 -1680 178 -1678
rect 187 -1674 188 -1672
rect 187 -1680 188 -1678
rect 191 -1674 192 -1672
rect 198 -1674 199 -1672
rect 198 -1680 199 -1678
rect 205 -1674 206 -1672
rect 205 -1680 206 -1678
rect 212 -1674 213 -1672
rect 212 -1680 213 -1678
rect 219 -1674 220 -1672
rect 219 -1680 220 -1678
rect 226 -1674 227 -1672
rect 226 -1680 227 -1678
rect 233 -1674 234 -1672
rect 233 -1680 234 -1678
rect 236 -1680 237 -1678
rect 243 -1680 244 -1678
rect 247 -1674 248 -1672
rect 247 -1680 248 -1678
rect 254 -1674 255 -1672
rect 254 -1680 255 -1678
rect 261 -1680 262 -1678
rect 264 -1680 265 -1678
rect 268 -1674 269 -1672
rect 268 -1680 269 -1678
rect 275 -1674 276 -1672
rect 275 -1680 276 -1678
rect 282 -1674 283 -1672
rect 282 -1680 283 -1678
rect 289 -1674 290 -1672
rect 292 -1674 293 -1672
rect 289 -1680 290 -1678
rect 292 -1680 293 -1678
rect 296 -1674 297 -1672
rect 299 -1674 300 -1672
rect 296 -1680 297 -1678
rect 306 -1680 307 -1678
rect 310 -1674 311 -1672
rect 310 -1680 311 -1678
rect 317 -1674 318 -1672
rect 317 -1680 318 -1678
rect 324 -1674 325 -1672
rect 324 -1680 325 -1678
rect 331 -1680 332 -1678
rect 334 -1680 335 -1678
rect 338 -1674 339 -1672
rect 345 -1674 346 -1672
rect 345 -1680 346 -1678
rect 352 -1680 353 -1678
rect 355 -1680 356 -1678
rect 359 -1674 360 -1672
rect 359 -1680 360 -1678
rect 362 -1680 363 -1678
rect 366 -1674 367 -1672
rect 369 -1674 370 -1672
rect 376 -1674 377 -1672
rect 373 -1680 374 -1678
rect 380 -1674 381 -1672
rect 380 -1680 381 -1678
rect 387 -1674 388 -1672
rect 390 -1680 391 -1678
rect 394 -1674 395 -1672
rect 394 -1680 395 -1678
rect 401 -1674 402 -1672
rect 401 -1680 402 -1678
rect 408 -1674 409 -1672
rect 408 -1680 409 -1678
rect 415 -1674 416 -1672
rect 415 -1680 416 -1678
rect 422 -1674 423 -1672
rect 422 -1680 423 -1678
rect 429 -1674 430 -1672
rect 429 -1680 430 -1678
rect 436 -1674 437 -1672
rect 436 -1680 437 -1678
rect 443 -1674 444 -1672
rect 443 -1680 444 -1678
rect 450 -1674 451 -1672
rect 450 -1680 451 -1678
rect 457 -1674 458 -1672
rect 457 -1680 458 -1678
rect 464 -1674 465 -1672
rect 464 -1680 465 -1678
rect 471 -1674 472 -1672
rect 471 -1680 472 -1678
rect 478 -1674 479 -1672
rect 478 -1680 479 -1678
rect 485 -1674 486 -1672
rect 485 -1680 486 -1678
rect 492 -1674 493 -1672
rect 492 -1680 493 -1678
rect 499 -1674 500 -1672
rect 499 -1680 500 -1678
rect 506 -1674 507 -1672
rect 506 -1680 507 -1678
rect 513 -1674 514 -1672
rect 513 -1680 514 -1678
rect 520 -1674 521 -1672
rect 520 -1680 521 -1678
rect 527 -1674 528 -1672
rect 527 -1680 528 -1678
rect 534 -1674 535 -1672
rect 534 -1680 535 -1678
rect 541 -1674 542 -1672
rect 541 -1680 542 -1678
rect 548 -1674 549 -1672
rect 548 -1680 549 -1678
rect 555 -1674 556 -1672
rect 555 -1680 556 -1678
rect 562 -1674 563 -1672
rect 562 -1680 563 -1678
rect 569 -1674 570 -1672
rect 569 -1680 570 -1678
rect 576 -1674 577 -1672
rect 576 -1680 577 -1678
rect 583 -1674 584 -1672
rect 583 -1680 584 -1678
rect 590 -1674 591 -1672
rect 590 -1680 591 -1678
rect 597 -1674 598 -1672
rect 597 -1680 598 -1678
rect 611 -1674 612 -1672
rect 611 -1680 612 -1678
rect 618 -1680 619 -1678
rect 621 -1680 622 -1678
rect 649 -1674 650 -1672
rect 649 -1680 650 -1678
rect 660 -1674 661 -1672
rect 660 -1680 661 -1678
rect 677 -1674 678 -1672
rect 681 -1674 682 -1672
rect 681 -1680 682 -1678
rect 9 -1731 10 -1729
rect 9 -1737 10 -1735
rect 16 -1731 17 -1729
rect 16 -1737 17 -1735
rect 23 -1731 24 -1729
rect 23 -1737 24 -1735
rect 30 -1731 31 -1729
rect 40 -1731 41 -1729
rect 44 -1731 45 -1729
rect 44 -1737 45 -1735
rect 51 -1731 52 -1729
rect 51 -1737 52 -1735
rect 58 -1731 59 -1729
rect 58 -1737 59 -1735
rect 65 -1731 66 -1729
rect 65 -1737 66 -1735
rect 72 -1731 73 -1729
rect 72 -1737 73 -1735
rect 79 -1731 80 -1729
rect 79 -1737 80 -1735
rect 86 -1731 87 -1729
rect 86 -1737 87 -1735
rect 93 -1737 94 -1735
rect 103 -1737 104 -1735
rect 107 -1731 108 -1729
rect 107 -1737 108 -1735
rect 114 -1731 115 -1729
rect 114 -1737 115 -1735
rect 121 -1731 122 -1729
rect 124 -1731 125 -1729
rect 128 -1731 129 -1729
rect 131 -1731 132 -1729
rect 135 -1731 136 -1729
rect 135 -1737 136 -1735
rect 142 -1731 143 -1729
rect 145 -1737 146 -1735
rect 152 -1737 153 -1735
rect 159 -1731 160 -1729
rect 159 -1737 160 -1735
rect 163 -1731 164 -1729
rect 163 -1737 164 -1735
rect 170 -1731 171 -1729
rect 170 -1737 171 -1735
rect 177 -1737 178 -1735
rect 184 -1731 185 -1729
rect 187 -1731 188 -1729
rect 191 -1731 192 -1729
rect 191 -1737 192 -1735
rect 198 -1731 199 -1729
rect 198 -1737 199 -1735
rect 208 -1737 209 -1735
rect 212 -1731 213 -1729
rect 212 -1737 213 -1735
rect 219 -1731 220 -1729
rect 219 -1737 220 -1735
rect 226 -1731 227 -1729
rect 226 -1737 227 -1735
rect 233 -1731 234 -1729
rect 233 -1737 234 -1735
rect 240 -1731 241 -1729
rect 243 -1737 244 -1735
rect 247 -1731 248 -1729
rect 250 -1731 251 -1729
rect 250 -1737 251 -1735
rect 257 -1731 258 -1729
rect 257 -1737 258 -1735
rect 261 -1731 262 -1729
rect 261 -1737 262 -1735
rect 268 -1731 269 -1729
rect 271 -1731 272 -1729
rect 268 -1737 269 -1735
rect 275 -1731 276 -1729
rect 275 -1737 276 -1735
rect 282 -1731 283 -1729
rect 282 -1737 283 -1735
rect 289 -1731 290 -1729
rect 292 -1737 293 -1735
rect 296 -1731 297 -1729
rect 296 -1737 297 -1735
rect 303 -1731 304 -1729
rect 303 -1737 304 -1735
rect 310 -1731 311 -1729
rect 313 -1731 314 -1729
rect 310 -1737 311 -1735
rect 317 -1731 318 -1729
rect 320 -1731 321 -1729
rect 324 -1731 325 -1729
rect 324 -1737 325 -1735
rect 331 -1731 332 -1729
rect 331 -1737 332 -1735
rect 338 -1731 339 -1729
rect 345 -1731 346 -1729
rect 345 -1737 346 -1735
rect 352 -1737 353 -1735
rect 355 -1737 356 -1735
rect 359 -1731 360 -1729
rect 362 -1737 363 -1735
rect 366 -1731 367 -1729
rect 366 -1737 367 -1735
rect 373 -1731 374 -1729
rect 376 -1731 377 -1729
rect 380 -1731 381 -1729
rect 380 -1737 381 -1735
rect 394 -1731 395 -1729
rect 394 -1737 395 -1735
rect 401 -1731 402 -1729
rect 401 -1737 402 -1735
rect 408 -1731 409 -1729
rect 408 -1737 409 -1735
rect 415 -1731 416 -1729
rect 415 -1737 416 -1735
rect 422 -1731 423 -1729
rect 422 -1737 423 -1735
rect 429 -1731 430 -1729
rect 429 -1737 430 -1735
rect 436 -1731 437 -1729
rect 436 -1737 437 -1735
rect 446 -1731 447 -1729
rect 457 -1731 458 -1729
rect 460 -1737 461 -1735
rect 464 -1731 465 -1729
rect 464 -1737 465 -1735
rect 471 -1731 472 -1729
rect 471 -1737 472 -1735
rect 478 -1731 479 -1729
rect 478 -1737 479 -1735
rect 485 -1731 486 -1729
rect 485 -1737 486 -1735
rect 492 -1731 493 -1729
rect 492 -1737 493 -1735
rect 499 -1731 500 -1729
rect 499 -1737 500 -1735
rect 520 -1731 521 -1729
rect 520 -1737 521 -1735
rect 527 -1731 528 -1729
rect 527 -1737 528 -1735
rect 555 -1731 556 -1729
rect 555 -1737 556 -1735
rect 579 -1731 580 -1729
rect 618 -1731 619 -1729
rect 618 -1737 619 -1735
rect 653 -1731 654 -1729
rect 653 -1737 654 -1735
rect 670 -1737 671 -1735
rect 674 -1731 675 -1729
rect 674 -1737 675 -1735
rect 37 -1772 38 -1770
rect 37 -1778 38 -1776
rect 51 -1772 52 -1770
rect 51 -1778 52 -1776
rect 61 -1778 62 -1776
rect 65 -1772 66 -1770
rect 65 -1778 66 -1776
rect 72 -1772 73 -1770
rect 72 -1778 73 -1776
rect 86 -1772 87 -1770
rect 86 -1778 87 -1776
rect 93 -1772 94 -1770
rect 93 -1778 94 -1776
rect 103 -1778 104 -1776
rect 107 -1772 108 -1770
rect 117 -1772 118 -1770
rect 117 -1778 118 -1776
rect 121 -1772 122 -1770
rect 124 -1772 125 -1770
rect 128 -1772 129 -1770
rect 128 -1778 129 -1776
rect 135 -1772 136 -1770
rect 135 -1778 136 -1776
rect 142 -1772 143 -1770
rect 142 -1778 143 -1776
rect 152 -1772 153 -1770
rect 156 -1772 157 -1770
rect 159 -1772 160 -1770
rect 156 -1778 157 -1776
rect 159 -1778 160 -1776
rect 163 -1772 164 -1770
rect 163 -1778 164 -1776
rect 173 -1772 174 -1770
rect 177 -1778 178 -1776
rect 184 -1778 185 -1776
rect 191 -1772 192 -1770
rect 191 -1778 192 -1776
rect 198 -1772 199 -1770
rect 198 -1778 199 -1776
rect 205 -1772 206 -1770
rect 212 -1778 213 -1776
rect 219 -1772 220 -1770
rect 219 -1778 220 -1776
rect 226 -1772 227 -1770
rect 226 -1778 227 -1776
rect 233 -1772 234 -1770
rect 233 -1778 234 -1776
rect 240 -1772 241 -1770
rect 240 -1778 241 -1776
rect 254 -1772 255 -1770
rect 261 -1772 262 -1770
rect 261 -1778 262 -1776
rect 268 -1772 269 -1770
rect 268 -1778 269 -1776
rect 275 -1772 276 -1770
rect 289 -1772 290 -1770
rect 289 -1778 290 -1776
rect 296 -1772 297 -1770
rect 296 -1778 297 -1776
rect 310 -1772 311 -1770
rect 310 -1778 311 -1776
rect 317 -1772 318 -1770
rect 317 -1778 318 -1776
rect 324 -1772 325 -1770
rect 324 -1778 325 -1776
rect 334 -1772 335 -1770
rect 334 -1778 335 -1776
rect 338 -1772 339 -1770
rect 338 -1778 339 -1776
rect 345 -1772 346 -1770
rect 345 -1778 346 -1776
rect 352 -1772 353 -1770
rect 352 -1778 353 -1776
rect 366 -1772 367 -1770
rect 366 -1778 367 -1776
rect 383 -1778 384 -1776
rect 404 -1772 405 -1770
rect 418 -1772 419 -1770
rect 418 -1778 419 -1776
rect 422 -1772 423 -1770
rect 422 -1778 423 -1776
rect 429 -1772 430 -1770
rect 429 -1778 430 -1776
rect 453 -1772 454 -1770
rect 460 -1772 461 -1770
rect 464 -1772 465 -1770
rect 464 -1778 465 -1776
rect 471 -1772 472 -1770
rect 471 -1778 472 -1776
rect 478 -1772 479 -1770
rect 478 -1778 479 -1776
rect 488 -1772 489 -1770
rect 485 -1778 486 -1776
rect 502 -1778 503 -1776
rect 513 -1772 514 -1770
rect 513 -1778 514 -1776
rect 520 -1772 521 -1770
rect 520 -1778 521 -1776
rect 527 -1772 528 -1770
rect 527 -1778 528 -1776
rect 534 -1772 535 -1770
rect 534 -1778 535 -1776
rect 541 -1778 542 -1776
rect 548 -1772 549 -1770
rect 548 -1778 549 -1776
rect 562 -1778 563 -1776
rect 614 -1778 615 -1776
rect 618 -1772 619 -1770
rect 618 -1778 619 -1776
rect 632 -1772 633 -1770
rect 632 -1778 633 -1776
rect 51 -1801 52 -1799
rect 51 -1807 52 -1805
rect 61 -1807 62 -1805
rect 89 -1801 90 -1799
rect 103 -1801 104 -1799
rect 110 -1801 111 -1799
rect 117 -1801 118 -1799
rect 124 -1801 125 -1799
rect 131 -1801 132 -1799
rect 135 -1801 136 -1799
rect 138 -1801 139 -1799
rect 142 -1801 143 -1799
rect 145 -1807 146 -1805
rect 149 -1801 150 -1799
rect 149 -1807 150 -1805
rect 156 -1801 157 -1799
rect 156 -1807 157 -1805
rect 173 -1801 174 -1799
rect 177 -1807 178 -1805
rect 180 -1807 181 -1805
rect 184 -1807 185 -1805
rect 205 -1801 206 -1799
rect 205 -1807 206 -1805
rect 233 -1801 234 -1799
rect 233 -1807 234 -1805
rect 247 -1801 248 -1799
rect 250 -1801 251 -1799
rect 254 -1801 255 -1799
rect 261 -1801 262 -1799
rect 264 -1801 265 -1799
rect 261 -1807 262 -1805
rect 271 -1807 272 -1805
rect 310 -1801 311 -1799
rect 352 -1801 353 -1799
rect 352 -1807 353 -1805
rect 373 -1801 374 -1799
rect 387 -1801 388 -1799
rect 411 -1801 412 -1799
rect 418 -1801 419 -1799
rect 418 -1807 419 -1805
rect 467 -1801 468 -1799
rect 471 -1801 472 -1799
rect 471 -1807 472 -1805
rect 478 -1807 479 -1805
rect 499 -1801 500 -1799
rect 520 -1801 521 -1799
rect 520 -1807 521 -1805
rect 527 -1807 528 -1805
rect 639 -1801 640 -1799
<< metal1 >>
rect 58 0 94 1
rect 114 0 143 1
rect 152 0 171 1
rect 177 0 213 1
rect 257 0 262 1
rect 124 -2 241 -1
rect 128 -4 136 -3
rect 156 -4 164 -3
rect 184 -4 192 -3
rect 198 -4 237 -3
rect 205 -6 339 -5
rect 44 -17 48 -16
rect 72 -17 94 -16
rect 103 -17 276 -16
rect 285 -17 346 -16
rect 79 -19 192 -18
rect 205 -19 318 -18
rect 338 -19 388 -18
rect 114 -21 132 -20
rect 177 -21 199 -20
rect 205 -21 325 -20
rect 124 -23 213 -22
rect 222 -23 241 -22
rect 247 -23 335 -22
rect 128 -25 136 -24
rect 149 -25 178 -24
rect 184 -25 220 -24
rect 240 -25 262 -24
rect 271 -25 353 -24
rect 93 -27 129 -26
rect 163 -27 199 -26
rect 212 -27 227 -26
rect 254 -27 283 -26
rect 289 -27 297 -26
rect 313 -27 339 -26
rect 170 -29 185 -28
rect 226 -29 234 -28
rect 142 -31 234 -30
rect 163 -33 171 -32
rect 16 -44 241 -43
rect 254 -44 342 -43
rect 345 -44 437 -43
rect 23 -46 118 -45
rect 128 -46 157 -45
rect 163 -46 171 -45
rect 191 -46 223 -45
rect 233 -46 311 -45
rect 317 -46 381 -45
rect 387 -46 409 -45
rect 44 -48 59 -47
rect 65 -48 108 -47
rect 114 -48 122 -47
rect 135 -48 143 -47
rect 156 -48 195 -47
rect 205 -48 220 -47
rect 247 -48 255 -47
rect 275 -48 332 -47
rect 338 -48 423 -47
rect 51 -50 346 -49
rect 352 -50 402 -49
rect 404 -50 416 -49
rect 61 -52 206 -51
rect 208 -52 227 -51
rect 268 -52 276 -51
rect 282 -52 318 -51
rect 324 -52 388 -51
rect 72 -54 153 -53
rect 170 -54 181 -53
rect 184 -54 227 -53
rect 296 -54 360 -53
rect 373 -54 395 -53
rect 82 -56 136 -55
rect 184 -56 241 -55
rect 299 -56 367 -55
rect 86 -58 178 -57
rect 212 -58 234 -57
rect 93 -60 325 -59
rect 93 -62 293 -61
rect 100 -64 111 -63
rect 177 -64 199 -63
rect 212 -64 272 -63
rect 198 -66 290 -65
rect 261 -68 272 -67
rect 23 -79 199 -78
rect 205 -79 507 -78
rect 37 -81 220 -80
rect 233 -81 248 -80
rect 250 -81 465 -80
rect 44 -83 297 -82
rect 303 -83 395 -82
rect 397 -83 458 -82
rect 58 -85 157 -84
rect 170 -85 206 -84
rect 208 -85 241 -84
rect 254 -85 269 -84
rect 275 -85 304 -84
rect 373 -85 430 -84
rect 436 -85 514 -84
rect 65 -87 153 -86
rect 156 -87 248 -86
rect 254 -87 318 -86
rect 345 -87 437 -86
rect 72 -89 115 -88
rect 121 -89 199 -88
rect 222 -89 318 -88
rect 338 -89 346 -88
rect 380 -89 472 -88
rect 79 -91 262 -90
rect 275 -91 311 -90
rect 387 -91 493 -90
rect 16 -93 262 -92
rect 285 -93 451 -92
rect 86 -95 101 -94
rect 107 -95 213 -94
rect 292 -95 423 -94
rect 93 -97 444 -96
rect 93 -99 283 -98
rect 310 -99 335 -98
rect 380 -99 423 -98
rect 128 -101 195 -100
rect 212 -101 307 -100
rect 401 -101 500 -100
rect 128 -103 300 -102
rect 359 -103 402 -102
rect 408 -103 486 -102
rect 135 -105 192 -104
rect 324 -105 360 -104
rect 366 -105 409 -104
rect 415 -105 479 -104
rect 149 -107 388 -106
rect 149 -109 164 -108
rect 173 -109 290 -108
rect 331 -109 367 -108
rect 373 -109 416 -108
rect 121 -111 290 -110
rect 331 -111 521 -110
rect 177 -113 234 -112
rect 187 -115 227 -114
rect 142 -117 227 -116
rect 142 -119 185 -118
rect 163 -121 188 -120
rect 12 -132 73 -131
rect 75 -132 507 -131
rect 520 -132 661 -131
rect 51 -134 178 -133
rect 180 -134 360 -133
rect 373 -134 377 -133
rect 383 -134 465 -133
rect 471 -134 619 -133
rect 58 -136 286 -135
rect 296 -136 332 -135
rect 334 -136 444 -135
rect 457 -136 584 -135
rect 58 -138 244 -137
rect 250 -138 269 -137
rect 282 -138 402 -137
rect 415 -138 570 -137
rect 79 -140 402 -139
rect 422 -140 444 -139
rect 478 -140 640 -139
rect 79 -142 104 -141
rect 121 -142 528 -141
rect 44 -144 122 -143
rect 128 -144 381 -143
rect 390 -144 654 -143
rect 44 -146 188 -145
rect 240 -146 276 -145
rect 282 -146 507 -145
rect 513 -146 521 -145
rect 89 -148 199 -147
rect 247 -148 276 -147
rect 292 -148 458 -147
rect 499 -148 633 -147
rect 93 -150 479 -149
rect 485 -150 500 -149
rect 93 -152 272 -151
rect 296 -152 325 -151
rect 327 -152 605 -151
rect 100 -154 563 -153
rect 100 -156 150 -155
rect 152 -156 535 -155
rect 128 -158 220 -157
rect 261 -158 416 -157
rect 422 -158 472 -157
rect 107 -160 262 -159
rect 303 -160 360 -159
rect 373 -160 451 -159
rect 107 -162 160 -161
rect 170 -162 549 -161
rect 117 -164 220 -163
rect 226 -164 304 -163
rect 341 -164 598 -163
rect 135 -166 612 -165
rect 138 -168 143 -167
rect 149 -168 465 -167
rect 142 -170 290 -169
rect 352 -170 493 -169
rect 156 -172 188 -171
rect 191 -172 353 -171
rect 376 -172 451 -171
rect 170 -174 234 -173
rect 289 -174 493 -173
rect 177 -176 591 -175
rect 180 -178 241 -177
rect 387 -178 514 -177
rect 191 -180 255 -179
rect 324 -180 388 -179
rect 394 -180 647 -179
rect 198 -182 626 -181
rect 205 -184 227 -183
rect 317 -184 395 -183
rect 408 -184 486 -183
rect 135 -186 318 -185
rect 408 -186 577 -185
rect 212 -188 234 -187
rect 429 -188 556 -187
rect 366 -190 430 -189
rect 436 -190 542 -189
rect 86 -192 437 -191
rect 345 -194 367 -193
rect 310 -196 346 -195
rect 33 -207 591 -206
rect 597 -207 668 -206
rect 51 -209 213 -208
rect 215 -209 605 -208
rect 65 -211 202 -210
rect 205 -211 241 -210
rect 243 -211 514 -210
rect 520 -211 605 -210
rect 79 -213 307 -212
rect 310 -213 325 -212
rect 338 -213 626 -212
rect 44 -215 325 -214
rect 366 -215 409 -214
rect 411 -215 507 -214
rect 513 -215 528 -214
rect 590 -215 633 -214
rect 89 -217 423 -216
rect 464 -217 521 -216
rect 527 -217 542 -216
rect 597 -217 640 -216
rect 100 -219 181 -218
rect 187 -219 227 -218
rect 254 -219 346 -218
rect 373 -219 542 -218
rect 625 -219 654 -218
rect 103 -221 178 -220
rect 198 -221 458 -220
rect 464 -221 486 -220
rect 632 -221 661 -220
rect 72 -223 199 -222
rect 208 -223 535 -222
rect 72 -225 83 -224
rect 114 -225 185 -224
rect 219 -225 227 -224
rect 247 -225 458 -224
rect 485 -225 563 -224
rect 58 -227 220 -226
rect 257 -227 360 -226
rect 373 -227 402 -226
rect 499 -227 563 -226
rect 58 -229 507 -228
rect 534 -229 556 -228
rect 114 -231 192 -230
rect 257 -231 577 -230
rect 121 -233 346 -232
rect 359 -233 381 -232
rect 387 -233 584 -232
rect 121 -235 584 -234
rect 124 -237 304 -236
rect 313 -237 549 -236
rect 65 -239 304 -238
rect 317 -239 402 -238
rect 548 -239 619 -238
rect 128 -241 381 -240
rect 387 -241 430 -240
rect 576 -241 619 -240
rect 128 -243 241 -242
rect 268 -243 612 -242
rect 135 -245 353 -244
rect 429 -245 472 -244
rect 100 -247 136 -246
rect 142 -247 164 -246
rect 170 -247 213 -246
rect 268 -247 500 -246
rect 93 -249 171 -248
rect 191 -249 251 -248
rect 275 -249 290 -248
rect 292 -249 395 -248
rect 443 -249 472 -248
rect 89 -251 395 -250
rect 436 -251 444 -250
rect 93 -253 297 -252
rect 299 -253 332 -252
rect 334 -253 612 -252
rect 107 -255 164 -254
rect 282 -255 570 -254
rect 107 -257 157 -256
rect 180 -257 570 -256
rect 142 -259 157 -258
rect 320 -259 451 -258
rect 149 -261 234 -260
rect 285 -261 451 -260
rect 23 -263 234 -262
rect 285 -263 416 -262
rect 425 -263 437 -262
rect 152 -265 262 -264
rect 282 -265 416 -264
rect 261 -267 279 -266
rect 331 -267 647 -266
rect 338 -269 367 -268
rect 44 -280 48 -279
rect 58 -280 213 -279
rect 247 -280 346 -279
rect 355 -280 388 -279
rect 390 -280 479 -279
rect 506 -280 619 -279
rect 667 -280 710 -279
rect 58 -282 255 -281
rect 261 -282 276 -281
rect 282 -282 311 -281
rect 317 -282 661 -281
rect 72 -284 178 -283
rect 187 -284 262 -283
rect 282 -284 339 -283
rect 341 -284 521 -283
rect 555 -284 640 -283
rect 72 -286 570 -285
rect 583 -286 640 -285
rect 89 -288 479 -287
rect 513 -288 675 -287
rect 89 -290 486 -289
rect 527 -290 570 -289
rect 590 -290 647 -289
rect 100 -292 654 -291
rect 107 -294 213 -293
rect 285 -294 486 -293
rect 492 -294 528 -293
rect 534 -294 584 -293
rect 604 -294 668 -293
rect 16 -296 605 -295
rect 107 -298 129 -297
rect 145 -298 160 -297
rect 163 -298 255 -297
rect 296 -298 626 -297
rect 54 -300 626 -299
rect 65 -302 297 -301
rect 299 -302 332 -301
rect 362 -302 514 -301
rect 541 -302 591 -301
rect 114 -304 129 -303
rect 149 -304 269 -303
rect 306 -304 633 -303
rect 114 -306 251 -305
rect 320 -306 430 -305
rect 450 -306 507 -305
rect 541 -306 563 -305
rect 30 -308 430 -307
rect 436 -308 451 -307
rect 464 -308 521 -307
rect 562 -308 612 -307
rect 30 -310 83 -309
rect 121 -310 388 -309
rect 415 -310 437 -309
rect 443 -310 465 -309
rect 499 -310 535 -309
rect 576 -310 612 -309
rect 23 -312 122 -311
rect 142 -312 269 -311
rect 320 -312 633 -311
rect 159 -314 381 -313
rect 408 -314 444 -313
rect 471 -314 577 -313
rect 65 -316 409 -315
rect 415 -316 423 -315
rect 457 -316 472 -315
rect 79 -318 458 -317
rect 51 -320 80 -319
rect 142 -320 381 -319
rect 394 -320 423 -319
rect 37 -322 52 -321
rect 170 -322 178 -321
rect 191 -322 335 -321
rect 352 -322 395 -321
rect 135 -324 171 -323
rect 191 -324 199 -323
rect 201 -324 304 -323
rect 324 -324 346 -323
rect 366 -324 374 -323
rect 135 -326 234 -325
rect 313 -326 374 -325
rect 184 -328 304 -327
rect 324 -328 500 -327
rect 149 -330 185 -329
rect 205 -330 318 -329
rect 369 -330 549 -329
rect 93 -332 206 -331
rect 233 -332 360 -331
rect 548 -332 598 -331
rect 93 -334 241 -333
rect 9 -345 661 -344
rect 709 -345 717 -344
rect 12 -347 66 -346
rect 68 -347 619 -346
rect 23 -349 129 -348
rect 142 -349 304 -348
rect 313 -349 367 -348
rect 467 -349 626 -348
rect 30 -351 80 -350
rect 89 -351 507 -350
rect 548 -351 619 -350
rect 37 -353 45 -352
rect 51 -353 482 -352
rect 506 -353 535 -352
rect 597 -353 633 -352
rect 37 -355 465 -354
rect 471 -355 661 -354
rect 44 -357 332 -356
rect 338 -357 444 -356
rect 450 -357 472 -356
rect 72 -359 101 -358
rect 117 -359 192 -358
rect 198 -359 248 -358
rect 282 -359 363 -358
rect 390 -359 535 -358
rect 75 -361 409 -360
rect 411 -361 626 -360
rect 79 -363 157 -362
rect 163 -363 213 -362
rect 226 -363 328 -362
rect 355 -363 654 -362
rect 86 -365 101 -364
rect 107 -365 164 -364
rect 177 -365 213 -364
rect 219 -365 227 -364
rect 233 -365 367 -364
rect 390 -365 416 -364
rect 443 -365 486 -364
rect 590 -365 654 -364
rect 86 -367 94 -366
rect 110 -367 220 -366
rect 233 -367 269 -366
rect 282 -367 342 -366
rect 359 -367 584 -366
rect 590 -367 612 -366
rect 58 -369 360 -368
rect 394 -369 416 -368
rect 450 -369 479 -368
rect 485 -369 514 -368
rect 583 -369 636 -368
rect 58 -371 157 -370
rect 201 -371 206 -370
rect 247 -371 255 -370
rect 268 -371 311 -370
rect 317 -371 381 -370
rect 457 -371 549 -370
rect 121 -373 192 -372
rect 254 -373 384 -372
rect 457 -373 521 -372
rect 121 -375 423 -374
rect 492 -375 514 -374
rect 128 -377 171 -376
rect 187 -377 206 -376
rect 296 -377 311 -376
rect 324 -377 675 -376
rect 114 -379 297 -378
rect 303 -379 346 -378
rect 352 -379 521 -378
rect 135 -381 178 -380
rect 334 -381 395 -380
rect 422 -381 528 -380
rect 135 -383 290 -382
rect 345 -383 374 -382
rect 380 -383 647 -382
rect 142 -385 150 -384
rect 170 -385 262 -384
rect 289 -385 430 -384
rect 492 -385 640 -384
rect 93 -387 150 -386
rect 261 -387 388 -386
rect 495 -387 528 -386
rect 562 -387 647 -386
rect 355 -389 612 -388
rect 373 -391 577 -390
rect 604 -391 640 -390
rect 541 -393 577 -392
rect 604 -393 668 -392
rect 243 -395 542 -394
rect 562 -395 570 -394
rect 324 -397 570 -396
rect 401 -399 668 -398
rect 401 -401 500 -400
rect 9 -412 97 -411
rect 100 -412 195 -411
rect 198 -412 244 -411
rect 268 -412 374 -411
rect 383 -412 528 -411
rect 562 -412 654 -411
rect 656 -412 661 -411
rect 716 -412 731 -411
rect 16 -414 80 -413
rect 93 -414 423 -413
rect 425 -414 577 -413
rect 597 -414 682 -413
rect 23 -416 83 -415
rect 114 -416 171 -415
rect 180 -416 640 -415
rect 30 -418 104 -417
rect 121 -418 577 -417
rect 583 -418 640 -417
rect 37 -420 111 -419
rect 156 -420 241 -419
rect 247 -420 269 -419
rect 282 -420 521 -419
rect 534 -420 563 -419
rect 569 -420 724 -419
rect 37 -422 52 -421
rect 58 -422 353 -421
rect 373 -422 423 -421
rect 432 -422 500 -421
rect 513 -422 570 -421
rect 604 -422 703 -421
rect 44 -424 94 -423
rect 100 -424 122 -423
rect 135 -424 241 -423
rect 303 -424 353 -423
rect 387 -424 454 -423
rect 464 -424 598 -423
rect 611 -424 689 -423
rect 44 -426 143 -425
rect 163 -426 339 -425
rect 390 -426 619 -425
rect 625 -426 675 -425
rect 58 -428 129 -427
rect 135 -428 206 -427
rect 219 -428 227 -427
rect 233 -428 283 -427
rect 296 -428 388 -427
rect 390 -428 528 -427
rect 541 -428 584 -427
rect 65 -430 108 -429
rect 149 -430 206 -429
rect 212 -430 234 -429
rect 313 -430 465 -429
rect 481 -430 633 -429
rect 68 -432 542 -431
rect 555 -432 605 -431
rect 72 -434 125 -433
rect 149 -434 286 -433
rect 324 -434 360 -433
rect 401 -434 535 -433
rect 72 -436 381 -435
rect 408 -436 647 -435
rect 86 -438 248 -437
rect 327 -438 549 -437
rect 590 -438 647 -437
rect 86 -440 255 -439
rect 331 -440 447 -439
rect 450 -440 514 -439
rect 170 -442 304 -441
rect 345 -442 381 -441
rect 411 -442 591 -441
rect 177 -444 213 -443
rect 254 -444 318 -443
rect 359 -444 419 -443
rect 436 -444 549 -443
rect 128 -446 178 -445
rect 184 -446 290 -445
rect 310 -446 346 -445
rect 366 -446 402 -445
rect 436 -446 626 -445
rect 184 -448 220 -447
rect 229 -448 318 -447
rect 439 -448 710 -447
rect 191 -450 297 -449
rect 443 -450 521 -449
rect 51 -452 192 -451
rect 198 -452 262 -451
rect 289 -452 395 -451
rect 492 -452 696 -451
rect 166 -454 262 -453
rect 394 -454 458 -453
rect 485 -454 493 -453
rect 502 -454 612 -453
rect 341 -456 458 -455
rect 506 -456 556 -455
rect 366 -458 486 -457
rect 471 -460 507 -459
rect 471 -462 668 -461
rect 478 -464 668 -463
rect 415 -466 479 -465
rect 58 -477 164 -476
rect 177 -477 605 -476
rect 639 -477 710 -476
rect 716 -477 731 -476
rect 75 -479 745 -478
rect 23 -481 76 -480
rect 79 -481 738 -480
rect 79 -483 136 -482
rect 145 -483 696 -482
rect 723 -483 780 -482
rect 93 -485 146 -484
rect 152 -485 206 -484
rect 219 -485 223 -484
rect 243 -485 346 -484
rect 359 -485 619 -484
rect 646 -485 724 -484
rect 37 -487 94 -486
rect 121 -487 192 -486
rect 219 -487 255 -486
rect 289 -487 451 -486
rect 555 -487 605 -486
rect 674 -487 717 -486
rect 121 -489 269 -488
rect 289 -489 332 -488
rect 345 -489 374 -488
rect 383 -489 416 -488
rect 422 -489 640 -488
rect 51 -491 332 -490
rect 352 -491 360 -490
rect 366 -491 549 -490
rect 555 -491 591 -490
rect 597 -491 661 -490
rect 16 -493 591 -492
rect 30 -495 52 -494
rect 124 -495 696 -494
rect 128 -497 269 -496
rect 390 -497 612 -496
rect 107 -499 129 -498
rect 135 -499 720 -498
rect 44 -501 108 -500
rect 149 -501 206 -500
rect 222 -501 255 -500
rect 394 -501 752 -500
rect 44 -503 115 -502
rect 180 -503 213 -502
rect 408 -503 437 -502
rect 439 -503 682 -502
rect 61 -505 115 -504
rect 187 -505 339 -504
rect 401 -505 409 -504
rect 411 -505 479 -504
rect 513 -505 549 -504
rect 562 -505 612 -504
rect 625 -505 682 -504
rect 65 -507 626 -506
rect 170 -509 563 -508
rect 576 -509 647 -508
rect 170 -511 283 -510
rect 303 -511 339 -510
rect 429 -511 654 -510
rect 191 -513 311 -512
rect 324 -513 402 -512
rect 432 -513 598 -512
rect 142 -515 311 -514
rect 317 -515 325 -514
rect 432 -515 668 -514
rect 212 -517 297 -516
rect 303 -517 731 -516
rect 226 -519 318 -518
rect 397 -519 668 -518
rect 226 -521 234 -520
rect 240 -521 297 -520
rect 443 -521 703 -520
rect 233 -523 353 -522
rect 387 -523 703 -522
rect 240 -525 374 -524
rect 443 -525 689 -524
rect 261 -527 388 -526
rect 478 -527 528 -526
rect 534 -527 577 -526
rect 583 -527 654 -526
rect 282 -529 370 -528
rect 453 -529 535 -528
rect 632 -529 689 -528
rect 9 -531 633 -530
rect 492 -533 584 -532
rect 446 -535 493 -534
rect 506 -535 528 -534
rect 261 -537 447 -536
rect 513 -537 542 -536
rect 320 -539 507 -538
rect 520 -539 675 -538
rect 499 -541 521 -540
rect 541 -541 570 -540
rect 464 -543 570 -542
rect 457 -545 465 -544
rect 485 -545 500 -544
rect 86 -547 458 -546
rect 471 -547 486 -546
rect 68 -549 472 -548
rect 26 -551 69 -550
rect 86 -551 164 -550
rect 16 -562 409 -561
rect 418 -562 724 -561
rect 779 -562 808 -561
rect 23 -564 55 -563
rect 58 -564 136 -563
rect 156 -564 178 -563
rect 187 -564 283 -563
rect 306 -564 325 -563
rect 355 -564 521 -563
rect 541 -564 545 -563
rect 23 -566 125 -565
rect 128 -566 157 -565
rect 166 -566 675 -565
rect 30 -568 97 -567
rect 100 -568 150 -567
rect 177 -568 188 -567
rect 205 -568 216 -567
rect 219 -568 318 -567
rect 366 -568 500 -567
rect 541 -568 577 -567
rect 33 -570 52 -569
rect 61 -570 626 -569
rect 44 -572 129 -571
rect 191 -572 318 -571
rect 369 -572 675 -571
rect 47 -574 654 -573
rect 51 -576 367 -575
rect 394 -576 647 -575
rect 65 -578 398 -577
rect 411 -578 500 -577
rect 544 -578 577 -577
rect 625 -578 689 -577
rect 65 -580 353 -579
rect 394 -580 752 -579
rect 72 -582 591 -581
rect 646 -582 696 -581
rect 72 -584 143 -583
rect 191 -584 199 -583
rect 212 -584 724 -583
rect 107 -586 185 -585
rect 212 -586 402 -585
rect 425 -586 535 -585
rect 590 -586 640 -585
rect 688 -586 731 -585
rect 114 -588 136 -587
rect 219 -588 311 -587
rect 338 -588 370 -587
rect 401 -588 416 -587
rect 429 -588 570 -587
rect 597 -588 696 -587
rect 730 -588 738 -587
rect 226 -590 521 -589
rect 569 -590 605 -589
rect 226 -592 262 -591
rect 275 -592 279 -591
rect 282 -592 297 -591
rect 310 -592 451 -591
rect 471 -592 738 -591
rect 233 -594 297 -593
rect 331 -594 416 -593
rect 429 -594 465 -593
rect 471 -594 493 -593
rect 604 -594 661 -593
rect 163 -596 661 -595
rect 233 -598 255 -597
rect 261 -598 388 -597
rect 432 -598 710 -597
rect 142 -600 710 -599
rect 184 -602 255 -601
rect 275 -602 654 -601
rect 236 -604 745 -603
rect 240 -606 248 -605
rect 289 -606 325 -605
rect 331 -606 374 -605
rect 387 -606 668 -605
rect 79 -608 241 -607
rect 247 -608 269 -607
rect 303 -608 374 -607
rect 390 -608 668 -607
rect 79 -610 171 -609
rect 198 -610 290 -609
rect 303 -610 346 -609
rect 348 -610 598 -609
rect 86 -612 171 -611
rect 268 -612 293 -611
rect 338 -612 458 -611
rect 464 -612 556 -611
rect 86 -614 104 -613
rect 320 -614 458 -613
rect 478 -614 535 -613
rect 555 -614 717 -613
rect 93 -616 346 -615
rect 352 -616 619 -615
rect 93 -618 206 -617
rect 383 -618 619 -617
rect 443 -620 612 -619
rect 446 -622 703 -621
rect 446 -624 640 -623
rect 450 -626 549 -625
rect 485 -628 612 -627
rect 485 -630 507 -629
rect 513 -630 703 -629
rect 478 -632 514 -631
rect 516 -632 717 -631
rect 506 -634 528 -633
rect 548 -634 584 -633
rect 380 -636 528 -635
rect 583 -636 633 -635
rect 359 -638 381 -637
rect 632 -638 682 -637
rect 359 -640 437 -639
rect 75 -642 437 -641
rect 425 -644 682 -643
rect 58 -655 97 -654
rect 100 -655 115 -654
rect 117 -655 157 -654
rect 166 -655 178 -654
rect 184 -655 241 -654
rect 254 -655 346 -654
rect 348 -655 451 -654
rect 474 -655 766 -654
rect 807 -655 829 -654
rect 9 -657 115 -656
rect 117 -657 199 -656
rect 212 -657 255 -656
rect 261 -657 279 -656
rect 282 -657 290 -656
rect 352 -657 416 -656
rect 418 -657 514 -656
rect 555 -657 773 -656
rect 16 -659 353 -658
rect 366 -659 535 -658
rect 597 -659 825 -658
rect 16 -661 73 -660
rect 86 -661 122 -660
rect 124 -661 433 -660
rect 443 -661 556 -660
rect 660 -661 696 -660
rect 709 -661 787 -660
rect 51 -663 101 -662
rect 107 -663 584 -662
rect 646 -663 696 -662
rect 716 -663 794 -662
rect 58 -665 801 -664
rect 65 -667 150 -666
rect 152 -667 244 -666
rect 261 -667 290 -666
rect 380 -667 388 -666
rect 408 -667 612 -666
rect 667 -667 710 -666
rect 730 -667 759 -666
rect 23 -669 66 -668
rect 86 -669 311 -668
rect 411 -669 808 -668
rect 23 -671 258 -670
rect 303 -671 381 -670
rect 422 -671 703 -670
rect 30 -673 412 -672
rect 429 -673 493 -672
rect 590 -673 612 -672
rect 618 -673 703 -672
rect 37 -675 409 -674
rect 443 -675 479 -674
rect 548 -675 591 -674
rect 604 -675 619 -674
rect 653 -675 668 -674
rect 674 -675 752 -674
rect 44 -677 654 -676
rect 681 -677 717 -676
rect 44 -679 94 -678
rect 107 -679 164 -678
rect 177 -679 402 -678
rect 439 -679 549 -678
rect 576 -679 605 -678
rect 681 -679 724 -678
rect 79 -681 304 -680
rect 310 -681 339 -680
rect 394 -681 423 -680
rect 457 -681 647 -680
rect 688 -681 780 -680
rect 79 -683 391 -682
rect 397 -683 577 -682
rect 632 -683 724 -682
rect 121 -685 528 -684
rect 625 -685 633 -684
rect 639 -685 689 -684
rect 128 -687 269 -686
rect 282 -687 395 -686
rect 467 -687 479 -686
rect 499 -687 640 -686
rect 131 -689 542 -688
rect 569 -689 626 -688
rect 135 -691 213 -690
rect 219 -691 339 -690
rect 359 -691 458 -690
rect 471 -691 535 -690
rect 124 -693 220 -692
rect 226 -693 269 -692
rect 292 -693 675 -692
rect 110 -695 227 -694
rect 236 -695 745 -694
rect 135 -697 146 -696
rect 156 -697 318 -696
rect 331 -697 402 -696
rect 436 -697 500 -696
rect 506 -697 542 -696
rect 142 -699 486 -698
rect 506 -699 738 -698
rect 47 -701 143 -700
rect 163 -701 563 -700
rect 166 -703 563 -702
rect 184 -705 276 -704
rect 296 -705 360 -704
rect 369 -705 738 -704
rect 173 -707 297 -706
rect 317 -707 815 -706
rect 198 -709 248 -708
rect 324 -709 370 -708
rect 446 -709 486 -708
rect 205 -711 584 -710
rect 170 -713 206 -712
rect 233 -713 276 -712
rect 324 -713 374 -712
rect 233 -715 521 -714
rect 240 -717 731 -716
rect 247 -719 430 -718
rect 464 -719 521 -718
rect 331 -721 528 -720
rect 334 -723 570 -722
rect 373 -725 437 -724
rect 40 -736 122 -735
rect 124 -736 731 -735
rect 817 -736 829 -735
rect 44 -738 69 -737
rect 72 -738 213 -737
rect 236 -738 465 -737
rect 467 -738 794 -737
rect 47 -740 66 -739
rect 72 -740 307 -739
rect 324 -740 465 -739
rect 474 -740 780 -739
rect 51 -742 584 -741
rect 597 -742 633 -741
rect 639 -742 815 -741
rect 58 -744 654 -743
rect 681 -744 780 -743
rect 58 -746 339 -745
rect 341 -746 808 -745
rect 75 -748 654 -747
rect 660 -748 682 -747
rect 96 -750 661 -749
rect 117 -752 703 -751
rect 142 -754 213 -753
rect 240 -754 825 -753
rect 79 -756 241 -755
rect 254 -756 269 -755
rect 289 -756 766 -755
rect 86 -758 269 -757
rect 282 -758 290 -757
rect 292 -758 486 -757
rect 506 -758 731 -757
rect 86 -760 234 -759
rect 275 -760 283 -759
rect 310 -760 507 -759
rect 583 -760 689 -759
rect 37 -762 311 -761
rect 324 -762 346 -761
rect 348 -762 794 -761
rect 37 -764 801 -763
rect 107 -766 234 -765
rect 331 -766 353 -765
rect 366 -766 703 -765
rect 107 -768 472 -767
rect 548 -768 689 -767
rect 82 -770 549 -769
rect 590 -770 766 -769
rect 135 -772 276 -771
rect 296 -772 332 -771
rect 352 -772 370 -771
rect 394 -772 493 -771
rect 600 -772 752 -771
rect 135 -774 367 -773
rect 387 -774 395 -773
rect 408 -774 444 -773
rect 450 -774 675 -773
rect 709 -774 752 -773
rect 142 -776 185 -775
rect 226 -776 346 -775
rect 408 -776 416 -775
rect 429 -776 521 -775
rect 632 -776 668 -775
rect 159 -778 773 -777
rect 163 -780 402 -779
rect 411 -780 626 -779
rect 639 -780 738 -779
rect 170 -782 206 -781
rect 296 -782 440 -781
rect 446 -782 675 -781
rect 198 -784 227 -783
rect 380 -784 416 -783
rect 436 -784 724 -783
rect 16 -786 724 -785
rect 198 -788 374 -787
rect 380 -788 745 -787
rect 205 -790 248 -789
rect 359 -790 374 -789
rect 404 -790 738 -789
rect 23 -792 248 -791
rect 338 -792 360 -791
rect 436 -792 745 -791
rect 23 -794 157 -793
rect 457 -794 486 -793
rect 492 -794 542 -793
rect 604 -794 668 -793
rect 93 -796 157 -795
rect 422 -796 458 -795
rect 471 -796 514 -795
rect 520 -796 577 -795
rect 625 -796 696 -795
rect 93 -798 262 -797
rect 453 -798 514 -797
rect 534 -798 542 -797
rect 562 -798 577 -797
rect 618 -798 696 -797
rect 16 -800 563 -799
rect 569 -800 605 -799
rect 646 -800 710 -799
rect 149 -802 423 -801
rect 499 -802 773 -801
rect 114 -804 150 -803
rect 261 -804 388 -803
rect 478 -804 500 -803
rect 527 -804 535 -803
rect 555 -804 570 -803
rect 646 -804 822 -803
rect 177 -806 528 -805
rect 555 -806 787 -805
rect 128 -808 178 -807
rect 219 -808 479 -807
rect 758 -808 787 -807
rect 30 -810 129 -809
rect 219 -810 318 -809
rect 716 -810 759 -809
rect 30 -812 188 -811
rect 271 -812 619 -811
rect 303 -814 318 -813
rect 390 -814 717 -813
rect 9 -825 94 -824
rect 96 -825 241 -824
rect 303 -825 773 -824
rect 23 -827 52 -826
rect 54 -827 363 -826
rect 369 -827 710 -826
rect 37 -829 724 -828
rect 37 -831 286 -830
rect 331 -831 745 -830
rect 26 -833 332 -832
rect 348 -833 528 -832
rect 530 -833 780 -832
rect 51 -835 213 -834
rect 352 -835 731 -834
rect 58 -837 241 -836
rect 359 -837 384 -836
rect 390 -837 766 -836
rect 58 -839 192 -838
rect 212 -839 255 -838
rect 373 -839 388 -838
rect 404 -839 570 -838
rect 590 -839 689 -838
rect 709 -839 759 -838
rect 30 -841 192 -840
rect 257 -841 374 -840
rect 380 -841 577 -840
rect 632 -841 636 -840
rect 681 -841 759 -840
rect 30 -843 101 -842
rect 128 -843 185 -842
rect 187 -843 283 -842
rect 306 -843 689 -842
rect 65 -845 654 -844
rect 65 -847 69 -846
rect 72 -847 108 -846
rect 114 -847 129 -846
rect 145 -847 738 -846
rect 16 -849 115 -848
rect 149 -849 318 -848
rect 324 -849 388 -848
rect 394 -849 405 -848
rect 411 -849 703 -848
rect 716 -849 738 -848
rect 44 -851 703 -850
rect 44 -853 248 -852
rect 310 -853 325 -852
rect 338 -853 577 -852
rect 611 -853 682 -852
rect 72 -855 199 -854
rect 219 -855 311 -854
rect 394 -855 409 -854
rect 422 -855 654 -854
rect 82 -857 507 -856
rect 537 -857 696 -856
rect 86 -859 199 -858
rect 226 -859 248 -858
rect 422 -859 563 -858
rect 569 -859 668 -858
rect 86 -861 122 -860
rect 149 -861 262 -860
rect 429 -861 486 -860
rect 555 -861 794 -860
rect 93 -863 143 -862
rect 152 -863 276 -862
rect 299 -863 430 -862
rect 436 -863 521 -862
rect 555 -863 619 -862
rect 632 -863 640 -862
rect 667 -863 752 -862
rect 107 -865 360 -864
rect 436 -865 479 -864
rect 485 -865 549 -864
rect 562 -865 661 -864
rect 121 -867 171 -866
rect 173 -867 297 -866
rect 306 -867 479 -866
rect 513 -867 661 -866
rect 142 -869 220 -868
rect 275 -869 444 -868
rect 450 -869 619 -868
rect 156 -871 160 -870
rect 163 -871 318 -870
rect 345 -871 521 -870
rect 156 -873 206 -872
rect 345 -873 416 -872
rect 443 -873 500 -872
rect 513 -873 605 -872
rect 117 -875 416 -874
rect 453 -875 493 -874
rect 597 -875 605 -874
rect 635 -875 640 -874
rect 163 -877 269 -876
rect 453 -877 787 -876
rect 170 -879 342 -878
rect 457 -879 500 -878
rect 135 -881 458 -880
rect 492 -881 542 -880
rect 135 -883 227 -882
rect 268 -883 290 -882
rect 541 -883 647 -882
rect 79 -885 290 -884
rect 583 -885 647 -884
rect 177 -887 353 -886
rect 583 -887 675 -886
rect 177 -889 234 -888
rect 674 -889 696 -888
rect 180 -891 262 -890
rect 233 -893 367 -892
rect 366 -895 465 -894
rect 464 -897 535 -896
rect 534 -899 598 -898
rect 2 -910 101 -909
rect 103 -910 234 -909
rect 240 -910 307 -909
rect 338 -910 353 -909
rect 359 -910 538 -909
rect 548 -910 563 -909
rect 576 -910 591 -909
rect 607 -910 682 -909
rect 695 -910 759 -909
rect 23 -912 500 -911
rect 509 -912 633 -911
rect 737 -912 752 -911
rect 26 -914 171 -913
rect 205 -914 255 -913
rect 257 -914 682 -913
rect 30 -916 146 -915
rect 205 -916 398 -915
rect 404 -916 647 -915
rect 30 -918 188 -917
rect 212 -918 290 -917
rect 296 -918 311 -917
rect 383 -918 395 -917
rect 408 -918 612 -917
rect 618 -918 633 -917
rect 37 -920 48 -919
rect 54 -920 689 -919
rect 40 -922 703 -921
rect 65 -924 146 -923
rect 156 -924 213 -923
rect 229 -924 591 -923
rect 597 -924 696 -923
rect 65 -926 556 -925
rect 576 -926 605 -925
rect 621 -926 710 -925
rect 72 -928 255 -927
rect 275 -928 703 -927
rect 72 -930 367 -929
rect 387 -930 451 -929
rect 478 -930 710 -929
rect 79 -932 174 -931
rect 219 -932 367 -931
rect 394 -932 661 -931
rect 688 -932 727 -931
rect 61 -934 80 -933
rect 86 -934 251 -933
rect 275 -934 346 -933
rect 362 -934 661 -933
rect 93 -936 153 -935
rect 156 -936 164 -935
rect 226 -936 388 -935
rect 415 -936 717 -935
rect 93 -938 199 -937
rect 233 -938 300 -937
rect 303 -938 363 -937
rect 450 -938 472 -937
rect 478 -938 528 -937
rect 534 -938 570 -937
rect 625 -938 629 -937
rect 44 -940 199 -939
rect 240 -940 269 -939
rect 278 -940 325 -939
rect 499 -940 647 -939
rect 44 -942 570 -941
rect 625 -942 640 -941
rect 107 -944 503 -943
rect 513 -944 528 -943
rect 555 -944 675 -943
rect 107 -946 353 -945
rect 513 -946 584 -945
rect 628 -946 640 -945
rect 114 -948 129 -947
rect 135 -948 472 -947
rect 520 -948 675 -947
rect 16 -950 129 -949
rect 163 -950 181 -949
rect 261 -950 346 -949
rect 520 -950 542 -949
rect 562 -950 605 -949
rect 16 -952 192 -951
rect 261 -952 412 -951
rect 100 -954 136 -953
rect 149 -954 192 -953
rect 282 -954 493 -953
rect 117 -956 248 -955
rect 285 -956 423 -955
rect 485 -956 493 -955
rect 121 -958 220 -957
rect 310 -958 654 -957
rect 58 -960 122 -959
rect 142 -960 423 -959
rect 653 -960 668 -959
rect 9 -962 59 -961
rect 149 -962 416 -961
rect 180 -964 458 -963
rect 324 -966 507 -965
rect 313 -968 507 -967
rect 331 -970 584 -969
rect 51 -972 332 -971
rect 373 -972 542 -971
rect 184 -974 374 -973
rect 401 -974 668 -973
rect 184 -976 269 -975
rect 401 -976 412 -975
rect 457 -976 465 -975
rect 429 -978 465 -977
rect 429 -980 444 -979
rect 380 -982 444 -981
rect 9 -993 185 -992
rect 187 -993 255 -992
rect 275 -993 356 -992
rect 404 -993 437 -992
rect 443 -993 451 -992
rect 464 -993 486 -992
rect 499 -993 507 -992
rect 520 -993 524 -992
rect 527 -993 731 -992
rect 751 -993 759 -992
rect 26 -995 66 -994
rect 79 -995 87 -994
rect 89 -995 612 -994
rect 618 -995 633 -994
rect 716 -995 724 -994
rect 30 -997 363 -996
rect 425 -997 528 -996
rect 604 -997 622 -996
rect 625 -997 633 -996
rect 709 -997 717 -996
rect 37 -999 143 -998
rect 149 -999 395 -998
rect 436 -999 458 -998
rect 464 -999 493 -998
rect 502 -999 577 -998
rect 695 -999 710 -998
rect 37 -1001 73 -1000
rect 79 -1001 430 -1000
rect 457 -1001 472 -1000
rect 478 -1001 507 -1000
rect 520 -1001 563 -1000
rect 695 -1001 703 -1000
rect 44 -1003 682 -1002
rect 688 -1003 703 -1002
rect 47 -1005 199 -1004
rect 205 -1005 447 -1004
rect 485 -1005 608 -1004
rect 674 -1005 689 -1004
rect 54 -1007 570 -1006
rect 660 -1007 675 -1006
rect 58 -1009 416 -1008
rect 488 -1009 577 -1008
rect 660 -1009 668 -1008
rect 68 -1011 479 -1010
rect 523 -1011 563 -1010
rect 569 -1011 584 -1010
rect 86 -1013 332 -1012
rect 352 -1013 472 -1012
rect 555 -1013 682 -1012
rect 93 -1015 185 -1014
rect 191 -1015 199 -1014
rect 205 -1015 346 -1014
rect 366 -1015 584 -1014
rect 2 -1017 346 -1016
rect 366 -1017 381 -1016
rect 383 -1017 430 -1016
rect 534 -1017 556 -1016
rect 93 -1019 101 -1018
rect 107 -1019 647 -1018
rect 16 -1021 108 -1020
rect 114 -1021 290 -1020
rect 292 -1021 598 -1020
rect 16 -1023 171 -1022
rect 180 -1023 374 -1022
rect 394 -1023 542 -1022
rect 100 -1025 213 -1024
rect 219 -1025 227 -1024
rect 240 -1025 314 -1024
rect 317 -1025 370 -1024
rect 373 -1025 514 -1024
rect 534 -1025 591 -1024
rect 23 -1027 591 -1026
rect 75 -1029 241 -1028
rect 247 -1029 262 -1028
rect 268 -1029 612 -1028
rect 117 -1031 220 -1030
rect 226 -1031 325 -1030
rect 331 -1031 360 -1030
rect 142 -1033 402 -1032
rect 156 -1035 171 -1034
rect 177 -1035 542 -1034
rect 128 -1037 178 -1036
rect 212 -1037 311 -1036
rect 317 -1037 339 -1036
rect 401 -1037 668 -1036
rect 103 -1039 129 -1038
rect 135 -1039 157 -1038
rect 163 -1039 192 -1038
rect 250 -1039 647 -1038
rect 121 -1041 164 -1040
rect 254 -1041 423 -1040
rect 30 -1043 122 -1042
rect 135 -1043 150 -1042
rect 261 -1043 297 -1042
rect 306 -1043 339 -1042
rect 422 -1043 514 -1042
rect 233 -1045 297 -1044
rect 310 -1045 626 -1044
rect 233 -1047 451 -1046
rect 268 -1049 409 -1048
rect 275 -1051 304 -1050
rect 320 -1051 388 -1050
rect 282 -1053 412 -1052
rect 303 -1055 493 -1054
rect 324 -1057 353 -1056
rect 387 -1057 398 -1056
rect 16 -1068 360 -1067
rect 362 -1068 696 -1067
rect 730 -1068 738 -1067
rect 751 -1068 755 -1067
rect 16 -1070 262 -1069
rect 268 -1070 290 -1069
rect 306 -1070 682 -1069
rect 754 -1070 794 -1069
rect 26 -1072 87 -1071
rect 89 -1072 174 -1071
rect 177 -1072 262 -1071
rect 310 -1072 346 -1071
rect 369 -1072 549 -1071
rect 597 -1072 731 -1071
rect 9 -1074 87 -1073
rect 107 -1074 304 -1073
rect 310 -1074 325 -1073
rect 327 -1074 374 -1073
rect 383 -1074 507 -1073
rect 509 -1074 682 -1073
rect 9 -1076 122 -1075
rect 156 -1076 188 -1075
rect 205 -1076 377 -1075
rect 394 -1076 440 -1075
rect 464 -1076 787 -1075
rect 30 -1078 472 -1077
rect 474 -1078 577 -1077
rect 604 -1078 654 -1077
rect 660 -1078 696 -1077
rect 37 -1080 139 -1079
rect 156 -1080 167 -1079
rect 170 -1080 272 -1079
rect 331 -1080 598 -1079
rect 632 -1080 654 -1079
rect 667 -1080 780 -1079
rect 44 -1082 220 -1081
rect 247 -1082 416 -1081
rect 418 -1082 724 -1081
rect 47 -1084 66 -1083
rect 72 -1084 136 -1083
rect 138 -1084 584 -1083
rect 625 -1084 668 -1083
rect 709 -1084 724 -1083
rect 23 -1086 66 -1085
rect 100 -1086 188 -1085
rect 198 -1086 220 -1085
rect 250 -1086 276 -1085
rect 345 -1086 426 -1085
rect 450 -1086 626 -1085
rect 632 -1086 675 -1085
rect 688 -1086 710 -1085
rect 58 -1088 108 -1087
rect 114 -1088 192 -1087
rect 208 -1088 255 -1087
rect 275 -1088 339 -1087
rect 380 -1088 605 -1087
rect 639 -1088 661 -1087
rect 58 -1090 143 -1089
rect 163 -1090 332 -1089
rect 380 -1090 741 -1089
rect 114 -1092 213 -1091
rect 387 -1092 416 -1091
rect 425 -1092 717 -1091
rect 79 -1094 388 -1093
rect 397 -1094 584 -1093
rect 611 -1094 640 -1093
rect 646 -1094 675 -1093
rect 117 -1096 297 -1095
rect 401 -1096 409 -1095
rect 436 -1096 451 -1095
rect 457 -1096 465 -1095
rect 471 -1096 717 -1095
rect 51 -1098 458 -1097
rect 499 -1098 815 -1097
rect 51 -1100 206 -1099
rect 212 -1100 318 -1099
rect 436 -1100 563 -1099
rect 618 -1100 647 -1099
rect 37 -1102 318 -1101
rect 513 -1102 549 -1101
rect 562 -1102 570 -1101
rect 103 -1104 500 -1103
rect 534 -1104 577 -1103
rect 121 -1106 423 -1105
rect 527 -1106 535 -1105
rect 128 -1108 143 -1107
rect 163 -1108 479 -1107
rect 527 -1108 556 -1107
rect 128 -1110 150 -1109
rect 177 -1110 283 -1109
rect 289 -1110 570 -1109
rect 79 -1112 150 -1111
rect 180 -1112 325 -1111
rect 429 -1112 479 -1111
rect 555 -1112 591 -1111
rect 184 -1114 199 -1113
rect 240 -1114 297 -1113
rect 366 -1114 591 -1113
rect 184 -1116 234 -1115
rect 240 -1116 248 -1115
rect 282 -1116 339 -1115
rect 366 -1116 514 -1115
rect 191 -1118 304 -1117
rect 429 -1118 444 -1117
rect 194 -1120 255 -1119
rect 443 -1120 493 -1119
rect 233 -1122 409 -1121
rect 485 -1122 493 -1121
rect 320 -1124 486 -1123
rect 9 -1135 328 -1134
rect 348 -1135 507 -1134
rect 509 -1135 703 -1134
rect 716 -1135 773 -1134
rect 793 -1135 801 -1134
rect 9 -1137 283 -1136
rect 310 -1137 321 -1136
rect 355 -1137 374 -1136
rect 422 -1137 594 -1136
rect 646 -1137 689 -1136
rect 740 -1137 794 -1136
rect 23 -1139 339 -1138
rect 366 -1139 549 -1138
rect 555 -1139 766 -1138
rect 26 -1141 640 -1140
rect 744 -1141 780 -1140
rect 30 -1143 598 -1142
rect 723 -1143 780 -1142
rect 37 -1145 188 -1144
rect 194 -1145 332 -1144
rect 341 -1145 598 -1144
rect 674 -1145 724 -1144
rect 751 -1145 759 -1144
rect 44 -1147 339 -1146
rect 373 -1147 514 -1146
rect 520 -1147 703 -1146
rect 44 -1149 430 -1148
rect 432 -1149 717 -1148
rect 54 -1151 458 -1150
rect 467 -1151 493 -1150
rect 534 -1151 612 -1150
rect 632 -1151 752 -1150
rect 72 -1153 248 -1152
rect 254 -1153 311 -1152
rect 324 -1153 367 -1152
rect 394 -1153 675 -1152
rect 695 -1153 759 -1152
rect 79 -1155 325 -1154
rect 331 -1155 381 -1154
rect 397 -1155 556 -1154
rect 562 -1155 633 -1154
rect 79 -1157 143 -1156
rect 145 -1157 209 -1156
rect 212 -1157 237 -1156
rect 247 -1157 258 -1156
rect 275 -1157 437 -1156
rect 443 -1157 563 -1156
rect 569 -1157 748 -1156
rect 16 -1159 276 -1158
rect 292 -1159 381 -1158
rect 401 -1159 493 -1158
rect 541 -1159 619 -1158
rect 16 -1161 164 -1160
rect 166 -1161 181 -1160
rect 187 -1161 458 -1160
rect 474 -1161 528 -1160
rect 548 -1161 787 -1160
rect 100 -1163 514 -1162
rect 569 -1163 815 -1162
rect 93 -1165 101 -1164
rect 114 -1165 682 -1164
rect 730 -1165 787 -1164
rect 93 -1167 391 -1166
rect 408 -1167 535 -1166
rect 576 -1167 640 -1166
rect 653 -1167 731 -1166
rect 117 -1169 283 -1168
rect 352 -1169 696 -1168
rect 117 -1171 192 -1170
rect 198 -1171 290 -1170
rect 296 -1171 353 -1170
rect 359 -1171 444 -1170
rect 450 -1171 521 -1170
rect 590 -1171 647 -1170
rect 121 -1173 150 -1172
rect 152 -1173 584 -1172
rect 625 -1173 682 -1172
rect 121 -1175 129 -1174
rect 135 -1175 584 -1174
rect 625 -1175 661 -1174
rect 51 -1177 129 -1176
rect 138 -1177 318 -1176
rect 429 -1177 472 -1176
rect 485 -1177 654 -1176
rect 33 -1179 486 -1178
rect 499 -1179 577 -1178
rect 51 -1181 738 -1180
rect 58 -1183 136 -1182
rect 177 -1183 370 -1182
rect 415 -1183 500 -1182
rect 58 -1185 69 -1184
rect 198 -1185 262 -1184
rect 296 -1185 426 -1184
rect 450 -1185 479 -1184
rect 65 -1187 416 -1186
rect 464 -1187 528 -1186
rect 65 -1189 73 -1188
rect 205 -1189 395 -1188
rect 471 -1189 605 -1188
rect 212 -1191 241 -1190
rect 250 -1191 605 -1190
rect 226 -1193 234 -1192
rect 240 -1193 405 -1192
rect 219 -1195 227 -1194
rect 261 -1195 269 -1194
rect 303 -1195 360 -1194
rect 369 -1195 388 -1194
rect 40 -1197 220 -1196
rect 268 -1197 412 -1196
rect 303 -1199 346 -1198
rect 345 -1201 668 -1200
rect 667 -1203 710 -1202
rect 478 -1205 710 -1204
rect 2 -1216 136 -1215
rect 184 -1216 199 -1215
rect 254 -1216 311 -1215
rect 317 -1216 444 -1215
rect 471 -1216 507 -1215
rect 541 -1216 647 -1215
rect 649 -1216 787 -1215
rect 789 -1216 801 -1215
rect 9 -1218 349 -1217
rect 362 -1218 598 -1217
rect 660 -1218 787 -1217
rect 9 -1220 31 -1219
rect 33 -1220 664 -1219
rect 667 -1220 738 -1219
rect 16 -1222 90 -1221
rect 128 -1222 395 -1221
rect 397 -1222 521 -1221
rect 593 -1222 731 -1221
rect 16 -1224 146 -1223
rect 198 -1224 381 -1223
rect 387 -1224 535 -1223
rect 681 -1224 731 -1223
rect 30 -1226 188 -1225
rect 254 -1226 328 -1225
rect 345 -1226 486 -1225
rect 506 -1226 612 -1225
rect 37 -1228 269 -1227
rect 278 -1228 591 -1227
rect 23 -1230 269 -1229
rect 282 -1230 346 -1229
rect 366 -1230 500 -1229
rect 520 -1230 577 -1229
rect 23 -1232 220 -1231
rect 247 -1232 500 -1231
rect 555 -1232 682 -1231
rect 51 -1234 59 -1233
rect 68 -1234 73 -1233
rect 75 -1234 437 -1233
rect 443 -1234 493 -1233
rect 555 -1234 654 -1233
rect 51 -1236 122 -1235
rect 128 -1236 339 -1235
rect 373 -1236 542 -1235
rect 576 -1236 605 -1235
rect 653 -1236 689 -1235
rect 54 -1238 493 -1237
rect 688 -1238 759 -1237
rect 58 -1240 241 -1239
rect 247 -1240 290 -1239
rect 317 -1240 423 -1239
rect 464 -1240 598 -1239
rect 758 -1240 780 -1239
rect 79 -1242 143 -1241
rect 145 -1242 192 -1241
rect 212 -1242 220 -1241
rect 240 -1242 353 -1241
rect 373 -1242 430 -1241
rect 464 -1242 514 -1241
rect 79 -1244 332 -1243
rect 334 -1244 605 -1243
rect 86 -1246 360 -1245
rect 390 -1246 633 -1245
rect 93 -1248 122 -1247
rect 135 -1248 206 -1247
rect 212 -1248 416 -1247
rect 422 -1248 451 -1247
rect 478 -1248 752 -1247
rect 93 -1250 178 -1249
rect 184 -1250 437 -1249
rect 450 -1250 668 -1249
rect 44 -1252 178 -1251
rect 191 -1252 304 -1251
rect 324 -1252 724 -1251
rect 44 -1254 73 -1253
rect 107 -1254 290 -1253
rect 324 -1254 458 -1253
rect 478 -1254 528 -1253
rect 632 -1254 780 -1253
rect 107 -1256 171 -1255
rect 205 -1256 227 -1255
rect 282 -1256 342 -1255
rect 401 -1256 549 -1255
rect 723 -1256 745 -1255
rect 65 -1258 171 -1257
rect 341 -1258 563 -1257
rect 744 -1258 773 -1257
rect 114 -1260 752 -1259
rect 772 -1260 794 -1259
rect 166 -1262 381 -1261
rect 401 -1262 766 -1261
rect 310 -1264 563 -1263
rect 404 -1266 612 -1265
rect 404 -1268 535 -1267
rect 548 -1268 619 -1267
rect 411 -1270 640 -1269
rect 411 -1272 703 -1271
rect 429 -1274 584 -1273
rect 639 -1274 696 -1273
rect 702 -1274 717 -1273
rect 457 -1276 486 -1275
rect 513 -1276 573 -1275
rect 646 -1276 717 -1275
rect 474 -1278 584 -1277
rect 695 -1278 710 -1277
rect 303 -1280 710 -1279
rect 481 -1282 783 -1281
rect 527 -1284 675 -1283
rect 569 -1286 619 -1285
rect 625 -1286 675 -1285
rect 275 -1288 626 -1287
rect 233 -1290 276 -1289
rect 233 -1292 262 -1291
rect 261 -1294 297 -1293
rect 296 -1296 409 -1295
rect 408 -1298 416 -1297
rect 2 -1309 349 -1308
rect 355 -1309 752 -1308
rect 782 -1309 801 -1308
rect 9 -1311 181 -1310
rect 191 -1311 314 -1310
rect 359 -1311 500 -1310
rect 516 -1311 675 -1310
rect 709 -1311 769 -1310
rect 9 -1313 321 -1312
rect 362 -1313 563 -1312
rect 565 -1313 706 -1312
rect 730 -1313 780 -1312
rect 30 -1315 34 -1314
rect 40 -1315 45 -1314
rect 65 -1315 528 -1314
rect 537 -1315 738 -1314
rect 30 -1317 129 -1316
rect 149 -1317 188 -1316
rect 198 -1317 353 -1316
rect 404 -1317 493 -1316
rect 527 -1317 556 -1316
rect 562 -1317 696 -1316
rect 44 -1319 465 -1318
rect 492 -1319 584 -1318
rect 590 -1319 710 -1318
rect 51 -1321 188 -1320
rect 198 -1321 206 -1320
rect 215 -1321 360 -1320
rect 408 -1321 703 -1320
rect 51 -1323 146 -1322
rect 149 -1323 157 -1322
rect 163 -1323 290 -1322
rect 296 -1323 367 -1322
rect 457 -1323 521 -1322
rect 534 -1323 591 -1322
rect 639 -1323 692 -1322
rect 702 -1323 724 -1322
rect 68 -1325 94 -1324
rect 114 -1325 202 -1324
rect 219 -1325 230 -1324
rect 268 -1325 290 -1324
rect 310 -1325 395 -1324
rect 429 -1325 535 -1324
rect 541 -1325 556 -1324
rect 572 -1325 759 -1324
rect 58 -1327 220 -1326
rect 226 -1327 248 -1326
rect 275 -1327 409 -1326
rect 457 -1327 479 -1326
rect 485 -1327 521 -1326
rect 541 -1327 549 -1326
rect 576 -1327 584 -1326
rect 639 -1327 654 -1326
rect 688 -1327 696 -1326
rect 744 -1327 759 -1326
rect 23 -1329 276 -1328
rect 296 -1329 577 -1328
rect 653 -1329 668 -1328
rect 23 -1331 416 -1330
rect 425 -1331 668 -1330
rect 65 -1333 94 -1332
rect 114 -1333 283 -1332
rect 345 -1333 416 -1332
rect 471 -1333 486 -1332
rect 506 -1333 549 -1332
rect 72 -1335 647 -1334
rect 75 -1337 430 -1336
rect 506 -1337 514 -1336
rect 82 -1339 108 -1338
rect 117 -1339 500 -1338
rect 107 -1341 185 -1340
rect 191 -1341 689 -1340
rect 117 -1343 143 -1342
rect 156 -1343 171 -1342
rect 177 -1343 248 -1342
rect 268 -1343 479 -1342
rect 16 -1345 171 -1344
rect 184 -1345 339 -1344
rect 352 -1345 374 -1344
rect 380 -1345 395 -1344
rect 464 -1345 514 -1344
rect 37 -1347 143 -1346
rect 163 -1347 437 -1346
rect 58 -1349 178 -1348
rect 233 -1349 283 -1348
rect 366 -1349 447 -1348
rect 86 -1351 234 -1350
rect 373 -1351 451 -1350
rect 121 -1353 129 -1352
rect 135 -1353 206 -1352
rect 380 -1353 598 -1352
rect 121 -1355 255 -1354
rect 387 -1355 472 -1354
rect 597 -1355 612 -1354
rect 135 -1357 335 -1356
rect 387 -1357 402 -1356
rect 422 -1357 437 -1356
rect 443 -1357 451 -1356
rect 611 -1357 626 -1356
rect 166 -1359 482 -1358
rect 254 -1361 318 -1360
rect 401 -1361 675 -1360
rect 212 -1363 318 -1362
rect 443 -1363 619 -1362
rect 33 -1365 213 -1364
rect 261 -1365 335 -1364
rect 618 -1365 661 -1364
rect 79 -1367 262 -1366
rect 303 -1367 423 -1366
rect 660 -1367 682 -1366
rect 79 -1369 605 -1368
rect 681 -1369 717 -1368
rect 303 -1371 325 -1370
rect 331 -1371 605 -1370
rect 240 -1373 325 -1372
rect 240 -1375 412 -1374
rect 9 -1386 143 -1385
rect 149 -1386 164 -1385
rect 170 -1386 213 -1385
rect 271 -1386 325 -1385
rect 338 -1386 346 -1385
rect 383 -1386 745 -1385
rect 758 -1386 783 -1385
rect 786 -1386 829 -1385
rect 16 -1388 181 -1387
rect 275 -1388 381 -1387
rect 411 -1388 738 -1387
rect 779 -1388 808 -1387
rect 37 -1390 136 -1389
rect 149 -1390 279 -1389
rect 296 -1390 430 -1389
rect 443 -1390 654 -1389
rect 674 -1390 731 -1389
rect 789 -1390 801 -1389
rect 44 -1392 216 -1391
rect 247 -1392 297 -1391
rect 310 -1392 332 -1391
rect 338 -1392 409 -1391
rect 443 -1392 510 -1391
rect 534 -1392 689 -1391
rect 695 -1392 773 -1391
rect 796 -1392 804 -1391
rect 44 -1394 108 -1393
rect 121 -1394 143 -1393
rect 156 -1394 171 -1393
rect 177 -1394 423 -1393
rect 457 -1394 836 -1393
rect 51 -1396 139 -1395
rect 163 -1396 185 -1395
rect 226 -1396 311 -1395
rect 324 -1396 353 -1395
rect 394 -1396 423 -1395
rect 450 -1396 458 -1395
rect 478 -1396 584 -1395
rect 590 -1396 703 -1395
rect 709 -1396 752 -1395
rect 51 -1398 388 -1397
rect 394 -1398 416 -1397
rect 488 -1398 528 -1397
rect 551 -1398 661 -1397
rect 674 -1398 682 -1397
rect 58 -1400 62 -1399
rect 75 -1400 167 -1399
rect 226 -1400 381 -1399
rect 404 -1400 710 -1399
rect 58 -1402 66 -1401
rect 75 -1402 206 -1401
rect 254 -1402 276 -1401
rect 303 -1402 388 -1401
rect 404 -1402 696 -1401
rect 61 -1404 66 -1403
rect 79 -1404 178 -1403
rect 205 -1404 300 -1403
rect 348 -1404 535 -1403
rect 555 -1404 717 -1403
rect 79 -1406 129 -1405
rect 261 -1406 304 -1405
rect 317 -1406 717 -1405
rect 86 -1408 101 -1407
rect 117 -1408 479 -1407
rect 506 -1408 626 -1407
rect 639 -1408 689 -1407
rect 89 -1410 248 -1409
rect 261 -1410 269 -1409
rect 282 -1410 318 -1409
rect 352 -1410 517 -1409
rect 520 -1410 591 -1409
rect 618 -1410 654 -1409
rect 93 -1412 612 -1411
rect 646 -1412 724 -1411
rect 30 -1414 94 -1413
rect 100 -1414 241 -1413
rect 359 -1414 451 -1413
rect 506 -1414 612 -1413
rect 23 -1416 31 -1415
rect 107 -1416 118 -1415
rect 128 -1416 199 -1415
rect 219 -1416 283 -1415
rect 359 -1416 374 -1415
rect 411 -1416 416 -1415
rect 432 -1416 556 -1415
rect 562 -1416 633 -1415
rect 23 -1418 472 -1417
rect 492 -1418 633 -1417
rect 198 -1420 290 -1419
rect 366 -1420 493 -1419
rect 513 -1420 619 -1419
rect 219 -1422 430 -1421
rect 439 -1422 514 -1421
rect 520 -1422 692 -1421
rect 233 -1424 290 -1423
rect 334 -1424 367 -1423
rect 527 -1424 549 -1423
rect 565 -1424 661 -1423
rect 191 -1426 234 -1425
rect 240 -1426 255 -1425
rect 268 -1426 374 -1425
rect 541 -1426 640 -1425
rect 191 -1428 766 -1427
rect 541 -1430 706 -1429
rect 548 -1432 682 -1431
rect 572 -1434 668 -1433
rect 583 -1436 605 -1435
rect 667 -1436 769 -1435
rect 485 -1438 605 -1437
rect 485 -1440 570 -1439
rect 597 -1440 647 -1439
rect 499 -1442 598 -1441
rect 436 -1444 500 -1443
rect 9 -1455 97 -1454
rect 128 -1455 549 -1454
rect 681 -1455 790 -1454
rect 800 -1455 815 -1454
rect 817 -1455 829 -1454
rect 9 -1457 780 -1456
rect 16 -1459 437 -1458
rect 439 -1459 633 -1458
rect 681 -1459 738 -1458
rect 768 -1459 808 -1458
rect 16 -1461 472 -1460
rect 474 -1461 752 -1460
rect 23 -1463 139 -1462
rect 156 -1463 724 -1462
rect 737 -1463 773 -1462
rect 23 -1465 164 -1464
rect 198 -1465 381 -1464
rect 394 -1465 423 -1464
rect 429 -1465 605 -1464
rect 632 -1465 668 -1464
rect 674 -1465 724 -1464
rect 30 -1467 185 -1466
rect 250 -1467 419 -1466
rect 422 -1467 493 -1466
rect 509 -1467 689 -1466
rect 30 -1469 181 -1468
rect 257 -1469 612 -1468
rect 667 -1469 717 -1468
rect 37 -1471 167 -1470
rect 268 -1471 297 -1470
rect 303 -1471 472 -1470
rect 523 -1471 626 -1470
rect 688 -1471 745 -1470
rect 44 -1473 118 -1472
rect 128 -1473 143 -1472
rect 159 -1473 409 -1472
rect 432 -1473 640 -1472
rect 54 -1475 717 -1474
rect 58 -1477 73 -1476
rect 79 -1477 83 -1476
rect 114 -1477 139 -1476
rect 142 -1477 178 -1476
rect 296 -1477 370 -1476
rect 383 -1477 612 -1476
rect 37 -1479 384 -1478
rect 401 -1479 458 -1478
rect 527 -1479 605 -1478
rect 44 -1481 178 -1480
rect 212 -1481 458 -1480
rect 464 -1481 528 -1480
rect 534 -1481 538 -1480
rect 541 -1481 626 -1480
rect 58 -1483 87 -1482
rect 135 -1483 157 -1482
rect 212 -1483 255 -1482
rect 306 -1483 731 -1482
rect 65 -1485 125 -1484
rect 331 -1485 346 -1484
rect 352 -1485 507 -1484
rect 513 -1485 542 -1484
rect 555 -1485 745 -1484
rect 65 -1487 150 -1486
rect 289 -1487 346 -1486
rect 359 -1487 430 -1486
rect 439 -1487 647 -1486
rect 79 -1489 101 -1488
rect 149 -1489 220 -1488
rect 289 -1489 374 -1488
rect 390 -1489 465 -1488
rect 478 -1489 514 -1488
rect 534 -1489 619 -1488
rect 646 -1489 836 -1488
rect 86 -1491 276 -1490
rect 317 -1491 353 -1490
rect 366 -1491 493 -1490
rect 555 -1491 584 -1490
rect 597 -1491 752 -1490
rect 170 -1493 220 -1492
rect 233 -1493 276 -1492
rect 282 -1493 318 -1492
rect 331 -1493 577 -1492
rect 597 -1493 731 -1492
rect 93 -1495 171 -1494
rect 191 -1495 374 -1494
rect 387 -1495 479 -1494
rect 562 -1495 675 -1494
rect 121 -1497 192 -1496
rect 233 -1497 272 -1496
rect 310 -1497 388 -1496
rect 397 -1497 577 -1496
rect 618 -1497 654 -1496
rect 107 -1499 122 -1498
rect 247 -1499 311 -1498
rect 334 -1499 661 -1498
rect 107 -1501 188 -1500
rect 198 -1501 248 -1500
rect 261 -1501 283 -1500
rect 338 -1501 402 -1500
rect 450 -1501 640 -1500
rect 653 -1501 696 -1500
rect 240 -1503 262 -1502
rect 324 -1503 339 -1502
rect 341 -1503 584 -1502
rect 660 -1503 703 -1502
rect 240 -1505 405 -1504
rect 450 -1505 500 -1504
rect 520 -1505 563 -1504
rect 324 -1507 444 -1506
rect 485 -1507 521 -1506
rect 537 -1507 696 -1506
rect 226 -1509 444 -1508
rect 205 -1511 227 -1510
rect 362 -1511 703 -1510
rect 366 -1513 710 -1512
rect 380 -1515 710 -1514
rect 415 -1517 500 -1516
rect 415 -1519 591 -1518
rect 569 -1521 591 -1520
rect 359 -1523 570 -1522
rect 12 -1534 17 -1533
rect 51 -1534 206 -1533
rect 208 -1534 262 -1533
rect 303 -1534 318 -1533
rect 331 -1534 437 -1533
rect 488 -1534 745 -1533
rect 16 -1536 213 -1535
rect 240 -1536 325 -1535
rect 338 -1536 472 -1535
rect 520 -1536 605 -1535
rect 618 -1536 668 -1535
rect 2 -1538 325 -1537
rect 341 -1538 668 -1537
rect 23 -1540 206 -1539
rect 212 -1540 290 -1539
rect 303 -1540 640 -1539
rect 23 -1542 346 -1541
rect 362 -1542 444 -1541
rect 471 -1542 703 -1541
rect 44 -1544 332 -1543
rect 341 -1544 500 -1543
rect 597 -1544 738 -1543
rect 44 -1546 570 -1545
rect 604 -1546 654 -1545
rect 51 -1548 129 -1547
rect 138 -1548 479 -1547
rect 499 -1548 752 -1547
rect 58 -1550 97 -1549
rect 103 -1550 192 -1549
rect 233 -1550 479 -1549
rect 569 -1550 633 -1549
rect 653 -1550 710 -1549
rect 58 -1552 171 -1551
rect 184 -1552 276 -1551
rect 278 -1552 598 -1551
rect 632 -1552 689 -1551
rect 72 -1554 101 -1553
rect 117 -1554 122 -1553
rect 128 -1554 321 -1553
rect 345 -1554 542 -1553
rect 79 -1556 90 -1555
rect 93 -1556 115 -1555
rect 121 -1556 297 -1555
rect 306 -1556 458 -1555
rect 82 -1558 255 -1557
rect 257 -1558 549 -1557
rect 86 -1560 269 -1559
rect 289 -1560 409 -1559
rect 415 -1560 647 -1559
rect 65 -1562 409 -1561
rect 415 -1562 423 -1561
rect 443 -1562 535 -1561
rect 548 -1562 601 -1561
rect 646 -1562 696 -1561
rect 30 -1564 66 -1563
rect 138 -1564 220 -1563
rect 247 -1564 402 -1563
rect 422 -1564 507 -1563
rect 534 -1564 612 -1563
rect 30 -1566 584 -1565
rect 611 -1566 661 -1565
rect 149 -1568 164 -1567
rect 170 -1568 237 -1567
rect 247 -1568 283 -1567
rect 296 -1568 514 -1567
rect 555 -1568 584 -1567
rect 660 -1568 717 -1567
rect 152 -1570 353 -1569
rect 362 -1570 542 -1569
rect 37 -1572 353 -1571
rect 366 -1572 493 -1571
rect 37 -1574 108 -1573
rect 184 -1574 199 -1573
rect 219 -1574 640 -1573
rect 9 -1576 108 -1575
rect 177 -1576 199 -1575
rect 250 -1576 374 -1575
rect 380 -1576 451 -1575
rect 457 -1576 577 -1575
rect 114 -1578 381 -1577
rect 387 -1578 675 -1577
rect 156 -1580 178 -1579
rect 187 -1580 192 -1579
rect 261 -1580 311 -1579
rect 313 -1580 430 -1579
rect 439 -1580 507 -1579
rect 674 -1580 724 -1579
rect 142 -1582 157 -1581
rect 275 -1582 374 -1581
rect 401 -1582 528 -1581
rect 282 -1584 311 -1583
rect 334 -1584 514 -1583
rect 306 -1586 528 -1585
rect 418 -1588 451 -1587
rect 485 -1588 577 -1587
rect 387 -1590 486 -1589
rect 492 -1590 591 -1589
rect 411 -1592 591 -1591
rect 429 -1594 465 -1593
rect 464 -1596 563 -1595
rect 562 -1598 626 -1597
rect 625 -1600 682 -1599
rect 681 -1602 731 -1601
rect 5 -1613 325 -1612
rect 359 -1613 472 -1612
rect 485 -1613 521 -1612
rect 558 -1613 647 -1612
rect 9 -1615 157 -1614
rect 187 -1615 199 -1614
rect 226 -1615 279 -1614
rect 317 -1615 500 -1614
rect 520 -1615 577 -1614
rect 625 -1615 650 -1614
rect 23 -1617 80 -1616
rect 82 -1617 640 -1616
rect 23 -1619 111 -1618
rect 114 -1619 300 -1618
rect 359 -1619 535 -1618
rect 30 -1621 325 -1620
rect 362 -1621 395 -1620
rect 401 -1621 409 -1620
rect 411 -1621 633 -1620
rect 30 -1623 220 -1622
rect 233 -1623 248 -1622
rect 254 -1623 318 -1622
rect 366 -1623 465 -1622
rect 478 -1623 500 -1622
rect 534 -1623 605 -1622
rect 16 -1625 465 -1624
rect 16 -1627 139 -1626
rect 152 -1627 255 -1626
rect 268 -1627 311 -1626
rect 373 -1627 479 -1626
rect 37 -1629 101 -1628
rect 128 -1629 157 -1628
rect 170 -1629 227 -1628
rect 240 -1629 269 -1628
rect 376 -1629 388 -1628
rect 394 -1629 507 -1628
rect 37 -1631 307 -1630
rect 380 -1631 472 -1630
rect 506 -1631 612 -1630
rect 65 -1633 276 -1632
rect 292 -1633 612 -1632
rect 58 -1635 66 -1634
rect 72 -1635 143 -1634
rect 173 -1635 199 -1634
rect 205 -1635 248 -1634
rect 275 -1635 353 -1634
rect 380 -1635 430 -1634
rect 436 -1635 458 -1634
rect 58 -1637 192 -1636
rect 205 -1637 370 -1636
rect 401 -1637 423 -1636
rect 429 -1637 451 -1636
rect 457 -1637 556 -1636
rect 47 -1639 192 -1638
rect 212 -1639 234 -1638
rect 296 -1639 388 -1638
rect 408 -1639 661 -1638
rect 51 -1641 423 -1640
rect 439 -1641 591 -1640
rect 660 -1641 675 -1640
rect 51 -1643 339 -1642
rect 443 -1643 598 -1642
rect 86 -1645 150 -1644
rect 184 -1645 220 -1644
rect 296 -1645 577 -1644
rect 597 -1645 682 -1644
rect 72 -1647 87 -1646
rect 89 -1647 654 -1646
rect 677 -1647 682 -1646
rect 93 -1649 118 -1648
rect 128 -1649 178 -1648
rect 194 -1649 591 -1648
rect 93 -1651 122 -1650
rect 135 -1651 178 -1650
rect 212 -1651 262 -1650
rect 331 -1651 339 -1650
rect 443 -1651 514 -1650
rect 107 -1653 136 -1652
rect 446 -1653 556 -1652
rect 114 -1655 171 -1654
rect 450 -1655 542 -1654
rect 121 -1657 290 -1656
rect 320 -1657 542 -1656
rect 282 -1659 290 -1658
rect 513 -1659 563 -1658
rect 282 -1661 416 -1660
rect 548 -1661 563 -1660
rect 345 -1663 416 -1662
rect 548 -1663 570 -1662
rect 345 -1665 493 -1664
rect 569 -1665 619 -1664
rect 492 -1667 528 -1666
rect 527 -1669 584 -1668
rect 583 -1671 668 -1670
rect 16 -1682 87 -1681
rect 107 -1682 160 -1681
rect 170 -1682 178 -1681
rect 187 -1682 423 -1681
rect 446 -1682 493 -1681
rect 506 -1682 654 -1681
rect 674 -1682 682 -1681
rect 16 -1684 94 -1683
rect 145 -1684 297 -1683
rect 306 -1684 472 -1683
rect 534 -1684 580 -1683
rect 649 -1684 661 -1683
rect 23 -1686 143 -1685
rect 156 -1686 192 -1685
rect 212 -1686 262 -1685
rect 264 -1686 465 -1685
rect 471 -1686 514 -1685
rect 548 -1686 622 -1685
rect 23 -1688 346 -1687
rect 352 -1688 591 -1687
rect 30 -1690 227 -1689
rect 243 -1690 325 -1689
rect 331 -1690 542 -1689
rect 569 -1690 619 -1689
rect 37 -1692 314 -1691
rect 317 -1692 360 -1691
rect 376 -1692 500 -1691
rect 597 -1692 619 -1691
rect 9 -1694 318 -1693
rect 320 -1694 409 -1693
rect 499 -1694 528 -1693
rect 9 -1696 129 -1695
rect 173 -1696 335 -1695
rect 338 -1696 577 -1695
rect 40 -1698 199 -1697
rect 212 -1698 276 -1697
rect 282 -1698 356 -1697
rect 390 -1698 444 -1697
rect 527 -1698 612 -1697
rect 44 -1700 132 -1699
rect 187 -1700 237 -1699
rect 247 -1700 290 -1699
rect 292 -1700 297 -1699
rect 310 -1700 360 -1699
rect 408 -1700 437 -1699
rect 47 -1702 59 -1701
rect 65 -1702 262 -1701
rect 271 -1702 465 -1701
rect 51 -1704 258 -1703
rect 275 -1704 395 -1703
rect 436 -1704 451 -1703
rect 58 -1706 521 -1705
rect 65 -1708 129 -1707
rect 198 -1708 234 -1707
rect 247 -1708 374 -1707
rect 380 -1708 395 -1707
rect 520 -1708 563 -1707
rect 72 -1710 125 -1709
rect 219 -1710 227 -1709
rect 250 -1710 493 -1709
rect 72 -1712 206 -1711
rect 254 -1712 325 -1711
rect 331 -1712 416 -1711
rect 79 -1714 290 -1713
rect 310 -1714 479 -1713
rect 79 -1716 269 -1715
rect 282 -1716 430 -1715
rect 86 -1718 115 -1717
rect 121 -1718 234 -1717
rect 240 -1718 479 -1717
rect 107 -1720 143 -1719
rect 149 -1720 220 -1719
rect 268 -1720 367 -1719
rect 373 -1720 423 -1719
rect 429 -1720 486 -1719
rect 114 -1722 136 -1721
rect 345 -1722 402 -1721
rect 485 -1722 556 -1721
rect 121 -1724 381 -1723
rect 401 -1724 458 -1723
rect 555 -1724 584 -1723
rect 135 -1726 164 -1725
rect 303 -1726 458 -1725
rect 163 -1728 185 -1727
rect 362 -1728 416 -1727
rect 16 -1739 153 -1738
rect 156 -1739 241 -1738
rect 254 -1739 258 -1738
rect 261 -1739 353 -1738
rect 418 -1739 535 -1738
rect 548 -1739 556 -1738
rect 632 -1739 654 -1738
rect 670 -1739 675 -1738
rect 23 -1741 363 -1740
rect 422 -1741 454 -1740
rect 460 -1741 521 -1740
rect 37 -1743 108 -1742
rect 114 -1743 178 -1742
rect 208 -1743 297 -1742
rect 331 -1743 353 -1742
rect 408 -1743 461 -1742
rect 471 -1743 514 -1742
rect 44 -1745 311 -1744
rect 334 -1745 493 -1744
rect 51 -1747 293 -1746
rect 296 -1747 367 -1746
rect 422 -1747 479 -1746
rect 51 -1749 136 -1748
rect 145 -1749 220 -1748
rect 226 -1749 244 -1748
rect 282 -1749 318 -1748
rect 338 -1749 402 -1748
rect 429 -1749 489 -1748
rect 58 -1751 356 -1750
rect 429 -1751 465 -1750
rect 471 -1751 528 -1750
rect 65 -1753 94 -1752
rect 117 -1753 206 -1752
rect 212 -1753 269 -1752
rect 289 -1753 325 -1752
rect 345 -1753 367 -1752
rect 394 -1753 465 -1752
rect 478 -1753 486 -1752
rect 499 -1753 528 -1752
rect 72 -1755 136 -1754
rect 152 -1755 192 -1754
rect 219 -1755 304 -1754
rect 310 -1755 405 -1754
rect 436 -1755 521 -1754
rect 72 -1757 80 -1756
rect 86 -1757 104 -1756
rect 124 -1757 143 -1756
rect 159 -1757 192 -1756
rect 268 -1757 381 -1756
rect 65 -1759 160 -1758
rect 163 -1759 227 -1758
rect 275 -1759 346 -1758
rect 86 -1761 122 -1760
rect 128 -1761 251 -1760
rect 324 -1761 416 -1760
rect 93 -1763 108 -1762
rect 163 -1763 262 -1762
rect 173 -1765 199 -1764
rect 233 -1765 276 -1764
rect 9 -1767 199 -1766
rect 170 -1769 234 -1768
rect 51 -1780 185 -1779
rect 198 -1780 251 -1779
rect 254 -1780 290 -1779
rect 317 -1780 384 -1779
rect 387 -1780 430 -1779
rect 464 -1780 486 -1779
rect 499 -1780 535 -1779
rect 541 -1780 549 -1779
rect 614 -1780 633 -1779
rect 51 -1782 62 -1781
rect 72 -1782 335 -1781
rect 345 -1782 412 -1781
rect 467 -1782 521 -1781
rect 618 -1782 640 -1781
rect 86 -1784 104 -1783
rect 110 -1784 213 -1783
rect 247 -1784 325 -1783
rect 352 -1784 419 -1783
rect 478 -1784 503 -1783
rect 513 -1784 563 -1783
rect 93 -1786 104 -1785
rect 117 -1786 129 -1785
rect 135 -1786 150 -1785
rect 156 -1786 227 -1785
rect 264 -1786 311 -1785
rect 338 -1786 353 -1785
rect 366 -1786 419 -1785
rect 520 -1786 528 -1785
rect 65 -1788 118 -1787
rect 124 -1788 241 -1787
rect 296 -1788 311 -1787
rect 373 -1788 423 -1787
rect 89 -1790 136 -1789
rect 138 -1790 157 -1789
rect 163 -1790 269 -1789
rect 142 -1792 160 -1791
rect 173 -1792 192 -1791
rect 205 -1792 220 -1791
rect 37 -1794 143 -1793
rect 177 -1794 234 -1793
rect 233 -1796 262 -1795
rect 131 -1798 262 -1797
rect 51 -1809 62 -1808
rect 145 -1809 206 -1808
rect 233 -1809 272 -1808
rect 352 -1809 419 -1808
rect 471 -1809 479 -1808
rect 520 -1809 528 -1808
rect 149 -1811 185 -1810
rect 156 -1813 178 -1812
rect 180 -1813 262 -1812
<< m2contact >>
rect 58 0 59 1
rect 93 0 94 1
rect 114 0 115 1
rect 142 0 143 1
rect 152 0 153 1
rect 170 0 171 1
rect 177 0 178 1
rect 212 0 213 1
rect 257 0 258 1
rect 261 0 262 1
rect 124 -2 125 -1
rect 240 -2 241 -1
rect 128 -4 129 -3
rect 135 -4 136 -3
rect 156 -4 157 -3
rect 163 -4 164 -3
rect 184 -4 185 -3
rect 191 -4 192 -3
rect 198 -4 199 -3
rect 236 -4 237 -3
rect 205 -6 206 -5
rect 338 -6 339 -5
rect 44 -17 45 -16
rect 47 -17 48 -16
rect 72 -17 73 -16
rect 93 -17 94 -16
rect 103 -17 104 -16
rect 275 -17 276 -16
rect 285 -17 286 -16
rect 345 -17 346 -16
rect 79 -19 80 -18
rect 191 -19 192 -18
rect 205 -19 206 -18
rect 317 -19 318 -18
rect 338 -19 339 -18
rect 387 -19 388 -18
rect 114 -21 115 -20
rect 131 -21 132 -20
rect 177 -21 178 -20
rect 198 -21 199 -20
rect 205 -21 206 -20
rect 324 -21 325 -20
rect 124 -23 125 -22
rect 212 -23 213 -22
rect 222 -23 223 -22
rect 240 -23 241 -22
rect 247 -23 248 -22
rect 334 -23 335 -22
rect 128 -25 129 -24
rect 135 -25 136 -24
rect 149 -25 150 -24
rect 177 -25 178 -24
rect 184 -25 185 -24
rect 219 -25 220 -24
rect 240 -25 241 -24
rect 261 -25 262 -24
rect 271 -25 272 -24
rect 352 -25 353 -24
rect 93 -27 94 -26
rect 128 -27 129 -26
rect 163 -27 164 -26
rect 198 -27 199 -26
rect 212 -27 213 -26
rect 226 -27 227 -26
rect 254 -27 255 -26
rect 282 -27 283 -26
rect 289 -27 290 -26
rect 296 -27 297 -26
rect 313 -27 314 -26
rect 338 -27 339 -26
rect 170 -29 171 -28
rect 184 -29 185 -28
rect 226 -29 227 -28
rect 233 -29 234 -28
rect 142 -31 143 -30
rect 233 -31 234 -30
rect 163 -33 164 -32
rect 170 -33 171 -32
rect 16 -44 17 -43
rect 240 -44 241 -43
rect 254 -44 255 -43
rect 341 -44 342 -43
rect 345 -44 346 -43
rect 436 -44 437 -43
rect 23 -46 24 -45
rect 117 -46 118 -45
rect 128 -46 129 -45
rect 156 -46 157 -45
rect 163 -46 164 -45
rect 170 -46 171 -45
rect 191 -46 192 -45
rect 222 -46 223 -45
rect 233 -46 234 -45
rect 310 -46 311 -45
rect 317 -46 318 -45
rect 380 -46 381 -45
rect 387 -46 388 -45
rect 408 -46 409 -45
rect 44 -48 45 -47
rect 58 -48 59 -47
rect 65 -48 66 -47
rect 107 -48 108 -47
rect 114 -48 115 -47
rect 121 -48 122 -47
rect 135 -48 136 -47
rect 142 -48 143 -47
rect 156 -48 157 -47
rect 194 -48 195 -47
rect 205 -48 206 -47
rect 219 -48 220 -47
rect 247 -48 248 -47
rect 254 -48 255 -47
rect 275 -48 276 -47
rect 331 -48 332 -47
rect 338 -48 339 -47
rect 422 -48 423 -47
rect 51 -50 52 -49
rect 345 -50 346 -49
rect 352 -50 353 -49
rect 401 -50 402 -49
rect 404 -50 405 -49
rect 415 -50 416 -49
rect 61 -52 62 -51
rect 205 -52 206 -51
rect 208 -52 209 -51
rect 226 -52 227 -51
rect 268 -52 269 -51
rect 275 -52 276 -51
rect 282 -52 283 -51
rect 317 -52 318 -51
rect 324 -52 325 -51
rect 387 -52 388 -51
rect 72 -54 73 -53
rect 152 -54 153 -53
rect 170 -54 171 -53
rect 180 -54 181 -53
rect 184 -54 185 -53
rect 226 -54 227 -53
rect 296 -54 297 -53
rect 359 -54 360 -53
rect 373 -54 374 -53
rect 394 -54 395 -53
rect 82 -56 83 -55
rect 135 -56 136 -55
rect 184 -56 185 -55
rect 240 -56 241 -55
rect 299 -56 300 -55
rect 366 -56 367 -55
rect 86 -58 87 -57
rect 177 -58 178 -57
rect 212 -58 213 -57
rect 233 -58 234 -57
rect 93 -60 94 -59
rect 324 -60 325 -59
rect 93 -62 94 -61
rect 292 -62 293 -61
rect 100 -64 101 -63
rect 110 -64 111 -63
rect 177 -64 178 -63
rect 198 -64 199 -63
rect 212 -64 213 -63
rect 271 -64 272 -63
rect 198 -66 199 -65
rect 289 -66 290 -65
rect 261 -68 262 -67
rect 271 -68 272 -67
rect 23 -79 24 -78
rect 198 -79 199 -78
rect 205 -79 206 -78
rect 506 -79 507 -78
rect 37 -81 38 -80
rect 219 -81 220 -80
rect 233 -81 234 -80
rect 247 -81 248 -80
rect 250 -81 251 -80
rect 464 -81 465 -80
rect 44 -83 45 -82
rect 296 -83 297 -82
rect 303 -83 304 -82
rect 394 -83 395 -82
rect 397 -83 398 -82
rect 457 -83 458 -82
rect 58 -85 59 -84
rect 156 -85 157 -84
rect 170 -85 171 -84
rect 205 -85 206 -84
rect 208 -85 209 -84
rect 240 -85 241 -84
rect 254 -85 255 -84
rect 268 -85 269 -84
rect 275 -85 276 -84
rect 303 -85 304 -84
rect 373 -85 374 -84
rect 429 -85 430 -84
rect 436 -85 437 -84
rect 513 -85 514 -84
rect 65 -87 66 -86
rect 152 -87 153 -86
rect 156 -87 157 -86
rect 247 -87 248 -86
rect 254 -87 255 -86
rect 317 -87 318 -86
rect 345 -87 346 -86
rect 436 -87 437 -86
rect 72 -89 73 -88
rect 114 -89 115 -88
rect 121 -89 122 -88
rect 198 -89 199 -88
rect 222 -89 223 -88
rect 317 -89 318 -88
rect 338 -89 339 -88
rect 345 -89 346 -88
rect 380 -89 381 -88
rect 471 -89 472 -88
rect 79 -91 80 -90
rect 261 -91 262 -90
rect 275 -91 276 -90
rect 310 -91 311 -90
rect 387 -91 388 -90
rect 492 -91 493 -90
rect 16 -93 17 -92
rect 261 -93 262 -92
rect 285 -93 286 -92
rect 450 -93 451 -92
rect 86 -95 87 -94
rect 100 -95 101 -94
rect 107 -95 108 -94
rect 212 -95 213 -94
rect 292 -95 293 -94
rect 422 -95 423 -94
rect 93 -97 94 -96
rect 443 -97 444 -96
rect 93 -99 94 -98
rect 282 -99 283 -98
rect 310 -99 311 -98
rect 334 -99 335 -98
rect 380 -99 381 -98
rect 422 -99 423 -98
rect 128 -101 129 -100
rect 194 -101 195 -100
rect 212 -101 213 -100
rect 306 -101 307 -100
rect 401 -101 402 -100
rect 499 -101 500 -100
rect 128 -103 129 -102
rect 299 -103 300 -102
rect 359 -103 360 -102
rect 401 -103 402 -102
rect 408 -103 409 -102
rect 485 -103 486 -102
rect 135 -105 136 -104
rect 191 -105 192 -104
rect 324 -105 325 -104
rect 359 -105 360 -104
rect 366 -105 367 -104
rect 408 -105 409 -104
rect 415 -105 416 -104
rect 478 -105 479 -104
rect 149 -107 150 -106
rect 387 -107 388 -106
rect 149 -109 150 -108
rect 163 -109 164 -108
rect 173 -109 174 -108
rect 289 -109 290 -108
rect 331 -109 332 -108
rect 366 -109 367 -108
rect 373 -109 374 -108
rect 415 -109 416 -108
rect 121 -111 122 -110
rect 289 -111 290 -110
rect 331 -111 332 -110
rect 520 -111 521 -110
rect 177 -113 178 -112
rect 233 -113 234 -112
rect 187 -115 188 -114
rect 226 -115 227 -114
rect 142 -117 143 -116
rect 226 -117 227 -116
rect 142 -119 143 -118
rect 184 -119 185 -118
rect 163 -121 164 -120
rect 187 -121 188 -120
rect 12 -132 13 -131
rect 72 -132 73 -131
rect 75 -132 76 -131
rect 506 -132 507 -131
rect 520 -132 521 -131
rect 660 -132 661 -131
rect 51 -134 52 -133
rect 177 -134 178 -133
rect 180 -134 181 -133
rect 359 -134 360 -133
rect 373 -134 374 -133
rect 376 -134 377 -133
rect 383 -134 384 -133
rect 464 -134 465 -133
rect 471 -134 472 -133
rect 618 -134 619 -133
rect 58 -136 59 -135
rect 285 -136 286 -135
rect 296 -136 297 -135
rect 331 -136 332 -135
rect 334 -136 335 -135
rect 443 -136 444 -135
rect 457 -136 458 -135
rect 583 -136 584 -135
rect 58 -138 59 -137
rect 243 -138 244 -137
rect 250 -138 251 -137
rect 268 -138 269 -137
rect 282 -138 283 -137
rect 401 -138 402 -137
rect 415 -138 416 -137
rect 569 -138 570 -137
rect 79 -140 80 -139
rect 401 -140 402 -139
rect 422 -140 423 -139
rect 443 -140 444 -139
rect 478 -140 479 -139
rect 639 -140 640 -139
rect 79 -142 80 -141
rect 103 -142 104 -141
rect 121 -142 122 -141
rect 527 -142 528 -141
rect 44 -144 45 -143
rect 121 -144 122 -143
rect 128 -144 129 -143
rect 380 -144 381 -143
rect 390 -144 391 -143
rect 653 -144 654 -143
rect 44 -146 45 -145
rect 187 -146 188 -145
rect 240 -146 241 -145
rect 275 -146 276 -145
rect 282 -146 283 -145
rect 506 -146 507 -145
rect 513 -146 514 -145
rect 520 -146 521 -145
rect 89 -148 90 -147
rect 198 -148 199 -147
rect 247 -148 248 -147
rect 275 -148 276 -147
rect 292 -148 293 -147
rect 457 -148 458 -147
rect 499 -148 500 -147
rect 632 -148 633 -147
rect 93 -150 94 -149
rect 478 -150 479 -149
rect 485 -150 486 -149
rect 499 -150 500 -149
rect 93 -152 94 -151
rect 271 -152 272 -151
rect 296 -152 297 -151
rect 324 -152 325 -151
rect 327 -152 328 -151
rect 604 -152 605 -151
rect 100 -154 101 -153
rect 562 -154 563 -153
rect 100 -156 101 -155
rect 149 -156 150 -155
rect 152 -156 153 -155
rect 534 -156 535 -155
rect 128 -158 129 -157
rect 219 -158 220 -157
rect 261 -158 262 -157
rect 415 -158 416 -157
rect 422 -158 423 -157
rect 471 -158 472 -157
rect 107 -160 108 -159
rect 261 -160 262 -159
rect 303 -160 304 -159
rect 359 -160 360 -159
rect 373 -160 374 -159
rect 450 -160 451 -159
rect 107 -162 108 -161
rect 159 -162 160 -161
rect 170 -162 171 -161
rect 548 -162 549 -161
rect 117 -164 118 -163
rect 219 -164 220 -163
rect 226 -164 227 -163
rect 303 -164 304 -163
rect 341 -164 342 -163
rect 597 -164 598 -163
rect 135 -166 136 -165
rect 611 -166 612 -165
rect 138 -168 139 -167
rect 142 -168 143 -167
rect 149 -168 150 -167
rect 464 -168 465 -167
rect 142 -170 143 -169
rect 289 -170 290 -169
rect 352 -170 353 -169
rect 492 -170 493 -169
rect 156 -172 157 -171
rect 187 -172 188 -171
rect 191 -172 192 -171
rect 352 -172 353 -171
rect 376 -172 377 -171
rect 450 -172 451 -171
rect 170 -174 171 -173
rect 233 -174 234 -173
rect 289 -174 290 -173
rect 492 -174 493 -173
rect 177 -176 178 -175
rect 590 -176 591 -175
rect 180 -178 181 -177
rect 240 -178 241 -177
rect 387 -178 388 -177
rect 513 -178 514 -177
rect 191 -180 192 -179
rect 254 -180 255 -179
rect 324 -180 325 -179
rect 387 -180 388 -179
rect 394 -180 395 -179
rect 646 -180 647 -179
rect 198 -182 199 -181
rect 625 -182 626 -181
rect 205 -184 206 -183
rect 226 -184 227 -183
rect 317 -184 318 -183
rect 394 -184 395 -183
rect 408 -184 409 -183
rect 485 -184 486 -183
rect 135 -186 136 -185
rect 317 -186 318 -185
rect 408 -186 409 -185
rect 576 -186 577 -185
rect 212 -188 213 -187
rect 233 -188 234 -187
rect 429 -188 430 -187
rect 555 -188 556 -187
rect 366 -190 367 -189
rect 429 -190 430 -189
rect 436 -190 437 -189
rect 541 -190 542 -189
rect 86 -192 87 -191
rect 436 -192 437 -191
rect 345 -194 346 -193
rect 366 -194 367 -193
rect 310 -196 311 -195
rect 345 -196 346 -195
rect 33 -207 34 -206
rect 590 -207 591 -206
rect 597 -207 598 -206
rect 667 -207 668 -206
rect 51 -209 52 -208
rect 212 -209 213 -208
rect 215 -209 216 -208
rect 604 -209 605 -208
rect 65 -211 66 -210
rect 201 -211 202 -210
rect 205 -211 206 -210
rect 240 -211 241 -210
rect 243 -211 244 -210
rect 513 -211 514 -210
rect 520 -211 521 -210
rect 604 -211 605 -210
rect 79 -213 80 -212
rect 306 -213 307 -212
rect 310 -213 311 -212
rect 324 -213 325 -212
rect 338 -213 339 -212
rect 625 -213 626 -212
rect 44 -215 45 -214
rect 324 -215 325 -214
rect 366 -215 367 -214
rect 408 -215 409 -214
rect 411 -215 412 -214
rect 506 -215 507 -214
rect 513 -215 514 -214
rect 527 -215 528 -214
rect 590 -215 591 -214
rect 632 -215 633 -214
rect 89 -217 90 -216
rect 422 -217 423 -216
rect 464 -217 465 -216
rect 520 -217 521 -216
rect 527 -217 528 -216
rect 541 -217 542 -216
rect 597 -217 598 -216
rect 639 -217 640 -216
rect 100 -219 101 -218
rect 180 -219 181 -218
rect 187 -219 188 -218
rect 226 -219 227 -218
rect 254 -219 255 -218
rect 345 -219 346 -218
rect 373 -219 374 -218
rect 541 -219 542 -218
rect 625 -219 626 -218
rect 653 -219 654 -218
rect 103 -221 104 -220
rect 177 -221 178 -220
rect 198 -221 199 -220
rect 457 -221 458 -220
rect 464 -221 465 -220
rect 485 -221 486 -220
rect 632 -221 633 -220
rect 660 -221 661 -220
rect 72 -223 73 -222
rect 198 -223 199 -222
rect 208 -223 209 -222
rect 534 -223 535 -222
rect 72 -225 73 -224
rect 82 -225 83 -224
rect 114 -225 115 -224
rect 184 -225 185 -224
rect 219 -225 220 -224
rect 226 -225 227 -224
rect 247 -225 248 -224
rect 457 -225 458 -224
rect 485 -225 486 -224
rect 562 -225 563 -224
rect 58 -227 59 -226
rect 219 -227 220 -226
rect 257 -227 258 -226
rect 359 -227 360 -226
rect 373 -227 374 -226
rect 401 -227 402 -226
rect 499 -227 500 -226
rect 562 -227 563 -226
rect 58 -229 59 -228
rect 506 -229 507 -228
rect 534 -229 535 -228
rect 555 -229 556 -228
rect 114 -231 115 -230
rect 191 -231 192 -230
rect 257 -231 258 -230
rect 576 -231 577 -230
rect 121 -233 122 -232
rect 345 -233 346 -232
rect 359 -233 360 -232
rect 380 -233 381 -232
rect 387 -233 388 -232
rect 583 -233 584 -232
rect 121 -235 122 -234
rect 583 -235 584 -234
rect 124 -237 125 -236
rect 303 -237 304 -236
rect 313 -237 314 -236
rect 548 -237 549 -236
rect 65 -239 66 -238
rect 303 -239 304 -238
rect 317 -239 318 -238
rect 401 -239 402 -238
rect 548 -239 549 -238
rect 618 -239 619 -238
rect 128 -241 129 -240
rect 380 -241 381 -240
rect 387 -241 388 -240
rect 429 -241 430 -240
rect 576 -241 577 -240
rect 618 -241 619 -240
rect 128 -243 129 -242
rect 240 -243 241 -242
rect 268 -243 269 -242
rect 611 -243 612 -242
rect 135 -245 136 -244
rect 352 -245 353 -244
rect 429 -245 430 -244
rect 471 -245 472 -244
rect 100 -247 101 -246
rect 135 -247 136 -246
rect 142 -247 143 -246
rect 163 -247 164 -246
rect 170 -247 171 -246
rect 212 -247 213 -246
rect 268 -247 269 -246
rect 499 -247 500 -246
rect 93 -249 94 -248
rect 170 -249 171 -248
rect 191 -249 192 -248
rect 250 -249 251 -248
rect 275 -249 276 -248
rect 289 -249 290 -248
rect 292 -249 293 -248
rect 394 -249 395 -248
rect 443 -249 444 -248
rect 471 -249 472 -248
rect 89 -251 90 -250
rect 394 -251 395 -250
rect 436 -251 437 -250
rect 443 -251 444 -250
rect 93 -253 94 -252
rect 296 -253 297 -252
rect 299 -253 300 -252
rect 331 -253 332 -252
rect 334 -253 335 -252
rect 611 -253 612 -252
rect 107 -255 108 -254
rect 163 -255 164 -254
rect 282 -255 283 -254
rect 569 -255 570 -254
rect 107 -257 108 -256
rect 156 -257 157 -256
rect 180 -257 181 -256
rect 569 -257 570 -256
rect 142 -259 143 -258
rect 156 -259 157 -258
rect 320 -259 321 -258
rect 450 -259 451 -258
rect 149 -261 150 -260
rect 233 -261 234 -260
rect 285 -261 286 -260
rect 450 -261 451 -260
rect 23 -263 24 -262
rect 233 -263 234 -262
rect 285 -263 286 -262
rect 415 -263 416 -262
rect 425 -263 426 -262
rect 436 -263 437 -262
rect 152 -265 153 -264
rect 261 -265 262 -264
rect 282 -265 283 -264
rect 415 -265 416 -264
rect 261 -267 262 -266
rect 278 -267 279 -266
rect 331 -267 332 -266
rect 646 -267 647 -266
rect 338 -269 339 -268
rect 366 -269 367 -268
rect 44 -280 45 -279
rect 47 -280 48 -279
rect 58 -280 59 -279
rect 212 -280 213 -279
rect 247 -280 248 -279
rect 345 -280 346 -279
rect 355 -280 356 -279
rect 387 -280 388 -279
rect 390 -280 391 -279
rect 478 -280 479 -279
rect 506 -280 507 -279
rect 618 -280 619 -279
rect 667 -280 668 -279
rect 709 -280 710 -279
rect 58 -282 59 -281
rect 254 -282 255 -281
rect 261 -282 262 -281
rect 275 -282 276 -281
rect 282 -282 283 -281
rect 310 -282 311 -281
rect 317 -282 318 -281
rect 660 -282 661 -281
rect 72 -284 73 -283
rect 177 -284 178 -283
rect 187 -284 188 -283
rect 261 -284 262 -283
rect 282 -284 283 -283
rect 338 -284 339 -283
rect 341 -284 342 -283
rect 520 -284 521 -283
rect 555 -284 556 -283
rect 639 -284 640 -283
rect 72 -286 73 -285
rect 569 -286 570 -285
rect 583 -286 584 -285
rect 639 -286 640 -285
rect 89 -288 90 -287
rect 478 -288 479 -287
rect 513 -288 514 -287
rect 674 -288 675 -287
rect 89 -290 90 -289
rect 485 -290 486 -289
rect 527 -290 528 -289
rect 569 -290 570 -289
rect 590 -290 591 -289
rect 646 -290 647 -289
rect 100 -292 101 -291
rect 653 -292 654 -291
rect 107 -294 108 -293
rect 212 -294 213 -293
rect 285 -294 286 -293
rect 485 -294 486 -293
rect 492 -294 493 -293
rect 527 -294 528 -293
rect 534 -294 535 -293
rect 583 -294 584 -293
rect 604 -294 605 -293
rect 667 -294 668 -293
rect 16 -296 17 -295
rect 604 -296 605 -295
rect 107 -298 108 -297
rect 128 -298 129 -297
rect 145 -298 146 -297
rect 159 -298 160 -297
rect 163 -298 164 -297
rect 254 -298 255 -297
rect 296 -298 297 -297
rect 625 -298 626 -297
rect 54 -300 55 -299
rect 625 -300 626 -299
rect 65 -302 66 -301
rect 296 -302 297 -301
rect 299 -302 300 -301
rect 331 -302 332 -301
rect 362 -302 363 -301
rect 513 -302 514 -301
rect 541 -302 542 -301
rect 590 -302 591 -301
rect 114 -304 115 -303
rect 128 -304 129 -303
rect 149 -304 150 -303
rect 268 -304 269 -303
rect 306 -304 307 -303
rect 632 -304 633 -303
rect 114 -306 115 -305
rect 250 -306 251 -305
rect 320 -306 321 -305
rect 429 -306 430 -305
rect 450 -306 451 -305
rect 506 -306 507 -305
rect 541 -306 542 -305
rect 562 -306 563 -305
rect 30 -308 31 -307
rect 429 -308 430 -307
rect 436 -308 437 -307
rect 450 -308 451 -307
rect 464 -308 465 -307
rect 520 -308 521 -307
rect 562 -308 563 -307
rect 611 -308 612 -307
rect 30 -310 31 -309
rect 82 -310 83 -309
rect 121 -310 122 -309
rect 387 -310 388 -309
rect 415 -310 416 -309
rect 436 -310 437 -309
rect 443 -310 444 -309
rect 464 -310 465 -309
rect 499 -310 500 -309
rect 534 -310 535 -309
rect 576 -310 577 -309
rect 611 -310 612 -309
rect 23 -312 24 -311
rect 121 -312 122 -311
rect 142 -312 143 -311
rect 268 -312 269 -311
rect 320 -312 321 -311
rect 632 -312 633 -311
rect 159 -314 160 -313
rect 380 -314 381 -313
rect 408 -314 409 -313
rect 443 -314 444 -313
rect 471 -314 472 -313
rect 576 -314 577 -313
rect 65 -316 66 -315
rect 408 -316 409 -315
rect 415 -316 416 -315
rect 422 -316 423 -315
rect 457 -316 458 -315
rect 471 -316 472 -315
rect 79 -318 80 -317
rect 457 -318 458 -317
rect 51 -320 52 -319
rect 79 -320 80 -319
rect 142 -320 143 -319
rect 380 -320 381 -319
rect 394 -320 395 -319
rect 422 -320 423 -319
rect 37 -322 38 -321
rect 51 -322 52 -321
rect 170 -322 171 -321
rect 177 -322 178 -321
rect 191 -322 192 -321
rect 334 -322 335 -321
rect 352 -322 353 -321
rect 394 -322 395 -321
rect 135 -324 136 -323
rect 170 -324 171 -323
rect 191 -324 192 -323
rect 198 -324 199 -323
rect 201 -324 202 -323
rect 303 -324 304 -323
rect 324 -324 325 -323
rect 345 -324 346 -323
rect 366 -324 367 -323
rect 373 -324 374 -323
rect 135 -326 136 -325
rect 233 -326 234 -325
rect 313 -326 314 -325
rect 373 -326 374 -325
rect 184 -328 185 -327
rect 303 -328 304 -327
rect 324 -328 325 -327
rect 499 -328 500 -327
rect 149 -330 150 -329
rect 184 -330 185 -329
rect 205 -330 206 -329
rect 317 -330 318 -329
rect 369 -330 370 -329
rect 548 -330 549 -329
rect 93 -332 94 -331
rect 205 -332 206 -331
rect 233 -332 234 -331
rect 359 -332 360 -331
rect 548 -332 549 -331
rect 597 -332 598 -331
rect 93 -334 94 -333
rect 240 -334 241 -333
rect 9 -345 10 -344
rect 660 -345 661 -344
rect 709 -345 710 -344
rect 716 -345 717 -344
rect 12 -347 13 -346
rect 65 -347 66 -346
rect 68 -347 69 -346
rect 618 -347 619 -346
rect 23 -349 24 -348
rect 128 -349 129 -348
rect 142 -349 143 -348
rect 303 -349 304 -348
rect 313 -349 314 -348
rect 366 -349 367 -348
rect 467 -349 468 -348
rect 625 -349 626 -348
rect 30 -351 31 -350
rect 79 -351 80 -350
rect 89 -351 90 -350
rect 506 -351 507 -350
rect 548 -351 549 -350
rect 618 -351 619 -350
rect 37 -353 38 -352
rect 44 -353 45 -352
rect 51 -353 52 -352
rect 481 -353 482 -352
rect 506 -353 507 -352
rect 534 -353 535 -352
rect 597 -353 598 -352
rect 632 -353 633 -352
rect 37 -355 38 -354
rect 464 -355 465 -354
rect 471 -355 472 -354
rect 660 -355 661 -354
rect 44 -357 45 -356
rect 331 -357 332 -356
rect 338 -357 339 -356
rect 443 -357 444 -356
rect 450 -357 451 -356
rect 471 -357 472 -356
rect 72 -359 73 -358
rect 100 -359 101 -358
rect 117 -359 118 -358
rect 191 -359 192 -358
rect 198 -359 199 -358
rect 247 -359 248 -358
rect 282 -359 283 -358
rect 362 -359 363 -358
rect 390 -359 391 -358
rect 534 -359 535 -358
rect 75 -361 76 -360
rect 408 -361 409 -360
rect 411 -361 412 -360
rect 625 -361 626 -360
rect 79 -363 80 -362
rect 156 -363 157 -362
rect 163 -363 164 -362
rect 212 -363 213 -362
rect 226 -363 227 -362
rect 327 -363 328 -362
rect 355 -363 356 -362
rect 653 -363 654 -362
rect 86 -365 87 -364
rect 100 -365 101 -364
rect 107 -365 108 -364
rect 163 -365 164 -364
rect 177 -365 178 -364
rect 212 -365 213 -364
rect 219 -365 220 -364
rect 226 -365 227 -364
rect 233 -365 234 -364
rect 366 -365 367 -364
rect 390 -365 391 -364
rect 415 -365 416 -364
rect 443 -365 444 -364
rect 485 -365 486 -364
rect 590 -365 591 -364
rect 653 -365 654 -364
rect 86 -367 87 -366
rect 93 -367 94 -366
rect 110 -367 111 -366
rect 219 -367 220 -366
rect 233 -367 234 -366
rect 268 -367 269 -366
rect 282 -367 283 -366
rect 341 -367 342 -366
rect 359 -367 360 -366
rect 583 -367 584 -366
rect 590 -367 591 -366
rect 611 -367 612 -366
rect 58 -369 59 -368
rect 359 -369 360 -368
rect 394 -369 395 -368
rect 415 -369 416 -368
rect 450 -369 451 -368
rect 478 -369 479 -368
rect 485 -369 486 -368
rect 513 -369 514 -368
rect 583 -369 584 -368
rect 635 -369 636 -368
rect 58 -371 59 -370
rect 156 -371 157 -370
rect 201 -371 202 -370
rect 205 -371 206 -370
rect 247 -371 248 -370
rect 254 -371 255 -370
rect 268 -371 269 -370
rect 310 -371 311 -370
rect 317 -371 318 -370
rect 380 -371 381 -370
rect 457 -371 458 -370
rect 548 -371 549 -370
rect 121 -373 122 -372
rect 191 -373 192 -372
rect 254 -373 255 -372
rect 383 -373 384 -372
rect 457 -373 458 -372
rect 520 -373 521 -372
rect 121 -375 122 -374
rect 422 -375 423 -374
rect 492 -375 493 -374
rect 513 -375 514 -374
rect 128 -377 129 -376
rect 170 -377 171 -376
rect 187 -377 188 -376
rect 205 -377 206 -376
rect 296 -377 297 -376
rect 310 -377 311 -376
rect 324 -377 325 -376
rect 674 -377 675 -376
rect 114 -379 115 -378
rect 296 -379 297 -378
rect 303 -379 304 -378
rect 345 -379 346 -378
rect 352 -379 353 -378
rect 520 -379 521 -378
rect 135 -381 136 -380
rect 177 -381 178 -380
rect 334 -381 335 -380
rect 394 -381 395 -380
rect 422 -381 423 -380
rect 527 -381 528 -380
rect 135 -383 136 -382
rect 289 -383 290 -382
rect 345 -383 346 -382
rect 373 -383 374 -382
rect 380 -383 381 -382
rect 646 -383 647 -382
rect 142 -385 143 -384
rect 149 -385 150 -384
rect 170 -385 171 -384
rect 261 -385 262 -384
rect 289 -385 290 -384
rect 429 -385 430 -384
rect 492 -385 493 -384
rect 639 -385 640 -384
rect 93 -387 94 -386
rect 149 -387 150 -386
rect 261 -387 262 -386
rect 387 -387 388 -386
rect 495 -387 496 -386
rect 527 -387 528 -386
rect 562 -387 563 -386
rect 646 -387 647 -386
rect 355 -389 356 -388
rect 611 -389 612 -388
rect 373 -391 374 -390
rect 576 -391 577 -390
rect 604 -391 605 -390
rect 639 -391 640 -390
rect 541 -393 542 -392
rect 576 -393 577 -392
rect 604 -393 605 -392
rect 667 -393 668 -392
rect 243 -395 244 -394
rect 541 -395 542 -394
rect 562 -395 563 -394
rect 569 -395 570 -394
rect 324 -397 325 -396
rect 569 -397 570 -396
rect 401 -399 402 -398
rect 667 -399 668 -398
rect 401 -401 402 -400
rect 499 -401 500 -400
rect 9 -412 10 -411
rect 96 -412 97 -411
rect 100 -412 101 -411
rect 194 -412 195 -411
rect 198 -412 199 -411
rect 243 -412 244 -411
rect 268 -412 269 -411
rect 373 -412 374 -411
rect 383 -412 384 -411
rect 527 -412 528 -411
rect 562 -412 563 -411
rect 653 -412 654 -411
rect 656 -412 657 -411
rect 660 -412 661 -411
rect 716 -412 717 -411
rect 730 -412 731 -411
rect 16 -414 17 -413
rect 79 -414 80 -413
rect 93 -414 94 -413
rect 422 -414 423 -413
rect 425 -414 426 -413
rect 576 -414 577 -413
rect 597 -414 598 -413
rect 681 -414 682 -413
rect 23 -416 24 -415
rect 82 -416 83 -415
rect 114 -416 115 -415
rect 170 -416 171 -415
rect 180 -416 181 -415
rect 639 -416 640 -415
rect 30 -418 31 -417
rect 103 -418 104 -417
rect 121 -418 122 -417
rect 576 -418 577 -417
rect 583 -418 584 -417
rect 639 -418 640 -417
rect 37 -420 38 -419
rect 110 -420 111 -419
rect 156 -420 157 -419
rect 240 -420 241 -419
rect 247 -420 248 -419
rect 268 -420 269 -419
rect 282 -420 283 -419
rect 520 -420 521 -419
rect 534 -420 535 -419
rect 562 -420 563 -419
rect 569 -420 570 -419
rect 723 -420 724 -419
rect 37 -422 38 -421
rect 51 -422 52 -421
rect 58 -422 59 -421
rect 352 -422 353 -421
rect 373 -422 374 -421
rect 422 -422 423 -421
rect 432 -422 433 -421
rect 499 -422 500 -421
rect 513 -422 514 -421
rect 569 -422 570 -421
rect 604 -422 605 -421
rect 702 -422 703 -421
rect 44 -424 45 -423
rect 93 -424 94 -423
rect 100 -424 101 -423
rect 121 -424 122 -423
rect 135 -424 136 -423
rect 240 -424 241 -423
rect 303 -424 304 -423
rect 352 -424 353 -423
rect 387 -424 388 -423
rect 453 -424 454 -423
rect 464 -424 465 -423
rect 597 -424 598 -423
rect 611 -424 612 -423
rect 688 -424 689 -423
rect 44 -426 45 -425
rect 142 -426 143 -425
rect 163 -426 164 -425
rect 338 -426 339 -425
rect 390 -426 391 -425
rect 618 -426 619 -425
rect 625 -426 626 -425
rect 674 -426 675 -425
rect 58 -428 59 -427
rect 128 -428 129 -427
rect 135 -428 136 -427
rect 205 -428 206 -427
rect 219 -428 220 -427
rect 226 -428 227 -427
rect 233 -428 234 -427
rect 282 -428 283 -427
rect 296 -428 297 -427
rect 387 -428 388 -427
rect 390 -428 391 -427
rect 527 -428 528 -427
rect 541 -428 542 -427
rect 583 -428 584 -427
rect 65 -430 66 -429
rect 107 -430 108 -429
rect 149 -430 150 -429
rect 205 -430 206 -429
rect 212 -430 213 -429
rect 233 -430 234 -429
rect 313 -430 314 -429
rect 464 -430 465 -429
rect 481 -430 482 -429
rect 632 -430 633 -429
rect 68 -432 69 -431
rect 541 -432 542 -431
rect 555 -432 556 -431
rect 604 -432 605 -431
rect 72 -434 73 -433
rect 124 -434 125 -433
rect 149 -434 150 -433
rect 285 -434 286 -433
rect 324 -434 325 -433
rect 359 -434 360 -433
rect 401 -434 402 -433
rect 534 -434 535 -433
rect 72 -436 73 -435
rect 380 -436 381 -435
rect 408 -436 409 -435
rect 646 -436 647 -435
rect 86 -438 87 -437
rect 247 -438 248 -437
rect 327 -438 328 -437
rect 548 -438 549 -437
rect 590 -438 591 -437
rect 646 -438 647 -437
rect 86 -440 87 -439
rect 254 -440 255 -439
rect 331 -440 332 -439
rect 446 -440 447 -439
rect 450 -440 451 -439
rect 513 -440 514 -439
rect 170 -442 171 -441
rect 303 -442 304 -441
rect 345 -442 346 -441
rect 380 -442 381 -441
rect 411 -442 412 -441
rect 590 -442 591 -441
rect 177 -444 178 -443
rect 212 -444 213 -443
rect 254 -444 255 -443
rect 317 -444 318 -443
rect 359 -444 360 -443
rect 418 -444 419 -443
rect 436 -444 437 -443
rect 548 -444 549 -443
rect 128 -446 129 -445
rect 177 -446 178 -445
rect 184 -446 185 -445
rect 289 -446 290 -445
rect 310 -446 311 -445
rect 345 -446 346 -445
rect 366 -446 367 -445
rect 401 -446 402 -445
rect 436 -446 437 -445
rect 625 -446 626 -445
rect 184 -448 185 -447
rect 219 -448 220 -447
rect 229 -448 230 -447
rect 317 -448 318 -447
rect 439 -448 440 -447
rect 709 -448 710 -447
rect 191 -450 192 -449
rect 296 -450 297 -449
rect 443 -450 444 -449
rect 520 -450 521 -449
rect 51 -452 52 -451
rect 191 -452 192 -451
rect 198 -452 199 -451
rect 261 -452 262 -451
rect 289 -452 290 -451
rect 394 -452 395 -451
rect 492 -452 493 -451
rect 695 -452 696 -451
rect 166 -454 167 -453
rect 261 -454 262 -453
rect 394 -454 395 -453
rect 457 -454 458 -453
rect 485 -454 486 -453
rect 492 -454 493 -453
rect 502 -454 503 -453
rect 611 -454 612 -453
rect 341 -456 342 -455
rect 457 -456 458 -455
rect 506 -456 507 -455
rect 555 -456 556 -455
rect 366 -458 367 -457
rect 485 -458 486 -457
rect 471 -460 472 -459
rect 506 -460 507 -459
rect 471 -462 472 -461
rect 667 -462 668 -461
rect 478 -464 479 -463
rect 667 -464 668 -463
rect 415 -466 416 -465
rect 478 -466 479 -465
rect 58 -477 59 -476
rect 163 -477 164 -476
rect 177 -477 178 -476
rect 604 -477 605 -476
rect 639 -477 640 -476
rect 709 -477 710 -476
rect 716 -477 717 -476
rect 730 -477 731 -476
rect 75 -479 76 -478
rect 744 -479 745 -478
rect 23 -481 24 -480
rect 75 -481 76 -480
rect 79 -481 80 -480
rect 737 -481 738 -480
rect 79 -483 80 -482
rect 135 -483 136 -482
rect 145 -483 146 -482
rect 695 -483 696 -482
rect 723 -483 724 -482
rect 779 -483 780 -482
rect 93 -485 94 -484
rect 145 -485 146 -484
rect 152 -485 153 -484
rect 205 -485 206 -484
rect 219 -485 220 -484
rect 222 -485 223 -484
rect 243 -485 244 -484
rect 345 -485 346 -484
rect 359 -485 360 -484
rect 618 -485 619 -484
rect 646 -485 647 -484
rect 723 -485 724 -484
rect 37 -487 38 -486
rect 93 -487 94 -486
rect 121 -487 122 -486
rect 191 -487 192 -486
rect 219 -487 220 -486
rect 254 -487 255 -486
rect 289 -487 290 -486
rect 450 -487 451 -486
rect 555 -487 556 -486
rect 604 -487 605 -486
rect 674 -487 675 -486
rect 716 -487 717 -486
rect 121 -489 122 -488
rect 268 -489 269 -488
rect 289 -489 290 -488
rect 331 -489 332 -488
rect 345 -489 346 -488
rect 373 -489 374 -488
rect 383 -489 384 -488
rect 415 -489 416 -488
rect 422 -489 423 -488
rect 639 -489 640 -488
rect 51 -491 52 -490
rect 331 -491 332 -490
rect 352 -491 353 -490
rect 359 -491 360 -490
rect 366 -491 367 -490
rect 548 -491 549 -490
rect 555 -491 556 -490
rect 590 -491 591 -490
rect 597 -491 598 -490
rect 660 -491 661 -490
rect 16 -493 17 -492
rect 590 -493 591 -492
rect 30 -495 31 -494
rect 51 -495 52 -494
rect 124 -495 125 -494
rect 695 -495 696 -494
rect 128 -497 129 -496
rect 268 -497 269 -496
rect 390 -497 391 -496
rect 611 -497 612 -496
rect 107 -499 108 -498
rect 128 -499 129 -498
rect 135 -499 136 -498
rect 719 -499 720 -498
rect 44 -501 45 -500
rect 107 -501 108 -500
rect 149 -501 150 -500
rect 205 -501 206 -500
rect 222 -501 223 -500
rect 254 -501 255 -500
rect 394 -501 395 -500
rect 751 -501 752 -500
rect 44 -503 45 -502
rect 114 -503 115 -502
rect 180 -503 181 -502
rect 212 -503 213 -502
rect 408 -503 409 -502
rect 436 -503 437 -502
rect 439 -503 440 -502
rect 681 -503 682 -502
rect 61 -505 62 -504
rect 114 -505 115 -504
rect 187 -505 188 -504
rect 338 -505 339 -504
rect 401 -505 402 -504
rect 408 -505 409 -504
rect 411 -505 412 -504
rect 478 -505 479 -504
rect 513 -505 514 -504
rect 548 -505 549 -504
rect 562 -505 563 -504
rect 611 -505 612 -504
rect 625 -505 626 -504
rect 681 -505 682 -504
rect 65 -507 66 -506
rect 625 -507 626 -506
rect 170 -509 171 -508
rect 562 -509 563 -508
rect 576 -509 577 -508
rect 646 -509 647 -508
rect 170 -511 171 -510
rect 282 -511 283 -510
rect 303 -511 304 -510
rect 338 -511 339 -510
rect 429 -511 430 -510
rect 653 -511 654 -510
rect 191 -513 192 -512
rect 310 -513 311 -512
rect 324 -513 325 -512
rect 401 -513 402 -512
rect 432 -513 433 -512
rect 597 -513 598 -512
rect 142 -515 143 -514
rect 310 -515 311 -514
rect 317 -515 318 -514
rect 324 -515 325 -514
rect 432 -515 433 -514
rect 667 -515 668 -514
rect 212 -517 213 -516
rect 296 -517 297 -516
rect 303 -517 304 -516
rect 730 -517 731 -516
rect 226 -519 227 -518
rect 317 -519 318 -518
rect 397 -519 398 -518
rect 667 -519 668 -518
rect 226 -521 227 -520
rect 233 -521 234 -520
rect 240 -521 241 -520
rect 296 -521 297 -520
rect 443 -521 444 -520
rect 702 -521 703 -520
rect 233 -523 234 -522
rect 352 -523 353 -522
rect 387 -523 388 -522
rect 702 -523 703 -522
rect 240 -525 241 -524
rect 373 -525 374 -524
rect 443 -525 444 -524
rect 688 -525 689 -524
rect 261 -527 262 -526
rect 387 -527 388 -526
rect 478 -527 479 -526
rect 527 -527 528 -526
rect 534 -527 535 -526
rect 576 -527 577 -526
rect 583 -527 584 -526
rect 653 -527 654 -526
rect 282 -529 283 -528
rect 369 -529 370 -528
rect 453 -529 454 -528
rect 534 -529 535 -528
rect 632 -529 633 -528
rect 688 -529 689 -528
rect 9 -531 10 -530
rect 632 -531 633 -530
rect 492 -533 493 -532
rect 583 -533 584 -532
rect 446 -535 447 -534
rect 492 -535 493 -534
rect 506 -535 507 -534
rect 527 -535 528 -534
rect 261 -537 262 -536
rect 446 -537 447 -536
rect 513 -537 514 -536
rect 541 -537 542 -536
rect 320 -539 321 -538
rect 506 -539 507 -538
rect 520 -539 521 -538
rect 674 -539 675 -538
rect 499 -541 500 -540
rect 520 -541 521 -540
rect 541 -541 542 -540
rect 569 -541 570 -540
rect 464 -543 465 -542
rect 569 -543 570 -542
rect 457 -545 458 -544
rect 464 -545 465 -544
rect 485 -545 486 -544
rect 499 -545 500 -544
rect 86 -547 87 -546
rect 457 -547 458 -546
rect 471 -547 472 -546
rect 485 -547 486 -546
rect 68 -549 69 -548
rect 471 -549 472 -548
rect 26 -551 27 -550
rect 68 -551 69 -550
rect 86 -551 87 -550
rect 163 -551 164 -550
rect 16 -562 17 -561
rect 408 -562 409 -561
rect 418 -562 419 -561
rect 723 -562 724 -561
rect 779 -562 780 -561
rect 807 -562 808 -561
rect 23 -564 24 -563
rect 54 -564 55 -563
rect 58 -564 59 -563
rect 135 -564 136 -563
rect 156 -564 157 -563
rect 177 -564 178 -563
rect 187 -564 188 -563
rect 282 -564 283 -563
rect 306 -564 307 -563
rect 324 -564 325 -563
rect 355 -564 356 -563
rect 520 -564 521 -563
rect 541 -564 542 -563
rect 544 -564 545 -563
rect 23 -566 24 -565
rect 124 -566 125 -565
rect 128 -566 129 -565
rect 156 -566 157 -565
rect 166 -566 167 -565
rect 674 -566 675 -565
rect 30 -568 31 -567
rect 96 -568 97 -567
rect 100 -568 101 -567
rect 149 -568 150 -567
rect 177 -568 178 -567
rect 187 -568 188 -567
rect 205 -568 206 -567
rect 215 -568 216 -567
rect 219 -568 220 -567
rect 317 -568 318 -567
rect 366 -568 367 -567
rect 499 -568 500 -567
rect 541 -568 542 -567
rect 576 -568 577 -567
rect 33 -570 34 -569
rect 51 -570 52 -569
rect 61 -570 62 -569
rect 625 -570 626 -569
rect 44 -572 45 -571
rect 128 -572 129 -571
rect 191 -572 192 -571
rect 317 -572 318 -571
rect 369 -572 370 -571
rect 674 -572 675 -571
rect 47 -574 48 -573
rect 653 -574 654 -573
rect 51 -576 52 -575
rect 366 -576 367 -575
rect 394 -576 395 -575
rect 646 -576 647 -575
rect 65 -578 66 -577
rect 397 -578 398 -577
rect 411 -578 412 -577
rect 499 -578 500 -577
rect 544 -578 545 -577
rect 576 -578 577 -577
rect 625 -578 626 -577
rect 688 -578 689 -577
rect 65 -580 66 -579
rect 352 -580 353 -579
rect 394 -580 395 -579
rect 751 -580 752 -579
rect 72 -582 73 -581
rect 590 -582 591 -581
rect 646 -582 647 -581
rect 695 -582 696 -581
rect 72 -584 73 -583
rect 142 -584 143 -583
rect 191 -584 192 -583
rect 198 -584 199 -583
rect 212 -584 213 -583
rect 723 -584 724 -583
rect 107 -586 108 -585
rect 184 -586 185 -585
rect 212 -586 213 -585
rect 401 -586 402 -585
rect 425 -586 426 -585
rect 534 -586 535 -585
rect 590 -586 591 -585
rect 639 -586 640 -585
rect 688 -586 689 -585
rect 730 -586 731 -585
rect 114 -588 115 -587
rect 135 -588 136 -587
rect 219 -588 220 -587
rect 310 -588 311 -587
rect 338 -588 339 -587
rect 369 -588 370 -587
rect 401 -588 402 -587
rect 415 -588 416 -587
rect 429 -588 430 -587
rect 569 -588 570 -587
rect 597 -588 598 -587
rect 695 -588 696 -587
rect 730 -588 731 -587
rect 737 -588 738 -587
rect 226 -590 227 -589
rect 520 -590 521 -589
rect 569 -590 570 -589
rect 604 -590 605 -589
rect 226 -592 227 -591
rect 261 -592 262 -591
rect 275 -592 276 -591
rect 278 -592 279 -591
rect 282 -592 283 -591
rect 296 -592 297 -591
rect 310 -592 311 -591
rect 450 -592 451 -591
rect 471 -592 472 -591
rect 737 -592 738 -591
rect 233 -594 234 -593
rect 296 -594 297 -593
rect 331 -594 332 -593
rect 415 -594 416 -593
rect 429 -594 430 -593
rect 464 -594 465 -593
rect 471 -594 472 -593
rect 492 -594 493 -593
rect 604 -594 605 -593
rect 660 -594 661 -593
rect 163 -596 164 -595
rect 660 -596 661 -595
rect 233 -598 234 -597
rect 254 -598 255 -597
rect 261 -598 262 -597
rect 387 -598 388 -597
rect 432 -598 433 -597
rect 709 -598 710 -597
rect 142 -600 143 -599
rect 709 -600 710 -599
rect 184 -602 185 -601
rect 254 -602 255 -601
rect 275 -602 276 -601
rect 653 -602 654 -601
rect 236 -604 237 -603
rect 744 -604 745 -603
rect 240 -606 241 -605
rect 247 -606 248 -605
rect 289 -606 290 -605
rect 324 -606 325 -605
rect 331 -606 332 -605
rect 373 -606 374 -605
rect 387 -606 388 -605
rect 667 -606 668 -605
rect 79 -608 80 -607
rect 240 -608 241 -607
rect 247 -608 248 -607
rect 268 -608 269 -607
rect 303 -608 304 -607
rect 373 -608 374 -607
rect 390 -608 391 -607
rect 667 -608 668 -607
rect 79 -610 80 -609
rect 170 -610 171 -609
rect 198 -610 199 -609
rect 289 -610 290 -609
rect 303 -610 304 -609
rect 345 -610 346 -609
rect 348 -610 349 -609
rect 597 -610 598 -609
rect 86 -612 87 -611
rect 170 -612 171 -611
rect 268 -612 269 -611
rect 292 -612 293 -611
rect 338 -612 339 -611
rect 457 -612 458 -611
rect 464 -612 465 -611
rect 555 -612 556 -611
rect 86 -614 87 -613
rect 103 -614 104 -613
rect 320 -614 321 -613
rect 457 -614 458 -613
rect 478 -614 479 -613
rect 534 -614 535 -613
rect 555 -614 556 -613
rect 716 -614 717 -613
rect 93 -616 94 -615
rect 345 -616 346 -615
rect 352 -616 353 -615
rect 618 -616 619 -615
rect 93 -618 94 -617
rect 205 -618 206 -617
rect 383 -618 384 -617
rect 618 -618 619 -617
rect 443 -620 444 -619
rect 611 -620 612 -619
rect 446 -622 447 -621
rect 702 -622 703 -621
rect 446 -624 447 -623
rect 639 -624 640 -623
rect 450 -626 451 -625
rect 548 -626 549 -625
rect 485 -628 486 -627
rect 611 -628 612 -627
rect 485 -630 486 -629
rect 506 -630 507 -629
rect 513 -630 514 -629
rect 702 -630 703 -629
rect 478 -632 479 -631
rect 513 -632 514 -631
rect 516 -632 517 -631
rect 716 -632 717 -631
rect 506 -634 507 -633
rect 527 -634 528 -633
rect 548 -634 549 -633
rect 583 -634 584 -633
rect 380 -636 381 -635
rect 527 -636 528 -635
rect 583 -636 584 -635
rect 632 -636 633 -635
rect 359 -638 360 -637
rect 380 -638 381 -637
rect 632 -638 633 -637
rect 681 -638 682 -637
rect 359 -640 360 -639
rect 436 -640 437 -639
rect 75 -642 76 -641
rect 436 -642 437 -641
rect 425 -644 426 -643
rect 681 -644 682 -643
rect 58 -655 59 -654
rect 96 -655 97 -654
rect 100 -655 101 -654
rect 114 -655 115 -654
rect 117 -655 118 -654
rect 156 -655 157 -654
rect 166 -655 167 -654
rect 177 -655 178 -654
rect 184 -655 185 -654
rect 240 -655 241 -654
rect 254 -655 255 -654
rect 345 -655 346 -654
rect 348 -655 349 -654
rect 450 -655 451 -654
rect 474 -655 475 -654
rect 765 -655 766 -654
rect 807 -655 808 -654
rect 828 -655 829 -654
rect 9 -657 10 -656
rect 114 -657 115 -656
rect 117 -657 118 -656
rect 198 -657 199 -656
rect 212 -657 213 -656
rect 254 -657 255 -656
rect 261 -657 262 -656
rect 278 -657 279 -656
rect 282 -657 283 -656
rect 289 -657 290 -656
rect 352 -657 353 -656
rect 415 -657 416 -656
rect 418 -657 419 -656
rect 513 -657 514 -656
rect 555 -657 556 -656
rect 772 -657 773 -656
rect 16 -659 17 -658
rect 352 -659 353 -658
rect 366 -659 367 -658
rect 534 -659 535 -658
rect 597 -659 598 -658
rect 824 -659 825 -658
rect 16 -661 17 -660
rect 72 -661 73 -660
rect 86 -661 87 -660
rect 121 -661 122 -660
rect 124 -661 125 -660
rect 432 -661 433 -660
rect 443 -661 444 -660
rect 555 -661 556 -660
rect 660 -661 661 -660
rect 695 -661 696 -660
rect 709 -661 710 -660
rect 786 -661 787 -660
rect 51 -663 52 -662
rect 100 -663 101 -662
rect 107 -663 108 -662
rect 583 -663 584 -662
rect 646 -663 647 -662
rect 695 -663 696 -662
rect 716 -663 717 -662
rect 793 -663 794 -662
rect 58 -665 59 -664
rect 800 -665 801 -664
rect 65 -667 66 -666
rect 149 -667 150 -666
rect 152 -667 153 -666
rect 243 -667 244 -666
rect 261 -667 262 -666
rect 289 -667 290 -666
rect 380 -667 381 -666
rect 387 -667 388 -666
rect 408 -667 409 -666
rect 611 -667 612 -666
rect 667 -667 668 -666
rect 709 -667 710 -666
rect 730 -667 731 -666
rect 758 -667 759 -666
rect 23 -669 24 -668
rect 65 -669 66 -668
rect 86 -669 87 -668
rect 310 -669 311 -668
rect 411 -669 412 -668
rect 807 -669 808 -668
rect 23 -671 24 -670
rect 257 -671 258 -670
rect 303 -671 304 -670
rect 380 -671 381 -670
rect 422 -671 423 -670
rect 702 -671 703 -670
rect 30 -673 31 -672
rect 411 -673 412 -672
rect 429 -673 430 -672
rect 492 -673 493 -672
rect 590 -673 591 -672
rect 611 -673 612 -672
rect 618 -673 619 -672
rect 702 -673 703 -672
rect 37 -675 38 -674
rect 408 -675 409 -674
rect 443 -675 444 -674
rect 478 -675 479 -674
rect 548 -675 549 -674
rect 590 -675 591 -674
rect 604 -675 605 -674
rect 618 -675 619 -674
rect 653 -675 654 -674
rect 667 -675 668 -674
rect 674 -675 675 -674
rect 751 -675 752 -674
rect 44 -677 45 -676
rect 653 -677 654 -676
rect 681 -677 682 -676
rect 716 -677 717 -676
rect 44 -679 45 -678
rect 93 -679 94 -678
rect 107 -679 108 -678
rect 163 -679 164 -678
rect 177 -679 178 -678
rect 401 -679 402 -678
rect 439 -679 440 -678
rect 548 -679 549 -678
rect 576 -679 577 -678
rect 604 -679 605 -678
rect 681 -679 682 -678
rect 723 -679 724 -678
rect 79 -681 80 -680
rect 303 -681 304 -680
rect 310 -681 311 -680
rect 338 -681 339 -680
rect 394 -681 395 -680
rect 422 -681 423 -680
rect 457 -681 458 -680
rect 646 -681 647 -680
rect 688 -681 689 -680
rect 779 -681 780 -680
rect 79 -683 80 -682
rect 390 -683 391 -682
rect 397 -683 398 -682
rect 576 -683 577 -682
rect 632 -683 633 -682
rect 723 -683 724 -682
rect 121 -685 122 -684
rect 527 -685 528 -684
rect 625 -685 626 -684
rect 632 -685 633 -684
rect 639 -685 640 -684
rect 688 -685 689 -684
rect 128 -687 129 -686
rect 268 -687 269 -686
rect 282 -687 283 -686
rect 394 -687 395 -686
rect 467 -687 468 -686
rect 478 -687 479 -686
rect 499 -687 500 -686
rect 639 -687 640 -686
rect 131 -689 132 -688
rect 541 -689 542 -688
rect 569 -689 570 -688
rect 625 -689 626 -688
rect 135 -691 136 -690
rect 212 -691 213 -690
rect 219 -691 220 -690
rect 338 -691 339 -690
rect 359 -691 360 -690
rect 457 -691 458 -690
rect 471 -691 472 -690
rect 534 -691 535 -690
rect 124 -693 125 -692
rect 219 -693 220 -692
rect 226 -693 227 -692
rect 268 -693 269 -692
rect 292 -693 293 -692
rect 674 -693 675 -692
rect 110 -695 111 -694
rect 226 -695 227 -694
rect 236 -695 237 -694
rect 744 -695 745 -694
rect 135 -697 136 -696
rect 145 -697 146 -696
rect 156 -697 157 -696
rect 317 -697 318 -696
rect 331 -697 332 -696
rect 401 -697 402 -696
rect 436 -697 437 -696
rect 499 -697 500 -696
rect 506 -697 507 -696
rect 541 -697 542 -696
rect 142 -699 143 -698
rect 485 -699 486 -698
rect 506 -699 507 -698
rect 737 -699 738 -698
rect 47 -701 48 -700
rect 142 -701 143 -700
rect 163 -701 164 -700
rect 562 -701 563 -700
rect 166 -703 167 -702
rect 562 -703 563 -702
rect 184 -705 185 -704
rect 275 -705 276 -704
rect 296 -705 297 -704
rect 359 -705 360 -704
rect 369 -705 370 -704
rect 737 -705 738 -704
rect 173 -707 174 -706
rect 296 -707 297 -706
rect 317 -707 318 -706
rect 814 -707 815 -706
rect 198 -709 199 -708
rect 247 -709 248 -708
rect 324 -709 325 -708
rect 369 -709 370 -708
rect 446 -709 447 -708
rect 485 -709 486 -708
rect 205 -711 206 -710
rect 583 -711 584 -710
rect 170 -713 171 -712
rect 205 -713 206 -712
rect 233 -713 234 -712
rect 275 -713 276 -712
rect 324 -713 325 -712
rect 373 -713 374 -712
rect 233 -715 234 -714
rect 520 -715 521 -714
rect 240 -717 241 -716
rect 730 -717 731 -716
rect 247 -719 248 -718
rect 429 -719 430 -718
rect 464 -719 465 -718
rect 520 -719 521 -718
rect 331 -721 332 -720
rect 527 -721 528 -720
rect 334 -723 335 -722
rect 569 -723 570 -722
rect 373 -725 374 -724
rect 436 -725 437 -724
rect 40 -736 41 -735
rect 121 -736 122 -735
rect 124 -736 125 -735
rect 730 -736 731 -735
rect 817 -736 818 -735
rect 828 -736 829 -735
rect 44 -738 45 -737
rect 68 -738 69 -737
rect 72 -738 73 -737
rect 212 -738 213 -737
rect 236 -738 237 -737
rect 464 -738 465 -737
rect 467 -738 468 -737
rect 793 -738 794 -737
rect 47 -740 48 -739
rect 65 -740 66 -739
rect 72 -740 73 -739
rect 306 -740 307 -739
rect 324 -740 325 -739
rect 464 -740 465 -739
rect 474 -740 475 -739
rect 779 -740 780 -739
rect 51 -742 52 -741
rect 583 -742 584 -741
rect 597 -742 598 -741
rect 632 -742 633 -741
rect 639 -742 640 -741
rect 814 -742 815 -741
rect 58 -744 59 -743
rect 653 -744 654 -743
rect 681 -744 682 -743
rect 779 -744 780 -743
rect 58 -746 59 -745
rect 338 -746 339 -745
rect 341 -746 342 -745
rect 807 -746 808 -745
rect 75 -748 76 -747
rect 653 -748 654 -747
rect 660 -748 661 -747
rect 681 -748 682 -747
rect 96 -750 97 -749
rect 660 -750 661 -749
rect 117 -752 118 -751
rect 702 -752 703 -751
rect 142 -754 143 -753
rect 212 -754 213 -753
rect 240 -754 241 -753
rect 824 -754 825 -753
rect 79 -756 80 -755
rect 240 -756 241 -755
rect 254 -756 255 -755
rect 268 -756 269 -755
rect 289 -756 290 -755
rect 765 -756 766 -755
rect 86 -758 87 -757
rect 268 -758 269 -757
rect 282 -758 283 -757
rect 289 -758 290 -757
rect 292 -758 293 -757
rect 485 -758 486 -757
rect 506 -758 507 -757
rect 730 -758 731 -757
rect 86 -760 87 -759
rect 233 -760 234 -759
rect 275 -760 276 -759
rect 282 -760 283 -759
rect 310 -760 311 -759
rect 506 -760 507 -759
rect 583 -760 584 -759
rect 688 -760 689 -759
rect 37 -762 38 -761
rect 310 -762 311 -761
rect 324 -762 325 -761
rect 345 -762 346 -761
rect 348 -762 349 -761
rect 793 -762 794 -761
rect 37 -764 38 -763
rect 800 -764 801 -763
rect 107 -766 108 -765
rect 233 -766 234 -765
rect 331 -766 332 -765
rect 352 -766 353 -765
rect 366 -766 367 -765
rect 702 -766 703 -765
rect 107 -768 108 -767
rect 471 -768 472 -767
rect 548 -768 549 -767
rect 688 -768 689 -767
rect 82 -770 83 -769
rect 548 -770 549 -769
rect 590 -770 591 -769
rect 765 -770 766 -769
rect 135 -772 136 -771
rect 275 -772 276 -771
rect 296 -772 297 -771
rect 331 -772 332 -771
rect 352 -772 353 -771
rect 369 -772 370 -771
rect 394 -772 395 -771
rect 492 -772 493 -771
rect 600 -772 601 -771
rect 751 -772 752 -771
rect 135 -774 136 -773
rect 366 -774 367 -773
rect 387 -774 388 -773
rect 394 -774 395 -773
rect 408 -774 409 -773
rect 443 -774 444 -773
rect 450 -774 451 -773
rect 674 -774 675 -773
rect 709 -774 710 -773
rect 751 -774 752 -773
rect 142 -776 143 -775
rect 184 -776 185 -775
rect 226 -776 227 -775
rect 345 -776 346 -775
rect 408 -776 409 -775
rect 415 -776 416 -775
rect 429 -776 430 -775
rect 520 -776 521 -775
rect 632 -776 633 -775
rect 667 -776 668 -775
rect 159 -778 160 -777
rect 772 -778 773 -777
rect 163 -780 164 -779
rect 401 -780 402 -779
rect 411 -780 412 -779
rect 625 -780 626 -779
rect 639 -780 640 -779
rect 737 -780 738 -779
rect 170 -782 171 -781
rect 205 -782 206 -781
rect 296 -782 297 -781
rect 439 -782 440 -781
rect 446 -782 447 -781
rect 674 -782 675 -781
rect 198 -784 199 -783
rect 226 -784 227 -783
rect 380 -784 381 -783
rect 415 -784 416 -783
rect 436 -784 437 -783
rect 723 -784 724 -783
rect 16 -786 17 -785
rect 723 -786 724 -785
rect 198 -788 199 -787
rect 373 -788 374 -787
rect 380 -788 381 -787
rect 744 -788 745 -787
rect 205 -790 206 -789
rect 247 -790 248 -789
rect 359 -790 360 -789
rect 373 -790 374 -789
rect 404 -790 405 -789
rect 737 -790 738 -789
rect 23 -792 24 -791
rect 247 -792 248 -791
rect 338 -792 339 -791
rect 359 -792 360 -791
rect 436 -792 437 -791
rect 744 -792 745 -791
rect 23 -794 24 -793
rect 156 -794 157 -793
rect 457 -794 458 -793
rect 485 -794 486 -793
rect 492 -794 493 -793
rect 541 -794 542 -793
rect 604 -794 605 -793
rect 667 -794 668 -793
rect 93 -796 94 -795
rect 156 -796 157 -795
rect 422 -796 423 -795
rect 457 -796 458 -795
rect 471 -796 472 -795
rect 513 -796 514 -795
rect 520 -796 521 -795
rect 576 -796 577 -795
rect 625 -796 626 -795
rect 695 -796 696 -795
rect 93 -798 94 -797
rect 261 -798 262 -797
rect 453 -798 454 -797
rect 513 -798 514 -797
rect 534 -798 535 -797
rect 541 -798 542 -797
rect 562 -798 563 -797
rect 576 -798 577 -797
rect 618 -798 619 -797
rect 695 -798 696 -797
rect 16 -800 17 -799
rect 562 -800 563 -799
rect 569 -800 570 -799
rect 604 -800 605 -799
rect 646 -800 647 -799
rect 709 -800 710 -799
rect 149 -802 150 -801
rect 422 -802 423 -801
rect 499 -802 500 -801
rect 772 -802 773 -801
rect 114 -804 115 -803
rect 149 -804 150 -803
rect 261 -804 262 -803
rect 387 -804 388 -803
rect 478 -804 479 -803
rect 499 -804 500 -803
rect 527 -804 528 -803
rect 534 -804 535 -803
rect 555 -804 556 -803
rect 569 -804 570 -803
rect 646 -804 647 -803
rect 821 -804 822 -803
rect 177 -806 178 -805
rect 527 -806 528 -805
rect 555 -806 556 -805
rect 786 -806 787 -805
rect 128 -808 129 -807
rect 177 -808 178 -807
rect 219 -808 220 -807
rect 478 -808 479 -807
rect 758 -808 759 -807
rect 786 -808 787 -807
rect 30 -810 31 -809
rect 128 -810 129 -809
rect 219 -810 220 -809
rect 317 -810 318 -809
rect 716 -810 717 -809
rect 758 -810 759 -809
rect 30 -812 31 -811
rect 187 -812 188 -811
rect 271 -812 272 -811
rect 618 -812 619 -811
rect 303 -814 304 -813
rect 317 -814 318 -813
rect 390 -814 391 -813
rect 716 -814 717 -813
rect 9 -825 10 -824
rect 93 -825 94 -824
rect 96 -825 97 -824
rect 240 -825 241 -824
rect 303 -825 304 -824
rect 772 -825 773 -824
rect 23 -827 24 -826
rect 51 -827 52 -826
rect 54 -827 55 -826
rect 362 -827 363 -826
rect 369 -827 370 -826
rect 709 -827 710 -826
rect 37 -829 38 -828
rect 723 -829 724 -828
rect 37 -831 38 -830
rect 285 -831 286 -830
rect 331 -831 332 -830
rect 744 -831 745 -830
rect 26 -833 27 -832
rect 331 -833 332 -832
rect 348 -833 349 -832
rect 527 -833 528 -832
rect 530 -833 531 -832
rect 779 -833 780 -832
rect 51 -835 52 -834
rect 212 -835 213 -834
rect 352 -835 353 -834
rect 730 -835 731 -834
rect 58 -837 59 -836
rect 240 -837 241 -836
rect 359 -837 360 -836
rect 383 -837 384 -836
rect 390 -837 391 -836
rect 765 -837 766 -836
rect 58 -839 59 -838
rect 191 -839 192 -838
rect 212 -839 213 -838
rect 254 -839 255 -838
rect 373 -839 374 -838
rect 387 -839 388 -838
rect 404 -839 405 -838
rect 569 -839 570 -838
rect 590 -839 591 -838
rect 688 -839 689 -838
rect 709 -839 710 -838
rect 758 -839 759 -838
rect 30 -841 31 -840
rect 191 -841 192 -840
rect 257 -841 258 -840
rect 373 -841 374 -840
rect 380 -841 381 -840
rect 576 -841 577 -840
rect 632 -841 633 -840
rect 635 -841 636 -840
rect 681 -841 682 -840
rect 758 -841 759 -840
rect 30 -843 31 -842
rect 100 -843 101 -842
rect 128 -843 129 -842
rect 184 -843 185 -842
rect 187 -843 188 -842
rect 282 -843 283 -842
rect 306 -843 307 -842
rect 688 -843 689 -842
rect 65 -845 66 -844
rect 653 -845 654 -844
rect 65 -847 66 -846
rect 68 -847 69 -846
rect 72 -847 73 -846
rect 107 -847 108 -846
rect 114 -847 115 -846
rect 128 -847 129 -846
rect 145 -847 146 -846
rect 737 -847 738 -846
rect 16 -849 17 -848
rect 114 -849 115 -848
rect 149 -849 150 -848
rect 317 -849 318 -848
rect 324 -849 325 -848
rect 387 -849 388 -848
rect 394 -849 395 -848
rect 404 -849 405 -848
rect 411 -849 412 -848
rect 702 -849 703 -848
rect 716 -849 717 -848
rect 737 -849 738 -848
rect 44 -851 45 -850
rect 702 -851 703 -850
rect 44 -853 45 -852
rect 247 -853 248 -852
rect 310 -853 311 -852
rect 324 -853 325 -852
rect 338 -853 339 -852
rect 576 -853 577 -852
rect 611 -853 612 -852
rect 681 -853 682 -852
rect 72 -855 73 -854
rect 198 -855 199 -854
rect 219 -855 220 -854
rect 310 -855 311 -854
rect 394 -855 395 -854
rect 408 -855 409 -854
rect 422 -855 423 -854
rect 653 -855 654 -854
rect 82 -857 83 -856
rect 506 -857 507 -856
rect 537 -857 538 -856
rect 695 -857 696 -856
rect 86 -859 87 -858
rect 198 -859 199 -858
rect 226 -859 227 -858
rect 247 -859 248 -858
rect 422 -859 423 -858
rect 562 -859 563 -858
rect 569 -859 570 -858
rect 667 -859 668 -858
rect 86 -861 87 -860
rect 121 -861 122 -860
rect 149 -861 150 -860
rect 261 -861 262 -860
rect 429 -861 430 -860
rect 485 -861 486 -860
rect 555 -861 556 -860
rect 793 -861 794 -860
rect 93 -863 94 -862
rect 142 -863 143 -862
rect 152 -863 153 -862
rect 275 -863 276 -862
rect 299 -863 300 -862
rect 429 -863 430 -862
rect 436 -863 437 -862
rect 520 -863 521 -862
rect 555 -863 556 -862
rect 618 -863 619 -862
rect 632 -863 633 -862
rect 639 -863 640 -862
rect 667 -863 668 -862
rect 751 -863 752 -862
rect 107 -865 108 -864
rect 359 -865 360 -864
rect 436 -865 437 -864
rect 478 -865 479 -864
rect 485 -865 486 -864
rect 548 -865 549 -864
rect 562 -865 563 -864
rect 660 -865 661 -864
rect 121 -867 122 -866
rect 170 -867 171 -866
rect 173 -867 174 -866
rect 296 -867 297 -866
rect 306 -867 307 -866
rect 478 -867 479 -866
rect 513 -867 514 -866
rect 660 -867 661 -866
rect 142 -869 143 -868
rect 219 -869 220 -868
rect 275 -869 276 -868
rect 443 -869 444 -868
rect 450 -869 451 -868
rect 618 -869 619 -868
rect 156 -871 157 -870
rect 159 -871 160 -870
rect 163 -871 164 -870
rect 317 -871 318 -870
rect 345 -871 346 -870
rect 520 -871 521 -870
rect 156 -873 157 -872
rect 205 -873 206 -872
rect 345 -873 346 -872
rect 415 -873 416 -872
rect 443 -873 444 -872
rect 499 -873 500 -872
rect 513 -873 514 -872
rect 604 -873 605 -872
rect 117 -875 118 -874
rect 415 -875 416 -874
rect 453 -875 454 -874
rect 492 -875 493 -874
rect 597 -875 598 -874
rect 604 -875 605 -874
rect 635 -875 636 -874
rect 639 -875 640 -874
rect 163 -877 164 -876
rect 268 -877 269 -876
rect 453 -877 454 -876
rect 786 -877 787 -876
rect 170 -879 171 -878
rect 341 -879 342 -878
rect 457 -879 458 -878
rect 499 -879 500 -878
rect 135 -881 136 -880
rect 457 -881 458 -880
rect 492 -881 493 -880
rect 541 -881 542 -880
rect 135 -883 136 -882
rect 226 -883 227 -882
rect 268 -883 269 -882
rect 289 -883 290 -882
rect 541 -883 542 -882
rect 646 -883 647 -882
rect 79 -885 80 -884
rect 289 -885 290 -884
rect 583 -885 584 -884
rect 646 -885 647 -884
rect 177 -887 178 -886
rect 352 -887 353 -886
rect 583 -887 584 -886
rect 674 -887 675 -886
rect 177 -889 178 -888
rect 233 -889 234 -888
rect 674 -889 675 -888
rect 695 -889 696 -888
rect 180 -891 181 -890
rect 261 -891 262 -890
rect 233 -893 234 -892
rect 366 -893 367 -892
rect 366 -895 367 -894
rect 464 -895 465 -894
rect 464 -897 465 -896
rect 534 -897 535 -896
rect 534 -899 535 -898
rect 597 -899 598 -898
rect 2 -910 3 -909
rect 100 -910 101 -909
rect 103 -910 104 -909
rect 233 -910 234 -909
rect 240 -910 241 -909
rect 306 -910 307 -909
rect 338 -910 339 -909
rect 352 -910 353 -909
rect 359 -910 360 -909
rect 537 -910 538 -909
rect 548 -910 549 -909
rect 562 -910 563 -909
rect 576 -910 577 -909
rect 590 -910 591 -909
rect 607 -910 608 -909
rect 681 -910 682 -909
rect 695 -910 696 -909
rect 758 -910 759 -909
rect 23 -912 24 -911
rect 499 -912 500 -911
rect 509 -912 510 -911
rect 632 -912 633 -911
rect 737 -912 738 -911
rect 751 -912 752 -911
rect 26 -914 27 -913
rect 170 -914 171 -913
rect 205 -914 206 -913
rect 254 -914 255 -913
rect 257 -914 258 -913
rect 681 -914 682 -913
rect 30 -916 31 -915
rect 145 -916 146 -915
rect 205 -916 206 -915
rect 397 -916 398 -915
rect 404 -916 405 -915
rect 646 -916 647 -915
rect 30 -918 31 -917
rect 187 -918 188 -917
rect 212 -918 213 -917
rect 289 -918 290 -917
rect 296 -918 297 -917
rect 310 -918 311 -917
rect 383 -918 384 -917
rect 394 -918 395 -917
rect 408 -918 409 -917
rect 611 -918 612 -917
rect 618 -918 619 -917
rect 632 -918 633 -917
rect 37 -920 38 -919
rect 47 -920 48 -919
rect 54 -920 55 -919
rect 688 -920 689 -919
rect 40 -922 41 -921
rect 702 -922 703 -921
rect 65 -924 66 -923
rect 145 -924 146 -923
rect 156 -924 157 -923
rect 212 -924 213 -923
rect 229 -924 230 -923
rect 590 -924 591 -923
rect 597 -924 598 -923
rect 695 -924 696 -923
rect 65 -926 66 -925
rect 555 -926 556 -925
rect 576 -926 577 -925
rect 604 -926 605 -925
rect 621 -926 622 -925
rect 709 -926 710 -925
rect 72 -928 73 -927
rect 254 -928 255 -927
rect 275 -928 276 -927
rect 702 -928 703 -927
rect 72 -930 73 -929
rect 366 -930 367 -929
rect 387 -930 388 -929
rect 450 -930 451 -929
rect 478 -930 479 -929
rect 709 -930 710 -929
rect 79 -932 80 -931
rect 173 -932 174 -931
rect 219 -932 220 -931
rect 366 -932 367 -931
rect 394 -932 395 -931
rect 660 -932 661 -931
rect 688 -932 689 -931
rect 726 -932 727 -931
rect 61 -934 62 -933
rect 79 -934 80 -933
rect 86 -934 87 -933
rect 250 -934 251 -933
rect 275 -934 276 -933
rect 345 -934 346 -933
rect 362 -934 363 -933
rect 660 -934 661 -933
rect 93 -936 94 -935
rect 152 -936 153 -935
rect 156 -936 157 -935
rect 163 -936 164 -935
rect 226 -936 227 -935
rect 387 -936 388 -935
rect 415 -936 416 -935
rect 716 -936 717 -935
rect 93 -938 94 -937
rect 198 -938 199 -937
rect 233 -938 234 -937
rect 299 -938 300 -937
rect 303 -938 304 -937
rect 362 -938 363 -937
rect 450 -938 451 -937
rect 471 -938 472 -937
rect 478 -938 479 -937
rect 527 -938 528 -937
rect 534 -938 535 -937
rect 569 -938 570 -937
rect 625 -938 626 -937
rect 628 -938 629 -937
rect 44 -940 45 -939
rect 198 -940 199 -939
rect 240 -940 241 -939
rect 268 -940 269 -939
rect 278 -940 279 -939
rect 324 -940 325 -939
rect 499 -940 500 -939
rect 646 -940 647 -939
rect 44 -942 45 -941
rect 569 -942 570 -941
rect 625 -942 626 -941
rect 639 -942 640 -941
rect 107 -944 108 -943
rect 502 -944 503 -943
rect 513 -944 514 -943
rect 527 -944 528 -943
rect 555 -944 556 -943
rect 674 -944 675 -943
rect 107 -946 108 -945
rect 352 -946 353 -945
rect 513 -946 514 -945
rect 583 -946 584 -945
rect 628 -946 629 -945
rect 639 -946 640 -945
rect 114 -948 115 -947
rect 128 -948 129 -947
rect 135 -948 136 -947
rect 471 -948 472 -947
rect 520 -948 521 -947
rect 674 -948 675 -947
rect 16 -950 17 -949
rect 128 -950 129 -949
rect 163 -950 164 -949
rect 180 -950 181 -949
rect 261 -950 262 -949
rect 345 -950 346 -949
rect 520 -950 521 -949
rect 541 -950 542 -949
rect 562 -950 563 -949
rect 604 -950 605 -949
rect 16 -952 17 -951
rect 191 -952 192 -951
rect 261 -952 262 -951
rect 411 -952 412 -951
rect 100 -954 101 -953
rect 135 -954 136 -953
rect 149 -954 150 -953
rect 191 -954 192 -953
rect 282 -954 283 -953
rect 492 -954 493 -953
rect 117 -956 118 -955
rect 247 -956 248 -955
rect 285 -956 286 -955
rect 422 -956 423 -955
rect 485 -956 486 -955
rect 492 -956 493 -955
rect 121 -958 122 -957
rect 219 -958 220 -957
rect 310 -958 311 -957
rect 653 -958 654 -957
rect 58 -960 59 -959
rect 121 -960 122 -959
rect 142 -960 143 -959
rect 422 -960 423 -959
rect 653 -960 654 -959
rect 667 -960 668 -959
rect 9 -962 10 -961
rect 58 -962 59 -961
rect 149 -962 150 -961
rect 415 -962 416 -961
rect 180 -964 181 -963
rect 457 -964 458 -963
rect 324 -966 325 -965
rect 506 -966 507 -965
rect 313 -968 314 -967
rect 506 -968 507 -967
rect 331 -970 332 -969
rect 583 -970 584 -969
rect 51 -972 52 -971
rect 331 -972 332 -971
rect 373 -972 374 -971
rect 541 -972 542 -971
rect 184 -974 185 -973
rect 373 -974 374 -973
rect 401 -974 402 -973
rect 667 -974 668 -973
rect 184 -976 185 -975
rect 268 -976 269 -975
rect 401 -976 402 -975
rect 411 -976 412 -975
rect 457 -976 458 -975
rect 464 -976 465 -975
rect 429 -978 430 -977
rect 464 -978 465 -977
rect 429 -980 430 -979
rect 443 -980 444 -979
rect 380 -982 381 -981
rect 443 -982 444 -981
rect 9 -993 10 -992
rect 184 -993 185 -992
rect 187 -993 188 -992
rect 254 -993 255 -992
rect 275 -993 276 -992
rect 355 -993 356 -992
rect 404 -993 405 -992
rect 436 -993 437 -992
rect 443 -993 444 -992
rect 450 -993 451 -992
rect 464 -993 465 -992
rect 485 -993 486 -992
rect 499 -993 500 -992
rect 506 -993 507 -992
rect 520 -993 521 -992
rect 523 -993 524 -992
rect 527 -993 528 -992
rect 730 -993 731 -992
rect 751 -993 752 -992
rect 758 -993 759 -992
rect 26 -995 27 -994
rect 65 -995 66 -994
rect 79 -995 80 -994
rect 86 -995 87 -994
rect 89 -995 90 -994
rect 611 -995 612 -994
rect 618 -995 619 -994
rect 632 -995 633 -994
rect 716 -995 717 -994
rect 723 -995 724 -994
rect 30 -997 31 -996
rect 362 -997 363 -996
rect 425 -997 426 -996
rect 527 -997 528 -996
rect 604 -997 605 -996
rect 621 -997 622 -996
rect 625 -997 626 -996
rect 632 -997 633 -996
rect 709 -997 710 -996
rect 716 -997 717 -996
rect 37 -999 38 -998
rect 142 -999 143 -998
rect 149 -999 150 -998
rect 394 -999 395 -998
rect 436 -999 437 -998
rect 457 -999 458 -998
rect 464 -999 465 -998
rect 492 -999 493 -998
rect 502 -999 503 -998
rect 576 -999 577 -998
rect 695 -999 696 -998
rect 709 -999 710 -998
rect 37 -1001 38 -1000
rect 72 -1001 73 -1000
rect 79 -1001 80 -1000
rect 429 -1001 430 -1000
rect 457 -1001 458 -1000
rect 471 -1001 472 -1000
rect 478 -1001 479 -1000
rect 506 -1001 507 -1000
rect 520 -1001 521 -1000
rect 562 -1001 563 -1000
rect 695 -1001 696 -1000
rect 702 -1001 703 -1000
rect 44 -1003 45 -1002
rect 681 -1003 682 -1002
rect 688 -1003 689 -1002
rect 702 -1003 703 -1002
rect 47 -1005 48 -1004
rect 198 -1005 199 -1004
rect 205 -1005 206 -1004
rect 446 -1005 447 -1004
rect 485 -1005 486 -1004
rect 607 -1005 608 -1004
rect 674 -1005 675 -1004
rect 688 -1005 689 -1004
rect 54 -1007 55 -1006
rect 569 -1007 570 -1006
rect 660 -1007 661 -1006
rect 674 -1007 675 -1006
rect 58 -1009 59 -1008
rect 415 -1009 416 -1008
rect 488 -1009 489 -1008
rect 576 -1009 577 -1008
rect 660 -1009 661 -1008
rect 667 -1009 668 -1008
rect 68 -1011 69 -1010
rect 478 -1011 479 -1010
rect 523 -1011 524 -1010
rect 562 -1011 563 -1010
rect 569 -1011 570 -1010
rect 583 -1011 584 -1010
rect 86 -1013 87 -1012
rect 331 -1013 332 -1012
rect 352 -1013 353 -1012
rect 471 -1013 472 -1012
rect 555 -1013 556 -1012
rect 681 -1013 682 -1012
rect 93 -1015 94 -1014
rect 184 -1015 185 -1014
rect 191 -1015 192 -1014
rect 198 -1015 199 -1014
rect 205 -1015 206 -1014
rect 345 -1015 346 -1014
rect 366 -1015 367 -1014
rect 583 -1015 584 -1014
rect 2 -1017 3 -1016
rect 345 -1017 346 -1016
rect 366 -1017 367 -1016
rect 380 -1017 381 -1016
rect 383 -1017 384 -1016
rect 429 -1017 430 -1016
rect 534 -1017 535 -1016
rect 555 -1017 556 -1016
rect 93 -1019 94 -1018
rect 100 -1019 101 -1018
rect 107 -1019 108 -1018
rect 646 -1019 647 -1018
rect 16 -1021 17 -1020
rect 107 -1021 108 -1020
rect 114 -1021 115 -1020
rect 289 -1021 290 -1020
rect 292 -1021 293 -1020
rect 597 -1021 598 -1020
rect 16 -1023 17 -1022
rect 170 -1023 171 -1022
rect 180 -1023 181 -1022
rect 373 -1023 374 -1022
rect 394 -1023 395 -1022
rect 541 -1023 542 -1022
rect 100 -1025 101 -1024
rect 212 -1025 213 -1024
rect 219 -1025 220 -1024
rect 226 -1025 227 -1024
rect 240 -1025 241 -1024
rect 313 -1025 314 -1024
rect 317 -1025 318 -1024
rect 369 -1025 370 -1024
rect 373 -1025 374 -1024
rect 513 -1025 514 -1024
rect 534 -1025 535 -1024
rect 590 -1025 591 -1024
rect 23 -1027 24 -1026
rect 590 -1027 591 -1026
rect 75 -1029 76 -1028
rect 240 -1029 241 -1028
rect 247 -1029 248 -1028
rect 261 -1029 262 -1028
rect 268 -1029 269 -1028
rect 611 -1029 612 -1028
rect 117 -1031 118 -1030
rect 219 -1031 220 -1030
rect 226 -1031 227 -1030
rect 324 -1031 325 -1030
rect 331 -1031 332 -1030
rect 359 -1031 360 -1030
rect 142 -1033 143 -1032
rect 401 -1033 402 -1032
rect 156 -1035 157 -1034
rect 170 -1035 171 -1034
rect 177 -1035 178 -1034
rect 541 -1035 542 -1034
rect 128 -1037 129 -1036
rect 177 -1037 178 -1036
rect 212 -1037 213 -1036
rect 310 -1037 311 -1036
rect 317 -1037 318 -1036
rect 338 -1037 339 -1036
rect 401 -1037 402 -1036
rect 667 -1037 668 -1036
rect 103 -1039 104 -1038
rect 128 -1039 129 -1038
rect 135 -1039 136 -1038
rect 156 -1039 157 -1038
rect 163 -1039 164 -1038
rect 191 -1039 192 -1038
rect 250 -1039 251 -1038
rect 646 -1039 647 -1038
rect 121 -1041 122 -1040
rect 163 -1041 164 -1040
rect 254 -1041 255 -1040
rect 422 -1041 423 -1040
rect 30 -1043 31 -1042
rect 121 -1043 122 -1042
rect 135 -1043 136 -1042
rect 149 -1043 150 -1042
rect 261 -1043 262 -1042
rect 296 -1043 297 -1042
rect 306 -1043 307 -1042
rect 338 -1043 339 -1042
rect 422 -1043 423 -1042
rect 513 -1043 514 -1042
rect 233 -1045 234 -1044
rect 296 -1045 297 -1044
rect 310 -1045 311 -1044
rect 625 -1045 626 -1044
rect 233 -1047 234 -1046
rect 450 -1047 451 -1046
rect 268 -1049 269 -1048
rect 408 -1049 409 -1048
rect 275 -1051 276 -1050
rect 303 -1051 304 -1050
rect 320 -1051 321 -1050
rect 387 -1051 388 -1050
rect 282 -1053 283 -1052
rect 411 -1053 412 -1052
rect 303 -1055 304 -1054
rect 492 -1055 493 -1054
rect 324 -1057 325 -1056
rect 352 -1057 353 -1056
rect 387 -1057 388 -1056
rect 397 -1057 398 -1056
rect 16 -1068 17 -1067
rect 359 -1068 360 -1067
rect 362 -1068 363 -1067
rect 695 -1068 696 -1067
rect 730 -1068 731 -1067
rect 737 -1068 738 -1067
rect 751 -1068 752 -1067
rect 754 -1068 755 -1067
rect 16 -1070 17 -1069
rect 261 -1070 262 -1069
rect 268 -1070 269 -1069
rect 289 -1070 290 -1069
rect 306 -1070 307 -1069
rect 681 -1070 682 -1069
rect 754 -1070 755 -1069
rect 793 -1070 794 -1069
rect 26 -1072 27 -1071
rect 86 -1072 87 -1071
rect 89 -1072 90 -1071
rect 173 -1072 174 -1071
rect 177 -1072 178 -1071
rect 261 -1072 262 -1071
rect 310 -1072 311 -1071
rect 345 -1072 346 -1071
rect 369 -1072 370 -1071
rect 548 -1072 549 -1071
rect 597 -1072 598 -1071
rect 730 -1072 731 -1071
rect 9 -1074 10 -1073
rect 86 -1074 87 -1073
rect 107 -1074 108 -1073
rect 303 -1074 304 -1073
rect 310 -1074 311 -1073
rect 324 -1074 325 -1073
rect 327 -1074 328 -1073
rect 373 -1074 374 -1073
rect 383 -1074 384 -1073
rect 506 -1074 507 -1073
rect 509 -1074 510 -1073
rect 681 -1074 682 -1073
rect 9 -1076 10 -1075
rect 121 -1076 122 -1075
rect 156 -1076 157 -1075
rect 187 -1076 188 -1075
rect 205 -1076 206 -1075
rect 376 -1076 377 -1075
rect 394 -1076 395 -1075
rect 439 -1076 440 -1075
rect 464 -1076 465 -1075
rect 786 -1076 787 -1075
rect 30 -1078 31 -1077
rect 471 -1078 472 -1077
rect 474 -1078 475 -1077
rect 576 -1078 577 -1077
rect 604 -1078 605 -1077
rect 653 -1078 654 -1077
rect 660 -1078 661 -1077
rect 695 -1078 696 -1077
rect 37 -1080 38 -1079
rect 138 -1080 139 -1079
rect 156 -1080 157 -1079
rect 166 -1080 167 -1079
rect 170 -1080 171 -1079
rect 271 -1080 272 -1079
rect 331 -1080 332 -1079
rect 597 -1080 598 -1079
rect 632 -1080 633 -1079
rect 653 -1080 654 -1079
rect 667 -1080 668 -1079
rect 779 -1080 780 -1079
rect 44 -1082 45 -1081
rect 219 -1082 220 -1081
rect 247 -1082 248 -1081
rect 415 -1082 416 -1081
rect 418 -1082 419 -1081
rect 723 -1082 724 -1081
rect 47 -1084 48 -1083
rect 65 -1084 66 -1083
rect 72 -1084 73 -1083
rect 135 -1084 136 -1083
rect 138 -1084 139 -1083
rect 583 -1084 584 -1083
rect 625 -1084 626 -1083
rect 667 -1084 668 -1083
rect 709 -1084 710 -1083
rect 723 -1084 724 -1083
rect 23 -1086 24 -1085
rect 65 -1086 66 -1085
rect 100 -1086 101 -1085
rect 187 -1086 188 -1085
rect 198 -1086 199 -1085
rect 219 -1086 220 -1085
rect 250 -1086 251 -1085
rect 275 -1086 276 -1085
rect 345 -1086 346 -1085
rect 425 -1086 426 -1085
rect 450 -1086 451 -1085
rect 625 -1086 626 -1085
rect 632 -1086 633 -1085
rect 674 -1086 675 -1085
rect 688 -1086 689 -1085
rect 709 -1086 710 -1085
rect 58 -1088 59 -1087
rect 107 -1088 108 -1087
rect 114 -1088 115 -1087
rect 191 -1088 192 -1087
rect 208 -1088 209 -1087
rect 254 -1088 255 -1087
rect 275 -1088 276 -1087
rect 338 -1088 339 -1087
rect 380 -1088 381 -1087
rect 604 -1088 605 -1087
rect 639 -1088 640 -1087
rect 660 -1088 661 -1087
rect 58 -1090 59 -1089
rect 142 -1090 143 -1089
rect 163 -1090 164 -1089
rect 331 -1090 332 -1089
rect 380 -1090 381 -1089
rect 740 -1090 741 -1089
rect 114 -1092 115 -1091
rect 212 -1092 213 -1091
rect 387 -1092 388 -1091
rect 415 -1092 416 -1091
rect 425 -1092 426 -1091
rect 716 -1092 717 -1091
rect 79 -1094 80 -1093
rect 387 -1094 388 -1093
rect 397 -1094 398 -1093
rect 583 -1094 584 -1093
rect 611 -1094 612 -1093
rect 639 -1094 640 -1093
rect 646 -1094 647 -1093
rect 674 -1094 675 -1093
rect 117 -1096 118 -1095
rect 296 -1096 297 -1095
rect 401 -1096 402 -1095
rect 408 -1096 409 -1095
rect 436 -1096 437 -1095
rect 450 -1096 451 -1095
rect 457 -1096 458 -1095
rect 464 -1096 465 -1095
rect 471 -1096 472 -1095
rect 716 -1096 717 -1095
rect 51 -1098 52 -1097
rect 457 -1098 458 -1097
rect 499 -1098 500 -1097
rect 814 -1098 815 -1097
rect 51 -1100 52 -1099
rect 205 -1100 206 -1099
rect 212 -1100 213 -1099
rect 317 -1100 318 -1099
rect 436 -1100 437 -1099
rect 562 -1100 563 -1099
rect 618 -1100 619 -1099
rect 646 -1100 647 -1099
rect 37 -1102 38 -1101
rect 317 -1102 318 -1101
rect 513 -1102 514 -1101
rect 548 -1102 549 -1101
rect 562 -1102 563 -1101
rect 569 -1102 570 -1101
rect 103 -1104 104 -1103
rect 499 -1104 500 -1103
rect 534 -1104 535 -1103
rect 576 -1104 577 -1103
rect 121 -1106 122 -1105
rect 422 -1106 423 -1105
rect 527 -1106 528 -1105
rect 534 -1106 535 -1105
rect 128 -1108 129 -1107
rect 142 -1108 143 -1107
rect 163 -1108 164 -1107
rect 478 -1108 479 -1107
rect 527 -1108 528 -1107
rect 555 -1108 556 -1107
rect 128 -1110 129 -1109
rect 149 -1110 150 -1109
rect 177 -1110 178 -1109
rect 282 -1110 283 -1109
rect 289 -1110 290 -1109
rect 569 -1110 570 -1109
rect 79 -1112 80 -1111
rect 149 -1112 150 -1111
rect 180 -1112 181 -1111
rect 324 -1112 325 -1111
rect 429 -1112 430 -1111
rect 478 -1112 479 -1111
rect 555 -1112 556 -1111
rect 590 -1112 591 -1111
rect 184 -1114 185 -1113
rect 198 -1114 199 -1113
rect 240 -1114 241 -1113
rect 296 -1114 297 -1113
rect 366 -1114 367 -1113
rect 590 -1114 591 -1113
rect 184 -1116 185 -1115
rect 233 -1116 234 -1115
rect 240 -1116 241 -1115
rect 247 -1116 248 -1115
rect 282 -1116 283 -1115
rect 338 -1116 339 -1115
rect 366 -1116 367 -1115
rect 513 -1116 514 -1115
rect 191 -1118 192 -1117
rect 303 -1118 304 -1117
rect 429 -1118 430 -1117
rect 443 -1118 444 -1117
rect 194 -1120 195 -1119
rect 254 -1120 255 -1119
rect 443 -1120 444 -1119
rect 492 -1120 493 -1119
rect 233 -1122 234 -1121
rect 408 -1122 409 -1121
rect 485 -1122 486 -1121
rect 492 -1122 493 -1121
rect 320 -1124 321 -1123
rect 485 -1124 486 -1123
rect 9 -1135 10 -1134
rect 327 -1135 328 -1134
rect 348 -1135 349 -1134
rect 506 -1135 507 -1134
rect 509 -1135 510 -1134
rect 702 -1135 703 -1134
rect 716 -1135 717 -1134
rect 772 -1135 773 -1134
rect 793 -1135 794 -1134
rect 800 -1135 801 -1134
rect 9 -1137 10 -1136
rect 282 -1137 283 -1136
rect 310 -1137 311 -1136
rect 320 -1137 321 -1136
rect 355 -1137 356 -1136
rect 373 -1137 374 -1136
rect 422 -1137 423 -1136
rect 593 -1137 594 -1136
rect 646 -1137 647 -1136
rect 688 -1137 689 -1136
rect 740 -1137 741 -1136
rect 793 -1137 794 -1136
rect 23 -1139 24 -1138
rect 338 -1139 339 -1138
rect 366 -1139 367 -1138
rect 548 -1139 549 -1138
rect 555 -1139 556 -1138
rect 765 -1139 766 -1138
rect 26 -1141 27 -1140
rect 639 -1141 640 -1140
rect 744 -1141 745 -1140
rect 779 -1141 780 -1140
rect 30 -1143 31 -1142
rect 597 -1143 598 -1142
rect 723 -1143 724 -1142
rect 779 -1143 780 -1142
rect 37 -1145 38 -1144
rect 187 -1145 188 -1144
rect 194 -1145 195 -1144
rect 331 -1145 332 -1144
rect 341 -1145 342 -1144
rect 597 -1145 598 -1144
rect 674 -1145 675 -1144
rect 723 -1145 724 -1144
rect 751 -1145 752 -1144
rect 758 -1145 759 -1144
rect 44 -1147 45 -1146
rect 338 -1147 339 -1146
rect 373 -1147 374 -1146
rect 513 -1147 514 -1146
rect 520 -1147 521 -1146
rect 702 -1147 703 -1146
rect 44 -1149 45 -1148
rect 429 -1149 430 -1148
rect 432 -1149 433 -1148
rect 716 -1149 717 -1148
rect 54 -1151 55 -1150
rect 457 -1151 458 -1150
rect 467 -1151 468 -1150
rect 492 -1151 493 -1150
rect 534 -1151 535 -1150
rect 611 -1151 612 -1150
rect 632 -1151 633 -1150
rect 751 -1151 752 -1150
rect 72 -1153 73 -1152
rect 247 -1153 248 -1152
rect 254 -1153 255 -1152
rect 310 -1153 311 -1152
rect 324 -1153 325 -1152
rect 366 -1153 367 -1152
rect 394 -1153 395 -1152
rect 674 -1153 675 -1152
rect 695 -1153 696 -1152
rect 758 -1153 759 -1152
rect 79 -1155 80 -1154
rect 324 -1155 325 -1154
rect 331 -1155 332 -1154
rect 380 -1155 381 -1154
rect 397 -1155 398 -1154
rect 555 -1155 556 -1154
rect 562 -1155 563 -1154
rect 632 -1155 633 -1154
rect 79 -1157 80 -1156
rect 142 -1157 143 -1156
rect 145 -1157 146 -1156
rect 208 -1157 209 -1156
rect 212 -1157 213 -1156
rect 236 -1157 237 -1156
rect 247 -1157 248 -1156
rect 257 -1157 258 -1156
rect 275 -1157 276 -1156
rect 436 -1157 437 -1156
rect 443 -1157 444 -1156
rect 562 -1157 563 -1156
rect 569 -1157 570 -1156
rect 747 -1157 748 -1156
rect 16 -1159 17 -1158
rect 275 -1159 276 -1158
rect 292 -1159 293 -1158
rect 380 -1159 381 -1158
rect 401 -1159 402 -1158
rect 492 -1159 493 -1158
rect 541 -1159 542 -1158
rect 618 -1159 619 -1158
rect 16 -1161 17 -1160
rect 163 -1161 164 -1160
rect 166 -1161 167 -1160
rect 180 -1161 181 -1160
rect 187 -1161 188 -1160
rect 457 -1161 458 -1160
rect 474 -1161 475 -1160
rect 527 -1161 528 -1160
rect 548 -1161 549 -1160
rect 786 -1161 787 -1160
rect 100 -1163 101 -1162
rect 513 -1163 514 -1162
rect 569 -1163 570 -1162
rect 814 -1163 815 -1162
rect 93 -1165 94 -1164
rect 100 -1165 101 -1164
rect 114 -1165 115 -1164
rect 681 -1165 682 -1164
rect 730 -1165 731 -1164
rect 786 -1165 787 -1164
rect 93 -1167 94 -1166
rect 390 -1167 391 -1166
rect 408 -1167 409 -1166
rect 534 -1167 535 -1166
rect 576 -1167 577 -1166
rect 639 -1167 640 -1166
rect 653 -1167 654 -1166
rect 730 -1167 731 -1166
rect 117 -1169 118 -1168
rect 282 -1169 283 -1168
rect 352 -1169 353 -1168
rect 695 -1169 696 -1168
rect 117 -1171 118 -1170
rect 191 -1171 192 -1170
rect 198 -1171 199 -1170
rect 289 -1171 290 -1170
rect 296 -1171 297 -1170
rect 352 -1171 353 -1170
rect 359 -1171 360 -1170
rect 443 -1171 444 -1170
rect 450 -1171 451 -1170
rect 520 -1171 521 -1170
rect 590 -1171 591 -1170
rect 646 -1171 647 -1170
rect 121 -1173 122 -1172
rect 149 -1173 150 -1172
rect 152 -1173 153 -1172
rect 583 -1173 584 -1172
rect 625 -1173 626 -1172
rect 681 -1173 682 -1172
rect 121 -1175 122 -1174
rect 128 -1175 129 -1174
rect 135 -1175 136 -1174
rect 583 -1175 584 -1174
rect 625 -1175 626 -1174
rect 660 -1175 661 -1174
rect 51 -1177 52 -1176
rect 128 -1177 129 -1176
rect 138 -1177 139 -1176
rect 317 -1177 318 -1176
rect 429 -1177 430 -1176
rect 471 -1177 472 -1176
rect 485 -1177 486 -1176
rect 653 -1177 654 -1176
rect 33 -1179 34 -1178
rect 485 -1179 486 -1178
rect 499 -1179 500 -1178
rect 576 -1179 577 -1178
rect 51 -1181 52 -1180
rect 737 -1181 738 -1180
rect 58 -1183 59 -1182
rect 135 -1183 136 -1182
rect 177 -1183 178 -1182
rect 369 -1183 370 -1182
rect 415 -1183 416 -1182
rect 499 -1183 500 -1182
rect 58 -1185 59 -1184
rect 68 -1185 69 -1184
rect 198 -1185 199 -1184
rect 261 -1185 262 -1184
rect 296 -1185 297 -1184
rect 425 -1185 426 -1184
rect 450 -1185 451 -1184
rect 478 -1185 479 -1184
rect 65 -1187 66 -1186
rect 415 -1187 416 -1186
rect 464 -1187 465 -1186
rect 527 -1187 528 -1186
rect 65 -1189 66 -1188
rect 72 -1189 73 -1188
rect 205 -1189 206 -1188
rect 394 -1189 395 -1188
rect 471 -1189 472 -1188
rect 604 -1189 605 -1188
rect 212 -1191 213 -1190
rect 240 -1191 241 -1190
rect 250 -1191 251 -1190
rect 604 -1191 605 -1190
rect 226 -1193 227 -1192
rect 233 -1193 234 -1192
rect 240 -1193 241 -1192
rect 404 -1193 405 -1192
rect 219 -1195 220 -1194
rect 226 -1195 227 -1194
rect 261 -1195 262 -1194
rect 268 -1195 269 -1194
rect 303 -1195 304 -1194
rect 359 -1195 360 -1194
rect 369 -1195 370 -1194
rect 387 -1195 388 -1194
rect 40 -1197 41 -1196
rect 219 -1197 220 -1196
rect 268 -1197 269 -1196
rect 411 -1197 412 -1196
rect 303 -1199 304 -1198
rect 345 -1199 346 -1198
rect 345 -1201 346 -1200
rect 667 -1201 668 -1200
rect 667 -1203 668 -1202
rect 709 -1203 710 -1202
rect 478 -1205 479 -1204
rect 709 -1205 710 -1204
rect 2 -1216 3 -1215
rect 135 -1216 136 -1215
rect 184 -1216 185 -1215
rect 198 -1216 199 -1215
rect 254 -1216 255 -1215
rect 310 -1216 311 -1215
rect 317 -1216 318 -1215
rect 443 -1216 444 -1215
rect 471 -1216 472 -1215
rect 506 -1216 507 -1215
rect 541 -1216 542 -1215
rect 646 -1216 647 -1215
rect 649 -1216 650 -1215
rect 786 -1216 787 -1215
rect 789 -1216 790 -1215
rect 800 -1216 801 -1215
rect 9 -1218 10 -1217
rect 348 -1218 349 -1217
rect 362 -1218 363 -1217
rect 597 -1218 598 -1217
rect 660 -1218 661 -1217
rect 786 -1218 787 -1217
rect 9 -1220 10 -1219
rect 30 -1220 31 -1219
rect 33 -1220 34 -1219
rect 663 -1220 664 -1219
rect 667 -1220 668 -1219
rect 737 -1220 738 -1219
rect 16 -1222 17 -1221
rect 89 -1222 90 -1221
rect 128 -1222 129 -1221
rect 394 -1222 395 -1221
rect 397 -1222 398 -1221
rect 520 -1222 521 -1221
rect 593 -1222 594 -1221
rect 730 -1222 731 -1221
rect 16 -1224 17 -1223
rect 145 -1224 146 -1223
rect 198 -1224 199 -1223
rect 380 -1224 381 -1223
rect 387 -1224 388 -1223
rect 534 -1224 535 -1223
rect 681 -1224 682 -1223
rect 730 -1224 731 -1223
rect 30 -1226 31 -1225
rect 187 -1226 188 -1225
rect 254 -1226 255 -1225
rect 327 -1226 328 -1225
rect 345 -1226 346 -1225
rect 485 -1226 486 -1225
rect 506 -1226 507 -1225
rect 611 -1226 612 -1225
rect 37 -1228 38 -1227
rect 268 -1228 269 -1227
rect 278 -1228 279 -1227
rect 590 -1228 591 -1227
rect 23 -1230 24 -1229
rect 268 -1230 269 -1229
rect 282 -1230 283 -1229
rect 345 -1230 346 -1229
rect 366 -1230 367 -1229
rect 499 -1230 500 -1229
rect 520 -1230 521 -1229
rect 576 -1230 577 -1229
rect 23 -1232 24 -1231
rect 219 -1232 220 -1231
rect 247 -1232 248 -1231
rect 499 -1232 500 -1231
rect 555 -1232 556 -1231
rect 681 -1232 682 -1231
rect 51 -1234 52 -1233
rect 58 -1234 59 -1233
rect 68 -1234 69 -1233
rect 72 -1234 73 -1233
rect 75 -1234 76 -1233
rect 436 -1234 437 -1233
rect 443 -1234 444 -1233
rect 492 -1234 493 -1233
rect 555 -1234 556 -1233
rect 653 -1234 654 -1233
rect 51 -1236 52 -1235
rect 121 -1236 122 -1235
rect 128 -1236 129 -1235
rect 338 -1236 339 -1235
rect 373 -1236 374 -1235
rect 541 -1236 542 -1235
rect 576 -1236 577 -1235
rect 604 -1236 605 -1235
rect 653 -1236 654 -1235
rect 688 -1236 689 -1235
rect 54 -1238 55 -1237
rect 492 -1238 493 -1237
rect 688 -1238 689 -1237
rect 758 -1238 759 -1237
rect 58 -1240 59 -1239
rect 240 -1240 241 -1239
rect 247 -1240 248 -1239
rect 289 -1240 290 -1239
rect 317 -1240 318 -1239
rect 422 -1240 423 -1239
rect 464 -1240 465 -1239
rect 597 -1240 598 -1239
rect 758 -1240 759 -1239
rect 779 -1240 780 -1239
rect 79 -1242 80 -1241
rect 142 -1242 143 -1241
rect 145 -1242 146 -1241
rect 191 -1242 192 -1241
rect 212 -1242 213 -1241
rect 219 -1242 220 -1241
rect 240 -1242 241 -1241
rect 352 -1242 353 -1241
rect 373 -1242 374 -1241
rect 429 -1242 430 -1241
rect 464 -1242 465 -1241
rect 513 -1242 514 -1241
rect 79 -1244 80 -1243
rect 331 -1244 332 -1243
rect 334 -1244 335 -1243
rect 604 -1244 605 -1243
rect 86 -1246 87 -1245
rect 359 -1246 360 -1245
rect 390 -1246 391 -1245
rect 632 -1246 633 -1245
rect 93 -1248 94 -1247
rect 121 -1248 122 -1247
rect 135 -1248 136 -1247
rect 205 -1248 206 -1247
rect 212 -1248 213 -1247
rect 415 -1248 416 -1247
rect 422 -1248 423 -1247
rect 450 -1248 451 -1247
rect 478 -1248 479 -1247
rect 751 -1248 752 -1247
rect 93 -1250 94 -1249
rect 177 -1250 178 -1249
rect 184 -1250 185 -1249
rect 436 -1250 437 -1249
rect 450 -1250 451 -1249
rect 667 -1250 668 -1249
rect 44 -1252 45 -1251
rect 177 -1252 178 -1251
rect 191 -1252 192 -1251
rect 303 -1252 304 -1251
rect 324 -1252 325 -1251
rect 723 -1252 724 -1251
rect 44 -1254 45 -1253
rect 72 -1254 73 -1253
rect 107 -1254 108 -1253
rect 289 -1254 290 -1253
rect 324 -1254 325 -1253
rect 457 -1254 458 -1253
rect 478 -1254 479 -1253
rect 527 -1254 528 -1253
rect 632 -1254 633 -1253
rect 779 -1254 780 -1253
rect 107 -1256 108 -1255
rect 170 -1256 171 -1255
rect 205 -1256 206 -1255
rect 226 -1256 227 -1255
rect 282 -1256 283 -1255
rect 341 -1256 342 -1255
rect 401 -1256 402 -1255
rect 548 -1256 549 -1255
rect 723 -1256 724 -1255
rect 744 -1256 745 -1255
rect 65 -1258 66 -1257
rect 170 -1258 171 -1257
rect 341 -1258 342 -1257
rect 562 -1258 563 -1257
rect 744 -1258 745 -1257
rect 772 -1258 773 -1257
rect 114 -1260 115 -1259
rect 751 -1260 752 -1259
rect 772 -1260 773 -1259
rect 793 -1260 794 -1259
rect 166 -1262 167 -1261
rect 380 -1262 381 -1261
rect 401 -1262 402 -1261
rect 765 -1262 766 -1261
rect 310 -1264 311 -1263
rect 562 -1264 563 -1263
rect 404 -1266 405 -1265
rect 611 -1266 612 -1265
rect 404 -1268 405 -1267
rect 534 -1268 535 -1267
rect 548 -1268 549 -1267
rect 618 -1268 619 -1267
rect 411 -1270 412 -1269
rect 639 -1270 640 -1269
rect 411 -1272 412 -1271
rect 702 -1272 703 -1271
rect 429 -1274 430 -1273
rect 583 -1274 584 -1273
rect 639 -1274 640 -1273
rect 695 -1274 696 -1273
rect 702 -1274 703 -1273
rect 716 -1274 717 -1273
rect 457 -1276 458 -1275
rect 485 -1276 486 -1275
rect 513 -1276 514 -1275
rect 572 -1276 573 -1275
rect 646 -1276 647 -1275
rect 716 -1276 717 -1275
rect 474 -1278 475 -1277
rect 583 -1278 584 -1277
rect 695 -1278 696 -1277
rect 709 -1278 710 -1277
rect 303 -1280 304 -1279
rect 709 -1280 710 -1279
rect 481 -1282 482 -1281
rect 782 -1282 783 -1281
rect 527 -1284 528 -1283
rect 674 -1284 675 -1283
rect 569 -1286 570 -1285
rect 618 -1286 619 -1285
rect 625 -1286 626 -1285
rect 674 -1286 675 -1285
rect 275 -1288 276 -1287
rect 625 -1288 626 -1287
rect 233 -1290 234 -1289
rect 275 -1290 276 -1289
rect 233 -1292 234 -1291
rect 261 -1292 262 -1291
rect 261 -1294 262 -1293
rect 296 -1294 297 -1293
rect 296 -1296 297 -1295
rect 408 -1296 409 -1295
rect 408 -1298 409 -1297
rect 415 -1298 416 -1297
rect 2 -1309 3 -1308
rect 348 -1309 349 -1308
rect 355 -1309 356 -1308
rect 751 -1309 752 -1308
rect 782 -1309 783 -1308
rect 800 -1309 801 -1308
rect 9 -1311 10 -1310
rect 180 -1311 181 -1310
rect 191 -1311 192 -1310
rect 313 -1311 314 -1310
rect 359 -1311 360 -1310
rect 499 -1311 500 -1310
rect 516 -1311 517 -1310
rect 674 -1311 675 -1310
rect 709 -1311 710 -1310
rect 768 -1311 769 -1310
rect 9 -1313 10 -1312
rect 320 -1313 321 -1312
rect 362 -1313 363 -1312
rect 562 -1313 563 -1312
rect 565 -1313 566 -1312
rect 705 -1313 706 -1312
rect 730 -1313 731 -1312
rect 779 -1313 780 -1312
rect 30 -1315 31 -1314
rect 33 -1315 34 -1314
rect 40 -1315 41 -1314
rect 44 -1315 45 -1314
rect 65 -1315 66 -1314
rect 527 -1315 528 -1314
rect 537 -1315 538 -1314
rect 737 -1315 738 -1314
rect 30 -1317 31 -1316
rect 128 -1317 129 -1316
rect 149 -1317 150 -1316
rect 187 -1317 188 -1316
rect 198 -1317 199 -1316
rect 352 -1317 353 -1316
rect 404 -1317 405 -1316
rect 492 -1317 493 -1316
rect 527 -1317 528 -1316
rect 555 -1317 556 -1316
rect 562 -1317 563 -1316
rect 695 -1317 696 -1316
rect 44 -1319 45 -1318
rect 464 -1319 465 -1318
rect 492 -1319 493 -1318
rect 583 -1319 584 -1318
rect 590 -1319 591 -1318
rect 709 -1319 710 -1318
rect 51 -1321 52 -1320
rect 187 -1321 188 -1320
rect 198 -1321 199 -1320
rect 205 -1321 206 -1320
rect 215 -1321 216 -1320
rect 359 -1321 360 -1320
rect 408 -1321 409 -1320
rect 702 -1321 703 -1320
rect 51 -1323 52 -1322
rect 145 -1323 146 -1322
rect 149 -1323 150 -1322
rect 156 -1323 157 -1322
rect 163 -1323 164 -1322
rect 289 -1323 290 -1322
rect 296 -1323 297 -1322
rect 366 -1323 367 -1322
rect 457 -1323 458 -1322
rect 520 -1323 521 -1322
rect 534 -1323 535 -1322
rect 590 -1323 591 -1322
rect 639 -1323 640 -1322
rect 691 -1323 692 -1322
rect 702 -1323 703 -1322
rect 723 -1323 724 -1322
rect 68 -1325 69 -1324
rect 93 -1325 94 -1324
rect 114 -1325 115 -1324
rect 201 -1325 202 -1324
rect 219 -1325 220 -1324
rect 229 -1325 230 -1324
rect 268 -1325 269 -1324
rect 289 -1325 290 -1324
rect 310 -1325 311 -1324
rect 394 -1325 395 -1324
rect 429 -1325 430 -1324
rect 534 -1325 535 -1324
rect 541 -1325 542 -1324
rect 555 -1325 556 -1324
rect 572 -1325 573 -1324
rect 758 -1325 759 -1324
rect 58 -1327 59 -1326
rect 219 -1327 220 -1326
rect 226 -1327 227 -1326
rect 247 -1327 248 -1326
rect 275 -1327 276 -1326
rect 408 -1327 409 -1326
rect 457 -1327 458 -1326
rect 478 -1327 479 -1326
rect 485 -1327 486 -1326
rect 520 -1327 521 -1326
rect 541 -1327 542 -1326
rect 548 -1327 549 -1326
rect 576 -1327 577 -1326
rect 583 -1327 584 -1326
rect 639 -1327 640 -1326
rect 653 -1327 654 -1326
rect 688 -1327 689 -1326
rect 695 -1327 696 -1326
rect 744 -1327 745 -1326
rect 758 -1327 759 -1326
rect 23 -1329 24 -1328
rect 275 -1329 276 -1328
rect 296 -1329 297 -1328
rect 576 -1329 577 -1328
rect 653 -1329 654 -1328
rect 667 -1329 668 -1328
rect 23 -1331 24 -1330
rect 415 -1331 416 -1330
rect 425 -1331 426 -1330
rect 667 -1331 668 -1330
rect 65 -1333 66 -1332
rect 93 -1333 94 -1332
rect 114 -1333 115 -1332
rect 282 -1333 283 -1332
rect 345 -1333 346 -1332
rect 415 -1333 416 -1332
rect 471 -1333 472 -1332
rect 485 -1333 486 -1332
rect 506 -1333 507 -1332
rect 548 -1333 549 -1332
rect 72 -1335 73 -1334
rect 646 -1335 647 -1334
rect 75 -1337 76 -1336
rect 429 -1337 430 -1336
rect 506 -1337 507 -1336
rect 513 -1337 514 -1336
rect 82 -1339 83 -1338
rect 107 -1339 108 -1338
rect 117 -1339 118 -1338
rect 499 -1339 500 -1338
rect 107 -1341 108 -1340
rect 184 -1341 185 -1340
rect 191 -1341 192 -1340
rect 688 -1341 689 -1340
rect 117 -1343 118 -1342
rect 142 -1343 143 -1342
rect 156 -1343 157 -1342
rect 170 -1343 171 -1342
rect 177 -1343 178 -1342
rect 247 -1343 248 -1342
rect 268 -1343 269 -1342
rect 478 -1343 479 -1342
rect 16 -1345 17 -1344
rect 170 -1345 171 -1344
rect 184 -1345 185 -1344
rect 338 -1345 339 -1344
rect 352 -1345 353 -1344
rect 373 -1345 374 -1344
rect 380 -1345 381 -1344
rect 394 -1345 395 -1344
rect 464 -1345 465 -1344
rect 513 -1345 514 -1344
rect 37 -1347 38 -1346
rect 142 -1347 143 -1346
rect 163 -1347 164 -1346
rect 436 -1347 437 -1346
rect 58 -1349 59 -1348
rect 177 -1349 178 -1348
rect 233 -1349 234 -1348
rect 282 -1349 283 -1348
rect 366 -1349 367 -1348
rect 446 -1349 447 -1348
rect 86 -1351 87 -1350
rect 233 -1351 234 -1350
rect 373 -1351 374 -1350
rect 450 -1351 451 -1350
rect 121 -1353 122 -1352
rect 128 -1353 129 -1352
rect 135 -1353 136 -1352
rect 205 -1353 206 -1352
rect 380 -1353 381 -1352
rect 597 -1353 598 -1352
rect 121 -1355 122 -1354
rect 254 -1355 255 -1354
rect 387 -1355 388 -1354
rect 471 -1355 472 -1354
rect 597 -1355 598 -1354
rect 611 -1355 612 -1354
rect 135 -1357 136 -1356
rect 334 -1357 335 -1356
rect 387 -1357 388 -1356
rect 401 -1357 402 -1356
rect 422 -1357 423 -1356
rect 436 -1357 437 -1356
rect 443 -1357 444 -1356
rect 450 -1357 451 -1356
rect 611 -1357 612 -1356
rect 625 -1357 626 -1356
rect 166 -1359 167 -1358
rect 481 -1359 482 -1358
rect 254 -1361 255 -1360
rect 317 -1361 318 -1360
rect 401 -1361 402 -1360
rect 674 -1361 675 -1360
rect 212 -1363 213 -1362
rect 317 -1363 318 -1362
rect 443 -1363 444 -1362
rect 618 -1363 619 -1362
rect 33 -1365 34 -1364
rect 212 -1365 213 -1364
rect 261 -1365 262 -1364
rect 334 -1365 335 -1364
rect 618 -1365 619 -1364
rect 660 -1365 661 -1364
rect 79 -1367 80 -1366
rect 261 -1367 262 -1366
rect 303 -1367 304 -1366
rect 422 -1367 423 -1366
rect 660 -1367 661 -1366
rect 681 -1367 682 -1366
rect 79 -1369 80 -1368
rect 604 -1369 605 -1368
rect 681 -1369 682 -1368
rect 716 -1369 717 -1368
rect 303 -1371 304 -1370
rect 324 -1371 325 -1370
rect 331 -1371 332 -1370
rect 604 -1371 605 -1370
rect 240 -1373 241 -1372
rect 324 -1373 325 -1372
rect 240 -1375 241 -1374
rect 411 -1375 412 -1374
rect 9 -1386 10 -1385
rect 142 -1386 143 -1385
rect 149 -1386 150 -1385
rect 163 -1386 164 -1385
rect 170 -1386 171 -1385
rect 212 -1386 213 -1385
rect 271 -1386 272 -1385
rect 324 -1386 325 -1385
rect 338 -1386 339 -1385
rect 345 -1386 346 -1385
rect 383 -1386 384 -1385
rect 744 -1386 745 -1385
rect 758 -1386 759 -1385
rect 782 -1386 783 -1385
rect 786 -1386 787 -1385
rect 828 -1386 829 -1385
rect 16 -1388 17 -1387
rect 180 -1388 181 -1387
rect 275 -1388 276 -1387
rect 380 -1388 381 -1387
rect 411 -1388 412 -1387
rect 737 -1388 738 -1387
rect 779 -1388 780 -1387
rect 807 -1388 808 -1387
rect 37 -1390 38 -1389
rect 135 -1390 136 -1389
rect 149 -1390 150 -1389
rect 278 -1390 279 -1389
rect 296 -1390 297 -1389
rect 429 -1390 430 -1389
rect 443 -1390 444 -1389
rect 653 -1390 654 -1389
rect 674 -1390 675 -1389
rect 730 -1390 731 -1389
rect 789 -1390 790 -1389
rect 800 -1390 801 -1389
rect 44 -1392 45 -1391
rect 215 -1392 216 -1391
rect 247 -1392 248 -1391
rect 296 -1392 297 -1391
rect 310 -1392 311 -1391
rect 331 -1392 332 -1391
rect 338 -1392 339 -1391
rect 408 -1392 409 -1391
rect 443 -1392 444 -1391
rect 509 -1392 510 -1391
rect 534 -1392 535 -1391
rect 688 -1392 689 -1391
rect 695 -1392 696 -1391
rect 772 -1392 773 -1391
rect 796 -1392 797 -1391
rect 803 -1392 804 -1391
rect 44 -1394 45 -1393
rect 107 -1394 108 -1393
rect 121 -1394 122 -1393
rect 142 -1394 143 -1393
rect 156 -1394 157 -1393
rect 170 -1394 171 -1393
rect 177 -1394 178 -1393
rect 422 -1394 423 -1393
rect 457 -1394 458 -1393
rect 835 -1394 836 -1393
rect 51 -1396 52 -1395
rect 138 -1396 139 -1395
rect 163 -1396 164 -1395
rect 184 -1396 185 -1395
rect 226 -1396 227 -1395
rect 310 -1396 311 -1395
rect 324 -1396 325 -1395
rect 352 -1396 353 -1395
rect 394 -1396 395 -1395
rect 422 -1396 423 -1395
rect 450 -1396 451 -1395
rect 457 -1396 458 -1395
rect 478 -1396 479 -1395
rect 583 -1396 584 -1395
rect 590 -1396 591 -1395
rect 702 -1396 703 -1395
rect 709 -1396 710 -1395
rect 751 -1396 752 -1395
rect 51 -1398 52 -1397
rect 387 -1398 388 -1397
rect 394 -1398 395 -1397
rect 415 -1398 416 -1397
rect 488 -1398 489 -1397
rect 527 -1398 528 -1397
rect 551 -1398 552 -1397
rect 660 -1398 661 -1397
rect 674 -1398 675 -1397
rect 681 -1398 682 -1397
rect 58 -1400 59 -1399
rect 61 -1400 62 -1399
rect 75 -1400 76 -1399
rect 166 -1400 167 -1399
rect 226 -1400 227 -1399
rect 380 -1400 381 -1399
rect 404 -1400 405 -1399
rect 709 -1400 710 -1399
rect 58 -1402 59 -1401
rect 65 -1402 66 -1401
rect 75 -1402 76 -1401
rect 205 -1402 206 -1401
rect 254 -1402 255 -1401
rect 275 -1402 276 -1401
rect 303 -1402 304 -1401
rect 387 -1402 388 -1401
rect 404 -1402 405 -1401
rect 695 -1402 696 -1401
rect 61 -1404 62 -1403
rect 65 -1404 66 -1403
rect 79 -1404 80 -1403
rect 177 -1404 178 -1403
rect 205 -1404 206 -1403
rect 299 -1404 300 -1403
rect 348 -1404 349 -1403
rect 534 -1404 535 -1403
rect 555 -1404 556 -1403
rect 716 -1404 717 -1403
rect 79 -1406 80 -1405
rect 128 -1406 129 -1405
rect 261 -1406 262 -1405
rect 303 -1406 304 -1405
rect 317 -1406 318 -1405
rect 716 -1406 717 -1405
rect 86 -1408 87 -1407
rect 100 -1408 101 -1407
rect 117 -1408 118 -1407
rect 478 -1408 479 -1407
rect 506 -1408 507 -1407
rect 625 -1408 626 -1407
rect 639 -1408 640 -1407
rect 688 -1408 689 -1407
rect 89 -1410 90 -1409
rect 247 -1410 248 -1409
rect 261 -1410 262 -1409
rect 268 -1410 269 -1409
rect 282 -1410 283 -1409
rect 317 -1410 318 -1409
rect 352 -1410 353 -1409
rect 516 -1410 517 -1409
rect 520 -1410 521 -1409
rect 590 -1410 591 -1409
rect 618 -1410 619 -1409
rect 653 -1410 654 -1409
rect 93 -1412 94 -1411
rect 611 -1412 612 -1411
rect 646 -1412 647 -1411
rect 723 -1412 724 -1411
rect 30 -1414 31 -1413
rect 93 -1414 94 -1413
rect 100 -1414 101 -1413
rect 240 -1414 241 -1413
rect 359 -1414 360 -1413
rect 450 -1414 451 -1413
rect 506 -1414 507 -1413
rect 611 -1414 612 -1413
rect 23 -1416 24 -1415
rect 30 -1416 31 -1415
rect 107 -1416 108 -1415
rect 117 -1416 118 -1415
rect 128 -1416 129 -1415
rect 198 -1416 199 -1415
rect 219 -1416 220 -1415
rect 282 -1416 283 -1415
rect 359 -1416 360 -1415
rect 373 -1416 374 -1415
rect 411 -1416 412 -1415
rect 415 -1416 416 -1415
rect 432 -1416 433 -1415
rect 555 -1416 556 -1415
rect 562 -1416 563 -1415
rect 632 -1416 633 -1415
rect 23 -1418 24 -1417
rect 471 -1418 472 -1417
rect 492 -1418 493 -1417
rect 632 -1418 633 -1417
rect 198 -1420 199 -1419
rect 289 -1420 290 -1419
rect 366 -1420 367 -1419
rect 492 -1420 493 -1419
rect 513 -1420 514 -1419
rect 618 -1420 619 -1419
rect 219 -1422 220 -1421
rect 429 -1422 430 -1421
rect 439 -1422 440 -1421
rect 513 -1422 514 -1421
rect 520 -1422 521 -1421
rect 691 -1422 692 -1421
rect 233 -1424 234 -1423
rect 289 -1424 290 -1423
rect 334 -1424 335 -1423
rect 366 -1424 367 -1423
rect 527 -1424 528 -1423
rect 548 -1424 549 -1423
rect 565 -1424 566 -1423
rect 660 -1424 661 -1423
rect 191 -1426 192 -1425
rect 233 -1426 234 -1425
rect 240 -1426 241 -1425
rect 254 -1426 255 -1425
rect 268 -1426 269 -1425
rect 373 -1426 374 -1425
rect 541 -1426 542 -1425
rect 639 -1426 640 -1425
rect 191 -1428 192 -1427
rect 765 -1428 766 -1427
rect 541 -1430 542 -1429
rect 705 -1430 706 -1429
rect 548 -1432 549 -1431
rect 681 -1432 682 -1431
rect 572 -1434 573 -1433
rect 667 -1434 668 -1433
rect 583 -1436 584 -1435
rect 604 -1436 605 -1435
rect 667 -1436 668 -1435
rect 768 -1436 769 -1435
rect 485 -1438 486 -1437
rect 604 -1438 605 -1437
rect 485 -1440 486 -1439
rect 569 -1440 570 -1439
rect 597 -1440 598 -1439
rect 646 -1440 647 -1439
rect 499 -1442 500 -1441
rect 597 -1442 598 -1441
rect 436 -1444 437 -1443
rect 499 -1444 500 -1443
rect 9 -1455 10 -1454
rect 96 -1455 97 -1454
rect 128 -1455 129 -1454
rect 548 -1455 549 -1454
rect 681 -1455 682 -1454
rect 789 -1455 790 -1454
rect 800 -1455 801 -1454
rect 814 -1455 815 -1454
rect 817 -1455 818 -1454
rect 828 -1455 829 -1454
rect 9 -1457 10 -1456
rect 779 -1457 780 -1456
rect 16 -1459 17 -1458
rect 436 -1459 437 -1458
rect 439 -1459 440 -1458
rect 632 -1459 633 -1458
rect 681 -1459 682 -1458
rect 737 -1459 738 -1458
rect 768 -1459 769 -1458
rect 807 -1459 808 -1458
rect 16 -1461 17 -1460
rect 471 -1461 472 -1460
rect 474 -1461 475 -1460
rect 751 -1461 752 -1460
rect 23 -1463 24 -1462
rect 138 -1463 139 -1462
rect 156 -1463 157 -1462
rect 723 -1463 724 -1462
rect 737 -1463 738 -1462
rect 772 -1463 773 -1462
rect 23 -1465 24 -1464
rect 163 -1465 164 -1464
rect 198 -1465 199 -1464
rect 380 -1465 381 -1464
rect 394 -1465 395 -1464
rect 422 -1465 423 -1464
rect 429 -1465 430 -1464
rect 604 -1465 605 -1464
rect 632 -1465 633 -1464
rect 667 -1465 668 -1464
rect 674 -1465 675 -1464
rect 723 -1465 724 -1464
rect 30 -1467 31 -1466
rect 184 -1467 185 -1466
rect 250 -1467 251 -1466
rect 418 -1467 419 -1466
rect 422 -1467 423 -1466
rect 492 -1467 493 -1466
rect 509 -1467 510 -1466
rect 688 -1467 689 -1466
rect 30 -1469 31 -1468
rect 180 -1469 181 -1468
rect 257 -1469 258 -1468
rect 611 -1469 612 -1468
rect 667 -1469 668 -1468
rect 716 -1469 717 -1468
rect 37 -1471 38 -1470
rect 166 -1471 167 -1470
rect 268 -1471 269 -1470
rect 296 -1471 297 -1470
rect 303 -1471 304 -1470
rect 471 -1471 472 -1470
rect 523 -1471 524 -1470
rect 625 -1471 626 -1470
rect 688 -1471 689 -1470
rect 744 -1471 745 -1470
rect 44 -1473 45 -1472
rect 117 -1473 118 -1472
rect 128 -1473 129 -1472
rect 142 -1473 143 -1472
rect 159 -1473 160 -1472
rect 408 -1473 409 -1472
rect 432 -1473 433 -1472
rect 639 -1473 640 -1472
rect 54 -1475 55 -1474
rect 716 -1475 717 -1474
rect 58 -1477 59 -1476
rect 72 -1477 73 -1476
rect 79 -1477 80 -1476
rect 82 -1477 83 -1476
rect 114 -1477 115 -1476
rect 138 -1477 139 -1476
rect 142 -1477 143 -1476
rect 177 -1477 178 -1476
rect 296 -1477 297 -1476
rect 369 -1477 370 -1476
rect 383 -1477 384 -1476
rect 611 -1477 612 -1476
rect 37 -1479 38 -1478
rect 383 -1479 384 -1478
rect 401 -1479 402 -1478
rect 457 -1479 458 -1478
rect 527 -1479 528 -1478
rect 604 -1479 605 -1478
rect 44 -1481 45 -1480
rect 177 -1481 178 -1480
rect 212 -1481 213 -1480
rect 457 -1481 458 -1480
rect 464 -1481 465 -1480
rect 527 -1481 528 -1480
rect 534 -1481 535 -1480
rect 537 -1481 538 -1480
rect 541 -1481 542 -1480
rect 625 -1481 626 -1480
rect 58 -1483 59 -1482
rect 86 -1483 87 -1482
rect 135 -1483 136 -1482
rect 156 -1483 157 -1482
rect 212 -1483 213 -1482
rect 254 -1483 255 -1482
rect 306 -1483 307 -1482
rect 730 -1483 731 -1482
rect 65 -1485 66 -1484
rect 124 -1485 125 -1484
rect 331 -1485 332 -1484
rect 345 -1485 346 -1484
rect 352 -1485 353 -1484
rect 506 -1485 507 -1484
rect 513 -1485 514 -1484
rect 541 -1485 542 -1484
rect 555 -1485 556 -1484
rect 744 -1485 745 -1484
rect 65 -1487 66 -1486
rect 149 -1487 150 -1486
rect 289 -1487 290 -1486
rect 345 -1487 346 -1486
rect 359 -1487 360 -1486
rect 429 -1487 430 -1486
rect 439 -1487 440 -1486
rect 646 -1487 647 -1486
rect 79 -1489 80 -1488
rect 100 -1489 101 -1488
rect 149 -1489 150 -1488
rect 219 -1489 220 -1488
rect 289 -1489 290 -1488
rect 373 -1489 374 -1488
rect 390 -1489 391 -1488
rect 464 -1489 465 -1488
rect 478 -1489 479 -1488
rect 513 -1489 514 -1488
rect 534 -1489 535 -1488
rect 618 -1489 619 -1488
rect 646 -1489 647 -1488
rect 835 -1489 836 -1488
rect 86 -1491 87 -1490
rect 275 -1491 276 -1490
rect 317 -1491 318 -1490
rect 352 -1491 353 -1490
rect 366 -1491 367 -1490
rect 492 -1491 493 -1490
rect 555 -1491 556 -1490
rect 583 -1491 584 -1490
rect 597 -1491 598 -1490
rect 751 -1491 752 -1490
rect 170 -1493 171 -1492
rect 219 -1493 220 -1492
rect 233 -1493 234 -1492
rect 275 -1493 276 -1492
rect 282 -1493 283 -1492
rect 317 -1493 318 -1492
rect 331 -1493 332 -1492
rect 576 -1493 577 -1492
rect 597 -1493 598 -1492
rect 730 -1493 731 -1492
rect 93 -1495 94 -1494
rect 170 -1495 171 -1494
rect 191 -1495 192 -1494
rect 373 -1495 374 -1494
rect 387 -1495 388 -1494
rect 478 -1495 479 -1494
rect 562 -1495 563 -1494
rect 674 -1495 675 -1494
rect 121 -1497 122 -1496
rect 191 -1497 192 -1496
rect 233 -1497 234 -1496
rect 271 -1497 272 -1496
rect 310 -1497 311 -1496
rect 387 -1497 388 -1496
rect 397 -1497 398 -1496
rect 576 -1497 577 -1496
rect 618 -1497 619 -1496
rect 653 -1497 654 -1496
rect 107 -1499 108 -1498
rect 121 -1499 122 -1498
rect 247 -1499 248 -1498
rect 310 -1499 311 -1498
rect 334 -1499 335 -1498
rect 660 -1499 661 -1498
rect 107 -1501 108 -1500
rect 187 -1501 188 -1500
rect 198 -1501 199 -1500
rect 247 -1501 248 -1500
rect 261 -1501 262 -1500
rect 282 -1501 283 -1500
rect 338 -1501 339 -1500
rect 401 -1501 402 -1500
rect 450 -1501 451 -1500
rect 639 -1501 640 -1500
rect 653 -1501 654 -1500
rect 695 -1501 696 -1500
rect 240 -1503 241 -1502
rect 261 -1503 262 -1502
rect 324 -1503 325 -1502
rect 338 -1503 339 -1502
rect 341 -1503 342 -1502
rect 583 -1503 584 -1502
rect 660 -1503 661 -1502
rect 702 -1503 703 -1502
rect 240 -1505 241 -1504
rect 404 -1505 405 -1504
rect 450 -1505 451 -1504
rect 499 -1505 500 -1504
rect 520 -1505 521 -1504
rect 562 -1505 563 -1504
rect 324 -1507 325 -1506
rect 443 -1507 444 -1506
rect 485 -1507 486 -1506
rect 520 -1507 521 -1506
rect 537 -1507 538 -1506
rect 695 -1507 696 -1506
rect 226 -1509 227 -1508
rect 443 -1509 444 -1508
rect 205 -1511 206 -1510
rect 226 -1511 227 -1510
rect 362 -1511 363 -1510
rect 702 -1511 703 -1510
rect 366 -1513 367 -1512
rect 709 -1513 710 -1512
rect 380 -1515 381 -1514
rect 709 -1515 710 -1514
rect 415 -1517 416 -1516
rect 499 -1517 500 -1516
rect 415 -1519 416 -1518
rect 590 -1519 591 -1518
rect 569 -1521 570 -1520
rect 590 -1521 591 -1520
rect 359 -1523 360 -1522
rect 569 -1523 570 -1522
rect 12 -1534 13 -1533
rect 16 -1534 17 -1533
rect 51 -1534 52 -1533
rect 205 -1534 206 -1533
rect 208 -1534 209 -1533
rect 261 -1534 262 -1533
rect 303 -1534 304 -1533
rect 317 -1534 318 -1533
rect 331 -1534 332 -1533
rect 436 -1534 437 -1533
rect 488 -1534 489 -1533
rect 744 -1534 745 -1533
rect 16 -1536 17 -1535
rect 212 -1536 213 -1535
rect 240 -1536 241 -1535
rect 324 -1536 325 -1535
rect 338 -1536 339 -1535
rect 471 -1536 472 -1535
rect 520 -1536 521 -1535
rect 604 -1536 605 -1535
rect 618 -1536 619 -1535
rect 667 -1536 668 -1535
rect 2 -1538 3 -1537
rect 324 -1538 325 -1537
rect 341 -1538 342 -1537
rect 667 -1538 668 -1537
rect 23 -1540 24 -1539
rect 205 -1540 206 -1539
rect 212 -1540 213 -1539
rect 289 -1540 290 -1539
rect 303 -1540 304 -1539
rect 639 -1540 640 -1539
rect 23 -1542 24 -1541
rect 345 -1542 346 -1541
rect 362 -1542 363 -1541
rect 443 -1542 444 -1541
rect 471 -1542 472 -1541
rect 702 -1542 703 -1541
rect 44 -1544 45 -1543
rect 331 -1544 332 -1543
rect 341 -1544 342 -1543
rect 499 -1544 500 -1543
rect 597 -1544 598 -1543
rect 737 -1544 738 -1543
rect 44 -1546 45 -1545
rect 569 -1546 570 -1545
rect 604 -1546 605 -1545
rect 653 -1546 654 -1545
rect 51 -1548 52 -1547
rect 128 -1548 129 -1547
rect 138 -1548 139 -1547
rect 478 -1548 479 -1547
rect 499 -1548 500 -1547
rect 751 -1548 752 -1547
rect 58 -1550 59 -1549
rect 96 -1550 97 -1549
rect 103 -1550 104 -1549
rect 191 -1550 192 -1549
rect 233 -1550 234 -1549
rect 478 -1550 479 -1549
rect 569 -1550 570 -1549
rect 632 -1550 633 -1549
rect 653 -1550 654 -1549
rect 709 -1550 710 -1549
rect 58 -1552 59 -1551
rect 170 -1552 171 -1551
rect 184 -1552 185 -1551
rect 275 -1552 276 -1551
rect 278 -1552 279 -1551
rect 597 -1552 598 -1551
rect 632 -1552 633 -1551
rect 688 -1552 689 -1551
rect 72 -1554 73 -1553
rect 100 -1554 101 -1553
rect 117 -1554 118 -1553
rect 121 -1554 122 -1553
rect 128 -1554 129 -1553
rect 320 -1554 321 -1553
rect 345 -1554 346 -1553
rect 541 -1554 542 -1553
rect 79 -1556 80 -1555
rect 89 -1556 90 -1555
rect 93 -1556 94 -1555
rect 114 -1556 115 -1555
rect 121 -1556 122 -1555
rect 296 -1556 297 -1555
rect 306 -1556 307 -1555
rect 457 -1556 458 -1555
rect 82 -1558 83 -1557
rect 254 -1558 255 -1557
rect 257 -1558 258 -1557
rect 548 -1558 549 -1557
rect 86 -1560 87 -1559
rect 268 -1560 269 -1559
rect 289 -1560 290 -1559
rect 408 -1560 409 -1559
rect 415 -1560 416 -1559
rect 646 -1560 647 -1559
rect 65 -1562 66 -1561
rect 408 -1562 409 -1561
rect 415 -1562 416 -1561
rect 422 -1562 423 -1561
rect 443 -1562 444 -1561
rect 534 -1562 535 -1561
rect 548 -1562 549 -1561
rect 600 -1562 601 -1561
rect 646 -1562 647 -1561
rect 695 -1562 696 -1561
rect 30 -1564 31 -1563
rect 65 -1564 66 -1563
rect 138 -1564 139 -1563
rect 219 -1564 220 -1563
rect 247 -1564 248 -1563
rect 401 -1564 402 -1563
rect 422 -1564 423 -1563
rect 506 -1564 507 -1563
rect 534 -1564 535 -1563
rect 611 -1564 612 -1563
rect 30 -1566 31 -1565
rect 583 -1566 584 -1565
rect 611 -1566 612 -1565
rect 660 -1566 661 -1565
rect 149 -1568 150 -1567
rect 163 -1568 164 -1567
rect 170 -1568 171 -1567
rect 236 -1568 237 -1567
rect 247 -1568 248 -1567
rect 282 -1568 283 -1567
rect 296 -1568 297 -1567
rect 513 -1568 514 -1567
rect 555 -1568 556 -1567
rect 583 -1568 584 -1567
rect 660 -1568 661 -1567
rect 716 -1568 717 -1567
rect 152 -1570 153 -1569
rect 352 -1570 353 -1569
rect 362 -1570 363 -1569
rect 541 -1570 542 -1569
rect 37 -1572 38 -1571
rect 352 -1572 353 -1571
rect 366 -1572 367 -1571
rect 492 -1572 493 -1571
rect 37 -1574 38 -1573
rect 107 -1574 108 -1573
rect 184 -1574 185 -1573
rect 198 -1574 199 -1573
rect 219 -1574 220 -1573
rect 639 -1574 640 -1573
rect 9 -1576 10 -1575
rect 107 -1576 108 -1575
rect 177 -1576 178 -1575
rect 198 -1576 199 -1575
rect 250 -1576 251 -1575
rect 373 -1576 374 -1575
rect 380 -1576 381 -1575
rect 450 -1576 451 -1575
rect 457 -1576 458 -1575
rect 576 -1576 577 -1575
rect 114 -1578 115 -1577
rect 380 -1578 381 -1577
rect 387 -1578 388 -1577
rect 674 -1578 675 -1577
rect 156 -1580 157 -1579
rect 177 -1580 178 -1579
rect 187 -1580 188 -1579
rect 191 -1580 192 -1579
rect 261 -1580 262 -1579
rect 310 -1580 311 -1579
rect 313 -1580 314 -1579
rect 429 -1580 430 -1579
rect 439 -1580 440 -1579
rect 506 -1580 507 -1579
rect 674 -1580 675 -1579
rect 723 -1580 724 -1579
rect 142 -1582 143 -1581
rect 156 -1582 157 -1581
rect 275 -1582 276 -1581
rect 373 -1582 374 -1581
rect 401 -1582 402 -1581
rect 527 -1582 528 -1581
rect 282 -1584 283 -1583
rect 310 -1584 311 -1583
rect 334 -1584 335 -1583
rect 513 -1584 514 -1583
rect 306 -1586 307 -1585
rect 527 -1586 528 -1585
rect 418 -1588 419 -1587
rect 450 -1588 451 -1587
rect 485 -1588 486 -1587
rect 576 -1588 577 -1587
rect 387 -1590 388 -1589
rect 485 -1590 486 -1589
rect 492 -1590 493 -1589
rect 590 -1590 591 -1589
rect 411 -1592 412 -1591
rect 590 -1592 591 -1591
rect 429 -1594 430 -1593
rect 464 -1594 465 -1593
rect 464 -1596 465 -1595
rect 562 -1596 563 -1595
rect 562 -1598 563 -1597
rect 625 -1598 626 -1597
rect 625 -1600 626 -1599
rect 681 -1600 682 -1599
rect 681 -1602 682 -1601
rect 730 -1602 731 -1601
rect 5 -1613 6 -1612
rect 324 -1613 325 -1612
rect 359 -1613 360 -1612
rect 471 -1613 472 -1612
rect 485 -1613 486 -1612
rect 520 -1613 521 -1612
rect 558 -1613 559 -1612
rect 646 -1613 647 -1612
rect 9 -1615 10 -1614
rect 156 -1615 157 -1614
rect 187 -1615 188 -1614
rect 198 -1615 199 -1614
rect 226 -1615 227 -1614
rect 278 -1615 279 -1614
rect 317 -1615 318 -1614
rect 499 -1615 500 -1614
rect 520 -1615 521 -1614
rect 576 -1615 577 -1614
rect 625 -1615 626 -1614
rect 649 -1615 650 -1614
rect 23 -1617 24 -1616
rect 79 -1617 80 -1616
rect 82 -1617 83 -1616
rect 639 -1617 640 -1616
rect 23 -1619 24 -1618
rect 110 -1619 111 -1618
rect 114 -1619 115 -1618
rect 299 -1619 300 -1618
rect 359 -1619 360 -1618
rect 534 -1619 535 -1618
rect 30 -1621 31 -1620
rect 324 -1621 325 -1620
rect 362 -1621 363 -1620
rect 394 -1621 395 -1620
rect 401 -1621 402 -1620
rect 408 -1621 409 -1620
rect 411 -1621 412 -1620
rect 632 -1621 633 -1620
rect 30 -1623 31 -1622
rect 219 -1623 220 -1622
rect 233 -1623 234 -1622
rect 247 -1623 248 -1622
rect 254 -1623 255 -1622
rect 317 -1623 318 -1622
rect 366 -1623 367 -1622
rect 464 -1623 465 -1622
rect 478 -1623 479 -1622
rect 499 -1623 500 -1622
rect 534 -1623 535 -1622
rect 604 -1623 605 -1622
rect 16 -1625 17 -1624
rect 464 -1625 465 -1624
rect 16 -1627 17 -1626
rect 138 -1627 139 -1626
rect 152 -1627 153 -1626
rect 254 -1627 255 -1626
rect 268 -1627 269 -1626
rect 310 -1627 311 -1626
rect 373 -1627 374 -1626
rect 478 -1627 479 -1626
rect 37 -1629 38 -1628
rect 100 -1629 101 -1628
rect 128 -1629 129 -1628
rect 156 -1629 157 -1628
rect 170 -1629 171 -1628
rect 226 -1629 227 -1628
rect 240 -1629 241 -1628
rect 268 -1629 269 -1628
rect 376 -1629 377 -1628
rect 387 -1629 388 -1628
rect 394 -1629 395 -1628
rect 506 -1629 507 -1628
rect 37 -1631 38 -1630
rect 306 -1631 307 -1630
rect 380 -1631 381 -1630
rect 471 -1631 472 -1630
rect 506 -1631 507 -1630
rect 611 -1631 612 -1630
rect 65 -1633 66 -1632
rect 275 -1633 276 -1632
rect 292 -1633 293 -1632
rect 611 -1633 612 -1632
rect 58 -1635 59 -1634
rect 65 -1635 66 -1634
rect 72 -1635 73 -1634
rect 142 -1635 143 -1634
rect 173 -1635 174 -1634
rect 198 -1635 199 -1634
rect 205 -1635 206 -1634
rect 247 -1635 248 -1634
rect 275 -1635 276 -1634
rect 352 -1635 353 -1634
rect 380 -1635 381 -1634
rect 429 -1635 430 -1634
rect 436 -1635 437 -1634
rect 457 -1635 458 -1634
rect 58 -1637 59 -1636
rect 191 -1637 192 -1636
rect 205 -1637 206 -1636
rect 369 -1637 370 -1636
rect 401 -1637 402 -1636
rect 422 -1637 423 -1636
rect 429 -1637 430 -1636
rect 450 -1637 451 -1636
rect 457 -1637 458 -1636
rect 555 -1637 556 -1636
rect 47 -1639 48 -1638
rect 191 -1639 192 -1638
rect 212 -1639 213 -1638
rect 233 -1639 234 -1638
rect 296 -1639 297 -1638
rect 387 -1639 388 -1638
rect 408 -1639 409 -1638
rect 660 -1639 661 -1638
rect 51 -1641 52 -1640
rect 422 -1641 423 -1640
rect 439 -1641 440 -1640
rect 590 -1641 591 -1640
rect 660 -1641 661 -1640
rect 674 -1641 675 -1640
rect 51 -1643 52 -1642
rect 338 -1643 339 -1642
rect 443 -1643 444 -1642
rect 597 -1643 598 -1642
rect 86 -1645 87 -1644
rect 149 -1645 150 -1644
rect 184 -1645 185 -1644
rect 219 -1645 220 -1644
rect 296 -1645 297 -1644
rect 576 -1645 577 -1644
rect 597 -1645 598 -1644
rect 681 -1645 682 -1644
rect 72 -1647 73 -1646
rect 86 -1647 87 -1646
rect 89 -1647 90 -1646
rect 653 -1647 654 -1646
rect 677 -1647 678 -1646
rect 681 -1647 682 -1646
rect 93 -1649 94 -1648
rect 117 -1649 118 -1648
rect 128 -1649 129 -1648
rect 177 -1649 178 -1648
rect 194 -1649 195 -1648
rect 590 -1649 591 -1648
rect 93 -1651 94 -1650
rect 121 -1651 122 -1650
rect 135 -1651 136 -1650
rect 177 -1651 178 -1650
rect 212 -1651 213 -1650
rect 261 -1651 262 -1650
rect 331 -1651 332 -1650
rect 338 -1651 339 -1650
rect 443 -1651 444 -1650
rect 513 -1651 514 -1650
rect 107 -1653 108 -1652
rect 135 -1653 136 -1652
rect 446 -1653 447 -1652
rect 555 -1653 556 -1652
rect 114 -1655 115 -1654
rect 170 -1655 171 -1654
rect 450 -1655 451 -1654
rect 541 -1655 542 -1654
rect 121 -1657 122 -1656
rect 289 -1657 290 -1656
rect 320 -1657 321 -1656
rect 541 -1657 542 -1656
rect 282 -1659 283 -1658
rect 289 -1659 290 -1658
rect 513 -1659 514 -1658
rect 562 -1659 563 -1658
rect 282 -1661 283 -1660
rect 415 -1661 416 -1660
rect 548 -1661 549 -1660
rect 562 -1661 563 -1660
rect 345 -1663 346 -1662
rect 415 -1663 416 -1662
rect 548 -1663 549 -1662
rect 569 -1663 570 -1662
rect 345 -1665 346 -1664
rect 492 -1665 493 -1664
rect 569 -1665 570 -1664
rect 618 -1665 619 -1664
rect 492 -1667 493 -1666
rect 527 -1667 528 -1666
rect 527 -1669 528 -1668
rect 583 -1669 584 -1668
rect 583 -1671 584 -1670
rect 667 -1671 668 -1670
rect 16 -1682 17 -1681
rect 86 -1682 87 -1681
rect 107 -1682 108 -1681
rect 159 -1682 160 -1681
rect 170 -1682 171 -1681
rect 177 -1682 178 -1681
rect 187 -1682 188 -1681
rect 422 -1682 423 -1681
rect 446 -1682 447 -1681
rect 492 -1682 493 -1681
rect 506 -1682 507 -1681
rect 653 -1682 654 -1681
rect 674 -1682 675 -1681
rect 681 -1682 682 -1681
rect 16 -1684 17 -1683
rect 93 -1684 94 -1683
rect 145 -1684 146 -1683
rect 296 -1684 297 -1683
rect 306 -1684 307 -1683
rect 471 -1684 472 -1683
rect 534 -1684 535 -1683
rect 579 -1684 580 -1683
rect 649 -1684 650 -1683
rect 660 -1684 661 -1683
rect 23 -1686 24 -1685
rect 142 -1686 143 -1685
rect 156 -1686 157 -1685
rect 191 -1686 192 -1685
rect 212 -1686 213 -1685
rect 261 -1686 262 -1685
rect 264 -1686 265 -1685
rect 464 -1686 465 -1685
rect 471 -1686 472 -1685
rect 513 -1686 514 -1685
rect 548 -1686 549 -1685
rect 621 -1686 622 -1685
rect 23 -1688 24 -1687
rect 345 -1688 346 -1687
rect 352 -1688 353 -1687
rect 590 -1688 591 -1687
rect 30 -1690 31 -1689
rect 226 -1690 227 -1689
rect 243 -1690 244 -1689
rect 324 -1690 325 -1689
rect 331 -1690 332 -1689
rect 541 -1690 542 -1689
rect 569 -1690 570 -1689
rect 618 -1690 619 -1689
rect 37 -1692 38 -1691
rect 313 -1692 314 -1691
rect 317 -1692 318 -1691
rect 359 -1692 360 -1691
rect 376 -1692 377 -1691
rect 499 -1692 500 -1691
rect 597 -1692 598 -1691
rect 618 -1692 619 -1691
rect 9 -1694 10 -1693
rect 317 -1694 318 -1693
rect 320 -1694 321 -1693
rect 408 -1694 409 -1693
rect 499 -1694 500 -1693
rect 527 -1694 528 -1693
rect 9 -1696 10 -1695
rect 128 -1696 129 -1695
rect 173 -1696 174 -1695
rect 334 -1696 335 -1695
rect 338 -1696 339 -1695
rect 576 -1696 577 -1695
rect 40 -1698 41 -1697
rect 198 -1698 199 -1697
rect 212 -1698 213 -1697
rect 275 -1698 276 -1697
rect 282 -1698 283 -1697
rect 355 -1698 356 -1697
rect 390 -1698 391 -1697
rect 443 -1698 444 -1697
rect 527 -1698 528 -1697
rect 611 -1698 612 -1697
rect 44 -1700 45 -1699
rect 131 -1700 132 -1699
rect 187 -1700 188 -1699
rect 236 -1700 237 -1699
rect 247 -1700 248 -1699
rect 289 -1700 290 -1699
rect 292 -1700 293 -1699
rect 296 -1700 297 -1699
rect 310 -1700 311 -1699
rect 359 -1700 360 -1699
rect 408 -1700 409 -1699
rect 436 -1700 437 -1699
rect 47 -1702 48 -1701
rect 58 -1702 59 -1701
rect 65 -1702 66 -1701
rect 261 -1702 262 -1701
rect 271 -1702 272 -1701
rect 464 -1702 465 -1701
rect 51 -1704 52 -1703
rect 257 -1704 258 -1703
rect 275 -1704 276 -1703
rect 394 -1704 395 -1703
rect 436 -1704 437 -1703
rect 450 -1704 451 -1703
rect 58 -1706 59 -1705
rect 520 -1706 521 -1705
rect 65 -1708 66 -1707
rect 128 -1708 129 -1707
rect 198 -1708 199 -1707
rect 233 -1708 234 -1707
rect 247 -1708 248 -1707
rect 373 -1708 374 -1707
rect 380 -1708 381 -1707
rect 394 -1708 395 -1707
rect 520 -1708 521 -1707
rect 562 -1708 563 -1707
rect 72 -1710 73 -1709
rect 124 -1710 125 -1709
rect 219 -1710 220 -1709
rect 226 -1710 227 -1709
rect 250 -1710 251 -1709
rect 492 -1710 493 -1709
rect 72 -1712 73 -1711
rect 205 -1712 206 -1711
rect 254 -1712 255 -1711
rect 324 -1712 325 -1711
rect 331 -1712 332 -1711
rect 415 -1712 416 -1711
rect 79 -1714 80 -1713
rect 289 -1714 290 -1713
rect 310 -1714 311 -1713
rect 478 -1714 479 -1713
rect 79 -1716 80 -1715
rect 268 -1716 269 -1715
rect 282 -1716 283 -1715
rect 429 -1716 430 -1715
rect 86 -1718 87 -1717
rect 114 -1718 115 -1717
rect 121 -1718 122 -1717
rect 233 -1718 234 -1717
rect 240 -1718 241 -1717
rect 478 -1718 479 -1717
rect 107 -1720 108 -1719
rect 142 -1720 143 -1719
rect 149 -1720 150 -1719
rect 219 -1720 220 -1719
rect 268 -1720 269 -1719
rect 366 -1720 367 -1719
rect 373 -1720 374 -1719
rect 422 -1720 423 -1719
rect 429 -1720 430 -1719
rect 485 -1720 486 -1719
rect 114 -1722 115 -1721
rect 135 -1722 136 -1721
rect 345 -1722 346 -1721
rect 401 -1722 402 -1721
rect 485 -1722 486 -1721
rect 555 -1722 556 -1721
rect 121 -1724 122 -1723
rect 380 -1724 381 -1723
rect 401 -1724 402 -1723
rect 457 -1724 458 -1723
rect 555 -1724 556 -1723
rect 583 -1724 584 -1723
rect 135 -1726 136 -1725
rect 163 -1726 164 -1725
rect 303 -1726 304 -1725
rect 457 -1726 458 -1725
rect 163 -1728 164 -1727
rect 184 -1728 185 -1727
rect 362 -1728 363 -1727
rect 415 -1728 416 -1727
rect 16 -1739 17 -1738
rect 152 -1739 153 -1738
rect 156 -1739 157 -1738
rect 240 -1739 241 -1738
rect 254 -1739 255 -1738
rect 257 -1739 258 -1738
rect 261 -1739 262 -1738
rect 352 -1739 353 -1738
rect 418 -1739 419 -1738
rect 534 -1739 535 -1738
rect 548 -1739 549 -1738
rect 555 -1739 556 -1738
rect 632 -1739 633 -1738
rect 653 -1739 654 -1738
rect 670 -1739 671 -1738
rect 674 -1739 675 -1738
rect 23 -1741 24 -1740
rect 362 -1741 363 -1740
rect 422 -1741 423 -1740
rect 453 -1741 454 -1740
rect 460 -1741 461 -1740
rect 520 -1741 521 -1740
rect 37 -1743 38 -1742
rect 107 -1743 108 -1742
rect 114 -1743 115 -1742
rect 177 -1743 178 -1742
rect 208 -1743 209 -1742
rect 296 -1743 297 -1742
rect 331 -1743 332 -1742
rect 352 -1743 353 -1742
rect 408 -1743 409 -1742
rect 460 -1743 461 -1742
rect 471 -1743 472 -1742
rect 513 -1743 514 -1742
rect 44 -1745 45 -1744
rect 310 -1745 311 -1744
rect 334 -1745 335 -1744
rect 492 -1745 493 -1744
rect 51 -1747 52 -1746
rect 292 -1747 293 -1746
rect 296 -1747 297 -1746
rect 366 -1747 367 -1746
rect 422 -1747 423 -1746
rect 478 -1747 479 -1746
rect 51 -1749 52 -1748
rect 135 -1749 136 -1748
rect 145 -1749 146 -1748
rect 219 -1749 220 -1748
rect 226 -1749 227 -1748
rect 243 -1749 244 -1748
rect 282 -1749 283 -1748
rect 317 -1749 318 -1748
rect 338 -1749 339 -1748
rect 401 -1749 402 -1748
rect 429 -1749 430 -1748
rect 488 -1749 489 -1748
rect 58 -1751 59 -1750
rect 355 -1751 356 -1750
rect 429 -1751 430 -1750
rect 464 -1751 465 -1750
rect 471 -1751 472 -1750
rect 527 -1751 528 -1750
rect 65 -1753 66 -1752
rect 93 -1753 94 -1752
rect 117 -1753 118 -1752
rect 205 -1753 206 -1752
rect 212 -1753 213 -1752
rect 268 -1753 269 -1752
rect 289 -1753 290 -1752
rect 324 -1753 325 -1752
rect 345 -1753 346 -1752
rect 366 -1753 367 -1752
rect 394 -1753 395 -1752
rect 464 -1753 465 -1752
rect 478 -1753 479 -1752
rect 485 -1753 486 -1752
rect 499 -1753 500 -1752
rect 527 -1753 528 -1752
rect 72 -1755 73 -1754
rect 135 -1755 136 -1754
rect 152 -1755 153 -1754
rect 191 -1755 192 -1754
rect 219 -1755 220 -1754
rect 303 -1755 304 -1754
rect 310 -1755 311 -1754
rect 404 -1755 405 -1754
rect 436 -1755 437 -1754
rect 520 -1755 521 -1754
rect 72 -1757 73 -1756
rect 79 -1757 80 -1756
rect 86 -1757 87 -1756
rect 103 -1757 104 -1756
rect 124 -1757 125 -1756
rect 142 -1757 143 -1756
rect 159 -1757 160 -1756
rect 191 -1757 192 -1756
rect 268 -1757 269 -1756
rect 380 -1757 381 -1756
rect 65 -1759 66 -1758
rect 159 -1759 160 -1758
rect 163 -1759 164 -1758
rect 226 -1759 227 -1758
rect 275 -1759 276 -1758
rect 345 -1759 346 -1758
rect 86 -1761 87 -1760
rect 121 -1761 122 -1760
rect 128 -1761 129 -1760
rect 250 -1761 251 -1760
rect 324 -1761 325 -1760
rect 415 -1761 416 -1760
rect 93 -1763 94 -1762
rect 107 -1763 108 -1762
rect 163 -1763 164 -1762
rect 261 -1763 262 -1762
rect 173 -1765 174 -1764
rect 198 -1765 199 -1764
rect 233 -1765 234 -1764
rect 275 -1765 276 -1764
rect 9 -1767 10 -1766
rect 198 -1767 199 -1766
rect 170 -1769 171 -1768
rect 233 -1769 234 -1768
rect 51 -1780 52 -1779
rect 184 -1780 185 -1779
rect 198 -1780 199 -1779
rect 250 -1780 251 -1779
rect 254 -1780 255 -1779
rect 289 -1780 290 -1779
rect 317 -1780 318 -1779
rect 383 -1780 384 -1779
rect 387 -1780 388 -1779
rect 429 -1780 430 -1779
rect 464 -1780 465 -1779
rect 485 -1780 486 -1779
rect 499 -1780 500 -1779
rect 534 -1780 535 -1779
rect 541 -1780 542 -1779
rect 548 -1780 549 -1779
rect 614 -1780 615 -1779
rect 632 -1780 633 -1779
rect 51 -1782 52 -1781
rect 61 -1782 62 -1781
rect 72 -1782 73 -1781
rect 334 -1782 335 -1781
rect 345 -1782 346 -1781
rect 411 -1782 412 -1781
rect 467 -1782 468 -1781
rect 520 -1782 521 -1781
rect 618 -1782 619 -1781
rect 639 -1782 640 -1781
rect 86 -1784 87 -1783
rect 103 -1784 104 -1783
rect 110 -1784 111 -1783
rect 212 -1784 213 -1783
rect 247 -1784 248 -1783
rect 324 -1784 325 -1783
rect 352 -1784 353 -1783
rect 418 -1784 419 -1783
rect 478 -1784 479 -1783
rect 502 -1784 503 -1783
rect 513 -1784 514 -1783
rect 562 -1784 563 -1783
rect 93 -1786 94 -1785
rect 103 -1786 104 -1785
rect 117 -1786 118 -1785
rect 128 -1786 129 -1785
rect 135 -1786 136 -1785
rect 149 -1786 150 -1785
rect 156 -1786 157 -1785
rect 226 -1786 227 -1785
rect 264 -1786 265 -1785
rect 310 -1786 311 -1785
rect 338 -1786 339 -1785
rect 352 -1786 353 -1785
rect 366 -1786 367 -1785
rect 418 -1786 419 -1785
rect 520 -1786 521 -1785
rect 527 -1786 528 -1785
rect 65 -1788 66 -1787
rect 117 -1788 118 -1787
rect 124 -1788 125 -1787
rect 240 -1788 241 -1787
rect 296 -1788 297 -1787
rect 310 -1788 311 -1787
rect 373 -1788 374 -1787
rect 422 -1788 423 -1787
rect 89 -1790 90 -1789
rect 135 -1790 136 -1789
rect 138 -1790 139 -1789
rect 156 -1790 157 -1789
rect 163 -1790 164 -1789
rect 268 -1790 269 -1789
rect 142 -1792 143 -1791
rect 159 -1792 160 -1791
rect 173 -1792 174 -1791
rect 191 -1792 192 -1791
rect 205 -1792 206 -1791
rect 219 -1792 220 -1791
rect 37 -1794 38 -1793
rect 142 -1794 143 -1793
rect 177 -1794 178 -1793
rect 233 -1794 234 -1793
rect 233 -1796 234 -1795
rect 261 -1796 262 -1795
rect 131 -1798 132 -1797
rect 261 -1798 262 -1797
rect 51 -1809 52 -1808
rect 61 -1809 62 -1808
rect 145 -1809 146 -1808
rect 205 -1809 206 -1808
rect 233 -1809 234 -1808
rect 271 -1809 272 -1808
rect 352 -1809 353 -1808
rect 418 -1809 419 -1808
rect 471 -1809 472 -1808
rect 478 -1809 479 -1808
rect 520 -1809 521 -1808
rect 527 -1809 528 -1808
rect 149 -1811 150 -1810
rect 184 -1811 185 -1810
rect 156 -1813 157 -1812
rect 177 -1813 178 -1812
rect 180 -1813 181 -1812
rect 261 -1813 262 -1812
<< metal2 >>
rect 58 -7 59 1
rect 93 -7 94 1
rect 114 -7 115 1
rect 142 -7 143 1
rect 152 -7 153 1
rect 170 -7 171 1
rect 177 -7 178 1
rect 212 -7 213 1
rect 257 -7 258 1
rect 261 -7 262 1
rect 124 -7 125 -1
rect 240 -7 241 -1
rect 128 -7 129 -3
rect 135 -7 136 -3
rect 156 -7 157 -3
rect 163 -7 164 -3
rect 184 -7 185 -3
rect 191 -7 192 -3
rect 198 -7 199 -3
rect 236 -7 237 -3
rect 205 -7 206 -5
rect 338 -7 339 -5
rect 44 -34 45 -16
rect 47 -17 48 -15
rect 72 -34 73 -16
rect 93 -17 94 -15
rect 103 -34 104 -16
rect 275 -34 276 -16
rect 285 -34 286 -16
rect 345 -34 346 -16
rect 79 -34 80 -18
rect 191 -34 192 -18
rect 205 -19 206 -15
rect 317 -34 318 -18
rect 338 -19 339 -15
rect 387 -34 388 -18
rect 114 -21 115 -15
rect 131 -34 132 -20
rect 177 -21 178 -15
rect 198 -21 199 -15
rect 205 -34 206 -20
rect 324 -34 325 -20
rect 124 -34 125 -22
rect 212 -23 213 -15
rect 222 -23 223 -15
rect 240 -23 241 -15
rect 247 -34 248 -22
rect 334 -34 335 -22
rect 128 -25 129 -15
rect 135 -34 136 -24
rect 149 -34 150 -24
rect 177 -34 178 -24
rect 184 -25 185 -15
rect 219 -34 220 -24
rect 240 -34 241 -24
rect 261 -25 262 -15
rect 271 -34 272 -24
rect 352 -34 353 -24
rect 93 -34 94 -26
rect 128 -34 129 -26
rect 163 -27 164 -15
rect 198 -34 199 -26
rect 212 -34 213 -26
rect 226 -27 227 -15
rect 254 -34 255 -26
rect 282 -34 283 -26
rect 289 -27 290 -15
rect 296 -34 297 -26
rect 313 -34 314 -26
rect 338 -34 339 -26
rect 170 -29 171 -15
rect 184 -34 185 -28
rect 226 -34 227 -28
rect 233 -29 234 -15
rect 142 -34 143 -30
rect 233 -34 234 -30
rect 163 -34 164 -32
rect 170 -34 171 -32
rect 16 -69 17 -43
rect 240 -44 241 -42
rect 254 -44 255 -42
rect 341 -69 342 -43
rect 345 -44 346 -42
rect 436 -69 437 -43
rect 23 -69 24 -45
rect 117 -46 118 -42
rect 128 -69 129 -45
rect 156 -46 157 -42
rect 163 -69 164 -45
rect 170 -46 171 -42
rect 191 -46 192 -42
rect 222 -69 223 -45
rect 233 -46 234 -42
rect 310 -69 311 -45
rect 317 -46 318 -42
rect 380 -69 381 -45
rect 387 -46 388 -42
rect 408 -69 409 -45
rect 44 -69 45 -47
rect 58 -69 59 -47
rect 65 -69 66 -47
rect 107 -48 108 -42
rect 114 -69 115 -47
rect 121 -69 122 -47
rect 135 -48 136 -42
rect 142 -69 143 -47
rect 156 -69 157 -47
rect 194 -69 195 -47
rect 205 -48 206 -42
rect 219 -48 220 -42
rect 247 -48 248 -42
rect 254 -69 255 -47
rect 275 -48 276 -42
rect 331 -69 332 -47
rect 338 -48 339 -42
rect 422 -69 423 -47
rect 51 -50 52 -42
rect 345 -69 346 -49
rect 352 -50 353 -42
rect 401 -69 402 -49
rect 404 -50 405 -42
rect 415 -69 416 -49
rect 61 -69 62 -51
rect 205 -69 206 -51
rect 208 -52 209 -42
rect 226 -52 227 -42
rect 268 -69 269 -51
rect 275 -69 276 -51
rect 282 -69 283 -51
rect 317 -69 318 -51
rect 324 -52 325 -42
rect 387 -69 388 -51
rect 72 -54 73 -42
rect 152 -69 153 -53
rect 170 -69 171 -53
rect 180 -69 181 -53
rect 184 -54 185 -42
rect 226 -69 227 -53
rect 296 -54 297 -42
rect 359 -69 360 -53
rect 373 -69 374 -53
rect 394 -69 395 -53
rect 82 -69 83 -55
rect 135 -69 136 -55
rect 184 -69 185 -55
rect 240 -69 241 -55
rect 299 -69 300 -55
rect 366 -69 367 -55
rect 86 -69 87 -57
rect 177 -58 178 -42
rect 212 -58 213 -42
rect 233 -69 234 -57
rect 93 -60 94 -42
rect 324 -69 325 -59
rect 93 -69 94 -61
rect 292 -62 293 -42
rect 100 -69 101 -63
rect 110 -69 111 -63
rect 177 -69 178 -63
rect 198 -64 199 -42
rect 212 -69 213 -63
rect 271 -64 272 -42
rect 198 -69 199 -65
rect 289 -69 290 -65
rect 261 -69 262 -67
rect 271 -69 272 -67
rect 23 -79 24 -77
rect 198 -79 199 -77
rect 205 -79 206 -77
rect 506 -122 507 -78
rect 37 -81 38 -77
rect 219 -122 220 -80
rect 233 -81 234 -77
rect 247 -81 248 -77
rect 250 -81 251 -77
rect 464 -122 465 -80
rect 44 -83 45 -77
rect 296 -122 297 -82
rect 303 -83 304 -77
rect 394 -122 395 -82
rect 397 -83 398 -77
rect 457 -122 458 -82
rect 58 -122 59 -84
rect 156 -85 157 -77
rect 170 -85 171 -77
rect 205 -122 206 -84
rect 208 -85 209 -77
rect 240 -85 241 -77
rect 254 -85 255 -77
rect 268 -122 269 -84
rect 275 -85 276 -77
rect 303 -122 304 -84
rect 373 -85 374 -77
rect 429 -122 430 -84
rect 436 -85 437 -77
rect 513 -122 514 -84
rect 65 -87 66 -77
rect 152 -87 153 -77
rect 156 -122 157 -86
rect 247 -122 248 -86
rect 254 -122 255 -86
rect 317 -87 318 -77
rect 345 -87 346 -77
rect 436 -122 437 -86
rect 72 -89 73 -77
rect 114 -122 115 -88
rect 121 -89 122 -77
rect 198 -122 199 -88
rect 222 -89 223 -77
rect 317 -122 318 -88
rect 338 -122 339 -88
rect 345 -122 346 -88
rect 380 -89 381 -77
rect 471 -122 472 -88
rect 79 -122 80 -90
rect 261 -91 262 -77
rect 275 -122 276 -90
rect 310 -91 311 -77
rect 387 -91 388 -77
rect 492 -122 493 -90
rect 16 -93 17 -77
rect 261 -122 262 -92
rect 285 -122 286 -92
rect 450 -122 451 -92
rect 86 -122 87 -94
rect 100 -95 101 -77
rect 107 -122 108 -94
rect 212 -95 213 -77
rect 292 -122 293 -94
rect 422 -95 423 -77
rect 93 -97 94 -77
rect 443 -122 444 -96
rect 93 -122 94 -98
rect 282 -122 283 -98
rect 310 -122 311 -98
rect 334 -122 335 -98
rect 380 -122 381 -98
rect 422 -122 423 -98
rect 128 -101 129 -77
rect 194 -101 195 -77
rect 212 -122 213 -100
rect 306 -101 307 -77
rect 401 -101 402 -77
rect 499 -122 500 -100
rect 128 -122 129 -102
rect 299 -103 300 -77
rect 359 -103 360 -77
rect 401 -122 402 -102
rect 408 -103 409 -77
rect 485 -122 486 -102
rect 135 -105 136 -77
rect 191 -122 192 -104
rect 324 -105 325 -77
rect 359 -122 360 -104
rect 366 -105 367 -77
rect 408 -122 409 -104
rect 415 -105 416 -77
rect 478 -122 479 -104
rect 149 -107 150 -77
rect 387 -122 388 -106
rect 149 -122 150 -108
rect 163 -109 164 -77
rect 173 -122 174 -108
rect 289 -109 290 -77
rect 331 -109 332 -77
rect 366 -122 367 -108
rect 373 -122 374 -108
rect 415 -122 416 -108
rect 121 -122 122 -110
rect 289 -122 290 -110
rect 331 -122 332 -110
rect 520 -122 521 -110
rect 177 -122 178 -112
rect 233 -122 234 -112
rect 187 -115 188 -77
rect 226 -115 227 -77
rect 142 -117 143 -77
rect 226 -122 227 -116
rect 142 -122 143 -118
rect 184 -119 185 -77
rect 163 -122 164 -120
rect 187 -122 188 -120
rect 12 -197 13 -131
rect 72 -197 73 -131
rect 75 -132 76 -130
rect 506 -132 507 -130
rect 520 -132 521 -130
rect 660 -197 661 -131
rect 51 -134 52 -130
rect 177 -134 178 -130
rect 180 -134 181 -130
rect 359 -134 360 -130
rect 373 -134 374 -130
rect 376 -172 377 -133
rect 383 -134 384 -130
rect 464 -134 465 -130
rect 471 -134 472 -130
rect 618 -197 619 -133
rect 58 -136 59 -130
rect 285 -197 286 -135
rect 296 -136 297 -130
rect 331 -197 332 -135
rect 334 -136 335 -130
rect 443 -136 444 -130
rect 457 -136 458 -130
rect 583 -197 584 -135
rect 58 -197 59 -137
rect 243 -138 244 -130
rect 250 -197 251 -137
rect 268 -138 269 -130
rect 282 -138 283 -130
rect 401 -138 402 -130
rect 415 -138 416 -130
rect 569 -197 570 -137
rect 65 -140 66 -130
rect 65 -197 66 -139
rect 65 -140 66 -130
rect 65 -197 66 -139
rect 79 -140 80 -130
rect 401 -197 402 -139
rect 422 -140 423 -130
rect 443 -197 444 -139
rect 478 -140 479 -130
rect 639 -197 640 -139
rect 79 -197 80 -141
rect 103 -142 104 -130
rect 121 -142 122 -130
rect 527 -197 528 -141
rect 44 -144 45 -130
rect 121 -197 122 -143
rect 128 -144 129 -130
rect 380 -197 381 -143
rect 390 -197 391 -143
rect 653 -197 654 -143
rect 44 -197 45 -145
rect 187 -146 188 -130
rect 240 -146 241 -130
rect 275 -146 276 -130
rect 282 -197 283 -145
rect 506 -197 507 -145
rect 513 -146 514 -130
rect 520 -197 521 -145
rect 89 -197 90 -147
rect 198 -148 199 -130
rect 247 -148 248 -130
rect 275 -197 276 -147
rect 292 -197 293 -147
rect 457 -197 458 -147
rect 499 -148 500 -130
rect 632 -197 633 -147
rect 93 -150 94 -130
rect 478 -197 479 -149
rect 485 -150 486 -130
rect 499 -197 500 -149
rect 93 -197 94 -151
rect 271 -197 272 -151
rect 296 -197 297 -151
rect 324 -152 325 -130
rect 327 -152 328 -130
rect 604 -197 605 -151
rect 100 -154 101 -130
rect 562 -197 563 -153
rect 100 -197 101 -155
rect 149 -156 150 -130
rect 152 -197 153 -155
rect 534 -197 535 -155
rect 128 -197 129 -157
rect 219 -158 220 -130
rect 261 -158 262 -130
rect 415 -197 416 -157
rect 422 -197 423 -157
rect 471 -197 472 -157
rect 107 -160 108 -130
rect 261 -197 262 -159
rect 303 -160 304 -130
rect 359 -197 360 -159
rect 373 -197 374 -159
rect 450 -160 451 -130
rect 107 -197 108 -161
rect 159 -162 160 -130
rect 163 -162 164 -130
rect 163 -197 164 -161
rect 163 -162 164 -130
rect 163 -197 164 -161
rect 170 -162 171 -130
rect 548 -197 549 -161
rect 117 -197 118 -163
rect 219 -197 220 -163
rect 226 -164 227 -130
rect 303 -197 304 -163
rect 341 -197 342 -163
rect 597 -197 598 -163
rect 135 -166 136 -130
rect 611 -197 612 -165
rect 138 -168 139 -130
rect 142 -168 143 -130
rect 149 -197 150 -167
rect 464 -197 465 -167
rect 142 -197 143 -169
rect 289 -170 290 -130
rect 352 -170 353 -130
rect 492 -170 493 -130
rect 156 -197 157 -171
rect 187 -197 188 -171
rect 191 -172 192 -130
rect 352 -197 353 -171
rect 450 -197 451 -171
rect 170 -197 171 -173
rect 233 -174 234 -130
rect 289 -197 290 -173
rect 492 -197 493 -173
rect 177 -197 178 -175
rect 590 -197 591 -175
rect 180 -197 181 -177
rect 240 -197 241 -177
rect 387 -178 388 -130
rect 513 -197 514 -177
rect 191 -197 192 -179
rect 254 -197 255 -179
rect 324 -197 325 -179
rect 387 -197 388 -179
rect 394 -180 395 -130
rect 646 -197 647 -179
rect 198 -197 199 -181
rect 625 -197 626 -181
rect 205 -184 206 -130
rect 226 -197 227 -183
rect 317 -184 318 -130
rect 394 -197 395 -183
rect 408 -184 409 -130
rect 485 -197 486 -183
rect 135 -197 136 -185
rect 317 -197 318 -185
rect 408 -197 409 -185
rect 576 -197 577 -185
rect 212 -188 213 -130
rect 233 -197 234 -187
rect 429 -188 430 -130
rect 555 -197 556 -187
rect 366 -190 367 -130
rect 429 -197 430 -189
rect 436 -190 437 -130
rect 541 -197 542 -189
rect 86 -192 87 -130
rect 436 -197 437 -191
rect 345 -194 346 -130
rect 366 -197 367 -193
rect 310 -196 311 -130
rect 345 -197 346 -195
rect 16 -207 17 -205
rect 16 -270 17 -206
rect 16 -207 17 -205
rect 16 -270 17 -206
rect 30 -207 31 -205
rect 30 -270 31 -206
rect 30 -207 31 -205
rect 30 -270 31 -206
rect 33 -207 34 -205
rect 590 -207 591 -205
rect 597 -207 598 -205
rect 667 -270 668 -206
rect 51 -270 52 -208
rect 212 -209 213 -205
rect 215 -209 216 -205
rect 604 -209 605 -205
rect 65 -211 66 -205
rect 201 -211 202 -205
rect 205 -270 206 -210
rect 240 -211 241 -205
rect 243 -270 244 -210
rect 513 -211 514 -205
rect 520 -211 521 -205
rect 604 -270 605 -210
rect 79 -213 80 -205
rect 306 -270 307 -212
rect 310 -270 311 -212
rect 324 -213 325 -205
rect 338 -213 339 -205
rect 625 -213 626 -205
rect 44 -215 45 -205
rect 324 -270 325 -214
rect 366 -215 367 -205
rect 408 -270 409 -214
rect 411 -215 412 -205
rect 506 -215 507 -205
rect 513 -270 514 -214
rect 527 -215 528 -205
rect 590 -270 591 -214
rect 632 -215 633 -205
rect 89 -217 90 -205
rect 422 -270 423 -216
rect 464 -217 465 -205
rect 520 -270 521 -216
rect 527 -270 528 -216
rect 541 -217 542 -205
rect 597 -270 598 -216
rect 639 -217 640 -205
rect 100 -219 101 -205
rect 180 -219 181 -205
rect 187 -219 188 -205
rect 226 -219 227 -205
rect 254 -219 255 -205
rect 345 -219 346 -205
rect 373 -219 374 -205
rect 541 -270 542 -218
rect 625 -270 626 -218
rect 653 -219 654 -205
rect 103 -270 104 -220
rect 177 -270 178 -220
rect 198 -221 199 -205
rect 457 -221 458 -205
rect 464 -270 465 -220
rect 485 -221 486 -205
rect 492 -221 493 -205
rect 492 -270 493 -220
rect 492 -221 493 -205
rect 492 -270 493 -220
rect 632 -270 633 -220
rect 660 -221 661 -205
rect 72 -223 73 -205
rect 198 -270 199 -222
rect 208 -223 209 -205
rect 534 -223 535 -205
rect 72 -270 73 -224
rect 82 -270 83 -224
rect 114 -225 115 -205
rect 184 -270 185 -224
rect 219 -225 220 -205
rect 226 -270 227 -224
rect 247 -225 248 -205
rect 457 -270 458 -224
rect 478 -225 479 -205
rect 478 -270 479 -224
rect 478 -225 479 -205
rect 478 -270 479 -224
rect 485 -270 486 -224
rect 562 -225 563 -205
rect 58 -227 59 -205
rect 219 -270 220 -226
rect 257 -227 258 -205
rect 359 -227 360 -205
rect 373 -270 374 -226
rect 401 -227 402 -205
rect 499 -227 500 -205
rect 562 -270 563 -226
rect 58 -270 59 -228
rect 506 -270 507 -228
rect 534 -270 535 -228
rect 555 -229 556 -205
rect 114 -270 115 -230
rect 191 -231 192 -205
rect 257 -270 258 -230
rect 576 -231 577 -205
rect 121 -233 122 -205
rect 345 -270 346 -232
rect 359 -270 360 -232
rect 380 -233 381 -205
rect 387 -233 388 -205
rect 583 -233 584 -205
rect 121 -270 122 -234
rect 583 -270 584 -234
rect 124 -270 125 -236
rect 303 -237 304 -205
rect 313 -237 314 -205
rect 548 -237 549 -205
rect 65 -270 66 -238
rect 303 -270 304 -238
rect 317 -239 318 -205
rect 401 -270 402 -238
rect 548 -270 549 -238
rect 618 -239 619 -205
rect 128 -241 129 -205
rect 380 -270 381 -240
rect 387 -270 388 -240
rect 429 -241 430 -205
rect 576 -270 577 -240
rect 618 -270 619 -240
rect 128 -270 129 -242
rect 240 -270 241 -242
rect 268 -243 269 -205
rect 611 -243 612 -205
rect 135 -245 136 -205
rect 352 -245 353 -205
rect 429 -270 430 -244
rect 471 -245 472 -205
rect 100 -270 101 -246
rect 135 -270 136 -246
rect 142 -247 143 -205
rect 163 -247 164 -205
rect 170 -247 171 -205
rect 212 -270 213 -246
rect 268 -270 269 -246
rect 499 -270 500 -246
rect 93 -249 94 -205
rect 170 -270 171 -248
rect 191 -270 192 -248
rect 250 -249 251 -205
rect 275 -249 276 -205
rect 289 -270 290 -248
rect 292 -249 293 -205
rect 394 -249 395 -205
rect 443 -249 444 -205
rect 471 -270 472 -248
rect 89 -270 90 -250
rect 394 -270 395 -250
rect 436 -251 437 -205
rect 443 -270 444 -250
rect 93 -270 94 -252
rect 296 -253 297 -205
rect 299 -270 300 -252
rect 331 -253 332 -205
rect 334 -270 335 -252
rect 611 -270 612 -252
rect 107 -255 108 -205
rect 163 -270 164 -254
rect 282 -255 283 -205
rect 569 -255 570 -205
rect 107 -270 108 -256
rect 156 -257 157 -205
rect 180 -270 181 -256
rect 569 -270 570 -256
rect 142 -270 143 -258
rect 156 -270 157 -258
rect 320 -270 321 -258
rect 450 -259 451 -205
rect 149 -270 150 -260
rect 233 -261 234 -205
rect 285 -261 286 -205
rect 450 -270 451 -260
rect 23 -263 24 -205
rect 233 -270 234 -262
rect 285 -270 286 -262
rect 415 -263 416 -205
rect 425 -263 426 -205
rect 436 -270 437 -262
rect 152 -265 153 -205
rect 261 -265 262 -205
rect 282 -270 283 -264
rect 415 -270 416 -264
rect 261 -270 262 -266
rect 278 -270 279 -266
rect 331 -270 332 -266
rect 646 -267 647 -205
rect 338 -270 339 -268
rect 366 -270 367 -268
rect 44 -280 45 -278
rect 47 -335 48 -279
rect 58 -280 59 -278
rect 212 -280 213 -278
rect 219 -280 220 -278
rect 219 -335 220 -279
rect 219 -280 220 -278
rect 219 -335 220 -279
rect 226 -280 227 -278
rect 226 -335 227 -279
rect 226 -280 227 -278
rect 226 -335 227 -279
rect 247 -335 248 -279
rect 345 -280 346 -278
rect 355 -280 356 -278
rect 387 -280 388 -278
rect 390 -335 391 -279
rect 478 -280 479 -278
rect 506 -280 507 -278
rect 618 -335 619 -279
rect 667 -280 668 -278
rect 709 -335 710 -279
rect 58 -335 59 -281
rect 254 -282 255 -278
rect 261 -282 262 -278
rect 275 -335 276 -281
rect 282 -282 283 -278
rect 310 -282 311 -278
rect 317 -282 318 -278
rect 660 -335 661 -281
rect 72 -284 73 -278
rect 177 -284 178 -278
rect 187 -335 188 -283
rect 261 -335 262 -283
rect 282 -335 283 -283
rect 338 -284 339 -278
rect 341 -335 342 -283
rect 520 -284 521 -278
rect 555 -335 556 -283
rect 639 -284 640 -278
rect 72 -335 73 -285
rect 569 -286 570 -278
rect 583 -286 584 -278
rect 639 -335 640 -285
rect 89 -288 90 -278
rect 478 -335 479 -287
rect 513 -288 514 -278
rect 674 -335 675 -287
rect 89 -335 90 -289
rect 485 -290 486 -278
rect 527 -290 528 -278
rect 569 -335 570 -289
rect 590 -290 591 -278
rect 646 -335 647 -289
rect 100 -292 101 -278
rect 653 -335 654 -291
rect 107 -294 108 -278
rect 212 -335 213 -293
rect 285 -294 286 -278
rect 485 -335 486 -293
rect 492 -294 493 -278
rect 527 -335 528 -293
rect 534 -294 535 -278
rect 583 -335 584 -293
rect 604 -294 605 -278
rect 667 -335 668 -293
rect 16 -335 17 -295
rect 604 -335 605 -295
rect 107 -335 108 -297
rect 128 -298 129 -278
rect 145 -335 146 -297
rect 159 -298 160 -278
rect 163 -298 164 -278
rect 254 -335 255 -297
rect 289 -298 290 -278
rect 289 -335 290 -297
rect 289 -298 290 -278
rect 289 -335 290 -297
rect 296 -298 297 -278
rect 625 -298 626 -278
rect 54 -335 55 -299
rect 625 -335 626 -299
rect 65 -302 66 -278
rect 296 -335 297 -301
rect 299 -302 300 -278
rect 331 -335 332 -301
rect 362 -335 363 -301
rect 513 -335 514 -301
rect 541 -302 542 -278
rect 590 -335 591 -301
rect 114 -304 115 -278
rect 128 -335 129 -303
rect 149 -304 150 -278
rect 268 -304 269 -278
rect 306 -304 307 -278
rect 632 -304 633 -278
rect 114 -335 115 -305
rect 250 -306 251 -278
rect 320 -306 321 -278
rect 429 -306 430 -278
rect 450 -306 451 -278
rect 506 -335 507 -305
rect 541 -335 542 -305
rect 562 -306 563 -278
rect 30 -308 31 -278
rect 429 -335 430 -307
rect 436 -308 437 -278
rect 450 -335 451 -307
rect 464 -308 465 -278
rect 520 -335 521 -307
rect 562 -335 563 -307
rect 611 -308 612 -278
rect 30 -335 31 -309
rect 82 -335 83 -309
rect 121 -310 122 -278
rect 387 -335 388 -309
rect 401 -310 402 -278
rect 401 -335 402 -309
rect 401 -310 402 -278
rect 401 -335 402 -309
rect 415 -310 416 -278
rect 436 -335 437 -309
rect 443 -310 444 -278
rect 464 -335 465 -309
rect 499 -310 500 -278
rect 534 -335 535 -309
rect 576 -310 577 -278
rect 611 -335 612 -309
rect 23 -335 24 -311
rect 121 -335 122 -311
rect 142 -312 143 -278
rect 268 -335 269 -311
rect 320 -335 321 -311
rect 632 -335 633 -311
rect 159 -335 160 -313
rect 380 -314 381 -278
rect 408 -314 409 -278
rect 443 -335 444 -313
rect 471 -314 472 -278
rect 576 -335 577 -313
rect 65 -335 66 -315
rect 408 -335 409 -315
rect 415 -335 416 -315
rect 422 -316 423 -278
rect 457 -316 458 -278
rect 471 -335 472 -315
rect 79 -318 80 -278
rect 457 -335 458 -317
rect 51 -320 52 -278
rect 79 -335 80 -319
rect 142 -335 143 -319
rect 380 -335 381 -319
rect 394 -320 395 -278
rect 422 -335 423 -319
rect 37 -335 38 -321
rect 51 -335 52 -321
rect 170 -322 171 -278
rect 177 -335 178 -321
rect 191 -322 192 -278
rect 334 -322 335 -278
rect 352 -322 353 -278
rect 394 -335 395 -321
rect 135 -324 136 -278
rect 170 -335 171 -323
rect 191 -335 192 -323
rect 198 -324 199 -278
rect 201 -335 202 -323
rect 303 -324 304 -278
rect 324 -324 325 -278
rect 345 -335 346 -323
rect 366 -335 367 -323
rect 373 -324 374 -278
rect 135 -335 136 -325
rect 233 -326 234 -278
rect 313 -335 314 -325
rect 373 -335 374 -325
rect 184 -328 185 -278
rect 303 -335 304 -327
rect 324 -335 325 -327
rect 499 -335 500 -327
rect 149 -335 150 -329
rect 184 -335 185 -329
rect 205 -330 206 -278
rect 317 -335 318 -329
rect 369 -330 370 -278
rect 548 -330 549 -278
rect 93 -332 94 -278
rect 205 -335 206 -331
rect 233 -335 234 -331
rect 359 -332 360 -278
rect 548 -335 549 -331
rect 597 -332 598 -278
rect 93 -335 94 -333
rect 240 -335 241 -333
rect 9 -345 10 -343
rect 660 -345 661 -343
rect 709 -345 710 -343
rect 716 -402 717 -344
rect 12 -347 13 -343
rect 65 -402 66 -346
rect 68 -347 69 -343
rect 618 -347 619 -343
rect 23 -402 24 -348
rect 128 -349 129 -343
rect 142 -349 143 -343
rect 303 -349 304 -343
rect 313 -349 314 -343
rect 366 -349 367 -343
rect 436 -349 437 -343
rect 436 -402 437 -348
rect 436 -349 437 -343
rect 436 -402 437 -348
rect 467 -402 468 -348
rect 625 -349 626 -343
rect 30 -402 31 -350
rect 79 -351 80 -343
rect 89 -351 90 -343
rect 506 -351 507 -343
rect 548 -351 549 -343
rect 618 -402 619 -350
rect 37 -353 38 -343
rect 44 -353 45 -343
rect 51 -402 52 -352
rect 481 -402 482 -352
rect 506 -402 507 -352
rect 534 -353 535 -343
rect 555 -353 556 -343
rect 555 -402 556 -352
rect 555 -353 556 -343
rect 555 -402 556 -352
rect 597 -402 598 -352
rect 632 -353 633 -343
rect 37 -402 38 -354
rect 464 -355 465 -343
rect 471 -355 472 -343
rect 660 -402 661 -354
rect 44 -402 45 -356
rect 331 -357 332 -343
rect 338 -402 339 -356
rect 443 -357 444 -343
rect 450 -357 451 -343
rect 471 -402 472 -356
rect 72 -402 73 -358
rect 100 -359 101 -343
rect 117 -402 118 -358
rect 191 -359 192 -343
rect 198 -402 199 -358
rect 247 -359 248 -343
rect 275 -359 276 -343
rect 275 -402 276 -358
rect 275 -359 276 -343
rect 275 -402 276 -358
rect 282 -359 283 -343
rect 362 -359 363 -343
rect 390 -359 391 -343
rect 534 -402 535 -358
rect 75 -361 76 -343
rect 408 -361 409 -343
rect 411 -402 412 -360
rect 625 -402 626 -360
rect 79 -402 80 -362
rect 156 -363 157 -343
rect 163 -363 164 -343
rect 212 -363 213 -343
rect 226 -363 227 -343
rect 327 -363 328 -343
rect 355 -363 356 -343
rect 653 -363 654 -343
rect 86 -365 87 -343
rect 100 -402 101 -364
rect 107 -365 108 -343
rect 163 -402 164 -364
rect 177 -365 178 -343
rect 212 -402 213 -364
rect 219 -365 220 -343
rect 226 -402 227 -364
rect 233 -365 234 -343
rect 366 -402 367 -364
rect 390 -402 391 -364
rect 415 -365 416 -343
rect 443 -402 444 -364
rect 485 -365 486 -343
rect 590 -365 591 -343
rect 653 -402 654 -364
rect 86 -402 87 -366
rect 93 -367 94 -343
rect 110 -402 111 -366
rect 219 -402 220 -366
rect 233 -402 234 -366
rect 268 -367 269 -343
rect 282 -402 283 -366
rect 341 -367 342 -343
rect 359 -367 360 -343
rect 583 -367 584 -343
rect 590 -402 591 -366
rect 611 -367 612 -343
rect 58 -369 59 -343
rect 359 -402 360 -368
rect 394 -369 395 -343
rect 415 -402 416 -368
rect 450 -402 451 -368
rect 478 -369 479 -343
rect 485 -402 486 -368
rect 513 -369 514 -343
rect 583 -402 584 -368
rect 635 -402 636 -368
rect 58 -402 59 -370
rect 156 -402 157 -370
rect 201 -371 202 -343
rect 205 -371 206 -343
rect 247 -402 248 -370
rect 254 -371 255 -343
rect 268 -402 269 -370
rect 310 -371 311 -343
rect 317 -402 318 -370
rect 380 -371 381 -343
rect 457 -371 458 -343
rect 548 -402 549 -370
rect 121 -373 122 -343
rect 191 -402 192 -372
rect 254 -402 255 -372
rect 383 -402 384 -372
rect 457 -402 458 -372
rect 520 -373 521 -343
rect 121 -402 122 -374
rect 422 -375 423 -343
rect 492 -375 493 -343
rect 513 -402 514 -374
rect 128 -402 129 -376
rect 170 -377 171 -343
rect 187 -402 188 -376
rect 205 -402 206 -376
rect 296 -377 297 -343
rect 310 -402 311 -376
rect 324 -377 325 -343
rect 674 -377 675 -343
rect 114 -379 115 -343
rect 296 -402 297 -378
rect 303 -402 304 -378
rect 345 -379 346 -343
rect 352 -379 353 -343
rect 520 -402 521 -378
rect 135 -381 136 -343
rect 177 -402 178 -380
rect 334 -402 335 -380
rect 394 -402 395 -380
rect 422 -402 423 -380
rect 527 -381 528 -343
rect 135 -402 136 -382
rect 289 -383 290 -343
rect 345 -402 346 -382
rect 373 -383 374 -343
rect 380 -402 381 -382
rect 646 -383 647 -343
rect 142 -402 143 -384
rect 149 -385 150 -343
rect 170 -402 171 -384
rect 261 -385 262 -343
rect 289 -402 290 -384
rect 429 -385 430 -343
rect 492 -402 493 -384
rect 639 -385 640 -343
rect 93 -402 94 -386
rect 149 -402 150 -386
rect 261 -402 262 -386
rect 387 -402 388 -386
rect 495 -387 496 -343
rect 527 -402 528 -386
rect 562 -387 563 -343
rect 646 -402 647 -386
rect 355 -402 356 -388
rect 611 -402 612 -388
rect 373 -402 374 -390
rect 576 -391 577 -343
rect 604 -391 605 -343
rect 639 -402 640 -390
rect 541 -393 542 -343
rect 576 -402 577 -392
rect 604 -402 605 -392
rect 667 -393 668 -343
rect 243 -402 244 -394
rect 541 -402 542 -394
rect 562 -402 563 -394
rect 569 -395 570 -343
rect 324 -402 325 -396
rect 569 -402 570 -396
rect 401 -399 402 -343
rect 667 -402 668 -398
rect 401 -402 402 -400
rect 499 -401 500 -343
rect 9 -467 10 -411
rect 96 -412 97 -410
rect 100 -412 101 -410
rect 194 -467 195 -411
rect 198 -412 199 -410
rect 243 -412 244 -410
rect 268 -412 269 -410
rect 373 -412 374 -410
rect 383 -412 384 -410
rect 527 -412 528 -410
rect 562 -412 563 -410
rect 653 -467 654 -411
rect 656 -412 657 -410
rect 660 -412 661 -410
rect 716 -412 717 -410
rect 730 -467 731 -411
rect 16 -467 17 -413
rect 79 -414 80 -410
rect 93 -414 94 -410
rect 422 -414 423 -410
rect 425 -467 426 -413
rect 576 -414 577 -410
rect 597 -414 598 -410
rect 681 -467 682 -413
rect 23 -416 24 -410
rect 82 -467 83 -415
rect 114 -467 115 -415
rect 170 -416 171 -410
rect 180 -467 181 -415
rect 639 -416 640 -410
rect 30 -467 31 -417
rect 103 -467 104 -417
rect 121 -418 122 -410
rect 576 -467 577 -417
rect 583 -418 584 -410
rect 639 -467 640 -417
rect 37 -420 38 -410
rect 110 -420 111 -410
rect 156 -467 157 -419
rect 240 -420 241 -410
rect 247 -420 248 -410
rect 268 -467 269 -419
rect 275 -420 276 -410
rect 275 -467 276 -419
rect 275 -420 276 -410
rect 275 -467 276 -419
rect 282 -420 283 -410
rect 520 -420 521 -410
rect 534 -420 535 -410
rect 562 -467 563 -419
rect 569 -420 570 -410
rect 723 -467 724 -419
rect 37 -467 38 -421
rect 51 -422 52 -410
rect 58 -422 59 -410
rect 352 -422 353 -410
rect 373 -467 374 -421
rect 422 -467 423 -421
rect 432 -422 433 -410
rect 499 -467 500 -421
rect 513 -422 514 -410
rect 569 -467 570 -421
rect 604 -422 605 -410
rect 702 -467 703 -421
rect 44 -424 45 -410
rect 93 -467 94 -423
rect 100 -467 101 -423
rect 121 -467 122 -423
rect 135 -424 136 -410
rect 240 -467 241 -423
rect 303 -424 304 -410
rect 352 -467 353 -423
rect 387 -424 388 -410
rect 453 -467 454 -423
rect 464 -424 465 -410
rect 597 -467 598 -423
rect 611 -424 612 -410
rect 688 -467 689 -423
rect 44 -467 45 -425
rect 142 -426 143 -410
rect 163 -426 164 -410
rect 338 -467 339 -425
rect 390 -426 391 -410
rect 618 -426 619 -410
rect 625 -426 626 -410
rect 674 -467 675 -425
rect 58 -467 59 -427
rect 128 -428 129 -410
rect 135 -467 136 -427
rect 205 -428 206 -410
rect 219 -428 220 -410
rect 226 -467 227 -427
rect 233 -428 234 -410
rect 282 -467 283 -427
rect 296 -428 297 -410
rect 387 -467 388 -427
rect 390 -467 391 -427
rect 527 -467 528 -427
rect 541 -428 542 -410
rect 583 -467 584 -427
rect 65 -467 66 -429
rect 107 -467 108 -429
rect 149 -430 150 -410
rect 205 -467 206 -429
rect 212 -430 213 -410
rect 233 -467 234 -429
rect 313 -467 314 -429
rect 464 -467 465 -429
rect 481 -430 482 -410
rect 632 -467 633 -429
rect 68 -432 69 -410
rect 541 -467 542 -431
rect 555 -432 556 -410
rect 604 -467 605 -431
rect 72 -434 73 -410
rect 124 -434 125 -410
rect 149 -467 150 -433
rect 285 -434 286 -410
rect 324 -467 325 -433
rect 359 -434 360 -410
rect 401 -434 402 -410
rect 534 -467 535 -433
rect 72 -467 73 -435
rect 380 -436 381 -410
rect 408 -467 409 -435
rect 646 -436 647 -410
rect 86 -438 87 -410
rect 247 -467 248 -437
rect 327 -438 328 -410
rect 548 -438 549 -410
rect 590 -438 591 -410
rect 646 -467 647 -437
rect 86 -467 87 -439
rect 254 -440 255 -410
rect 331 -467 332 -439
rect 446 -467 447 -439
rect 450 -440 451 -410
rect 513 -467 514 -439
rect 170 -467 171 -441
rect 303 -467 304 -441
rect 345 -442 346 -410
rect 380 -467 381 -441
rect 411 -467 412 -441
rect 590 -467 591 -441
rect 177 -444 178 -410
rect 212 -467 213 -443
rect 254 -467 255 -443
rect 317 -444 318 -410
rect 359 -467 360 -443
rect 418 -467 419 -443
rect 436 -444 437 -410
rect 548 -467 549 -443
rect 128 -467 129 -445
rect 177 -467 178 -445
rect 184 -446 185 -410
rect 289 -446 290 -410
rect 310 -446 311 -410
rect 345 -467 346 -445
rect 366 -446 367 -410
rect 401 -467 402 -445
rect 436 -467 437 -445
rect 625 -467 626 -445
rect 184 -467 185 -447
rect 219 -467 220 -447
rect 229 -448 230 -410
rect 317 -467 318 -447
rect 439 -467 440 -447
rect 709 -467 710 -447
rect 191 -450 192 -410
rect 296 -467 297 -449
rect 443 -450 444 -410
rect 520 -467 521 -449
rect 51 -467 52 -451
rect 191 -467 192 -451
rect 198 -467 199 -451
rect 261 -452 262 -410
rect 289 -467 290 -451
rect 394 -452 395 -410
rect 492 -452 493 -410
rect 695 -467 696 -451
rect 166 -467 167 -453
rect 261 -467 262 -453
rect 394 -467 395 -453
rect 457 -454 458 -410
rect 485 -454 486 -410
rect 492 -467 493 -453
rect 502 -454 503 -410
rect 611 -467 612 -453
rect 341 -456 342 -410
rect 457 -467 458 -455
rect 506 -456 507 -410
rect 555 -467 556 -455
rect 366 -467 367 -457
rect 485 -467 486 -457
rect 471 -460 472 -410
rect 506 -467 507 -459
rect 471 -467 472 -461
rect 667 -462 668 -410
rect 478 -464 479 -410
rect 667 -467 668 -463
rect 415 -466 416 -410
rect 478 -467 479 -465
rect 58 -477 59 -475
rect 163 -477 164 -475
rect 177 -477 178 -475
rect 604 -477 605 -475
rect 639 -477 640 -475
rect 709 -552 710 -476
rect 716 -477 717 -475
rect 730 -477 731 -475
rect 75 -479 76 -475
rect 744 -552 745 -478
rect 23 -552 24 -480
rect 75 -552 76 -480
rect 79 -481 80 -475
rect 737 -552 738 -480
rect 79 -552 80 -482
rect 135 -483 136 -475
rect 145 -483 146 -475
rect 695 -483 696 -475
rect 723 -483 724 -475
rect 779 -552 780 -482
rect 93 -485 94 -475
rect 145 -552 146 -484
rect 152 -552 153 -484
rect 205 -485 206 -475
rect 219 -485 220 -475
rect 222 -501 223 -484
rect 243 -552 244 -484
rect 345 -485 346 -475
rect 359 -485 360 -475
rect 618 -552 619 -484
rect 646 -485 647 -475
rect 723 -552 724 -484
rect 37 -487 38 -475
rect 93 -552 94 -486
rect 121 -487 122 -475
rect 191 -487 192 -475
rect 198 -487 199 -475
rect 198 -552 199 -486
rect 198 -487 199 -475
rect 198 -552 199 -486
rect 219 -552 220 -486
rect 254 -487 255 -475
rect 275 -487 276 -475
rect 275 -552 276 -486
rect 275 -487 276 -475
rect 275 -552 276 -486
rect 289 -487 290 -475
rect 450 -552 451 -486
rect 555 -487 556 -475
rect 604 -552 605 -486
rect 674 -487 675 -475
rect 716 -552 717 -486
rect 121 -552 122 -488
rect 268 -489 269 -475
rect 289 -552 290 -488
rect 331 -489 332 -475
rect 345 -552 346 -488
rect 373 -489 374 -475
rect 383 -489 384 -475
rect 415 -552 416 -488
rect 422 -552 423 -488
rect 639 -552 640 -488
rect 51 -491 52 -475
rect 331 -552 332 -490
rect 352 -491 353 -475
rect 359 -552 360 -490
rect 366 -491 367 -475
rect 548 -491 549 -475
rect 555 -552 556 -490
rect 590 -491 591 -475
rect 597 -491 598 -475
rect 660 -552 661 -490
rect 16 -493 17 -475
rect 590 -552 591 -492
rect 30 -495 31 -475
rect 51 -552 52 -494
rect 124 -552 125 -494
rect 695 -552 696 -494
rect 128 -497 129 -475
rect 268 -552 269 -496
rect 390 -497 391 -475
rect 611 -497 612 -475
rect 107 -499 108 -475
rect 128 -552 129 -498
rect 135 -552 136 -498
rect 719 -499 720 -475
rect 44 -501 45 -475
rect 107 -552 108 -500
rect 149 -501 150 -475
rect 205 -552 206 -500
rect 254 -552 255 -500
rect 394 -501 395 -475
rect 751 -552 752 -500
rect 44 -552 45 -502
rect 114 -503 115 -475
rect 156 -503 157 -475
rect 156 -552 157 -502
rect 156 -503 157 -475
rect 156 -552 157 -502
rect 180 -503 181 -475
rect 212 -503 213 -475
rect 247 -503 248 -475
rect 247 -552 248 -502
rect 247 -503 248 -475
rect 247 -552 248 -502
rect 408 -503 409 -475
rect 436 -552 437 -502
rect 439 -503 440 -475
rect 681 -503 682 -475
rect 61 -552 62 -504
rect 114 -552 115 -504
rect 187 -505 188 -475
rect 338 -505 339 -475
rect 401 -505 402 -475
rect 408 -552 409 -504
rect 411 -505 412 -475
rect 478 -505 479 -475
rect 513 -505 514 -475
rect 548 -552 549 -504
rect 562 -505 563 -475
rect 611 -552 612 -504
rect 625 -505 626 -475
rect 681 -552 682 -504
rect 65 -552 66 -506
rect 625 -552 626 -506
rect 170 -509 171 -475
rect 562 -552 563 -508
rect 576 -509 577 -475
rect 646 -552 647 -508
rect 170 -552 171 -510
rect 282 -511 283 -475
rect 303 -511 304 -475
rect 338 -552 339 -510
rect 429 -511 430 -475
rect 653 -511 654 -475
rect 191 -552 192 -512
rect 310 -513 311 -475
rect 324 -513 325 -475
rect 401 -552 402 -512
rect 432 -513 433 -475
rect 597 -552 598 -512
rect 142 -515 143 -475
rect 310 -552 311 -514
rect 317 -515 318 -475
rect 324 -552 325 -514
rect 432 -552 433 -514
rect 667 -515 668 -475
rect 212 -552 213 -516
rect 296 -517 297 -475
rect 303 -552 304 -516
rect 730 -552 731 -516
rect 226 -519 227 -475
rect 317 -552 318 -518
rect 397 -552 398 -518
rect 667 -552 668 -518
rect 226 -552 227 -520
rect 233 -521 234 -475
rect 240 -521 241 -475
rect 296 -552 297 -520
rect 443 -521 444 -475
rect 702 -521 703 -475
rect 233 -552 234 -522
rect 352 -552 353 -522
rect 387 -523 388 -475
rect 702 -552 703 -522
rect 240 -552 241 -524
rect 373 -552 374 -524
rect 443 -552 444 -524
rect 688 -525 689 -475
rect 261 -527 262 -475
rect 387 -552 388 -526
rect 478 -552 479 -526
rect 527 -527 528 -475
rect 534 -527 535 -475
rect 576 -552 577 -526
rect 583 -527 584 -475
rect 653 -552 654 -526
rect 282 -552 283 -528
rect 369 -552 370 -528
rect 453 -529 454 -475
rect 534 -552 535 -528
rect 632 -529 633 -475
rect 688 -552 689 -528
rect 9 -531 10 -475
rect 632 -552 633 -530
rect 492 -533 493 -475
rect 583 -552 584 -532
rect 446 -535 447 -475
rect 492 -552 493 -534
rect 506 -535 507 -475
rect 527 -552 528 -534
rect 261 -552 262 -536
rect 446 -552 447 -536
rect 513 -552 514 -536
rect 541 -537 542 -475
rect 320 -552 321 -538
rect 506 -552 507 -538
rect 520 -539 521 -475
rect 674 -552 675 -538
rect 499 -541 500 -475
rect 520 -552 521 -540
rect 541 -552 542 -540
rect 569 -541 570 -475
rect 464 -543 465 -475
rect 569 -552 570 -542
rect 457 -545 458 -475
rect 464 -552 465 -544
rect 485 -545 486 -475
rect 499 -552 500 -544
rect 86 -547 87 -475
rect 457 -552 458 -546
rect 471 -547 472 -475
rect 485 -552 486 -546
rect 68 -549 69 -475
rect 471 -552 472 -548
rect 26 -551 27 -475
rect 68 -552 69 -550
rect 86 -552 87 -550
rect 163 -552 164 -550
rect 16 -645 17 -561
rect 408 -562 409 -560
rect 418 -645 419 -561
rect 723 -562 724 -560
rect 779 -562 780 -560
rect 807 -645 808 -561
rect 23 -564 24 -560
rect 54 -564 55 -560
rect 58 -645 59 -563
rect 135 -564 136 -560
rect 156 -564 157 -560
rect 177 -564 178 -560
rect 187 -564 188 -560
rect 282 -564 283 -560
rect 306 -564 307 -560
rect 324 -564 325 -560
rect 355 -645 356 -563
rect 520 -564 521 -560
rect 541 -564 542 -560
rect 544 -578 545 -563
rect 562 -564 563 -560
rect 562 -645 563 -563
rect 562 -564 563 -560
rect 562 -645 563 -563
rect 23 -645 24 -565
rect 124 -645 125 -565
rect 128 -566 129 -560
rect 156 -645 157 -565
rect 166 -566 167 -560
rect 674 -566 675 -560
rect 30 -645 31 -567
rect 96 -645 97 -567
rect 100 -645 101 -567
rect 149 -645 150 -567
rect 177 -645 178 -567
rect 187 -645 188 -567
rect 205 -568 206 -560
rect 215 -568 216 -560
rect 219 -568 220 -560
rect 317 -568 318 -560
rect 366 -568 367 -560
rect 499 -568 500 -560
rect 541 -645 542 -567
rect 576 -568 577 -560
rect 33 -645 34 -569
rect 51 -570 52 -560
rect 61 -570 62 -560
rect 625 -570 626 -560
rect 40 -572 41 -560
rect 40 -645 41 -571
rect 40 -572 41 -560
rect 40 -645 41 -571
rect 44 -572 45 -560
rect 128 -645 129 -571
rect 191 -572 192 -560
rect 317 -645 318 -571
rect 369 -572 370 -560
rect 674 -645 675 -571
rect 47 -645 48 -573
rect 653 -574 654 -560
rect 51 -645 52 -575
rect 366 -645 367 -575
rect 394 -576 395 -560
rect 646 -576 647 -560
rect 65 -578 66 -560
rect 397 -578 398 -560
rect 411 -645 412 -577
rect 499 -645 500 -577
rect 576 -645 577 -577
rect 625 -645 626 -577
rect 688 -578 689 -560
rect 65 -645 66 -579
rect 352 -580 353 -560
rect 394 -645 395 -579
rect 751 -580 752 -560
rect 72 -582 73 -560
rect 590 -582 591 -560
rect 646 -645 647 -581
rect 695 -582 696 -560
rect 72 -645 73 -583
rect 142 -584 143 -560
rect 191 -645 192 -583
rect 198 -584 199 -560
rect 212 -584 213 -560
rect 723 -645 724 -583
rect 107 -586 108 -560
rect 184 -586 185 -560
rect 212 -645 213 -585
rect 401 -586 402 -560
rect 425 -586 426 -560
rect 534 -586 535 -560
rect 590 -645 591 -585
rect 639 -586 640 -560
rect 688 -645 689 -585
rect 730 -586 731 -560
rect 114 -588 115 -560
rect 135 -645 136 -587
rect 219 -645 220 -587
rect 310 -588 311 -560
rect 338 -588 339 -560
rect 369 -645 370 -587
rect 401 -645 402 -587
rect 415 -588 416 -560
rect 429 -588 430 -560
rect 569 -588 570 -560
rect 597 -588 598 -560
rect 695 -645 696 -587
rect 730 -645 731 -587
rect 737 -588 738 -560
rect 226 -590 227 -560
rect 520 -645 521 -589
rect 569 -645 570 -589
rect 604 -590 605 -560
rect 226 -645 227 -591
rect 261 -592 262 -560
rect 275 -592 276 -560
rect 278 -645 279 -591
rect 282 -645 283 -591
rect 296 -592 297 -560
rect 310 -645 311 -591
rect 450 -592 451 -560
rect 471 -592 472 -560
rect 737 -645 738 -591
rect 233 -594 234 -560
rect 296 -645 297 -593
rect 331 -594 332 -560
rect 415 -645 416 -593
rect 429 -645 430 -593
rect 464 -594 465 -560
rect 471 -645 472 -593
rect 492 -594 493 -560
rect 604 -645 605 -593
rect 660 -594 661 -560
rect 163 -596 164 -560
rect 660 -645 661 -595
rect 233 -645 234 -597
rect 254 -598 255 -560
rect 261 -645 262 -597
rect 387 -598 388 -560
rect 432 -598 433 -560
rect 709 -598 710 -560
rect 142 -645 143 -599
rect 709 -645 710 -599
rect 184 -645 185 -601
rect 254 -645 255 -601
rect 275 -645 276 -601
rect 653 -645 654 -601
rect 236 -604 237 -560
rect 744 -604 745 -560
rect 240 -606 241 -560
rect 247 -606 248 -560
rect 289 -606 290 -560
rect 324 -645 325 -605
rect 331 -645 332 -605
rect 373 -606 374 -560
rect 387 -645 388 -605
rect 667 -606 668 -560
rect 79 -608 80 -560
rect 240 -645 241 -607
rect 247 -645 248 -607
rect 268 -608 269 -560
rect 303 -608 304 -560
rect 373 -645 374 -607
rect 390 -645 391 -607
rect 667 -645 668 -607
rect 79 -645 80 -609
rect 170 -610 171 -560
rect 198 -645 199 -609
rect 289 -645 290 -609
rect 303 -645 304 -609
rect 345 -610 346 -560
rect 348 -645 349 -609
rect 597 -645 598 -609
rect 86 -612 87 -560
rect 170 -645 171 -611
rect 268 -645 269 -611
rect 292 -645 293 -611
rect 338 -645 339 -611
rect 457 -612 458 -560
rect 464 -645 465 -611
rect 555 -612 556 -560
rect 86 -645 87 -613
rect 103 -614 104 -560
rect 320 -614 321 -560
rect 457 -645 458 -613
rect 478 -614 479 -560
rect 534 -645 535 -613
rect 555 -645 556 -613
rect 716 -614 717 -560
rect 93 -616 94 -560
rect 345 -645 346 -615
rect 352 -645 353 -615
rect 618 -616 619 -560
rect 93 -645 94 -617
rect 205 -645 206 -617
rect 383 -618 384 -560
rect 618 -645 619 -617
rect 443 -645 444 -619
rect 611 -620 612 -560
rect 446 -622 447 -560
rect 702 -622 703 -560
rect 446 -645 447 -623
rect 639 -645 640 -623
rect 450 -645 451 -625
rect 548 -626 549 -560
rect 485 -628 486 -560
rect 611 -645 612 -627
rect 485 -645 486 -629
rect 506 -630 507 -560
rect 513 -630 514 -560
rect 702 -645 703 -629
rect 478 -645 479 -631
rect 513 -645 514 -631
rect 516 -645 517 -631
rect 716 -645 717 -631
rect 506 -645 507 -633
rect 527 -634 528 -560
rect 548 -645 549 -633
rect 583 -634 584 -560
rect 380 -636 381 -560
rect 527 -645 528 -635
rect 583 -645 584 -635
rect 632 -636 633 -560
rect 359 -638 360 -560
rect 380 -645 381 -637
rect 632 -645 633 -637
rect 681 -638 682 -560
rect 359 -645 360 -639
rect 436 -640 437 -560
rect 75 -642 76 -560
rect 436 -645 437 -641
rect 425 -645 426 -643
rect 681 -645 682 -643
rect 58 -655 59 -653
rect 96 -726 97 -654
rect 100 -655 101 -653
rect 114 -655 115 -653
rect 117 -655 118 -653
rect 156 -655 157 -653
rect 166 -655 167 -653
rect 177 -655 178 -653
rect 184 -655 185 -653
rect 240 -655 241 -653
rect 254 -655 255 -653
rect 345 -726 346 -654
rect 348 -655 349 -653
rect 450 -655 451 -653
rect 474 -726 475 -654
rect 765 -726 766 -654
rect 807 -655 808 -653
rect 828 -726 829 -654
rect 9 -726 10 -656
rect 114 -726 115 -656
rect 117 -726 118 -656
rect 198 -657 199 -653
rect 212 -657 213 -653
rect 254 -726 255 -656
rect 261 -657 262 -653
rect 278 -657 279 -653
rect 282 -657 283 -653
rect 289 -657 290 -653
rect 352 -657 353 -653
rect 415 -726 416 -656
rect 418 -657 419 -653
rect 513 -726 514 -656
rect 555 -657 556 -653
rect 772 -726 773 -656
rect 16 -659 17 -653
rect 352 -726 353 -658
rect 366 -659 367 -653
rect 534 -659 535 -653
rect 597 -659 598 -653
rect 824 -726 825 -658
rect 16 -726 17 -660
rect 72 -661 73 -653
rect 86 -661 87 -653
rect 121 -661 122 -653
rect 124 -661 125 -653
rect 432 -726 433 -660
rect 443 -661 444 -653
rect 555 -726 556 -660
rect 660 -726 661 -660
rect 695 -661 696 -653
rect 709 -661 710 -653
rect 786 -726 787 -660
rect 51 -663 52 -653
rect 100 -726 101 -662
rect 107 -663 108 -653
rect 583 -663 584 -653
rect 646 -663 647 -653
rect 695 -726 696 -662
rect 716 -663 717 -653
rect 793 -726 794 -662
rect 58 -726 59 -664
rect 800 -726 801 -664
rect 65 -667 66 -653
rect 149 -726 150 -666
rect 152 -667 153 -653
rect 243 -726 244 -666
rect 261 -726 262 -666
rect 289 -726 290 -666
rect 380 -667 381 -653
rect 387 -726 388 -666
rect 408 -667 409 -653
rect 611 -667 612 -653
rect 667 -667 668 -653
rect 709 -726 710 -666
rect 730 -667 731 -653
rect 758 -726 759 -666
rect 23 -669 24 -653
rect 65 -726 66 -668
rect 86 -726 87 -668
rect 310 -669 311 -653
rect 411 -669 412 -653
rect 807 -726 808 -668
rect 23 -726 24 -670
rect 257 -726 258 -670
rect 303 -671 304 -653
rect 380 -726 381 -670
rect 422 -671 423 -653
rect 702 -671 703 -653
rect 30 -726 31 -672
rect 411 -726 412 -672
rect 429 -673 430 -653
rect 492 -726 493 -672
rect 590 -673 591 -653
rect 611 -726 612 -672
rect 618 -673 619 -653
rect 702 -726 703 -672
rect 37 -726 38 -674
rect 408 -726 409 -674
rect 443 -726 444 -674
rect 478 -675 479 -653
rect 548 -675 549 -653
rect 590 -726 591 -674
rect 604 -675 605 -653
rect 618 -726 619 -674
rect 653 -675 654 -653
rect 667 -726 668 -674
rect 674 -675 675 -653
rect 751 -726 752 -674
rect 44 -677 45 -653
rect 653 -726 654 -676
rect 681 -677 682 -653
rect 716 -726 717 -676
rect 44 -726 45 -678
rect 93 -726 94 -678
rect 107 -726 108 -678
rect 163 -679 164 -653
rect 177 -726 178 -678
rect 401 -679 402 -653
rect 439 -726 440 -678
rect 548 -726 549 -678
rect 576 -679 577 -653
rect 604 -726 605 -678
rect 681 -726 682 -678
rect 723 -679 724 -653
rect 79 -681 80 -653
rect 303 -726 304 -680
rect 310 -726 311 -680
rect 338 -681 339 -653
rect 394 -681 395 -653
rect 422 -726 423 -680
rect 457 -681 458 -653
rect 646 -726 647 -680
rect 688 -681 689 -653
rect 779 -726 780 -680
rect 79 -726 80 -682
rect 390 -683 391 -653
rect 397 -726 398 -682
rect 576 -726 577 -682
rect 632 -683 633 -653
rect 723 -726 724 -682
rect 121 -726 122 -684
rect 527 -685 528 -653
rect 625 -685 626 -653
rect 632 -726 633 -684
rect 639 -685 640 -653
rect 688 -726 689 -684
rect 128 -726 129 -686
rect 268 -687 269 -653
rect 282 -726 283 -686
rect 394 -726 395 -686
rect 467 -726 468 -686
rect 478 -726 479 -686
rect 499 -687 500 -653
rect 639 -726 640 -686
rect 131 -689 132 -653
rect 541 -689 542 -653
rect 569 -689 570 -653
rect 625 -726 626 -688
rect 135 -691 136 -653
rect 212 -726 213 -690
rect 219 -691 220 -653
rect 338 -726 339 -690
rect 359 -691 360 -653
rect 457 -726 458 -690
rect 471 -691 472 -653
rect 534 -726 535 -690
rect 124 -726 125 -692
rect 219 -726 220 -692
rect 226 -693 227 -653
rect 268 -726 269 -692
rect 292 -693 293 -653
rect 674 -726 675 -692
rect 110 -695 111 -653
rect 226 -726 227 -694
rect 236 -726 237 -694
rect 744 -726 745 -694
rect 135 -726 136 -696
rect 145 -697 146 -653
rect 156 -726 157 -696
rect 317 -697 318 -653
rect 331 -697 332 -653
rect 401 -726 402 -696
rect 436 -697 437 -653
rect 499 -726 500 -696
rect 506 -697 507 -653
rect 541 -726 542 -696
rect 142 -699 143 -653
rect 485 -699 486 -653
rect 506 -726 507 -698
rect 737 -699 738 -653
rect 47 -701 48 -653
rect 142 -726 143 -700
rect 163 -726 164 -700
rect 562 -701 563 -653
rect 166 -726 167 -702
rect 562 -726 563 -702
rect 184 -726 185 -704
rect 275 -705 276 -653
rect 296 -705 297 -653
rect 359 -726 360 -704
rect 369 -705 370 -653
rect 737 -726 738 -704
rect 173 -726 174 -706
rect 296 -726 297 -706
rect 317 -726 318 -706
rect 814 -726 815 -706
rect 191 -709 192 -653
rect 191 -726 192 -708
rect 191 -709 192 -653
rect 191 -726 192 -708
rect 198 -726 199 -708
rect 247 -709 248 -653
rect 324 -709 325 -653
rect 369 -726 370 -708
rect 446 -709 447 -653
rect 485 -726 486 -708
rect 205 -711 206 -653
rect 583 -726 584 -710
rect 170 -713 171 -653
rect 205 -726 206 -712
rect 233 -713 234 -653
rect 275 -726 276 -712
rect 324 -726 325 -712
rect 373 -713 374 -653
rect 233 -726 234 -714
rect 520 -715 521 -653
rect 240 -726 241 -716
rect 730 -726 731 -716
rect 247 -726 248 -718
rect 429 -726 430 -718
rect 464 -719 465 -653
rect 520 -726 521 -718
rect 331 -726 332 -720
rect 527 -726 528 -720
rect 334 -726 335 -722
rect 569 -726 570 -722
rect 373 -726 374 -724
rect 436 -726 437 -724
rect 9 -736 10 -734
rect 9 -815 10 -735
rect 9 -736 10 -734
rect 9 -815 10 -735
rect 40 -815 41 -735
rect 121 -815 122 -735
rect 124 -736 125 -734
rect 730 -736 731 -734
rect 817 -736 818 -734
rect 828 -736 829 -734
rect 44 -738 45 -734
rect 68 -738 69 -734
rect 72 -738 73 -734
rect 212 -738 213 -734
rect 236 -738 237 -734
rect 464 -738 465 -734
rect 467 -738 468 -734
rect 793 -738 794 -734
rect 47 -815 48 -739
rect 65 -740 66 -734
rect 72 -815 73 -739
rect 306 -815 307 -739
rect 324 -740 325 -734
rect 464 -815 465 -739
rect 474 -740 475 -734
rect 779 -740 780 -734
rect 51 -742 52 -734
rect 583 -742 584 -734
rect 597 -815 598 -741
rect 632 -742 633 -734
rect 639 -742 640 -734
rect 814 -742 815 -734
rect 58 -744 59 -734
rect 653 -744 654 -734
rect 681 -744 682 -734
rect 779 -815 780 -743
rect 58 -815 59 -745
rect 338 -746 339 -734
rect 341 -815 342 -745
rect 807 -746 808 -734
rect 75 -748 76 -734
rect 653 -815 654 -747
rect 660 -748 661 -734
rect 681 -815 682 -747
rect 96 -815 97 -749
rect 660 -815 661 -749
rect 100 -752 101 -734
rect 100 -815 101 -751
rect 100 -752 101 -734
rect 100 -815 101 -751
rect 117 -752 118 -734
rect 702 -752 703 -734
rect 142 -754 143 -734
rect 212 -815 213 -753
rect 240 -754 241 -734
rect 824 -754 825 -734
rect 79 -756 80 -734
rect 240 -815 241 -755
rect 254 -815 255 -755
rect 268 -756 269 -734
rect 289 -756 290 -734
rect 765 -756 766 -734
rect 86 -758 87 -734
rect 268 -815 269 -757
rect 282 -758 283 -734
rect 289 -815 290 -757
rect 292 -758 293 -734
rect 485 -758 486 -734
rect 506 -758 507 -734
rect 730 -815 731 -757
rect 86 -815 87 -759
rect 233 -760 234 -734
rect 275 -760 276 -734
rect 282 -815 283 -759
rect 310 -760 311 -734
rect 506 -815 507 -759
rect 583 -815 584 -759
rect 688 -760 689 -734
rect 37 -762 38 -734
rect 310 -815 311 -761
rect 324 -815 325 -761
rect 345 -762 346 -734
rect 348 -815 349 -761
rect 793 -815 794 -761
rect 37 -815 38 -763
rect 800 -764 801 -734
rect 107 -766 108 -734
rect 233 -815 234 -765
rect 331 -766 332 -734
rect 352 -766 353 -734
rect 366 -766 367 -734
rect 702 -815 703 -765
rect 107 -815 108 -767
rect 471 -768 472 -734
rect 548 -768 549 -734
rect 688 -815 689 -767
rect 82 -815 83 -769
rect 548 -815 549 -769
rect 590 -770 591 -734
rect 765 -815 766 -769
rect 135 -772 136 -734
rect 275 -815 276 -771
rect 296 -772 297 -734
rect 331 -815 332 -771
rect 352 -815 353 -771
rect 369 -815 370 -771
rect 394 -772 395 -734
rect 492 -772 493 -734
rect 600 -772 601 -734
rect 751 -772 752 -734
rect 135 -815 136 -773
rect 366 -815 367 -773
rect 387 -774 388 -734
rect 394 -815 395 -773
rect 408 -774 409 -734
rect 443 -774 444 -734
rect 450 -774 451 -734
rect 674 -774 675 -734
rect 709 -774 710 -734
rect 751 -815 752 -773
rect 142 -815 143 -775
rect 184 -776 185 -734
rect 191 -776 192 -734
rect 191 -815 192 -775
rect 191 -776 192 -734
rect 191 -815 192 -775
rect 226 -776 227 -734
rect 345 -815 346 -775
rect 408 -815 409 -775
rect 415 -776 416 -734
rect 429 -776 430 -734
rect 520 -776 521 -734
rect 611 -776 612 -734
rect 611 -815 612 -775
rect 611 -776 612 -734
rect 611 -815 612 -775
rect 632 -815 633 -775
rect 667 -776 668 -734
rect 159 -778 160 -734
rect 772 -778 773 -734
rect 163 -815 164 -779
rect 401 -780 402 -734
rect 411 -780 412 -734
rect 625 -780 626 -734
rect 639 -815 640 -779
rect 737 -780 738 -734
rect 170 -815 171 -781
rect 205 -782 206 -734
rect 296 -815 297 -781
rect 439 -815 440 -781
rect 446 -815 447 -781
rect 674 -815 675 -781
rect 198 -784 199 -734
rect 226 -815 227 -783
rect 380 -784 381 -734
rect 415 -815 416 -783
rect 436 -784 437 -734
rect 723 -784 724 -734
rect 16 -786 17 -734
rect 723 -815 724 -785
rect 198 -815 199 -787
rect 373 -788 374 -734
rect 380 -815 381 -787
rect 744 -788 745 -734
rect 205 -815 206 -789
rect 247 -790 248 -734
rect 359 -790 360 -734
rect 373 -815 374 -789
rect 404 -815 405 -789
rect 737 -815 738 -789
rect 23 -792 24 -734
rect 247 -815 248 -791
rect 338 -815 339 -791
rect 359 -815 360 -791
rect 436 -815 437 -791
rect 744 -815 745 -791
rect 23 -815 24 -793
rect 156 -794 157 -734
rect 457 -794 458 -734
rect 485 -815 486 -793
rect 492 -815 493 -793
rect 541 -794 542 -734
rect 604 -794 605 -734
rect 667 -815 668 -793
rect 93 -796 94 -734
rect 156 -815 157 -795
rect 422 -796 423 -734
rect 457 -815 458 -795
rect 471 -815 472 -795
rect 513 -796 514 -734
rect 520 -815 521 -795
rect 576 -796 577 -734
rect 625 -815 626 -795
rect 695 -796 696 -734
rect 93 -815 94 -797
rect 261 -798 262 -734
rect 453 -815 454 -797
rect 513 -815 514 -797
rect 534 -798 535 -734
rect 541 -815 542 -797
rect 562 -798 563 -734
rect 576 -815 577 -797
rect 618 -798 619 -734
rect 695 -815 696 -797
rect 16 -815 17 -799
rect 562 -815 563 -799
rect 569 -800 570 -734
rect 604 -815 605 -799
rect 646 -800 647 -734
rect 709 -815 710 -799
rect 149 -802 150 -734
rect 422 -815 423 -801
rect 499 -802 500 -734
rect 772 -815 773 -801
rect 114 -815 115 -803
rect 149 -815 150 -803
rect 261 -815 262 -803
rect 387 -815 388 -803
rect 478 -804 479 -734
rect 499 -815 500 -803
rect 527 -804 528 -734
rect 534 -815 535 -803
rect 555 -804 556 -734
rect 569 -815 570 -803
rect 646 -815 647 -803
rect 821 -804 822 -734
rect 177 -806 178 -734
rect 527 -815 528 -805
rect 555 -815 556 -805
rect 786 -806 787 -734
rect 128 -808 129 -734
rect 177 -815 178 -807
rect 219 -808 220 -734
rect 478 -815 479 -807
rect 758 -808 759 -734
rect 786 -815 787 -807
rect 30 -810 31 -734
rect 128 -815 129 -809
rect 219 -815 220 -809
rect 317 -810 318 -734
rect 716 -810 717 -734
rect 758 -815 759 -809
rect 30 -815 31 -811
rect 187 -815 188 -811
rect 271 -815 272 -811
rect 618 -815 619 -811
rect 303 -814 304 -734
rect 317 -815 318 -813
rect 390 -815 391 -813
rect 716 -815 717 -813
rect 9 -825 10 -823
rect 93 -825 94 -823
rect 96 -825 97 -823
rect 240 -825 241 -823
rect 303 -825 304 -823
rect 772 -825 773 -823
rect 23 -827 24 -823
rect 51 -827 52 -823
rect 54 -900 55 -826
rect 362 -900 363 -826
rect 369 -827 370 -823
rect 709 -827 710 -823
rect 37 -829 38 -823
rect 723 -829 724 -823
rect 37 -900 38 -830
rect 285 -900 286 -830
rect 331 -831 332 -823
rect 744 -831 745 -823
rect 26 -900 27 -832
rect 331 -900 332 -832
rect 348 -833 349 -823
rect 527 -833 528 -823
rect 530 -900 531 -832
rect 779 -833 780 -823
rect 51 -900 52 -834
rect 212 -835 213 -823
rect 352 -835 353 -823
rect 730 -835 731 -823
rect 58 -837 59 -823
rect 240 -900 241 -836
rect 359 -837 360 -823
rect 383 -837 384 -823
rect 390 -837 391 -823
rect 765 -837 766 -823
rect 58 -900 59 -838
rect 191 -839 192 -823
rect 212 -900 213 -838
rect 254 -839 255 -823
rect 373 -839 374 -823
rect 387 -839 388 -823
rect 404 -839 405 -823
rect 569 -839 570 -823
rect 590 -839 591 -823
rect 688 -839 689 -823
rect 709 -900 710 -838
rect 758 -839 759 -823
rect 30 -841 31 -823
rect 191 -900 192 -840
rect 257 -900 258 -840
rect 373 -900 374 -840
rect 380 -900 381 -840
rect 576 -841 577 -823
rect 625 -841 626 -823
rect 625 -900 626 -840
rect 625 -841 626 -823
rect 625 -900 626 -840
rect 632 -841 633 -823
rect 635 -841 636 -823
rect 681 -841 682 -823
rect 758 -900 759 -840
rect 30 -900 31 -842
rect 100 -843 101 -823
rect 128 -843 129 -823
rect 184 -900 185 -842
rect 187 -843 188 -823
rect 282 -843 283 -823
rect 306 -843 307 -823
rect 688 -900 689 -842
rect 65 -845 66 -823
rect 653 -845 654 -823
rect 65 -900 66 -846
rect 68 -847 69 -823
rect 72 -847 73 -823
rect 107 -847 108 -823
rect 114 -847 115 -823
rect 128 -900 129 -846
rect 145 -900 146 -846
rect 737 -847 738 -823
rect 16 -900 17 -848
rect 114 -900 115 -848
rect 149 -849 150 -823
rect 317 -849 318 -823
rect 324 -849 325 -823
rect 387 -900 388 -848
rect 394 -849 395 -823
rect 404 -900 405 -848
rect 411 -900 412 -848
rect 702 -849 703 -823
rect 716 -849 717 -823
rect 737 -900 738 -848
rect 44 -851 45 -823
rect 702 -900 703 -850
rect 44 -900 45 -852
rect 247 -853 248 -823
rect 310 -853 311 -823
rect 324 -900 325 -852
rect 338 -853 339 -823
rect 576 -900 577 -852
rect 611 -853 612 -823
rect 681 -900 682 -852
rect 72 -900 73 -854
rect 198 -855 199 -823
rect 219 -855 220 -823
rect 310 -900 311 -854
rect 394 -900 395 -854
rect 408 -855 409 -823
rect 422 -855 423 -823
rect 653 -900 654 -854
rect 82 -857 83 -823
rect 506 -857 507 -823
rect 537 -900 538 -856
rect 695 -857 696 -823
rect 86 -859 87 -823
rect 198 -900 199 -858
rect 226 -859 227 -823
rect 247 -900 248 -858
rect 422 -900 423 -858
rect 562 -859 563 -823
rect 569 -900 570 -858
rect 667 -859 668 -823
rect 86 -900 87 -860
rect 121 -861 122 -823
rect 149 -900 150 -860
rect 261 -861 262 -823
rect 429 -861 430 -823
rect 485 -861 486 -823
rect 555 -861 556 -823
rect 793 -861 794 -823
rect 93 -900 94 -862
rect 142 -863 143 -823
rect 152 -863 153 -823
rect 275 -863 276 -823
rect 299 -900 300 -862
rect 429 -900 430 -862
rect 436 -863 437 -823
rect 520 -863 521 -823
rect 555 -900 556 -862
rect 618 -863 619 -823
rect 632 -900 633 -862
rect 639 -863 640 -823
rect 667 -900 668 -862
rect 751 -863 752 -823
rect 107 -900 108 -864
rect 359 -900 360 -864
rect 436 -900 437 -864
rect 478 -865 479 -823
rect 485 -900 486 -864
rect 548 -865 549 -823
rect 562 -900 563 -864
rect 660 -865 661 -823
rect 121 -900 122 -866
rect 170 -867 171 -823
rect 173 -900 174 -866
rect 296 -867 297 -823
rect 306 -900 307 -866
rect 478 -900 479 -866
rect 513 -867 514 -823
rect 660 -900 661 -866
rect 142 -900 143 -868
rect 219 -900 220 -868
rect 275 -900 276 -868
rect 443 -869 444 -823
rect 450 -900 451 -868
rect 618 -900 619 -868
rect 156 -871 157 -823
rect 159 -875 160 -870
rect 163 -871 164 -823
rect 317 -900 318 -870
rect 345 -871 346 -823
rect 520 -900 521 -870
rect 156 -900 157 -872
rect 345 -900 346 -872
rect 415 -873 416 -823
rect 443 -900 444 -872
rect 499 -873 500 -823
rect 513 -900 514 -872
rect 604 -873 605 -823
rect 117 -900 118 -874
rect 415 -900 416 -874
rect 453 -875 454 -823
rect 492 -875 493 -823
rect 597 -875 598 -823
rect 604 -900 605 -874
rect 635 -900 636 -874
rect 639 -900 640 -874
rect 163 -900 164 -876
rect 268 -877 269 -823
rect 453 -900 454 -876
rect 786 -877 787 -823
rect 170 -900 171 -878
rect 341 -900 342 -878
rect 457 -879 458 -823
rect 499 -900 500 -878
rect 135 -881 136 -823
rect 457 -900 458 -880
rect 471 -881 472 -823
rect 471 -900 472 -880
rect 471 -881 472 -823
rect 471 -900 472 -880
rect 492 -900 493 -880
rect 541 -881 542 -823
rect 135 -900 136 -882
rect 226 -900 227 -882
rect 268 -900 269 -882
rect 289 -883 290 -823
rect 541 -900 542 -882
rect 646 -883 647 -823
rect 79 -900 80 -884
rect 289 -900 290 -884
rect 583 -885 584 -823
rect 646 -900 647 -884
rect 177 -887 178 -823
rect 352 -900 353 -886
rect 583 -900 584 -886
rect 674 -887 675 -823
rect 177 -900 178 -888
rect 233 -889 234 -823
rect 674 -900 675 -888
rect 695 -900 696 -888
rect 180 -900 181 -890
rect 261 -900 262 -890
rect 233 -900 234 -892
rect 366 -893 367 -823
rect 366 -900 367 -894
rect 464 -895 465 -823
rect 464 -900 465 -896
rect 534 -897 535 -823
rect 534 -900 535 -898
rect 597 -900 598 -898
rect 2 -983 3 -909
rect 100 -910 101 -908
rect 103 -910 104 -908
rect 233 -910 234 -908
rect 240 -910 241 -908
rect 306 -910 307 -908
rect 317 -910 318 -908
rect 317 -983 318 -909
rect 317 -910 318 -908
rect 317 -983 318 -909
rect 338 -983 339 -909
rect 352 -910 353 -908
rect 359 -983 360 -909
rect 537 -910 538 -908
rect 548 -983 549 -909
rect 562 -910 563 -908
rect 576 -910 577 -908
rect 590 -910 591 -908
rect 607 -983 608 -909
rect 681 -910 682 -908
rect 695 -910 696 -908
rect 758 -910 759 -908
rect 23 -912 24 -908
rect 499 -912 500 -908
rect 509 -912 510 -908
rect 632 -912 633 -908
rect 737 -912 738 -908
rect 751 -983 752 -911
rect 26 -983 27 -913
rect 170 -983 171 -913
rect 205 -914 206 -908
rect 254 -914 255 -908
rect 257 -914 258 -908
rect 681 -983 682 -913
rect 30 -916 31 -908
rect 145 -916 146 -908
rect 205 -983 206 -915
rect 397 -983 398 -915
rect 404 -916 405 -908
rect 646 -916 647 -908
rect 30 -983 31 -917
rect 187 -983 188 -917
rect 212 -918 213 -908
rect 289 -983 290 -917
rect 296 -983 297 -917
rect 310 -918 311 -908
rect 383 -983 384 -917
rect 394 -918 395 -908
rect 408 -983 409 -917
rect 611 -983 612 -917
rect 618 -918 619 -908
rect 632 -983 633 -917
rect 37 -983 38 -919
rect 47 -983 48 -919
rect 54 -983 55 -919
rect 688 -920 689 -908
rect 40 -922 41 -908
rect 702 -922 703 -908
rect 65 -924 66 -908
rect 145 -983 146 -923
rect 156 -924 157 -908
rect 212 -983 213 -923
rect 229 -983 230 -923
rect 590 -983 591 -923
rect 597 -924 598 -908
rect 695 -983 696 -923
rect 65 -983 66 -925
rect 555 -926 556 -908
rect 576 -983 577 -925
rect 604 -926 605 -908
rect 621 -983 622 -925
rect 709 -926 710 -908
rect 72 -928 73 -908
rect 254 -983 255 -927
rect 275 -928 276 -908
rect 702 -983 703 -927
rect 72 -983 73 -929
rect 366 -930 367 -908
rect 387 -930 388 -908
rect 450 -930 451 -908
rect 478 -930 479 -908
rect 709 -983 710 -929
rect 79 -932 80 -908
rect 173 -932 174 -908
rect 219 -932 220 -908
rect 366 -983 367 -931
rect 394 -983 395 -931
rect 660 -932 661 -908
rect 688 -983 689 -931
rect 726 -983 727 -931
rect 61 -983 62 -933
rect 79 -983 80 -933
rect 86 -934 87 -908
rect 250 -983 251 -933
rect 275 -983 276 -933
rect 345 -934 346 -908
rect 362 -934 363 -908
rect 660 -983 661 -933
rect 93 -936 94 -908
rect 152 -983 153 -935
rect 156 -983 157 -935
rect 163 -936 164 -908
rect 226 -936 227 -908
rect 387 -983 388 -935
rect 415 -936 416 -908
rect 716 -983 717 -935
rect 93 -983 94 -937
rect 198 -938 199 -908
rect 233 -983 234 -937
rect 299 -938 300 -908
rect 303 -983 304 -937
rect 362 -983 363 -937
rect 436 -938 437 -908
rect 436 -983 437 -937
rect 436 -938 437 -908
rect 436 -983 437 -937
rect 450 -983 451 -937
rect 471 -938 472 -908
rect 478 -983 479 -937
rect 527 -938 528 -908
rect 534 -983 535 -937
rect 569 -938 570 -908
rect 625 -938 626 -908
rect 628 -946 629 -937
rect 44 -940 45 -908
rect 198 -983 199 -939
rect 240 -983 241 -939
rect 268 -940 269 -908
rect 278 -940 279 -908
rect 324 -940 325 -908
rect 499 -983 500 -939
rect 646 -983 647 -939
rect 44 -983 45 -941
rect 569 -983 570 -941
rect 625 -983 626 -941
rect 639 -942 640 -908
rect 107 -944 108 -908
rect 502 -983 503 -943
rect 513 -944 514 -908
rect 527 -983 528 -943
rect 555 -983 556 -943
rect 674 -944 675 -908
rect 107 -983 108 -945
rect 352 -983 353 -945
rect 513 -983 514 -945
rect 583 -946 584 -908
rect 639 -983 640 -945
rect 114 -983 115 -947
rect 128 -948 129 -908
rect 135 -948 136 -908
rect 471 -983 472 -947
rect 520 -948 521 -908
rect 674 -983 675 -947
rect 16 -950 17 -908
rect 128 -983 129 -949
rect 163 -983 164 -949
rect 180 -950 181 -908
rect 261 -950 262 -908
rect 345 -983 346 -949
rect 520 -983 521 -949
rect 541 -950 542 -908
rect 562 -983 563 -949
rect 604 -983 605 -949
rect 16 -983 17 -951
rect 191 -952 192 -908
rect 261 -983 262 -951
rect 411 -952 412 -908
rect 100 -983 101 -953
rect 135 -983 136 -953
rect 149 -954 150 -908
rect 191 -983 192 -953
rect 282 -983 283 -953
rect 492 -954 493 -908
rect 117 -956 118 -908
rect 247 -956 248 -908
rect 285 -956 286 -908
rect 422 -956 423 -908
rect 485 -956 486 -908
rect 492 -983 493 -955
rect 121 -958 122 -908
rect 219 -983 220 -957
rect 310 -983 311 -957
rect 653 -958 654 -908
rect 58 -960 59 -908
rect 121 -983 122 -959
rect 142 -983 143 -959
rect 422 -983 423 -959
rect 653 -983 654 -959
rect 667 -960 668 -908
rect 9 -962 10 -908
rect 58 -983 59 -961
rect 149 -983 150 -961
rect 415 -983 416 -961
rect 180 -983 181 -963
rect 457 -964 458 -908
rect 324 -983 325 -965
rect 506 -966 507 -908
rect 313 -983 314 -967
rect 506 -983 507 -967
rect 331 -970 332 -908
rect 583 -983 584 -969
rect 51 -983 52 -971
rect 331 -983 332 -971
rect 373 -972 374 -908
rect 541 -983 542 -971
rect 184 -974 185 -908
rect 373 -983 374 -973
rect 401 -974 402 -908
rect 667 -983 668 -973
rect 184 -983 185 -975
rect 268 -983 269 -975
rect 401 -983 402 -975
rect 411 -983 412 -975
rect 457 -983 458 -975
rect 464 -976 465 -908
rect 429 -978 430 -908
rect 464 -983 465 -977
rect 429 -983 430 -979
rect 443 -980 444 -908
rect 380 -982 381 -908
rect 443 -983 444 -981
rect 9 -993 10 -991
rect 184 -993 185 -991
rect 187 -993 188 -991
rect 254 -993 255 -991
rect 275 -993 276 -991
rect 355 -1058 356 -992
rect 404 -1058 405 -992
rect 436 -993 437 -991
rect 443 -1058 444 -992
rect 450 -993 451 -991
rect 464 -993 465 -991
rect 485 -993 486 -991
rect 499 -1058 500 -992
rect 506 -993 507 -991
rect 520 -993 521 -991
rect 523 -1011 524 -992
rect 527 -993 528 -991
rect 730 -1058 731 -992
rect 751 -993 752 -991
rect 758 -1058 759 -992
rect 26 -995 27 -991
rect 65 -1058 66 -994
rect 79 -995 80 -991
rect 86 -995 87 -991
rect 89 -995 90 -991
rect 611 -995 612 -991
rect 618 -1058 619 -994
rect 632 -995 633 -991
rect 639 -995 640 -991
rect 639 -1058 640 -994
rect 639 -995 640 -991
rect 639 -1058 640 -994
rect 653 -995 654 -991
rect 653 -1058 654 -994
rect 653 -995 654 -991
rect 653 -1058 654 -994
rect 716 -995 717 -991
rect 723 -1058 724 -994
rect 30 -997 31 -991
rect 362 -1058 363 -996
rect 425 -1058 426 -996
rect 527 -1058 528 -996
rect 548 -997 549 -991
rect 548 -1058 549 -996
rect 548 -997 549 -991
rect 548 -1058 549 -996
rect 604 -997 605 -991
rect 621 -997 622 -991
rect 625 -997 626 -991
rect 632 -1058 633 -996
rect 709 -997 710 -991
rect 716 -1058 717 -996
rect 37 -999 38 -991
rect 142 -999 143 -991
rect 149 -999 150 -991
rect 394 -999 395 -991
rect 436 -1058 437 -998
rect 457 -999 458 -991
rect 464 -1058 465 -998
rect 492 -999 493 -991
rect 502 -999 503 -991
rect 576 -999 577 -991
rect 695 -999 696 -991
rect 709 -1058 710 -998
rect 37 -1058 38 -1000
rect 72 -1001 73 -991
rect 79 -1058 80 -1000
rect 429 -1001 430 -991
rect 457 -1058 458 -1000
rect 471 -1001 472 -991
rect 478 -1001 479 -991
rect 506 -1058 507 -1000
rect 520 -1058 521 -1000
rect 562 -1001 563 -991
rect 695 -1058 696 -1000
rect 702 -1001 703 -991
rect 44 -1003 45 -991
rect 681 -1003 682 -991
rect 688 -1003 689 -991
rect 702 -1058 703 -1002
rect 47 -1005 48 -991
rect 198 -1005 199 -991
rect 205 -1005 206 -991
rect 446 -1005 447 -991
rect 485 -1058 486 -1004
rect 607 -1005 608 -991
rect 674 -1005 675 -991
rect 688 -1058 689 -1004
rect 54 -1058 55 -1006
rect 569 -1007 570 -991
rect 660 -1007 661 -991
rect 674 -1058 675 -1006
rect 58 -1058 59 -1008
rect 415 -1009 416 -991
rect 488 -1009 489 -991
rect 576 -1058 577 -1008
rect 660 -1058 661 -1008
rect 667 -1009 668 -991
rect 68 -1011 69 -991
rect 478 -1058 479 -1010
rect 562 -1058 563 -1010
rect 569 -1058 570 -1010
rect 583 -1011 584 -991
rect 86 -1058 87 -1012
rect 331 -1013 332 -991
rect 352 -1013 353 -991
rect 471 -1058 472 -1012
rect 555 -1013 556 -991
rect 681 -1058 682 -1012
rect 93 -1015 94 -991
rect 184 -1058 185 -1014
rect 191 -1015 192 -991
rect 198 -1058 199 -1014
rect 205 -1058 206 -1014
rect 345 -1015 346 -991
rect 366 -1015 367 -991
rect 583 -1058 584 -1014
rect 2 -1017 3 -991
rect 345 -1058 346 -1016
rect 366 -1058 367 -1016
rect 380 -1058 381 -1016
rect 383 -1017 384 -991
rect 429 -1058 430 -1016
rect 534 -1017 535 -991
rect 555 -1058 556 -1016
rect 93 -1058 94 -1018
rect 100 -1019 101 -991
rect 107 -1019 108 -991
rect 646 -1019 647 -991
rect 16 -1021 17 -991
rect 107 -1058 108 -1020
rect 114 -1021 115 -991
rect 289 -1058 290 -1020
rect 292 -1021 293 -991
rect 597 -1058 598 -1020
rect 16 -1058 17 -1022
rect 170 -1023 171 -991
rect 180 -1023 181 -991
rect 373 -1023 374 -991
rect 394 -1058 395 -1022
rect 541 -1023 542 -991
rect 100 -1058 101 -1024
rect 212 -1025 213 -991
rect 219 -1025 220 -991
rect 226 -1025 227 -991
rect 240 -1025 241 -991
rect 313 -1025 314 -991
rect 317 -1025 318 -991
rect 369 -1058 370 -1024
rect 373 -1058 374 -1024
rect 513 -1025 514 -991
rect 534 -1058 535 -1024
rect 590 -1025 591 -991
rect 23 -1058 24 -1026
rect 590 -1058 591 -1026
rect 75 -1058 76 -1028
rect 240 -1058 241 -1028
rect 247 -1058 248 -1028
rect 261 -1029 262 -991
rect 268 -1029 269 -991
rect 611 -1058 612 -1028
rect 117 -1058 118 -1030
rect 219 -1058 220 -1030
rect 226 -1058 227 -1030
rect 324 -1031 325 -991
rect 331 -1058 332 -1030
rect 359 -1058 360 -1030
rect 142 -1058 143 -1032
rect 401 -1033 402 -991
rect 156 -1035 157 -991
rect 170 -1058 171 -1034
rect 177 -1035 178 -991
rect 541 -1058 542 -1034
rect 128 -1037 129 -991
rect 177 -1058 178 -1036
rect 212 -1058 213 -1036
rect 310 -1037 311 -991
rect 317 -1058 318 -1036
rect 338 -1037 339 -991
rect 401 -1058 402 -1036
rect 667 -1058 668 -1036
rect 103 -1058 104 -1038
rect 128 -1058 129 -1038
rect 135 -1039 136 -991
rect 156 -1058 157 -1038
rect 163 -1039 164 -991
rect 191 -1058 192 -1038
rect 250 -1039 251 -991
rect 646 -1058 647 -1038
rect 121 -1041 122 -991
rect 163 -1058 164 -1040
rect 254 -1058 255 -1040
rect 422 -1041 423 -991
rect 30 -1058 31 -1042
rect 121 -1058 122 -1042
rect 135 -1058 136 -1042
rect 149 -1058 150 -1042
rect 261 -1058 262 -1042
rect 296 -1043 297 -991
rect 306 -1058 307 -1042
rect 338 -1058 339 -1042
rect 422 -1058 423 -1042
rect 513 -1058 514 -1042
rect 233 -1045 234 -991
rect 296 -1058 297 -1044
rect 310 -1058 311 -1044
rect 625 -1058 626 -1044
rect 233 -1058 234 -1046
rect 450 -1058 451 -1046
rect 268 -1058 269 -1048
rect 408 -1058 409 -1048
rect 275 -1058 276 -1050
rect 303 -1051 304 -991
rect 320 -1058 321 -1050
rect 387 -1051 388 -991
rect 282 -1053 283 -991
rect 411 -1053 412 -991
rect 303 -1058 304 -1054
rect 492 -1058 493 -1054
rect 324 -1058 325 -1056
rect 352 -1058 353 -1056
rect 387 -1058 388 -1056
rect 397 -1057 398 -991
rect 16 -1068 17 -1066
rect 359 -1125 360 -1067
rect 362 -1068 363 -1066
rect 695 -1068 696 -1066
rect 702 -1068 703 -1066
rect 702 -1125 703 -1067
rect 702 -1068 703 -1066
rect 702 -1125 703 -1067
rect 730 -1068 731 -1066
rect 737 -1125 738 -1067
rect 751 -1125 752 -1067
rect 754 -1068 755 -1066
rect 758 -1068 759 -1066
rect 758 -1125 759 -1067
rect 758 -1068 759 -1066
rect 758 -1125 759 -1067
rect 16 -1125 17 -1069
rect 261 -1070 262 -1066
rect 268 -1125 269 -1069
rect 289 -1070 290 -1066
rect 306 -1070 307 -1066
rect 681 -1070 682 -1066
rect 754 -1125 755 -1069
rect 793 -1125 794 -1069
rect 26 -1072 27 -1066
rect 86 -1072 87 -1066
rect 89 -1125 90 -1071
rect 173 -1072 174 -1066
rect 177 -1072 178 -1066
rect 261 -1125 262 -1071
rect 310 -1072 311 -1066
rect 345 -1072 346 -1066
rect 369 -1125 370 -1071
rect 548 -1072 549 -1066
rect 597 -1072 598 -1066
rect 730 -1125 731 -1071
rect 9 -1074 10 -1066
rect 86 -1125 87 -1073
rect 93 -1074 94 -1066
rect 93 -1125 94 -1073
rect 93 -1074 94 -1066
rect 93 -1125 94 -1073
rect 107 -1074 108 -1066
rect 303 -1074 304 -1066
rect 310 -1125 311 -1073
rect 324 -1074 325 -1066
rect 327 -1125 328 -1073
rect 373 -1125 374 -1073
rect 383 -1125 384 -1073
rect 506 -1074 507 -1066
rect 509 -1125 510 -1073
rect 681 -1125 682 -1073
rect 9 -1125 10 -1075
rect 121 -1076 122 -1066
rect 156 -1076 157 -1066
rect 187 -1076 188 -1066
rect 205 -1076 206 -1066
rect 376 -1076 377 -1066
rect 394 -1125 395 -1075
rect 439 -1125 440 -1075
rect 464 -1076 465 -1066
rect 786 -1125 787 -1075
rect 30 -1078 31 -1066
rect 471 -1078 472 -1066
rect 474 -1125 475 -1077
rect 576 -1078 577 -1066
rect 604 -1078 605 -1066
rect 653 -1078 654 -1066
rect 660 -1078 661 -1066
rect 695 -1125 696 -1077
rect 37 -1080 38 -1066
rect 138 -1080 139 -1066
rect 156 -1125 157 -1079
rect 166 -1125 167 -1079
rect 170 -1125 171 -1079
rect 271 -1080 272 -1066
rect 331 -1080 332 -1066
rect 597 -1125 598 -1079
rect 632 -1080 633 -1066
rect 653 -1125 654 -1079
rect 667 -1080 668 -1066
rect 779 -1125 780 -1079
rect 44 -1125 45 -1081
rect 219 -1082 220 -1066
rect 226 -1082 227 -1066
rect 226 -1125 227 -1081
rect 226 -1082 227 -1066
rect 226 -1125 227 -1081
rect 247 -1082 248 -1066
rect 415 -1082 416 -1066
rect 418 -1082 419 -1066
rect 723 -1082 724 -1066
rect 47 -1084 48 -1066
rect 65 -1084 66 -1066
rect 72 -1125 73 -1083
rect 135 -1084 136 -1066
rect 138 -1125 139 -1083
rect 583 -1084 584 -1066
rect 625 -1084 626 -1066
rect 667 -1125 668 -1083
rect 709 -1084 710 -1066
rect 723 -1125 724 -1083
rect 23 -1125 24 -1085
rect 65 -1125 66 -1085
rect 100 -1125 101 -1085
rect 187 -1125 188 -1085
rect 198 -1086 199 -1066
rect 219 -1125 220 -1085
rect 250 -1125 251 -1085
rect 275 -1086 276 -1066
rect 345 -1125 346 -1085
rect 425 -1086 426 -1066
rect 450 -1086 451 -1066
rect 625 -1125 626 -1085
rect 632 -1125 633 -1085
rect 674 -1086 675 -1066
rect 688 -1086 689 -1066
rect 709 -1125 710 -1085
rect 58 -1088 59 -1066
rect 107 -1125 108 -1087
rect 114 -1088 115 -1066
rect 191 -1088 192 -1066
rect 208 -1125 209 -1087
rect 254 -1088 255 -1066
rect 275 -1125 276 -1087
rect 338 -1088 339 -1066
rect 380 -1088 381 -1066
rect 604 -1125 605 -1087
rect 639 -1088 640 -1066
rect 660 -1125 661 -1087
rect 58 -1125 59 -1089
rect 142 -1090 143 -1066
rect 163 -1090 164 -1066
rect 331 -1125 332 -1089
rect 380 -1125 381 -1089
rect 740 -1125 741 -1089
rect 114 -1125 115 -1091
rect 212 -1092 213 -1066
rect 387 -1092 388 -1066
rect 415 -1125 416 -1091
rect 425 -1125 426 -1091
rect 716 -1092 717 -1066
rect 79 -1094 80 -1066
rect 387 -1125 388 -1093
rect 397 -1094 398 -1066
rect 583 -1125 584 -1093
rect 611 -1094 612 -1066
rect 639 -1125 640 -1093
rect 646 -1094 647 -1066
rect 674 -1125 675 -1093
rect 117 -1125 118 -1095
rect 296 -1096 297 -1066
rect 401 -1125 402 -1095
rect 408 -1096 409 -1066
rect 436 -1096 437 -1066
rect 450 -1125 451 -1095
rect 457 -1096 458 -1066
rect 464 -1125 465 -1095
rect 471 -1125 472 -1095
rect 716 -1125 717 -1095
rect 51 -1098 52 -1066
rect 457 -1125 458 -1097
rect 499 -1098 500 -1066
rect 814 -1125 815 -1097
rect 51 -1125 52 -1099
rect 205 -1125 206 -1099
rect 212 -1125 213 -1099
rect 317 -1100 318 -1066
rect 436 -1125 437 -1099
rect 562 -1100 563 -1066
rect 618 -1100 619 -1066
rect 646 -1125 647 -1099
rect 37 -1125 38 -1101
rect 317 -1125 318 -1101
rect 513 -1102 514 -1066
rect 548 -1125 549 -1101
rect 562 -1125 563 -1101
rect 569 -1102 570 -1066
rect 103 -1104 104 -1066
rect 499 -1125 500 -1103
rect 520 -1104 521 -1066
rect 520 -1125 521 -1103
rect 520 -1104 521 -1066
rect 520 -1125 521 -1103
rect 534 -1104 535 -1066
rect 576 -1125 577 -1103
rect 121 -1125 122 -1105
rect 422 -1125 423 -1105
rect 527 -1106 528 -1066
rect 534 -1125 535 -1105
rect 541 -1106 542 -1066
rect 541 -1125 542 -1105
rect 541 -1106 542 -1066
rect 541 -1125 542 -1105
rect 128 -1108 129 -1066
rect 142 -1125 143 -1107
rect 163 -1125 164 -1107
rect 478 -1108 479 -1066
rect 527 -1125 528 -1107
rect 555 -1108 556 -1066
rect 128 -1125 129 -1109
rect 149 -1110 150 -1066
rect 177 -1125 178 -1109
rect 282 -1110 283 -1066
rect 289 -1125 290 -1109
rect 569 -1125 570 -1109
rect 79 -1125 80 -1111
rect 149 -1125 150 -1111
rect 180 -1125 181 -1111
rect 324 -1125 325 -1111
rect 429 -1112 430 -1066
rect 478 -1125 479 -1111
rect 555 -1125 556 -1111
rect 590 -1112 591 -1066
rect 184 -1114 185 -1066
rect 198 -1125 199 -1113
rect 240 -1114 241 -1066
rect 296 -1125 297 -1113
rect 366 -1114 367 -1066
rect 590 -1125 591 -1113
rect 184 -1125 185 -1115
rect 233 -1116 234 -1066
rect 240 -1125 241 -1115
rect 247 -1125 248 -1115
rect 282 -1125 283 -1115
rect 338 -1125 339 -1115
rect 366 -1125 367 -1115
rect 513 -1125 514 -1115
rect 191 -1125 192 -1117
rect 303 -1125 304 -1117
rect 429 -1125 430 -1117
rect 443 -1118 444 -1066
rect 194 -1125 195 -1119
rect 254 -1125 255 -1119
rect 443 -1125 444 -1119
rect 492 -1120 493 -1066
rect 233 -1125 234 -1121
rect 408 -1125 409 -1121
rect 485 -1122 486 -1066
rect 492 -1125 493 -1121
rect 320 -1125 321 -1123
rect 485 -1125 486 -1123
rect 9 -1135 10 -1133
rect 327 -1135 328 -1133
rect 348 -1206 349 -1134
rect 506 -1206 507 -1134
rect 509 -1135 510 -1133
rect 702 -1135 703 -1133
rect 716 -1135 717 -1133
rect 772 -1206 773 -1134
rect 793 -1135 794 -1133
rect 800 -1206 801 -1134
rect 9 -1206 10 -1136
rect 282 -1137 283 -1133
rect 310 -1137 311 -1133
rect 320 -1206 321 -1136
rect 355 -1137 356 -1133
rect 373 -1137 374 -1133
rect 422 -1206 423 -1136
rect 593 -1206 594 -1136
rect 646 -1137 647 -1133
rect 688 -1206 689 -1136
rect 740 -1137 741 -1133
rect 793 -1206 794 -1136
rect 23 -1206 24 -1138
rect 338 -1139 339 -1133
rect 366 -1139 367 -1133
rect 548 -1139 549 -1133
rect 555 -1139 556 -1133
rect 765 -1206 766 -1138
rect 26 -1141 27 -1133
rect 639 -1141 640 -1133
rect 744 -1206 745 -1140
rect 779 -1141 780 -1133
rect 30 -1206 31 -1142
rect 597 -1143 598 -1133
rect 723 -1143 724 -1133
rect 779 -1206 780 -1142
rect 37 -1145 38 -1133
rect 187 -1145 188 -1133
rect 194 -1145 195 -1133
rect 331 -1145 332 -1133
rect 341 -1206 342 -1144
rect 597 -1206 598 -1144
rect 674 -1145 675 -1133
rect 723 -1206 724 -1144
rect 751 -1145 752 -1133
rect 758 -1145 759 -1133
rect 44 -1147 45 -1133
rect 338 -1206 339 -1146
rect 373 -1206 374 -1146
rect 513 -1147 514 -1133
rect 520 -1147 521 -1133
rect 702 -1206 703 -1146
rect 44 -1206 45 -1148
rect 429 -1149 430 -1133
rect 432 -1149 433 -1133
rect 716 -1206 717 -1148
rect 54 -1206 55 -1150
rect 457 -1151 458 -1133
rect 467 -1206 468 -1150
rect 492 -1151 493 -1133
rect 534 -1151 535 -1133
rect 611 -1206 612 -1150
rect 632 -1151 633 -1133
rect 751 -1206 752 -1150
rect 72 -1153 73 -1133
rect 247 -1153 248 -1133
rect 254 -1153 255 -1133
rect 310 -1206 311 -1152
rect 324 -1153 325 -1133
rect 366 -1206 367 -1152
rect 394 -1153 395 -1133
rect 674 -1206 675 -1152
rect 695 -1153 696 -1133
rect 758 -1206 759 -1152
rect 79 -1155 80 -1133
rect 324 -1206 325 -1154
rect 331 -1206 332 -1154
rect 380 -1155 381 -1133
rect 397 -1206 398 -1154
rect 555 -1206 556 -1154
rect 562 -1155 563 -1133
rect 632 -1206 633 -1154
rect 79 -1206 80 -1156
rect 142 -1157 143 -1133
rect 145 -1206 146 -1156
rect 208 -1157 209 -1133
rect 212 -1157 213 -1133
rect 236 -1206 237 -1156
rect 247 -1206 248 -1156
rect 257 -1206 258 -1156
rect 275 -1157 276 -1133
rect 436 -1206 437 -1156
rect 443 -1157 444 -1133
rect 562 -1206 563 -1156
rect 569 -1157 570 -1133
rect 747 -1157 748 -1133
rect 16 -1159 17 -1133
rect 275 -1206 276 -1158
rect 292 -1159 293 -1133
rect 380 -1206 381 -1158
rect 401 -1159 402 -1133
rect 492 -1206 493 -1158
rect 541 -1159 542 -1133
rect 618 -1206 619 -1158
rect 16 -1206 17 -1160
rect 163 -1161 164 -1133
rect 166 -1206 167 -1160
rect 180 -1161 181 -1133
rect 187 -1206 188 -1160
rect 457 -1206 458 -1160
rect 474 -1161 475 -1133
rect 527 -1161 528 -1133
rect 548 -1206 549 -1160
rect 786 -1161 787 -1133
rect 100 -1163 101 -1133
rect 513 -1206 514 -1162
rect 569 -1206 570 -1162
rect 814 -1163 815 -1133
rect 93 -1165 94 -1133
rect 100 -1206 101 -1164
rect 107 -1165 108 -1133
rect 107 -1206 108 -1164
rect 107 -1165 108 -1133
rect 107 -1206 108 -1164
rect 114 -1165 115 -1133
rect 681 -1165 682 -1133
rect 730 -1165 731 -1133
rect 786 -1206 787 -1164
rect 93 -1206 94 -1166
rect 390 -1206 391 -1166
rect 408 -1167 409 -1133
rect 534 -1206 535 -1166
rect 576 -1167 577 -1133
rect 639 -1206 640 -1166
rect 653 -1167 654 -1133
rect 730 -1206 731 -1166
rect 117 -1169 118 -1133
rect 282 -1206 283 -1168
rect 352 -1169 353 -1133
rect 695 -1206 696 -1168
rect 117 -1206 118 -1170
rect 191 -1206 192 -1170
rect 198 -1171 199 -1133
rect 289 -1206 290 -1170
rect 296 -1171 297 -1133
rect 352 -1206 353 -1170
rect 359 -1171 360 -1133
rect 443 -1206 444 -1170
rect 450 -1171 451 -1133
rect 520 -1206 521 -1170
rect 590 -1171 591 -1133
rect 646 -1206 647 -1170
rect 121 -1173 122 -1133
rect 149 -1206 150 -1172
rect 152 -1173 153 -1133
rect 583 -1173 584 -1133
rect 625 -1173 626 -1133
rect 681 -1206 682 -1172
rect 121 -1206 122 -1174
rect 128 -1175 129 -1133
rect 135 -1175 136 -1133
rect 583 -1206 584 -1174
rect 625 -1206 626 -1174
rect 660 -1175 661 -1133
rect 51 -1177 52 -1133
rect 128 -1206 129 -1176
rect 138 -1177 139 -1133
rect 317 -1177 318 -1133
rect 429 -1206 430 -1176
rect 471 -1177 472 -1133
rect 485 -1177 486 -1133
rect 653 -1206 654 -1176
rect 33 -1206 34 -1178
rect 485 -1206 486 -1178
rect 499 -1179 500 -1133
rect 576 -1206 577 -1178
rect 51 -1206 52 -1180
rect 737 -1181 738 -1133
rect 58 -1183 59 -1133
rect 135 -1206 136 -1182
rect 156 -1183 157 -1133
rect 156 -1206 157 -1182
rect 156 -1183 157 -1133
rect 156 -1206 157 -1182
rect 170 -1183 171 -1133
rect 170 -1206 171 -1182
rect 170 -1183 171 -1133
rect 170 -1206 171 -1182
rect 177 -1206 178 -1182
rect 369 -1183 370 -1133
rect 415 -1183 416 -1133
rect 499 -1206 500 -1182
rect 58 -1206 59 -1184
rect 68 -1206 69 -1184
rect 198 -1206 199 -1184
rect 261 -1185 262 -1133
rect 296 -1206 297 -1184
rect 425 -1185 426 -1133
rect 450 -1206 451 -1184
rect 478 -1185 479 -1133
rect 65 -1187 66 -1133
rect 415 -1206 416 -1186
rect 464 -1187 465 -1133
rect 527 -1206 528 -1186
rect 65 -1206 66 -1188
rect 72 -1206 73 -1188
rect 205 -1206 206 -1188
rect 394 -1206 395 -1188
rect 471 -1206 472 -1188
rect 604 -1189 605 -1133
rect 212 -1206 213 -1190
rect 240 -1191 241 -1133
rect 250 -1191 251 -1133
rect 604 -1206 605 -1190
rect 226 -1193 227 -1133
rect 233 -1193 234 -1133
rect 240 -1206 241 -1192
rect 404 -1206 405 -1192
rect 219 -1195 220 -1133
rect 226 -1206 227 -1194
rect 261 -1206 262 -1194
rect 268 -1195 269 -1133
rect 303 -1195 304 -1133
rect 359 -1206 360 -1194
rect 369 -1206 370 -1194
rect 387 -1195 388 -1133
rect 40 -1206 41 -1196
rect 219 -1206 220 -1196
rect 268 -1206 269 -1196
rect 411 -1206 412 -1196
rect 303 -1206 304 -1198
rect 345 -1199 346 -1133
rect 345 -1206 346 -1200
rect 667 -1201 668 -1133
rect 667 -1206 668 -1202
rect 709 -1203 710 -1133
rect 478 -1206 479 -1204
rect 709 -1206 710 -1204
rect 2 -1299 3 -1215
rect 135 -1216 136 -1214
rect 149 -1216 150 -1214
rect 149 -1299 150 -1215
rect 149 -1216 150 -1214
rect 149 -1299 150 -1215
rect 156 -1216 157 -1214
rect 156 -1299 157 -1215
rect 156 -1216 157 -1214
rect 156 -1299 157 -1215
rect 184 -1216 185 -1214
rect 198 -1216 199 -1214
rect 254 -1216 255 -1214
rect 310 -1216 311 -1214
rect 317 -1216 318 -1214
rect 443 -1216 444 -1214
rect 471 -1299 472 -1215
rect 506 -1216 507 -1214
rect 541 -1216 542 -1214
rect 646 -1216 647 -1214
rect 649 -1299 650 -1215
rect 786 -1216 787 -1214
rect 789 -1299 790 -1215
rect 800 -1216 801 -1214
rect 9 -1218 10 -1214
rect 348 -1218 349 -1214
rect 362 -1299 363 -1217
rect 597 -1218 598 -1214
rect 660 -1299 661 -1217
rect 786 -1299 787 -1217
rect 9 -1299 10 -1219
rect 30 -1220 31 -1214
rect 33 -1220 34 -1214
rect 663 -1220 664 -1214
rect 667 -1220 668 -1214
rect 737 -1299 738 -1219
rect 16 -1222 17 -1214
rect 89 -1222 90 -1214
rect 100 -1222 101 -1214
rect 100 -1299 101 -1221
rect 100 -1222 101 -1214
rect 100 -1299 101 -1221
rect 128 -1222 129 -1214
rect 394 -1299 395 -1221
rect 397 -1222 398 -1214
rect 520 -1222 521 -1214
rect 593 -1222 594 -1214
rect 730 -1222 731 -1214
rect 16 -1299 17 -1223
rect 145 -1224 146 -1214
rect 198 -1299 199 -1223
rect 380 -1224 381 -1214
rect 387 -1299 388 -1223
rect 534 -1224 535 -1214
rect 681 -1224 682 -1214
rect 730 -1299 731 -1223
rect 30 -1299 31 -1225
rect 187 -1299 188 -1225
rect 254 -1299 255 -1225
rect 327 -1226 328 -1214
rect 345 -1226 346 -1214
rect 485 -1226 486 -1214
rect 506 -1299 507 -1225
rect 611 -1226 612 -1214
rect 37 -1299 38 -1227
rect 268 -1228 269 -1214
rect 278 -1228 279 -1214
rect 590 -1299 591 -1227
rect 23 -1230 24 -1214
rect 268 -1299 269 -1229
rect 282 -1230 283 -1214
rect 345 -1299 346 -1229
rect 366 -1230 367 -1214
rect 499 -1230 500 -1214
rect 520 -1299 521 -1229
rect 576 -1230 577 -1214
rect 23 -1299 24 -1231
rect 219 -1232 220 -1214
rect 247 -1232 248 -1214
rect 499 -1299 500 -1231
rect 555 -1232 556 -1214
rect 681 -1299 682 -1231
rect 51 -1234 52 -1214
rect 58 -1234 59 -1214
rect 68 -1234 69 -1214
rect 72 -1234 73 -1214
rect 75 -1299 76 -1233
rect 436 -1234 437 -1214
rect 443 -1299 444 -1233
rect 492 -1234 493 -1214
rect 555 -1299 556 -1233
rect 653 -1234 654 -1214
rect 51 -1299 52 -1235
rect 121 -1236 122 -1214
rect 128 -1299 129 -1235
rect 338 -1299 339 -1235
rect 373 -1236 374 -1214
rect 541 -1299 542 -1235
rect 576 -1299 577 -1235
rect 604 -1236 605 -1214
rect 653 -1299 654 -1235
rect 688 -1236 689 -1214
rect 54 -1238 55 -1214
rect 492 -1299 493 -1237
rect 688 -1299 689 -1237
rect 758 -1238 759 -1214
rect 58 -1299 59 -1239
rect 240 -1240 241 -1214
rect 247 -1299 248 -1239
rect 289 -1240 290 -1214
rect 317 -1299 318 -1239
rect 422 -1240 423 -1214
rect 464 -1240 465 -1214
rect 597 -1299 598 -1239
rect 758 -1299 759 -1239
rect 779 -1240 780 -1214
rect 79 -1242 80 -1214
rect 142 -1242 143 -1214
rect 145 -1299 146 -1241
rect 191 -1242 192 -1214
rect 212 -1242 213 -1214
rect 219 -1299 220 -1241
rect 240 -1299 241 -1241
rect 352 -1242 353 -1214
rect 373 -1299 374 -1241
rect 429 -1242 430 -1214
rect 464 -1299 465 -1241
rect 513 -1242 514 -1214
rect 79 -1299 80 -1243
rect 331 -1244 332 -1214
rect 334 -1299 335 -1243
rect 604 -1299 605 -1243
rect 86 -1299 87 -1245
rect 359 -1246 360 -1214
rect 390 -1246 391 -1214
rect 632 -1246 633 -1214
rect 93 -1248 94 -1214
rect 121 -1299 122 -1247
rect 135 -1299 136 -1247
rect 205 -1248 206 -1214
rect 212 -1299 213 -1247
rect 415 -1248 416 -1214
rect 422 -1299 423 -1247
rect 450 -1248 451 -1214
rect 478 -1248 479 -1214
rect 751 -1248 752 -1214
rect 93 -1299 94 -1249
rect 177 -1250 178 -1214
rect 184 -1299 185 -1249
rect 436 -1299 437 -1249
rect 450 -1299 451 -1249
rect 667 -1299 668 -1249
rect 44 -1252 45 -1214
rect 177 -1299 178 -1251
rect 191 -1299 192 -1251
rect 303 -1252 304 -1214
rect 324 -1252 325 -1214
rect 723 -1252 724 -1214
rect 44 -1299 45 -1253
rect 72 -1299 73 -1253
rect 107 -1254 108 -1214
rect 289 -1299 290 -1253
rect 324 -1299 325 -1253
rect 457 -1254 458 -1214
rect 478 -1299 479 -1253
rect 527 -1254 528 -1214
rect 632 -1299 633 -1253
rect 779 -1299 780 -1253
rect 107 -1299 108 -1255
rect 170 -1256 171 -1214
rect 205 -1299 206 -1255
rect 226 -1256 227 -1214
rect 282 -1299 283 -1255
rect 341 -1256 342 -1214
rect 401 -1256 402 -1214
rect 548 -1256 549 -1214
rect 723 -1299 724 -1255
rect 744 -1256 745 -1214
rect 65 -1299 66 -1257
rect 170 -1299 171 -1257
rect 341 -1299 342 -1257
rect 562 -1258 563 -1214
rect 744 -1299 745 -1257
rect 772 -1258 773 -1214
rect 114 -1260 115 -1214
rect 751 -1299 752 -1259
rect 772 -1299 773 -1259
rect 793 -1260 794 -1214
rect 166 -1299 167 -1261
rect 380 -1299 381 -1261
rect 401 -1299 402 -1261
rect 765 -1262 766 -1214
rect 310 -1299 311 -1263
rect 562 -1299 563 -1263
rect 404 -1266 405 -1214
rect 611 -1299 612 -1265
rect 404 -1299 405 -1267
rect 534 -1299 535 -1267
rect 548 -1299 549 -1267
rect 618 -1268 619 -1214
rect 411 -1270 412 -1214
rect 639 -1270 640 -1214
rect 411 -1299 412 -1271
rect 702 -1272 703 -1214
rect 429 -1299 430 -1273
rect 583 -1274 584 -1214
rect 639 -1299 640 -1273
rect 695 -1274 696 -1214
rect 702 -1299 703 -1273
rect 716 -1274 717 -1214
rect 457 -1299 458 -1275
rect 485 -1299 486 -1275
rect 513 -1299 514 -1275
rect 572 -1299 573 -1275
rect 646 -1299 647 -1275
rect 716 -1299 717 -1275
rect 474 -1278 475 -1214
rect 583 -1299 584 -1277
rect 695 -1299 696 -1277
rect 709 -1278 710 -1214
rect 303 -1299 304 -1279
rect 709 -1299 710 -1279
rect 481 -1282 482 -1214
rect 782 -1299 783 -1281
rect 527 -1299 528 -1283
rect 674 -1284 675 -1214
rect 569 -1286 570 -1214
rect 618 -1299 619 -1285
rect 625 -1286 626 -1214
rect 674 -1299 675 -1285
rect 275 -1288 276 -1214
rect 625 -1299 626 -1287
rect 233 -1290 234 -1214
rect 275 -1299 276 -1289
rect 233 -1299 234 -1291
rect 261 -1292 262 -1214
rect 261 -1299 262 -1293
rect 296 -1294 297 -1214
rect 296 -1299 297 -1295
rect 408 -1296 409 -1214
rect 408 -1299 409 -1297
rect 415 -1299 416 -1297
rect 2 -1309 3 -1307
rect 348 -1376 349 -1308
rect 355 -1309 356 -1307
rect 751 -1309 752 -1307
rect 782 -1309 783 -1307
rect 800 -1376 801 -1308
rect 9 -1311 10 -1307
rect 180 -1376 181 -1310
rect 191 -1311 192 -1307
rect 313 -1311 314 -1307
rect 359 -1311 360 -1307
rect 499 -1311 500 -1307
rect 516 -1376 517 -1310
rect 674 -1311 675 -1307
rect 709 -1311 710 -1307
rect 768 -1311 769 -1307
rect 9 -1376 10 -1312
rect 320 -1376 321 -1312
rect 362 -1313 363 -1307
rect 562 -1313 563 -1307
rect 565 -1376 566 -1312
rect 705 -1376 706 -1312
rect 730 -1313 731 -1307
rect 779 -1376 780 -1312
rect 30 -1315 31 -1307
rect 33 -1365 34 -1314
rect 40 -1376 41 -1314
rect 44 -1315 45 -1307
rect 65 -1315 66 -1307
rect 527 -1315 528 -1307
rect 537 -1315 538 -1307
rect 737 -1315 738 -1307
rect 30 -1376 31 -1316
rect 128 -1317 129 -1307
rect 149 -1317 150 -1307
rect 187 -1317 188 -1307
rect 198 -1317 199 -1307
rect 352 -1317 353 -1307
rect 404 -1376 405 -1316
rect 492 -1317 493 -1307
rect 527 -1376 528 -1316
rect 555 -1317 556 -1307
rect 562 -1376 563 -1316
rect 695 -1317 696 -1307
rect 44 -1376 45 -1318
rect 464 -1319 465 -1307
rect 492 -1376 493 -1318
rect 583 -1319 584 -1307
rect 590 -1319 591 -1307
rect 709 -1376 710 -1318
rect 51 -1321 52 -1307
rect 187 -1376 188 -1320
rect 198 -1376 199 -1320
rect 205 -1321 206 -1307
rect 215 -1376 216 -1320
rect 359 -1376 360 -1320
rect 408 -1321 409 -1307
rect 702 -1321 703 -1307
rect 51 -1376 52 -1322
rect 145 -1376 146 -1322
rect 149 -1376 150 -1322
rect 156 -1323 157 -1307
rect 163 -1323 164 -1307
rect 289 -1323 290 -1307
rect 296 -1323 297 -1307
rect 366 -1323 367 -1307
rect 457 -1323 458 -1307
rect 520 -1323 521 -1307
rect 534 -1323 535 -1307
rect 590 -1376 591 -1322
rect 632 -1323 633 -1307
rect 632 -1376 633 -1322
rect 632 -1323 633 -1307
rect 632 -1376 633 -1322
rect 639 -1323 640 -1307
rect 691 -1376 692 -1322
rect 702 -1376 703 -1322
rect 723 -1323 724 -1307
rect 68 -1325 69 -1307
rect 93 -1325 94 -1307
rect 100 -1325 101 -1307
rect 100 -1376 101 -1324
rect 100 -1325 101 -1307
rect 100 -1376 101 -1324
rect 114 -1325 115 -1307
rect 201 -1325 202 -1307
rect 219 -1325 220 -1307
rect 229 -1325 230 -1307
rect 268 -1325 269 -1307
rect 289 -1376 290 -1324
rect 310 -1376 311 -1324
rect 394 -1325 395 -1307
rect 429 -1325 430 -1307
rect 534 -1376 535 -1324
rect 541 -1325 542 -1307
rect 555 -1376 556 -1324
rect 572 -1325 573 -1307
rect 758 -1325 759 -1307
rect 58 -1327 59 -1307
rect 219 -1376 220 -1326
rect 226 -1376 227 -1326
rect 247 -1327 248 -1307
rect 275 -1327 276 -1307
rect 408 -1376 409 -1326
rect 457 -1376 458 -1326
rect 478 -1327 479 -1307
rect 485 -1327 486 -1307
rect 520 -1376 521 -1326
rect 541 -1376 542 -1326
rect 548 -1327 549 -1307
rect 576 -1327 577 -1307
rect 583 -1376 584 -1326
rect 639 -1376 640 -1326
rect 653 -1327 654 -1307
rect 688 -1327 689 -1307
rect 695 -1376 696 -1326
rect 744 -1327 745 -1307
rect 758 -1376 759 -1326
rect 23 -1329 24 -1307
rect 275 -1376 276 -1328
rect 296 -1376 297 -1328
rect 576 -1376 577 -1328
rect 653 -1376 654 -1328
rect 667 -1329 668 -1307
rect 23 -1376 24 -1330
rect 415 -1331 416 -1307
rect 425 -1331 426 -1307
rect 667 -1376 668 -1330
rect 65 -1376 66 -1332
rect 93 -1376 94 -1332
rect 114 -1376 115 -1332
rect 282 -1333 283 -1307
rect 345 -1333 346 -1307
rect 415 -1376 416 -1332
rect 471 -1333 472 -1307
rect 485 -1376 486 -1332
rect 506 -1333 507 -1307
rect 548 -1376 549 -1332
rect 72 -1376 73 -1334
rect 646 -1376 647 -1334
rect 75 -1337 76 -1307
rect 429 -1376 430 -1336
rect 506 -1376 507 -1336
rect 513 -1337 514 -1307
rect 82 -1376 83 -1338
rect 107 -1339 108 -1307
rect 117 -1339 118 -1307
rect 499 -1376 500 -1338
rect 107 -1376 108 -1340
rect 184 -1341 185 -1307
rect 191 -1376 192 -1340
rect 688 -1376 689 -1340
rect 117 -1376 118 -1342
rect 142 -1343 143 -1307
rect 156 -1376 157 -1342
rect 170 -1343 171 -1307
rect 177 -1343 178 -1307
rect 247 -1376 248 -1342
rect 268 -1376 269 -1342
rect 478 -1376 479 -1342
rect 16 -1345 17 -1307
rect 170 -1376 171 -1344
rect 184 -1376 185 -1344
rect 338 -1376 339 -1344
rect 352 -1376 353 -1344
rect 373 -1345 374 -1307
rect 380 -1345 381 -1307
rect 394 -1376 395 -1344
rect 464 -1376 465 -1344
rect 513 -1376 514 -1344
rect 37 -1347 38 -1307
rect 142 -1376 143 -1346
rect 163 -1376 164 -1346
rect 436 -1347 437 -1307
rect 58 -1376 59 -1348
rect 177 -1376 178 -1348
rect 233 -1349 234 -1307
rect 282 -1376 283 -1348
rect 366 -1376 367 -1348
rect 446 -1376 447 -1348
rect 86 -1351 87 -1307
rect 233 -1376 234 -1350
rect 373 -1376 374 -1350
rect 450 -1351 451 -1307
rect 121 -1353 122 -1307
rect 128 -1376 129 -1352
rect 135 -1353 136 -1307
rect 205 -1376 206 -1352
rect 380 -1376 381 -1352
rect 597 -1353 598 -1307
rect 121 -1376 122 -1354
rect 254 -1355 255 -1307
rect 387 -1355 388 -1307
rect 471 -1376 472 -1354
rect 597 -1376 598 -1354
rect 611 -1355 612 -1307
rect 135 -1376 136 -1356
rect 334 -1357 335 -1307
rect 387 -1376 388 -1356
rect 401 -1357 402 -1307
rect 422 -1357 423 -1307
rect 436 -1376 437 -1356
rect 443 -1357 444 -1307
rect 450 -1376 451 -1356
rect 611 -1376 612 -1356
rect 625 -1357 626 -1307
rect 166 -1359 167 -1307
rect 481 -1376 482 -1358
rect 254 -1376 255 -1360
rect 317 -1361 318 -1307
rect 401 -1376 402 -1360
rect 674 -1376 675 -1360
rect 212 -1363 213 -1307
rect 317 -1376 318 -1362
rect 443 -1376 444 -1362
rect 618 -1363 619 -1307
rect 212 -1376 213 -1364
rect 261 -1365 262 -1307
rect 334 -1376 335 -1364
rect 618 -1376 619 -1364
rect 660 -1365 661 -1307
rect 79 -1367 80 -1307
rect 261 -1376 262 -1366
rect 303 -1367 304 -1307
rect 422 -1376 423 -1366
rect 660 -1376 661 -1366
rect 681 -1367 682 -1307
rect 79 -1376 80 -1368
rect 604 -1369 605 -1307
rect 681 -1376 682 -1368
rect 716 -1369 717 -1307
rect 303 -1376 304 -1370
rect 324 -1371 325 -1307
rect 331 -1376 332 -1370
rect 604 -1376 605 -1370
rect 240 -1373 241 -1307
rect 324 -1376 325 -1372
rect 240 -1376 241 -1374
rect 411 -1375 412 -1307
rect 9 -1445 10 -1385
rect 142 -1386 143 -1384
rect 149 -1386 150 -1384
rect 163 -1386 164 -1384
rect 170 -1386 171 -1384
rect 212 -1445 213 -1385
rect 271 -1445 272 -1385
rect 324 -1386 325 -1384
rect 338 -1386 339 -1384
rect 345 -1445 346 -1385
rect 383 -1445 384 -1385
rect 744 -1445 745 -1385
rect 758 -1386 759 -1384
rect 782 -1445 783 -1385
rect 786 -1445 787 -1385
rect 828 -1445 829 -1385
rect 16 -1445 17 -1387
rect 180 -1388 181 -1384
rect 275 -1388 276 -1384
rect 380 -1388 381 -1384
rect 411 -1388 412 -1384
rect 737 -1445 738 -1387
rect 779 -1388 780 -1384
rect 807 -1445 808 -1387
rect 37 -1445 38 -1389
rect 135 -1390 136 -1384
rect 149 -1445 150 -1389
rect 278 -1390 279 -1384
rect 296 -1390 297 -1384
rect 429 -1390 430 -1384
rect 443 -1390 444 -1384
rect 653 -1390 654 -1384
rect 674 -1390 675 -1384
rect 730 -1445 731 -1389
rect 789 -1445 790 -1389
rect 800 -1390 801 -1384
rect 44 -1392 45 -1384
rect 215 -1392 216 -1384
rect 247 -1392 248 -1384
rect 296 -1445 297 -1391
rect 310 -1392 311 -1384
rect 331 -1392 332 -1384
rect 338 -1445 339 -1391
rect 408 -1392 409 -1384
rect 443 -1445 444 -1391
rect 509 -1445 510 -1391
rect 534 -1392 535 -1384
rect 688 -1392 689 -1384
rect 695 -1392 696 -1384
rect 772 -1445 773 -1391
rect 796 -1445 797 -1391
rect 803 -1445 804 -1391
rect 44 -1445 45 -1393
rect 107 -1394 108 -1384
rect 121 -1394 122 -1384
rect 142 -1445 143 -1393
rect 156 -1394 157 -1384
rect 170 -1445 171 -1393
rect 177 -1394 178 -1384
rect 422 -1394 423 -1384
rect 457 -1394 458 -1384
rect 835 -1445 836 -1393
rect 51 -1396 52 -1384
rect 138 -1445 139 -1395
rect 163 -1445 164 -1395
rect 184 -1396 185 -1384
rect 226 -1396 227 -1384
rect 310 -1445 311 -1395
rect 324 -1445 325 -1395
rect 352 -1396 353 -1384
rect 394 -1396 395 -1384
rect 422 -1445 423 -1395
rect 450 -1396 451 -1384
rect 457 -1445 458 -1395
rect 464 -1396 465 -1384
rect 464 -1445 465 -1395
rect 464 -1396 465 -1384
rect 464 -1445 465 -1395
rect 478 -1396 479 -1384
rect 583 -1396 584 -1384
rect 590 -1396 591 -1384
rect 702 -1445 703 -1395
rect 709 -1396 710 -1384
rect 751 -1445 752 -1395
rect 51 -1445 52 -1397
rect 387 -1398 388 -1384
rect 394 -1445 395 -1397
rect 415 -1398 416 -1384
rect 488 -1445 489 -1397
rect 527 -1398 528 -1384
rect 551 -1445 552 -1397
rect 660 -1398 661 -1384
rect 674 -1445 675 -1397
rect 681 -1398 682 -1384
rect 58 -1400 59 -1384
rect 61 -1404 62 -1399
rect 75 -1400 76 -1384
rect 166 -1400 167 -1384
rect 226 -1445 227 -1399
rect 380 -1445 381 -1399
rect 404 -1400 405 -1384
rect 709 -1445 710 -1399
rect 58 -1445 59 -1401
rect 65 -1402 66 -1384
rect 75 -1445 76 -1401
rect 205 -1402 206 -1384
rect 254 -1402 255 -1384
rect 275 -1445 276 -1401
rect 303 -1402 304 -1384
rect 387 -1445 388 -1401
rect 404 -1445 405 -1401
rect 695 -1445 696 -1401
rect 65 -1445 66 -1403
rect 79 -1404 80 -1384
rect 177 -1445 178 -1403
rect 205 -1445 206 -1403
rect 299 -1404 300 -1384
rect 348 -1404 349 -1384
rect 534 -1445 535 -1403
rect 555 -1404 556 -1384
rect 716 -1404 717 -1384
rect 79 -1445 80 -1405
rect 128 -1406 129 -1384
rect 261 -1406 262 -1384
rect 303 -1445 304 -1405
rect 317 -1406 318 -1384
rect 716 -1445 717 -1405
rect 86 -1445 87 -1407
rect 100 -1408 101 -1384
rect 117 -1408 118 -1384
rect 478 -1445 479 -1407
rect 506 -1408 507 -1384
rect 625 -1445 626 -1407
rect 639 -1408 640 -1384
rect 688 -1445 689 -1407
rect 89 -1410 90 -1384
rect 247 -1445 248 -1409
rect 261 -1445 262 -1409
rect 268 -1410 269 -1384
rect 282 -1410 283 -1384
rect 317 -1445 318 -1409
rect 352 -1445 353 -1409
rect 516 -1410 517 -1384
rect 520 -1410 521 -1384
rect 590 -1445 591 -1409
rect 618 -1410 619 -1384
rect 653 -1445 654 -1409
rect 93 -1412 94 -1384
rect 611 -1412 612 -1384
rect 646 -1412 647 -1384
rect 723 -1445 724 -1411
rect 30 -1414 31 -1384
rect 93 -1445 94 -1413
rect 100 -1445 101 -1413
rect 240 -1414 241 -1384
rect 359 -1414 360 -1384
rect 450 -1445 451 -1413
rect 506 -1445 507 -1413
rect 611 -1445 612 -1413
rect 23 -1416 24 -1384
rect 30 -1445 31 -1415
rect 107 -1445 108 -1415
rect 117 -1445 118 -1415
rect 128 -1445 129 -1415
rect 198 -1416 199 -1384
rect 219 -1416 220 -1384
rect 282 -1445 283 -1415
rect 359 -1445 360 -1415
rect 373 -1416 374 -1384
rect 411 -1445 412 -1415
rect 415 -1445 416 -1415
rect 432 -1445 433 -1415
rect 555 -1445 556 -1415
rect 562 -1445 563 -1415
rect 632 -1416 633 -1384
rect 23 -1445 24 -1417
rect 471 -1418 472 -1384
rect 492 -1418 493 -1384
rect 632 -1445 633 -1417
rect 198 -1445 199 -1419
rect 289 -1420 290 -1384
rect 366 -1420 367 -1384
rect 492 -1445 493 -1419
rect 513 -1420 514 -1384
rect 618 -1445 619 -1419
rect 219 -1445 220 -1421
rect 429 -1445 430 -1421
rect 439 -1445 440 -1421
rect 513 -1445 514 -1421
rect 520 -1445 521 -1421
rect 691 -1422 692 -1384
rect 233 -1424 234 -1384
rect 289 -1445 290 -1423
rect 334 -1445 335 -1423
rect 366 -1445 367 -1423
rect 527 -1445 528 -1423
rect 548 -1424 549 -1384
rect 565 -1424 566 -1384
rect 660 -1445 661 -1423
rect 191 -1426 192 -1384
rect 233 -1445 234 -1425
rect 240 -1445 241 -1425
rect 254 -1445 255 -1425
rect 268 -1445 269 -1425
rect 373 -1445 374 -1425
rect 541 -1426 542 -1384
rect 639 -1445 640 -1425
rect 191 -1445 192 -1427
rect 765 -1445 766 -1427
rect 541 -1445 542 -1429
rect 705 -1430 706 -1384
rect 548 -1445 549 -1431
rect 681 -1445 682 -1431
rect 572 -1434 573 -1384
rect 667 -1434 668 -1384
rect 576 -1436 577 -1384
rect 576 -1445 577 -1435
rect 576 -1436 577 -1384
rect 576 -1445 577 -1435
rect 583 -1445 584 -1435
rect 604 -1436 605 -1384
rect 667 -1445 668 -1435
rect 768 -1445 769 -1435
rect 485 -1438 486 -1384
rect 604 -1445 605 -1437
rect 485 -1445 486 -1439
rect 569 -1445 570 -1439
rect 597 -1440 598 -1384
rect 646 -1445 647 -1439
rect 499 -1442 500 -1384
rect 597 -1445 598 -1441
rect 436 -1444 437 -1384
rect 499 -1445 500 -1443
rect 9 -1455 10 -1453
rect 96 -1524 97 -1454
rect 128 -1455 129 -1453
rect 548 -1524 549 -1454
rect 681 -1455 682 -1453
rect 789 -1455 790 -1453
rect 800 -1455 801 -1453
rect 814 -1455 815 -1453
rect 817 -1455 818 -1453
rect 828 -1455 829 -1453
rect 9 -1524 10 -1456
rect 779 -1457 780 -1453
rect 16 -1459 17 -1453
rect 436 -1524 437 -1458
rect 439 -1459 440 -1453
rect 632 -1459 633 -1453
rect 681 -1524 682 -1458
rect 737 -1459 738 -1453
rect 768 -1459 769 -1453
rect 807 -1459 808 -1453
rect 16 -1524 17 -1460
rect 471 -1461 472 -1453
rect 474 -1461 475 -1453
rect 751 -1461 752 -1453
rect 23 -1463 24 -1453
rect 138 -1463 139 -1453
rect 156 -1463 157 -1453
rect 723 -1463 724 -1453
rect 737 -1524 738 -1462
rect 772 -1463 773 -1453
rect 23 -1524 24 -1464
rect 163 -1465 164 -1453
rect 198 -1465 199 -1453
rect 380 -1465 381 -1453
rect 394 -1524 395 -1464
rect 422 -1465 423 -1453
rect 429 -1465 430 -1453
rect 604 -1465 605 -1453
rect 632 -1524 633 -1464
rect 667 -1465 668 -1453
rect 674 -1465 675 -1453
rect 723 -1524 724 -1464
rect 30 -1467 31 -1453
rect 184 -1467 185 -1453
rect 250 -1524 251 -1466
rect 418 -1524 419 -1466
rect 422 -1524 423 -1466
rect 492 -1467 493 -1453
rect 509 -1467 510 -1453
rect 688 -1467 689 -1453
rect 30 -1524 31 -1468
rect 180 -1524 181 -1468
rect 257 -1524 258 -1468
rect 611 -1469 612 -1453
rect 667 -1524 668 -1468
rect 716 -1469 717 -1453
rect 37 -1471 38 -1453
rect 166 -1524 167 -1470
rect 268 -1524 269 -1470
rect 296 -1471 297 -1453
rect 303 -1471 304 -1453
rect 471 -1524 472 -1470
rect 523 -1524 524 -1470
rect 625 -1471 626 -1453
rect 688 -1524 689 -1470
rect 744 -1471 745 -1453
rect 44 -1473 45 -1453
rect 117 -1473 118 -1453
rect 128 -1524 129 -1472
rect 142 -1473 143 -1453
rect 159 -1473 160 -1453
rect 408 -1524 409 -1472
rect 432 -1473 433 -1453
rect 639 -1473 640 -1453
rect 54 -1524 55 -1474
rect 716 -1524 717 -1474
rect 58 -1477 59 -1453
rect 72 -1524 73 -1476
rect 79 -1477 80 -1453
rect 82 -1507 83 -1476
rect 114 -1524 115 -1476
rect 138 -1524 139 -1476
rect 142 -1524 143 -1476
rect 177 -1477 178 -1453
rect 296 -1524 297 -1476
rect 369 -1524 370 -1476
rect 383 -1477 384 -1453
rect 611 -1524 612 -1476
rect 37 -1524 38 -1478
rect 383 -1524 384 -1478
rect 401 -1479 402 -1453
rect 457 -1479 458 -1453
rect 527 -1479 528 -1453
rect 604 -1524 605 -1478
rect 44 -1524 45 -1480
rect 177 -1524 178 -1480
rect 212 -1481 213 -1453
rect 457 -1524 458 -1480
rect 464 -1481 465 -1453
rect 527 -1524 528 -1480
rect 534 -1481 535 -1453
rect 537 -1481 538 -1453
rect 541 -1481 542 -1453
rect 625 -1524 626 -1480
rect 58 -1524 59 -1482
rect 86 -1483 87 -1453
rect 135 -1483 136 -1453
rect 156 -1524 157 -1482
rect 212 -1524 213 -1482
rect 254 -1483 255 -1453
rect 306 -1524 307 -1482
rect 730 -1483 731 -1453
rect 65 -1485 66 -1453
rect 124 -1485 125 -1453
rect 331 -1485 332 -1453
rect 345 -1485 346 -1453
rect 352 -1485 353 -1453
rect 506 -1524 507 -1484
rect 513 -1485 514 -1453
rect 541 -1524 542 -1484
rect 555 -1485 556 -1453
rect 744 -1524 745 -1484
rect 65 -1524 66 -1486
rect 149 -1487 150 -1453
rect 289 -1487 290 -1453
rect 345 -1524 346 -1486
rect 359 -1487 360 -1453
rect 429 -1524 430 -1486
rect 439 -1524 440 -1486
rect 646 -1487 647 -1453
rect 79 -1524 80 -1488
rect 149 -1524 150 -1488
rect 219 -1489 220 -1453
rect 289 -1524 290 -1488
rect 373 -1489 374 -1453
rect 390 -1524 391 -1488
rect 464 -1524 465 -1488
rect 478 -1489 479 -1453
rect 513 -1524 514 -1488
rect 534 -1524 535 -1488
rect 618 -1489 619 -1453
rect 646 -1524 647 -1488
rect 835 -1489 836 -1453
rect 86 -1524 87 -1490
rect 275 -1491 276 -1453
rect 317 -1491 318 -1453
rect 352 -1524 353 -1490
rect 366 -1491 367 -1453
rect 492 -1524 493 -1490
rect 555 -1524 556 -1490
rect 583 -1491 584 -1453
rect 597 -1491 598 -1453
rect 751 -1524 752 -1490
rect 170 -1493 171 -1453
rect 219 -1524 220 -1492
rect 233 -1493 234 -1453
rect 275 -1524 276 -1492
rect 282 -1493 283 -1453
rect 317 -1524 318 -1492
rect 331 -1524 332 -1492
rect 576 -1493 577 -1453
rect 597 -1524 598 -1492
rect 730 -1524 731 -1492
rect 93 -1495 94 -1453
rect 170 -1524 171 -1494
rect 191 -1495 192 -1453
rect 373 -1524 374 -1494
rect 387 -1495 388 -1453
rect 478 -1524 479 -1494
rect 562 -1495 563 -1453
rect 674 -1524 675 -1494
rect 121 -1497 122 -1453
rect 191 -1524 192 -1496
rect 233 -1524 234 -1496
rect 271 -1497 272 -1453
rect 310 -1497 311 -1453
rect 387 -1524 388 -1496
rect 397 -1497 398 -1453
rect 576 -1524 577 -1496
rect 618 -1524 619 -1496
rect 653 -1497 654 -1453
rect 107 -1499 108 -1453
rect 121 -1524 122 -1498
rect 247 -1499 248 -1453
rect 310 -1524 311 -1498
rect 334 -1499 335 -1453
rect 660 -1499 661 -1453
rect 107 -1524 108 -1500
rect 187 -1501 188 -1453
rect 198 -1524 199 -1500
rect 247 -1524 248 -1500
rect 261 -1501 262 -1453
rect 282 -1524 283 -1500
rect 338 -1501 339 -1453
rect 401 -1524 402 -1500
rect 450 -1501 451 -1453
rect 639 -1524 640 -1500
rect 653 -1524 654 -1500
rect 695 -1501 696 -1453
rect 240 -1503 241 -1453
rect 261 -1524 262 -1502
rect 324 -1503 325 -1453
rect 338 -1524 339 -1502
rect 341 -1524 342 -1502
rect 583 -1524 584 -1502
rect 660 -1524 661 -1502
rect 702 -1503 703 -1453
rect 240 -1524 241 -1504
rect 404 -1505 405 -1453
rect 450 -1524 451 -1504
rect 499 -1505 500 -1453
rect 520 -1505 521 -1453
rect 562 -1524 563 -1504
rect 324 -1524 325 -1506
rect 443 -1507 444 -1453
rect 485 -1524 486 -1506
rect 520 -1524 521 -1506
rect 537 -1524 538 -1506
rect 695 -1524 696 -1506
rect 226 -1509 227 -1453
rect 443 -1524 444 -1508
rect 205 -1511 206 -1453
rect 226 -1524 227 -1510
rect 362 -1524 363 -1510
rect 702 -1524 703 -1510
rect 366 -1524 367 -1512
rect 709 -1513 710 -1453
rect 380 -1524 381 -1514
rect 709 -1524 710 -1514
rect 415 -1517 416 -1453
rect 499 -1524 500 -1516
rect 415 -1524 416 -1518
rect 590 -1519 591 -1453
rect 569 -1521 570 -1453
rect 590 -1524 591 -1520
rect 359 -1524 360 -1522
rect 569 -1524 570 -1522
rect 12 -1603 13 -1533
rect 16 -1534 17 -1532
rect 51 -1534 52 -1532
rect 205 -1534 206 -1532
rect 208 -1534 209 -1532
rect 261 -1534 262 -1532
rect 303 -1534 304 -1532
rect 317 -1534 318 -1532
rect 331 -1534 332 -1532
rect 436 -1603 437 -1533
rect 488 -1603 489 -1533
rect 744 -1534 745 -1532
rect 16 -1603 17 -1535
rect 212 -1536 213 -1532
rect 226 -1536 227 -1532
rect 226 -1603 227 -1535
rect 226 -1536 227 -1532
rect 226 -1603 227 -1535
rect 240 -1603 241 -1535
rect 324 -1536 325 -1532
rect 338 -1536 339 -1532
rect 471 -1536 472 -1532
rect 520 -1603 521 -1535
rect 604 -1536 605 -1532
rect 618 -1603 619 -1535
rect 667 -1536 668 -1532
rect 2 -1538 3 -1532
rect 324 -1603 325 -1537
rect 341 -1538 342 -1532
rect 667 -1603 668 -1537
rect 23 -1540 24 -1532
rect 205 -1603 206 -1539
rect 212 -1603 213 -1539
rect 289 -1540 290 -1532
rect 303 -1603 304 -1539
rect 639 -1540 640 -1532
rect 23 -1603 24 -1541
rect 345 -1542 346 -1532
rect 362 -1542 363 -1532
rect 443 -1542 444 -1532
rect 471 -1603 472 -1541
rect 702 -1542 703 -1532
rect 44 -1544 45 -1532
rect 331 -1603 332 -1543
rect 341 -1603 342 -1543
rect 499 -1544 500 -1532
rect 597 -1544 598 -1532
rect 737 -1544 738 -1532
rect 44 -1603 45 -1545
rect 569 -1546 570 -1532
rect 604 -1603 605 -1545
rect 653 -1546 654 -1532
rect 51 -1603 52 -1547
rect 128 -1548 129 -1532
rect 138 -1548 139 -1532
rect 478 -1548 479 -1532
rect 499 -1603 500 -1547
rect 751 -1548 752 -1532
rect 58 -1550 59 -1532
rect 96 -1550 97 -1532
rect 103 -1603 104 -1549
rect 191 -1550 192 -1532
rect 233 -1603 234 -1549
rect 478 -1603 479 -1549
rect 569 -1603 570 -1549
rect 632 -1550 633 -1532
rect 653 -1603 654 -1549
rect 709 -1550 710 -1532
rect 58 -1603 59 -1551
rect 170 -1552 171 -1532
rect 184 -1552 185 -1532
rect 275 -1552 276 -1532
rect 278 -1603 279 -1551
rect 597 -1603 598 -1551
rect 632 -1603 633 -1551
rect 688 -1552 689 -1532
rect 72 -1603 73 -1553
rect 100 -1554 101 -1532
rect 117 -1603 118 -1553
rect 121 -1554 122 -1532
rect 128 -1603 129 -1553
rect 320 -1603 321 -1553
rect 345 -1603 346 -1553
rect 541 -1554 542 -1532
rect 79 -1556 80 -1532
rect 89 -1603 90 -1555
rect 93 -1603 94 -1555
rect 114 -1556 115 -1532
rect 121 -1603 122 -1555
rect 296 -1556 297 -1532
rect 306 -1556 307 -1532
rect 457 -1556 458 -1532
rect 82 -1603 83 -1557
rect 254 -1603 255 -1557
rect 257 -1558 258 -1532
rect 548 -1558 549 -1532
rect 86 -1560 87 -1532
rect 268 -1603 269 -1559
rect 289 -1603 290 -1559
rect 408 -1560 409 -1532
rect 415 -1560 416 -1532
rect 646 -1560 647 -1532
rect 65 -1562 66 -1532
rect 408 -1603 409 -1561
rect 415 -1603 416 -1561
rect 422 -1562 423 -1532
rect 443 -1603 444 -1561
rect 534 -1562 535 -1532
rect 548 -1603 549 -1561
rect 600 -1562 601 -1532
rect 646 -1603 647 -1561
rect 695 -1562 696 -1532
rect 30 -1564 31 -1532
rect 65 -1603 66 -1563
rect 138 -1603 139 -1563
rect 219 -1564 220 -1532
rect 247 -1564 248 -1532
rect 401 -1564 402 -1532
rect 422 -1603 423 -1563
rect 506 -1564 507 -1532
rect 534 -1603 535 -1563
rect 611 -1564 612 -1532
rect 30 -1603 31 -1565
rect 583 -1566 584 -1532
rect 611 -1603 612 -1565
rect 660 -1566 661 -1532
rect 149 -1568 150 -1532
rect 163 -1603 164 -1567
rect 170 -1603 171 -1567
rect 236 -1603 237 -1567
rect 247 -1603 248 -1567
rect 282 -1568 283 -1532
rect 296 -1603 297 -1567
rect 513 -1568 514 -1532
rect 555 -1568 556 -1532
rect 583 -1603 584 -1567
rect 660 -1603 661 -1567
rect 716 -1568 717 -1532
rect 152 -1603 153 -1569
rect 352 -1570 353 -1532
rect 362 -1603 363 -1569
rect 541 -1603 542 -1569
rect 37 -1572 38 -1532
rect 352 -1603 353 -1571
rect 366 -1603 367 -1571
rect 492 -1572 493 -1532
rect 37 -1603 38 -1573
rect 107 -1574 108 -1532
rect 184 -1603 185 -1573
rect 198 -1574 199 -1532
rect 219 -1603 220 -1573
rect 639 -1603 640 -1573
rect 9 -1576 10 -1532
rect 107 -1603 108 -1575
rect 177 -1576 178 -1532
rect 198 -1603 199 -1575
rect 250 -1576 251 -1532
rect 373 -1576 374 -1532
rect 380 -1576 381 -1532
rect 450 -1576 451 -1532
rect 457 -1603 458 -1575
rect 576 -1576 577 -1532
rect 114 -1603 115 -1577
rect 380 -1603 381 -1577
rect 387 -1578 388 -1532
rect 674 -1578 675 -1532
rect 156 -1580 157 -1532
rect 177 -1603 178 -1579
rect 187 -1580 188 -1532
rect 191 -1603 192 -1579
rect 261 -1603 262 -1579
rect 310 -1580 311 -1532
rect 313 -1603 314 -1579
rect 429 -1580 430 -1532
rect 439 -1580 440 -1532
rect 506 -1603 507 -1579
rect 674 -1603 675 -1579
rect 723 -1580 724 -1532
rect 142 -1582 143 -1532
rect 156 -1603 157 -1581
rect 275 -1603 276 -1581
rect 373 -1603 374 -1581
rect 394 -1582 395 -1532
rect 394 -1603 395 -1581
rect 394 -1582 395 -1532
rect 394 -1603 395 -1581
rect 401 -1603 402 -1581
rect 527 -1582 528 -1532
rect 282 -1603 283 -1583
rect 310 -1603 311 -1583
rect 334 -1584 335 -1532
rect 513 -1603 514 -1583
rect 306 -1603 307 -1585
rect 527 -1603 528 -1585
rect 418 -1588 419 -1532
rect 450 -1603 451 -1587
rect 485 -1588 486 -1532
rect 576 -1603 577 -1587
rect 387 -1603 388 -1589
rect 485 -1603 486 -1589
rect 492 -1603 493 -1589
rect 590 -1590 591 -1532
rect 411 -1603 412 -1591
rect 590 -1603 591 -1591
rect 429 -1603 430 -1593
rect 464 -1594 465 -1532
rect 464 -1603 465 -1595
rect 562 -1596 563 -1532
rect 562 -1603 563 -1597
rect 625 -1598 626 -1532
rect 625 -1603 626 -1599
rect 681 -1600 682 -1532
rect 681 -1603 682 -1601
rect 730 -1602 731 -1532
rect 5 -1613 6 -1611
rect 324 -1613 325 -1611
rect 359 -1613 360 -1611
rect 471 -1613 472 -1611
rect 485 -1672 486 -1612
rect 520 -1613 521 -1611
rect 558 -1613 559 -1611
rect 646 -1613 647 -1611
rect 9 -1672 10 -1614
rect 156 -1615 157 -1611
rect 163 -1615 164 -1611
rect 163 -1672 164 -1614
rect 163 -1615 164 -1611
rect 163 -1672 164 -1614
rect 187 -1672 188 -1614
rect 198 -1615 199 -1611
rect 226 -1615 227 -1611
rect 278 -1615 279 -1611
rect 317 -1615 318 -1611
rect 499 -1615 500 -1611
rect 520 -1672 521 -1614
rect 576 -1615 577 -1611
rect 625 -1615 626 -1611
rect 649 -1672 650 -1614
rect 23 -1617 24 -1611
rect 79 -1672 80 -1616
rect 82 -1617 83 -1611
rect 639 -1617 640 -1611
rect 23 -1672 24 -1618
rect 110 -1672 111 -1618
rect 114 -1619 115 -1611
rect 299 -1672 300 -1618
rect 359 -1672 360 -1618
rect 534 -1619 535 -1611
rect 30 -1621 31 -1611
rect 324 -1672 325 -1620
rect 362 -1621 363 -1611
rect 394 -1621 395 -1611
rect 401 -1621 402 -1611
rect 408 -1621 409 -1611
rect 411 -1621 412 -1611
rect 632 -1621 633 -1611
rect 30 -1672 31 -1622
rect 219 -1623 220 -1611
rect 233 -1623 234 -1611
rect 247 -1623 248 -1611
rect 254 -1623 255 -1611
rect 317 -1672 318 -1622
rect 366 -1672 367 -1622
rect 464 -1623 465 -1611
rect 478 -1623 479 -1611
rect 499 -1672 500 -1622
rect 534 -1672 535 -1622
rect 604 -1623 605 -1611
rect 16 -1625 17 -1611
rect 464 -1672 465 -1624
rect 16 -1672 17 -1626
rect 138 -1627 139 -1611
rect 152 -1627 153 -1611
rect 254 -1672 255 -1626
rect 268 -1627 269 -1611
rect 310 -1672 311 -1626
rect 373 -1627 374 -1611
rect 478 -1672 479 -1626
rect 37 -1629 38 -1611
rect 100 -1672 101 -1628
rect 128 -1629 129 -1611
rect 156 -1672 157 -1628
rect 170 -1629 171 -1611
rect 226 -1672 227 -1628
rect 240 -1629 241 -1611
rect 268 -1672 269 -1628
rect 376 -1672 377 -1628
rect 387 -1629 388 -1611
rect 394 -1672 395 -1628
rect 506 -1629 507 -1611
rect 37 -1672 38 -1630
rect 306 -1631 307 -1611
rect 380 -1631 381 -1611
rect 471 -1672 472 -1630
rect 506 -1672 507 -1630
rect 611 -1631 612 -1611
rect 65 -1633 66 -1611
rect 275 -1633 276 -1611
rect 292 -1672 293 -1632
rect 611 -1672 612 -1632
rect 58 -1635 59 -1611
rect 65 -1672 66 -1634
rect 72 -1635 73 -1611
rect 142 -1635 143 -1611
rect 173 -1672 174 -1634
rect 198 -1672 199 -1634
rect 205 -1635 206 -1611
rect 247 -1672 248 -1634
rect 275 -1672 276 -1634
rect 352 -1635 353 -1611
rect 380 -1672 381 -1634
rect 429 -1635 430 -1611
rect 436 -1672 437 -1634
rect 457 -1635 458 -1611
rect 58 -1672 59 -1636
rect 191 -1637 192 -1611
rect 205 -1672 206 -1636
rect 369 -1672 370 -1636
rect 401 -1672 402 -1636
rect 422 -1637 423 -1611
rect 429 -1672 430 -1636
rect 450 -1637 451 -1611
rect 457 -1672 458 -1636
rect 555 -1637 556 -1611
rect 47 -1639 48 -1611
rect 191 -1672 192 -1638
rect 212 -1639 213 -1611
rect 233 -1672 234 -1638
rect 296 -1639 297 -1611
rect 387 -1672 388 -1638
rect 408 -1672 409 -1638
rect 660 -1639 661 -1611
rect 51 -1641 52 -1611
rect 422 -1672 423 -1640
rect 439 -1641 440 -1611
rect 590 -1641 591 -1611
rect 660 -1672 661 -1640
rect 674 -1641 675 -1611
rect 51 -1672 52 -1642
rect 338 -1643 339 -1611
rect 443 -1643 444 -1611
rect 597 -1643 598 -1611
rect 86 -1645 87 -1611
rect 149 -1672 150 -1644
rect 184 -1645 185 -1611
rect 219 -1672 220 -1644
rect 296 -1672 297 -1644
rect 576 -1672 577 -1644
rect 597 -1672 598 -1644
rect 681 -1645 682 -1611
rect 72 -1672 73 -1646
rect 86 -1672 87 -1646
rect 89 -1647 90 -1611
rect 653 -1647 654 -1611
rect 677 -1672 678 -1646
rect 681 -1672 682 -1646
rect 93 -1649 94 -1611
rect 117 -1672 118 -1648
rect 128 -1672 129 -1648
rect 177 -1649 178 -1611
rect 194 -1649 195 -1611
rect 590 -1672 591 -1648
rect 93 -1672 94 -1650
rect 121 -1651 122 -1611
rect 135 -1651 136 -1611
rect 177 -1672 178 -1650
rect 212 -1672 213 -1650
rect 261 -1651 262 -1611
rect 331 -1651 332 -1611
rect 338 -1672 339 -1650
rect 443 -1672 444 -1650
rect 513 -1651 514 -1611
rect 107 -1653 108 -1611
rect 135 -1672 136 -1652
rect 446 -1653 447 -1611
rect 555 -1672 556 -1652
rect 114 -1672 115 -1654
rect 170 -1672 171 -1654
rect 450 -1672 451 -1654
rect 541 -1655 542 -1611
rect 121 -1672 122 -1656
rect 289 -1657 290 -1611
rect 320 -1657 321 -1611
rect 541 -1672 542 -1656
rect 282 -1659 283 -1611
rect 289 -1672 290 -1658
rect 513 -1672 514 -1658
rect 562 -1659 563 -1611
rect 282 -1672 283 -1660
rect 415 -1661 416 -1611
rect 548 -1661 549 -1611
rect 562 -1672 563 -1660
rect 345 -1663 346 -1611
rect 415 -1672 416 -1662
rect 548 -1672 549 -1662
rect 569 -1663 570 -1611
rect 345 -1672 346 -1664
rect 492 -1665 493 -1611
rect 569 -1672 570 -1664
rect 618 -1665 619 -1611
rect 492 -1672 493 -1666
rect 527 -1667 528 -1611
rect 527 -1672 528 -1668
rect 583 -1669 584 -1611
rect 583 -1672 584 -1670
rect 667 -1671 668 -1611
rect 16 -1682 17 -1680
rect 86 -1682 87 -1680
rect 107 -1682 108 -1680
rect 159 -1729 160 -1681
rect 170 -1729 171 -1681
rect 177 -1682 178 -1680
rect 187 -1682 188 -1680
rect 422 -1682 423 -1680
rect 446 -1729 447 -1681
rect 492 -1682 493 -1680
rect 506 -1682 507 -1680
rect 653 -1729 654 -1681
rect 674 -1729 675 -1681
rect 681 -1682 682 -1680
rect 16 -1729 17 -1683
rect 93 -1684 94 -1680
rect 145 -1684 146 -1680
rect 296 -1684 297 -1680
rect 306 -1684 307 -1680
rect 471 -1684 472 -1680
rect 534 -1684 535 -1680
rect 579 -1729 580 -1683
rect 649 -1684 650 -1680
rect 660 -1684 661 -1680
rect 23 -1686 24 -1680
rect 142 -1686 143 -1680
rect 156 -1686 157 -1680
rect 191 -1729 192 -1685
rect 212 -1686 213 -1680
rect 261 -1686 262 -1680
rect 264 -1686 265 -1680
rect 464 -1686 465 -1680
rect 471 -1729 472 -1685
rect 513 -1686 514 -1680
rect 548 -1686 549 -1680
rect 621 -1686 622 -1680
rect 23 -1729 24 -1687
rect 345 -1688 346 -1680
rect 352 -1688 353 -1680
rect 590 -1688 591 -1680
rect 30 -1729 31 -1689
rect 226 -1690 227 -1680
rect 243 -1690 244 -1680
rect 324 -1690 325 -1680
rect 331 -1690 332 -1680
rect 541 -1690 542 -1680
rect 569 -1690 570 -1680
rect 618 -1690 619 -1680
rect 37 -1692 38 -1680
rect 313 -1729 314 -1691
rect 317 -1692 318 -1680
rect 359 -1692 360 -1680
rect 376 -1729 377 -1691
rect 499 -1692 500 -1680
rect 597 -1692 598 -1680
rect 618 -1729 619 -1691
rect 9 -1694 10 -1680
rect 317 -1729 318 -1693
rect 320 -1729 321 -1693
rect 408 -1694 409 -1680
rect 499 -1729 500 -1693
rect 527 -1694 528 -1680
rect 9 -1729 10 -1695
rect 128 -1696 129 -1680
rect 173 -1696 174 -1680
rect 334 -1696 335 -1680
rect 338 -1729 339 -1695
rect 576 -1696 577 -1680
rect 40 -1729 41 -1697
rect 198 -1698 199 -1680
rect 212 -1729 213 -1697
rect 275 -1698 276 -1680
rect 282 -1698 283 -1680
rect 355 -1698 356 -1680
rect 390 -1698 391 -1680
rect 443 -1698 444 -1680
rect 527 -1729 528 -1697
rect 611 -1698 612 -1680
rect 44 -1729 45 -1699
rect 131 -1729 132 -1699
rect 187 -1729 188 -1699
rect 236 -1700 237 -1680
rect 247 -1700 248 -1680
rect 289 -1700 290 -1680
rect 292 -1700 293 -1680
rect 296 -1729 297 -1699
rect 310 -1700 311 -1680
rect 359 -1729 360 -1699
rect 408 -1729 409 -1699
rect 436 -1700 437 -1680
rect 47 -1702 48 -1680
rect 58 -1702 59 -1680
rect 65 -1702 66 -1680
rect 261 -1729 262 -1701
rect 271 -1729 272 -1701
rect 464 -1729 465 -1701
rect 51 -1729 52 -1703
rect 257 -1729 258 -1703
rect 275 -1729 276 -1703
rect 394 -1704 395 -1680
rect 436 -1729 437 -1703
rect 450 -1704 451 -1680
rect 58 -1729 59 -1705
rect 520 -1706 521 -1680
rect 65 -1729 66 -1707
rect 128 -1729 129 -1707
rect 198 -1729 199 -1707
rect 233 -1708 234 -1680
rect 247 -1729 248 -1707
rect 373 -1708 374 -1680
rect 380 -1708 381 -1680
rect 394 -1729 395 -1707
rect 520 -1729 521 -1707
rect 562 -1708 563 -1680
rect 72 -1710 73 -1680
rect 124 -1729 125 -1709
rect 219 -1710 220 -1680
rect 226 -1729 227 -1709
rect 250 -1729 251 -1709
rect 492 -1729 493 -1709
rect 72 -1729 73 -1711
rect 205 -1712 206 -1680
rect 254 -1712 255 -1680
rect 324 -1729 325 -1711
rect 331 -1729 332 -1711
rect 415 -1712 416 -1680
rect 79 -1714 80 -1680
rect 289 -1729 290 -1713
rect 310 -1729 311 -1713
rect 478 -1714 479 -1680
rect 79 -1729 80 -1715
rect 268 -1716 269 -1680
rect 282 -1729 283 -1715
rect 429 -1716 430 -1680
rect 86 -1729 87 -1717
rect 114 -1718 115 -1680
rect 121 -1718 122 -1680
rect 233 -1729 234 -1717
rect 240 -1729 241 -1717
rect 478 -1729 479 -1717
rect 107 -1729 108 -1719
rect 142 -1729 143 -1719
rect 149 -1720 150 -1680
rect 219 -1729 220 -1719
rect 268 -1729 269 -1719
rect 366 -1729 367 -1719
rect 373 -1729 374 -1719
rect 422 -1729 423 -1719
rect 429 -1729 430 -1719
rect 485 -1720 486 -1680
rect 114 -1729 115 -1721
rect 135 -1722 136 -1680
rect 345 -1729 346 -1721
rect 401 -1722 402 -1680
rect 485 -1729 486 -1721
rect 555 -1722 556 -1680
rect 121 -1729 122 -1723
rect 380 -1729 381 -1723
rect 401 -1729 402 -1723
rect 457 -1724 458 -1680
rect 555 -1729 556 -1723
rect 583 -1724 584 -1680
rect 135 -1729 136 -1725
rect 163 -1726 164 -1680
rect 303 -1729 304 -1725
rect 457 -1729 458 -1725
rect 163 -1729 164 -1727
rect 184 -1729 185 -1727
rect 362 -1728 363 -1680
rect 415 -1729 416 -1727
rect 16 -1739 17 -1737
rect 152 -1739 153 -1737
rect 156 -1770 157 -1738
rect 240 -1770 241 -1738
rect 254 -1770 255 -1738
rect 257 -1739 258 -1737
rect 261 -1739 262 -1737
rect 352 -1739 353 -1737
rect 418 -1770 419 -1738
rect 534 -1770 535 -1738
rect 548 -1770 549 -1738
rect 555 -1739 556 -1737
rect 618 -1739 619 -1737
rect 618 -1770 619 -1738
rect 618 -1739 619 -1737
rect 618 -1770 619 -1738
rect 632 -1770 633 -1738
rect 653 -1739 654 -1737
rect 670 -1739 671 -1737
rect 674 -1739 675 -1737
rect 23 -1741 24 -1737
rect 362 -1741 363 -1737
rect 422 -1741 423 -1737
rect 453 -1770 454 -1740
rect 460 -1741 461 -1737
rect 520 -1741 521 -1737
rect 37 -1770 38 -1742
rect 107 -1743 108 -1737
rect 114 -1743 115 -1737
rect 177 -1743 178 -1737
rect 208 -1743 209 -1737
rect 296 -1743 297 -1737
rect 331 -1743 332 -1737
rect 352 -1770 353 -1742
rect 408 -1743 409 -1737
rect 460 -1770 461 -1742
rect 471 -1743 472 -1737
rect 513 -1770 514 -1742
rect 44 -1745 45 -1737
rect 310 -1745 311 -1737
rect 334 -1770 335 -1744
rect 492 -1745 493 -1737
rect 51 -1747 52 -1737
rect 292 -1747 293 -1737
rect 296 -1770 297 -1746
rect 366 -1747 367 -1737
rect 422 -1770 423 -1746
rect 478 -1747 479 -1737
rect 51 -1770 52 -1748
rect 135 -1749 136 -1737
rect 145 -1749 146 -1737
rect 219 -1749 220 -1737
rect 226 -1749 227 -1737
rect 243 -1749 244 -1737
rect 282 -1749 283 -1737
rect 317 -1770 318 -1748
rect 338 -1770 339 -1748
rect 401 -1749 402 -1737
rect 429 -1749 430 -1737
rect 488 -1770 489 -1748
rect 58 -1751 59 -1737
rect 355 -1751 356 -1737
rect 429 -1770 430 -1750
rect 464 -1751 465 -1737
rect 471 -1770 472 -1750
rect 527 -1751 528 -1737
rect 65 -1753 66 -1737
rect 93 -1753 94 -1737
rect 117 -1770 118 -1752
rect 205 -1770 206 -1752
rect 212 -1753 213 -1737
rect 268 -1753 269 -1737
rect 289 -1770 290 -1752
rect 324 -1753 325 -1737
rect 345 -1753 346 -1737
rect 366 -1770 367 -1752
rect 394 -1753 395 -1737
rect 464 -1770 465 -1752
rect 478 -1770 479 -1752
rect 485 -1753 486 -1737
rect 499 -1753 500 -1737
rect 527 -1770 528 -1752
rect 72 -1755 73 -1737
rect 135 -1770 136 -1754
rect 152 -1770 153 -1754
rect 191 -1755 192 -1737
rect 219 -1770 220 -1754
rect 303 -1755 304 -1737
rect 310 -1770 311 -1754
rect 404 -1770 405 -1754
rect 436 -1755 437 -1737
rect 520 -1770 521 -1754
rect 72 -1770 73 -1756
rect 79 -1757 80 -1737
rect 86 -1757 87 -1737
rect 103 -1757 104 -1737
rect 124 -1770 125 -1756
rect 142 -1770 143 -1756
rect 159 -1757 160 -1737
rect 191 -1770 192 -1756
rect 268 -1770 269 -1756
rect 380 -1757 381 -1737
rect 65 -1770 66 -1758
rect 159 -1770 160 -1758
rect 163 -1759 164 -1737
rect 226 -1770 227 -1758
rect 275 -1759 276 -1737
rect 345 -1770 346 -1758
rect 86 -1770 87 -1760
rect 121 -1770 122 -1760
rect 128 -1770 129 -1760
rect 250 -1761 251 -1737
rect 324 -1770 325 -1760
rect 415 -1761 416 -1737
rect 93 -1770 94 -1762
rect 107 -1770 108 -1762
rect 163 -1770 164 -1762
rect 261 -1770 262 -1762
rect 173 -1770 174 -1764
rect 198 -1765 199 -1737
rect 233 -1765 234 -1737
rect 275 -1770 276 -1764
rect 9 -1767 10 -1737
rect 198 -1770 199 -1766
rect 170 -1769 171 -1737
rect 233 -1770 234 -1768
rect 51 -1780 52 -1778
rect 184 -1780 185 -1778
rect 198 -1780 199 -1778
rect 250 -1799 251 -1779
rect 254 -1799 255 -1779
rect 289 -1780 290 -1778
rect 317 -1780 318 -1778
rect 383 -1780 384 -1778
rect 387 -1799 388 -1779
rect 429 -1780 430 -1778
rect 464 -1780 465 -1778
rect 485 -1780 486 -1778
rect 499 -1799 500 -1779
rect 534 -1780 535 -1778
rect 541 -1780 542 -1778
rect 548 -1780 549 -1778
rect 614 -1780 615 -1778
rect 632 -1780 633 -1778
rect 51 -1799 52 -1781
rect 61 -1782 62 -1778
rect 72 -1782 73 -1778
rect 334 -1782 335 -1778
rect 345 -1782 346 -1778
rect 411 -1799 412 -1781
rect 467 -1799 468 -1781
rect 520 -1782 521 -1778
rect 618 -1782 619 -1778
rect 639 -1799 640 -1781
rect 86 -1784 87 -1778
rect 103 -1784 104 -1778
rect 110 -1799 111 -1783
rect 212 -1784 213 -1778
rect 247 -1799 248 -1783
rect 324 -1784 325 -1778
rect 352 -1784 353 -1778
rect 418 -1784 419 -1778
rect 471 -1784 472 -1778
rect 471 -1799 472 -1783
rect 471 -1784 472 -1778
rect 471 -1799 472 -1783
rect 478 -1784 479 -1778
rect 502 -1784 503 -1778
rect 513 -1784 514 -1778
rect 562 -1784 563 -1778
rect 93 -1786 94 -1778
rect 103 -1799 104 -1785
rect 117 -1786 118 -1778
rect 128 -1786 129 -1778
rect 135 -1786 136 -1778
rect 149 -1799 150 -1785
rect 156 -1786 157 -1778
rect 226 -1786 227 -1778
rect 264 -1799 265 -1785
rect 310 -1786 311 -1778
rect 338 -1786 339 -1778
rect 352 -1799 353 -1785
rect 366 -1786 367 -1778
rect 418 -1799 419 -1785
rect 520 -1799 521 -1785
rect 527 -1786 528 -1778
rect 65 -1788 66 -1778
rect 117 -1799 118 -1787
rect 124 -1799 125 -1787
rect 240 -1788 241 -1778
rect 296 -1788 297 -1778
rect 310 -1799 311 -1787
rect 373 -1799 374 -1787
rect 422 -1788 423 -1778
rect 89 -1799 90 -1789
rect 135 -1799 136 -1789
rect 138 -1799 139 -1789
rect 156 -1799 157 -1789
rect 163 -1790 164 -1778
rect 268 -1790 269 -1778
rect 142 -1792 143 -1778
rect 159 -1792 160 -1778
rect 173 -1799 174 -1791
rect 191 -1792 192 -1778
rect 205 -1799 206 -1791
rect 219 -1792 220 -1778
rect 37 -1794 38 -1778
rect 142 -1799 143 -1793
rect 177 -1794 178 -1778
rect 233 -1794 234 -1778
rect 233 -1799 234 -1795
rect 261 -1796 262 -1778
rect 131 -1799 132 -1797
rect 261 -1799 262 -1797
rect 51 -1809 52 -1807
rect 61 -1809 62 -1807
rect 145 -1809 146 -1807
rect 205 -1809 206 -1807
rect 233 -1809 234 -1807
rect 271 -1809 272 -1807
rect 352 -1809 353 -1807
rect 418 -1809 419 -1807
rect 471 -1809 472 -1807
rect 478 -1809 479 -1807
rect 520 -1809 521 -1807
rect 527 -1809 528 -1807
rect 149 -1811 150 -1807
rect 184 -1811 185 -1807
rect 156 -1813 157 -1807
rect 177 -1813 178 -1807
rect 180 -1813 181 -1807
rect 261 -1813 262 -1807
<< labels >>
rlabel pdiffusion 3 -12 3 -12 0 cellNo=21
rlabel pdiffusion 10 -12 10 -12 0 cellNo=140
rlabel pdiffusion 17 -12 17 -12 0 cellNo=105
rlabel pdiffusion 24 -12 24 -12 0 cellNo=174
rlabel pdiffusion 31 -12 31 -12 0 cellNo=276
rlabel pdiffusion 38 -12 38 -12 0 cellNo=604
rlabel pdiffusion 45 -12 45 -12 0 cellNo=198
rlabel pdiffusion 52 -12 52 -12 0 cellNo=410
rlabel pdiffusion 59 -12 59 -12 0 cellNo=681
rlabel pdiffusion 94 -12 94 -12 0 feedthrough
rlabel pdiffusion 115 -12 115 -12 0 feedthrough
rlabel pdiffusion 122 -12 122 -12 0 cellNo=96
rlabel pdiffusion 129 -12 129 -12 0 feedthrough
rlabel pdiffusion 136 -12 136 -12 0 cellNo=115
rlabel pdiffusion 143 -12 143 -12 0 cellNo=192
rlabel pdiffusion 150 -12 150 -12 0 cellNo=80
rlabel pdiffusion 157 -12 157 -12 0 cellNo=7
rlabel pdiffusion 164 -12 164 -12 0 feedthrough
rlabel pdiffusion 171 -12 171 -12 0 feedthrough
rlabel pdiffusion 178 -12 178 -12 0 cellNo=321
rlabel pdiffusion 185 -12 185 -12 0 feedthrough
rlabel pdiffusion 192 -12 192 -12 0 cellNo=126
rlabel pdiffusion 199 -12 199 -12 0 feedthrough
rlabel pdiffusion 206 -12 206 -12 0 feedthrough
rlabel pdiffusion 213 -12 213 -12 0 feedthrough
rlabel pdiffusion 220 -12 220 -12 0 cellNo=336
rlabel pdiffusion 227 -12 227 -12 0 cellNo=261
rlabel pdiffusion 234 -12 234 -12 0 cellNo=358
rlabel pdiffusion 241 -12 241 -12 0 feedthrough
rlabel pdiffusion 255 -12 255 -12 0 cellNo=361
rlabel pdiffusion 262 -12 262 -12 0 feedthrough
rlabel pdiffusion 290 -12 290 -12 0 cellNo=616
rlabel pdiffusion 339 -12 339 -12 0 cellNo=371
rlabel pdiffusion 3 -39 3 -39 0 cellNo=180
rlabel pdiffusion 10 -39 10 -39 0 cellNo=339
rlabel pdiffusion 17 -39 17 -39 0 cellNo=221
rlabel pdiffusion 31 -39 31 -39 0 cellNo=402
rlabel pdiffusion 38 -39 38 -39 0 cellNo=663
rlabel pdiffusion 45 -39 45 -39 0 cellNo=64
rlabel pdiffusion 52 -39 52 -39 0 cellNo=392
rlabel pdiffusion 66 -39 66 -39 0 cellNo=717
rlabel pdiffusion 73 -39 73 -39 0 feedthrough
rlabel pdiffusion 80 -39 80 -39 0 cellNo=175
rlabel pdiffusion 94 -39 94 -39 0 feedthrough
rlabel pdiffusion 101 -39 101 -39 0 cellNo=91
rlabel pdiffusion 108 -39 108 -39 0 cellNo=168
rlabel pdiffusion 115 -39 115 -39 0 cellNo=513
rlabel pdiffusion 122 -39 122 -39 0 cellNo=277
rlabel pdiffusion 129 -39 129 -39 0 cellNo=716
rlabel pdiffusion 136 -39 136 -39 0 feedthrough
rlabel pdiffusion 143 -39 143 -39 0 cellNo=449
rlabel pdiffusion 150 -39 150 -39 0 cellNo=208
rlabel pdiffusion 157 -39 157 -39 0 cellNo=701
rlabel pdiffusion 164 -39 164 -39 0 cellNo=107
rlabel pdiffusion 171 -39 171 -39 0 feedthrough
rlabel pdiffusion 178 -39 178 -39 0 feedthrough
rlabel pdiffusion 185 -39 185 -39 0 feedthrough
rlabel pdiffusion 192 -39 192 -39 0 feedthrough
rlabel pdiffusion 199 -39 199 -39 0 feedthrough
rlabel pdiffusion 206 -39 206 -39 0 cellNo=55
rlabel pdiffusion 213 -39 213 -39 0 feedthrough
rlabel pdiffusion 220 -39 220 -39 0 feedthrough
rlabel pdiffusion 227 -39 227 -39 0 feedthrough
rlabel pdiffusion 234 -39 234 -39 0 feedthrough
rlabel pdiffusion 241 -39 241 -39 0 feedthrough
rlabel pdiffusion 248 -39 248 -39 0 feedthrough
rlabel pdiffusion 255 -39 255 -39 0 feedthrough
rlabel pdiffusion 269 -39 269 -39 0 cellNo=661
rlabel pdiffusion 276 -39 276 -39 0 feedthrough
rlabel pdiffusion 283 -39 283 -39 0 cellNo=178
rlabel pdiffusion 290 -39 290 -39 0 cellNo=45
rlabel pdiffusion 297 -39 297 -39 0 feedthrough
rlabel pdiffusion 311 -39 311 -39 0 cellNo=628
rlabel pdiffusion 318 -39 318 -39 0 feedthrough
rlabel pdiffusion 325 -39 325 -39 0 feedthrough
rlabel pdiffusion 332 -39 332 -39 0 cellNo=58
rlabel pdiffusion 339 -39 339 -39 0 feedthrough
rlabel pdiffusion 346 -39 346 -39 0 feedthrough
rlabel pdiffusion 353 -39 353 -39 0 feedthrough
rlabel pdiffusion 388 -39 388 -39 0 feedthrough
rlabel pdiffusion 402 -39 402 -39 0 cellNo=611
rlabel pdiffusion 3 -74 3 -74 0 cellNo=88
rlabel pdiffusion 17 -74 17 -74 0 feedthrough
rlabel pdiffusion 24 -74 24 -74 0 feedthrough
rlabel pdiffusion 31 -74 31 -74 0 cellNo=253
rlabel pdiffusion 38 -74 38 -74 0 cellNo=82
rlabel pdiffusion 45 -74 45 -74 0 feedthrough
rlabel pdiffusion 52 -74 52 -74 0 cellNo=325
rlabel pdiffusion 59 -74 59 -74 0 cellNo=605
rlabel pdiffusion 66 -74 66 -74 0 feedthrough
rlabel pdiffusion 73 -74 73 -74 0 cellNo=566
rlabel pdiffusion 80 -74 80 -74 0 cellNo=22
rlabel pdiffusion 87 -74 87 -74 0 cellNo=559
rlabel pdiffusion 94 -74 94 -74 0 feedthrough
rlabel pdiffusion 101 -74 101 -74 0 feedthrough
rlabel pdiffusion 108 -74 108 -74 0 cellNo=120
rlabel pdiffusion 115 -74 115 -74 0 cellNo=574
rlabel pdiffusion 122 -74 122 -74 0 feedthrough
rlabel pdiffusion 129 -74 129 -74 0 feedthrough
rlabel pdiffusion 136 -74 136 -74 0 feedthrough
rlabel pdiffusion 143 -74 143 -74 0 feedthrough
rlabel pdiffusion 150 -74 150 -74 0 cellNo=379
rlabel pdiffusion 157 -74 157 -74 0 feedthrough
rlabel pdiffusion 164 -74 164 -74 0 feedthrough
rlabel pdiffusion 171 -74 171 -74 0 feedthrough
rlabel pdiffusion 178 -74 178 -74 0 cellNo=218
rlabel pdiffusion 185 -74 185 -74 0 cellNo=390
rlabel pdiffusion 192 -74 192 -74 0 cellNo=102
rlabel pdiffusion 199 -74 199 -74 0 cellNo=322
rlabel pdiffusion 206 -74 206 -74 0 cellNo=548
rlabel pdiffusion 213 -74 213 -74 0 feedthrough
rlabel pdiffusion 220 -74 220 -74 0 cellNo=121
rlabel pdiffusion 227 -74 227 -74 0 feedthrough
rlabel pdiffusion 234 -74 234 -74 0 feedthrough
rlabel pdiffusion 241 -74 241 -74 0 feedthrough
rlabel pdiffusion 248 -74 248 -74 0 cellNo=543
rlabel pdiffusion 255 -74 255 -74 0 feedthrough
rlabel pdiffusion 262 -74 262 -74 0 cellNo=67
rlabel pdiffusion 269 -74 269 -74 0 cellNo=153
rlabel pdiffusion 276 -74 276 -74 0 feedthrough
rlabel pdiffusion 283 -74 283 -74 0 cellNo=507
rlabel pdiffusion 290 -74 290 -74 0 feedthrough
rlabel pdiffusion 297 -74 297 -74 0 cellNo=561
rlabel pdiffusion 304 -74 304 -74 0 cellNo=579
rlabel pdiffusion 311 -74 311 -74 0 feedthrough
rlabel pdiffusion 318 -74 318 -74 0 feedthrough
rlabel pdiffusion 325 -74 325 -74 0 feedthrough
rlabel pdiffusion 332 -74 332 -74 0 feedthrough
rlabel pdiffusion 339 -74 339 -74 0 cellNo=329
rlabel pdiffusion 346 -74 346 -74 0 feedthrough
rlabel pdiffusion 353 -74 353 -74 0 cellNo=511
rlabel pdiffusion 360 -74 360 -74 0 feedthrough
rlabel pdiffusion 367 -74 367 -74 0 feedthrough
rlabel pdiffusion 374 -74 374 -74 0 feedthrough
rlabel pdiffusion 381 -74 381 -74 0 feedthrough
rlabel pdiffusion 388 -74 388 -74 0 feedthrough
rlabel pdiffusion 395 -74 395 -74 0 cellNo=650
rlabel pdiffusion 402 -74 402 -74 0 feedthrough
rlabel pdiffusion 409 -74 409 -74 0 feedthrough
rlabel pdiffusion 416 -74 416 -74 0 feedthrough
rlabel pdiffusion 423 -74 423 -74 0 feedthrough
rlabel pdiffusion 430 -74 430 -74 0 cellNo=310
rlabel pdiffusion 437 -74 437 -74 0 feedthrough
rlabel pdiffusion 3 -127 3 -127 0 cellNo=25
rlabel pdiffusion 10 -127 10 -127 0 cellNo=291
rlabel pdiffusion 17 -127 17 -127 0 cellNo=412
rlabel pdiffusion 24 -127 24 -127 0 cellNo=331
rlabel pdiffusion 31 -127 31 -127 0 cellNo=130
rlabel pdiffusion 38 -127 38 -127 0 cellNo=237
rlabel pdiffusion 45 -127 45 -127 0 cellNo=191
rlabel pdiffusion 52 -127 52 -127 0 cellNo=81
rlabel pdiffusion 59 -127 59 -127 0 feedthrough
rlabel pdiffusion 66 -127 66 -127 0 cellNo=199
rlabel pdiffusion 73 -127 73 -127 0 cellNo=63
rlabel pdiffusion 80 -127 80 -127 0 feedthrough
rlabel pdiffusion 87 -127 87 -127 0 feedthrough
rlabel pdiffusion 94 -127 94 -127 0 feedthrough
rlabel pdiffusion 101 -127 101 -127 0 cellNo=287
rlabel pdiffusion 108 -127 108 -127 0 feedthrough
rlabel pdiffusion 115 -127 115 -127 0 cellNo=70
rlabel pdiffusion 122 -127 122 -127 0 feedthrough
rlabel pdiffusion 129 -127 129 -127 0 feedthrough
rlabel pdiffusion 136 -127 136 -127 0 cellNo=593
rlabel pdiffusion 143 -127 143 -127 0 feedthrough
rlabel pdiffusion 150 -127 150 -127 0 feedthrough
rlabel pdiffusion 157 -127 157 -127 0 cellNo=664
rlabel pdiffusion 164 -127 164 -127 0 feedthrough
rlabel pdiffusion 171 -127 171 -127 0 cellNo=50
rlabel pdiffusion 178 -127 178 -127 0 cellNo=360
rlabel pdiffusion 185 -127 185 -127 0 cellNo=476
rlabel pdiffusion 192 -127 192 -127 0 feedthrough
rlabel pdiffusion 199 -127 199 -127 0 feedthrough
rlabel pdiffusion 206 -127 206 -127 0 feedthrough
rlabel pdiffusion 213 -127 213 -127 0 feedthrough
rlabel pdiffusion 220 -127 220 -127 0 feedthrough
rlabel pdiffusion 227 -127 227 -127 0 feedthrough
rlabel pdiffusion 234 -127 234 -127 0 feedthrough
rlabel pdiffusion 241 -127 241 -127 0 cellNo=420
rlabel pdiffusion 248 -127 248 -127 0 feedthrough
rlabel pdiffusion 255 -127 255 -127 0 cellNo=213
rlabel pdiffusion 262 -127 262 -127 0 feedthrough
rlabel pdiffusion 269 -127 269 -127 0 feedthrough
rlabel pdiffusion 276 -127 276 -127 0 feedthrough
rlabel pdiffusion 283 -127 283 -127 0 cellNo=501
rlabel pdiffusion 290 -127 290 -127 0 cellNo=28
rlabel pdiffusion 297 -127 297 -127 0 feedthrough
rlabel pdiffusion 304 -127 304 -127 0 feedthrough
rlabel pdiffusion 311 -127 311 -127 0 feedthrough
rlabel pdiffusion 318 -127 318 -127 0 feedthrough
rlabel pdiffusion 325 -127 325 -127 0 cellNo=639
rlabel pdiffusion 332 -127 332 -127 0 cellNo=555
rlabel pdiffusion 339 -127 339 -127 0 cellNo=57
rlabel pdiffusion 346 -127 346 -127 0 feedthrough
rlabel pdiffusion 353 -127 353 -127 0 cellNo=374
rlabel pdiffusion 360 -127 360 -127 0 feedthrough
rlabel pdiffusion 367 -127 367 -127 0 feedthrough
rlabel pdiffusion 374 -127 374 -127 0 cellNo=534
rlabel pdiffusion 381 -127 381 -127 0 cellNo=377
rlabel pdiffusion 388 -127 388 -127 0 feedthrough
rlabel pdiffusion 395 -127 395 -127 0 feedthrough
rlabel pdiffusion 402 -127 402 -127 0 feedthrough
rlabel pdiffusion 409 -127 409 -127 0 feedthrough
rlabel pdiffusion 416 -127 416 -127 0 feedthrough
rlabel pdiffusion 423 -127 423 -127 0 feedthrough
rlabel pdiffusion 430 -127 430 -127 0 feedthrough
rlabel pdiffusion 437 -127 437 -127 0 feedthrough
rlabel pdiffusion 444 -127 444 -127 0 feedthrough
rlabel pdiffusion 451 -127 451 -127 0 feedthrough
rlabel pdiffusion 458 -127 458 -127 0 feedthrough
rlabel pdiffusion 465 -127 465 -127 0 feedthrough
rlabel pdiffusion 472 -127 472 -127 0 feedthrough
rlabel pdiffusion 479 -127 479 -127 0 feedthrough
rlabel pdiffusion 486 -127 486 -127 0 feedthrough
rlabel pdiffusion 493 -127 493 -127 0 feedthrough
rlabel pdiffusion 500 -127 500 -127 0 feedthrough
rlabel pdiffusion 507 -127 507 -127 0 feedthrough
rlabel pdiffusion 514 -127 514 -127 0 feedthrough
rlabel pdiffusion 521 -127 521 -127 0 feedthrough
rlabel pdiffusion 3 -202 3 -202 0 cellNo=177
rlabel pdiffusion 10 -202 10 -202 0 cellNo=244
rlabel pdiffusion 17 -202 17 -202 0 cellNo=565
rlabel pdiffusion 24 -202 24 -202 0 cellNo=660
rlabel pdiffusion 31 -202 31 -202 0 cellNo=505
rlabel pdiffusion 38 -202 38 -202 0 cellNo=247
rlabel pdiffusion 45 -202 45 -202 0 feedthrough
rlabel pdiffusion 52 -202 52 -202 0 cellNo=629
rlabel pdiffusion 59 -202 59 -202 0 feedthrough
rlabel pdiffusion 66 -202 66 -202 0 feedthrough
rlabel pdiffusion 73 -202 73 -202 0 feedthrough
rlabel pdiffusion 80 -202 80 -202 0 feedthrough
rlabel pdiffusion 87 -202 87 -202 0 cellNo=196
rlabel pdiffusion 94 -202 94 -202 0 feedthrough
rlabel pdiffusion 101 -202 101 -202 0 feedthrough
rlabel pdiffusion 108 -202 108 -202 0 feedthrough
rlabel pdiffusion 115 -202 115 -202 0 cellNo=298
rlabel pdiffusion 122 -202 122 -202 0 feedthrough
rlabel pdiffusion 129 -202 129 -202 0 feedthrough
rlabel pdiffusion 136 -202 136 -202 0 cellNo=472
rlabel pdiffusion 143 -202 143 -202 0 cellNo=84
rlabel pdiffusion 150 -202 150 -202 0 cellNo=571
rlabel pdiffusion 157 -202 157 -202 0 feedthrough
rlabel pdiffusion 164 -202 164 -202 0 feedthrough
rlabel pdiffusion 171 -202 171 -202 0 feedthrough
rlabel pdiffusion 178 -202 178 -202 0 cellNo=231
rlabel pdiffusion 185 -202 185 -202 0 cellNo=264
rlabel pdiffusion 192 -202 192 -202 0 feedthrough
rlabel pdiffusion 199 -202 199 -202 0 cellNo=459
rlabel pdiffusion 206 -202 206 -202 0 cellNo=17
rlabel pdiffusion 213 -202 213 -202 0 cellNo=111
rlabel pdiffusion 220 -202 220 -202 0 feedthrough
rlabel pdiffusion 227 -202 227 -202 0 feedthrough
rlabel pdiffusion 234 -202 234 -202 0 feedthrough
rlabel pdiffusion 241 -202 241 -202 0 feedthrough
rlabel pdiffusion 248 -202 248 -202 0 cellNo=149
rlabel pdiffusion 255 -202 255 -202 0 cellNo=590
rlabel pdiffusion 262 -202 262 -202 0 feedthrough
rlabel pdiffusion 269 -202 269 -202 0 cellNo=473
rlabel pdiffusion 276 -202 276 -202 0 feedthrough
rlabel pdiffusion 283 -202 283 -202 0 cellNo=141
rlabel pdiffusion 290 -202 290 -202 0 cellNo=489
rlabel pdiffusion 297 -202 297 -202 0 feedthrough
rlabel pdiffusion 304 -202 304 -202 0 feedthrough
rlabel pdiffusion 311 -202 311 -202 0 cellNo=452
rlabel pdiffusion 318 -202 318 -202 0 feedthrough
rlabel pdiffusion 325 -202 325 -202 0 feedthrough
rlabel pdiffusion 332 -202 332 -202 0 feedthrough
rlabel pdiffusion 339 -202 339 -202 0 cellNo=514
rlabel pdiffusion 346 -202 346 -202 0 feedthrough
rlabel pdiffusion 353 -202 353 -202 0 feedthrough
rlabel pdiffusion 360 -202 360 -202 0 feedthrough
rlabel pdiffusion 367 -202 367 -202 0 feedthrough
rlabel pdiffusion 374 -202 374 -202 0 feedthrough
rlabel pdiffusion 381 -202 381 -202 0 feedthrough
rlabel pdiffusion 388 -202 388 -202 0 cellNo=290
rlabel pdiffusion 395 -202 395 -202 0 feedthrough
rlabel pdiffusion 402 -202 402 -202 0 feedthrough
rlabel pdiffusion 409 -202 409 -202 0 cellNo=61
rlabel pdiffusion 416 -202 416 -202 0 feedthrough
rlabel pdiffusion 423 -202 423 -202 0 cellNo=458
rlabel pdiffusion 430 -202 430 -202 0 feedthrough
rlabel pdiffusion 437 -202 437 -202 0 feedthrough
rlabel pdiffusion 444 -202 444 -202 0 feedthrough
rlabel pdiffusion 451 -202 451 -202 0 feedthrough
rlabel pdiffusion 458 -202 458 -202 0 feedthrough
rlabel pdiffusion 465 -202 465 -202 0 feedthrough
rlabel pdiffusion 472 -202 472 -202 0 feedthrough
rlabel pdiffusion 479 -202 479 -202 0 feedthrough
rlabel pdiffusion 486 -202 486 -202 0 feedthrough
rlabel pdiffusion 493 -202 493 -202 0 feedthrough
rlabel pdiffusion 500 -202 500 -202 0 feedthrough
rlabel pdiffusion 507 -202 507 -202 0 feedthrough
rlabel pdiffusion 514 -202 514 -202 0 feedthrough
rlabel pdiffusion 521 -202 521 -202 0 feedthrough
rlabel pdiffusion 528 -202 528 -202 0 feedthrough
rlabel pdiffusion 535 -202 535 -202 0 feedthrough
rlabel pdiffusion 542 -202 542 -202 0 feedthrough
rlabel pdiffusion 549 -202 549 -202 0 feedthrough
rlabel pdiffusion 556 -202 556 -202 0 feedthrough
rlabel pdiffusion 563 -202 563 -202 0 feedthrough
rlabel pdiffusion 570 -202 570 -202 0 feedthrough
rlabel pdiffusion 577 -202 577 -202 0 feedthrough
rlabel pdiffusion 584 -202 584 -202 0 feedthrough
rlabel pdiffusion 591 -202 591 -202 0 feedthrough
rlabel pdiffusion 598 -202 598 -202 0 feedthrough
rlabel pdiffusion 605 -202 605 -202 0 feedthrough
rlabel pdiffusion 612 -202 612 -202 0 feedthrough
rlabel pdiffusion 619 -202 619 -202 0 feedthrough
rlabel pdiffusion 626 -202 626 -202 0 feedthrough
rlabel pdiffusion 633 -202 633 -202 0 feedthrough
rlabel pdiffusion 640 -202 640 -202 0 feedthrough
rlabel pdiffusion 647 -202 647 -202 0 feedthrough
rlabel pdiffusion 654 -202 654 -202 0 feedthrough
rlabel pdiffusion 661 -202 661 -202 0 feedthrough
rlabel pdiffusion 3 -275 3 -275 0 cellNo=99
rlabel pdiffusion 10 -275 10 -275 0 cellNo=439
rlabel pdiffusion 17 -275 17 -275 0 cellNo=299
rlabel pdiffusion 24 -275 24 -275 0 cellNo=355
rlabel pdiffusion 31 -275 31 -275 0 feedthrough
rlabel pdiffusion 38 -275 38 -275 0 cellNo=496
rlabel pdiffusion 45 -275 45 -275 0 cellNo=300
rlabel pdiffusion 52 -275 52 -275 0 feedthrough
rlabel pdiffusion 59 -275 59 -275 0 cellNo=258
rlabel pdiffusion 66 -275 66 -275 0 feedthrough
rlabel pdiffusion 73 -275 73 -275 0 feedthrough
rlabel pdiffusion 80 -275 80 -275 0 cellNo=494
rlabel pdiffusion 87 -275 87 -275 0 cellNo=408
rlabel pdiffusion 94 -275 94 -275 0 feedthrough
rlabel pdiffusion 101 -275 101 -275 0 cellNo=348
rlabel pdiffusion 108 -275 108 -275 0 feedthrough
rlabel pdiffusion 115 -275 115 -275 0 feedthrough
rlabel pdiffusion 122 -275 122 -275 0 cellNo=376
rlabel pdiffusion 129 -275 129 -275 0 feedthrough
rlabel pdiffusion 136 -275 136 -275 0 feedthrough
rlabel pdiffusion 143 -275 143 -275 0 feedthrough
rlabel pdiffusion 150 -275 150 -275 0 feedthrough
rlabel pdiffusion 157 -275 157 -275 0 cellNo=705
rlabel pdiffusion 164 -275 164 -275 0 feedthrough
rlabel pdiffusion 171 -275 171 -275 0 feedthrough
rlabel pdiffusion 178 -275 178 -275 0 cellNo=13
rlabel pdiffusion 185 -275 185 -275 0 feedthrough
rlabel pdiffusion 192 -275 192 -275 0 feedthrough
rlabel pdiffusion 199 -275 199 -275 0 feedthrough
rlabel pdiffusion 206 -275 206 -275 0 feedthrough
rlabel pdiffusion 213 -275 213 -275 0 feedthrough
rlabel pdiffusion 220 -275 220 -275 0 feedthrough
rlabel pdiffusion 227 -275 227 -275 0 feedthrough
rlabel pdiffusion 234 -275 234 -275 0 feedthrough
rlabel pdiffusion 241 -275 241 -275 0 cellNo=34
rlabel pdiffusion 248 -275 248 -275 0 cellNo=450
rlabel pdiffusion 255 -275 255 -275 0 cellNo=343
rlabel pdiffusion 262 -275 262 -275 0 feedthrough
rlabel pdiffusion 269 -275 269 -275 0 cellNo=414
rlabel pdiffusion 276 -275 276 -275 0 cellNo=455
rlabel pdiffusion 283 -275 283 -275 0 cellNo=131
rlabel pdiffusion 290 -275 290 -275 0 feedthrough
rlabel pdiffusion 297 -275 297 -275 0 cellNo=195
rlabel pdiffusion 304 -275 304 -275 0 cellNo=506
rlabel pdiffusion 311 -275 311 -275 0 feedthrough
rlabel pdiffusion 318 -275 318 -275 0 cellNo=375
rlabel pdiffusion 325 -275 325 -275 0 feedthrough
rlabel pdiffusion 332 -275 332 -275 0 cellNo=690
rlabel pdiffusion 339 -275 339 -275 0 feedthrough
rlabel pdiffusion 346 -275 346 -275 0 feedthrough
rlabel pdiffusion 353 -275 353 -275 0 cellNo=667
rlabel pdiffusion 360 -275 360 -275 0 feedthrough
rlabel pdiffusion 367 -275 367 -275 0 cellNo=328
rlabel pdiffusion 374 -275 374 -275 0 feedthrough
rlabel pdiffusion 381 -275 381 -275 0 feedthrough
rlabel pdiffusion 388 -275 388 -275 0 feedthrough
rlabel pdiffusion 395 -275 395 -275 0 feedthrough
rlabel pdiffusion 402 -275 402 -275 0 feedthrough
rlabel pdiffusion 409 -275 409 -275 0 feedthrough
rlabel pdiffusion 416 -275 416 -275 0 feedthrough
rlabel pdiffusion 423 -275 423 -275 0 feedthrough
rlabel pdiffusion 430 -275 430 -275 0 feedthrough
rlabel pdiffusion 437 -275 437 -275 0 feedthrough
rlabel pdiffusion 444 -275 444 -275 0 feedthrough
rlabel pdiffusion 451 -275 451 -275 0 feedthrough
rlabel pdiffusion 458 -275 458 -275 0 feedthrough
rlabel pdiffusion 465 -275 465 -275 0 feedthrough
rlabel pdiffusion 472 -275 472 -275 0 feedthrough
rlabel pdiffusion 479 -275 479 -275 0 feedthrough
rlabel pdiffusion 486 -275 486 -275 0 feedthrough
rlabel pdiffusion 493 -275 493 -275 0 feedthrough
rlabel pdiffusion 500 -275 500 -275 0 feedthrough
rlabel pdiffusion 507 -275 507 -275 0 feedthrough
rlabel pdiffusion 514 -275 514 -275 0 feedthrough
rlabel pdiffusion 521 -275 521 -275 0 feedthrough
rlabel pdiffusion 528 -275 528 -275 0 feedthrough
rlabel pdiffusion 535 -275 535 -275 0 feedthrough
rlabel pdiffusion 542 -275 542 -275 0 feedthrough
rlabel pdiffusion 549 -275 549 -275 0 feedthrough
rlabel pdiffusion 563 -275 563 -275 0 feedthrough
rlabel pdiffusion 570 -275 570 -275 0 feedthrough
rlabel pdiffusion 577 -275 577 -275 0 feedthrough
rlabel pdiffusion 584 -275 584 -275 0 feedthrough
rlabel pdiffusion 591 -275 591 -275 0 feedthrough
rlabel pdiffusion 598 -275 598 -275 0 feedthrough
rlabel pdiffusion 605 -275 605 -275 0 feedthrough
rlabel pdiffusion 612 -275 612 -275 0 feedthrough
rlabel pdiffusion 619 -275 619 -275 0 cellNo=170
rlabel pdiffusion 626 -275 626 -275 0 feedthrough
rlabel pdiffusion 633 -275 633 -275 0 feedthrough
rlabel pdiffusion 640 -275 640 -275 0 cellNo=42
rlabel pdiffusion 668 -275 668 -275 0 feedthrough
rlabel pdiffusion 3 -340 3 -340 0 cellNo=474
rlabel pdiffusion 10 -340 10 -340 0 cellNo=426
rlabel pdiffusion 17 -340 17 -340 0 cellNo=148
rlabel pdiffusion 24 -340 24 -340 0 cellNo=330
rlabel pdiffusion 31 -340 31 -340 0 cellNo=280
rlabel pdiffusion 38 -340 38 -340 0 feedthrough
rlabel pdiffusion 45 -340 45 -340 0 cellNo=12
rlabel pdiffusion 52 -340 52 -340 0 cellNo=288
rlabel pdiffusion 59 -340 59 -340 0 feedthrough
rlabel pdiffusion 66 -340 66 -340 0 cellNo=146
rlabel pdiffusion 73 -340 73 -340 0 cellNo=152
rlabel pdiffusion 80 -340 80 -340 0 cellNo=490
rlabel pdiffusion 87 -340 87 -340 0 cellNo=110
rlabel pdiffusion 94 -340 94 -340 0 feedthrough
rlabel pdiffusion 101 -340 101 -340 0 cellNo=296
rlabel pdiffusion 108 -340 108 -340 0 feedthrough
rlabel pdiffusion 115 -340 115 -340 0 feedthrough
rlabel pdiffusion 122 -340 122 -340 0 feedthrough
rlabel pdiffusion 129 -340 129 -340 0 feedthrough
rlabel pdiffusion 136 -340 136 -340 0 cellNo=157
rlabel pdiffusion 143 -340 143 -340 0 cellNo=538
rlabel pdiffusion 150 -340 150 -340 0 feedthrough
rlabel pdiffusion 157 -340 157 -340 0 cellNo=172
rlabel pdiffusion 164 -340 164 -340 0 cellNo=689
rlabel pdiffusion 171 -340 171 -340 0 feedthrough
rlabel pdiffusion 178 -340 178 -340 0 feedthrough
rlabel pdiffusion 185 -340 185 -340 0 cellNo=428
rlabel pdiffusion 192 -340 192 -340 0 feedthrough
rlabel pdiffusion 199 -340 199 -340 0 cellNo=159
rlabel pdiffusion 206 -340 206 -340 0 feedthrough
rlabel pdiffusion 213 -340 213 -340 0 feedthrough
rlabel pdiffusion 220 -340 220 -340 0 feedthrough
rlabel pdiffusion 227 -340 227 -340 0 feedthrough
rlabel pdiffusion 234 -340 234 -340 0 feedthrough
rlabel pdiffusion 241 -340 241 -340 0 cellNo=240
rlabel pdiffusion 248 -340 248 -340 0 feedthrough
rlabel pdiffusion 255 -340 255 -340 0 feedthrough
rlabel pdiffusion 262 -340 262 -340 0 feedthrough
rlabel pdiffusion 269 -340 269 -340 0 feedthrough
rlabel pdiffusion 276 -340 276 -340 0 feedthrough
rlabel pdiffusion 283 -340 283 -340 0 feedthrough
rlabel pdiffusion 290 -340 290 -340 0 feedthrough
rlabel pdiffusion 297 -340 297 -340 0 feedthrough
rlabel pdiffusion 304 -340 304 -340 0 feedthrough
rlabel pdiffusion 311 -340 311 -340 0 cellNo=6
rlabel pdiffusion 318 -340 318 -340 0 cellNo=89
rlabel pdiffusion 325 -340 325 -340 0 cellNo=211
rlabel pdiffusion 332 -340 332 -340 0 feedthrough
rlabel pdiffusion 339 -340 339 -340 0 cellNo=69
rlabel pdiffusion 346 -340 346 -340 0 feedthrough
rlabel pdiffusion 353 -340 353 -340 0 cellNo=268
rlabel pdiffusion 360 -340 360 -340 0 cellNo=457
rlabel pdiffusion 367 -340 367 -340 0 feedthrough
rlabel pdiffusion 374 -340 374 -340 0 feedthrough
rlabel pdiffusion 381 -340 381 -340 0 feedthrough
rlabel pdiffusion 388 -340 388 -340 0 cellNo=186
rlabel pdiffusion 395 -340 395 -340 0 feedthrough
rlabel pdiffusion 402 -340 402 -340 0 feedthrough
rlabel pdiffusion 409 -340 409 -340 0 feedthrough
rlabel pdiffusion 416 -340 416 -340 0 feedthrough
rlabel pdiffusion 423 -340 423 -340 0 feedthrough
rlabel pdiffusion 430 -340 430 -340 0 feedthrough
rlabel pdiffusion 437 -340 437 -340 0 feedthrough
rlabel pdiffusion 444 -340 444 -340 0 feedthrough
rlabel pdiffusion 451 -340 451 -340 0 feedthrough
rlabel pdiffusion 458 -340 458 -340 0 feedthrough
rlabel pdiffusion 465 -340 465 -340 0 feedthrough
rlabel pdiffusion 472 -340 472 -340 0 feedthrough
rlabel pdiffusion 479 -340 479 -340 0 feedthrough
rlabel pdiffusion 486 -340 486 -340 0 feedthrough
rlabel pdiffusion 493 -340 493 -340 0 cellNo=295
rlabel pdiffusion 500 -340 500 -340 0 feedthrough
rlabel pdiffusion 507 -340 507 -340 0 feedthrough
rlabel pdiffusion 514 -340 514 -340 0 feedthrough
rlabel pdiffusion 521 -340 521 -340 0 feedthrough
rlabel pdiffusion 528 -340 528 -340 0 feedthrough
rlabel pdiffusion 535 -340 535 -340 0 feedthrough
rlabel pdiffusion 542 -340 542 -340 0 feedthrough
rlabel pdiffusion 549 -340 549 -340 0 feedthrough
rlabel pdiffusion 556 -340 556 -340 0 feedthrough
rlabel pdiffusion 563 -340 563 -340 0 feedthrough
rlabel pdiffusion 570 -340 570 -340 0 feedthrough
rlabel pdiffusion 577 -340 577 -340 0 feedthrough
rlabel pdiffusion 584 -340 584 -340 0 feedthrough
rlabel pdiffusion 591 -340 591 -340 0 feedthrough
rlabel pdiffusion 605 -340 605 -340 0 feedthrough
rlabel pdiffusion 612 -340 612 -340 0 feedthrough
rlabel pdiffusion 619 -340 619 -340 0 feedthrough
rlabel pdiffusion 626 -340 626 -340 0 feedthrough
rlabel pdiffusion 633 -340 633 -340 0 feedthrough
rlabel pdiffusion 640 -340 640 -340 0 feedthrough
rlabel pdiffusion 647 -340 647 -340 0 feedthrough
rlabel pdiffusion 654 -340 654 -340 0 feedthrough
rlabel pdiffusion 661 -340 661 -340 0 feedthrough
rlabel pdiffusion 668 -340 668 -340 0 feedthrough
rlabel pdiffusion 675 -340 675 -340 0 feedthrough
rlabel pdiffusion 710 -340 710 -340 0 feedthrough
rlabel pdiffusion 3 -407 3 -407 0 cellNo=100
rlabel pdiffusion 10 -407 10 -407 0 cellNo=228
rlabel pdiffusion 24 -407 24 -407 0 feedthrough
rlabel pdiffusion 31 -407 31 -407 0 cellNo=524
rlabel pdiffusion 38 -407 38 -407 0 feedthrough
rlabel pdiffusion 45 -407 45 -407 0 feedthrough
rlabel pdiffusion 52 -407 52 -407 0 feedthrough
rlabel pdiffusion 59 -407 59 -407 0 feedthrough
rlabel pdiffusion 66 -407 66 -407 0 cellNo=598
rlabel pdiffusion 73 -407 73 -407 0 feedthrough
rlabel pdiffusion 80 -407 80 -407 0 feedthrough
rlabel pdiffusion 87 -407 87 -407 0 feedthrough
rlabel pdiffusion 94 -407 94 -407 0 cellNo=229
rlabel pdiffusion 101 -407 101 -407 0 feedthrough
rlabel pdiffusion 108 -407 108 -407 0 cellNo=52
rlabel pdiffusion 115 -407 115 -407 0 cellNo=251
rlabel pdiffusion 122 -407 122 -407 0 cellNo=133
rlabel pdiffusion 129 -407 129 -407 0 feedthrough
rlabel pdiffusion 136 -407 136 -407 0 feedthrough
rlabel pdiffusion 143 -407 143 -407 0 feedthrough
rlabel pdiffusion 150 -407 150 -407 0 feedthrough
rlabel pdiffusion 157 -407 157 -407 0 cellNo=239
rlabel pdiffusion 164 -407 164 -407 0 feedthrough
rlabel pdiffusion 171 -407 171 -407 0 feedthrough
rlabel pdiffusion 178 -407 178 -407 0 feedthrough
rlabel pdiffusion 185 -407 185 -407 0 cellNo=640
rlabel pdiffusion 192 -407 192 -407 0 feedthrough
rlabel pdiffusion 199 -407 199 -407 0 feedthrough
rlabel pdiffusion 206 -407 206 -407 0 feedthrough
rlabel pdiffusion 213 -407 213 -407 0 feedthrough
rlabel pdiffusion 220 -407 220 -407 0 feedthrough
rlabel pdiffusion 227 -407 227 -407 0 cellNo=350
rlabel pdiffusion 234 -407 234 -407 0 feedthrough
rlabel pdiffusion 241 -407 241 -407 0 cellNo=124
rlabel pdiffusion 248 -407 248 -407 0 feedthrough
rlabel pdiffusion 255 -407 255 -407 0 feedthrough
rlabel pdiffusion 262 -407 262 -407 0 feedthrough
rlabel pdiffusion 269 -407 269 -407 0 feedthrough
rlabel pdiffusion 276 -407 276 -407 0 feedthrough
rlabel pdiffusion 283 -407 283 -407 0 cellNo=596
rlabel pdiffusion 290 -407 290 -407 0 feedthrough
rlabel pdiffusion 297 -407 297 -407 0 feedthrough
rlabel pdiffusion 304 -407 304 -407 0 feedthrough
rlabel pdiffusion 311 -407 311 -407 0 feedthrough
rlabel pdiffusion 318 -407 318 -407 0 feedthrough
rlabel pdiffusion 325 -407 325 -407 0 cellNo=623
rlabel pdiffusion 332 -407 332 -407 0 cellNo=521
rlabel pdiffusion 339 -407 339 -407 0 cellNo=5
rlabel pdiffusion 346 -407 346 -407 0 feedthrough
rlabel pdiffusion 353 -407 353 -407 0 cellNo=357
rlabel pdiffusion 360 -407 360 -407 0 feedthrough
rlabel pdiffusion 367 -407 367 -407 0 feedthrough
rlabel pdiffusion 374 -407 374 -407 0 cellNo=51
rlabel pdiffusion 381 -407 381 -407 0 cellNo=29
rlabel pdiffusion 388 -407 388 -407 0 cellNo=535
rlabel pdiffusion 395 -407 395 -407 0 feedthrough
rlabel pdiffusion 402 -407 402 -407 0 feedthrough
rlabel pdiffusion 409 -407 409 -407 0 cellNo=558
rlabel pdiffusion 416 -407 416 -407 0 feedthrough
rlabel pdiffusion 423 -407 423 -407 0 feedthrough
rlabel pdiffusion 430 -407 430 -407 0 cellNo=315
rlabel pdiffusion 437 -407 437 -407 0 feedthrough
rlabel pdiffusion 444 -407 444 -407 0 feedthrough
rlabel pdiffusion 451 -407 451 -407 0 feedthrough
rlabel pdiffusion 458 -407 458 -407 0 feedthrough
rlabel pdiffusion 465 -407 465 -407 0 cellNo=435
rlabel pdiffusion 472 -407 472 -407 0 feedthrough
rlabel pdiffusion 479 -407 479 -407 0 cellNo=363
rlabel pdiffusion 486 -407 486 -407 0 feedthrough
rlabel pdiffusion 493 -407 493 -407 0 feedthrough
rlabel pdiffusion 500 -407 500 -407 0 cellNo=292
rlabel pdiffusion 507 -407 507 -407 0 feedthrough
rlabel pdiffusion 514 -407 514 -407 0 feedthrough
rlabel pdiffusion 521 -407 521 -407 0 feedthrough
rlabel pdiffusion 528 -407 528 -407 0 feedthrough
rlabel pdiffusion 535 -407 535 -407 0 feedthrough
rlabel pdiffusion 542 -407 542 -407 0 feedthrough
rlabel pdiffusion 549 -407 549 -407 0 feedthrough
rlabel pdiffusion 556 -407 556 -407 0 feedthrough
rlabel pdiffusion 563 -407 563 -407 0 feedthrough
rlabel pdiffusion 570 -407 570 -407 0 feedthrough
rlabel pdiffusion 577 -407 577 -407 0 feedthrough
rlabel pdiffusion 584 -407 584 -407 0 feedthrough
rlabel pdiffusion 591 -407 591 -407 0 feedthrough
rlabel pdiffusion 598 -407 598 -407 0 feedthrough
rlabel pdiffusion 605 -407 605 -407 0 feedthrough
rlabel pdiffusion 612 -407 612 -407 0 feedthrough
rlabel pdiffusion 619 -407 619 -407 0 feedthrough
rlabel pdiffusion 626 -407 626 -407 0 feedthrough
rlabel pdiffusion 633 -407 633 -407 0 cellNo=302
rlabel pdiffusion 640 -407 640 -407 0 feedthrough
rlabel pdiffusion 647 -407 647 -407 0 feedthrough
rlabel pdiffusion 654 -407 654 -407 0 cellNo=238
rlabel pdiffusion 661 -407 661 -407 0 feedthrough
rlabel pdiffusion 668 -407 668 -407 0 feedthrough
rlabel pdiffusion 717 -407 717 -407 0 feedthrough
rlabel pdiffusion 3 -472 3 -472 0 cellNo=114
rlabel pdiffusion 10 -472 10 -472 0 feedthrough
rlabel pdiffusion 17 -472 17 -472 0 feedthrough
rlabel pdiffusion 24 -472 24 -472 0 cellNo=520
rlabel pdiffusion 31 -472 31 -472 0 feedthrough
rlabel pdiffusion 38 -472 38 -472 0 feedthrough
rlabel pdiffusion 45 -472 45 -472 0 feedthrough
rlabel pdiffusion 52 -472 52 -472 0 feedthrough
rlabel pdiffusion 59 -472 59 -472 0 feedthrough
rlabel pdiffusion 66 -472 66 -472 0 cellNo=413
rlabel pdiffusion 73 -472 73 -472 0 cellNo=537
rlabel pdiffusion 80 -472 80 -472 0 cellNo=206
rlabel pdiffusion 87 -472 87 -472 0 feedthrough
rlabel pdiffusion 94 -472 94 -472 0 feedthrough
rlabel pdiffusion 101 -472 101 -472 0 cellNo=386
rlabel pdiffusion 108 -472 108 -472 0 feedthrough
rlabel pdiffusion 115 -472 115 -472 0 feedthrough
rlabel pdiffusion 122 -472 122 -472 0 feedthrough
rlabel pdiffusion 129 -472 129 -472 0 feedthrough
rlabel pdiffusion 136 -472 136 -472 0 feedthrough
rlabel pdiffusion 143 -472 143 -472 0 cellNo=351
rlabel pdiffusion 150 -472 150 -472 0 feedthrough
rlabel pdiffusion 157 -472 157 -472 0 feedthrough
rlabel pdiffusion 164 -472 164 -472 0 cellNo=451
rlabel pdiffusion 171 -472 171 -472 0 cellNo=1
rlabel pdiffusion 178 -472 178 -472 0 cellNo=189
rlabel pdiffusion 185 -472 185 -472 0 cellNo=359
rlabel pdiffusion 192 -472 192 -472 0 cellNo=65
rlabel pdiffusion 199 -472 199 -472 0 feedthrough
rlabel pdiffusion 206 -472 206 -472 0 feedthrough
rlabel pdiffusion 213 -472 213 -472 0 feedthrough
rlabel pdiffusion 220 -472 220 -472 0 feedthrough
rlabel pdiffusion 227 -472 227 -472 0 feedthrough
rlabel pdiffusion 234 -472 234 -472 0 feedthrough
rlabel pdiffusion 241 -472 241 -472 0 feedthrough
rlabel pdiffusion 248 -472 248 -472 0 feedthrough
rlabel pdiffusion 255 -472 255 -472 0 feedthrough
rlabel pdiffusion 262 -472 262 -472 0 feedthrough
rlabel pdiffusion 269 -472 269 -472 0 feedthrough
rlabel pdiffusion 276 -472 276 -472 0 feedthrough
rlabel pdiffusion 283 -472 283 -472 0 feedthrough
rlabel pdiffusion 290 -472 290 -472 0 feedthrough
rlabel pdiffusion 297 -472 297 -472 0 feedthrough
rlabel pdiffusion 304 -472 304 -472 0 feedthrough
rlabel pdiffusion 311 -472 311 -472 0 cellNo=122
rlabel pdiffusion 318 -472 318 -472 0 feedthrough
rlabel pdiffusion 325 -472 325 -472 0 feedthrough
rlabel pdiffusion 332 -472 332 -472 0 feedthrough
rlabel pdiffusion 339 -472 339 -472 0 feedthrough
rlabel pdiffusion 346 -472 346 -472 0 feedthrough
rlabel pdiffusion 353 -472 353 -472 0 feedthrough
rlabel pdiffusion 360 -472 360 -472 0 cellNo=383
rlabel pdiffusion 367 -472 367 -472 0 cellNo=179
rlabel pdiffusion 374 -472 374 -472 0 feedthrough
rlabel pdiffusion 381 -472 381 -472 0 cellNo=306
rlabel pdiffusion 388 -472 388 -472 0 cellNo=85
rlabel pdiffusion 395 -472 395 -472 0 cellNo=112
rlabel pdiffusion 402 -472 402 -472 0 feedthrough
rlabel pdiffusion 409 -472 409 -472 0 cellNo=72
rlabel pdiffusion 416 -472 416 -472 0 cellNo=137
rlabel pdiffusion 423 -472 423 -472 0 cellNo=15
rlabel pdiffusion 430 -472 430 -472 0 cellNo=128
rlabel pdiffusion 437 -472 437 -472 0 cellNo=197
rlabel pdiffusion 444 -472 444 -472 0 cellNo=98
rlabel pdiffusion 451 -472 451 -472 0 cellNo=147
rlabel pdiffusion 458 -472 458 -472 0 feedthrough
rlabel pdiffusion 465 -472 465 -472 0 feedthrough
rlabel pdiffusion 472 -472 472 -472 0 feedthrough
rlabel pdiffusion 479 -472 479 -472 0 feedthrough
rlabel pdiffusion 486 -472 486 -472 0 feedthrough
rlabel pdiffusion 493 -472 493 -472 0 feedthrough
rlabel pdiffusion 500 -472 500 -472 0 feedthrough
rlabel pdiffusion 507 -472 507 -472 0 feedthrough
rlabel pdiffusion 514 -472 514 -472 0 feedthrough
rlabel pdiffusion 521 -472 521 -472 0 feedthrough
rlabel pdiffusion 528 -472 528 -472 0 feedthrough
rlabel pdiffusion 535 -472 535 -472 0 feedthrough
rlabel pdiffusion 542 -472 542 -472 0 feedthrough
rlabel pdiffusion 549 -472 549 -472 0 feedthrough
rlabel pdiffusion 556 -472 556 -472 0 feedthrough
rlabel pdiffusion 563 -472 563 -472 0 feedthrough
rlabel pdiffusion 570 -472 570 -472 0 feedthrough
rlabel pdiffusion 577 -472 577 -472 0 feedthrough
rlabel pdiffusion 584 -472 584 -472 0 feedthrough
rlabel pdiffusion 591 -472 591 -472 0 feedthrough
rlabel pdiffusion 598 -472 598 -472 0 feedthrough
rlabel pdiffusion 605 -472 605 -472 0 feedthrough
rlabel pdiffusion 612 -472 612 -472 0 feedthrough
rlabel pdiffusion 626 -472 626 -472 0 feedthrough
rlabel pdiffusion 633 -472 633 -472 0 feedthrough
rlabel pdiffusion 640 -472 640 -472 0 feedthrough
rlabel pdiffusion 647 -472 647 -472 0 feedthrough
rlabel pdiffusion 654 -472 654 -472 0 feedthrough
rlabel pdiffusion 668 -472 668 -472 0 feedthrough
rlabel pdiffusion 675 -472 675 -472 0 feedthrough
rlabel pdiffusion 682 -472 682 -472 0 feedthrough
rlabel pdiffusion 689 -472 689 -472 0 feedthrough
rlabel pdiffusion 696 -472 696 -472 0 feedthrough
rlabel pdiffusion 703 -472 703 -472 0 feedthrough
rlabel pdiffusion 710 -472 710 -472 0 cellNo=560
rlabel pdiffusion 717 -472 717 -472 0 cellNo=73
rlabel pdiffusion 724 -472 724 -472 0 feedthrough
rlabel pdiffusion 731 -472 731 -472 0 feedthrough
rlabel pdiffusion 3 -557 3 -557 0 cellNo=235
rlabel pdiffusion 10 -557 10 -557 0 cellNo=384
rlabel pdiffusion 17 -557 17 -557 0 cellNo=720
rlabel pdiffusion 24 -557 24 -557 0 feedthrough
rlabel pdiffusion 31 -557 31 -557 0 cellNo=620
rlabel pdiffusion 38 -557 38 -557 0 cellNo=117
rlabel pdiffusion 45 -557 45 -557 0 feedthrough
rlabel pdiffusion 52 -557 52 -557 0 cellNo=185
rlabel pdiffusion 59 -557 59 -557 0 cellNo=164
rlabel pdiffusion 66 -557 66 -557 0 cellNo=36
rlabel pdiffusion 73 -557 73 -557 0 cellNo=552
rlabel pdiffusion 80 -557 80 -557 0 feedthrough
rlabel pdiffusion 87 -557 87 -557 0 feedthrough
rlabel pdiffusion 94 -557 94 -557 0 feedthrough
rlabel pdiffusion 101 -557 101 -557 0 cellNo=304
rlabel pdiffusion 108 -557 108 -557 0 feedthrough
rlabel pdiffusion 115 -557 115 -557 0 feedthrough
rlabel pdiffusion 122 -557 122 -557 0 cellNo=305
rlabel pdiffusion 129 -557 129 -557 0 feedthrough
rlabel pdiffusion 136 -557 136 -557 0 feedthrough
rlabel pdiffusion 143 -557 143 -557 0 cellNo=403
rlabel pdiffusion 150 -557 150 -557 0 cellNo=66
rlabel pdiffusion 157 -557 157 -557 0 feedthrough
rlabel pdiffusion 164 -557 164 -557 0 cellNo=674
rlabel pdiffusion 171 -557 171 -557 0 feedthrough
rlabel pdiffusion 178 -557 178 -557 0 cellNo=483
rlabel pdiffusion 185 -557 185 -557 0 cellNo=632
rlabel pdiffusion 192 -557 192 -557 0 feedthrough
rlabel pdiffusion 199 -557 199 -557 0 feedthrough
rlabel pdiffusion 206 -557 206 -557 0 feedthrough
rlabel pdiffusion 213 -557 213 -557 0 cellNo=567
rlabel pdiffusion 220 -557 220 -557 0 feedthrough
rlabel pdiffusion 227 -557 227 -557 0 feedthrough
rlabel pdiffusion 234 -557 234 -557 0 cellNo=641
rlabel pdiffusion 241 -557 241 -557 0 cellNo=9
rlabel pdiffusion 248 -557 248 -557 0 feedthrough
rlabel pdiffusion 255 -557 255 -557 0 feedthrough
rlabel pdiffusion 262 -557 262 -557 0 feedthrough
rlabel pdiffusion 269 -557 269 -557 0 feedthrough
rlabel pdiffusion 276 -557 276 -557 0 feedthrough
rlabel pdiffusion 283 -557 283 -557 0 feedthrough
rlabel pdiffusion 290 -557 290 -557 0 feedthrough
rlabel pdiffusion 297 -557 297 -557 0 feedthrough
rlabel pdiffusion 304 -557 304 -557 0 cellNo=104
rlabel pdiffusion 311 -557 311 -557 0 feedthrough
rlabel pdiffusion 318 -557 318 -557 0 cellNo=547
rlabel pdiffusion 325 -557 325 -557 0 feedthrough
rlabel pdiffusion 332 -557 332 -557 0 feedthrough
rlabel pdiffusion 339 -557 339 -557 0 feedthrough
rlabel pdiffusion 346 -557 346 -557 0 feedthrough
rlabel pdiffusion 353 -557 353 -557 0 feedthrough
rlabel pdiffusion 360 -557 360 -557 0 feedthrough
rlabel pdiffusion 367 -557 367 -557 0 cellNo=592
rlabel pdiffusion 374 -557 374 -557 0 feedthrough
rlabel pdiffusion 381 -557 381 -557 0 cellNo=95
rlabel pdiffusion 388 -557 388 -557 0 feedthrough
rlabel pdiffusion 395 -557 395 -557 0 cellNo=466
rlabel pdiffusion 402 -557 402 -557 0 feedthrough
rlabel pdiffusion 409 -557 409 -557 0 feedthrough
rlabel pdiffusion 416 -557 416 -557 0 feedthrough
rlabel pdiffusion 423 -557 423 -557 0 cellNo=504
rlabel pdiffusion 430 -557 430 -557 0 cellNo=395
rlabel pdiffusion 437 -557 437 -557 0 feedthrough
rlabel pdiffusion 444 -557 444 -557 0 cellNo=462
rlabel pdiffusion 451 -557 451 -557 0 feedthrough
rlabel pdiffusion 458 -557 458 -557 0 feedthrough
rlabel pdiffusion 465 -557 465 -557 0 feedthrough
rlabel pdiffusion 472 -557 472 -557 0 feedthrough
rlabel pdiffusion 479 -557 479 -557 0 feedthrough
rlabel pdiffusion 486 -557 486 -557 0 feedthrough
rlabel pdiffusion 493 -557 493 -557 0 feedthrough
rlabel pdiffusion 500 -557 500 -557 0 feedthrough
rlabel pdiffusion 507 -557 507 -557 0 feedthrough
rlabel pdiffusion 514 -557 514 -557 0 feedthrough
rlabel pdiffusion 521 -557 521 -557 0 feedthrough
rlabel pdiffusion 528 -557 528 -557 0 feedthrough
rlabel pdiffusion 535 -557 535 -557 0 feedthrough
rlabel pdiffusion 542 -557 542 -557 0 feedthrough
rlabel pdiffusion 549 -557 549 -557 0 feedthrough
rlabel pdiffusion 556 -557 556 -557 0 feedthrough
rlabel pdiffusion 563 -557 563 -557 0 feedthrough
rlabel pdiffusion 570 -557 570 -557 0 feedthrough
rlabel pdiffusion 577 -557 577 -557 0 feedthrough
rlabel pdiffusion 584 -557 584 -557 0 feedthrough
rlabel pdiffusion 591 -557 591 -557 0 feedthrough
rlabel pdiffusion 598 -557 598 -557 0 feedthrough
rlabel pdiffusion 605 -557 605 -557 0 feedthrough
rlabel pdiffusion 612 -557 612 -557 0 feedthrough
rlabel pdiffusion 619 -557 619 -557 0 feedthrough
rlabel pdiffusion 626 -557 626 -557 0 feedthrough
rlabel pdiffusion 633 -557 633 -557 0 feedthrough
rlabel pdiffusion 640 -557 640 -557 0 feedthrough
rlabel pdiffusion 647 -557 647 -557 0 feedthrough
rlabel pdiffusion 654 -557 654 -557 0 feedthrough
rlabel pdiffusion 661 -557 661 -557 0 feedthrough
rlabel pdiffusion 668 -557 668 -557 0 feedthrough
rlabel pdiffusion 675 -557 675 -557 0 feedthrough
rlabel pdiffusion 682 -557 682 -557 0 feedthrough
rlabel pdiffusion 689 -557 689 -557 0 feedthrough
rlabel pdiffusion 696 -557 696 -557 0 feedthrough
rlabel pdiffusion 703 -557 703 -557 0 feedthrough
rlabel pdiffusion 710 -557 710 -557 0 feedthrough
rlabel pdiffusion 717 -557 717 -557 0 feedthrough
rlabel pdiffusion 724 -557 724 -557 0 feedthrough
rlabel pdiffusion 731 -557 731 -557 0 feedthrough
rlabel pdiffusion 738 -557 738 -557 0 feedthrough
rlabel pdiffusion 745 -557 745 -557 0 feedthrough
rlabel pdiffusion 752 -557 752 -557 0 feedthrough
rlabel pdiffusion 780 -557 780 -557 0 feedthrough
rlabel pdiffusion 3 -650 3 -650 0 cellNo=381
rlabel pdiffusion 10 -650 10 -650 0 cellNo=441
rlabel pdiffusion 17 -650 17 -650 0 feedthrough
rlabel pdiffusion 24 -650 24 -650 0 feedthrough
rlabel pdiffusion 31 -650 31 -650 0 cellNo=94
rlabel pdiffusion 38 -650 38 -650 0 cellNo=320
rlabel pdiffusion 45 -650 45 -650 0 cellNo=307
rlabel pdiffusion 52 -650 52 -650 0 feedthrough
rlabel pdiffusion 59 -650 59 -650 0 feedthrough
rlabel pdiffusion 66 -650 66 -650 0 feedthrough
rlabel pdiffusion 73 -650 73 -650 0 feedthrough
rlabel pdiffusion 80 -650 80 -650 0 feedthrough
rlabel pdiffusion 87 -650 87 -650 0 feedthrough
rlabel pdiffusion 94 -650 94 -650 0 cellNo=303
rlabel pdiffusion 101 -650 101 -650 0 feedthrough
rlabel pdiffusion 108 -650 108 -650 0 cellNo=270
rlabel pdiffusion 115 -650 115 -650 0 cellNo=214
rlabel pdiffusion 122 -650 122 -650 0 cellNo=250
rlabel pdiffusion 129 -650 129 -650 0 cellNo=135
rlabel pdiffusion 136 -650 136 -650 0 feedthrough
rlabel pdiffusion 143 -650 143 -650 0 cellNo=529
rlabel pdiffusion 150 -650 150 -650 0 cellNo=138
rlabel pdiffusion 157 -650 157 -650 0 feedthrough
rlabel pdiffusion 164 -650 164 -650 0 cellNo=83
rlabel pdiffusion 171 -650 171 -650 0 feedthrough
rlabel pdiffusion 178 -650 178 -650 0 feedthrough
rlabel pdiffusion 185 -650 185 -650 0 cellNo=165
rlabel pdiffusion 192 -650 192 -650 0 feedthrough
rlabel pdiffusion 199 -650 199 -650 0 feedthrough
rlabel pdiffusion 206 -650 206 -650 0 feedthrough
rlabel pdiffusion 213 -650 213 -650 0 feedthrough
rlabel pdiffusion 220 -650 220 -650 0 feedthrough
rlabel pdiffusion 227 -650 227 -650 0 feedthrough
rlabel pdiffusion 234 -650 234 -650 0 feedthrough
rlabel pdiffusion 241 -650 241 -650 0 feedthrough
rlabel pdiffusion 248 -650 248 -650 0 feedthrough
rlabel pdiffusion 255 -650 255 -650 0 feedthrough
rlabel pdiffusion 262 -650 262 -650 0 feedthrough
rlabel pdiffusion 269 -650 269 -650 0 feedthrough
rlabel pdiffusion 276 -650 276 -650 0 cellNo=692
rlabel pdiffusion 283 -650 283 -650 0 feedthrough
rlabel pdiffusion 290 -650 290 -650 0 cellNo=260
rlabel pdiffusion 297 -650 297 -650 0 feedthrough
rlabel pdiffusion 304 -650 304 -650 0 feedthrough
rlabel pdiffusion 311 -650 311 -650 0 feedthrough
rlabel pdiffusion 318 -650 318 -650 0 feedthrough
rlabel pdiffusion 325 -650 325 -650 0 feedthrough
rlabel pdiffusion 332 -650 332 -650 0 feedthrough
rlabel pdiffusion 339 -650 339 -650 0 feedthrough
rlabel pdiffusion 346 -650 346 -650 0 cellNo=676
rlabel pdiffusion 353 -650 353 -650 0 cellNo=263
rlabel pdiffusion 360 -650 360 -650 0 feedthrough
rlabel pdiffusion 367 -650 367 -650 0 cellNo=269
rlabel pdiffusion 374 -650 374 -650 0 feedthrough
rlabel pdiffusion 381 -650 381 -650 0 feedthrough
rlabel pdiffusion 388 -650 388 -650 0 cellNo=388
rlabel pdiffusion 395 -650 395 -650 0 cellNo=314
rlabel pdiffusion 402 -650 402 -650 0 feedthrough
rlabel pdiffusion 409 -650 409 -650 0 cellNo=27
rlabel pdiffusion 416 -650 416 -650 0 cellNo=432
rlabel pdiffusion 423 -650 423 -650 0 cellNo=142
rlabel pdiffusion 430 -650 430 -650 0 feedthrough
rlabel pdiffusion 437 -650 437 -650 0 feedthrough
rlabel pdiffusion 444 -650 444 -650 0 cellNo=255
rlabel pdiffusion 451 -650 451 -650 0 feedthrough
rlabel pdiffusion 458 -650 458 -650 0 feedthrough
rlabel pdiffusion 465 -650 465 -650 0 feedthrough
rlabel pdiffusion 472 -650 472 -650 0 feedthrough
rlabel pdiffusion 479 -650 479 -650 0 feedthrough
rlabel pdiffusion 486 -650 486 -650 0 feedthrough
rlabel pdiffusion 500 -650 500 -650 0 feedthrough
rlabel pdiffusion 507 -650 507 -650 0 feedthrough
rlabel pdiffusion 514 -650 514 -650 0 cellNo=338
rlabel pdiffusion 521 -650 521 -650 0 feedthrough
rlabel pdiffusion 528 -650 528 -650 0 feedthrough
rlabel pdiffusion 535 -650 535 -650 0 feedthrough
rlabel pdiffusion 542 -650 542 -650 0 feedthrough
rlabel pdiffusion 549 -650 549 -650 0 feedthrough
rlabel pdiffusion 556 -650 556 -650 0 feedthrough
rlabel pdiffusion 563 -650 563 -650 0 feedthrough
rlabel pdiffusion 570 -650 570 -650 0 feedthrough
rlabel pdiffusion 577 -650 577 -650 0 feedthrough
rlabel pdiffusion 584 -650 584 -650 0 feedthrough
rlabel pdiffusion 591 -650 591 -650 0 feedthrough
rlabel pdiffusion 598 -650 598 -650 0 feedthrough
rlabel pdiffusion 605 -650 605 -650 0 feedthrough
rlabel pdiffusion 612 -650 612 -650 0 feedthrough
rlabel pdiffusion 619 -650 619 -650 0 feedthrough
rlabel pdiffusion 626 -650 626 -650 0 feedthrough
rlabel pdiffusion 633 -650 633 -650 0 feedthrough
rlabel pdiffusion 640 -650 640 -650 0 feedthrough
rlabel pdiffusion 647 -650 647 -650 0 feedthrough
rlabel pdiffusion 654 -650 654 -650 0 feedthrough
rlabel pdiffusion 661 -650 661 -650 0 cellNo=576
rlabel pdiffusion 668 -650 668 -650 0 feedthrough
rlabel pdiffusion 675 -650 675 -650 0 feedthrough
rlabel pdiffusion 682 -650 682 -650 0 feedthrough
rlabel pdiffusion 689 -650 689 -650 0 feedthrough
rlabel pdiffusion 696 -650 696 -650 0 feedthrough
rlabel pdiffusion 703 -650 703 -650 0 feedthrough
rlabel pdiffusion 710 -650 710 -650 0 feedthrough
rlabel pdiffusion 717 -650 717 -650 0 feedthrough
rlabel pdiffusion 724 -650 724 -650 0 feedthrough
rlabel pdiffusion 731 -650 731 -650 0 feedthrough
rlabel pdiffusion 738 -650 738 -650 0 feedthrough
rlabel pdiffusion 808 -650 808 -650 0 feedthrough
rlabel pdiffusion 3 -731 3 -731 0 cellNo=411
rlabel pdiffusion 10 -731 10 -731 0 feedthrough
rlabel pdiffusion 17 -731 17 -731 0 feedthrough
rlabel pdiffusion 24 -731 24 -731 0 feedthrough
rlabel pdiffusion 31 -731 31 -731 0 feedthrough
rlabel pdiffusion 38 -731 38 -731 0 feedthrough
rlabel pdiffusion 45 -731 45 -731 0 feedthrough
rlabel pdiffusion 52 -731 52 -731 0 cellNo=573
rlabel pdiffusion 59 -731 59 -731 0 cellNo=207
rlabel pdiffusion 66 -731 66 -731 0 cellNo=539
rlabel pdiffusion 73 -731 73 -731 0 cellNo=38
rlabel pdiffusion 80 -731 80 -731 0 feedthrough
rlabel pdiffusion 87 -731 87 -731 0 feedthrough
rlabel pdiffusion 94 -731 94 -731 0 cellNo=706
rlabel pdiffusion 101 -731 101 -731 0 feedthrough
rlabel pdiffusion 108 -731 108 -731 0 feedthrough
rlabel pdiffusion 115 -731 115 -731 0 cellNo=694
rlabel pdiffusion 122 -731 122 -731 0 cellNo=19
rlabel pdiffusion 129 -731 129 -731 0 feedthrough
rlabel pdiffusion 136 -731 136 -731 0 feedthrough
rlabel pdiffusion 143 -731 143 -731 0 feedthrough
rlabel pdiffusion 150 -731 150 -731 0 feedthrough
rlabel pdiffusion 157 -731 157 -731 0 cellNo=658
rlabel pdiffusion 164 -731 164 -731 0 cellNo=609
rlabel pdiffusion 171 -731 171 -731 0 cellNo=509
rlabel pdiffusion 178 -731 178 -731 0 feedthrough
rlabel pdiffusion 185 -731 185 -731 0 feedthrough
rlabel pdiffusion 192 -731 192 -731 0 feedthrough
rlabel pdiffusion 199 -731 199 -731 0 feedthrough
rlabel pdiffusion 206 -731 206 -731 0 feedthrough
rlabel pdiffusion 213 -731 213 -731 0 feedthrough
rlabel pdiffusion 220 -731 220 -731 0 feedthrough
rlabel pdiffusion 227 -731 227 -731 0 feedthrough
rlabel pdiffusion 234 -731 234 -731 0 cellNo=40
rlabel pdiffusion 241 -731 241 -731 0 cellNo=103
rlabel pdiffusion 248 -731 248 -731 0 feedthrough
rlabel pdiffusion 255 -731 255 -731 0 cellNo=481
rlabel pdiffusion 262 -731 262 -731 0 feedthrough
rlabel pdiffusion 269 -731 269 -731 0 feedthrough
rlabel pdiffusion 276 -731 276 -731 0 feedthrough
rlabel pdiffusion 283 -731 283 -731 0 feedthrough
rlabel pdiffusion 290 -731 290 -731 0 cellNo=508
rlabel pdiffusion 297 -731 297 -731 0 feedthrough
rlabel pdiffusion 304 -731 304 -731 0 feedthrough
rlabel pdiffusion 311 -731 311 -731 0 feedthrough
rlabel pdiffusion 318 -731 318 -731 0 feedthrough
rlabel pdiffusion 325 -731 325 -731 0 feedthrough
rlabel pdiffusion 332 -731 332 -731 0 cellNo=71
rlabel pdiffusion 339 -731 339 -731 0 feedthrough
rlabel pdiffusion 346 -731 346 -731 0 feedthrough
rlabel pdiffusion 353 -731 353 -731 0 feedthrough
rlabel pdiffusion 360 -731 360 -731 0 feedthrough
rlabel pdiffusion 367 -731 367 -731 0 cellNo=62
rlabel pdiffusion 374 -731 374 -731 0 feedthrough
rlabel pdiffusion 381 -731 381 -731 0 feedthrough
rlabel pdiffusion 388 -731 388 -731 0 feedthrough
rlabel pdiffusion 395 -731 395 -731 0 cellNo=440
rlabel pdiffusion 402 -731 402 -731 0 feedthrough
rlabel pdiffusion 409 -731 409 -731 0 cellNo=498
rlabel pdiffusion 416 -731 416 -731 0 feedthrough
rlabel pdiffusion 423 -731 423 -731 0 feedthrough
rlabel pdiffusion 430 -731 430 -731 0 cellNo=430
rlabel pdiffusion 437 -731 437 -731 0 cellNo=399
rlabel pdiffusion 444 -731 444 -731 0 feedthrough
rlabel pdiffusion 451 -731 451 -731 0 cellNo=279
rlabel pdiffusion 458 -731 458 -731 0 feedthrough
rlabel pdiffusion 465 -731 465 -731 0 cellNo=648
rlabel pdiffusion 472 -731 472 -731 0 cellNo=132
rlabel pdiffusion 479 -731 479 -731 0 feedthrough
rlabel pdiffusion 486 -731 486 -731 0 feedthrough
rlabel pdiffusion 493 -731 493 -731 0 feedthrough
rlabel pdiffusion 500 -731 500 -731 0 feedthrough
rlabel pdiffusion 507 -731 507 -731 0 feedthrough
rlabel pdiffusion 514 -731 514 -731 0 feedthrough
rlabel pdiffusion 521 -731 521 -731 0 feedthrough
rlabel pdiffusion 528 -731 528 -731 0 feedthrough
rlabel pdiffusion 535 -731 535 -731 0 feedthrough
rlabel pdiffusion 542 -731 542 -731 0 feedthrough
rlabel pdiffusion 549 -731 549 -731 0 feedthrough
rlabel pdiffusion 556 -731 556 -731 0 feedthrough
rlabel pdiffusion 563 -731 563 -731 0 feedthrough
rlabel pdiffusion 570 -731 570 -731 0 feedthrough
rlabel pdiffusion 577 -731 577 -731 0 feedthrough
rlabel pdiffusion 584 -731 584 -731 0 feedthrough
rlabel pdiffusion 591 -731 591 -731 0 feedthrough
rlabel pdiffusion 598 -731 598 -731 0 cellNo=202
rlabel pdiffusion 605 -731 605 -731 0 feedthrough
rlabel pdiffusion 612 -731 612 -731 0 feedthrough
rlabel pdiffusion 619 -731 619 -731 0 feedthrough
rlabel pdiffusion 626 -731 626 -731 0 feedthrough
rlabel pdiffusion 633 -731 633 -731 0 feedthrough
rlabel pdiffusion 640 -731 640 -731 0 feedthrough
rlabel pdiffusion 647 -731 647 -731 0 feedthrough
rlabel pdiffusion 654 -731 654 -731 0 feedthrough
rlabel pdiffusion 661 -731 661 -731 0 feedthrough
rlabel pdiffusion 668 -731 668 -731 0 feedthrough
rlabel pdiffusion 675 -731 675 -731 0 feedthrough
rlabel pdiffusion 682 -731 682 -731 0 feedthrough
rlabel pdiffusion 689 -731 689 -731 0 feedthrough
rlabel pdiffusion 696 -731 696 -731 0 feedthrough
rlabel pdiffusion 703 -731 703 -731 0 feedthrough
rlabel pdiffusion 710 -731 710 -731 0 feedthrough
rlabel pdiffusion 717 -731 717 -731 0 feedthrough
rlabel pdiffusion 724 -731 724 -731 0 feedthrough
rlabel pdiffusion 731 -731 731 -731 0 feedthrough
rlabel pdiffusion 738 -731 738 -731 0 feedthrough
rlabel pdiffusion 745 -731 745 -731 0 feedthrough
rlabel pdiffusion 752 -731 752 -731 0 feedthrough
rlabel pdiffusion 759 -731 759 -731 0 feedthrough
rlabel pdiffusion 766 -731 766 -731 0 feedthrough
rlabel pdiffusion 773 -731 773 -731 0 feedthrough
rlabel pdiffusion 780 -731 780 -731 0 feedthrough
rlabel pdiffusion 787 -731 787 -731 0 feedthrough
rlabel pdiffusion 794 -731 794 -731 0 feedthrough
rlabel pdiffusion 801 -731 801 -731 0 feedthrough
rlabel pdiffusion 808 -731 808 -731 0 feedthrough
rlabel pdiffusion 815 -731 815 -731 0 cellNo=323
rlabel pdiffusion 822 -731 822 -731 0 cellNo=354
rlabel pdiffusion 829 -731 829 -731 0 feedthrough
rlabel pdiffusion 3 -820 3 -820 0 cellNo=554
rlabel pdiffusion 10 -820 10 -820 0 feedthrough
rlabel pdiffusion 17 -820 17 -820 0 cellNo=587
rlabel pdiffusion 24 -820 24 -820 0 feedthrough
rlabel pdiffusion 31 -820 31 -820 0 feedthrough
rlabel pdiffusion 38 -820 38 -820 0 cellNo=31
rlabel pdiffusion 45 -820 45 -820 0 cellNo=60
rlabel pdiffusion 52 -820 52 -820 0 cellNo=394
rlabel pdiffusion 59 -820 59 -820 0 feedthrough
rlabel pdiffusion 66 -820 66 -820 0 cellNo=68
rlabel pdiffusion 73 -820 73 -820 0 cellNo=367
rlabel pdiffusion 80 -820 80 -820 0 cellNo=181
rlabel pdiffusion 87 -820 87 -820 0 feedthrough
rlabel pdiffusion 94 -820 94 -820 0 cellNo=453
rlabel pdiffusion 101 -820 101 -820 0 feedthrough
rlabel pdiffusion 108 -820 108 -820 0 feedthrough
rlabel pdiffusion 115 -820 115 -820 0 feedthrough
rlabel pdiffusion 122 -820 122 -820 0 feedthrough
rlabel pdiffusion 129 -820 129 -820 0 feedthrough
rlabel pdiffusion 136 -820 136 -820 0 feedthrough
rlabel pdiffusion 143 -820 143 -820 0 feedthrough
rlabel pdiffusion 150 -820 150 -820 0 cellNo=16
rlabel pdiffusion 157 -820 157 -820 0 feedthrough
rlabel pdiffusion 164 -820 164 -820 0 feedthrough
rlabel pdiffusion 171 -820 171 -820 0 feedthrough
rlabel pdiffusion 178 -820 178 -820 0 feedthrough
rlabel pdiffusion 185 -820 185 -820 0 cellNo=90
rlabel pdiffusion 192 -820 192 -820 0 feedthrough
rlabel pdiffusion 199 -820 199 -820 0 feedthrough
rlabel pdiffusion 206 -820 206 -820 0 feedthrough
rlabel pdiffusion 213 -820 213 -820 0 feedthrough
rlabel pdiffusion 220 -820 220 -820 0 feedthrough
rlabel pdiffusion 227 -820 227 -820 0 feedthrough
rlabel pdiffusion 234 -820 234 -820 0 feedthrough
rlabel pdiffusion 241 -820 241 -820 0 feedthrough
rlabel pdiffusion 248 -820 248 -820 0 feedthrough
rlabel pdiffusion 255 -820 255 -820 0 feedthrough
rlabel pdiffusion 262 -820 262 -820 0 feedthrough
rlabel pdiffusion 269 -820 269 -820 0 cellNo=352
rlabel pdiffusion 276 -820 276 -820 0 feedthrough
rlabel pdiffusion 283 -820 283 -820 0 feedthrough
rlabel pdiffusion 290 -820 290 -820 0 feedthrough
rlabel pdiffusion 297 -820 297 -820 0 feedthrough
rlabel pdiffusion 304 -820 304 -820 0 cellNo=347
rlabel pdiffusion 311 -820 311 -820 0 feedthrough
rlabel pdiffusion 318 -820 318 -820 0 feedthrough
rlabel pdiffusion 325 -820 325 -820 0 feedthrough
rlabel pdiffusion 332 -820 332 -820 0 cellNo=478
rlabel pdiffusion 339 -820 339 -820 0 cellNo=665
rlabel pdiffusion 346 -820 346 -820 0 cellNo=672
rlabel pdiffusion 353 -820 353 -820 0 cellNo=77
rlabel pdiffusion 360 -820 360 -820 0 feedthrough
rlabel pdiffusion 367 -820 367 -820 0 cellNo=447
rlabel pdiffusion 374 -820 374 -820 0 feedthrough
rlabel pdiffusion 381 -820 381 -820 0 cellNo=418
rlabel pdiffusion 388 -820 388 -820 0 cellNo=312
rlabel pdiffusion 395 -820 395 -820 0 feedthrough
rlabel pdiffusion 402 -820 402 -820 0 cellNo=109
rlabel pdiffusion 409 -820 409 -820 0 feedthrough
rlabel pdiffusion 416 -820 416 -820 0 feedthrough
rlabel pdiffusion 423 -820 423 -820 0 feedthrough
rlabel pdiffusion 430 -820 430 -820 0 cellNo=215
rlabel pdiffusion 437 -820 437 -820 0 cellNo=627
rlabel pdiffusion 444 -820 444 -820 0 cellNo=345
rlabel pdiffusion 451 -820 451 -820 0 cellNo=154
rlabel pdiffusion 458 -820 458 -820 0 feedthrough
rlabel pdiffusion 465 -820 465 -820 0 feedthrough
rlabel pdiffusion 472 -820 472 -820 0 feedthrough
rlabel pdiffusion 479 -820 479 -820 0 feedthrough
rlabel pdiffusion 486 -820 486 -820 0 feedthrough
rlabel pdiffusion 493 -820 493 -820 0 feedthrough
rlabel pdiffusion 500 -820 500 -820 0 feedthrough
rlabel pdiffusion 507 -820 507 -820 0 feedthrough
rlabel pdiffusion 514 -820 514 -820 0 feedthrough
rlabel pdiffusion 521 -820 521 -820 0 feedthrough
rlabel pdiffusion 528 -820 528 -820 0 feedthrough
rlabel pdiffusion 535 -820 535 -820 0 feedthrough
rlabel pdiffusion 542 -820 542 -820 0 feedthrough
rlabel pdiffusion 549 -820 549 -820 0 feedthrough
rlabel pdiffusion 556 -820 556 -820 0 cellNo=516
rlabel pdiffusion 563 -820 563 -820 0 feedthrough
rlabel pdiffusion 570 -820 570 -820 0 feedthrough
rlabel pdiffusion 577 -820 577 -820 0 feedthrough
rlabel pdiffusion 584 -820 584 -820 0 feedthrough
rlabel pdiffusion 591 -820 591 -820 0 cellNo=273
rlabel pdiffusion 598 -820 598 -820 0 feedthrough
rlabel pdiffusion 605 -820 605 -820 0 feedthrough
rlabel pdiffusion 612 -820 612 -820 0 feedthrough
rlabel pdiffusion 619 -820 619 -820 0 feedthrough
rlabel pdiffusion 626 -820 626 -820 0 feedthrough
rlabel pdiffusion 633 -820 633 -820 0 feedthrough
rlabel pdiffusion 640 -820 640 -820 0 feedthrough
rlabel pdiffusion 647 -820 647 -820 0 feedthrough
rlabel pdiffusion 654 -820 654 -820 0 feedthrough
rlabel pdiffusion 661 -820 661 -820 0 feedthrough
rlabel pdiffusion 668 -820 668 -820 0 feedthrough
rlabel pdiffusion 675 -820 675 -820 0 feedthrough
rlabel pdiffusion 682 -820 682 -820 0 feedthrough
rlabel pdiffusion 689 -820 689 -820 0 feedthrough
rlabel pdiffusion 696 -820 696 -820 0 feedthrough
rlabel pdiffusion 703 -820 703 -820 0 feedthrough
rlabel pdiffusion 710 -820 710 -820 0 feedthrough
rlabel pdiffusion 717 -820 717 -820 0 feedthrough
rlabel pdiffusion 724 -820 724 -820 0 feedthrough
rlabel pdiffusion 731 -820 731 -820 0 feedthrough
rlabel pdiffusion 738 -820 738 -820 0 feedthrough
rlabel pdiffusion 745 -820 745 -820 0 feedthrough
rlabel pdiffusion 752 -820 752 -820 0 feedthrough
rlabel pdiffusion 759 -820 759 -820 0 feedthrough
rlabel pdiffusion 766 -820 766 -820 0 feedthrough
rlabel pdiffusion 773 -820 773 -820 0 feedthrough
rlabel pdiffusion 780 -820 780 -820 0 feedthrough
rlabel pdiffusion 787 -820 787 -820 0 feedthrough
rlabel pdiffusion 794 -820 794 -820 0 feedthrough
rlabel pdiffusion 3 -905 3 -905 0 cellNo=591
rlabel pdiffusion 10 -905 10 -905 0 cellNo=419
rlabel pdiffusion 17 -905 17 -905 0 feedthrough
rlabel pdiffusion 24 -905 24 -905 0 cellNo=23
rlabel pdiffusion 31 -905 31 -905 0 feedthrough
rlabel pdiffusion 38 -905 38 -905 0 cellNo=225
rlabel pdiffusion 45 -905 45 -905 0 feedthrough
rlabel pdiffusion 52 -905 52 -905 0 cellNo=631
rlabel pdiffusion 59 -905 59 -905 0 feedthrough
rlabel pdiffusion 66 -905 66 -905 0 feedthrough
rlabel pdiffusion 73 -905 73 -905 0 feedthrough
rlabel pdiffusion 80 -905 80 -905 0 feedthrough
rlabel pdiffusion 87 -905 87 -905 0 feedthrough
rlabel pdiffusion 94 -905 94 -905 0 feedthrough
rlabel pdiffusion 101 -905 101 -905 0 cellNo=33
rlabel pdiffusion 108 -905 108 -905 0 feedthrough
rlabel pdiffusion 115 -905 115 -905 0 cellNo=317
rlabel pdiffusion 122 -905 122 -905 0 feedthrough
rlabel pdiffusion 129 -905 129 -905 0 feedthrough
rlabel pdiffusion 136 -905 136 -905 0 cellNo=259
rlabel pdiffusion 143 -905 143 -905 0 cellNo=275
rlabel pdiffusion 150 -905 150 -905 0 feedthrough
rlabel pdiffusion 157 -905 157 -905 0 feedthrough
rlabel pdiffusion 164 -905 164 -905 0 feedthrough
rlabel pdiffusion 171 -905 171 -905 0 cellNo=582
rlabel pdiffusion 178 -905 178 -905 0 cellNo=519
rlabel pdiffusion 185 -905 185 -905 0 feedthrough
rlabel pdiffusion 192 -905 192 -905 0 feedthrough
rlabel pdiffusion 199 -905 199 -905 0 feedthrough
rlabel pdiffusion 206 -905 206 -905 0 feedthrough
rlabel pdiffusion 213 -905 213 -905 0 feedthrough
rlabel pdiffusion 220 -905 220 -905 0 feedthrough
rlabel pdiffusion 227 -905 227 -905 0 feedthrough
rlabel pdiffusion 234 -905 234 -905 0 feedthrough
rlabel pdiffusion 241 -905 241 -905 0 feedthrough
rlabel pdiffusion 248 -905 248 -905 0 feedthrough
rlabel pdiffusion 255 -905 255 -905 0 cellNo=337
rlabel pdiffusion 262 -905 262 -905 0 feedthrough
rlabel pdiffusion 269 -905 269 -905 0 feedthrough
rlabel pdiffusion 276 -905 276 -905 0 cellNo=79
rlabel pdiffusion 283 -905 283 -905 0 cellNo=491
rlabel pdiffusion 290 -905 290 -905 0 cellNo=217
rlabel pdiffusion 297 -905 297 -905 0 cellNo=438
rlabel pdiffusion 304 -905 304 -905 0 cellNo=378
rlabel pdiffusion 311 -905 311 -905 0 feedthrough
rlabel pdiffusion 318 -905 318 -905 0 feedthrough
rlabel pdiffusion 325 -905 325 -905 0 feedthrough
rlabel pdiffusion 332 -905 332 -905 0 feedthrough
rlabel pdiffusion 339 -905 339 -905 0 cellNo=324
rlabel pdiffusion 346 -905 346 -905 0 feedthrough
rlabel pdiffusion 353 -905 353 -905 0 feedthrough
rlabel pdiffusion 360 -905 360 -905 0 cellNo=703
rlabel pdiffusion 367 -905 367 -905 0 feedthrough
rlabel pdiffusion 374 -905 374 -905 0 feedthrough
rlabel pdiffusion 381 -905 381 -905 0 feedthrough
rlabel pdiffusion 388 -905 388 -905 0 feedthrough
rlabel pdiffusion 395 -905 395 -905 0 feedthrough
rlabel pdiffusion 402 -905 402 -905 0 cellNo=123
rlabel pdiffusion 409 -905 409 -905 0 cellNo=563
rlabel pdiffusion 416 -905 416 -905 0 feedthrough
rlabel pdiffusion 423 -905 423 -905 0 feedthrough
rlabel pdiffusion 430 -905 430 -905 0 feedthrough
rlabel pdiffusion 437 -905 437 -905 0 feedthrough
rlabel pdiffusion 444 -905 444 -905 0 feedthrough
rlabel pdiffusion 451 -905 451 -905 0 cellNo=544
rlabel pdiffusion 458 -905 458 -905 0 feedthrough
rlabel pdiffusion 465 -905 465 -905 0 feedthrough
rlabel pdiffusion 472 -905 472 -905 0 feedthrough
rlabel pdiffusion 479 -905 479 -905 0 feedthrough
rlabel pdiffusion 486 -905 486 -905 0 feedthrough
rlabel pdiffusion 493 -905 493 -905 0 feedthrough
rlabel pdiffusion 500 -905 500 -905 0 feedthrough
rlabel pdiffusion 507 -905 507 -905 0 cellNo=143
rlabel pdiffusion 514 -905 514 -905 0 feedthrough
rlabel pdiffusion 521 -905 521 -905 0 feedthrough
rlabel pdiffusion 528 -905 528 -905 0 cellNo=422
rlabel pdiffusion 535 -905 535 -905 0 cellNo=369
rlabel pdiffusion 542 -905 542 -905 0 feedthrough
rlabel pdiffusion 556 -905 556 -905 0 feedthrough
rlabel pdiffusion 563 -905 563 -905 0 feedthrough
rlabel pdiffusion 570 -905 570 -905 0 feedthrough
rlabel pdiffusion 577 -905 577 -905 0 feedthrough
rlabel pdiffusion 584 -905 584 -905 0 feedthrough
rlabel pdiffusion 591 -905 591 -905 0 cellNo=460
rlabel pdiffusion 598 -905 598 -905 0 feedthrough
rlabel pdiffusion 605 -905 605 -905 0 feedthrough
rlabel pdiffusion 619 -905 619 -905 0 feedthrough
rlabel pdiffusion 626 -905 626 -905 0 feedthrough
rlabel pdiffusion 633 -905 633 -905 0 feedthrough
rlabel pdiffusion 640 -905 640 -905 0 feedthrough
rlabel pdiffusion 647 -905 647 -905 0 feedthrough
rlabel pdiffusion 654 -905 654 -905 0 feedthrough
rlabel pdiffusion 661 -905 661 -905 0 feedthrough
rlabel pdiffusion 668 -905 668 -905 0 feedthrough
rlabel pdiffusion 675 -905 675 -905 0 feedthrough
rlabel pdiffusion 682 -905 682 -905 0 feedthrough
rlabel pdiffusion 689 -905 689 -905 0 feedthrough
rlabel pdiffusion 696 -905 696 -905 0 cellNo=380
rlabel pdiffusion 703 -905 703 -905 0 feedthrough
rlabel pdiffusion 710 -905 710 -905 0 feedthrough
rlabel pdiffusion 738 -905 738 -905 0 feedthrough
rlabel pdiffusion 759 -905 759 -905 0 feedthrough
rlabel pdiffusion 3 -988 3 -988 0 feedthrough
rlabel pdiffusion 10 -988 10 -988 0 cellNo=53
rlabel pdiffusion 17 -988 17 -988 0 feedthrough
rlabel pdiffusion 24 -988 24 -988 0 cellNo=583
rlabel pdiffusion 31 -988 31 -988 0 feedthrough
rlabel pdiffusion 38 -988 38 -988 0 feedthrough
rlabel pdiffusion 45 -988 45 -988 0 cellNo=471
rlabel pdiffusion 52 -988 52 -988 0 cellNo=219
rlabel pdiffusion 59 -988 59 -988 0 cellNo=645
rlabel pdiffusion 66 -988 66 -988 0 cellNo=116
rlabel pdiffusion 73 -988 73 -988 0 feedthrough
rlabel pdiffusion 80 -988 80 -988 0 feedthrough
rlabel pdiffusion 87 -988 87 -988 0 cellNo=515
rlabel pdiffusion 94 -988 94 -988 0 feedthrough
rlabel pdiffusion 101 -988 101 -988 0 feedthrough
rlabel pdiffusion 108 -988 108 -988 0 cellNo=311
rlabel pdiffusion 115 -988 115 -988 0 feedthrough
rlabel pdiffusion 122 -988 122 -988 0 feedthrough
rlabel pdiffusion 129 -988 129 -988 0 feedthrough
rlabel pdiffusion 136 -988 136 -988 0 cellNo=278
rlabel pdiffusion 143 -988 143 -988 0 cellNo=493
rlabel pdiffusion 150 -988 150 -988 0 cellNo=75
rlabel pdiffusion 157 -988 157 -988 0 feedthrough
rlabel pdiffusion 164 -988 164 -988 0 feedthrough
rlabel pdiffusion 171 -988 171 -988 0 feedthrough
rlabel pdiffusion 178 -988 178 -988 0 cellNo=249
rlabel pdiffusion 185 -988 185 -988 0 cellNo=93
rlabel pdiffusion 192 -988 192 -988 0 feedthrough
rlabel pdiffusion 199 -988 199 -988 0 feedthrough
rlabel pdiffusion 206 -988 206 -988 0 feedthrough
rlabel pdiffusion 213 -988 213 -988 0 feedthrough
rlabel pdiffusion 220 -988 220 -988 0 feedthrough
rlabel pdiffusion 227 -988 227 -988 0 cellNo=125
rlabel pdiffusion 234 -988 234 -988 0 feedthrough
rlabel pdiffusion 241 -988 241 -988 0 feedthrough
rlabel pdiffusion 248 -988 248 -988 0 cellNo=368
rlabel pdiffusion 255 -988 255 -988 0 feedthrough
rlabel pdiffusion 262 -988 262 -988 0 feedthrough
rlabel pdiffusion 269 -988 269 -988 0 feedthrough
rlabel pdiffusion 276 -988 276 -988 0 feedthrough
rlabel pdiffusion 283 -988 283 -988 0 feedthrough
rlabel pdiffusion 290 -988 290 -988 0 cellNo=586
rlabel pdiffusion 297 -988 297 -988 0 feedthrough
rlabel pdiffusion 304 -988 304 -988 0 feedthrough
rlabel pdiffusion 311 -988 311 -988 0 cellNo=401
rlabel pdiffusion 318 -988 318 -988 0 feedthrough
rlabel pdiffusion 325 -988 325 -988 0 feedthrough
rlabel pdiffusion 332 -988 332 -988 0 feedthrough
rlabel pdiffusion 339 -988 339 -988 0 feedthrough
rlabel pdiffusion 346 -988 346 -988 0 feedthrough
rlabel pdiffusion 353 -988 353 -988 0 feedthrough
rlabel pdiffusion 360 -988 360 -988 0 cellNo=223
rlabel pdiffusion 367 -988 367 -988 0 feedthrough
rlabel pdiffusion 374 -988 374 -988 0 feedthrough
rlabel pdiffusion 381 -988 381 -988 0 cellNo=510
rlabel pdiffusion 388 -988 388 -988 0 feedthrough
rlabel pdiffusion 395 -988 395 -988 0 cellNo=119
rlabel pdiffusion 402 -988 402 -988 0 feedthrough
rlabel pdiffusion 409 -988 409 -988 0 cellNo=606
rlabel pdiffusion 416 -988 416 -988 0 feedthrough
rlabel pdiffusion 423 -988 423 -988 0 feedthrough
rlabel pdiffusion 430 -988 430 -988 0 feedthrough
rlabel pdiffusion 437 -988 437 -988 0 feedthrough
rlabel pdiffusion 444 -988 444 -988 0 cellNo=267
rlabel pdiffusion 451 -988 451 -988 0 feedthrough
rlabel pdiffusion 458 -988 458 -988 0 feedthrough
rlabel pdiffusion 465 -988 465 -988 0 feedthrough
rlabel pdiffusion 472 -988 472 -988 0 feedthrough
rlabel pdiffusion 479 -988 479 -988 0 feedthrough
rlabel pdiffusion 486 -988 486 -988 0 cellNo=318
rlabel pdiffusion 493 -988 493 -988 0 feedthrough
rlabel pdiffusion 500 -988 500 -988 0 cellNo=47
rlabel pdiffusion 507 -988 507 -988 0 feedthrough
rlabel pdiffusion 514 -988 514 -988 0 feedthrough
rlabel pdiffusion 521 -988 521 -988 0 feedthrough
rlabel pdiffusion 528 -988 528 -988 0 feedthrough
rlabel pdiffusion 535 -988 535 -988 0 feedthrough
rlabel pdiffusion 542 -988 542 -988 0 feedthrough
rlabel pdiffusion 549 -988 549 -988 0 feedthrough
rlabel pdiffusion 556 -988 556 -988 0 feedthrough
rlabel pdiffusion 563 -988 563 -988 0 feedthrough
rlabel pdiffusion 570 -988 570 -988 0 feedthrough
rlabel pdiffusion 577 -988 577 -988 0 feedthrough
rlabel pdiffusion 584 -988 584 -988 0 feedthrough
rlabel pdiffusion 591 -988 591 -988 0 feedthrough
rlabel pdiffusion 605 -988 605 -988 0 cellNo=642
rlabel pdiffusion 612 -988 612 -988 0 feedthrough
rlabel pdiffusion 619 -988 619 -988 0 cellNo=230
rlabel pdiffusion 626 -988 626 -988 0 feedthrough
rlabel pdiffusion 633 -988 633 -988 0 feedthrough
rlabel pdiffusion 640 -988 640 -988 0 feedthrough
rlabel pdiffusion 647 -988 647 -988 0 feedthrough
rlabel pdiffusion 654 -988 654 -988 0 feedthrough
rlabel pdiffusion 661 -988 661 -988 0 feedthrough
rlabel pdiffusion 668 -988 668 -988 0 feedthrough
rlabel pdiffusion 675 -988 675 -988 0 feedthrough
rlabel pdiffusion 682 -988 682 -988 0 feedthrough
rlabel pdiffusion 689 -988 689 -988 0 feedthrough
rlabel pdiffusion 696 -988 696 -988 0 feedthrough
rlabel pdiffusion 703 -988 703 -988 0 feedthrough
rlabel pdiffusion 710 -988 710 -988 0 feedthrough
rlabel pdiffusion 717 -988 717 -988 0 feedthrough
rlabel pdiffusion 724 -988 724 -988 0 cellNo=525
rlabel pdiffusion 752 -988 752 -988 0 feedthrough
rlabel pdiffusion 10 -1063 10 -1063 0 cellNo=344
rlabel pdiffusion 17 -1063 17 -1063 0 feedthrough
rlabel pdiffusion 24 -1063 24 -1063 0 cellNo=536
rlabel pdiffusion 31 -1063 31 -1063 0 cellNo=234
rlabel pdiffusion 38 -1063 38 -1063 0 feedthrough
rlabel pdiffusion 45 -1063 45 -1063 0 cellNo=14
rlabel pdiffusion 52 -1063 52 -1063 0 cellNo=625
rlabel pdiffusion 59 -1063 59 -1063 0 feedthrough
rlabel pdiffusion 66 -1063 66 -1063 0 feedthrough
rlabel pdiffusion 73 -1063 73 -1063 0 cellNo=46
rlabel pdiffusion 80 -1063 80 -1063 0 feedthrough
rlabel pdiffusion 87 -1063 87 -1063 0 feedthrough
rlabel pdiffusion 94 -1063 94 -1063 0 feedthrough
rlabel pdiffusion 101 -1063 101 -1063 0 cellNo=601
rlabel pdiffusion 108 -1063 108 -1063 0 feedthrough
rlabel pdiffusion 115 -1063 115 -1063 0 cellNo=341
rlabel pdiffusion 122 -1063 122 -1063 0 feedthrough
rlabel pdiffusion 129 -1063 129 -1063 0 feedthrough
rlabel pdiffusion 136 -1063 136 -1063 0 cellNo=393
rlabel pdiffusion 143 -1063 143 -1063 0 feedthrough
rlabel pdiffusion 150 -1063 150 -1063 0 feedthrough
rlabel pdiffusion 157 -1063 157 -1063 0 feedthrough
rlabel pdiffusion 164 -1063 164 -1063 0 feedthrough
rlabel pdiffusion 171 -1063 171 -1063 0 cellNo=528
rlabel pdiffusion 178 -1063 178 -1063 0 feedthrough
rlabel pdiffusion 185 -1063 185 -1063 0 cellNo=166
rlabel pdiffusion 192 -1063 192 -1063 0 feedthrough
rlabel pdiffusion 199 -1063 199 -1063 0 feedthrough
rlabel pdiffusion 206 -1063 206 -1063 0 feedthrough
rlabel pdiffusion 213 -1063 213 -1063 0 feedthrough
rlabel pdiffusion 220 -1063 220 -1063 0 feedthrough
rlabel pdiffusion 227 -1063 227 -1063 0 feedthrough
rlabel pdiffusion 234 -1063 234 -1063 0 feedthrough
rlabel pdiffusion 241 -1063 241 -1063 0 feedthrough
rlabel pdiffusion 248 -1063 248 -1063 0 feedthrough
rlabel pdiffusion 255 -1063 255 -1063 0 feedthrough
rlabel pdiffusion 262 -1063 262 -1063 0 feedthrough
rlabel pdiffusion 269 -1063 269 -1063 0 cellNo=687
rlabel pdiffusion 276 -1063 276 -1063 0 feedthrough
rlabel pdiffusion 283 -1063 283 -1063 0 cellNo=397
rlabel pdiffusion 290 -1063 290 -1063 0 feedthrough
rlabel pdiffusion 297 -1063 297 -1063 0 feedthrough
rlabel pdiffusion 304 -1063 304 -1063 0 cellNo=129
rlabel pdiffusion 311 -1063 311 -1063 0 cellNo=335
rlabel pdiffusion 318 -1063 318 -1063 0 cellNo=437
rlabel pdiffusion 325 -1063 325 -1063 0 feedthrough
rlabel pdiffusion 332 -1063 332 -1063 0 feedthrough
rlabel pdiffusion 339 -1063 339 -1063 0 feedthrough
rlabel pdiffusion 346 -1063 346 -1063 0 feedthrough
rlabel pdiffusion 353 -1063 353 -1063 0 cellNo=436
rlabel pdiffusion 360 -1063 360 -1063 0 cellNo=43
rlabel pdiffusion 367 -1063 367 -1063 0 cellNo=256
rlabel pdiffusion 374 -1063 374 -1063 0 cellNo=35
rlabel pdiffusion 381 -1063 381 -1063 0 feedthrough
rlabel pdiffusion 388 -1063 388 -1063 0 feedthrough
rlabel pdiffusion 395 -1063 395 -1063 0 cellNo=434
rlabel pdiffusion 402 -1063 402 -1063 0 cellNo=293
rlabel pdiffusion 409 -1063 409 -1063 0 feedthrough
rlabel pdiffusion 416 -1063 416 -1063 0 cellNo=464
rlabel pdiffusion 423 -1063 423 -1063 0 cellNo=602
rlabel pdiffusion 430 -1063 430 -1063 0 feedthrough
rlabel pdiffusion 437 -1063 437 -1063 0 feedthrough
rlabel pdiffusion 444 -1063 444 -1063 0 feedthrough
rlabel pdiffusion 451 -1063 451 -1063 0 cellNo=118
rlabel pdiffusion 458 -1063 458 -1063 0 feedthrough
rlabel pdiffusion 465 -1063 465 -1063 0 feedthrough
rlabel pdiffusion 472 -1063 472 -1063 0 feedthrough
rlabel pdiffusion 479 -1063 479 -1063 0 feedthrough
rlabel pdiffusion 486 -1063 486 -1063 0 feedthrough
rlabel pdiffusion 493 -1063 493 -1063 0 feedthrough
rlabel pdiffusion 500 -1063 500 -1063 0 feedthrough
rlabel pdiffusion 507 -1063 507 -1063 0 feedthrough
rlabel pdiffusion 514 -1063 514 -1063 0 feedthrough
rlabel pdiffusion 521 -1063 521 -1063 0 feedthrough
rlabel pdiffusion 528 -1063 528 -1063 0 feedthrough
rlabel pdiffusion 535 -1063 535 -1063 0 feedthrough
rlabel pdiffusion 542 -1063 542 -1063 0 feedthrough
rlabel pdiffusion 549 -1063 549 -1063 0 feedthrough
rlabel pdiffusion 556 -1063 556 -1063 0 feedthrough
rlabel pdiffusion 563 -1063 563 -1063 0 feedthrough
rlabel pdiffusion 570 -1063 570 -1063 0 feedthrough
rlabel pdiffusion 577 -1063 577 -1063 0 feedthrough
rlabel pdiffusion 584 -1063 584 -1063 0 feedthrough
rlabel pdiffusion 591 -1063 591 -1063 0 feedthrough
rlabel pdiffusion 598 -1063 598 -1063 0 feedthrough
rlabel pdiffusion 605 -1063 605 -1063 0 cellNo=342
rlabel pdiffusion 612 -1063 612 -1063 0 feedthrough
rlabel pdiffusion 619 -1063 619 -1063 0 feedthrough
rlabel pdiffusion 626 -1063 626 -1063 0 feedthrough
rlabel pdiffusion 633 -1063 633 -1063 0 feedthrough
rlabel pdiffusion 640 -1063 640 -1063 0 feedthrough
rlabel pdiffusion 647 -1063 647 -1063 0 feedthrough
rlabel pdiffusion 654 -1063 654 -1063 0 feedthrough
rlabel pdiffusion 661 -1063 661 -1063 0 feedthrough
rlabel pdiffusion 668 -1063 668 -1063 0 feedthrough
rlabel pdiffusion 675 -1063 675 -1063 0 feedthrough
rlabel pdiffusion 682 -1063 682 -1063 0 feedthrough
rlabel pdiffusion 689 -1063 689 -1063 0 feedthrough
rlabel pdiffusion 696 -1063 696 -1063 0 feedthrough
rlabel pdiffusion 703 -1063 703 -1063 0 feedthrough
rlabel pdiffusion 710 -1063 710 -1063 0 feedthrough
rlabel pdiffusion 717 -1063 717 -1063 0 feedthrough
rlabel pdiffusion 724 -1063 724 -1063 0 feedthrough
rlabel pdiffusion 731 -1063 731 -1063 0 feedthrough
rlabel pdiffusion 752 -1063 752 -1063 0 cellNo=715
rlabel pdiffusion 759 -1063 759 -1063 0 feedthrough
rlabel pdiffusion 10 -1130 10 -1130 0 feedthrough
rlabel pdiffusion 17 -1130 17 -1130 0 feedthrough
rlabel pdiffusion 24 -1130 24 -1130 0 cellNo=711
rlabel pdiffusion 38 -1130 38 -1130 0 feedthrough
rlabel pdiffusion 45 -1130 45 -1130 0 feedthrough
rlabel pdiffusion 52 -1130 52 -1130 0 feedthrough
rlabel pdiffusion 59 -1130 59 -1130 0 feedthrough
rlabel pdiffusion 66 -1130 66 -1130 0 feedthrough
rlabel pdiffusion 73 -1130 73 -1130 0 feedthrough
rlabel pdiffusion 80 -1130 80 -1130 0 feedthrough
rlabel pdiffusion 87 -1130 87 -1130 0 cellNo=712
rlabel pdiffusion 94 -1130 94 -1130 0 feedthrough
rlabel pdiffusion 101 -1130 101 -1130 0 feedthrough
rlabel pdiffusion 108 -1130 108 -1130 0 feedthrough
rlabel pdiffusion 115 -1130 115 -1130 0 cellNo=200
rlabel pdiffusion 122 -1130 122 -1130 0 feedthrough
rlabel pdiffusion 129 -1130 129 -1130 0 feedthrough
rlabel pdiffusion 136 -1130 136 -1130 0 cellNo=160
rlabel pdiffusion 143 -1130 143 -1130 0 feedthrough
rlabel pdiffusion 150 -1130 150 -1130 0 cellNo=406
rlabel pdiffusion 157 -1130 157 -1130 0 feedthrough
rlabel pdiffusion 164 -1130 164 -1130 0 cellNo=556
rlabel pdiffusion 171 -1130 171 -1130 0 feedthrough
rlabel pdiffusion 178 -1130 178 -1130 0 cellNo=101
rlabel pdiffusion 185 -1130 185 -1130 0 cellNo=531
rlabel pdiffusion 192 -1130 192 -1130 0 cellNo=463
rlabel pdiffusion 199 -1130 199 -1130 0 feedthrough
rlabel pdiffusion 206 -1130 206 -1130 0 cellNo=485
rlabel pdiffusion 213 -1130 213 -1130 0 feedthrough
rlabel pdiffusion 220 -1130 220 -1130 0 feedthrough
rlabel pdiffusion 227 -1130 227 -1130 0 feedthrough
rlabel pdiffusion 234 -1130 234 -1130 0 cellNo=184
rlabel pdiffusion 241 -1130 241 -1130 0 feedthrough
rlabel pdiffusion 248 -1130 248 -1130 0 cellNo=610
rlabel pdiffusion 255 -1130 255 -1130 0 feedthrough
rlabel pdiffusion 262 -1130 262 -1130 0 feedthrough
rlabel pdiffusion 269 -1130 269 -1130 0 feedthrough
rlabel pdiffusion 276 -1130 276 -1130 0 feedthrough
rlabel pdiffusion 283 -1130 283 -1130 0 cellNo=557
rlabel pdiffusion 290 -1130 290 -1130 0 cellNo=621
rlabel pdiffusion 297 -1130 297 -1130 0 feedthrough
rlabel pdiffusion 304 -1130 304 -1130 0 feedthrough
rlabel pdiffusion 311 -1130 311 -1130 0 feedthrough
rlabel pdiffusion 318 -1130 318 -1130 0 cellNo=527
rlabel pdiffusion 325 -1130 325 -1130 0 cellNo=49
rlabel pdiffusion 332 -1130 332 -1130 0 feedthrough
rlabel pdiffusion 339 -1130 339 -1130 0 feedthrough
rlabel pdiffusion 346 -1130 346 -1130 0 feedthrough
rlabel pdiffusion 353 -1130 353 -1130 0 cellNo=673
rlabel pdiffusion 360 -1130 360 -1130 0 feedthrough
rlabel pdiffusion 367 -1130 367 -1130 0 cellNo=163
rlabel pdiffusion 374 -1130 374 -1130 0 feedthrough
rlabel pdiffusion 381 -1130 381 -1130 0 cellNo=662
rlabel pdiffusion 388 -1130 388 -1130 0 feedthrough
rlabel pdiffusion 395 -1130 395 -1130 0 feedthrough
rlabel pdiffusion 402 -1130 402 -1130 0 feedthrough
rlabel pdiffusion 409 -1130 409 -1130 0 feedthrough
rlabel pdiffusion 416 -1130 416 -1130 0 feedthrough
rlabel pdiffusion 423 -1130 423 -1130 0 cellNo=545
rlabel pdiffusion 430 -1130 430 -1130 0 cellNo=334
rlabel pdiffusion 437 -1130 437 -1130 0 cellNo=546
rlabel pdiffusion 444 -1130 444 -1130 0 feedthrough
rlabel pdiffusion 451 -1130 451 -1130 0 feedthrough
rlabel pdiffusion 458 -1130 458 -1130 0 feedthrough
rlabel pdiffusion 465 -1130 465 -1130 0 feedthrough
rlabel pdiffusion 472 -1130 472 -1130 0 cellNo=633
rlabel pdiffusion 479 -1130 479 -1130 0 feedthrough
rlabel pdiffusion 486 -1130 486 -1130 0 feedthrough
rlabel pdiffusion 493 -1130 493 -1130 0 feedthrough
rlabel pdiffusion 500 -1130 500 -1130 0 feedthrough
rlabel pdiffusion 507 -1130 507 -1130 0 cellNo=373
rlabel pdiffusion 514 -1130 514 -1130 0 feedthrough
rlabel pdiffusion 521 -1130 521 -1130 0 feedthrough
rlabel pdiffusion 528 -1130 528 -1130 0 feedthrough
rlabel pdiffusion 535 -1130 535 -1130 0 feedthrough
rlabel pdiffusion 542 -1130 542 -1130 0 feedthrough
rlabel pdiffusion 549 -1130 549 -1130 0 feedthrough
rlabel pdiffusion 556 -1130 556 -1130 0 feedthrough
rlabel pdiffusion 563 -1130 563 -1130 0 feedthrough
rlabel pdiffusion 570 -1130 570 -1130 0 feedthrough
rlabel pdiffusion 577 -1130 577 -1130 0 feedthrough
rlabel pdiffusion 584 -1130 584 -1130 0 feedthrough
rlabel pdiffusion 591 -1130 591 -1130 0 feedthrough
rlabel pdiffusion 598 -1130 598 -1130 0 feedthrough
rlabel pdiffusion 605 -1130 605 -1130 0 feedthrough
rlabel pdiffusion 626 -1130 626 -1130 0 feedthrough
rlabel pdiffusion 633 -1130 633 -1130 0 feedthrough
rlabel pdiffusion 640 -1130 640 -1130 0 feedthrough
rlabel pdiffusion 647 -1130 647 -1130 0 feedthrough
rlabel pdiffusion 654 -1130 654 -1130 0 feedthrough
rlabel pdiffusion 661 -1130 661 -1130 0 feedthrough
rlabel pdiffusion 668 -1130 668 -1130 0 feedthrough
rlabel pdiffusion 675 -1130 675 -1130 0 feedthrough
rlabel pdiffusion 682 -1130 682 -1130 0 feedthrough
rlabel pdiffusion 696 -1130 696 -1130 0 feedthrough
rlabel pdiffusion 703 -1130 703 -1130 0 feedthrough
rlabel pdiffusion 710 -1130 710 -1130 0 feedthrough
rlabel pdiffusion 717 -1130 717 -1130 0 feedthrough
rlabel pdiffusion 724 -1130 724 -1130 0 feedthrough
rlabel pdiffusion 731 -1130 731 -1130 0 feedthrough
rlabel pdiffusion 738 -1130 738 -1130 0 cellNo=448
rlabel pdiffusion 745 -1130 745 -1130 0 cellNo=600
rlabel pdiffusion 752 -1130 752 -1130 0 cellNo=475
rlabel pdiffusion 759 -1130 759 -1130 0 feedthrough
rlabel pdiffusion 780 -1130 780 -1130 0 feedthrough
rlabel pdiffusion 787 -1130 787 -1130 0 feedthrough
rlabel pdiffusion 794 -1130 794 -1130 0 feedthrough
rlabel pdiffusion 815 -1130 815 -1130 0 feedthrough
rlabel pdiffusion 10 -1211 10 -1211 0 feedthrough
rlabel pdiffusion 17 -1211 17 -1211 0 feedthrough
rlabel pdiffusion 24 -1211 24 -1211 0 feedthrough
rlabel pdiffusion 31 -1211 31 -1211 0 cellNo=708
rlabel pdiffusion 38 -1211 38 -1211 0 cellNo=499
rlabel pdiffusion 45 -1211 45 -1211 0 feedthrough
rlabel pdiffusion 52 -1211 52 -1211 0 cellNo=265
rlabel pdiffusion 59 -1211 59 -1211 0 feedthrough
rlabel pdiffusion 66 -1211 66 -1211 0 cellNo=48
rlabel pdiffusion 73 -1211 73 -1211 0 feedthrough
rlabel pdiffusion 80 -1211 80 -1211 0 feedthrough
rlabel pdiffusion 87 -1211 87 -1211 0 cellNo=257
rlabel pdiffusion 94 -1211 94 -1211 0 feedthrough
rlabel pdiffusion 101 -1211 101 -1211 0 feedthrough
rlabel pdiffusion 108 -1211 108 -1211 0 feedthrough
rlabel pdiffusion 115 -1211 115 -1211 0 cellNo=156
rlabel pdiffusion 122 -1211 122 -1211 0 feedthrough
rlabel pdiffusion 129 -1211 129 -1211 0 feedthrough
rlabel pdiffusion 136 -1211 136 -1211 0 feedthrough
rlabel pdiffusion 143 -1211 143 -1211 0 cellNo=319
rlabel pdiffusion 150 -1211 150 -1211 0 feedthrough
rlabel pdiffusion 157 -1211 157 -1211 0 feedthrough
rlabel pdiffusion 164 -1211 164 -1211 0 cellNo=541
rlabel pdiffusion 171 -1211 171 -1211 0 feedthrough
rlabel pdiffusion 178 -1211 178 -1211 0 feedthrough
rlabel pdiffusion 185 -1211 185 -1211 0 cellNo=699
rlabel pdiffusion 192 -1211 192 -1211 0 feedthrough
rlabel pdiffusion 199 -1211 199 -1211 0 feedthrough
rlabel pdiffusion 206 -1211 206 -1211 0 feedthrough
rlabel pdiffusion 213 -1211 213 -1211 0 feedthrough
rlabel pdiffusion 220 -1211 220 -1211 0 feedthrough
rlabel pdiffusion 227 -1211 227 -1211 0 feedthrough
rlabel pdiffusion 234 -1211 234 -1211 0 cellNo=484
rlabel pdiffusion 241 -1211 241 -1211 0 feedthrough
rlabel pdiffusion 248 -1211 248 -1211 0 feedthrough
rlabel pdiffusion 255 -1211 255 -1211 0 cellNo=173
rlabel pdiffusion 262 -1211 262 -1211 0 feedthrough
rlabel pdiffusion 269 -1211 269 -1211 0 feedthrough
rlabel pdiffusion 276 -1211 276 -1211 0 cellNo=682
rlabel pdiffusion 283 -1211 283 -1211 0 feedthrough
rlabel pdiffusion 290 -1211 290 -1211 0 feedthrough
rlabel pdiffusion 297 -1211 297 -1211 0 feedthrough
rlabel pdiffusion 304 -1211 304 -1211 0 feedthrough
rlabel pdiffusion 311 -1211 311 -1211 0 feedthrough
rlabel pdiffusion 318 -1211 318 -1211 0 cellNo=171
rlabel pdiffusion 325 -1211 325 -1211 0 cellNo=398
rlabel pdiffusion 332 -1211 332 -1211 0 feedthrough
rlabel pdiffusion 339 -1211 339 -1211 0 cellNo=286
rlabel pdiffusion 346 -1211 346 -1211 0 cellNo=151
rlabel pdiffusion 353 -1211 353 -1211 0 feedthrough
rlabel pdiffusion 360 -1211 360 -1211 0 feedthrough
rlabel pdiffusion 367 -1211 367 -1211 0 cellNo=272
rlabel pdiffusion 374 -1211 374 -1211 0 feedthrough
rlabel pdiffusion 381 -1211 381 -1211 0 feedthrough
rlabel pdiffusion 388 -1211 388 -1211 0 cellNo=488
rlabel pdiffusion 395 -1211 395 -1211 0 cellNo=454
rlabel pdiffusion 402 -1211 402 -1211 0 cellNo=203
rlabel pdiffusion 409 -1211 409 -1211 0 cellNo=161
rlabel pdiffusion 416 -1211 416 -1211 0 feedthrough
rlabel pdiffusion 423 -1211 423 -1211 0 feedthrough
rlabel pdiffusion 430 -1211 430 -1211 0 feedthrough
rlabel pdiffusion 437 -1211 437 -1211 0 feedthrough
rlabel pdiffusion 444 -1211 444 -1211 0 feedthrough
rlabel pdiffusion 451 -1211 451 -1211 0 feedthrough
rlabel pdiffusion 458 -1211 458 -1211 0 feedthrough
rlabel pdiffusion 465 -1211 465 -1211 0 cellNo=427
rlabel pdiffusion 472 -1211 472 -1211 0 cellNo=227
rlabel pdiffusion 479 -1211 479 -1211 0 cellNo=710
rlabel pdiffusion 486 -1211 486 -1211 0 feedthrough
rlabel pdiffusion 493 -1211 493 -1211 0 feedthrough
rlabel pdiffusion 500 -1211 500 -1211 0 feedthrough
rlabel pdiffusion 507 -1211 507 -1211 0 feedthrough
rlabel pdiffusion 514 -1211 514 -1211 0 feedthrough
rlabel pdiffusion 521 -1211 521 -1211 0 feedthrough
rlabel pdiffusion 528 -1211 528 -1211 0 feedthrough
rlabel pdiffusion 535 -1211 535 -1211 0 feedthrough
rlabel pdiffusion 542 -1211 542 -1211 0 cellNo=297
rlabel pdiffusion 549 -1211 549 -1211 0 feedthrough
rlabel pdiffusion 556 -1211 556 -1211 0 feedthrough
rlabel pdiffusion 563 -1211 563 -1211 0 feedthrough
rlabel pdiffusion 570 -1211 570 -1211 0 feedthrough
rlabel pdiffusion 577 -1211 577 -1211 0 feedthrough
rlabel pdiffusion 584 -1211 584 -1211 0 feedthrough
rlabel pdiffusion 591 -1211 591 -1211 0 cellNo=26
rlabel pdiffusion 598 -1211 598 -1211 0 feedthrough
rlabel pdiffusion 605 -1211 605 -1211 0 feedthrough
rlabel pdiffusion 612 -1211 612 -1211 0 feedthrough
rlabel pdiffusion 619 -1211 619 -1211 0 feedthrough
rlabel pdiffusion 626 -1211 626 -1211 0 feedthrough
rlabel pdiffusion 633 -1211 633 -1211 0 feedthrough
rlabel pdiffusion 640 -1211 640 -1211 0 feedthrough
rlabel pdiffusion 647 -1211 647 -1211 0 feedthrough
rlabel pdiffusion 654 -1211 654 -1211 0 feedthrough
rlabel pdiffusion 661 -1211 661 -1211 0 cellNo=477
rlabel pdiffusion 668 -1211 668 -1211 0 feedthrough
rlabel pdiffusion 675 -1211 675 -1211 0 feedthrough
rlabel pdiffusion 682 -1211 682 -1211 0 feedthrough
rlabel pdiffusion 689 -1211 689 -1211 0 feedthrough
rlabel pdiffusion 696 -1211 696 -1211 0 feedthrough
rlabel pdiffusion 703 -1211 703 -1211 0 feedthrough
rlabel pdiffusion 710 -1211 710 -1211 0 feedthrough
rlabel pdiffusion 717 -1211 717 -1211 0 feedthrough
rlabel pdiffusion 724 -1211 724 -1211 0 feedthrough
rlabel pdiffusion 731 -1211 731 -1211 0 feedthrough
rlabel pdiffusion 745 -1211 745 -1211 0 feedthrough
rlabel pdiffusion 752 -1211 752 -1211 0 feedthrough
rlabel pdiffusion 759 -1211 759 -1211 0 feedthrough
rlabel pdiffusion 766 -1211 766 -1211 0 feedthrough
rlabel pdiffusion 773 -1211 773 -1211 0 feedthrough
rlabel pdiffusion 780 -1211 780 -1211 0 feedthrough
rlabel pdiffusion 787 -1211 787 -1211 0 feedthrough
rlabel pdiffusion 794 -1211 794 -1211 0 feedthrough
rlabel pdiffusion 801 -1211 801 -1211 0 feedthrough
rlabel pdiffusion 3 -1304 3 -1304 0 feedthrough
rlabel pdiffusion 10 -1304 10 -1304 0 feedthrough
rlabel pdiffusion 17 -1304 17 -1304 0 feedthrough
rlabel pdiffusion 24 -1304 24 -1304 0 feedthrough
rlabel pdiffusion 31 -1304 31 -1304 0 feedthrough
rlabel pdiffusion 38 -1304 38 -1304 0 feedthrough
rlabel pdiffusion 45 -1304 45 -1304 0 feedthrough
rlabel pdiffusion 52 -1304 52 -1304 0 feedthrough
rlabel pdiffusion 59 -1304 59 -1304 0 feedthrough
rlabel pdiffusion 66 -1304 66 -1304 0 cellNo=332
rlabel pdiffusion 73 -1304 73 -1304 0 cellNo=415
rlabel pdiffusion 80 -1304 80 -1304 0 feedthrough
rlabel pdiffusion 87 -1304 87 -1304 0 feedthrough
rlabel pdiffusion 94 -1304 94 -1304 0 feedthrough
rlabel pdiffusion 101 -1304 101 -1304 0 feedthrough
rlabel pdiffusion 108 -1304 108 -1304 0 feedthrough
rlabel pdiffusion 115 -1304 115 -1304 0 cellNo=423
rlabel pdiffusion 122 -1304 122 -1304 0 feedthrough
rlabel pdiffusion 129 -1304 129 -1304 0 feedthrough
rlabel pdiffusion 136 -1304 136 -1304 0 feedthrough
rlabel pdiffusion 143 -1304 143 -1304 0 cellNo=8
rlabel pdiffusion 150 -1304 150 -1304 0 feedthrough
rlabel pdiffusion 157 -1304 157 -1304 0 feedthrough
rlabel pdiffusion 164 -1304 164 -1304 0 cellNo=619
rlabel pdiffusion 171 -1304 171 -1304 0 feedthrough
rlabel pdiffusion 178 -1304 178 -1304 0 feedthrough
rlabel pdiffusion 185 -1304 185 -1304 0 cellNo=446
rlabel pdiffusion 192 -1304 192 -1304 0 feedthrough
rlabel pdiffusion 199 -1304 199 -1304 0 cellNo=194
rlabel pdiffusion 206 -1304 206 -1304 0 feedthrough
rlabel pdiffusion 213 -1304 213 -1304 0 feedthrough
rlabel pdiffusion 220 -1304 220 -1304 0 feedthrough
rlabel pdiffusion 227 -1304 227 -1304 0 cellNo=127
rlabel pdiffusion 234 -1304 234 -1304 0 feedthrough
rlabel pdiffusion 241 -1304 241 -1304 0 feedthrough
rlabel pdiffusion 248 -1304 248 -1304 0 feedthrough
rlabel pdiffusion 255 -1304 255 -1304 0 feedthrough
rlabel pdiffusion 262 -1304 262 -1304 0 feedthrough
rlabel pdiffusion 269 -1304 269 -1304 0 feedthrough
rlabel pdiffusion 276 -1304 276 -1304 0 feedthrough
rlabel pdiffusion 283 -1304 283 -1304 0 feedthrough
rlabel pdiffusion 290 -1304 290 -1304 0 feedthrough
rlabel pdiffusion 297 -1304 297 -1304 0 feedthrough
rlabel pdiffusion 304 -1304 304 -1304 0 cellNo=24
rlabel pdiffusion 311 -1304 311 -1304 0 cellNo=271
rlabel pdiffusion 318 -1304 318 -1304 0 feedthrough
rlabel pdiffusion 325 -1304 325 -1304 0 feedthrough
rlabel pdiffusion 332 -1304 332 -1304 0 cellNo=54
rlabel pdiffusion 339 -1304 339 -1304 0 cellNo=709
rlabel pdiffusion 346 -1304 346 -1304 0 feedthrough
rlabel pdiffusion 353 -1304 353 -1304 0 cellNo=32
rlabel pdiffusion 360 -1304 360 -1304 0 cellNo=656
rlabel pdiffusion 367 -1304 367 -1304 0 cellNo=615
rlabel pdiffusion 374 -1304 374 -1304 0 feedthrough
rlabel pdiffusion 381 -1304 381 -1304 0 feedthrough
rlabel pdiffusion 388 -1304 388 -1304 0 feedthrough
rlabel pdiffusion 395 -1304 395 -1304 0 feedthrough
rlabel pdiffusion 402 -1304 402 -1304 0 cellNo=340
rlabel pdiffusion 409 -1304 409 -1304 0 cellNo=553
rlabel pdiffusion 416 -1304 416 -1304 0 feedthrough
rlabel pdiffusion 423 -1304 423 -1304 0 cellNo=59
rlabel pdiffusion 430 -1304 430 -1304 0 feedthrough
rlabel pdiffusion 437 -1304 437 -1304 0 feedthrough
rlabel pdiffusion 444 -1304 444 -1304 0 feedthrough
rlabel pdiffusion 451 -1304 451 -1304 0 cellNo=262
rlabel pdiffusion 458 -1304 458 -1304 0 cellNo=254
rlabel pdiffusion 465 -1304 465 -1304 0 feedthrough
rlabel pdiffusion 472 -1304 472 -1304 0 feedthrough
rlabel pdiffusion 479 -1304 479 -1304 0 feedthrough
rlabel pdiffusion 486 -1304 486 -1304 0 feedthrough
rlabel pdiffusion 493 -1304 493 -1304 0 feedthrough
rlabel pdiffusion 500 -1304 500 -1304 0 feedthrough
rlabel pdiffusion 507 -1304 507 -1304 0 feedthrough
rlabel pdiffusion 514 -1304 514 -1304 0 feedthrough
rlabel pdiffusion 521 -1304 521 -1304 0 feedthrough
rlabel pdiffusion 528 -1304 528 -1304 0 feedthrough
rlabel pdiffusion 535 -1304 535 -1304 0 cellNo=585
rlabel pdiffusion 542 -1304 542 -1304 0 feedthrough
rlabel pdiffusion 549 -1304 549 -1304 0 feedthrough
rlabel pdiffusion 556 -1304 556 -1304 0 feedthrough
rlabel pdiffusion 563 -1304 563 -1304 0 feedthrough
rlabel pdiffusion 570 -1304 570 -1304 0 cellNo=326
rlabel pdiffusion 577 -1304 577 -1304 0 feedthrough
rlabel pdiffusion 584 -1304 584 -1304 0 feedthrough
rlabel pdiffusion 591 -1304 591 -1304 0 feedthrough
rlabel pdiffusion 598 -1304 598 -1304 0 feedthrough
rlabel pdiffusion 605 -1304 605 -1304 0 feedthrough
rlabel pdiffusion 612 -1304 612 -1304 0 feedthrough
rlabel pdiffusion 619 -1304 619 -1304 0 feedthrough
rlabel pdiffusion 626 -1304 626 -1304 0 feedthrough
rlabel pdiffusion 633 -1304 633 -1304 0 feedthrough
rlabel pdiffusion 640 -1304 640 -1304 0 feedthrough
rlabel pdiffusion 647 -1304 647 -1304 0 cellNo=356
rlabel pdiffusion 654 -1304 654 -1304 0 feedthrough
rlabel pdiffusion 661 -1304 661 -1304 0 feedthrough
rlabel pdiffusion 668 -1304 668 -1304 0 feedthrough
rlabel pdiffusion 675 -1304 675 -1304 0 feedthrough
rlabel pdiffusion 682 -1304 682 -1304 0 feedthrough
rlabel pdiffusion 689 -1304 689 -1304 0 feedthrough
rlabel pdiffusion 696 -1304 696 -1304 0 feedthrough
rlabel pdiffusion 703 -1304 703 -1304 0 feedthrough
rlabel pdiffusion 710 -1304 710 -1304 0 feedthrough
rlabel pdiffusion 717 -1304 717 -1304 0 feedthrough
rlabel pdiffusion 724 -1304 724 -1304 0 feedthrough
rlabel pdiffusion 731 -1304 731 -1304 0 feedthrough
rlabel pdiffusion 738 -1304 738 -1304 0 feedthrough
rlabel pdiffusion 745 -1304 745 -1304 0 feedthrough
rlabel pdiffusion 752 -1304 752 -1304 0 feedthrough
rlabel pdiffusion 759 -1304 759 -1304 0 feedthrough
rlabel pdiffusion 766 -1304 766 -1304 0 cellNo=568
rlabel pdiffusion 773 -1304 773 -1304 0 cellNo=584
rlabel pdiffusion 780 -1304 780 -1304 0 cellNo=236
rlabel pdiffusion 787 -1304 787 -1304 0 cellNo=391
rlabel pdiffusion 10 -1381 10 -1381 0 cellNo=580
rlabel pdiffusion 24 -1381 24 -1381 0 feedthrough
rlabel pdiffusion 31 -1381 31 -1381 0 feedthrough
rlabel pdiffusion 38 -1381 38 -1381 0 cellNo=700
rlabel pdiffusion 45 -1381 45 -1381 0 feedthrough
rlabel pdiffusion 52 -1381 52 -1381 0 feedthrough
rlabel pdiffusion 59 -1381 59 -1381 0 feedthrough
rlabel pdiffusion 66 -1381 66 -1381 0 feedthrough
rlabel pdiffusion 73 -1381 73 -1381 0 cellNo=500
rlabel pdiffusion 80 -1381 80 -1381 0 cellNo=301
rlabel pdiffusion 87 -1381 87 -1381 0 cellNo=404
rlabel pdiffusion 94 -1381 94 -1381 0 cellNo=465
rlabel pdiffusion 101 -1381 101 -1381 0 feedthrough
rlabel pdiffusion 108 -1381 108 -1381 0 feedthrough
rlabel pdiffusion 115 -1381 115 -1381 0 cellNo=182
rlabel pdiffusion 122 -1381 122 -1381 0 feedthrough
rlabel pdiffusion 129 -1381 129 -1381 0 feedthrough
rlabel pdiffusion 136 -1381 136 -1381 0 feedthrough
rlabel pdiffusion 143 -1381 143 -1381 0 cellNo=613
rlabel pdiffusion 150 -1381 150 -1381 0 feedthrough
rlabel pdiffusion 157 -1381 157 -1381 0 feedthrough
rlabel pdiffusion 164 -1381 164 -1381 0 cellNo=653
rlabel pdiffusion 171 -1381 171 -1381 0 feedthrough
rlabel pdiffusion 178 -1381 178 -1381 0 cellNo=232
rlabel pdiffusion 185 -1381 185 -1381 0 cellNo=316
rlabel pdiffusion 192 -1381 192 -1381 0 feedthrough
rlabel pdiffusion 199 -1381 199 -1381 0 feedthrough
rlabel pdiffusion 206 -1381 206 -1381 0 feedthrough
rlabel pdiffusion 213 -1381 213 -1381 0 cellNo=597
rlabel pdiffusion 220 -1381 220 -1381 0 feedthrough
rlabel pdiffusion 227 -1381 227 -1381 0 feedthrough
rlabel pdiffusion 234 -1381 234 -1381 0 feedthrough
rlabel pdiffusion 241 -1381 241 -1381 0 feedthrough
rlabel pdiffusion 248 -1381 248 -1381 0 feedthrough
rlabel pdiffusion 255 -1381 255 -1381 0 feedthrough
rlabel pdiffusion 262 -1381 262 -1381 0 feedthrough
rlabel pdiffusion 269 -1381 269 -1381 0 feedthrough
rlabel pdiffusion 276 -1381 276 -1381 0 cellNo=41
rlabel pdiffusion 283 -1381 283 -1381 0 feedthrough
rlabel pdiffusion 290 -1381 290 -1381 0 feedthrough
rlabel pdiffusion 297 -1381 297 -1381 0 cellNo=39
rlabel pdiffusion 304 -1381 304 -1381 0 feedthrough
rlabel pdiffusion 311 -1381 311 -1381 0 feedthrough
rlabel pdiffusion 318 -1381 318 -1381 0 cellNo=444
rlabel pdiffusion 325 -1381 325 -1381 0 feedthrough
rlabel pdiffusion 332 -1381 332 -1381 0 cellNo=162
rlabel pdiffusion 339 -1381 339 -1381 0 feedthrough
rlabel pdiffusion 346 -1381 346 -1381 0 cellNo=289
rlabel pdiffusion 353 -1381 353 -1381 0 feedthrough
rlabel pdiffusion 360 -1381 360 -1381 0 feedthrough
rlabel pdiffusion 367 -1381 367 -1381 0 feedthrough
rlabel pdiffusion 374 -1381 374 -1381 0 feedthrough
rlabel pdiffusion 381 -1381 381 -1381 0 feedthrough
rlabel pdiffusion 388 -1381 388 -1381 0 feedthrough
rlabel pdiffusion 395 -1381 395 -1381 0 feedthrough
rlabel pdiffusion 402 -1381 402 -1381 0 cellNo=651
rlabel pdiffusion 409 -1381 409 -1381 0 cellNo=209
rlabel pdiffusion 416 -1381 416 -1381 0 feedthrough
rlabel pdiffusion 423 -1381 423 -1381 0 feedthrough
rlabel pdiffusion 430 -1381 430 -1381 0 feedthrough
rlabel pdiffusion 437 -1381 437 -1381 0 feedthrough
rlabel pdiffusion 444 -1381 444 -1381 0 cellNo=167
rlabel pdiffusion 451 -1381 451 -1381 0 feedthrough
rlabel pdiffusion 458 -1381 458 -1381 0 feedthrough
rlabel pdiffusion 465 -1381 465 -1381 0 feedthrough
rlabel pdiffusion 472 -1381 472 -1381 0 feedthrough
rlabel pdiffusion 479 -1381 479 -1381 0 cellNo=78
rlabel pdiffusion 486 -1381 486 -1381 0 feedthrough
rlabel pdiffusion 493 -1381 493 -1381 0 feedthrough
rlabel pdiffusion 500 -1381 500 -1381 0 feedthrough
rlabel pdiffusion 507 -1381 507 -1381 0 feedthrough
rlabel pdiffusion 514 -1381 514 -1381 0 cellNo=220
rlabel pdiffusion 521 -1381 521 -1381 0 feedthrough
rlabel pdiffusion 528 -1381 528 -1381 0 feedthrough
rlabel pdiffusion 535 -1381 535 -1381 0 feedthrough
rlabel pdiffusion 542 -1381 542 -1381 0 feedthrough
rlabel pdiffusion 549 -1381 549 -1381 0 feedthrough
rlabel pdiffusion 556 -1381 556 -1381 0 feedthrough
rlabel pdiffusion 563 -1381 563 -1381 0 cellNo=482
rlabel pdiffusion 570 -1381 570 -1381 0 cellNo=193
rlabel pdiffusion 577 -1381 577 -1381 0 feedthrough
rlabel pdiffusion 584 -1381 584 -1381 0 feedthrough
rlabel pdiffusion 591 -1381 591 -1381 0 feedthrough
rlabel pdiffusion 598 -1381 598 -1381 0 feedthrough
rlabel pdiffusion 605 -1381 605 -1381 0 feedthrough
rlabel pdiffusion 612 -1381 612 -1381 0 feedthrough
rlabel pdiffusion 619 -1381 619 -1381 0 feedthrough
rlabel pdiffusion 633 -1381 633 -1381 0 feedthrough
rlabel pdiffusion 640 -1381 640 -1381 0 feedthrough
rlabel pdiffusion 647 -1381 647 -1381 0 feedthrough
rlabel pdiffusion 654 -1381 654 -1381 0 feedthrough
rlabel pdiffusion 661 -1381 661 -1381 0 feedthrough
rlabel pdiffusion 668 -1381 668 -1381 0 feedthrough
rlabel pdiffusion 675 -1381 675 -1381 0 feedthrough
rlabel pdiffusion 682 -1381 682 -1381 0 feedthrough
rlabel pdiffusion 689 -1381 689 -1381 0 cellNo=468
rlabel pdiffusion 696 -1381 696 -1381 0 feedthrough
rlabel pdiffusion 703 -1381 703 -1381 0 cellNo=387
rlabel pdiffusion 710 -1381 710 -1381 0 feedthrough
rlabel pdiffusion 717 -1381 717 -1381 0 cellNo=353
rlabel pdiffusion 759 -1381 759 -1381 0 feedthrough
rlabel pdiffusion 780 -1381 780 -1381 0 feedthrough
rlabel pdiffusion 801 -1381 801 -1381 0 feedthrough
rlabel pdiffusion 10 -1450 10 -1450 0 feedthrough
rlabel pdiffusion 17 -1450 17 -1450 0 feedthrough
rlabel pdiffusion 24 -1450 24 -1450 0 feedthrough
rlabel pdiffusion 31 -1450 31 -1450 0 feedthrough
rlabel pdiffusion 38 -1450 38 -1450 0 feedthrough
rlabel pdiffusion 45 -1450 45 -1450 0 feedthrough
rlabel pdiffusion 52 -1450 52 -1450 0 cellNo=113
rlabel pdiffusion 59 -1450 59 -1450 0 feedthrough
rlabel pdiffusion 66 -1450 66 -1450 0 feedthrough
rlabel pdiffusion 73 -1450 73 -1450 0 cellNo=637
rlabel pdiffusion 80 -1450 80 -1450 0 feedthrough
rlabel pdiffusion 87 -1450 87 -1450 0 feedthrough
rlabel pdiffusion 94 -1450 94 -1450 0 feedthrough
rlabel pdiffusion 101 -1450 101 -1450 0 cellNo=365
rlabel pdiffusion 108 -1450 108 -1450 0 feedthrough
rlabel pdiffusion 115 -1450 115 -1450 0 cellNo=333
rlabel pdiffusion 122 -1450 122 -1450 0 cellNo=678
rlabel pdiffusion 129 -1450 129 -1450 0 feedthrough
rlabel pdiffusion 136 -1450 136 -1450 0 cellNo=675
rlabel pdiffusion 143 -1450 143 -1450 0 feedthrough
rlabel pdiffusion 150 -1450 150 -1450 0 feedthrough
rlabel pdiffusion 157 -1450 157 -1450 0 cellNo=106
rlabel pdiffusion 164 -1450 164 -1450 0 feedthrough
rlabel pdiffusion 171 -1450 171 -1450 0 feedthrough
rlabel pdiffusion 178 -1450 178 -1450 0 feedthrough
rlabel pdiffusion 185 -1450 185 -1450 0 cellNo=686
rlabel pdiffusion 192 -1450 192 -1450 0 feedthrough
rlabel pdiffusion 199 -1450 199 -1450 0 feedthrough
rlabel pdiffusion 206 -1450 206 -1450 0 feedthrough
rlabel pdiffusion 213 -1450 213 -1450 0 feedthrough
rlabel pdiffusion 220 -1450 220 -1450 0 feedthrough
rlabel pdiffusion 227 -1450 227 -1450 0 feedthrough
rlabel pdiffusion 234 -1450 234 -1450 0 feedthrough
rlabel pdiffusion 241 -1450 241 -1450 0 feedthrough
rlabel pdiffusion 248 -1450 248 -1450 0 feedthrough
rlabel pdiffusion 255 -1450 255 -1450 0 cellNo=282
rlabel pdiffusion 262 -1450 262 -1450 0 feedthrough
rlabel pdiffusion 269 -1450 269 -1450 0 cellNo=479
rlabel pdiffusion 276 -1450 276 -1450 0 feedthrough
rlabel pdiffusion 283 -1450 283 -1450 0 feedthrough
rlabel pdiffusion 290 -1450 290 -1450 0 feedthrough
rlabel pdiffusion 297 -1450 297 -1450 0 feedthrough
rlabel pdiffusion 304 -1450 304 -1450 0 feedthrough
rlabel pdiffusion 311 -1450 311 -1450 0 feedthrough
rlabel pdiffusion 318 -1450 318 -1450 0 feedthrough
rlabel pdiffusion 325 -1450 325 -1450 0 feedthrough
rlabel pdiffusion 332 -1450 332 -1450 0 cellNo=243
rlabel pdiffusion 339 -1450 339 -1450 0 feedthrough
rlabel pdiffusion 346 -1450 346 -1450 0 feedthrough
rlabel pdiffusion 353 -1450 353 -1450 0 feedthrough
rlabel pdiffusion 360 -1450 360 -1450 0 feedthrough
rlabel pdiffusion 367 -1450 367 -1450 0 feedthrough
rlabel pdiffusion 374 -1450 374 -1450 0 feedthrough
rlabel pdiffusion 381 -1450 381 -1450 0 cellNo=417
rlabel pdiffusion 388 -1450 388 -1450 0 feedthrough
rlabel pdiffusion 395 -1450 395 -1450 0 cellNo=150
rlabel pdiffusion 402 -1450 402 -1450 0 cellNo=569
rlabel pdiffusion 409 -1450 409 -1450 0 cellNo=589
rlabel pdiffusion 416 -1450 416 -1450 0 feedthrough
rlabel pdiffusion 423 -1450 423 -1450 0 feedthrough
rlabel pdiffusion 430 -1450 430 -1450 0 cellNo=294
rlabel pdiffusion 437 -1450 437 -1450 0 cellNo=467
rlabel pdiffusion 444 -1450 444 -1450 0 feedthrough
rlabel pdiffusion 451 -1450 451 -1450 0 feedthrough
rlabel pdiffusion 458 -1450 458 -1450 0 feedthrough
rlabel pdiffusion 465 -1450 465 -1450 0 feedthrough
rlabel pdiffusion 472 -1450 472 -1450 0 cellNo=523
rlabel pdiffusion 479 -1450 479 -1450 0 feedthrough
rlabel pdiffusion 486 -1450 486 -1450 0 cellNo=285
rlabel pdiffusion 493 -1450 493 -1450 0 feedthrough
rlabel pdiffusion 500 -1450 500 -1450 0 feedthrough
rlabel pdiffusion 507 -1450 507 -1450 0 cellNo=274
rlabel pdiffusion 514 -1450 514 -1450 0 feedthrough
rlabel pdiffusion 521 -1450 521 -1450 0 feedthrough
rlabel pdiffusion 528 -1450 528 -1450 0 feedthrough
rlabel pdiffusion 535 -1450 535 -1450 0 feedthrough
rlabel pdiffusion 542 -1450 542 -1450 0 feedthrough
rlabel pdiffusion 549 -1450 549 -1450 0 cellNo=542
rlabel pdiffusion 556 -1450 556 -1450 0 feedthrough
rlabel pdiffusion 563 -1450 563 -1450 0 feedthrough
rlabel pdiffusion 570 -1450 570 -1450 0 feedthrough
rlabel pdiffusion 577 -1450 577 -1450 0 feedthrough
rlabel pdiffusion 584 -1450 584 -1450 0 feedthrough
rlabel pdiffusion 591 -1450 591 -1450 0 feedthrough
rlabel pdiffusion 598 -1450 598 -1450 0 feedthrough
rlabel pdiffusion 605 -1450 605 -1450 0 feedthrough
rlabel pdiffusion 612 -1450 612 -1450 0 feedthrough
rlabel pdiffusion 619 -1450 619 -1450 0 feedthrough
rlabel pdiffusion 626 -1450 626 -1450 0 feedthrough
rlabel pdiffusion 633 -1450 633 -1450 0 feedthrough
rlabel pdiffusion 640 -1450 640 -1450 0 feedthrough
rlabel pdiffusion 647 -1450 647 -1450 0 feedthrough
rlabel pdiffusion 654 -1450 654 -1450 0 feedthrough
rlabel pdiffusion 661 -1450 661 -1450 0 feedthrough
rlabel pdiffusion 668 -1450 668 -1450 0 feedthrough
rlabel pdiffusion 675 -1450 675 -1450 0 feedthrough
rlabel pdiffusion 682 -1450 682 -1450 0 feedthrough
rlabel pdiffusion 689 -1450 689 -1450 0 feedthrough
rlabel pdiffusion 696 -1450 696 -1450 0 feedthrough
rlabel pdiffusion 703 -1450 703 -1450 0 feedthrough
rlabel pdiffusion 710 -1450 710 -1450 0 feedthrough
rlabel pdiffusion 717 -1450 717 -1450 0 feedthrough
rlabel pdiffusion 724 -1450 724 -1450 0 feedthrough
rlabel pdiffusion 731 -1450 731 -1450 0 feedthrough
rlabel pdiffusion 738 -1450 738 -1450 0 feedthrough
rlabel pdiffusion 745 -1450 745 -1450 0 feedthrough
rlabel pdiffusion 752 -1450 752 -1450 0 feedthrough
rlabel pdiffusion 766 -1450 766 -1450 0 cellNo=666
rlabel pdiffusion 773 -1450 773 -1450 0 feedthrough
rlabel pdiffusion 780 -1450 780 -1450 0 cellNo=670
rlabel pdiffusion 787 -1450 787 -1450 0 cellNo=385
rlabel pdiffusion 794 -1450 794 -1450 0 cellNo=549
rlabel pdiffusion 801 -1450 801 -1450 0 cellNo=108
rlabel pdiffusion 808 -1450 808 -1450 0 feedthrough
rlabel pdiffusion 815 -1450 815 -1450 0 cellNo=226
rlabel pdiffusion 829 -1450 829 -1450 0 feedthrough
rlabel pdiffusion 836 -1450 836 -1450 0 feedthrough
rlabel pdiffusion 3 -1529 3 -1529 0 cellNo=409
rlabel pdiffusion 10 -1529 10 -1529 0 feedthrough
rlabel pdiffusion 17 -1529 17 -1529 0 feedthrough
rlabel pdiffusion 24 -1529 24 -1529 0 feedthrough
rlabel pdiffusion 31 -1529 31 -1529 0 feedthrough
rlabel pdiffusion 38 -1529 38 -1529 0 feedthrough
rlabel pdiffusion 45 -1529 45 -1529 0 feedthrough
rlabel pdiffusion 52 -1529 52 -1529 0 cellNo=87
rlabel pdiffusion 59 -1529 59 -1529 0 feedthrough
rlabel pdiffusion 66 -1529 66 -1529 0 feedthrough
rlabel pdiffusion 73 -1529 73 -1529 0 cellNo=10
rlabel pdiffusion 80 -1529 80 -1529 0 feedthrough
rlabel pdiffusion 87 -1529 87 -1529 0 feedthrough
rlabel pdiffusion 94 -1529 94 -1529 0 cellNo=691
rlabel pdiffusion 101 -1529 101 -1529 0 feedthrough
rlabel pdiffusion 108 -1529 108 -1529 0 feedthrough
rlabel pdiffusion 115 -1529 115 -1529 0 feedthrough
rlabel pdiffusion 122 -1529 122 -1529 0 feedthrough
rlabel pdiffusion 129 -1529 129 -1529 0 feedthrough
rlabel pdiffusion 136 -1529 136 -1529 0 cellNo=595
rlabel pdiffusion 143 -1529 143 -1529 0 feedthrough
rlabel pdiffusion 150 -1529 150 -1529 0 feedthrough
rlabel pdiffusion 157 -1529 157 -1529 0 feedthrough
rlabel pdiffusion 164 -1529 164 -1529 0 cellNo=2
rlabel pdiffusion 171 -1529 171 -1529 0 cellNo=144
rlabel pdiffusion 178 -1529 178 -1529 0 cellNo=188
rlabel pdiffusion 185 -1529 185 -1529 0 cellNo=578
rlabel pdiffusion 192 -1529 192 -1529 0 feedthrough
rlabel pdiffusion 199 -1529 199 -1529 0 feedthrough
rlabel pdiffusion 206 -1529 206 -1529 0 cellNo=346
rlabel pdiffusion 213 -1529 213 -1529 0 feedthrough
rlabel pdiffusion 220 -1529 220 -1529 0 feedthrough
rlabel pdiffusion 227 -1529 227 -1529 0 feedthrough
rlabel pdiffusion 234 -1529 234 -1529 0 cellNo=480
rlabel pdiffusion 241 -1529 241 -1529 0 cellNo=222
rlabel pdiffusion 248 -1529 248 -1529 0 cellNo=659
rlabel pdiffusion 255 -1529 255 -1529 0 cellNo=657
rlabel pdiffusion 262 -1529 262 -1529 0 feedthrough
rlabel pdiffusion 269 -1529 269 -1529 0 cellNo=245
rlabel pdiffusion 276 -1529 276 -1529 0 feedthrough
rlabel pdiffusion 283 -1529 283 -1529 0 feedthrough
rlabel pdiffusion 290 -1529 290 -1529 0 feedthrough
rlabel pdiffusion 297 -1529 297 -1529 0 feedthrough
rlabel pdiffusion 304 -1529 304 -1529 0 cellNo=461
rlabel pdiffusion 311 -1529 311 -1529 0 feedthrough
rlabel pdiffusion 318 -1529 318 -1529 0 feedthrough
rlabel pdiffusion 325 -1529 325 -1529 0 feedthrough
rlabel pdiffusion 332 -1529 332 -1529 0 cellNo=212
rlabel pdiffusion 339 -1529 339 -1529 0 cellNo=224
rlabel pdiffusion 346 -1529 346 -1529 0 feedthrough
rlabel pdiffusion 353 -1529 353 -1529 0 feedthrough
rlabel pdiffusion 360 -1529 360 -1529 0 cellNo=431
rlabel pdiffusion 367 -1529 367 -1529 0 cellNo=308
rlabel pdiffusion 374 -1529 374 -1529 0 feedthrough
rlabel pdiffusion 381 -1529 381 -1529 0 cellNo=702
rlabel pdiffusion 388 -1529 388 -1529 0 cellNo=502
rlabel pdiffusion 395 -1529 395 -1529 0 feedthrough
rlabel pdiffusion 402 -1529 402 -1529 0 feedthrough
rlabel pdiffusion 409 -1529 409 -1529 0 feedthrough
rlabel pdiffusion 416 -1529 416 -1529 0 cellNo=248
rlabel pdiffusion 423 -1529 423 -1529 0 feedthrough
rlabel pdiffusion 430 -1529 430 -1529 0 feedthrough
rlabel pdiffusion 437 -1529 437 -1529 0 cellNo=492
rlabel pdiffusion 444 -1529 444 -1529 0 feedthrough
rlabel pdiffusion 451 -1529 451 -1529 0 feedthrough
rlabel pdiffusion 458 -1529 458 -1529 0 feedthrough
rlabel pdiffusion 465 -1529 465 -1529 0 feedthrough
rlabel pdiffusion 472 -1529 472 -1529 0 feedthrough
rlabel pdiffusion 479 -1529 479 -1529 0 feedthrough
rlabel pdiffusion 486 -1529 486 -1529 0 feedthrough
rlabel pdiffusion 493 -1529 493 -1529 0 feedthrough
rlabel pdiffusion 500 -1529 500 -1529 0 feedthrough
rlabel pdiffusion 507 -1529 507 -1529 0 feedthrough
rlabel pdiffusion 514 -1529 514 -1529 0 feedthrough
rlabel pdiffusion 521 -1529 521 -1529 0 cellNo=668
rlabel pdiffusion 528 -1529 528 -1529 0 feedthrough
rlabel pdiffusion 535 -1529 535 -1529 0 feedthrough
rlabel pdiffusion 542 -1529 542 -1529 0 feedthrough
rlabel pdiffusion 549 -1529 549 -1529 0 feedthrough
rlabel pdiffusion 556 -1529 556 -1529 0 feedthrough
rlabel pdiffusion 563 -1529 563 -1529 0 feedthrough
rlabel pdiffusion 570 -1529 570 -1529 0 feedthrough
rlabel pdiffusion 577 -1529 577 -1529 0 feedthrough
rlabel pdiffusion 584 -1529 584 -1529 0 feedthrough
rlabel pdiffusion 591 -1529 591 -1529 0 feedthrough
rlabel pdiffusion 598 -1529 598 -1529 0 cellNo=649
rlabel pdiffusion 605 -1529 605 -1529 0 feedthrough
rlabel pdiffusion 612 -1529 612 -1529 0 feedthrough
rlabel pdiffusion 619 -1529 619 -1529 0 cellNo=487
rlabel pdiffusion 626 -1529 626 -1529 0 feedthrough
rlabel pdiffusion 633 -1529 633 -1529 0 feedthrough
rlabel pdiffusion 640 -1529 640 -1529 0 feedthrough
rlabel pdiffusion 647 -1529 647 -1529 0 feedthrough
rlabel pdiffusion 654 -1529 654 -1529 0 feedthrough
rlabel pdiffusion 661 -1529 661 -1529 0 feedthrough
rlabel pdiffusion 668 -1529 668 -1529 0 feedthrough
rlabel pdiffusion 675 -1529 675 -1529 0 feedthrough
rlabel pdiffusion 682 -1529 682 -1529 0 feedthrough
rlabel pdiffusion 689 -1529 689 -1529 0 feedthrough
rlabel pdiffusion 696 -1529 696 -1529 0 feedthrough
rlabel pdiffusion 703 -1529 703 -1529 0 feedthrough
rlabel pdiffusion 710 -1529 710 -1529 0 feedthrough
rlabel pdiffusion 717 -1529 717 -1529 0 feedthrough
rlabel pdiffusion 724 -1529 724 -1529 0 feedthrough
rlabel pdiffusion 731 -1529 731 -1529 0 feedthrough
rlabel pdiffusion 738 -1529 738 -1529 0 feedthrough
rlabel pdiffusion 745 -1529 745 -1529 0 feedthrough
rlabel pdiffusion 752 -1529 752 -1529 0 feedthrough
rlabel pdiffusion 3 -1608 3 -1608 0 cellNo=210
rlabel pdiffusion 10 -1608 10 -1608 0 cellNo=252
rlabel pdiffusion 17 -1608 17 -1608 0 feedthrough
rlabel pdiffusion 24 -1608 24 -1608 0 feedthrough
rlabel pdiffusion 31 -1608 31 -1608 0 cellNo=704
rlabel pdiffusion 38 -1608 38 -1608 0 feedthrough
rlabel pdiffusion 45 -1608 45 -1608 0 cellNo=503
rlabel pdiffusion 52 -1608 52 -1608 0 feedthrough
rlabel pdiffusion 59 -1608 59 -1608 0 feedthrough
rlabel pdiffusion 66 -1608 66 -1608 0 feedthrough
rlabel pdiffusion 73 -1608 73 -1608 0 feedthrough
rlabel pdiffusion 80 -1608 80 -1608 0 cellNo=532
rlabel pdiffusion 87 -1608 87 -1608 0 cellNo=719
rlabel pdiffusion 94 -1608 94 -1608 0 feedthrough
rlabel pdiffusion 101 -1608 101 -1608 0 cellNo=37
rlabel pdiffusion 108 -1608 108 -1608 0 feedthrough
rlabel pdiffusion 115 -1608 115 -1608 0 cellNo=679
rlabel pdiffusion 122 -1608 122 -1608 0 feedthrough
rlabel pdiffusion 129 -1608 129 -1608 0 feedthrough
rlabel pdiffusion 136 -1608 136 -1608 0 cellNo=416
rlabel pdiffusion 143 -1608 143 -1608 0 cellNo=530
rlabel pdiffusion 150 -1608 150 -1608 0 cellNo=577
rlabel pdiffusion 157 -1608 157 -1608 0 feedthrough
rlabel pdiffusion 164 -1608 164 -1608 0 feedthrough
rlabel pdiffusion 171 -1608 171 -1608 0 feedthrough
rlabel pdiffusion 178 -1608 178 -1608 0 feedthrough
rlabel pdiffusion 185 -1608 185 -1608 0 feedthrough
rlabel pdiffusion 192 -1608 192 -1608 0 cellNo=638
rlabel pdiffusion 199 -1608 199 -1608 0 feedthrough
rlabel pdiffusion 206 -1608 206 -1608 0 feedthrough
rlabel pdiffusion 213 -1608 213 -1608 0 feedthrough
rlabel pdiffusion 220 -1608 220 -1608 0 cellNo=626
rlabel pdiffusion 227 -1608 227 -1608 0 feedthrough
rlabel pdiffusion 234 -1608 234 -1608 0 cellNo=693
rlabel pdiffusion 241 -1608 241 -1608 0 feedthrough
rlabel pdiffusion 248 -1608 248 -1608 0 feedthrough
rlabel pdiffusion 255 -1608 255 -1608 0 feedthrough
rlabel pdiffusion 262 -1608 262 -1608 0 feedthrough
rlabel pdiffusion 269 -1608 269 -1608 0 feedthrough
rlabel pdiffusion 276 -1608 276 -1608 0 cellNo=266
rlabel pdiffusion 283 -1608 283 -1608 0 feedthrough
rlabel pdiffusion 290 -1608 290 -1608 0 feedthrough
rlabel pdiffusion 297 -1608 297 -1608 0 feedthrough
rlabel pdiffusion 304 -1608 304 -1608 0 cellNo=216
rlabel pdiffusion 311 -1608 311 -1608 0 cellNo=382
rlabel pdiffusion 318 -1608 318 -1608 0 cellNo=425
rlabel pdiffusion 325 -1608 325 -1608 0 feedthrough
rlabel pdiffusion 332 -1608 332 -1608 0 feedthrough
rlabel pdiffusion 339 -1608 339 -1608 0 cellNo=495
rlabel pdiffusion 346 -1608 346 -1608 0 feedthrough
rlabel pdiffusion 353 -1608 353 -1608 0 feedthrough
rlabel pdiffusion 360 -1608 360 -1608 0 cellNo=327
rlabel pdiffusion 367 -1608 367 -1608 0 cellNo=364
rlabel pdiffusion 374 -1608 374 -1608 0 feedthrough
rlabel pdiffusion 381 -1608 381 -1608 0 feedthrough
rlabel pdiffusion 388 -1608 388 -1608 0 feedthrough
rlabel pdiffusion 395 -1608 395 -1608 0 feedthrough
rlabel pdiffusion 402 -1608 402 -1608 0 feedthrough
rlabel pdiffusion 409 -1608 409 -1608 0 cellNo=313
rlabel pdiffusion 416 -1608 416 -1608 0 feedthrough
rlabel pdiffusion 423 -1608 423 -1608 0 feedthrough
rlabel pdiffusion 430 -1608 430 -1608 0 feedthrough
rlabel pdiffusion 437 -1608 437 -1608 0 cellNo=76
rlabel pdiffusion 444 -1608 444 -1608 0 cellNo=155
rlabel pdiffusion 451 -1608 451 -1608 0 feedthrough
rlabel pdiffusion 458 -1608 458 -1608 0 feedthrough
rlabel pdiffusion 465 -1608 465 -1608 0 feedthrough
rlabel pdiffusion 472 -1608 472 -1608 0 cellNo=389
rlabel pdiffusion 479 -1608 479 -1608 0 feedthrough
rlabel pdiffusion 486 -1608 486 -1608 0 cellNo=570
rlabel pdiffusion 493 -1608 493 -1608 0 feedthrough
rlabel pdiffusion 500 -1608 500 -1608 0 feedthrough
rlabel pdiffusion 507 -1608 507 -1608 0 feedthrough
rlabel pdiffusion 514 -1608 514 -1608 0 feedthrough
rlabel pdiffusion 521 -1608 521 -1608 0 feedthrough
rlabel pdiffusion 528 -1608 528 -1608 0 feedthrough
rlabel pdiffusion 535 -1608 535 -1608 0 feedthrough
rlabel pdiffusion 542 -1608 542 -1608 0 feedthrough
rlabel pdiffusion 549 -1608 549 -1608 0 feedthrough
rlabel pdiffusion 556 -1608 556 -1608 0 cellNo=30
rlabel pdiffusion 563 -1608 563 -1608 0 feedthrough
rlabel pdiffusion 570 -1608 570 -1608 0 feedthrough
rlabel pdiffusion 577 -1608 577 -1608 0 feedthrough
rlabel pdiffusion 584 -1608 584 -1608 0 feedthrough
rlabel pdiffusion 591 -1608 591 -1608 0 feedthrough
rlabel pdiffusion 598 -1608 598 -1608 0 feedthrough
rlabel pdiffusion 605 -1608 605 -1608 0 feedthrough
rlabel pdiffusion 612 -1608 612 -1608 0 feedthrough
rlabel pdiffusion 619 -1608 619 -1608 0 feedthrough
rlabel pdiffusion 626 -1608 626 -1608 0 feedthrough
rlabel pdiffusion 633 -1608 633 -1608 0 feedthrough
rlabel pdiffusion 640 -1608 640 -1608 0 feedthrough
rlabel pdiffusion 647 -1608 647 -1608 0 feedthrough
rlabel pdiffusion 654 -1608 654 -1608 0 feedthrough
rlabel pdiffusion 661 -1608 661 -1608 0 feedthrough
rlabel pdiffusion 668 -1608 668 -1608 0 feedthrough
rlabel pdiffusion 675 -1608 675 -1608 0 feedthrough
rlabel pdiffusion 682 -1608 682 -1608 0 feedthrough
rlabel pdiffusion 10 -1677 10 -1677 0 feedthrough
rlabel pdiffusion 17 -1677 17 -1677 0 feedthrough
rlabel pdiffusion 24 -1677 24 -1677 0 feedthrough
rlabel pdiffusion 31 -1677 31 -1677 0 cellNo=183
rlabel pdiffusion 38 -1677 38 -1677 0 feedthrough
rlabel pdiffusion 45 -1677 45 -1677 0 cellNo=634
rlabel pdiffusion 52 -1677 52 -1677 0 cellNo=74
rlabel pdiffusion 59 -1677 59 -1677 0 feedthrough
rlabel pdiffusion 66 -1677 66 -1677 0 feedthrough
rlabel pdiffusion 73 -1677 73 -1677 0 feedthrough
rlabel pdiffusion 80 -1677 80 -1677 0 feedthrough
rlabel pdiffusion 87 -1677 87 -1677 0 cellNo=396
rlabel pdiffusion 94 -1677 94 -1677 0 feedthrough
rlabel pdiffusion 101 -1677 101 -1677 0 cellNo=614
rlabel pdiffusion 108 -1677 108 -1677 0 cellNo=518
rlabel pdiffusion 115 -1677 115 -1677 0 cellNo=20
rlabel pdiffusion 122 -1677 122 -1677 0 feedthrough
rlabel pdiffusion 129 -1677 129 -1677 0 feedthrough
rlabel pdiffusion 136 -1677 136 -1677 0 feedthrough
rlabel pdiffusion 143 -1677 143 -1677 0 cellNo=11
rlabel pdiffusion 150 -1677 150 -1677 0 feedthrough
rlabel pdiffusion 157 -1677 157 -1677 0 feedthrough
rlabel pdiffusion 164 -1677 164 -1677 0 feedthrough
rlabel pdiffusion 171 -1677 171 -1677 0 cellNo=349
rlabel pdiffusion 178 -1677 178 -1677 0 feedthrough
rlabel pdiffusion 185 -1677 185 -1677 0 cellNo=684
rlabel pdiffusion 192 -1677 192 -1677 0 cellNo=594
rlabel pdiffusion 199 -1677 199 -1677 0 feedthrough
rlabel pdiffusion 206 -1677 206 -1677 0 feedthrough
rlabel pdiffusion 213 -1677 213 -1677 0 feedthrough
rlabel pdiffusion 220 -1677 220 -1677 0 feedthrough
rlabel pdiffusion 227 -1677 227 -1677 0 feedthrough
rlabel pdiffusion 234 -1677 234 -1677 0 cellNo=400
rlabel pdiffusion 241 -1677 241 -1677 0 cellNo=204
rlabel pdiffusion 248 -1677 248 -1677 0 feedthrough
rlabel pdiffusion 255 -1677 255 -1677 0 feedthrough
rlabel pdiffusion 262 -1677 262 -1677 0 cellNo=522
rlabel pdiffusion 269 -1677 269 -1677 0 feedthrough
rlabel pdiffusion 276 -1677 276 -1677 0 feedthrough
rlabel pdiffusion 283 -1677 283 -1677 0 feedthrough
rlabel pdiffusion 290 -1677 290 -1677 0 cellNo=644
rlabel pdiffusion 297 -1677 297 -1677 0 cellNo=654
rlabel pdiffusion 304 -1677 304 -1677 0 cellNo=362
rlabel pdiffusion 311 -1677 311 -1677 0 feedthrough
rlabel pdiffusion 318 -1677 318 -1677 0 feedthrough
rlabel pdiffusion 325 -1677 325 -1677 0 feedthrough
rlabel pdiffusion 332 -1677 332 -1677 0 cellNo=680
rlabel pdiffusion 339 -1677 339 -1677 0 cellNo=18
rlabel pdiffusion 346 -1677 346 -1677 0 feedthrough
rlabel pdiffusion 353 -1677 353 -1677 0 cellNo=617
rlabel pdiffusion 360 -1677 360 -1677 0 cellNo=145
rlabel pdiffusion 367 -1677 367 -1677 0 cellNo=309
rlabel pdiffusion 374 -1677 374 -1677 0 cellNo=233
rlabel pdiffusion 381 -1677 381 -1677 0 feedthrough
rlabel pdiffusion 388 -1677 388 -1677 0 cellNo=696
rlabel pdiffusion 395 -1677 395 -1677 0 feedthrough
rlabel pdiffusion 402 -1677 402 -1677 0 feedthrough
rlabel pdiffusion 409 -1677 409 -1677 0 feedthrough
rlabel pdiffusion 416 -1677 416 -1677 0 feedthrough
rlabel pdiffusion 423 -1677 423 -1677 0 feedthrough
rlabel pdiffusion 430 -1677 430 -1677 0 feedthrough
rlabel pdiffusion 437 -1677 437 -1677 0 feedthrough
rlabel pdiffusion 444 -1677 444 -1677 0 feedthrough
rlabel pdiffusion 451 -1677 451 -1677 0 feedthrough
rlabel pdiffusion 458 -1677 458 -1677 0 feedthrough
rlabel pdiffusion 465 -1677 465 -1677 0 feedthrough
rlabel pdiffusion 472 -1677 472 -1677 0 feedthrough
rlabel pdiffusion 479 -1677 479 -1677 0 feedthrough
rlabel pdiffusion 486 -1677 486 -1677 0 feedthrough
rlabel pdiffusion 493 -1677 493 -1677 0 feedthrough
rlabel pdiffusion 500 -1677 500 -1677 0 feedthrough
rlabel pdiffusion 507 -1677 507 -1677 0 feedthrough
rlabel pdiffusion 514 -1677 514 -1677 0 feedthrough
rlabel pdiffusion 521 -1677 521 -1677 0 feedthrough
rlabel pdiffusion 528 -1677 528 -1677 0 feedthrough
rlabel pdiffusion 535 -1677 535 -1677 0 feedthrough
rlabel pdiffusion 542 -1677 542 -1677 0 feedthrough
rlabel pdiffusion 549 -1677 549 -1677 0 feedthrough
rlabel pdiffusion 556 -1677 556 -1677 0 feedthrough
rlabel pdiffusion 563 -1677 563 -1677 0 feedthrough
rlabel pdiffusion 570 -1677 570 -1677 0 feedthrough
rlabel pdiffusion 577 -1677 577 -1677 0 feedthrough
rlabel pdiffusion 584 -1677 584 -1677 0 feedthrough
rlabel pdiffusion 591 -1677 591 -1677 0 feedthrough
rlabel pdiffusion 598 -1677 598 -1677 0 feedthrough
rlabel pdiffusion 612 -1677 612 -1677 0 feedthrough
rlabel pdiffusion 619 -1677 619 -1677 0 cellNo=572
rlabel pdiffusion 647 -1677 647 -1677 0 cellNo=366
rlabel pdiffusion 661 -1677 661 -1677 0 feedthrough
rlabel pdiffusion 675 -1677 675 -1677 0 cellNo=517
rlabel pdiffusion 682 -1677 682 -1677 0 feedthrough
rlabel pdiffusion 10 -1734 10 -1734 0 feedthrough
rlabel pdiffusion 17 -1734 17 -1734 0 feedthrough
rlabel pdiffusion 24 -1734 24 -1734 0 feedthrough
rlabel pdiffusion 31 -1734 31 -1734 0 cellNo=669
rlabel pdiffusion 38 -1734 38 -1734 0 cellNo=551
rlabel pdiffusion 45 -1734 45 -1734 0 feedthrough
rlabel pdiffusion 52 -1734 52 -1734 0 feedthrough
rlabel pdiffusion 59 -1734 59 -1734 0 feedthrough
rlabel pdiffusion 66 -1734 66 -1734 0 feedthrough
rlabel pdiffusion 73 -1734 73 -1734 0 feedthrough
rlabel pdiffusion 80 -1734 80 -1734 0 feedthrough
rlabel pdiffusion 87 -1734 87 -1734 0 feedthrough
rlabel pdiffusion 94 -1734 94 -1734 0 cellNo=588
rlabel pdiffusion 101 -1734 101 -1734 0 cellNo=56
rlabel pdiffusion 108 -1734 108 -1734 0 feedthrough
rlabel pdiffusion 115 -1734 115 -1734 0 feedthrough
rlabel pdiffusion 122 -1734 122 -1734 0 cellNo=643
rlabel pdiffusion 129 -1734 129 -1734 0 cellNo=372
rlabel pdiffusion 136 -1734 136 -1734 0 feedthrough
rlabel pdiffusion 143 -1734 143 -1734 0 cellNo=187
rlabel pdiffusion 150 -1734 150 -1734 0 cellNo=241
rlabel pdiffusion 157 -1734 157 -1734 0 cellNo=486
rlabel pdiffusion 164 -1734 164 -1734 0 feedthrough
rlabel pdiffusion 171 -1734 171 -1734 0 feedthrough
rlabel pdiffusion 178 -1734 178 -1734 0 cellNo=139
rlabel pdiffusion 185 -1734 185 -1734 0 cellNo=630
rlabel pdiffusion 192 -1734 192 -1734 0 feedthrough
rlabel pdiffusion 199 -1734 199 -1734 0 feedthrough
rlabel pdiffusion 206 -1734 206 -1734 0 cellNo=246
rlabel pdiffusion 213 -1734 213 -1734 0 feedthrough
rlabel pdiffusion 220 -1734 220 -1734 0 feedthrough
rlabel pdiffusion 227 -1734 227 -1734 0 feedthrough
rlabel pdiffusion 234 -1734 234 -1734 0 feedthrough
rlabel pdiffusion 241 -1734 241 -1734 0 cellNo=205
rlabel pdiffusion 248 -1734 248 -1734 0 cellNo=97
rlabel pdiffusion 255 -1734 255 -1734 0 cellNo=624
rlabel pdiffusion 262 -1734 262 -1734 0 feedthrough
rlabel pdiffusion 269 -1734 269 -1734 0 cellNo=607
rlabel pdiffusion 276 -1734 276 -1734 0 feedthrough
rlabel pdiffusion 283 -1734 283 -1734 0 feedthrough
rlabel pdiffusion 290 -1734 290 -1734 0 cellNo=698
rlabel pdiffusion 297 -1734 297 -1734 0 feedthrough
rlabel pdiffusion 304 -1734 304 -1734 0 feedthrough
rlabel pdiffusion 311 -1734 311 -1734 0 cellNo=677
rlabel pdiffusion 318 -1734 318 -1734 0 cellNo=652
rlabel pdiffusion 325 -1734 325 -1734 0 feedthrough
rlabel pdiffusion 332 -1734 332 -1734 0 feedthrough
rlabel pdiffusion 339 -1734 339 -1734 0 cellNo=688
rlabel pdiffusion 346 -1734 346 -1734 0 feedthrough
rlabel pdiffusion 353 -1734 353 -1734 0 cellNo=575
rlabel pdiffusion 360 -1734 360 -1734 0 cellNo=433
rlabel pdiffusion 367 -1734 367 -1734 0 feedthrough
rlabel pdiffusion 374 -1734 374 -1734 0 cellNo=697
rlabel pdiffusion 381 -1734 381 -1734 0 feedthrough
rlabel pdiffusion 395 -1734 395 -1734 0 feedthrough
rlabel pdiffusion 402 -1734 402 -1734 0 feedthrough
rlabel pdiffusion 409 -1734 409 -1734 0 feedthrough
rlabel pdiffusion 416 -1734 416 -1734 0 feedthrough
rlabel pdiffusion 423 -1734 423 -1734 0 feedthrough
rlabel pdiffusion 430 -1734 430 -1734 0 feedthrough
rlabel pdiffusion 437 -1734 437 -1734 0 feedthrough
rlabel pdiffusion 444 -1734 444 -1734 0 cellNo=421
rlabel pdiffusion 458 -1734 458 -1734 0 cellNo=608
rlabel pdiffusion 465 -1734 465 -1734 0 feedthrough
rlabel pdiffusion 472 -1734 472 -1734 0 feedthrough
rlabel pdiffusion 479 -1734 479 -1734 0 feedthrough
rlabel pdiffusion 486 -1734 486 -1734 0 feedthrough
rlabel pdiffusion 493 -1734 493 -1734 0 feedthrough
rlabel pdiffusion 500 -1734 500 -1734 0 feedthrough
rlabel pdiffusion 521 -1734 521 -1734 0 feedthrough
rlabel pdiffusion 528 -1734 528 -1734 0 feedthrough
rlabel pdiffusion 556 -1734 556 -1734 0 feedthrough
rlabel pdiffusion 577 -1734 577 -1734 0 cellNo=429
rlabel pdiffusion 619 -1734 619 -1734 0 feedthrough
rlabel pdiffusion 654 -1734 654 -1734 0 feedthrough
rlabel pdiffusion 668 -1734 668 -1734 0 cellNo=550
rlabel pdiffusion 675 -1734 675 -1734 0 feedthrough
rlabel pdiffusion 38 -1775 38 -1775 0 feedthrough
rlabel pdiffusion 52 -1775 52 -1775 0 feedthrough
rlabel pdiffusion 59 -1775 59 -1775 0 cellNo=636
rlabel pdiffusion 66 -1775 66 -1775 0 feedthrough
rlabel pdiffusion 73 -1775 73 -1775 0 feedthrough
rlabel pdiffusion 87 -1775 87 -1775 0 feedthrough
rlabel pdiffusion 94 -1775 94 -1775 0 feedthrough
rlabel pdiffusion 101 -1775 101 -1775 0 cellNo=4
rlabel pdiffusion 108 -1775 108 -1775 0 cellNo=169
rlabel pdiffusion 115 -1775 115 -1775 0 cellNo=647
rlabel pdiffusion 122 -1775 122 -1775 0 cellNo=526
rlabel pdiffusion 129 -1775 129 -1775 0 feedthrough
rlabel pdiffusion 136 -1775 136 -1775 0 feedthrough
rlabel pdiffusion 143 -1775 143 -1775 0 feedthrough
rlabel pdiffusion 150 -1775 150 -1775 0 cellNo=622
rlabel pdiffusion 157 -1775 157 -1775 0 cellNo=713
rlabel pdiffusion 164 -1775 164 -1775 0 cellNo=512
rlabel pdiffusion 171 -1775 171 -1775 0 cellNo=176
rlabel pdiffusion 178 -1775 178 -1775 0 cellNo=86
rlabel pdiffusion 185 -1775 185 -1775 0 cellNo=456
rlabel pdiffusion 192 -1775 192 -1775 0 feedthrough
rlabel pdiffusion 199 -1775 199 -1775 0 feedthrough
rlabel pdiffusion 206 -1775 206 -1775 0 cellNo=695
rlabel pdiffusion 213 -1775 213 -1775 0 cellNo=445
rlabel pdiffusion 220 -1775 220 -1775 0 feedthrough
rlabel pdiffusion 227 -1775 227 -1775 0 feedthrough
rlabel pdiffusion 234 -1775 234 -1775 0 feedthrough
rlabel pdiffusion 241 -1775 241 -1775 0 feedthrough
rlabel pdiffusion 255 -1775 255 -1775 0 cellNo=134
rlabel pdiffusion 262 -1775 262 -1775 0 feedthrough
rlabel pdiffusion 269 -1775 269 -1775 0 feedthrough
rlabel pdiffusion 276 -1775 276 -1775 0 cellNo=283
rlabel pdiffusion 290 -1775 290 -1775 0 feedthrough
rlabel pdiffusion 297 -1775 297 -1775 0 feedthrough
rlabel pdiffusion 311 -1775 311 -1775 0 feedthrough
rlabel pdiffusion 318 -1775 318 -1775 0 feedthrough
rlabel pdiffusion 325 -1775 325 -1775 0 feedthrough
rlabel pdiffusion 332 -1775 332 -1775 0 cellNo=685
rlabel pdiffusion 339 -1775 339 -1775 0 feedthrough
rlabel pdiffusion 346 -1775 346 -1775 0 feedthrough
rlabel pdiffusion 353 -1775 353 -1775 0 feedthrough
rlabel pdiffusion 367 -1775 367 -1775 0 feedthrough
rlabel pdiffusion 381 -1775 381 -1775 0 cellNo=618
rlabel pdiffusion 402 -1775 402 -1775 0 cellNo=424
rlabel pdiffusion 416 -1775 416 -1775 0 cellNo=599
rlabel pdiffusion 423 -1775 423 -1775 0 feedthrough
rlabel pdiffusion 430 -1775 430 -1775 0 feedthrough
rlabel pdiffusion 451 -1775 451 -1775 0 cellNo=533
rlabel pdiffusion 458 -1775 458 -1775 0 cellNo=562
rlabel pdiffusion 465 -1775 465 -1775 0 feedthrough
rlabel pdiffusion 472 -1775 472 -1775 0 feedthrough
rlabel pdiffusion 479 -1775 479 -1775 0 feedthrough
rlabel pdiffusion 486 -1775 486 -1775 0 cellNo=540
rlabel pdiffusion 500 -1775 500 -1775 0 cellNo=603
rlabel pdiffusion 514 -1775 514 -1775 0 feedthrough
rlabel pdiffusion 521 -1775 521 -1775 0 feedthrough
rlabel pdiffusion 528 -1775 528 -1775 0 feedthrough
rlabel pdiffusion 535 -1775 535 -1775 0 feedthrough
rlabel pdiffusion 542 -1775 542 -1775 0 cellNo=370
rlabel pdiffusion 549 -1775 549 -1775 0 feedthrough
rlabel pdiffusion 563 -1775 563 -1775 0 cellNo=201
rlabel pdiffusion 612 -1775 612 -1775 0 cellNo=190
rlabel pdiffusion 619 -1775 619 -1775 0 feedthrough
rlabel pdiffusion 633 -1775 633 -1775 0 feedthrough
rlabel pdiffusion 52 -1804 52 -1804 0 feedthrough
rlabel pdiffusion 59 -1804 59 -1804 0 cellNo=581
rlabel pdiffusion 87 -1804 87 -1804 0 cellNo=44
rlabel pdiffusion 101 -1804 101 -1804 0 cellNo=655
rlabel pdiffusion 108 -1804 108 -1804 0 cellNo=683
rlabel pdiffusion 115 -1804 115 -1804 0 cellNo=469
rlabel pdiffusion 122 -1804 122 -1804 0 cellNo=470
rlabel pdiffusion 129 -1804 129 -1804 0 cellNo=284
rlabel pdiffusion 136 -1804 136 -1804 0 cellNo=281
rlabel pdiffusion 143 -1804 143 -1804 0 cellNo=714
rlabel pdiffusion 150 -1804 150 -1804 0 feedthrough
rlabel pdiffusion 157 -1804 157 -1804 0 feedthrough
rlabel pdiffusion 171 -1804 171 -1804 0 cellNo=158
rlabel pdiffusion 178 -1804 178 -1804 0 cellNo=564
rlabel pdiffusion 185 -1804 185 -1804 0 cellNo=497
rlabel pdiffusion 206 -1804 206 -1804 0 feedthrough
rlabel pdiffusion 234 -1804 234 -1804 0 feedthrough
rlabel pdiffusion 248 -1804 248 -1804 0 cellNo=718
rlabel pdiffusion 255 -1804 255 -1804 0 cellNo=242
rlabel pdiffusion 262 -1804 262 -1804 0 cellNo=407
rlabel pdiffusion 269 -1804 269 -1804 0 cellNo=646
rlabel pdiffusion 311 -1804 311 -1804 0 cellNo=92
rlabel pdiffusion 353 -1804 353 -1804 0 feedthrough
rlabel pdiffusion 374 -1804 374 -1804 0 cellNo=405
rlabel pdiffusion 388 -1804 388 -1804 0 cellNo=3
rlabel pdiffusion 409 -1804 409 -1804 0 cellNo=136
rlabel pdiffusion 416 -1804 416 -1804 0 cellNo=707
rlabel pdiffusion 465 -1804 465 -1804 0 cellNo=443
rlabel pdiffusion 472 -1804 472 -1804 0 feedthrough
rlabel pdiffusion 479 -1804 479 -1804 0 cellNo=442
rlabel pdiffusion 500 -1804 500 -1804 0 cellNo=635
rlabel pdiffusion 521 -1804 521 -1804 0 feedthrough
rlabel pdiffusion 528 -1804 528 -1804 0 cellNo=671
rlabel pdiffusion 640 -1804 640 -1804 0 cellNo=612
rlabel polysilicon 47 -14 47 -14 0 4
rlabel polysilicon 58 -8 58 -8 0 1
rlabel polysilicon 93 -8 93 -8 0 1
rlabel polysilicon 93 -14 93 -14 0 3
rlabel polysilicon 114 -8 114 -8 0 1
rlabel polysilicon 114 -14 114 -14 0 3
rlabel polysilicon 124 -8 124 -8 0 2
rlabel polysilicon 128 -8 128 -8 0 1
rlabel polysilicon 128 -14 128 -14 0 3
rlabel polysilicon 135 -8 135 -8 0 1
rlabel polysilicon 142 -8 142 -8 0 1
rlabel polysilicon 152 -8 152 -8 0 2
rlabel polysilicon 156 -8 156 -8 0 1
rlabel polysilicon 163 -8 163 -8 0 1
rlabel polysilicon 163 -14 163 -14 0 3
rlabel polysilicon 170 -8 170 -8 0 1
rlabel polysilicon 170 -14 170 -14 0 3
rlabel polysilicon 177 -8 177 -8 0 1
rlabel polysilicon 177 -14 177 -14 0 3
rlabel polysilicon 184 -8 184 -8 0 1
rlabel polysilicon 184 -14 184 -14 0 3
rlabel polysilicon 191 -8 191 -8 0 1
rlabel polysilicon 198 -8 198 -8 0 1
rlabel polysilicon 198 -14 198 -14 0 3
rlabel polysilicon 205 -8 205 -8 0 1
rlabel polysilicon 205 -14 205 -14 0 3
rlabel polysilicon 212 -8 212 -8 0 1
rlabel polysilicon 212 -14 212 -14 0 3
rlabel polysilicon 222 -14 222 -14 0 4
rlabel polysilicon 226 -14 226 -14 0 3
rlabel polysilicon 236 -8 236 -8 0 2
rlabel polysilicon 233 -14 233 -14 0 3
rlabel polysilicon 240 -8 240 -8 0 1
rlabel polysilicon 240 -14 240 -14 0 3
rlabel polysilicon 257 -8 257 -8 0 2
rlabel polysilicon 261 -8 261 -8 0 1
rlabel polysilicon 261 -14 261 -14 0 3
rlabel polysilicon 289 -14 289 -14 0 3
rlabel polysilicon 338 -8 338 -8 0 1
rlabel polysilicon 338 -14 338 -14 0 3
rlabel polysilicon 44 -35 44 -35 0 1
rlabel polysilicon 51 -41 51 -41 0 3
rlabel polysilicon 72 -35 72 -35 0 1
rlabel polysilicon 72 -41 72 -41 0 3
rlabel polysilicon 79 -35 79 -35 0 1
rlabel polysilicon 93 -35 93 -35 0 1
rlabel polysilicon 93 -41 93 -41 0 3
rlabel polysilicon 103 -35 103 -35 0 2
rlabel polysilicon 107 -41 107 -41 0 3
rlabel polysilicon 117 -41 117 -41 0 4
rlabel polysilicon 124 -35 124 -35 0 2
rlabel polysilicon 128 -35 128 -35 0 1
rlabel polysilicon 131 -35 131 -35 0 2
rlabel polysilicon 135 -35 135 -35 0 1
rlabel polysilicon 135 -41 135 -41 0 3
rlabel polysilicon 142 -35 142 -35 0 1
rlabel polysilicon 149 -35 149 -35 0 1
rlabel polysilicon 156 -41 156 -41 0 3
rlabel polysilicon 163 -35 163 -35 0 1
rlabel polysilicon 170 -35 170 -35 0 1
rlabel polysilicon 170 -41 170 -41 0 3
rlabel polysilicon 177 -35 177 -35 0 1
rlabel polysilicon 177 -41 177 -41 0 3
rlabel polysilicon 184 -35 184 -35 0 1
rlabel polysilicon 184 -41 184 -41 0 3
rlabel polysilicon 191 -35 191 -35 0 1
rlabel polysilicon 191 -41 191 -41 0 3
rlabel polysilicon 198 -35 198 -35 0 1
rlabel polysilicon 198 -41 198 -41 0 3
rlabel polysilicon 205 -35 205 -35 0 1
rlabel polysilicon 205 -41 205 -41 0 3
rlabel polysilicon 208 -41 208 -41 0 4
rlabel polysilicon 212 -35 212 -35 0 1
rlabel polysilicon 212 -41 212 -41 0 3
rlabel polysilicon 219 -35 219 -35 0 1
rlabel polysilicon 219 -41 219 -41 0 3
rlabel polysilicon 226 -35 226 -35 0 1
rlabel polysilicon 226 -41 226 -41 0 3
rlabel polysilicon 233 -35 233 -35 0 1
rlabel polysilicon 233 -41 233 -41 0 3
rlabel polysilicon 240 -35 240 -35 0 1
rlabel polysilicon 240 -41 240 -41 0 3
rlabel polysilicon 247 -35 247 -35 0 1
rlabel polysilicon 247 -41 247 -41 0 3
rlabel polysilicon 254 -35 254 -35 0 1
rlabel polysilicon 254 -41 254 -41 0 3
rlabel polysilicon 271 -35 271 -35 0 2
rlabel polysilicon 271 -41 271 -41 0 4
rlabel polysilicon 275 -35 275 -35 0 1
rlabel polysilicon 275 -41 275 -41 0 3
rlabel polysilicon 282 -35 282 -35 0 1
rlabel polysilicon 285 -35 285 -35 0 2
rlabel polysilicon 292 -41 292 -41 0 4
rlabel polysilicon 296 -35 296 -35 0 1
rlabel polysilicon 296 -41 296 -41 0 3
rlabel polysilicon 313 -35 313 -35 0 2
rlabel polysilicon 317 -35 317 -35 0 1
rlabel polysilicon 317 -41 317 -41 0 3
rlabel polysilicon 324 -35 324 -35 0 1
rlabel polysilicon 324 -41 324 -41 0 3
rlabel polysilicon 334 -35 334 -35 0 2
rlabel polysilicon 338 -35 338 -35 0 1
rlabel polysilicon 338 -41 338 -41 0 3
rlabel polysilicon 345 -35 345 -35 0 1
rlabel polysilicon 345 -41 345 -41 0 3
rlabel polysilicon 352 -35 352 -35 0 1
rlabel polysilicon 352 -41 352 -41 0 3
rlabel polysilicon 387 -35 387 -35 0 1
rlabel polysilicon 387 -41 387 -41 0 3
rlabel polysilicon 404 -41 404 -41 0 4
rlabel polysilicon 16 -70 16 -70 0 1
rlabel polysilicon 16 -76 16 -76 0 3
rlabel polysilicon 23 -70 23 -70 0 1
rlabel polysilicon 23 -76 23 -76 0 3
rlabel polysilicon 37 -76 37 -76 0 3
rlabel polysilicon 44 -70 44 -70 0 1
rlabel polysilicon 44 -76 44 -76 0 3
rlabel polysilicon 58 -70 58 -70 0 1
rlabel polysilicon 61 -70 61 -70 0 2
rlabel polysilicon 65 -70 65 -70 0 1
rlabel polysilicon 65 -76 65 -76 0 3
rlabel polysilicon 72 -76 72 -76 0 3
rlabel polysilicon 82 -70 82 -70 0 2
rlabel polysilicon 86 -70 86 -70 0 1
rlabel polysilicon 93 -70 93 -70 0 1
rlabel polysilicon 93 -76 93 -76 0 3
rlabel polysilicon 100 -70 100 -70 0 1
rlabel polysilicon 100 -76 100 -76 0 3
rlabel polysilicon 110 -70 110 -70 0 2
rlabel polysilicon 114 -70 114 -70 0 1
rlabel polysilicon 121 -70 121 -70 0 1
rlabel polysilicon 121 -76 121 -76 0 3
rlabel polysilicon 128 -70 128 -70 0 1
rlabel polysilicon 128 -76 128 -76 0 3
rlabel polysilicon 135 -70 135 -70 0 1
rlabel polysilicon 135 -76 135 -76 0 3
rlabel polysilicon 142 -70 142 -70 0 1
rlabel polysilicon 142 -76 142 -76 0 3
rlabel polysilicon 152 -70 152 -70 0 2
rlabel polysilicon 149 -76 149 -76 0 3
rlabel polysilicon 152 -76 152 -76 0 4
rlabel polysilicon 156 -70 156 -70 0 1
rlabel polysilicon 156 -76 156 -76 0 3
rlabel polysilicon 163 -70 163 -70 0 1
rlabel polysilicon 163 -76 163 -76 0 3
rlabel polysilicon 170 -70 170 -70 0 1
rlabel polysilicon 170 -76 170 -76 0 3
rlabel polysilicon 177 -70 177 -70 0 1
rlabel polysilicon 180 -70 180 -70 0 2
rlabel polysilicon 184 -70 184 -70 0 1
rlabel polysilicon 184 -76 184 -76 0 3
rlabel polysilicon 187 -76 187 -76 0 4
rlabel polysilicon 194 -70 194 -70 0 2
rlabel polysilicon 194 -76 194 -76 0 4
rlabel polysilicon 198 -70 198 -70 0 1
rlabel polysilicon 198 -76 198 -76 0 3
rlabel polysilicon 205 -70 205 -70 0 1
rlabel polysilicon 205 -76 205 -76 0 3
rlabel polysilicon 208 -76 208 -76 0 4
rlabel polysilicon 212 -70 212 -70 0 1
rlabel polysilicon 212 -76 212 -76 0 3
rlabel polysilicon 222 -70 222 -70 0 2
rlabel polysilicon 222 -76 222 -76 0 4
rlabel polysilicon 226 -70 226 -70 0 1
rlabel polysilicon 226 -76 226 -76 0 3
rlabel polysilicon 233 -70 233 -70 0 1
rlabel polysilicon 233 -76 233 -76 0 3
rlabel polysilicon 240 -70 240 -70 0 1
rlabel polysilicon 240 -76 240 -76 0 3
rlabel polysilicon 247 -76 247 -76 0 3
rlabel polysilicon 250 -76 250 -76 0 4
rlabel polysilicon 254 -70 254 -70 0 1
rlabel polysilicon 254 -76 254 -76 0 3
rlabel polysilicon 261 -70 261 -70 0 1
rlabel polysilicon 261 -76 261 -76 0 3
rlabel polysilicon 268 -70 268 -70 0 1
rlabel polysilicon 271 -70 271 -70 0 2
rlabel polysilicon 275 -70 275 -70 0 1
rlabel polysilicon 275 -76 275 -76 0 3
rlabel polysilicon 282 -70 282 -70 0 1
rlabel polysilicon 289 -70 289 -70 0 1
rlabel polysilicon 289 -76 289 -76 0 3
rlabel polysilicon 299 -70 299 -70 0 2
rlabel polysilicon 299 -76 299 -76 0 4
rlabel polysilicon 303 -76 303 -76 0 3
rlabel polysilicon 306 -76 306 -76 0 4
rlabel polysilicon 310 -70 310 -70 0 1
rlabel polysilicon 310 -76 310 -76 0 3
rlabel polysilicon 317 -70 317 -70 0 1
rlabel polysilicon 317 -76 317 -76 0 3
rlabel polysilicon 324 -70 324 -70 0 1
rlabel polysilicon 324 -76 324 -76 0 3
rlabel polysilicon 331 -70 331 -70 0 1
rlabel polysilicon 331 -76 331 -76 0 3
rlabel polysilicon 341 -70 341 -70 0 2
rlabel polysilicon 345 -70 345 -70 0 1
rlabel polysilicon 345 -76 345 -76 0 3
rlabel polysilicon 359 -70 359 -70 0 1
rlabel polysilicon 359 -76 359 -76 0 3
rlabel polysilicon 366 -70 366 -70 0 1
rlabel polysilicon 366 -76 366 -76 0 3
rlabel polysilicon 373 -70 373 -70 0 1
rlabel polysilicon 373 -76 373 -76 0 3
rlabel polysilicon 380 -70 380 -70 0 1
rlabel polysilicon 380 -76 380 -76 0 3
rlabel polysilicon 387 -70 387 -70 0 1
rlabel polysilicon 387 -76 387 -76 0 3
rlabel polysilicon 394 -70 394 -70 0 1
rlabel polysilicon 397 -76 397 -76 0 4
rlabel polysilicon 401 -70 401 -70 0 1
rlabel polysilicon 401 -76 401 -76 0 3
rlabel polysilicon 408 -70 408 -70 0 1
rlabel polysilicon 408 -76 408 -76 0 3
rlabel polysilicon 415 -70 415 -70 0 1
rlabel polysilicon 415 -76 415 -76 0 3
rlabel polysilicon 422 -70 422 -70 0 1
rlabel polysilicon 422 -76 422 -76 0 3
rlabel polysilicon 436 -70 436 -70 0 1
rlabel polysilicon 436 -76 436 -76 0 3
rlabel polysilicon 44 -129 44 -129 0 3
rlabel polysilicon 51 -129 51 -129 0 3
rlabel polysilicon 58 -123 58 -123 0 1
rlabel polysilicon 58 -129 58 -129 0 3
rlabel polysilicon 65 -129 65 -129 0 3
rlabel polysilicon 75 -129 75 -129 0 4
rlabel polysilicon 79 -123 79 -123 0 1
rlabel polysilicon 79 -129 79 -129 0 3
rlabel polysilicon 86 -123 86 -123 0 1
rlabel polysilicon 86 -129 86 -129 0 3
rlabel polysilicon 93 -123 93 -123 0 1
rlabel polysilicon 93 -129 93 -129 0 3
rlabel polysilicon 100 -129 100 -129 0 3
rlabel polysilicon 103 -129 103 -129 0 4
rlabel polysilicon 107 -123 107 -123 0 1
rlabel polysilicon 107 -129 107 -129 0 3
rlabel polysilicon 114 -123 114 -123 0 1
rlabel polysilicon 121 -123 121 -123 0 1
rlabel polysilicon 121 -129 121 -129 0 3
rlabel polysilicon 128 -123 128 -123 0 1
rlabel polysilicon 128 -129 128 -129 0 3
rlabel polysilicon 135 -129 135 -129 0 3
rlabel polysilicon 138 -129 138 -129 0 4
rlabel polysilicon 142 -123 142 -123 0 1
rlabel polysilicon 142 -129 142 -129 0 3
rlabel polysilicon 149 -123 149 -123 0 1
rlabel polysilicon 149 -129 149 -129 0 3
rlabel polysilicon 156 -123 156 -123 0 1
rlabel polysilicon 159 -129 159 -129 0 4
rlabel polysilicon 163 -123 163 -123 0 1
rlabel polysilicon 163 -129 163 -129 0 3
rlabel polysilicon 173 -123 173 -123 0 2
rlabel polysilicon 170 -129 170 -129 0 3
rlabel polysilicon 177 -123 177 -123 0 1
rlabel polysilicon 177 -129 177 -129 0 3
rlabel polysilicon 180 -129 180 -129 0 4
rlabel polysilicon 187 -123 187 -123 0 2
rlabel polysilicon 187 -129 187 -129 0 4
rlabel polysilicon 191 -123 191 -123 0 1
rlabel polysilicon 191 -129 191 -129 0 3
rlabel polysilicon 198 -123 198 -123 0 1
rlabel polysilicon 198 -129 198 -129 0 3
rlabel polysilicon 205 -123 205 -123 0 1
rlabel polysilicon 205 -129 205 -129 0 3
rlabel polysilicon 212 -123 212 -123 0 1
rlabel polysilicon 212 -129 212 -129 0 3
rlabel polysilicon 219 -123 219 -123 0 1
rlabel polysilicon 219 -129 219 -129 0 3
rlabel polysilicon 226 -123 226 -123 0 1
rlabel polysilicon 226 -129 226 -129 0 3
rlabel polysilicon 233 -123 233 -123 0 1
rlabel polysilicon 233 -129 233 -129 0 3
rlabel polysilicon 240 -129 240 -129 0 3
rlabel polysilicon 243 -129 243 -129 0 4
rlabel polysilicon 247 -123 247 -123 0 1
rlabel polysilicon 247 -129 247 -129 0 3
rlabel polysilicon 254 -123 254 -123 0 1
rlabel polysilicon 261 -123 261 -123 0 1
rlabel polysilicon 261 -129 261 -129 0 3
rlabel polysilicon 268 -123 268 -123 0 1
rlabel polysilicon 268 -129 268 -129 0 3
rlabel polysilicon 275 -123 275 -123 0 1
rlabel polysilicon 275 -129 275 -129 0 3
rlabel polysilicon 282 -123 282 -123 0 1
rlabel polysilicon 285 -123 285 -123 0 2
rlabel polysilicon 282 -129 282 -129 0 3
rlabel polysilicon 289 -123 289 -123 0 1
rlabel polysilicon 292 -123 292 -123 0 2
rlabel polysilicon 289 -129 289 -129 0 3
rlabel polysilicon 296 -123 296 -123 0 1
rlabel polysilicon 296 -129 296 -129 0 3
rlabel polysilicon 303 -123 303 -123 0 1
rlabel polysilicon 303 -129 303 -129 0 3
rlabel polysilicon 310 -123 310 -123 0 1
rlabel polysilicon 310 -129 310 -129 0 3
rlabel polysilicon 317 -123 317 -123 0 1
rlabel polysilicon 317 -129 317 -129 0 3
rlabel polysilicon 324 -129 324 -129 0 3
rlabel polysilicon 327 -129 327 -129 0 4
rlabel polysilicon 331 -123 331 -123 0 1
rlabel polysilicon 334 -123 334 -123 0 2
rlabel polysilicon 334 -129 334 -129 0 4
rlabel polysilicon 338 -123 338 -123 0 1
rlabel polysilicon 345 -123 345 -123 0 1
rlabel polysilicon 345 -129 345 -129 0 3
rlabel polysilicon 352 -129 352 -129 0 3
rlabel polysilicon 359 -123 359 -123 0 1
rlabel polysilicon 359 -129 359 -129 0 3
rlabel polysilicon 366 -123 366 -123 0 1
rlabel polysilicon 366 -129 366 -129 0 3
rlabel polysilicon 373 -123 373 -123 0 1
rlabel polysilicon 373 -129 373 -129 0 3
rlabel polysilicon 380 -123 380 -123 0 1
rlabel polysilicon 383 -129 383 -129 0 4
rlabel polysilicon 387 -123 387 -123 0 1
rlabel polysilicon 387 -129 387 -129 0 3
rlabel polysilicon 394 -123 394 -123 0 1
rlabel polysilicon 394 -129 394 -129 0 3
rlabel polysilicon 401 -123 401 -123 0 1
rlabel polysilicon 401 -129 401 -129 0 3
rlabel polysilicon 408 -123 408 -123 0 1
rlabel polysilicon 408 -129 408 -129 0 3
rlabel polysilicon 415 -123 415 -123 0 1
rlabel polysilicon 415 -129 415 -129 0 3
rlabel polysilicon 422 -123 422 -123 0 1
rlabel polysilicon 422 -129 422 -129 0 3
rlabel polysilicon 429 -123 429 -123 0 1
rlabel polysilicon 429 -129 429 -129 0 3
rlabel polysilicon 436 -123 436 -123 0 1
rlabel polysilicon 436 -129 436 -129 0 3
rlabel polysilicon 443 -123 443 -123 0 1
rlabel polysilicon 443 -129 443 -129 0 3
rlabel polysilicon 450 -123 450 -123 0 1
rlabel polysilicon 450 -129 450 -129 0 3
rlabel polysilicon 457 -123 457 -123 0 1
rlabel polysilicon 457 -129 457 -129 0 3
rlabel polysilicon 464 -123 464 -123 0 1
rlabel polysilicon 464 -129 464 -129 0 3
rlabel polysilicon 471 -123 471 -123 0 1
rlabel polysilicon 471 -129 471 -129 0 3
rlabel polysilicon 478 -123 478 -123 0 1
rlabel polysilicon 478 -129 478 -129 0 3
rlabel polysilicon 485 -123 485 -123 0 1
rlabel polysilicon 485 -129 485 -129 0 3
rlabel polysilicon 492 -123 492 -123 0 1
rlabel polysilicon 492 -129 492 -129 0 3
rlabel polysilicon 499 -123 499 -123 0 1
rlabel polysilicon 499 -129 499 -129 0 3
rlabel polysilicon 506 -123 506 -123 0 1
rlabel polysilicon 506 -129 506 -129 0 3
rlabel polysilicon 513 -123 513 -123 0 1
rlabel polysilicon 513 -129 513 -129 0 3
rlabel polysilicon 520 -123 520 -123 0 1
rlabel polysilicon 520 -129 520 -129 0 3
rlabel polysilicon 12 -198 12 -198 0 2
rlabel polysilicon 16 -204 16 -204 0 3
rlabel polysilicon 23 -204 23 -204 0 3
rlabel polysilicon 30 -204 30 -204 0 3
rlabel polysilicon 33 -204 33 -204 0 4
rlabel polysilicon 44 -198 44 -198 0 1
rlabel polysilicon 44 -204 44 -204 0 3
rlabel polysilicon 58 -198 58 -198 0 1
rlabel polysilicon 58 -204 58 -204 0 3
rlabel polysilicon 65 -198 65 -198 0 1
rlabel polysilicon 65 -204 65 -204 0 3
rlabel polysilicon 72 -198 72 -198 0 1
rlabel polysilicon 72 -204 72 -204 0 3
rlabel polysilicon 79 -198 79 -198 0 1
rlabel polysilicon 79 -204 79 -204 0 3
rlabel polysilicon 89 -198 89 -198 0 2
rlabel polysilicon 89 -204 89 -204 0 4
rlabel polysilicon 93 -198 93 -198 0 1
rlabel polysilicon 93 -204 93 -204 0 3
rlabel polysilicon 100 -198 100 -198 0 1
rlabel polysilicon 100 -204 100 -204 0 3
rlabel polysilicon 107 -198 107 -198 0 1
rlabel polysilicon 107 -204 107 -204 0 3
rlabel polysilicon 117 -198 117 -198 0 2
rlabel polysilicon 114 -204 114 -204 0 3
rlabel polysilicon 121 -198 121 -198 0 1
rlabel polysilicon 121 -204 121 -204 0 3
rlabel polysilicon 128 -198 128 -198 0 1
rlabel polysilicon 128 -204 128 -204 0 3
rlabel polysilicon 135 -198 135 -198 0 1
rlabel polysilicon 135 -204 135 -204 0 3
rlabel polysilicon 142 -198 142 -198 0 1
rlabel polysilicon 142 -204 142 -204 0 3
rlabel polysilicon 149 -198 149 -198 0 1
rlabel polysilicon 152 -198 152 -198 0 2
rlabel polysilicon 152 -204 152 -204 0 4
rlabel polysilicon 156 -198 156 -198 0 1
rlabel polysilicon 156 -204 156 -204 0 3
rlabel polysilicon 163 -198 163 -198 0 1
rlabel polysilicon 163 -204 163 -204 0 3
rlabel polysilicon 170 -198 170 -198 0 1
rlabel polysilicon 170 -204 170 -204 0 3
rlabel polysilicon 177 -198 177 -198 0 1
rlabel polysilicon 180 -198 180 -198 0 2
rlabel polysilicon 180 -204 180 -204 0 4
rlabel polysilicon 187 -198 187 -198 0 2
rlabel polysilicon 187 -204 187 -204 0 4
rlabel polysilicon 191 -198 191 -198 0 1
rlabel polysilicon 191 -204 191 -204 0 3
rlabel polysilicon 198 -198 198 -198 0 1
rlabel polysilicon 198 -204 198 -204 0 3
rlabel polysilicon 201 -204 201 -204 0 4
rlabel polysilicon 208 -204 208 -204 0 4
rlabel polysilicon 212 -204 212 -204 0 3
rlabel polysilicon 215 -204 215 -204 0 4
rlabel polysilicon 219 -198 219 -198 0 1
rlabel polysilicon 219 -204 219 -204 0 3
rlabel polysilicon 226 -198 226 -198 0 1
rlabel polysilicon 226 -204 226 -204 0 3
rlabel polysilicon 233 -198 233 -198 0 1
rlabel polysilicon 233 -204 233 -204 0 3
rlabel polysilicon 240 -198 240 -198 0 1
rlabel polysilicon 240 -204 240 -204 0 3
rlabel polysilicon 250 -198 250 -198 0 2
rlabel polysilicon 247 -204 247 -204 0 3
rlabel polysilicon 250 -204 250 -204 0 4
rlabel polysilicon 254 -198 254 -198 0 1
rlabel polysilicon 254 -204 254 -204 0 3
rlabel polysilicon 257 -204 257 -204 0 4
rlabel polysilicon 261 -198 261 -198 0 1
rlabel polysilicon 261 -204 261 -204 0 3
rlabel polysilicon 271 -198 271 -198 0 2
rlabel polysilicon 268 -204 268 -204 0 3
rlabel polysilicon 275 -198 275 -198 0 1
rlabel polysilicon 275 -204 275 -204 0 3
rlabel polysilicon 282 -198 282 -198 0 1
rlabel polysilicon 285 -198 285 -198 0 2
rlabel polysilicon 282 -204 282 -204 0 3
rlabel polysilicon 285 -204 285 -204 0 4
rlabel polysilicon 289 -198 289 -198 0 1
rlabel polysilicon 292 -198 292 -198 0 2
rlabel polysilicon 292 -204 292 -204 0 4
rlabel polysilicon 296 -198 296 -198 0 1
rlabel polysilicon 296 -204 296 -204 0 3
rlabel polysilicon 303 -198 303 -198 0 1
rlabel polysilicon 303 -204 303 -204 0 3
rlabel polysilicon 313 -204 313 -204 0 4
rlabel polysilicon 317 -198 317 -198 0 1
rlabel polysilicon 317 -204 317 -204 0 3
rlabel polysilicon 324 -198 324 -198 0 1
rlabel polysilicon 324 -204 324 -204 0 3
rlabel polysilicon 331 -198 331 -198 0 1
rlabel polysilicon 331 -204 331 -204 0 3
rlabel polysilicon 341 -198 341 -198 0 2
rlabel polysilicon 338 -204 338 -204 0 3
rlabel polysilicon 345 -198 345 -198 0 1
rlabel polysilicon 345 -204 345 -204 0 3
rlabel polysilicon 352 -198 352 -198 0 1
rlabel polysilicon 352 -204 352 -204 0 3
rlabel polysilicon 359 -198 359 -198 0 1
rlabel polysilicon 359 -204 359 -204 0 3
rlabel polysilicon 366 -198 366 -198 0 1
rlabel polysilicon 366 -204 366 -204 0 3
rlabel polysilicon 373 -198 373 -198 0 1
rlabel polysilicon 373 -204 373 -204 0 3
rlabel polysilicon 380 -198 380 -198 0 1
rlabel polysilicon 380 -204 380 -204 0 3
rlabel polysilicon 387 -198 387 -198 0 1
rlabel polysilicon 390 -198 390 -198 0 2
rlabel polysilicon 387 -204 387 -204 0 3
rlabel polysilicon 394 -198 394 -198 0 1
rlabel polysilicon 394 -204 394 -204 0 3
rlabel polysilicon 401 -198 401 -198 0 1
rlabel polysilicon 401 -204 401 -204 0 3
rlabel polysilicon 408 -198 408 -198 0 1
rlabel polysilicon 411 -204 411 -204 0 4
rlabel polysilicon 415 -198 415 -198 0 1
rlabel polysilicon 415 -204 415 -204 0 3
rlabel polysilicon 422 -198 422 -198 0 1
rlabel polysilicon 425 -204 425 -204 0 4
rlabel polysilicon 429 -198 429 -198 0 1
rlabel polysilicon 429 -204 429 -204 0 3
rlabel polysilicon 436 -198 436 -198 0 1
rlabel polysilicon 436 -204 436 -204 0 3
rlabel polysilicon 443 -198 443 -198 0 1
rlabel polysilicon 443 -204 443 -204 0 3
rlabel polysilicon 450 -198 450 -198 0 1
rlabel polysilicon 450 -204 450 -204 0 3
rlabel polysilicon 457 -198 457 -198 0 1
rlabel polysilicon 457 -204 457 -204 0 3
rlabel polysilicon 464 -198 464 -198 0 1
rlabel polysilicon 464 -204 464 -204 0 3
rlabel polysilicon 471 -198 471 -198 0 1
rlabel polysilicon 471 -204 471 -204 0 3
rlabel polysilicon 478 -198 478 -198 0 1
rlabel polysilicon 478 -204 478 -204 0 3
rlabel polysilicon 485 -198 485 -198 0 1
rlabel polysilicon 485 -204 485 -204 0 3
rlabel polysilicon 492 -198 492 -198 0 1
rlabel polysilicon 492 -204 492 -204 0 3
rlabel polysilicon 499 -198 499 -198 0 1
rlabel polysilicon 499 -204 499 -204 0 3
rlabel polysilicon 506 -198 506 -198 0 1
rlabel polysilicon 506 -204 506 -204 0 3
rlabel polysilicon 513 -198 513 -198 0 1
rlabel polysilicon 513 -204 513 -204 0 3
rlabel polysilicon 520 -198 520 -198 0 1
rlabel polysilicon 520 -204 520 -204 0 3
rlabel polysilicon 527 -198 527 -198 0 1
rlabel polysilicon 527 -204 527 -204 0 3
rlabel polysilicon 534 -198 534 -198 0 1
rlabel polysilicon 534 -204 534 -204 0 3
rlabel polysilicon 541 -198 541 -198 0 1
rlabel polysilicon 541 -204 541 -204 0 3
rlabel polysilicon 548 -198 548 -198 0 1
rlabel polysilicon 548 -204 548 -204 0 3
rlabel polysilicon 555 -198 555 -198 0 1
rlabel polysilicon 555 -204 555 -204 0 3
rlabel polysilicon 562 -198 562 -198 0 1
rlabel polysilicon 562 -204 562 -204 0 3
rlabel polysilicon 569 -198 569 -198 0 1
rlabel polysilicon 569 -204 569 -204 0 3
rlabel polysilicon 576 -198 576 -198 0 1
rlabel polysilicon 576 -204 576 -204 0 3
rlabel polysilicon 583 -198 583 -198 0 1
rlabel polysilicon 583 -204 583 -204 0 3
rlabel polysilicon 590 -198 590 -198 0 1
rlabel polysilicon 590 -204 590 -204 0 3
rlabel polysilicon 597 -198 597 -198 0 1
rlabel polysilicon 597 -204 597 -204 0 3
rlabel polysilicon 604 -198 604 -198 0 1
rlabel polysilicon 604 -204 604 -204 0 3
rlabel polysilicon 611 -198 611 -198 0 1
rlabel polysilicon 611 -204 611 -204 0 3
rlabel polysilicon 618 -198 618 -198 0 1
rlabel polysilicon 618 -204 618 -204 0 3
rlabel polysilicon 625 -198 625 -198 0 1
rlabel polysilicon 625 -204 625 -204 0 3
rlabel polysilicon 632 -198 632 -198 0 1
rlabel polysilicon 632 -204 632 -204 0 3
rlabel polysilicon 639 -198 639 -198 0 1
rlabel polysilicon 639 -204 639 -204 0 3
rlabel polysilicon 646 -198 646 -198 0 1
rlabel polysilicon 646 -204 646 -204 0 3
rlabel polysilicon 653 -198 653 -198 0 1
rlabel polysilicon 653 -204 653 -204 0 3
rlabel polysilicon 660 -198 660 -198 0 1
rlabel polysilicon 660 -204 660 -204 0 3
rlabel polysilicon 16 -271 16 -271 0 1
rlabel polysilicon 30 -271 30 -271 0 1
rlabel polysilicon 30 -277 30 -277 0 3
rlabel polysilicon 44 -277 44 -277 0 3
rlabel polysilicon 51 -271 51 -271 0 1
rlabel polysilicon 51 -277 51 -277 0 3
rlabel polysilicon 58 -271 58 -271 0 1
rlabel polysilicon 58 -277 58 -277 0 3
rlabel polysilicon 65 -271 65 -271 0 1
rlabel polysilicon 65 -277 65 -277 0 3
rlabel polysilicon 72 -271 72 -271 0 1
rlabel polysilicon 72 -277 72 -277 0 3
rlabel polysilicon 82 -271 82 -271 0 2
rlabel polysilicon 79 -277 79 -277 0 3
rlabel polysilicon 89 -271 89 -271 0 2
rlabel polysilicon 89 -277 89 -277 0 4
rlabel polysilicon 93 -271 93 -271 0 1
rlabel polysilicon 93 -277 93 -277 0 3
rlabel polysilicon 100 -271 100 -271 0 1
rlabel polysilicon 103 -271 103 -271 0 2
rlabel polysilicon 100 -277 100 -277 0 3
rlabel polysilicon 107 -271 107 -271 0 1
rlabel polysilicon 107 -277 107 -277 0 3
rlabel polysilicon 114 -271 114 -271 0 1
rlabel polysilicon 114 -277 114 -277 0 3
rlabel polysilicon 121 -271 121 -271 0 1
rlabel polysilicon 124 -271 124 -271 0 2
rlabel polysilicon 121 -277 121 -277 0 3
rlabel polysilicon 128 -271 128 -271 0 1
rlabel polysilicon 128 -277 128 -277 0 3
rlabel polysilicon 135 -271 135 -271 0 1
rlabel polysilicon 135 -277 135 -277 0 3
rlabel polysilicon 142 -271 142 -271 0 1
rlabel polysilicon 142 -277 142 -277 0 3
rlabel polysilicon 149 -271 149 -271 0 1
rlabel polysilicon 149 -277 149 -277 0 3
rlabel polysilicon 156 -271 156 -271 0 1
rlabel polysilicon 159 -277 159 -277 0 4
rlabel polysilicon 163 -271 163 -271 0 1
rlabel polysilicon 163 -277 163 -277 0 3
rlabel polysilicon 170 -271 170 -271 0 1
rlabel polysilicon 170 -277 170 -277 0 3
rlabel polysilicon 177 -271 177 -271 0 1
rlabel polysilicon 180 -271 180 -271 0 2
rlabel polysilicon 177 -277 177 -277 0 3
rlabel polysilicon 184 -271 184 -271 0 1
rlabel polysilicon 184 -277 184 -277 0 3
rlabel polysilicon 191 -271 191 -271 0 1
rlabel polysilicon 191 -277 191 -277 0 3
rlabel polysilicon 198 -271 198 -271 0 1
rlabel polysilicon 198 -277 198 -277 0 3
rlabel polysilicon 205 -271 205 -271 0 1
rlabel polysilicon 205 -277 205 -277 0 3
rlabel polysilicon 212 -271 212 -271 0 1
rlabel polysilicon 212 -277 212 -277 0 3
rlabel polysilicon 219 -271 219 -271 0 1
rlabel polysilicon 219 -277 219 -277 0 3
rlabel polysilicon 226 -271 226 -271 0 1
rlabel polysilicon 226 -277 226 -277 0 3
rlabel polysilicon 233 -271 233 -271 0 1
rlabel polysilicon 233 -277 233 -277 0 3
rlabel polysilicon 240 -271 240 -271 0 1
rlabel polysilicon 243 -271 243 -271 0 2
rlabel polysilicon 250 -277 250 -277 0 4
rlabel polysilicon 257 -271 257 -271 0 2
rlabel polysilicon 254 -277 254 -277 0 3
rlabel polysilicon 261 -271 261 -271 0 1
rlabel polysilicon 261 -277 261 -277 0 3
rlabel polysilicon 268 -271 268 -271 0 1
rlabel polysilicon 268 -277 268 -277 0 3
rlabel polysilicon 278 -271 278 -271 0 2
rlabel polysilicon 282 -271 282 -271 0 1
rlabel polysilicon 285 -271 285 -271 0 2
rlabel polysilicon 282 -277 282 -277 0 3
rlabel polysilicon 285 -277 285 -277 0 4
rlabel polysilicon 289 -271 289 -271 0 1
rlabel polysilicon 289 -277 289 -277 0 3
rlabel polysilicon 299 -271 299 -271 0 2
rlabel polysilicon 296 -277 296 -277 0 3
rlabel polysilicon 299 -277 299 -277 0 4
rlabel polysilicon 303 -271 303 -271 0 1
rlabel polysilicon 306 -271 306 -271 0 2
rlabel polysilicon 303 -277 303 -277 0 3
rlabel polysilicon 306 -277 306 -277 0 4
rlabel polysilicon 310 -271 310 -271 0 1
rlabel polysilicon 310 -277 310 -277 0 3
rlabel polysilicon 320 -271 320 -271 0 2
rlabel polysilicon 317 -277 317 -277 0 3
rlabel polysilicon 320 -277 320 -277 0 4
rlabel polysilicon 324 -271 324 -271 0 1
rlabel polysilicon 324 -277 324 -277 0 3
rlabel polysilicon 331 -271 331 -271 0 1
rlabel polysilicon 334 -271 334 -271 0 2
rlabel polysilicon 334 -277 334 -277 0 4
rlabel polysilicon 338 -271 338 -271 0 1
rlabel polysilicon 338 -277 338 -277 0 3
rlabel polysilicon 345 -271 345 -271 0 1
rlabel polysilicon 345 -277 345 -277 0 3
rlabel polysilicon 352 -277 352 -277 0 3
rlabel polysilicon 355 -277 355 -277 0 4
rlabel polysilicon 359 -271 359 -271 0 1
rlabel polysilicon 359 -277 359 -277 0 3
rlabel polysilicon 366 -271 366 -271 0 1
rlabel polysilicon 369 -277 369 -277 0 4
rlabel polysilicon 373 -271 373 -271 0 1
rlabel polysilicon 373 -277 373 -277 0 3
rlabel polysilicon 380 -271 380 -271 0 1
rlabel polysilicon 380 -277 380 -277 0 3
rlabel polysilicon 387 -271 387 -271 0 1
rlabel polysilicon 387 -277 387 -277 0 3
rlabel polysilicon 394 -271 394 -271 0 1
rlabel polysilicon 394 -277 394 -277 0 3
rlabel polysilicon 401 -271 401 -271 0 1
rlabel polysilicon 401 -277 401 -277 0 3
rlabel polysilicon 408 -271 408 -271 0 1
rlabel polysilicon 408 -277 408 -277 0 3
rlabel polysilicon 415 -271 415 -271 0 1
rlabel polysilicon 415 -277 415 -277 0 3
rlabel polysilicon 422 -271 422 -271 0 1
rlabel polysilicon 422 -277 422 -277 0 3
rlabel polysilicon 429 -271 429 -271 0 1
rlabel polysilicon 429 -277 429 -277 0 3
rlabel polysilicon 436 -271 436 -271 0 1
rlabel polysilicon 436 -277 436 -277 0 3
rlabel polysilicon 443 -271 443 -271 0 1
rlabel polysilicon 443 -277 443 -277 0 3
rlabel polysilicon 450 -271 450 -271 0 1
rlabel polysilicon 450 -277 450 -277 0 3
rlabel polysilicon 457 -271 457 -271 0 1
rlabel polysilicon 457 -277 457 -277 0 3
rlabel polysilicon 464 -271 464 -271 0 1
rlabel polysilicon 464 -277 464 -277 0 3
rlabel polysilicon 471 -271 471 -271 0 1
rlabel polysilicon 471 -277 471 -277 0 3
rlabel polysilicon 478 -271 478 -271 0 1
rlabel polysilicon 478 -277 478 -277 0 3
rlabel polysilicon 485 -271 485 -271 0 1
rlabel polysilicon 485 -277 485 -277 0 3
rlabel polysilicon 492 -271 492 -271 0 1
rlabel polysilicon 492 -277 492 -277 0 3
rlabel polysilicon 499 -271 499 -271 0 1
rlabel polysilicon 499 -277 499 -277 0 3
rlabel polysilicon 506 -271 506 -271 0 1
rlabel polysilicon 506 -277 506 -277 0 3
rlabel polysilicon 513 -271 513 -271 0 1
rlabel polysilicon 513 -277 513 -277 0 3
rlabel polysilicon 520 -271 520 -271 0 1
rlabel polysilicon 520 -277 520 -277 0 3
rlabel polysilicon 527 -271 527 -271 0 1
rlabel polysilicon 527 -277 527 -277 0 3
rlabel polysilicon 534 -271 534 -271 0 1
rlabel polysilicon 534 -277 534 -277 0 3
rlabel polysilicon 541 -271 541 -271 0 1
rlabel polysilicon 541 -277 541 -277 0 3
rlabel polysilicon 548 -271 548 -271 0 1
rlabel polysilicon 548 -277 548 -277 0 3
rlabel polysilicon 562 -271 562 -271 0 1
rlabel polysilicon 562 -277 562 -277 0 3
rlabel polysilicon 569 -271 569 -271 0 1
rlabel polysilicon 569 -277 569 -277 0 3
rlabel polysilicon 576 -271 576 -271 0 1
rlabel polysilicon 576 -277 576 -277 0 3
rlabel polysilicon 583 -271 583 -271 0 1
rlabel polysilicon 583 -277 583 -277 0 3
rlabel polysilicon 590 -271 590 -271 0 1
rlabel polysilicon 590 -277 590 -277 0 3
rlabel polysilicon 597 -271 597 -271 0 1
rlabel polysilicon 597 -277 597 -277 0 3
rlabel polysilicon 604 -271 604 -271 0 1
rlabel polysilicon 604 -277 604 -277 0 3
rlabel polysilicon 611 -271 611 -271 0 1
rlabel polysilicon 611 -277 611 -277 0 3
rlabel polysilicon 618 -271 618 -271 0 1
rlabel polysilicon 625 -271 625 -271 0 1
rlabel polysilicon 625 -277 625 -277 0 3
rlabel polysilicon 632 -271 632 -271 0 1
rlabel polysilicon 632 -277 632 -277 0 3
rlabel polysilicon 639 -277 639 -277 0 3
rlabel polysilicon 667 -271 667 -271 0 1
rlabel polysilicon 667 -277 667 -277 0 3
rlabel polysilicon 9 -342 9 -342 0 3
rlabel polysilicon 12 -342 12 -342 0 4
rlabel polysilicon 16 -336 16 -336 0 1
rlabel polysilicon 23 -336 23 -336 0 1
rlabel polysilicon 30 -336 30 -336 0 1
rlabel polysilicon 37 -336 37 -336 0 1
rlabel polysilicon 37 -342 37 -342 0 3
rlabel polysilicon 47 -336 47 -336 0 2
rlabel polysilicon 44 -342 44 -342 0 3
rlabel polysilicon 51 -336 51 -336 0 1
rlabel polysilicon 54 -336 54 -336 0 2
rlabel polysilicon 58 -336 58 -336 0 1
rlabel polysilicon 58 -342 58 -342 0 3
rlabel polysilicon 65 -336 65 -336 0 1
rlabel polysilicon 68 -342 68 -342 0 4
rlabel polysilicon 72 -336 72 -336 0 1
rlabel polysilicon 75 -342 75 -342 0 4
rlabel polysilicon 79 -336 79 -336 0 1
rlabel polysilicon 82 -336 82 -336 0 2
rlabel polysilicon 79 -342 79 -342 0 3
rlabel polysilicon 89 -336 89 -336 0 2
rlabel polysilicon 86 -342 86 -342 0 3
rlabel polysilicon 89 -342 89 -342 0 4
rlabel polysilicon 93 -336 93 -336 0 1
rlabel polysilicon 93 -342 93 -342 0 3
rlabel polysilicon 100 -342 100 -342 0 3
rlabel polysilicon 107 -336 107 -336 0 1
rlabel polysilicon 107 -342 107 -342 0 3
rlabel polysilicon 114 -336 114 -336 0 1
rlabel polysilicon 114 -342 114 -342 0 3
rlabel polysilicon 121 -336 121 -336 0 1
rlabel polysilicon 121 -342 121 -342 0 3
rlabel polysilicon 128 -336 128 -336 0 1
rlabel polysilicon 128 -342 128 -342 0 3
rlabel polysilicon 135 -336 135 -336 0 1
rlabel polysilicon 135 -342 135 -342 0 3
rlabel polysilicon 142 -336 142 -336 0 1
rlabel polysilicon 145 -336 145 -336 0 2
rlabel polysilicon 142 -342 142 -342 0 3
rlabel polysilicon 149 -336 149 -336 0 1
rlabel polysilicon 149 -342 149 -342 0 3
rlabel polysilicon 159 -336 159 -336 0 2
rlabel polysilicon 156 -342 156 -342 0 3
rlabel polysilicon 163 -342 163 -342 0 3
rlabel polysilicon 170 -336 170 -336 0 1
rlabel polysilicon 170 -342 170 -342 0 3
rlabel polysilicon 177 -336 177 -336 0 1
rlabel polysilicon 177 -342 177 -342 0 3
rlabel polysilicon 184 -336 184 -336 0 1
rlabel polysilicon 187 -336 187 -336 0 2
rlabel polysilicon 191 -336 191 -336 0 1
rlabel polysilicon 191 -342 191 -342 0 3
rlabel polysilicon 201 -336 201 -336 0 2
rlabel polysilicon 201 -342 201 -342 0 4
rlabel polysilicon 205 -336 205 -336 0 1
rlabel polysilicon 205 -342 205 -342 0 3
rlabel polysilicon 212 -336 212 -336 0 1
rlabel polysilicon 212 -342 212 -342 0 3
rlabel polysilicon 219 -336 219 -336 0 1
rlabel polysilicon 219 -342 219 -342 0 3
rlabel polysilicon 226 -336 226 -336 0 1
rlabel polysilicon 226 -342 226 -342 0 3
rlabel polysilicon 233 -336 233 -336 0 1
rlabel polysilicon 233 -342 233 -342 0 3
rlabel polysilicon 240 -336 240 -336 0 1
rlabel polysilicon 247 -336 247 -336 0 1
rlabel polysilicon 247 -342 247 -342 0 3
rlabel polysilicon 254 -336 254 -336 0 1
rlabel polysilicon 254 -342 254 -342 0 3
rlabel polysilicon 261 -336 261 -336 0 1
rlabel polysilicon 261 -342 261 -342 0 3
rlabel polysilicon 268 -336 268 -336 0 1
rlabel polysilicon 268 -342 268 -342 0 3
rlabel polysilicon 275 -336 275 -336 0 1
rlabel polysilicon 275 -342 275 -342 0 3
rlabel polysilicon 282 -336 282 -336 0 1
rlabel polysilicon 282 -342 282 -342 0 3
rlabel polysilicon 289 -336 289 -336 0 1
rlabel polysilicon 289 -342 289 -342 0 3
rlabel polysilicon 296 -336 296 -336 0 1
rlabel polysilicon 296 -342 296 -342 0 3
rlabel polysilicon 303 -336 303 -336 0 1
rlabel polysilicon 303 -342 303 -342 0 3
rlabel polysilicon 313 -336 313 -336 0 2
rlabel polysilicon 310 -342 310 -342 0 3
rlabel polysilicon 313 -342 313 -342 0 4
rlabel polysilicon 317 -336 317 -336 0 1
rlabel polysilicon 320 -336 320 -336 0 2
rlabel polysilicon 324 -336 324 -336 0 1
rlabel polysilicon 324 -342 324 -342 0 3
rlabel polysilicon 327 -342 327 -342 0 4
rlabel polysilicon 331 -336 331 -336 0 1
rlabel polysilicon 331 -342 331 -342 0 3
rlabel polysilicon 341 -336 341 -336 0 2
rlabel polysilicon 341 -342 341 -342 0 4
rlabel polysilicon 345 -336 345 -336 0 1
rlabel polysilicon 345 -342 345 -342 0 3
rlabel polysilicon 352 -342 352 -342 0 3
rlabel polysilicon 355 -342 355 -342 0 4
rlabel polysilicon 362 -336 362 -336 0 2
rlabel polysilicon 359 -342 359 -342 0 3
rlabel polysilicon 362 -342 362 -342 0 4
rlabel polysilicon 366 -336 366 -336 0 1
rlabel polysilicon 366 -342 366 -342 0 3
rlabel polysilicon 373 -336 373 -336 0 1
rlabel polysilicon 373 -342 373 -342 0 3
rlabel polysilicon 380 -336 380 -336 0 1
rlabel polysilicon 380 -342 380 -342 0 3
rlabel polysilicon 387 -336 387 -336 0 1
rlabel polysilicon 390 -336 390 -336 0 2
rlabel polysilicon 390 -342 390 -342 0 4
rlabel polysilicon 394 -336 394 -336 0 1
rlabel polysilicon 394 -342 394 -342 0 3
rlabel polysilicon 401 -336 401 -336 0 1
rlabel polysilicon 401 -342 401 -342 0 3
rlabel polysilicon 408 -336 408 -336 0 1
rlabel polysilicon 408 -342 408 -342 0 3
rlabel polysilicon 415 -336 415 -336 0 1
rlabel polysilicon 415 -342 415 -342 0 3
rlabel polysilicon 422 -336 422 -336 0 1
rlabel polysilicon 422 -342 422 -342 0 3
rlabel polysilicon 429 -336 429 -336 0 1
rlabel polysilicon 429 -342 429 -342 0 3
rlabel polysilicon 436 -336 436 -336 0 1
rlabel polysilicon 436 -342 436 -342 0 3
rlabel polysilicon 443 -336 443 -336 0 1
rlabel polysilicon 443 -342 443 -342 0 3
rlabel polysilicon 450 -336 450 -336 0 1
rlabel polysilicon 450 -342 450 -342 0 3
rlabel polysilicon 457 -336 457 -336 0 1
rlabel polysilicon 457 -342 457 -342 0 3
rlabel polysilicon 464 -336 464 -336 0 1
rlabel polysilicon 464 -342 464 -342 0 3
rlabel polysilicon 471 -336 471 -336 0 1
rlabel polysilicon 471 -342 471 -342 0 3
rlabel polysilicon 478 -336 478 -336 0 1
rlabel polysilicon 478 -342 478 -342 0 3
rlabel polysilicon 485 -336 485 -336 0 1
rlabel polysilicon 485 -342 485 -342 0 3
rlabel polysilicon 492 -342 492 -342 0 3
rlabel polysilicon 495 -342 495 -342 0 4
rlabel polysilicon 499 -336 499 -336 0 1
rlabel polysilicon 499 -342 499 -342 0 3
rlabel polysilicon 506 -336 506 -336 0 1
rlabel polysilicon 506 -342 506 -342 0 3
rlabel polysilicon 513 -336 513 -336 0 1
rlabel polysilicon 513 -342 513 -342 0 3
rlabel polysilicon 520 -336 520 -336 0 1
rlabel polysilicon 520 -342 520 -342 0 3
rlabel polysilicon 527 -336 527 -336 0 1
rlabel polysilicon 527 -342 527 -342 0 3
rlabel polysilicon 534 -336 534 -336 0 1
rlabel polysilicon 534 -342 534 -342 0 3
rlabel polysilicon 541 -336 541 -336 0 1
rlabel polysilicon 541 -342 541 -342 0 3
rlabel polysilicon 548 -336 548 -336 0 1
rlabel polysilicon 548 -342 548 -342 0 3
rlabel polysilicon 555 -336 555 -336 0 1
rlabel polysilicon 555 -342 555 -342 0 3
rlabel polysilicon 562 -336 562 -336 0 1
rlabel polysilicon 562 -342 562 -342 0 3
rlabel polysilicon 569 -336 569 -336 0 1
rlabel polysilicon 569 -342 569 -342 0 3
rlabel polysilicon 576 -336 576 -336 0 1
rlabel polysilicon 576 -342 576 -342 0 3
rlabel polysilicon 583 -336 583 -336 0 1
rlabel polysilicon 583 -342 583 -342 0 3
rlabel polysilicon 590 -336 590 -336 0 1
rlabel polysilicon 590 -342 590 -342 0 3
rlabel polysilicon 604 -336 604 -336 0 1
rlabel polysilicon 604 -342 604 -342 0 3
rlabel polysilicon 611 -336 611 -336 0 1
rlabel polysilicon 611 -342 611 -342 0 3
rlabel polysilicon 618 -336 618 -336 0 1
rlabel polysilicon 618 -342 618 -342 0 3
rlabel polysilicon 625 -336 625 -336 0 1
rlabel polysilicon 625 -342 625 -342 0 3
rlabel polysilicon 632 -336 632 -336 0 1
rlabel polysilicon 632 -342 632 -342 0 3
rlabel polysilicon 639 -336 639 -336 0 1
rlabel polysilicon 639 -342 639 -342 0 3
rlabel polysilicon 646 -336 646 -336 0 1
rlabel polysilicon 646 -342 646 -342 0 3
rlabel polysilicon 653 -336 653 -336 0 1
rlabel polysilicon 653 -342 653 -342 0 3
rlabel polysilicon 660 -336 660 -336 0 1
rlabel polysilicon 660 -342 660 -342 0 3
rlabel polysilicon 667 -336 667 -336 0 1
rlabel polysilicon 667 -342 667 -342 0 3
rlabel polysilicon 674 -336 674 -336 0 1
rlabel polysilicon 674 -342 674 -342 0 3
rlabel polysilicon 709 -336 709 -336 0 1
rlabel polysilicon 709 -342 709 -342 0 3
rlabel polysilicon 23 -403 23 -403 0 1
rlabel polysilicon 23 -409 23 -409 0 3
rlabel polysilicon 30 -403 30 -403 0 1
rlabel polysilicon 37 -403 37 -403 0 1
rlabel polysilicon 37 -409 37 -409 0 3
rlabel polysilicon 44 -403 44 -403 0 1
rlabel polysilicon 44 -409 44 -409 0 3
rlabel polysilicon 51 -403 51 -403 0 1
rlabel polysilicon 51 -409 51 -409 0 3
rlabel polysilicon 58 -403 58 -403 0 1
rlabel polysilicon 58 -409 58 -409 0 3
rlabel polysilicon 65 -403 65 -403 0 1
rlabel polysilicon 68 -409 68 -409 0 4
rlabel polysilicon 72 -403 72 -403 0 1
rlabel polysilicon 72 -409 72 -409 0 3
rlabel polysilicon 79 -403 79 -403 0 1
rlabel polysilicon 79 -409 79 -409 0 3
rlabel polysilicon 86 -403 86 -403 0 1
rlabel polysilicon 86 -409 86 -409 0 3
rlabel polysilicon 93 -403 93 -403 0 1
rlabel polysilicon 93 -409 93 -409 0 3
rlabel polysilicon 96 -409 96 -409 0 4
rlabel polysilicon 100 -403 100 -403 0 1
rlabel polysilicon 100 -409 100 -409 0 3
rlabel polysilicon 110 -403 110 -403 0 2
rlabel polysilicon 110 -409 110 -409 0 4
rlabel polysilicon 117 -403 117 -403 0 2
rlabel polysilicon 121 -403 121 -403 0 1
rlabel polysilicon 121 -409 121 -409 0 3
rlabel polysilicon 124 -409 124 -409 0 4
rlabel polysilicon 128 -403 128 -403 0 1
rlabel polysilicon 128 -409 128 -409 0 3
rlabel polysilicon 135 -403 135 -403 0 1
rlabel polysilicon 135 -409 135 -409 0 3
rlabel polysilicon 142 -403 142 -403 0 1
rlabel polysilicon 142 -409 142 -409 0 3
rlabel polysilicon 149 -403 149 -403 0 1
rlabel polysilicon 149 -409 149 -409 0 3
rlabel polysilicon 156 -403 156 -403 0 1
rlabel polysilicon 163 -403 163 -403 0 1
rlabel polysilicon 163 -409 163 -409 0 3
rlabel polysilicon 170 -403 170 -403 0 1
rlabel polysilicon 170 -409 170 -409 0 3
rlabel polysilicon 177 -403 177 -403 0 1
rlabel polysilicon 177 -409 177 -409 0 3
rlabel polysilicon 187 -403 187 -403 0 2
rlabel polysilicon 184 -409 184 -409 0 3
rlabel polysilicon 191 -403 191 -403 0 1
rlabel polysilicon 191 -409 191 -409 0 3
rlabel polysilicon 198 -403 198 -403 0 1
rlabel polysilicon 198 -409 198 -409 0 3
rlabel polysilicon 205 -403 205 -403 0 1
rlabel polysilicon 205 -409 205 -409 0 3
rlabel polysilicon 212 -403 212 -403 0 1
rlabel polysilicon 212 -409 212 -409 0 3
rlabel polysilicon 219 -403 219 -403 0 1
rlabel polysilicon 219 -409 219 -409 0 3
rlabel polysilicon 226 -403 226 -403 0 1
rlabel polysilicon 229 -409 229 -409 0 4
rlabel polysilicon 233 -403 233 -403 0 1
rlabel polysilicon 233 -409 233 -409 0 3
rlabel polysilicon 243 -403 243 -403 0 2
rlabel polysilicon 240 -409 240 -409 0 3
rlabel polysilicon 243 -409 243 -409 0 4
rlabel polysilicon 247 -403 247 -403 0 1
rlabel polysilicon 247 -409 247 -409 0 3
rlabel polysilicon 254 -403 254 -403 0 1
rlabel polysilicon 254 -409 254 -409 0 3
rlabel polysilicon 261 -403 261 -403 0 1
rlabel polysilicon 261 -409 261 -409 0 3
rlabel polysilicon 268 -403 268 -403 0 1
rlabel polysilicon 268 -409 268 -409 0 3
rlabel polysilicon 275 -403 275 -403 0 1
rlabel polysilicon 275 -409 275 -409 0 3
rlabel polysilicon 282 -403 282 -403 0 1
rlabel polysilicon 282 -409 282 -409 0 3
rlabel polysilicon 285 -409 285 -409 0 4
rlabel polysilicon 289 -403 289 -403 0 1
rlabel polysilicon 289 -409 289 -409 0 3
rlabel polysilicon 296 -403 296 -403 0 1
rlabel polysilicon 296 -409 296 -409 0 3
rlabel polysilicon 303 -403 303 -403 0 1
rlabel polysilicon 303 -409 303 -409 0 3
rlabel polysilicon 310 -403 310 -403 0 1
rlabel polysilicon 310 -409 310 -409 0 3
rlabel polysilicon 317 -403 317 -403 0 1
rlabel polysilicon 317 -409 317 -409 0 3
rlabel polysilicon 324 -403 324 -403 0 1
rlabel polysilicon 327 -409 327 -409 0 4
rlabel polysilicon 334 -403 334 -403 0 2
rlabel polysilicon 338 -403 338 -403 0 1
rlabel polysilicon 341 -409 341 -409 0 4
rlabel polysilicon 345 -403 345 -403 0 1
rlabel polysilicon 345 -409 345 -409 0 3
rlabel polysilicon 355 -403 355 -403 0 2
rlabel polysilicon 352 -409 352 -409 0 3
rlabel polysilicon 359 -403 359 -403 0 1
rlabel polysilicon 359 -409 359 -409 0 3
rlabel polysilicon 366 -403 366 -403 0 1
rlabel polysilicon 366 -409 366 -409 0 3
rlabel polysilicon 373 -403 373 -403 0 1
rlabel polysilicon 373 -409 373 -409 0 3
rlabel polysilicon 380 -403 380 -403 0 1
rlabel polysilicon 383 -403 383 -403 0 2
rlabel polysilicon 380 -409 380 -409 0 3
rlabel polysilicon 383 -409 383 -409 0 4
rlabel polysilicon 387 -403 387 -403 0 1
rlabel polysilicon 390 -403 390 -403 0 2
rlabel polysilicon 387 -409 387 -409 0 3
rlabel polysilicon 390 -409 390 -409 0 4
rlabel polysilicon 394 -403 394 -403 0 1
rlabel polysilicon 394 -409 394 -409 0 3
rlabel polysilicon 401 -403 401 -403 0 1
rlabel polysilicon 401 -409 401 -409 0 3
rlabel polysilicon 411 -403 411 -403 0 2
rlabel polysilicon 415 -403 415 -403 0 1
rlabel polysilicon 415 -409 415 -409 0 3
rlabel polysilicon 422 -403 422 -403 0 1
rlabel polysilicon 422 -409 422 -409 0 3
rlabel polysilicon 432 -409 432 -409 0 4
rlabel polysilicon 436 -403 436 -403 0 1
rlabel polysilicon 436 -409 436 -409 0 3
rlabel polysilicon 443 -403 443 -403 0 1
rlabel polysilicon 443 -409 443 -409 0 3
rlabel polysilicon 450 -403 450 -403 0 1
rlabel polysilicon 450 -409 450 -409 0 3
rlabel polysilicon 457 -403 457 -403 0 1
rlabel polysilicon 457 -409 457 -409 0 3
rlabel polysilicon 467 -403 467 -403 0 2
rlabel polysilicon 464 -409 464 -409 0 3
rlabel polysilicon 471 -403 471 -403 0 1
rlabel polysilicon 471 -409 471 -409 0 3
rlabel polysilicon 481 -403 481 -403 0 2
rlabel polysilicon 478 -409 478 -409 0 3
rlabel polysilicon 481 -409 481 -409 0 4
rlabel polysilicon 485 -403 485 -403 0 1
rlabel polysilicon 485 -409 485 -409 0 3
rlabel polysilicon 492 -403 492 -403 0 1
rlabel polysilicon 492 -409 492 -409 0 3
rlabel polysilicon 502 -409 502 -409 0 4
rlabel polysilicon 506 -403 506 -403 0 1
rlabel polysilicon 506 -409 506 -409 0 3
rlabel polysilicon 513 -403 513 -403 0 1
rlabel polysilicon 513 -409 513 -409 0 3
rlabel polysilicon 520 -403 520 -403 0 1
rlabel polysilicon 520 -409 520 -409 0 3
rlabel polysilicon 527 -403 527 -403 0 1
rlabel polysilicon 527 -409 527 -409 0 3
rlabel polysilicon 534 -403 534 -403 0 1
rlabel polysilicon 534 -409 534 -409 0 3
rlabel polysilicon 541 -403 541 -403 0 1
rlabel polysilicon 541 -409 541 -409 0 3
rlabel polysilicon 548 -403 548 -403 0 1
rlabel polysilicon 548 -409 548 -409 0 3
rlabel polysilicon 555 -403 555 -403 0 1
rlabel polysilicon 555 -409 555 -409 0 3
rlabel polysilicon 562 -403 562 -403 0 1
rlabel polysilicon 562 -409 562 -409 0 3
rlabel polysilicon 569 -403 569 -403 0 1
rlabel polysilicon 569 -409 569 -409 0 3
rlabel polysilicon 576 -403 576 -403 0 1
rlabel polysilicon 576 -409 576 -409 0 3
rlabel polysilicon 583 -403 583 -403 0 1
rlabel polysilicon 583 -409 583 -409 0 3
rlabel polysilicon 590 -403 590 -403 0 1
rlabel polysilicon 590 -409 590 -409 0 3
rlabel polysilicon 597 -403 597 -403 0 1
rlabel polysilicon 597 -409 597 -409 0 3
rlabel polysilicon 604 -403 604 -403 0 1
rlabel polysilicon 604 -409 604 -409 0 3
rlabel polysilicon 611 -403 611 -403 0 1
rlabel polysilicon 611 -409 611 -409 0 3
rlabel polysilicon 618 -403 618 -403 0 1
rlabel polysilicon 618 -409 618 -409 0 3
rlabel polysilicon 625 -403 625 -403 0 1
rlabel polysilicon 625 -409 625 -409 0 3
rlabel polysilicon 635 -403 635 -403 0 2
rlabel polysilicon 639 -403 639 -403 0 1
rlabel polysilicon 639 -409 639 -409 0 3
rlabel polysilicon 646 -403 646 -403 0 1
rlabel polysilicon 646 -409 646 -409 0 3
rlabel polysilicon 653 -403 653 -403 0 1
rlabel polysilicon 656 -409 656 -409 0 4
rlabel polysilicon 660 -403 660 -403 0 1
rlabel polysilicon 660 -409 660 -409 0 3
rlabel polysilicon 667 -403 667 -403 0 1
rlabel polysilicon 667 -409 667 -409 0 3
rlabel polysilicon 716 -403 716 -403 0 1
rlabel polysilicon 716 -409 716 -409 0 3
rlabel polysilicon 9 -468 9 -468 0 1
rlabel polysilicon 9 -474 9 -474 0 3
rlabel polysilicon 16 -468 16 -468 0 1
rlabel polysilicon 16 -474 16 -474 0 3
rlabel polysilicon 26 -474 26 -474 0 4
rlabel polysilicon 30 -468 30 -468 0 1
rlabel polysilicon 30 -474 30 -474 0 3
rlabel polysilicon 37 -468 37 -468 0 1
rlabel polysilicon 37 -474 37 -474 0 3
rlabel polysilicon 44 -468 44 -468 0 1
rlabel polysilicon 44 -474 44 -474 0 3
rlabel polysilicon 51 -468 51 -468 0 1
rlabel polysilicon 51 -474 51 -474 0 3
rlabel polysilicon 58 -468 58 -468 0 1
rlabel polysilicon 58 -474 58 -474 0 3
rlabel polysilicon 65 -468 65 -468 0 1
rlabel polysilicon 68 -474 68 -474 0 4
rlabel polysilicon 72 -468 72 -468 0 1
rlabel polysilicon 75 -474 75 -474 0 4
rlabel polysilicon 82 -468 82 -468 0 2
rlabel polysilicon 79 -474 79 -474 0 3
rlabel polysilicon 86 -468 86 -468 0 1
rlabel polysilicon 86 -474 86 -474 0 3
rlabel polysilicon 93 -468 93 -468 0 1
rlabel polysilicon 93 -474 93 -474 0 3
rlabel polysilicon 100 -468 100 -468 0 1
rlabel polysilicon 103 -468 103 -468 0 2
rlabel polysilicon 107 -468 107 -468 0 1
rlabel polysilicon 107 -474 107 -474 0 3
rlabel polysilicon 114 -468 114 -468 0 1
rlabel polysilicon 114 -474 114 -474 0 3
rlabel polysilicon 121 -468 121 -468 0 1
rlabel polysilicon 121 -474 121 -474 0 3
rlabel polysilicon 128 -468 128 -468 0 1
rlabel polysilicon 128 -474 128 -474 0 3
rlabel polysilicon 135 -468 135 -468 0 1
rlabel polysilicon 135 -474 135 -474 0 3
rlabel polysilicon 142 -474 142 -474 0 3
rlabel polysilicon 145 -474 145 -474 0 4
rlabel polysilicon 149 -468 149 -468 0 1
rlabel polysilicon 149 -474 149 -474 0 3
rlabel polysilicon 156 -468 156 -468 0 1
rlabel polysilicon 156 -474 156 -474 0 3
rlabel polysilicon 166 -468 166 -468 0 2
rlabel polysilicon 163 -474 163 -474 0 3
rlabel polysilicon 170 -468 170 -468 0 1
rlabel polysilicon 170 -474 170 -474 0 3
rlabel polysilicon 177 -468 177 -468 0 1
rlabel polysilicon 180 -468 180 -468 0 2
rlabel polysilicon 177 -474 177 -474 0 3
rlabel polysilicon 180 -474 180 -474 0 4
rlabel polysilicon 184 -468 184 -468 0 1
rlabel polysilicon 187 -474 187 -474 0 4
rlabel polysilicon 191 -468 191 -468 0 1
rlabel polysilicon 194 -468 194 -468 0 2
rlabel polysilicon 191 -474 191 -474 0 3
rlabel polysilicon 198 -468 198 -468 0 1
rlabel polysilicon 198 -474 198 -474 0 3
rlabel polysilicon 205 -468 205 -468 0 1
rlabel polysilicon 205 -474 205 -474 0 3
rlabel polysilicon 212 -468 212 -468 0 1
rlabel polysilicon 212 -474 212 -474 0 3
rlabel polysilicon 219 -468 219 -468 0 1
rlabel polysilicon 219 -474 219 -474 0 3
rlabel polysilicon 226 -468 226 -468 0 1
rlabel polysilicon 226 -474 226 -474 0 3
rlabel polysilicon 233 -468 233 -468 0 1
rlabel polysilicon 233 -474 233 -474 0 3
rlabel polysilicon 240 -468 240 -468 0 1
rlabel polysilicon 240 -474 240 -474 0 3
rlabel polysilicon 247 -468 247 -468 0 1
rlabel polysilicon 247 -474 247 -474 0 3
rlabel polysilicon 254 -468 254 -468 0 1
rlabel polysilicon 254 -474 254 -474 0 3
rlabel polysilicon 261 -468 261 -468 0 1
rlabel polysilicon 261 -474 261 -474 0 3
rlabel polysilicon 268 -468 268 -468 0 1
rlabel polysilicon 268 -474 268 -474 0 3
rlabel polysilicon 275 -468 275 -468 0 1
rlabel polysilicon 275 -474 275 -474 0 3
rlabel polysilicon 282 -468 282 -468 0 1
rlabel polysilicon 282 -474 282 -474 0 3
rlabel polysilicon 289 -468 289 -468 0 1
rlabel polysilicon 289 -474 289 -474 0 3
rlabel polysilicon 296 -468 296 -468 0 1
rlabel polysilicon 296 -474 296 -474 0 3
rlabel polysilicon 303 -468 303 -468 0 1
rlabel polysilicon 303 -474 303 -474 0 3
rlabel polysilicon 313 -468 313 -468 0 2
rlabel polysilicon 310 -474 310 -474 0 3
rlabel polysilicon 317 -468 317 -468 0 1
rlabel polysilicon 317 -474 317 -474 0 3
rlabel polysilicon 324 -468 324 -468 0 1
rlabel polysilicon 324 -474 324 -474 0 3
rlabel polysilicon 331 -468 331 -468 0 1
rlabel polysilicon 331 -474 331 -474 0 3
rlabel polysilicon 338 -468 338 -468 0 1
rlabel polysilicon 338 -474 338 -474 0 3
rlabel polysilicon 345 -468 345 -468 0 1
rlabel polysilicon 345 -474 345 -474 0 3
rlabel polysilicon 352 -468 352 -468 0 1
rlabel polysilicon 352 -474 352 -474 0 3
rlabel polysilicon 359 -468 359 -468 0 1
rlabel polysilicon 359 -474 359 -474 0 3
rlabel polysilicon 366 -468 366 -468 0 1
rlabel polysilicon 366 -474 366 -474 0 3
rlabel polysilicon 373 -468 373 -468 0 1
rlabel polysilicon 373 -474 373 -474 0 3
rlabel polysilicon 380 -468 380 -468 0 1
rlabel polysilicon 383 -474 383 -474 0 4
rlabel polysilicon 387 -468 387 -468 0 1
rlabel polysilicon 390 -468 390 -468 0 2
rlabel polysilicon 387 -474 387 -474 0 3
rlabel polysilicon 390 -474 390 -474 0 4
rlabel polysilicon 394 -468 394 -468 0 1
rlabel polysilicon 394 -474 394 -474 0 3
rlabel polysilicon 401 -468 401 -468 0 1
rlabel polysilicon 401 -474 401 -474 0 3
rlabel polysilicon 408 -468 408 -468 0 1
rlabel polysilicon 411 -468 411 -468 0 2
rlabel polysilicon 408 -474 408 -474 0 3
rlabel polysilicon 411 -474 411 -474 0 4
rlabel polysilicon 418 -468 418 -468 0 2
rlabel polysilicon 422 -468 422 -468 0 1
rlabel polysilicon 425 -468 425 -468 0 2
rlabel polysilicon 429 -474 429 -474 0 3
rlabel polysilicon 432 -474 432 -474 0 4
rlabel polysilicon 436 -468 436 -468 0 1
rlabel polysilicon 439 -468 439 -468 0 2
rlabel polysilicon 439 -474 439 -474 0 4
rlabel polysilicon 446 -468 446 -468 0 2
rlabel polysilicon 443 -474 443 -474 0 3
rlabel polysilicon 446 -474 446 -474 0 4
rlabel polysilicon 453 -468 453 -468 0 2
rlabel polysilicon 453 -474 453 -474 0 4
rlabel polysilicon 457 -468 457 -468 0 1
rlabel polysilicon 457 -474 457 -474 0 3
rlabel polysilicon 464 -468 464 -468 0 1
rlabel polysilicon 464 -474 464 -474 0 3
rlabel polysilicon 471 -468 471 -468 0 1
rlabel polysilicon 471 -474 471 -474 0 3
rlabel polysilicon 478 -468 478 -468 0 1
rlabel polysilicon 478 -474 478 -474 0 3
rlabel polysilicon 485 -468 485 -468 0 1
rlabel polysilicon 485 -474 485 -474 0 3
rlabel polysilicon 492 -468 492 -468 0 1
rlabel polysilicon 492 -474 492 -474 0 3
rlabel polysilicon 499 -468 499 -468 0 1
rlabel polysilicon 499 -474 499 -474 0 3
rlabel polysilicon 506 -468 506 -468 0 1
rlabel polysilicon 506 -474 506 -474 0 3
rlabel polysilicon 513 -468 513 -468 0 1
rlabel polysilicon 513 -474 513 -474 0 3
rlabel polysilicon 520 -468 520 -468 0 1
rlabel polysilicon 520 -474 520 -474 0 3
rlabel polysilicon 527 -468 527 -468 0 1
rlabel polysilicon 527 -474 527 -474 0 3
rlabel polysilicon 534 -468 534 -468 0 1
rlabel polysilicon 534 -474 534 -474 0 3
rlabel polysilicon 541 -468 541 -468 0 1
rlabel polysilicon 541 -474 541 -474 0 3
rlabel polysilicon 548 -468 548 -468 0 1
rlabel polysilicon 548 -474 548 -474 0 3
rlabel polysilicon 555 -468 555 -468 0 1
rlabel polysilicon 555 -474 555 -474 0 3
rlabel polysilicon 562 -468 562 -468 0 1
rlabel polysilicon 562 -474 562 -474 0 3
rlabel polysilicon 569 -468 569 -468 0 1
rlabel polysilicon 569 -474 569 -474 0 3
rlabel polysilicon 576 -468 576 -468 0 1
rlabel polysilicon 576 -474 576 -474 0 3
rlabel polysilicon 583 -468 583 -468 0 1
rlabel polysilicon 583 -474 583 -474 0 3
rlabel polysilicon 590 -468 590 -468 0 1
rlabel polysilicon 590 -474 590 -474 0 3
rlabel polysilicon 597 -468 597 -468 0 1
rlabel polysilicon 597 -474 597 -474 0 3
rlabel polysilicon 604 -468 604 -468 0 1
rlabel polysilicon 604 -474 604 -474 0 3
rlabel polysilicon 611 -468 611 -468 0 1
rlabel polysilicon 611 -474 611 -474 0 3
rlabel polysilicon 625 -468 625 -468 0 1
rlabel polysilicon 625 -474 625 -474 0 3
rlabel polysilicon 632 -468 632 -468 0 1
rlabel polysilicon 632 -474 632 -474 0 3
rlabel polysilicon 639 -468 639 -468 0 1
rlabel polysilicon 639 -474 639 -474 0 3
rlabel polysilicon 646 -468 646 -468 0 1
rlabel polysilicon 646 -474 646 -474 0 3
rlabel polysilicon 653 -468 653 -468 0 1
rlabel polysilicon 653 -474 653 -474 0 3
rlabel polysilicon 667 -468 667 -468 0 1
rlabel polysilicon 667 -474 667 -474 0 3
rlabel polysilicon 674 -468 674 -468 0 1
rlabel polysilicon 674 -474 674 -474 0 3
rlabel polysilicon 681 -468 681 -468 0 1
rlabel polysilicon 681 -474 681 -474 0 3
rlabel polysilicon 688 -468 688 -468 0 1
rlabel polysilicon 688 -474 688 -474 0 3
rlabel polysilicon 695 -468 695 -468 0 1
rlabel polysilicon 695 -474 695 -474 0 3
rlabel polysilicon 702 -468 702 -468 0 1
rlabel polysilicon 702 -474 702 -474 0 3
rlabel polysilicon 709 -468 709 -468 0 1
rlabel polysilicon 716 -474 716 -474 0 3
rlabel polysilicon 719 -474 719 -474 0 4
rlabel polysilicon 723 -468 723 -468 0 1
rlabel polysilicon 723 -474 723 -474 0 3
rlabel polysilicon 730 -468 730 -468 0 1
rlabel polysilicon 730 -474 730 -474 0 3
rlabel polysilicon 23 -553 23 -553 0 1
rlabel polysilicon 23 -559 23 -559 0 3
rlabel polysilicon 40 -559 40 -559 0 4
rlabel polysilicon 44 -553 44 -553 0 1
rlabel polysilicon 44 -559 44 -559 0 3
rlabel polysilicon 51 -553 51 -553 0 1
rlabel polysilicon 51 -559 51 -559 0 3
rlabel polysilicon 54 -559 54 -559 0 4
rlabel polysilicon 61 -553 61 -553 0 2
rlabel polysilicon 61 -559 61 -559 0 4
rlabel polysilicon 65 -553 65 -553 0 1
rlabel polysilicon 68 -553 68 -553 0 2
rlabel polysilicon 65 -559 65 -559 0 3
rlabel polysilicon 75 -553 75 -553 0 2
rlabel polysilicon 72 -559 72 -559 0 3
rlabel polysilicon 75 -559 75 -559 0 4
rlabel polysilicon 79 -553 79 -553 0 1
rlabel polysilicon 79 -559 79 -559 0 3
rlabel polysilicon 86 -553 86 -553 0 1
rlabel polysilicon 86 -559 86 -559 0 3
rlabel polysilicon 93 -553 93 -553 0 1
rlabel polysilicon 93 -559 93 -559 0 3
rlabel polysilicon 103 -559 103 -559 0 4
rlabel polysilicon 107 -553 107 -553 0 1
rlabel polysilicon 107 -559 107 -559 0 3
rlabel polysilicon 114 -553 114 -553 0 1
rlabel polysilicon 114 -559 114 -559 0 3
rlabel polysilicon 121 -553 121 -553 0 1
rlabel polysilicon 124 -553 124 -553 0 2
rlabel polysilicon 128 -553 128 -553 0 1
rlabel polysilicon 128 -559 128 -559 0 3
rlabel polysilicon 135 -553 135 -553 0 1
rlabel polysilicon 135 -559 135 -559 0 3
rlabel polysilicon 145 -553 145 -553 0 2
rlabel polysilicon 142 -559 142 -559 0 3
rlabel polysilicon 152 -553 152 -553 0 2
rlabel polysilicon 156 -553 156 -553 0 1
rlabel polysilicon 156 -559 156 -559 0 3
rlabel polysilicon 163 -553 163 -553 0 1
rlabel polysilicon 163 -559 163 -559 0 3
rlabel polysilicon 166 -559 166 -559 0 4
rlabel polysilicon 170 -553 170 -553 0 1
rlabel polysilicon 170 -559 170 -559 0 3
rlabel polysilicon 177 -559 177 -559 0 3
rlabel polysilicon 184 -559 184 -559 0 3
rlabel polysilicon 187 -559 187 -559 0 4
rlabel polysilicon 191 -553 191 -553 0 1
rlabel polysilicon 191 -559 191 -559 0 3
rlabel polysilicon 198 -553 198 -553 0 1
rlabel polysilicon 198 -559 198 -559 0 3
rlabel polysilicon 205 -553 205 -553 0 1
rlabel polysilicon 205 -559 205 -559 0 3
rlabel polysilicon 212 -553 212 -553 0 1
rlabel polysilicon 212 -559 212 -559 0 3
rlabel polysilicon 215 -559 215 -559 0 4
rlabel polysilicon 219 -553 219 -553 0 1
rlabel polysilicon 219 -559 219 -559 0 3
rlabel polysilicon 226 -553 226 -553 0 1
rlabel polysilicon 226 -559 226 -559 0 3
rlabel polysilicon 233 -553 233 -553 0 1
rlabel polysilicon 233 -559 233 -559 0 3
rlabel polysilicon 236 -559 236 -559 0 4
rlabel polysilicon 240 -553 240 -553 0 1
rlabel polysilicon 243 -553 243 -553 0 2
rlabel polysilicon 240 -559 240 -559 0 3
rlabel polysilicon 247 -553 247 -553 0 1
rlabel polysilicon 247 -559 247 -559 0 3
rlabel polysilicon 254 -553 254 -553 0 1
rlabel polysilicon 254 -559 254 -559 0 3
rlabel polysilicon 261 -553 261 -553 0 1
rlabel polysilicon 261 -559 261 -559 0 3
rlabel polysilicon 268 -553 268 -553 0 1
rlabel polysilicon 268 -559 268 -559 0 3
rlabel polysilicon 275 -553 275 -553 0 1
rlabel polysilicon 275 -559 275 -559 0 3
rlabel polysilicon 282 -553 282 -553 0 1
rlabel polysilicon 282 -559 282 -559 0 3
rlabel polysilicon 289 -553 289 -553 0 1
rlabel polysilicon 289 -559 289 -559 0 3
rlabel polysilicon 296 -553 296 -553 0 1
rlabel polysilicon 296 -559 296 -559 0 3
rlabel polysilicon 303 -553 303 -553 0 1
rlabel polysilicon 303 -559 303 -559 0 3
rlabel polysilicon 306 -559 306 -559 0 4
rlabel polysilicon 310 -553 310 -553 0 1
rlabel polysilicon 310 -559 310 -559 0 3
rlabel polysilicon 317 -553 317 -553 0 1
rlabel polysilicon 320 -553 320 -553 0 2
rlabel polysilicon 317 -559 317 -559 0 3
rlabel polysilicon 320 -559 320 -559 0 4
rlabel polysilicon 324 -553 324 -553 0 1
rlabel polysilicon 324 -559 324 -559 0 3
rlabel polysilicon 331 -553 331 -553 0 1
rlabel polysilicon 331 -559 331 -559 0 3
rlabel polysilicon 338 -553 338 -553 0 1
rlabel polysilicon 338 -559 338 -559 0 3
rlabel polysilicon 345 -553 345 -553 0 1
rlabel polysilicon 345 -559 345 -559 0 3
rlabel polysilicon 352 -553 352 -553 0 1
rlabel polysilicon 352 -559 352 -559 0 3
rlabel polysilicon 359 -553 359 -553 0 1
rlabel polysilicon 359 -559 359 -559 0 3
rlabel polysilicon 369 -553 369 -553 0 2
rlabel polysilicon 366 -559 366 -559 0 3
rlabel polysilicon 369 -559 369 -559 0 4
rlabel polysilicon 373 -553 373 -553 0 1
rlabel polysilicon 373 -559 373 -559 0 3
rlabel polysilicon 380 -559 380 -559 0 3
rlabel polysilicon 383 -559 383 -559 0 4
rlabel polysilicon 387 -553 387 -553 0 1
rlabel polysilicon 387 -559 387 -559 0 3
rlabel polysilicon 397 -553 397 -553 0 2
rlabel polysilicon 394 -559 394 -559 0 3
rlabel polysilicon 397 -559 397 -559 0 4
rlabel polysilicon 401 -553 401 -553 0 1
rlabel polysilicon 401 -559 401 -559 0 3
rlabel polysilicon 408 -553 408 -553 0 1
rlabel polysilicon 408 -559 408 -559 0 3
rlabel polysilicon 415 -553 415 -553 0 1
rlabel polysilicon 415 -559 415 -559 0 3
rlabel polysilicon 422 -553 422 -553 0 1
rlabel polysilicon 425 -559 425 -559 0 4
rlabel polysilicon 432 -553 432 -553 0 2
rlabel polysilicon 429 -559 429 -559 0 3
rlabel polysilicon 432 -559 432 -559 0 4
rlabel polysilicon 436 -553 436 -553 0 1
rlabel polysilicon 436 -559 436 -559 0 3
rlabel polysilicon 443 -553 443 -553 0 1
rlabel polysilicon 446 -553 446 -553 0 2
rlabel polysilicon 446 -559 446 -559 0 4
rlabel polysilicon 450 -553 450 -553 0 1
rlabel polysilicon 450 -559 450 -559 0 3
rlabel polysilicon 457 -553 457 -553 0 1
rlabel polysilicon 457 -559 457 -559 0 3
rlabel polysilicon 464 -553 464 -553 0 1
rlabel polysilicon 464 -559 464 -559 0 3
rlabel polysilicon 471 -553 471 -553 0 1
rlabel polysilicon 471 -559 471 -559 0 3
rlabel polysilicon 478 -553 478 -553 0 1
rlabel polysilicon 478 -559 478 -559 0 3
rlabel polysilicon 485 -553 485 -553 0 1
rlabel polysilicon 485 -559 485 -559 0 3
rlabel polysilicon 492 -553 492 -553 0 1
rlabel polysilicon 492 -559 492 -559 0 3
rlabel polysilicon 499 -553 499 -553 0 1
rlabel polysilicon 499 -559 499 -559 0 3
rlabel polysilicon 506 -553 506 -553 0 1
rlabel polysilicon 506 -559 506 -559 0 3
rlabel polysilicon 513 -553 513 -553 0 1
rlabel polysilicon 513 -559 513 -559 0 3
rlabel polysilicon 520 -553 520 -553 0 1
rlabel polysilicon 520 -559 520 -559 0 3
rlabel polysilicon 527 -553 527 -553 0 1
rlabel polysilicon 527 -559 527 -559 0 3
rlabel polysilicon 534 -553 534 -553 0 1
rlabel polysilicon 534 -559 534 -559 0 3
rlabel polysilicon 541 -553 541 -553 0 1
rlabel polysilicon 541 -559 541 -559 0 3
rlabel polysilicon 548 -553 548 -553 0 1
rlabel polysilicon 548 -559 548 -559 0 3
rlabel polysilicon 555 -553 555 -553 0 1
rlabel polysilicon 555 -559 555 -559 0 3
rlabel polysilicon 562 -553 562 -553 0 1
rlabel polysilicon 562 -559 562 -559 0 3
rlabel polysilicon 569 -553 569 -553 0 1
rlabel polysilicon 569 -559 569 -559 0 3
rlabel polysilicon 576 -553 576 -553 0 1
rlabel polysilicon 576 -559 576 -559 0 3
rlabel polysilicon 583 -553 583 -553 0 1
rlabel polysilicon 583 -559 583 -559 0 3
rlabel polysilicon 590 -553 590 -553 0 1
rlabel polysilicon 590 -559 590 -559 0 3
rlabel polysilicon 597 -553 597 -553 0 1
rlabel polysilicon 597 -559 597 -559 0 3
rlabel polysilicon 604 -553 604 -553 0 1
rlabel polysilicon 604 -559 604 -559 0 3
rlabel polysilicon 611 -553 611 -553 0 1
rlabel polysilicon 611 -559 611 -559 0 3
rlabel polysilicon 618 -553 618 -553 0 1
rlabel polysilicon 618 -559 618 -559 0 3
rlabel polysilicon 625 -553 625 -553 0 1
rlabel polysilicon 625 -559 625 -559 0 3
rlabel polysilicon 632 -553 632 -553 0 1
rlabel polysilicon 632 -559 632 -559 0 3
rlabel polysilicon 639 -553 639 -553 0 1
rlabel polysilicon 639 -559 639 -559 0 3
rlabel polysilicon 646 -553 646 -553 0 1
rlabel polysilicon 646 -559 646 -559 0 3
rlabel polysilicon 653 -553 653 -553 0 1
rlabel polysilicon 653 -559 653 -559 0 3
rlabel polysilicon 660 -553 660 -553 0 1
rlabel polysilicon 660 -559 660 -559 0 3
rlabel polysilicon 667 -553 667 -553 0 1
rlabel polysilicon 667 -559 667 -559 0 3
rlabel polysilicon 674 -553 674 -553 0 1
rlabel polysilicon 674 -559 674 -559 0 3
rlabel polysilicon 681 -553 681 -553 0 1
rlabel polysilicon 681 -559 681 -559 0 3
rlabel polysilicon 688 -553 688 -553 0 1
rlabel polysilicon 688 -559 688 -559 0 3
rlabel polysilicon 695 -553 695 -553 0 1
rlabel polysilicon 695 -559 695 -559 0 3
rlabel polysilicon 702 -553 702 -553 0 1
rlabel polysilicon 702 -559 702 -559 0 3
rlabel polysilicon 709 -553 709 -553 0 1
rlabel polysilicon 709 -559 709 -559 0 3
rlabel polysilicon 716 -553 716 -553 0 1
rlabel polysilicon 716 -559 716 -559 0 3
rlabel polysilicon 723 -553 723 -553 0 1
rlabel polysilicon 723 -559 723 -559 0 3
rlabel polysilicon 730 -553 730 -553 0 1
rlabel polysilicon 730 -559 730 -559 0 3
rlabel polysilicon 737 -553 737 -553 0 1
rlabel polysilicon 737 -559 737 -559 0 3
rlabel polysilicon 744 -553 744 -553 0 1
rlabel polysilicon 744 -559 744 -559 0 3
rlabel polysilicon 751 -553 751 -553 0 1
rlabel polysilicon 751 -559 751 -559 0 3
rlabel polysilicon 779 -553 779 -553 0 1
rlabel polysilicon 779 -559 779 -559 0 3
rlabel polysilicon 16 -646 16 -646 0 1
rlabel polysilicon 16 -652 16 -652 0 3
rlabel polysilicon 23 -646 23 -646 0 1
rlabel polysilicon 23 -652 23 -652 0 3
rlabel polysilicon 30 -646 30 -646 0 1
rlabel polysilicon 33 -646 33 -646 0 2
rlabel polysilicon 40 -646 40 -646 0 2
rlabel polysilicon 47 -646 47 -646 0 2
rlabel polysilicon 44 -652 44 -652 0 3
rlabel polysilicon 47 -652 47 -652 0 4
rlabel polysilicon 51 -646 51 -646 0 1
rlabel polysilicon 51 -652 51 -652 0 3
rlabel polysilicon 58 -646 58 -646 0 1
rlabel polysilicon 58 -652 58 -652 0 3
rlabel polysilicon 65 -646 65 -646 0 1
rlabel polysilicon 65 -652 65 -652 0 3
rlabel polysilicon 72 -646 72 -646 0 1
rlabel polysilicon 72 -652 72 -652 0 3
rlabel polysilicon 79 -646 79 -646 0 1
rlabel polysilicon 79 -652 79 -652 0 3
rlabel polysilicon 86 -646 86 -646 0 1
rlabel polysilicon 86 -652 86 -652 0 3
rlabel polysilicon 93 -646 93 -646 0 1
rlabel polysilicon 96 -646 96 -646 0 2
rlabel polysilicon 100 -646 100 -646 0 1
rlabel polysilicon 100 -652 100 -652 0 3
rlabel polysilicon 107 -652 107 -652 0 3
rlabel polysilicon 110 -652 110 -652 0 4
rlabel polysilicon 114 -652 114 -652 0 3
rlabel polysilicon 117 -652 117 -652 0 4
rlabel polysilicon 124 -646 124 -646 0 2
rlabel polysilicon 121 -652 121 -652 0 3
rlabel polysilicon 124 -652 124 -652 0 4
rlabel polysilicon 128 -646 128 -646 0 1
rlabel polysilicon 131 -652 131 -652 0 4
rlabel polysilicon 135 -646 135 -646 0 1
rlabel polysilicon 135 -652 135 -652 0 3
rlabel polysilicon 142 -646 142 -646 0 1
rlabel polysilicon 142 -652 142 -652 0 3
rlabel polysilicon 145 -652 145 -652 0 4
rlabel polysilicon 149 -646 149 -646 0 1
rlabel polysilicon 152 -652 152 -652 0 4
rlabel polysilicon 156 -646 156 -646 0 1
rlabel polysilicon 156 -652 156 -652 0 3
rlabel polysilicon 163 -652 163 -652 0 3
rlabel polysilicon 166 -652 166 -652 0 4
rlabel polysilicon 170 -646 170 -646 0 1
rlabel polysilicon 170 -652 170 -652 0 3
rlabel polysilicon 177 -646 177 -646 0 1
rlabel polysilicon 177 -652 177 -652 0 3
rlabel polysilicon 184 -646 184 -646 0 1
rlabel polysilicon 187 -646 187 -646 0 2
rlabel polysilicon 184 -652 184 -652 0 3
rlabel polysilicon 191 -646 191 -646 0 1
rlabel polysilicon 191 -652 191 -652 0 3
rlabel polysilicon 198 -646 198 -646 0 1
rlabel polysilicon 198 -652 198 -652 0 3
rlabel polysilicon 205 -646 205 -646 0 1
rlabel polysilicon 205 -652 205 -652 0 3
rlabel polysilicon 212 -646 212 -646 0 1
rlabel polysilicon 212 -652 212 -652 0 3
rlabel polysilicon 219 -646 219 -646 0 1
rlabel polysilicon 219 -652 219 -652 0 3
rlabel polysilicon 226 -646 226 -646 0 1
rlabel polysilicon 226 -652 226 -652 0 3
rlabel polysilicon 233 -646 233 -646 0 1
rlabel polysilicon 233 -652 233 -652 0 3
rlabel polysilicon 240 -646 240 -646 0 1
rlabel polysilicon 240 -652 240 -652 0 3
rlabel polysilicon 247 -646 247 -646 0 1
rlabel polysilicon 247 -652 247 -652 0 3
rlabel polysilicon 254 -646 254 -646 0 1
rlabel polysilicon 254 -652 254 -652 0 3
rlabel polysilicon 261 -646 261 -646 0 1
rlabel polysilicon 261 -652 261 -652 0 3
rlabel polysilicon 268 -646 268 -646 0 1
rlabel polysilicon 268 -652 268 -652 0 3
rlabel polysilicon 275 -646 275 -646 0 1
rlabel polysilicon 278 -646 278 -646 0 2
rlabel polysilicon 275 -652 275 -652 0 3
rlabel polysilicon 278 -652 278 -652 0 4
rlabel polysilicon 282 -646 282 -646 0 1
rlabel polysilicon 282 -652 282 -652 0 3
rlabel polysilicon 289 -646 289 -646 0 1
rlabel polysilicon 292 -646 292 -646 0 2
rlabel polysilicon 289 -652 289 -652 0 3
rlabel polysilicon 292 -652 292 -652 0 4
rlabel polysilicon 296 -646 296 -646 0 1
rlabel polysilicon 296 -652 296 -652 0 3
rlabel polysilicon 303 -646 303 -646 0 1
rlabel polysilicon 303 -652 303 -652 0 3
rlabel polysilicon 310 -646 310 -646 0 1
rlabel polysilicon 310 -652 310 -652 0 3
rlabel polysilicon 317 -646 317 -646 0 1
rlabel polysilicon 317 -652 317 -652 0 3
rlabel polysilicon 324 -646 324 -646 0 1
rlabel polysilicon 324 -652 324 -652 0 3
rlabel polysilicon 331 -646 331 -646 0 1
rlabel polysilicon 331 -652 331 -652 0 3
rlabel polysilicon 338 -646 338 -646 0 1
rlabel polysilicon 338 -652 338 -652 0 3
rlabel polysilicon 345 -646 345 -646 0 1
rlabel polysilicon 348 -646 348 -646 0 2
rlabel polysilicon 348 -652 348 -652 0 4
rlabel polysilicon 352 -646 352 -646 0 1
rlabel polysilicon 355 -646 355 -646 0 2
rlabel polysilicon 352 -652 352 -652 0 3
rlabel polysilicon 359 -646 359 -646 0 1
rlabel polysilicon 359 -652 359 -652 0 3
rlabel polysilicon 366 -646 366 -646 0 1
rlabel polysilicon 369 -646 369 -646 0 2
rlabel polysilicon 366 -652 366 -652 0 3
rlabel polysilicon 369 -652 369 -652 0 4
rlabel polysilicon 373 -646 373 -646 0 1
rlabel polysilicon 373 -652 373 -652 0 3
rlabel polysilicon 380 -646 380 -646 0 1
rlabel polysilicon 380 -652 380 -652 0 3
rlabel polysilicon 387 -646 387 -646 0 1
rlabel polysilicon 390 -646 390 -646 0 2
rlabel polysilicon 390 -652 390 -652 0 4
rlabel polysilicon 394 -646 394 -646 0 1
rlabel polysilicon 394 -652 394 -652 0 3
rlabel polysilicon 401 -646 401 -646 0 1
rlabel polysilicon 401 -652 401 -652 0 3
rlabel polysilicon 411 -646 411 -646 0 2
rlabel polysilicon 408 -652 408 -652 0 3
rlabel polysilicon 411 -652 411 -652 0 4
rlabel polysilicon 415 -646 415 -646 0 1
rlabel polysilicon 418 -646 418 -646 0 2
rlabel polysilicon 418 -652 418 -652 0 4
rlabel polysilicon 425 -646 425 -646 0 2
rlabel polysilicon 422 -652 422 -652 0 3
rlabel polysilicon 429 -646 429 -646 0 1
rlabel polysilicon 429 -652 429 -652 0 3
rlabel polysilicon 436 -646 436 -646 0 1
rlabel polysilicon 436 -652 436 -652 0 3
rlabel polysilicon 443 -646 443 -646 0 1
rlabel polysilicon 446 -646 446 -646 0 2
rlabel polysilicon 443 -652 443 -652 0 3
rlabel polysilicon 446 -652 446 -652 0 4
rlabel polysilicon 450 -646 450 -646 0 1
rlabel polysilicon 450 -652 450 -652 0 3
rlabel polysilicon 457 -646 457 -646 0 1
rlabel polysilicon 457 -652 457 -652 0 3
rlabel polysilicon 464 -646 464 -646 0 1
rlabel polysilicon 464 -652 464 -652 0 3
rlabel polysilicon 471 -646 471 -646 0 1
rlabel polysilicon 471 -652 471 -652 0 3
rlabel polysilicon 478 -646 478 -646 0 1
rlabel polysilicon 478 -652 478 -652 0 3
rlabel polysilicon 485 -646 485 -646 0 1
rlabel polysilicon 485 -652 485 -652 0 3
rlabel polysilicon 499 -646 499 -646 0 1
rlabel polysilicon 499 -652 499 -652 0 3
rlabel polysilicon 506 -646 506 -646 0 1
rlabel polysilicon 506 -652 506 -652 0 3
rlabel polysilicon 513 -646 513 -646 0 1
rlabel polysilicon 516 -646 516 -646 0 2
rlabel polysilicon 520 -646 520 -646 0 1
rlabel polysilicon 520 -652 520 -652 0 3
rlabel polysilicon 527 -646 527 -646 0 1
rlabel polysilicon 527 -652 527 -652 0 3
rlabel polysilicon 534 -646 534 -646 0 1
rlabel polysilicon 534 -652 534 -652 0 3
rlabel polysilicon 541 -646 541 -646 0 1
rlabel polysilicon 541 -652 541 -652 0 3
rlabel polysilicon 548 -646 548 -646 0 1
rlabel polysilicon 548 -652 548 -652 0 3
rlabel polysilicon 555 -646 555 -646 0 1
rlabel polysilicon 555 -652 555 -652 0 3
rlabel polysilicon 562 -646 562 -646 0 1
rlabel polysilicon 562 -652 562 -652 0 3
rlabel polysilicon 569 -646 569 -646 0 1
rlabel polysilicon 569 -652 569 -652 0 3
rlabel polysilicon 576 -646 576 -646 0 1
rlabel polysilicon 576 -652 576 -652 0 3
rlabel polysilicon 583 -646 583 -646 0 1
rlabel polysilicon 583 -652 583 -652 0 3
rlabel polysilicon 590 -646 590 -646 0 1
rlabel polysilicon 590 -652 590 -652 0 3
rlabel polysilicon 597 -646 597 -646 0 1
rlabel polysilicon 597 -652 597 -652 0 3
rlabel polysilicon 604 -646 604 -646 0 1
rlabel polysilicon 604 -652 604 -652 0 3
rlabel polysilicon 611 -646 611 -646 0 1
rlabel polysilicon 611 -652 611 -652 0 3
rlabel polysilicon 618 -646 618 -646 0 1
rlabel polysilicon 618 -652 618 -652 0 3
rlabel polysilicon 625 -646 625 -646 0 1
rlabel polysilicon 625 -652 625 -652 0 3
rlabel polysilicon 632 -646 632 -646 0 1
rlabel polysilicon 632 -652 632 -652 0 3
rlabel polysilicon 639 -646 639 -646 0 1
rlabel polysilicon 639 -652 639 -652 0 3
rlabel polysilicon 646 -646 646 -646 0 1
rlabel polysilicon 646 -652 646 -652 0 3
rlabel polysilicon 653 -646 653 -646 0 1
rlabel polysilicon 653 -652 653 -652 0 3
rlabel polysilicon 660 -646 660 -646 0 1
rlabel polysilicon 667 -646 667 -646 0 1
rlabel polysilicon 667 -652 667 -652 0 3
rlabel polysilicon 674 -646 674 -646 0 1
rlabel polysilicon 674 -652 674 -652 0 3
rlabel polysilicon 681 -646 681 -646 0 1
rlabel polysilicon 681 -652 681 -652 0 3
rlabel polysilicon 688 -646 688 -646 0 1
rlabel polysilicon 688 -652 688 -652 0 3
rlabel polysilicon 695 -646 695 -646 0 1
rlabel polysilicon 695 -652 695 -652 0 3
rlabel polysilicon 702 -646 702 -646 0 1
rlabel polysilicon 702 -652 702 -652 0 3
rlabel polysilicon 709 -646 709 -646 0 1
rlabel polysilicon 709 -652 709 -652 0 3
rlabel polysilicon 716 -646 716 -646 0 1
rlabel polysilicon 716 -652 716 -652 0 3
rlabel polysilicon 723 -646 723 -646 0 1
rlabel polysilicon 723 -652 723 -652 0 3
rlabel polysilicon 730 -646 730 -646 0 1
rlabel polysilicon 730 -652 730 -652 0 3
rlabel polysilicon 737 -646 737 -646 0 1
rlabel polysilicon 737 -652 737 -652 0 3
rlabel polysilicon 807 -646 807 -646 0 1
rlabel polysilicon 807 -652 807 -652 0 3
rlabel polysilicon 9 -727 9 -727 0 1
rlabel polysilicon 9 -733 9 -733 0 3
rlabel polysilicon 16 -727 16 -727 0 1
rlabel polysilicon 16 -733 16 -733 0 3
rlabel polysilicon 23 -727 23 -727 0 1
rlabel polysilicon 23 -733 23 -733 0 3
rlabel polysilicon 30 -727 30 -727 0 1
rlabel polysilicon 30 -733 30 -733 0 3
rlabel polysilicon 37 -727 37 -727 0 1
rlabel polysilicon 37 -733 37 -733 0 3
rlabel polysilicon 44 -727 44 -727 0 1
rlabel polysilicon 44 -733 44 -733 0 3
rlabel polysilicon 51 -733 51 -733 0 3
rlabel polysilicon 58 -727 58 -727 0 1
rlabel polysilicon 58 -733 58 -733 0 3
rlabel polysilicon 65 -727 65 -727 0 1
rlabel polysilicon 65 -733 65 -733 0 3
rlabel polysilicon 68 -733 68 -733 0 4
rlabel polysilicon 72 -733 72 -733 0 3
rlabel polysilicon 75 -733 75 -733 0 4
rlabel polysilicon 79 -727 79 -727 0 1
rlabel polysilicon 79 -733 79 -733 0 3
rlabel polysilicon 86 -727 86 -727 0 1
rlabel polysilicon 86 -733 86 -733 0 3
rlabel polysilicon 93 -727 93 -727 0 1
rlabel polysilicon 96 -727 96 -727 0 2
rlabel polysilicon 93 -733 93 -733 0 3
rlabel polysilicon 100 -727 100 -727 0 1
rlabel polysilicon 100 -733 100 -733 0 3
rlabel polysilicon 107 -727 107 -727 0 1
rlabel polysilicon 107 -733 107 -733 0 3
rlabel polysilicon 114 -727 114 -727 0 1
rlabel polysilicon 117 -727 117 -727 0 2
rlabel polysilicon 117 -733 117 -733 0 4
rlabel polysilicon 121 -727 121 -727 0 1
rlabel polysilicon 124 -727 124 -727 0 2
rlabel polysilicon 124 -733 124 -733 0 4
rlabel polysilicon 128 -727 128 -727 0 1
rlabel polysilicon 128 -733 128 -733 0 3
rlabel polysilicon 135 -727 135 -727 0 1
rlabel polysilicon 135 -733 135 -733 0 3
rlabel polysilicon 142 -727 142 -727 0 1
rlabel polysilicon 142 -733 142 -733 0 3
rlabel polysilicon 149 -727 149 -727 0 1
rlabel polysilicon 149 -733 149 -733 0 3
rlabel polysilicon 156 -727 156 -727 0 1
rlabel polysilicon 156 -733 156 -733 0 3
rlabel polysilicon 159 -733 159 -733 0 4
rlabel polysilicon 163 -727 163 -727 0 1
rlabel polysilicon 166 -727 166 -727 0 2
rlabel polysilicon 173 -727 173 -727 0 2
rlabel polysilicon 177 -727 177 -727 0 1
rlabel polysilicon 177 -733 177 -733 0 3
rlabel polysilicon 184 -727 184 -727 0 1
rlabel polysilicon 184 -733 184 -733 0 3
rlabel polysilicon 191 -727 191 -727 0 1
rlabel polysilicon 191 -733 191 -733 0 3
rlabel polysilicon 198 -727 198 -727 0 1
rlabel polysilicon 198 -733 198 -733 0 3
rlabel polysilicon 205 -727 205 -727 0 1
rlabel polysilicon 205 -733 205 -733 0 3
rlabel polysilicon 212 -727 212 -727 0 1
rlabel polysilicon 212 -733 212 -733 0 3
rlabel polysilicon 219 -727 219 -727 0 1
rlabel polysilicon 219 -733 219 -733 0 3
rlabel polysilicon 226 -727 226 -727 0 1
rlabel polysilicon 226 -733 226 -733 0 3
rlabel polysilicon 233 -727 233 -727 0 1
rlabel polysilicon 236 -727 236 -727 0 2
rlabel polysilicon 233 -733 233 -733 0 3
rlabel polysilicon 236 -733 236 -733 0 4
rlabel polysilicon 240 -727 240 -727 0 1
rlabel polysilicon 243 -727 243 -727 0 2
rlabel polysilicon 240 -733 240 -733 0 3
rlabel polysilicon 247 -727 247 -727 0 1
rlabel polysilicon 247 -733 247 -733 0 3
rlabel polysilicon 254 -727 254 -727 0 1
rlabel polysilicon 257 -727 257 -727 0 2
rlabel polysilicon 261 -727 261 -727 0 1
rlabel polysilicon 261 -733 261 -733 0 3
rlabel polysilicon 268 -727 268 -727 0 1
rlabel polysilicon 268 -733 268 -733 0 3
rlabel polysilicon 275 -727 275 -727 0 1
rlabel polysilicon 275 -733 275 -733 0 3
rlabel polysilicon 282 -727 282 -727 0 1
rlabel polysilicon 282 -733 282 -733 0 3
rlabel polysilicon 289 -727 289 -727 0 1
rlabel polysilicon 289 -733 289 -733 0 3
rlabel polysilicon 292 -733 292 -733 0 4
rlabel polysilicon 296 -727 296 -727 0 1
rlabel polysilicon 296 -733 296 -733 0 3
rlabel polysilicon 303 -727 303 -727 0 1
rlabel polysilicon 303 -733 303 -733 0 3
rlabel polysilicon 310 -727 310 -727 0 1
rlabel polysilicon 310 -733 310 -733 0 3
rlabel polysilicon 317 -727 317 -727 0 1
rlabel polysilicon 317 -733 317 -733 0 3
rlabel polysilicon 324 -727 324 -727 0 1
rlabel polysilicon 324 -733 324 -733 0 3
rlabel polysilicon 331 -727 331 -727 0 1
rlabel polysilicon 334 -727 334 -727 0 2
rlabel polysilicon 331 -733 331 -733 0 3
rlabel polysilicon 338 -727 338 -727 0 1
rlabel polysilicon 338 -733 338 -733 0 3
rlabel polysilicon 345 -727 345 -727 0 1
rlabel polysilicon 345 -733 345 -733 0 3
rlabel polysilicon 352 -727 352 -727 0 1
rlabel polysilicon 352 -733 352 -733 0 3
rlabel polysilicon 359 -727 359 -727 0 1
rlabel polysilicon 359 -733 359 -733 0 3
rlabel polysilicon 369 -727 369 -727 0 2
rlabel polysilicon 366 -733 366 -733 0 3
rlabel polysilicon 373 -727 373 -727 0 1
rlabel polysilicon 373 -733 373 -733 0 3
rlabel polysilicon 380 -727 380 -727 0 1
rlabel polysilicon 380 -733 380 -733 0 3
rlabel polysilicon 387 -727 387 -727 0 1
rlabel polysilicon 387 -733 387 -733 0 3
rlabel polysilicon 394 -727 394 -727 0 1
rlabel polysilicon 397 -727 397 -727 0 2
rlabel polysilicon 394 -733 394 -733 0 3
rlabel polysilicon 401 -727 401 -727 0 1
rlabel polysilicon 401 -733 401 -733 0 3
rlabel polysilicon 408 -727 408 -727 0 1
rlabel polysilicon 411 -727 411 -727 0 2
rlabel polysilicon 408 -733 408 -733 0 3
rlabel polysilicon 411 -733 411 -733 0 4
rlabel polysilicon 415 -727 415 -727 0 1
rlabel polysilicon 415 -733 415 -733 0 3
rlabel polysilicon 422 -727 422 -727 0 1
rlabel polysilicon 422 -733 422 -733 0 3
rlabel polysilicon 429 -727 429 -727 0 1
rlabel polysilicon 432 -727 432 -727 0 2
rlabel polysilicon 429 -733 429 -733 0 3
rlabel polysilicon 436 -727 436 -727 0 1
rlabel polysilicon 439 -727 439 -727 0 2
rlabel polysilicon 436 -733 436 -733 0 3
rlabel polysilicon 443 -727 443 -727 0 1
rlabel polysilicon 443 -733 443 -733 0 3
rlabel polysilicon 450 -733 450 -733 0 3
rlabel polysilicon 457 -727 457 -727 0 1
rlabel polysilicon 457 -733 457 -733 0 3
rlabel polysilicon 467 -727 467 -727 0 2
rlabel polysilicon 464 -733 464 -733 0 3
rlabel polysilicon 467 -733 467 -733 0 4
rlabel polysilicon 474 -727 474 -727 0 2
rlabel polysilicon 471 -733 471 -733 0 3
rlabel polysilicon 474 -733 474 -733 0 4
rlabel polysilicon 478 -727 478 -727 0 1
rlabel polysilicon 478 -733 478 -733 0 3
rlabel polysilicon 485 -727 485 -727 0 1
rlabel polysilicon 485 -733 485 -733 0 3
rlabel polysilicon 492 -727 492 -727 0 1
rlabel polysilicon 492 -733 492 -733 0 3
rlabel polysilicon 499 -727 499 -727 0 1
rlabel polysilicon 499 -733 499 -733 0 3
rlabel polysilicon 506 -727 506 -727 0 1
rlabel polysilicon 506 -733 506 -733 0 3
rlabel polysilicon 513 -727 513 -727 0 1
rlabel polysilicon 513 -733 513 -733 0 3
rlabel polysilicon 520 -727 520 -727 0 1
rlabel polysilicon 520 -733 520 -733 0 3
rlabel polysilicon 527 -727 527 -727 0 1
rlabel polysilicon 527 -733 527 -733 0 3
rlabel polysilicon 534 -727 534 -727 0 1
rlabel polysilicon 534 -733 534 -733 0 3
rlabel polysilicon 541 -727 541 -727 0 1
rlabel polysilicon 541 -733 541 -733 0 3
rlabel polysilicon 548 -727 548 -727 0 1
rlabel polysilicon 548 -733 548 -733 0 3
rlabel polysilicon 555 -727 555 -727 0 1
rlabel polysilicon 555 -733 555 -733 0 3
rlabel polysilicon 562 -727 562 -727 0 1
rlabel polysilicon 562 -733 562 -733 0 3
rlabel polysilicon 569 -727 569 -727 0 1
rlabel polysilicon 569 -733 569 -733 0 3
rlabel polysilicon 576 -727 576 -727 0 1
rlabel polysilicon 576 -733 576 -733 0 3
rlabel polysilicon 583 -727 583 -727 0 1
rlabel polysilicon 583 -733 583 -733 0 3
rlabel polysilicon 590 -727 590 -727 0 1
rlabel polysilicon 590 -733 590 -733 0 3
rlabel polysilicon 600 -733 600 -733 0 4
rlabel polysilicon 604 -727 604 -727 0 1
rlabel polysilicon 604 -733 604 -733 0 3
rlabel polysilicon 611 -727 611 -727 0 1
rlabel polysilicon 611 -733 611 -733 0 3
rlabel polysilicon 618 -727 618 -727 0 1
rlabel polysilicon 618 -733 618 -733 0 3
rlabel polysilicon 625 -727 625 -727 0 1
rlabel polysilicon 625 -733 625 -733 0 3
rlabel polysilicon 632 -727 632 -727 0 1
rlabel polysilicon 632 -733 632 -733 0 3
rlabel polysilicon 639 -727 639 -727 0 1
rlabel polysilicon 639 -733 639 -733 0 3
rlabel polysilicon 646 -727 646 -727 0 1
rlabel polysilicon 646 -733 646 -733 0 3
rlabel polysilicon 653 -727 653 -727 0 1
rlabel polysilicon 653 -733 653 -733 0 3
rlabel polysilicon 660 -727 660 -727 0 1
rlabel polysilicon 660 -733 660 -733 0 3
rlabel polysilicon 667 -727 667 -727 0 1
rlabel polysilicon 667 -733 667 -733 0 3
rlabel polysilicon 674 -727 674 -727 0 1
rlabel polysilicon 674 -733 674 -733 0 3
rlabel polysilicon 681 -727 681 -727 0 1
rlabel polysilicon 681 -733 681 -733 0 3
rlabel polysilicon 688 -727 688 -727 0 1
rlabel polysilicon 688 -733 688 -733 0 3
rlabel polysilicon 695 -727 695 -727 0 1
rlabel polysilicon 695 -733 695 -733 0 3
rlabel polysilicon 702 -727 702 -727 0 1
rlabel polysilicon 702 -733 702 -733 0 3
rlabel polysilicon 709 -727 709 -727 0 1
rlabel polysilicon 709 -733 709 -733 0 3
rlabel polysilicon 716 -727 716 -727 0 1
rlabel polysilicon 716 -733 716 -733 0 3
rlabel polysilicon 723 -727 723 -727 0 1
rlabel polysilicon 723 -733 723 -733 0 3
rlabel polysilicon 730 -727 730 -727 0 1
rlabel polysilicon 730 -733 730 -733 0 3
rlabel polysilicon 737 -727 737 -727 0 1
rlabel polysilicon 737 -733 737 -733 0 3
rlabel polysilicon 744 -727 744 -727 0 1
rlabel polysilicon 744 -733 744 -733 0 3
rlabel polysilicon 751 -727 751 -727 0 1
rlabel polysilicon 751 -733 751 -733 0 3
rlabel polysilicon 758 -727 758 -727 0 1
rlabel polysilicon 758 -733 758 -733 0 3
rlabel polysilicon 765 -727 765 -727 0 1
rlabel polysilicon 765 -733 765 -733 0 3
rlabel polysilicon 772 -727 772 -727 0 1
rlabel polysilicon 772 -733 772 -733 0 3
rlabel polysilicon 779 -727 779 -727 0 1
rlabel polysilicon 779 -733 779 -733 0 3
rlabel polysilicon 786 -727 786 -727 0 1
rlabel polysilicon 786 -733 786 -733 0 3
rlabel polysilicon 793 -727 793 -727 0 1
rlabel polysilicon 793 -733 793 -733 0 3
rlabel polysilicon 800 -727 800 -727 0 1
rlabel polysilicon 800 -733 800 -733 0 3
rlabel polysilicon 807 -727 807 -727 0 1
rlabel polysilicon 807 -733 807 -733 0 3
rlabel polysilicon 814 -727 814 -727 0 1
rlabel polysilicon 814 -733 814 -733 0 3
rlabel polysilicon 817 -733 817 -733 0 4
rlabel polysilicon 824 -727 824 -727 0 2
rlabel polysilicon 821 -733 821 -733 0 3
rlabel polysilicon 824 -733 824 -733 0 4
rlabel polysilicon 828 -727 828 -727 0 1
rlabel polysilicon 828 -733 828 -733 0 3
rlabel polysilicon 9 -816 9 -816 0 1
rlabel polysilicon 9 -822 9 -822 0 3
rlabel polysilicon 16 -816 16 -816 0 1
rlabel polysilicon 23 -816 23 -816 0 1
rlabel polysilicon 23 -822 23 -822 0 3
rlabel polysilicon 30 -816 30 -816 0 1
rlabel polysilicon 30 -822 30 -822 0 3
rlabel polysilicon 37 -816 37 -816 0 1
rlabel polysilicon 40 -816 40 -816 0 2
rlabel polysilicon 37 -822 37 -822 0 3
rlabel polysilicon 47 -816 47 -816 0 2
rlabel polysilicon 44 -822 44 -822 0 3
rlabel polysilicon 51 -822 51 -822 0 3
rlabel polysilicon 58 -816 58 -816 0 1
rlabel polysilicon 58 -822 58 -822 0 3
rlabel polysilicon 65 -822 65 -822 0 3
rlabel polysilicon 68 -822 68 -822 0 4
rlabel polysilicon 72 -816 72 -816 0 1
rlabel polysilicon 72 -822 72 -822 0 3
rlabel polysilicon 82 -816 82 -816 0 2
rlabel polysilicon 82 -822 82 -822 0 4
rlabel polysilicon 86 -816 86 -816 0 1
rlabel polysilicon 86 -822 86 -822 0 3
rlabel polysilicon 93 -816 93 -816 0 1
rlabel polysilicon 96 -816 96 -816 0 2
rlabel polysilicon 93 -822 93 -822 0 3
rlabel polysilicon 96 -822 96 -822 0 4
rlabel polysilicon 100 -816 100 -816 0 1
rlabel polysilicon 100 -822 100 -822 0 3
rlabel polysilicon 107 -816 107 -816 0 1
rlabel polysilicon 107 -822 107 -822 0 3
rlabel polysilicon 114 -816 114 -816 0 1
rlabel polysilicon 114 -822 114 -822 0 3
rlabel polysilicon 121 -816 121 -816 0 1
rlabel polysilicon 121 -822 121 -822 0 3
rlabel polysilicon 128 -816 128 -816 0 1
rlabel polysilicon 128 -822 128 -822 0 3
rlabel polysilicon 135 -816 135 -816 0 1
rlabel polysilicon 135 -822 135 -822 0 3
rlabel polysilicon 142 -816 142 -816 0 1
rlabel polysilicon 142 -822 142 -822 0 3
rlabel polysilicon 149 -816 149 -816 0 1
rlabel polysilicon 149 -822 149 -822 0 3
rlabel polysilicon 152 -822 152 -822 0 4
rlabel polysilicon 156 -816 156 -816 0 1
rlabel polysilicon 156 -822 156 -822 0 3
rlabel polysilicon 163 -816 163 -816 0 1
rlabel polysilicon 163 -822 163 -822 0 3
rlabel polysilicon 170 -816 170 -816 0 1
rlabel polysilicon 170 -822 170 -822 0 3
rlabel polysilicon 177 -816 177 -816 0 1
rlabel polysilicon 177 -822 177 -822 0 3
rlabel polysilicon 187 -816 187 -816 0 2
rlabel polysilicon 187 -822 187 -822 0 4
rlabel polysilicon 191 -816 191 -816 0 1
rlabel polysilicon 191 -822 191 -822 0 3
rlabel polysilicon 198 -816 198 -816 0 1
rlabel polysilicon 198 -822 198 -822 0 3
rlabel polysilicon 205 -816 205 -816 0 1
rlabel polysilicon 212 -816 212 -816 0 1
rlabel polysilicon 212 -822 212 -822 0 3
rlabel polysilicon 219 -816 219 -816 0 1
rlabel polysilicon 219 -822 219 -822 0 3
rlabel polysilicon 226 -816 226 -816 0 1
rlabel polysilicon 226 -822 226 -822 0 3
rlabel polysilicon 233 -816 233 -816 0 1
rlabel polysilicon 233 -822 233 -822 0 3
rlabel polysilicon 240 -816 240 -816 0 1
rlabel polysilicon 240 -822 240 -822 0 3
rlabel polysilicon 247 -816 247 -816 0 1
rlabel polysilicon 247 -822 247 -822 0 3
rlabel polysilicon 254 -816 254 -816 0 1
rlabel polysilicon 254 -822 254 -822 0 3
rlabel polysilicon 261 -816 261 -816 0 1
rlabel polysilicon 261 -822 261 -822 0 3
rlabel polysilicon 268 -816 268 -816 0 1
rlabel polysilicon 271 -816 271 -816 0 2
rlabel polysilicon 268 -822 268 -822 0 3
rlabel polysilicon 275 -816 275 -816 0 1
rlabel polysilicon 275 -822 275 -822 0 3
rlabel polysilicon 282 -816 282 -816 0 1
rlabel polysilicon 282 -822 282 -822 0 3
rlabel polysilicon 289 -816 289 -816 0 1
rlabel polysilicon 289 -822 289 -822 0 3
rlabel polysilicon 296 -816 296 -816 0 1
rlabel polysilicon 296 -822 296 -822 0 3
rlabel polysilicon 306 -816 306 -816 0 2
rlabel polysilicon 303 -822 303 -822 0 3
rlabel polysilicon 306 -822 306 -822 0 4
rlabel polysilicon 310 -816 310 -816 0 1
rlabel polysilicon 310 -822 310 -822 0 3
rlabel polysilicon 317 -816 317 -816 0 1
rlabel polysilicon 317 -822 317 -822 0 3
rlabel polysilicon 324 -816 324 -816 0 1
rlabel polysilicon 324 -822 324 -822 0 3
rlabel polysilicon 331 -816 331 -816 0 1
rlabel polysilicon 331 -822 331 -822 0 3
rlabel polysilicon 338 -816 338 -816 0 1
rlabel polysilicon 341 -816 341 -816 0 2
rlabel polysilicon 338 -822 338 -822 0 3
rlabel polysilicon 345 -816 345 -816 0 1
rlabel polysilicon 348 -816 348 -816 0 2
rlabel polysilicon 345 -822 345 -822 0 3
rlabel polysilicon 348 -822 348 -822 0 4
rlabel polysilicon 352 -816 352 -816 0 1
rlabel polysilicon 352 -822 352 -822 0 3
rlabel polysilicon 359 -816 359 -816 0 1
rlabel polysilicon 359 -822 359 -822 0 3
rlabel polysilicon 366 -816 366 -816 0 1
rlabel polysilicon 369 -816 369 -816 0 2
rlabel polysilicon 366 -822 366 -822 0 3
rlabel polysilicon 369 -822 369 -822 0 4
rlabel polysilicon 373 -816 373 -816 0 1
rlabel polysilicon 373 -822 373 -822 0 3
rlabel polysilicon 380 -816 380 -816 0 1
rlabel polysilicon 383 -822 383 -822 0 4
rlabel polysilicon 387 -816 387 -816 0 1
rlabel polysilicon 390 -816 390 -816 0 2
rlabel polysilicon 387 -822 387 -822 0 3
rlabel polysilicon 390 -822 390 -822 0 4
rlabel polysilicon 394 -816 394 -816 0 1
rlabel polysilicon 394 -822 394 -822 0 3
rlabel polysilicon 404 -816 404 -816 0 2
rlabel polysilicon 404 -822 404 -822 0 4
rlabel polysilicon 408 -816 408 -816 0 1
rlabel polysilicon 408 -822 408 -822 0 3
rlabel polysilicon 415 -816 415 -816 0 1
rlabel polysilicon 415 -822 415 -822 0 3
rlabel polysilicon 422 -816 422 -816 0 1
rlabel polysilicon 422 -822 422 -822 0 3
rlabel polysilicon 429 -822 429 -822 0 3
rlabel polysilicon 436 -816 436 -816 0 1
rlabel polysilicon 439 -816 439 -816 0 2
rlabel polysilicon 436 -822 436 -822 0 3
rlabel polysilicon 446 -816 446 -816 0 2
rlabel polysilicon 443 -822 443 -822 0 3
rlabel polysilicon 453 -816 453 -816 0 2
rlabel polysilicon 453 -822 453 -822 0 4
rlabel polysilicon 457 -816 457 -816 0 1
rlabel polysilicon 457 -822 457 -822 0 3
rlabel polysilicon 464 -816 464 -816 0 1
rlabel polysilicon 464 -822 464 -822 0 3
rlabel polysilicon 471 -816 471 -816 0 1
rlabel polysilicon 471 -822 471 -822 0 3
rlabel polysilicon 478 -816 478 -816 0 1
rlabel polysilicon 478 -822 478 -822 0 3
rlabel polysilicon 485 -816 485 -816 0 1
rlabel polysilicon 485 -822 485 -822 0 3
rlabel polysilicon 492 -816 492 -816 0 1
rlabel polysilicon 492 -822 492 -822 0 3
rlabel polysilicon 499 -816 499 -816 0 1
rlabel polysilicon 499 -822 499 -822 0 3
rlabel polysilicon 506 -816 506 -816 0 1
rlabel polysilicon 506 -822 506 -822 0 3
rlabel polysilicon 513 -816 513 -816 0 1
rlabel polysilicon 513 -822 513 -822 0 3
rlabel polysilicon 520 -816 520 -816 0 1
rlabel polysilicon 520 -822 520 -822 0 3
rlabel polysilicon 527 -816 527 -816 0 1
rlabel polysilicon 527 -822 527 -822 0 3
rlabel polysilicon 534 -816 534 -816 0 1
rlabel polysilicon 534 -822 534 -822 0 3
rlabel polysilicon 541 -816 541 -816 0 1
rlabel polysilicon 541 -822 541 -822 0 3
rlabel polysilicon 548 -816 548 -816 0 1
rlabel polysilicon 548 -822 548 -822 0 3
rlabel polysilicon 555 -816 555 -816 0 1
rlabel polysilicon 555 -822 555 -822 0 3
rlabel polysilicon 562 -816 562 -816 0 1
rlabel polysilicon 562 -822 562 -822 0 3
rlabel polysilicon 569 -816 569 -816 0 1
rlabel polysilicon 569 -822 569 -822 0 3
rlabel polysilicon 576 -816 576 -816 0 1
rlabel polysilicon 576 -822 576 -822 0 3
rlabel polysilicon 583 -816 583 -816 0 1
rlabel polysilicon 583 -822 583 -822 0 3
rlabel polysilicon 590 -822 590 -822 0 3
rlabel polysilicon 597 -816 597 -816 0 1
rlabel polysilicon 597 -822 597 -822 0 3
rlabel polysilicon 604 -816 604 -816 0 1
rlabel polysilicon 604 -822 604 -822 0 3
rlabel polysilicon 611 -816 611 -816 0 1
rlabel polysilicon 611 -822 611 -822 0 3
rlabel polysilicon 618 -816 618 -816 0 1
rlabel polysilicon 618 -822 618 -822 0 3
rlabel polysilicon 625 -816 625 -816 0 1
rlabel polysilicon 625 -822 625 -822 0 3
rlabel polysilicon 632 -816 632 -816 0 1
rlabel polysilicon 632 -822 632 -822 0 3
rlabel polysilicon 635 -822 635 -822 0 4
rlabel polysilicon 639 -816 639 -816 0 1
rlabel polysilicon 639 -822 639 -822 0 3
rlabel polysilicon 646 -816 646 -816 0 1
rlabel polysilicon 646 -822 646 -822 0 3
rlabel polysilicon 653 -816 653 -816 0 1
rlabel polysilicon 653 -822 653 -822 0 3
rlabel polysilicon 660 -816 660 -816 0 1
rlabel polysilicon 660 -822 660 -822 0 3
rlabel polysilicon 667 -816 667 -816 0 1
rlabel polysilicon 667 -822 667 -822 0 3
rlabel polysilicon 674 -816 674 -816 0 1
rlabel polysilicon 674 -822 674 -822 0 3
rlabel polysilicon 681 -816 681 -816 0 1
rlabel polysilicon 681 -822 681 -822 0 3
rlabel polysilicon 688 -816 688 -816 0 1
rlabel polysilicon 688 -822 688 -822 0 3
rlabel polysilicon 695 -816 695 -816 0 1
rlabel polysilicon 695 -822 695 -822 0 3
rlabel polysilicon 702 -816 702 -816 0 1
rlabel polysilicon 702 -822 702 -822 0 3
rlabel polysilicon 709 -816 709 -816 0 1
rlabel polysilicon 709 -822 709 -822 0 3
rlabel polysilicon 716 -816 716 -816 0 1
rlabel polysilicon 716 -822 716 -822 0 3
rlabel polysilicon 723 -816 723 -816 0 1
rlabel polysilicon 723 -822 723 -822 0 3
rlabel polysilicon 730 -816 730 -816 0 1
rlabel polysilicon 730 -822 730 -822 0 3
rlabel polysilicon 737 -816 737 -816 0 1
rlabel polysilicon 737 -822 737 -822 0 3
rlabel polysilicon 744 -816 744 -816 0 1
rlabel polysilicon 744 -822 744 -822 0 3
rlabel polysilicon 751 -816 751 -816 0 1
rlabel polysilicon 751 -822 751 -822 0 3
rlabel polysilicon 758 -816 758 -816 0 1
rlabel polysilicon 758 -822 758 -822 0 3
rlabel polysilicon 765 -816 765 -816 0 1
rlabel polysilicon 765 -822 765 -822 0 3
rlabel polysilicon 772 -816 772 -816 0 1
rlabel polysilicon 772 -822 772 -822 0 3
rlabel polysilicon 779 -816 779 -816 0 1
rlabel polysilicon 779 -822 779 -822 0 3
rlabel polysilicon 786 -816 786 -816 0 1
rlabel polysilicon 786 -822 786 -822 0 3
rlabel polysilicon 793 -816 793 -816 0 1
rlabel polysilicon 793 -822 793 -822 0 3
rlabel polysilicon 9 -907 9 -907 0 3
rlabel polysilicon 16 -901 16 -901 0 1
rlabel polysilicon 16 -907 16 -907 0 3
rlabel polysilicon 26 -901 26 -901 0 2
rlabel polysilicon 23 -907 23 -907 0 3
rlabel polysilicon 30 -901 30 -901 0 1
rlabel polysilicon 30 -907 30 -907 0 3
rlabel polysilicon 37 -901 37 -901 0 1
rlabel polysilicon 40 -907 40 -907 0 4
rlabel polysilicon 44 -901 44 -901 0 1
rlabel polysilicon 44 -907 44 -907 0 3
rlabel polysilicon 51 -901 51 -901 0 1
rlabel polysilicon 54 -901 54 -901 0 2
rlabel polysilicon 58 -901 58 -901 0 1
rlabel polysilicon 58 -907 58 -907 0 3
rlabel polysilicon 65 -901 65 -901 0 1
rlabel polysilicon 65 -907 65 -907 0 3
rlabel polysilicon 72 -901 72 -901 0 1
rlabel polysilicon 72 -907 72 -907 0 3
rlabel polysilicon 79 -901 79 -901 0 1
rlabel polysilicon 79 -907 79 -907 0 3
rlabel polysilicon 86 -901 86 -901 0 1
rlabel polysilicon 86 -907 86 -907 0 3
rlabel polysilicon 93 -901 93 -901 0 1
rlabel polysilicon 93 -907 93 -907 0 3
rlabel polysilicon 100 -907 100 -907 0 3
rlabel polysilicon 103 -907 103 -907 0 4
rlabel polysilicon 107 -901 107 -901 0 1
rlabel polysilicon 107 -907 107 -907 0 3
rlabel polysilicon 114 -901 114 -901 0 1
rlabel polysilicon 117 -901 117 -901 0 2
rlabel polysilicon 117 -907 117 -907 0 4
rlabel polysilicon 121 -901 121 -901 0 1
rlabel polysilicon 121 -907 121 -907 0 3
rlabel polysilicon 128 -901 128 -901 0 1
rlabel polysilicon 128 -907 128 -907 0 3
rlabel polysilicon 135 -901 135 -901 0 1
rlabel polysilicon 135 -907 135 -907 0 3
rlabel polysilicon 142 -901 142 -901 0 1
rlabel polysilicon 145 -901 145 -901 0 2
rlabel polysilicon 145 -907 145 -907 0 4
rlabel polysilicon 149 -901 149 -901 0 1
rlabel polysilicon 149 -907 149 -907 0 3
rlabel polysilicon 156 -901 156 -901 0 1
rlabel polysilicon 156 -907 156 -907 0 3
rlabel polysilicon 163 -901 163 -901 0 1
rlabel polysilicon 163 -907 163 -907 0 3
rlabel polysilicon 170 -901 170 -901 0 1
rlabel polysilicon 173 -901 173 -901 0 2
rlabel polysilicon 173 -907 173 -907 0 4
rlabel polysilicon 177 -901 177 -901 0 1
rlabel polysilicon 180 -901 180 -901 0 2
rlabel polysilicon 180 -907 180 -907 0 4
rlabel polysilicon 184 -901 184 -901 0 1
rlabel polysilicon 184 -907 184 -907 0 3
rlabel polysilicon 191 -901 191 -901 0 1
rlabel polysilicon 191 -907 191 -907 0 3
rlabel polysilicon 198 -901 198 -901 0 1
rlabel polysilicon 198 -907 198 -907 0 3
rlabel polysilicon 205 -907 205 -907 0 3
rlabel polysilicon 212 -901 212 -901 0 1
rlabel polysilicon 212 -907 212 -907 0 3
rlabel polysilicon 219 -901 219 -901 0 1
rlabel polysilicon 219 -907 219 -907 0 3
rlabel polysilicon 226 -901 226 -901 0 1
rlabel polysilicon 226 -907 226 -907 0 3
rlabel polysilicon 233 -901 233 -901 0 1
rlabel polysilicon 233 -907 233 -907 0 3
rlabel polysilicon 240 -901 240 -901 0 1
rlabel polysilicon 240 -907 240 -907 0 3
rlabel polysilicon 247 -901 247 -901 0 1
rlabel polysilicon 247 -907 247 -907 0 3
rlabel polysilicon 257 -901 257 -901 0 2
rlabel polysilicon 254 -907 254 -907 0 3
rlabel polysilicon 257 -907 257 -907 0 4
rlabel polysilicon 261 -901 261 -901 0 1
rlabel polysilicon 261 -907 261 -907 0 3
rlabel polysilicon 268 -901 268 -901 0 1
rlabel polysilicon 268 -907 268 -907 0 3
rlabel polysilicon 275 -901 275 -901 0 1
rlabel polysilicon 275 -907 275 -907 0 3
rlabel polysilicon 278 -907 278 -907 0 4
rlabel polysilicon 285 -901 285 -901 0 2
rlabel polysilicon 285 -907 285 -907 0 4
rlabel polysilicon 289 -901 289 -901 0 1
rlabel polysilicon 299 -901 299 -901 0 2
rlabel polysilicon 299 -907 299 -907 0 4
rlabel polysilicon 306 -901 306 -901 0 2
rlabel polysilicon 306 -907 306 -907 0 4
rlabel polysilicon 310 -901 310 -901 0 1
rlabel polysilicon 310 -907 310 -907 0 3
rlabel polysilicon 317 -901 317 -901 0 1
rlabel polysilicon 317 -907 317 -907 0 3
rlabel polysilicon 324 -901 324 -901 0 1
rlabel polysilicon 324 -907 324 -907 0 3
rlabel polysilicon 331 -901 331 -901 0 1
rlabel polysilicon 331 -907 331 -907 0 3
rlabel polysilicon 341 -901 341 -901 0 2
rlabel polysilicon 345 -901 345 -901 0 1
rlabel polysilicon 345 -907 345 -907 0 3
rlabel polysilicon 352 -901 352 -901 0 1
rlabel polysilicon 352 -907 352 -907 0 3
rlabel polysilicon 359 -901 359 -901 0 1
rlabel polysilicon 362 -901 362 -901 0 2
rlabel polysilicon 362 -907 362 -907 0 4
rlabel polysilicon 366 -901 366 -901 0 1
rlabel polysilicon 366 -907 366 -907 0 3
rlabel polysilicon 373 -901 373 -901 0 1
rlabel polysilicon 373 -907 373 -907 0 3
rlabel polysilicon 380 -901 380 -901 0 1
rlabel polysilicon 380 -907 380 -907 0 3
rlabel polysilicon 387 -901 387 -901 0 1
rlabel polysilicon 387 -907 387 -907 0 3
rlabel polysilicon 394 -901 394 -901 0 1
rlabel polysilicon 394 -907 394 -907 0 3
rlabel polysilicon 404 -901 404 -901 0 2
rlabel polysilicon 401 -907 401 -907 0 3
rlabel polysilicon 404 -907 404 -907 0 4
rlabel polysilicon 411 -901 411 -901 0 2
rlabel polysilicon 411 -907 411 -907 0 4
rlabel polysilicon 415 -901 415 -901 0 1
rlabel polysilicon 415 -907 415 -907 0 3
rlabel polysilicon 422 -901 422 -901 0 1
rlabel polysilicon 422 -907 422 -907 0 3
rlabel polysilicon 429 -901 429 -901 0 1
rlabel polysilicon 429 -907 429 -907 0 3
rlabel polysilicon 436 -901 436 -901 0 1
rlabel polysilicon 436 -907 436 -907 0 3
rlabel polysilicon 443 -901 443 -901 0 1
rlabel polysilicon 443 -907 443 -907 0 3
rlabel polysilicon 450 -901 450 -901 0 1
rlabel polysilicon 453 -901 453 -901 0 2
rlabel polysilicon 450 -907 450 -907 0 3
rlabel polysilicon 457 -901 457 -901 0 1
rlabel polysilicon 457 -907 457 -907 0 3
rlabel polysilicon 464 -901 464 -901 0 1
rlabel polysilicon 464 -907 464 -907 0 3
rlabel polysilicon 471 -901 471 -901 0 1
rlabel polysilicon 471 -907 471 -907 0 3
rlabel polysilicon 478 -901 478 -901 0 1
rlabel polysilicon 478 -907 478 -907 0 3
rlabel polysilicon 485 -901 485 -901 0 1
rlabel polysilicon 485 -907 485 -907 0 3
rlabel polysilicon 492 -901 492 -901 0 1
rlabel polysilicon 492 -907 492 -907 0 3
rlabel polysilicon 499 -901 499 -901 0 1
rlabel polysilicon 499 -907 499 -907 0 3
rlabel polysilicon 506 -907 506 -907 0 3
rlabel polysilicon 509 -907 509 -907 0 4
rlabel polysilicon 513 -901 513 -901 0 1
rlabel polysilicon 513 -907 513 -907 0 3
rlabel polysilicon 520 -901 520 -901 0 1
rlabel polysilicon 520 -907 520 -907 0 3
rlabel polysilicon 530 -901 530 -901 0 2
rlabel polysilicon 527 -907 527 -907 0 3
rlabel polysilicon 534 -901 534 -901 0 1
rlabel polysilicon 537 -901 537 -901 0 2
rlabel polysilicon 537 -907 537 -907 0 4
rlabel polysilicon 541 -901 541 -901 0 1
rlabel polysilicon 541 -907 541 -907 0 3
rlabel polysilicon 555 -901 555 -901 0 1
rlabel polysilicon 555 -907 555 -907 0 3
rlabel polysilicon 562 -901 562 -901 0 1
rlabel polysilicon 562 -907 562 -907 0 3
rlabel polysilicon 569 -901 569 -901 0 1
rlabel polysilicon 569 -907 569 -907 0 3
rlabel polysilicon 576 -901 576 -901 0 1
rlabel polysilicon 576 -907 576 -907 0 3
rlabel polysilicon 583 -901 583 -901 0 1
rlabel polysilicon 583 -907 583 -907 0 3
rlabel polysilicon 590 -907 590 -907 0 3
rlabel polysilicon 597 -901 597 -901 0 1
rlabel polysilicon 597 -907 597 -907 0 3
rlabel polysilicon 604 -901 604 -901 0 1
rlabel polysilicon 604 -907 604 -907 0 3
rlabel polysilicon 618 -901 618 -901 0 1
rlabel polysilicon 618 -907 618 -907 0 3
rlabel polysilicon 625 -901 625 -901 0 1
rlabel polysilicon 625 -907 625 -907 0 3
rlabel polysilicon 632 -901 632 -901 0 1
rlabel polysilicon 635 -901 635 -901 0 2
rlabel polysilicon 632 -907 632 -907 0 3
rlabel polysilicon 639 -901 639 -901 0 1
rlabel polysilicon 639 -907 639 -907 0 3
rlabel polysilicon 646 -901 646 -901 0 1
rlabel polysilicon 646 -907 646 -907 0 3
rlabel polysilicon 653 -901 653 -901 0 1
rlabel polysilicon 653 -907 653 -907 0 3
rlabel polysilicon 660 -901 660 -901 0 1
rlabel polysilicon 660 -907 660 -907 0 3
rlabel polysilicon 667 -901 667 -901 0 1
rlabel polysilicon 667 -907 667 -907 0 3
rlabel polysilicon 674 -901 674 -901 0 1
rlabel polysilicon 674 -907 674 -907 0 3
rlabel polysilicon 681 -901 681 -901 0 1
rlabel polysilicon 681 -907 681 -907 0 3
rlabel polysilicon 688 -901 688 -901 0 1
rlabel polysilicon 688 -907 688 -907 0 3
rlabel polysilicon 695 -901 695 -901 0 1
rlabel polysilicon 695 -907 695 -907 0 3
rlabel polysilicon 702 -901 702 -901 0 1
rlabel polysilicon 702 -907 702 -907 0 3
rlabel polysilicon 709 -901 709 -901 0 1
rlabel polysilicon 709 -907 709 -907 0 3
rlabel polysilicon 737 -901 737 -901 0 1
rlabel polysilicon 737 -907 737 -907 0 3
rlabel polysilicon 758 -901 758 -901 0 1
rlabel polysilicon 758 -907 758 -907 0 3
rlabel polysilicon 2 -984 2 -984 0 1
rlabel polysilicon 2 -990 2 -990 0 3
rlabel polysilicon 9 -990 9 -990 0 3
rlabel polysilicon 16 -984 16 -984 0 1
rlabel polysilicon 16 -990 16 -990 0 3
rlabel polysilicon 26 -984 26 -984 0 2
rlabel polysilicon 26 -990 26 -990 0 4
rlabel polysilicon 30 -984 30 -984 0 1
rlabel polysilicon 30 -990 30 -990 0 3
rlabel polysilicon 37 -984 37 -984 0 1
rlabel polysilicon 37 -990 37 -990 0 3
rlabel polysilicon 44 -984 44 -984 0 1
rlabel polysilicon 47 -984 47 -984 0 2
rlabel polysilicon 44 -990 44 -990 0 3
rlabel polysilicon 47 -990 47 -990 0 4
rlabel polysilicon 51 -984 51 -984 0 1
rlabel polysilicon 54 -984 54 -984 0 2
rlabel polysilicon 58 -984 58 -984 0 1
rlabel polysilicon 61 -984 61 -984 0 2
rlabel polysilicon 65 -984 65 -984 0 1
rlabel polysilicon 68 -990 68 -990 0 4
rlabel polysilicon 72 -984 72 -984 0 1
rlabel polysilicon 72 -990 72 -990 0 3
rlabel polysilicon 79 -984 79 -984 0 1
rlabel polysilicon 79 -990 79 -990 0 3
rlabel polysilicon 86 -990 86 -990 0 3
rlabel polysilicon 89 -990 89 -990 0 4
rlabel polysilicon 93 -984 93 -984 0 1
rlabel polysilicon 93 -990 93 -990 0 3
rlabel polysilicon 100 -984 100 -984 0 1
rlabel polysilicon 100 -990 100 -990 0 3
rlabel polysilicon 107 -984 107 -984 0 1
rlabel polysilicon 107 -990 107 -990 0 3
rlabel polysilicon 114 -984 114 -984 0 1
rlabel polysilicon 114 -990 114 -990 0 3
rlabel polysilicon 121 -984 121 -984 0 1
rlabel polysilicon 121 -990 121 -990 0 3
rlabel polysilicon 128 -984 128 -984 0 1
rlabel polysilicon 128 -990 128 -990 0 3
rlabel polysilicon 135 -984 135 -984 0 1
rlabel polysilicon 135 -990 135 -990 0 3
rlabel polysilicon 142 -984 142 -984 0 1
rlabel polysilicon 145 -984 145 -984 0 2
rlabel polysilicon 142 -990 142 -990 0 3
rlabel polysilicon 149 -984 149 -984 0 1
rlabel polysilicon 152 -984 152 -984 0 2
rlabel polysilicon 149 -990 149 -990 0 3
rlabel polysilicon 156 -984 156 -984 0 1
rlabel polysilicon 156 -990 156 -990 0 3
rlabel polysilicon 163 -984 163 -984 0 1
rlabel polysilicon 163 -990 163 -990 0 3
rlabel polysilicon 170 -984 170 -984 0 1
rlabel polysilicon 170 -990 170 -990 0 3
rlabel polysilicon 180 -984 180 -984 0 2
rlabel polysilicon 177 -990 177 -990 0 3
rlabel polysilicon 180 -990 180 -990 0 4
rlabel polysilicon 184 -984 184 -984 0 1
rlabel polysilicon 187 -984 187 -984 0 2
rlabel polysilicon 184 -990 184 -990 0 3
rlabel polysilicon 187 -990 187 -990 0 4
rlabel polysilicon 191 -984 191 -984 0 1
rlabel polysilicon 191 -990 191 -990 0 3
rlabel polysilicon 198 -984 198 -984 0 1
rlabel polysilicon 198 -990 198 -990 0 3
rlabel polysilicon 205 -984 205 -984 0 1
rlabel polysilicon 205 -990 205 -990 0 3
rlabel polysilicon 212 -984 212 -984 0 1
rlabel polysilicon 212 -990 212 -990 0 3
rlabel polysilicon 219 -984 219 -984 0 1
rlabel polysilicon 219 -990 219 -990 0 3
rlabel polysilicon 229 -984 229 -984 0 2
rlabel polysilicon 226 -990 226 -990 0 3
rlabel polysilicon 233 -984 233 -984 0 1
rlabel polysilicon 233 -990 233 -990 0 3
rlabel polysilicon 240 -984 240 -984 0 1
rlabel polysilicon 240 -990 240 -990 0 3
rlabel polysilicon 250 -984 250 -984 0 2
rlabel polysilicon 250 -990 250 -990 0 4
rlabel polysilicon 254 -984 254 -984 0 1
rlabel polysilicon 254 -990 254 -990 0 3
rlabel polysilicon 261 -984 261 -984 0 1
rlabel polysilicon 261 -990 261 -990 0 3
rlabel polysilicon 268 -984 268 -984 0 1
rlabel polysilicon 268 -990 268 -990 0 3
rlabel polysilicon 275 -984 275 -984 0 1
rlabel polysilicon 275 -990 275 -990 0 3
rlabel polysilicon 282 -984 282 -984 0 1
rlabel polysilicon 282 -990 282 -990 0 3
rlabel polysilicon 289 -984 289 -984 0 1
rlabel polysilicon 292 -990 292 -990 0 4
rlabel polysilicon 296 -984 296 -984 0 1
rlabel polysilicon 296 -990 296 -990 0 3
rlabel polysilicon 303 -984 303 -984 0 1
rlabel polysilicon 303 -990 303 -990 0 3
rlabel polysilicon 310 -984 310 -984 0 1
rlabel polysilicon 313 -984 313 -984 0 2
rlabel polysilicon 310 -990 310 -990 0 3
rlabel polysilicon 313 -990 313 -990 0 4
rlabel polysilicon 317 -984 317 -984 0 1
rlabel polysilicon 317 -990 317 -990 0 3
rlabel polysilicon 324 -984 324 -984 0 1
rlabel polysilicon 324 -990 324 -990 0 3
rlabel polysilicon 331 -984 331 -984 0 1
rlabel polysilicon 331 -990 331 -990 0 3
rlabel polysilicon 338 -984 338 -984 0 1
rlabel polysilicon 338 -990 338 -990 0 3
rlabel polysilicon 345 -984 345 -984 0 1
rlabel polysilicon 345 -990 345 -990 0 3
rlabel polysilicon 352 -984 352 -984 0 1
rlabel polysilicon 352 -990 352 -990 0 3
rlabel polysilicon 359 -984 359 -984 0 1
rlabel polysilicon 362 -984 362 -984 0 2
rlabel polysilicon 366 -984 366 -984 0 1
rlabel polysilicon 366 -990 366 -990 0 3
rlabel polysilicon 373 -984 373 -984 0 1
rlabel polysilicon 373 -990 373 -990 0 3
rlabel polysilicon 383 -984 383 -984 0 2
rlabel polysilicon 383 -990 383 -990 0 4
rlabel polysilicon 387 -984 387 -984 0 1
rlabel polysilicon 387 -990 387 -990 0 3
rlabel polysilicon 394 -984 394 -984 0 1
rlabel polysilicon 397 -984 397 -984 0 2
rlabel polysilicon 394 -990 394 -990 0 3
rlabel polysilicon 397 -990 397 -990 0 4
rlabel polysilicon 401 -984 401 -984 0 1
rlabel polysilicon 401 -990 401 -990 0 3
rlabel polysilicon 408 -984 408 -984 0 1
rlabel polysilicon 411 -984 411 -984 0 2
rlabel polysilicon 411 -990 411 -990 0 4
rlabel polysilicon 415 -984 415 -984 0 1
rlabel polysilicon 415 -990 415 -990 0 3
rlabel polysilicon 422 -984 422 -984 0 1
rlabel polysilicon 422 -990 422 -990 0 3
rlabel polysilicon 429 -984 429 -984 0 1
rlabel polysilicon 429 -990 429 -990 0 3
rlabel polysilicon 436 -984 436 -984 0 1
rlabel polysilicon 436 -990 436 -990 0 3
rlabel polysilicon 443 -984 443 -984 0 1
rlabel polysilicon 446 -990 446 -990 0 4
rlabel polysilicon 450 -984 450 -984 0 1
rlabel polysilicon 450 -990 450 -990 0 3
rlabel polysilicon 457 -984 457 -984 0 1
rlabel polysilicon 457 -990 457 -990 0 3
rlabel polysilicon 464 -984 464 -984 0 1
rlabel polysilicon 464 -990 464 -990 0 3
rlabel polysilicon 471 -984 471 -984 0 1
rlabel polysilicon 471 -990 471 -990 0 3
rlabel polysilicon 478 -984 478 -984 0 1
rlabel polysilicon 478 -990 478 -990 0 3
rlabel polysilicon 485 -990 485 -990 0 3
rlabel polysilicon 488 -990 488 -990 0 4
rlabel polysilicon 492 -984 492 -984 0 1
rlabel polysilicon 492 -990 492 -990 0 3
rlabel polysilicon 499 -984 499 -984 0 1
rlabel polysilicon 502 -984 502 -984 0 2
rlabel polysilicon 502 -990 502 -990 0 4
rlabel polysilicon 506 -984 506 -984 0 1
rlabel polysilicon 506 -990 506 -990 0 3
rlabel polysilicon 513 -984 513 -984 0 1
rlabel polysilicon 513 -990 513 -990 0 3
rlabel polysilicon 520 -984 520 -984 0 1
rlabel polysilicon 520 -990 520 -990 0 3
rlabel polysilicon 527 -984 527 -984 0 1
rlabel polysilicon 527 -990 527 -990 0 3
rlabel polysilicon 534 -984 534 -984 0 1
rlabel polysilicon 534 -990 534 -990 0 3
rlabel polysilicon 541 -984 541 -984 0 1
rlabel polysilicon 541 -990 541 -990 0 3
rlabel polysilicon 548 -984 548 -984 0 1
rlabel polysilicon 548 -990 548 -990 0 3
rlabel polysilicon 555 -984 555 -984 0 1
rlabel polysilicon 555 -990 555 -990 0 3
rlabel polysilicon 562 -984 562 -984 0 1
rlabel polysilicon 562 -990 562 -990 0 3
rlabel polysilicon 569 -984 569 -984 0 1
rlabel polysilicon 569 -990 569 -990 0 3
rlabel polysilicon 576 -984 576 -984 0 1
rlabel polysilicon 576 -990 576 -990 0 3
rlabel polysilicon 583 -984 583 -984 0 1
rlabel polysilicon 583 -990 583 -990 0 3
rlabel polysilicon 590 -984 590 -984 0 1
rlabel polysilicon 590 -990 590 -990 0 3
rlabel polysilicon 604 -984 604 -984 0 1
rlabel polysilicon 607 -984 607 -984 0 2
rlabel polysilicon 604 -990 604 -990 0 3
rlabel polysilicon 607 -990 607 -990 0 4
rlabel polysilicon 611 -984 611 -984 0 1
rlabel polysilicon 611 -990 611 -990 0 3
rlabel polysilicon 621 -984 621 -984 0 2
rlabel polysilicon 621 -990 621 -990 0 4
rlabel polysilicon 625 -984 625 -984 0 1
rlabel polysilicon 625 -990 625 -990 0 3
rlabel polysilicon 632 -984 632 -984 0 1
rlabel polysilicon 632 -990 632 -990 0 3
rlabel polysilicon 639 -984 639 -984 0 1
rlabel polysilicon 639 -990 639 -990 0 3
rlabel polysilicon 646 -984 646 -984 0 1
rlabel polysilicon 646 -990 646 -990 0 3
rlabel polysilicon 653 -984 653 -984 0 1
rlabel polysilicon 653 -990 653 -990 0 3
rlabel polysilicon 660 -984 660 -984 0 1
rlabel polysilicon 660 -990 660 -990 0 3
rlabel polysilicon 667 -984 667 -984 0 1
rlabel polysilicon 667 -990 667 -990 0 3
rlabel polysilicon 674 -984 674 -984 0 1
rlabel polysilicon 674 -990 674 -990 0 3
rlabel polysilicon 681 -984 681 -984 0 1
rlabel polysilicon 681 -990 681 -990 0 3
rlabel polysilicon 688 -984 688 -984 0 1
rlabel polysilicon 688 -990 688 -990 0 3
rlabel polysilicon 695 -984 695 -984 0 1
rlabel polysilicon 695 -990 695 -990 0 3
rlabel polysilicon 702 -984 702 -984 0 1
rlabel polysilicon 702 -990 702 -990 0 3
rlabel polysilicon 709 -984 709 -984 0 1
rlabel polysilicon 709 -990 709 -990 0 3
rlabel polysilicon 716 -984 716 -984 0 1
rlabel polysilicon 716 -990 716 -990 0 3
rlabel polysilicon 726 -984 726 -984 0 2
rlabel polysilicon 751 -984 751 -984 0 1
rlabel polysilicon 751 -990 751 -990 0 3
rlabel polysilicon 9 -1065 9 -1065 0 3
rlabel polysilicon 16 -1059 16 -1059 0 1
rlabel polysilicon 16 -1065 16 -1065 0 3
rlabel polysilicon 23 -1059 23 -1059 0 1
rlabel polysilicon 26 -1065 26 -1065 0 4
rlabel polysilicon 30 -1059 30 -1059 0 1
rlabel polysilicon 30 -1065 30 -1065 0 3
rlabel polysilicon 37 -1059 37 -1059 0 1
rlabel polysilicon 37 -1065 37 -1065 0 3
rlabel polysilicon 47 -1065 47 -1065 0 4
rlabel polysilicon 54 -1059 54 -1059 0 2
rlabel polysilicon 51 -1065 51 -1065 0 3
rlabel polysilicon 58 -1059 58 -1059 0 1
rlabel polysilicon 58 -1065 58 -1065 0 3
rlabel polysilicon 65 -1059 65 -1059 0 1
rlabel polysilicon 65 -1065 65 -1065 0 3
rlabel polysilicon 75 -1059 75 -1059 0 2
rlabel polysilicon 79 -1059 79 -1059 0 1
rlabel polysilicon 79 -1065 79 -1065 0 3
rlabel polysilicon 86 -1059 86 -1059 0 1
rlabel polysilicon 86 -1065 86 -1065 0 3
rlabel polysilicon 93 -1059 93 -1059 0 1
rlabel polysilicon 93 -1065 93 -1065 0 3
rlabel polysilicon 100 -1059 100 -1059 0 1
rlabel polysilicon 103 -1059 103 -1059 0 2
rlabel polysilicon 103 -1065 103 -1065 0 4
rlabel polysilicon 107 -1059 107 -1059 0 1
rlabel polysilicon 107 -1065 107 -1065 0 3
rlabel polysilicon 117 -1059 117 -1059 0 2
rlabel polysilicon 114 -1065 114 -1065 0 3
rlabel polysilicon 121 -1059 121 -1059 0 1
rlabel polysilicon 121 -1065 121 -1065 0 3
rlabel polysilicon 128 -1059 128 -1059 0 1
rlabel polysilicon 128 -1065 128 -1065 0 3
rlabel polysilicon 135 -1059 135 -1059 0 1
rlabel polysilicon 135 -1065 135 -1065 0 3
rlabel polysilicon 138 -1065 138 -1065 0 4
rlabel polysilicon 142 -1059 142 -1059 0 1
rlabel polysilicon 142 -1065 142 -1065 0 3
rlabel polysilicon 149 -1059 149 -1059 0 1
rlabel polysilicon 149 -1065 149 -1065 0 3
rlabel polysilicon 156 -1059 156 -1059 0 1
rlabel polysilicon 156 -1065 156 -1065 0 3
rlabel polysilicon 163 -1059 163 -1059 0 1
rlabel polysilicon 163 -1065 163 -1065 0 3
rlabel polysilicon 170 -1059 170 -1059 0 1
rlabel polysilicon 173 -1065 173 -1065 0 4
rlabel polysilicon 177 -1059 177 -1059 0 1
rlabel polysilicon 177 -1065 177 -1065 0 3
rlabel polysilicon 184 -1059 184 -1059 0 1
rlabel polysilicon 184 -1065 184 -1065 0 3
rlabel polysilicon 187 -1065 187 -1065 0 4
rlabel polysilicon 191 -1059 191 -1059 0 1
rlabel polysilicon 191 -1065 191 -1065 0 3
rlabel polysilicon 198 -1059 198 -1059 0 1
rlabel polysilicon 198 -1065 198 -1065 0 3
rlabel polysilicon 205 -1059 205 -1059 0 1
rlabel polysilicon 205 -1065 205 -1065 0 3
rlabel polysilicon 212 -1059 212 -1059 0 1
rlabel polysilicon 212 -1065 212 -1065 0 3
rlabel polysilicon 219 -1059 219 -1059 0 1
rlabel polysilicon 219 -1065 219 -1065 0 3
rlabel polysilicon 226 -1059 226 -1059 0 1
rlabel polysilicon 226 -1065 226 -1065 0 3
rlabel polysilicon 233 -1059 233 -1059 0 1
rlabel polysilicon 233 -1065 233 -1065 0 3
rlabel polysilicon 240 -1059 240 -1059 0 1
rlabel polysilicon 240 -1065 240 -1065 0 3
rlabel polysilicon 247 -1059 247 -1059 0 1
rlabel polysilicon 247 -1065 247 -1065 0 3
rlabel polysilicon 254 -1059 254 -1059 0 1
rlabel polysilicon 254 -1065 254 -1065 0 3
rlabel polysilicon 261 -1059 261 -1059 0 1
rlabel polysilicon 261 -1065 261 -1065 0 3
rlabel polysilicon 268 -1059 268 -1059 0 1
rlabel polysilicon 271 -1065 271 -1065 0 4
rlabel polysilicon 275 -1059 275 -1059 0 1
rlabel polysilicon 275 -1065 275 -1065 0 3
rlabel polysilicon 282 -1065 282 -1065 0 3
rlabel polysilicon 289 -1059 289 -1059 0 1
rlabel polysilicon 289 -1065 289 -1065 0 3
rlabel polysilicon 296 -1059 296 -1059 0 1
rlabel polysilicon 296 -1065 296 -1065 0 3
rlabel polysilicon 303 -1059 303 -1059 0 1
rlabel polysilicon 306 -1059 306 -1059 0 2
rlabel polysilicon 303 -1065 303 -1065 0 3
rlabel polysilicon 306 -1065 306 -1065 0 4
rlabel polysilicon 310 -1059 310 -1059 0 1
rlabel polysilicon 310 -1065 310 -1065 0 3
rlabel polysilicon 317 -1059 317 -1059 0 1
rlabel polysilicon 320 -1059 320 -1059 0 2
rlabel polysilicon 317 -1065 317 -1065 0 3
rlabel polysilicon 324 -1059 324 -1059 0 1
rlabel polysilicon 324 -1065 324 -1065 0 3
rlabel polysilicon 331 -1059 331 -1059 0 1
rlabel polysilicon 331 -1065 331 -1065 0 3
rlabel polysilicon 338 -1059 338 -1059 0 1
rlabel polysilicon 338 -1065 338 -1065 0 3
rlabel polysilicon 345 -1059 345 -1059 0 1
rlabel polysilicon 345 -1065 345 -1065 0 3
rlabel polysilicon 352 -1059 352 -1059 0 1
rlabel polysilicon 355 -1059 355 -1059 0 2
rlabel polysilicon 359 -1059 359 -1059 0 1
rlabel polysilicon 362 -1059 362 -1059 0 2
rlabel polysilicon 362 -1065 362 -1065 0 4
rlabel polysilicon 366 -1059 366 -1059 0 1
rlabel polysilicon 369 -1059 369 -1059 0 2
rlabel polysilicon 366 -1065 366 -1065 0 3
rlabel polysilicon 373 -1059 373 -1059 0 1
rlabel polysilicon 376 -1065 376 -1065 0 4
rlabel polysilicon 380 -1059 380 -1059 0 1
rlabel polysilicon 380 -1065 380 -1065 0 3
rlabel polysilicon 387 -1059 387 -1059 0 1
rlabel polysilicon 387 -1065 387 -1065 0 3
rlabel polysilicon 394 -1059 394 -1059 0 1
rlabel polysilicon 397 -1065 397 -1065 0 4
rlabel polysilicon 401 -1059 401 -1059 0 1
rlabel polysilicon 404 -1059 404 -1059 0 2
rlabel polysilicon 408 -1059 408 -1059 0 1
rlabel polysilicon 408 -1065 408 -1065 0 3
rlabel polysilicon 415 -1065 415 -1065 0 3
rlabel polysilicon 418 -1065 418 -1065 0 4
rlabel polysilicon 422 -1059 422 -1059 0 1
rlabel polysilicon 425 -1059 425 -1059 0 2
rlabel polysilicon 425 -1065 425 -1065 0 4
rlabel polysilicon 429 -1059 429 -1059 0 1
rlabel polysilicon 429 -1065 429 -1065 0 3
rlabel polysilicon 436 -1059 436 -1059 0 1
rlabel polysilicon 436 -1065 436 -1065 0 3
rlabel polysilicon 443 -1059 443 -1059 0 1
rlabel polysilicon 443 -1065 443 -1065 0 3
rlabel polysilicon 450 -1059 450 -1059 0 1
rlabel polysilicon 450 -1065 450 -1065 0 3
rlabel polysilicon 457 -1059 457 -1059 0 1
rlabel polysilicon 457 -1065 457 -1065 0 3
rlabel polysilicon 464 -1059 464 -1059 0 1
rlabel polysilicon 464 -1065 464 -1065 0 3
rlabel polysilicon 471 -1059 471 -1059 0 1
rlabel polysilicon 471 -1065 471 -1065 0 3
rlabel polysilicon 478 -1059 478 -1059 0 1
rlabel polysilicon 478 -1065 478 -1065 0 3
rlabel polysilicon 485 -1059 485 -1059 0 1
rlabel polysilicon 485 -1065 485 -1065 0 3
rlabel polysilicon 492 -1059 492 -1059 0 1
rlabel polysilicon 492 -1065 492 -1065 0 3
rlabel polysilicon 499 -1059 499 -1059 0 1
rlabel polysilicon 499 -1065 499 -1065 0 3
rlabel polysilicon 506 -1059 506 -1059 0 1
rlabel polysilicon 506 -1065 506 -1065 0 3
rlabel polysilicon 513 -1059 513 -1059 0 1
rlabel polysilicon 513 -1065 513 -1065 0 3
rlabel polysilicon 520 -1059 520 -1059 0 1
rlabel polysilicon 520 -1065 520 -1065 0 3
rlabel polysilicon 527 -1059 527 -1059 0 1
rlabel polysilicon 527 -1065 527 -1065 0 3
rlabel polysilicon 534 -1059 534 -1059 0 1
rlabel polysilicon 534 -1065 534 -1065 0 3
rlabel polysilicon 541 -1059 541 -1059 0 1
rlabel polysilicon 541 -1065 541 -1065 0 3
rlabel polysilicon 548 -1059 548 -1059 0 1
rlabel polysilicon 548 -1065 548 -1065 0 3
rlabel polysilicon 555 -1059 555 -1059 0 1
rlabel polysilicon 555 -1065 555 -1065 0 3
rlabel polysilicon 562 -1059 562 -1059 0 1
rlabel polysilicon 562 -1065 562 -1065 0 3
rlabel polysilicon 569 -1059 569 -1059 0 1
rlabel polysilicon 569 -1065 569 -1065 0 3
rlabel polysilicon 576 -1059 576 -1059 0 1
rlabel polysilicon 576 -1065 576 -1065 0 3
rlabel polysilicon 583 -1059 583 -1059 0 1
rlabel polysilicon 583 -1065 583 -1065 0 3
rlabel polysilicon 590 -1059 590 -1059 0 1
rlabel polysilicon 590 -1065 590 -1065 0 3
rlabel polysilicon 597 -1059 597 -1059 0 1
rlabel polysilicon 597 -1065 597 -1065 0 3
rlabel polysilicon 604 -1065 604 -1065 0 3
rlabel polysilicon 611 -1059 611 -1059 0 1
rlabel polysilicon 611 -1065 611 -1065 0 3
rlabel polysilicon 618 -1059 618 -1059 0 1
rlabel polysilicon 618 -1065 618 -1065 0 3
rlabel polysilicon 625 -1059 625 -1059 0 1
rlabel polysilicon 625 -1065 625 -1065 0 3
rlabel polysilicon 632 -1059 632 -1059 0 1
rlabel polysilicon 632 -1065 632 -1065 0 3
rlabel polysilicon 639 -1059 639 -1059 0 1
rlabel polysilicon 639 -1065 639 -1065 0 3
rlabel polysilicon 646 -1059 646 -1059 0 1
rlabel polysilicon 646 -1065 646 -1065 0 3
rlabel polysilicon 653 -1059 653 -1059 0 1
rlabel polysilicon 653 -1065 653 -1065 0 3
rlabel polysilicon 660 -1059 660 -1059 0 1
rlabel polysilicon 660 -1065 660 -1065 0 3
rlabel polysilicon 667 -1059 667 -1059 0 1
rlabel polysilicon 667 -1065 667 -1065 0 3
rlabel polysilicon 674 -1059 674 -1059 0 1
rlabel polysilicon 674 -1065 674 -1065 0 3
rlabel polysilicon 681 -1059 681 -1059 0 1
rlabel polysilicon 681 -1065 681 -1065 0 3
rlabel polysilicon 688 -1059 688 -1059 0 1
rlabel polysilicon 688 -1065 688 -1065 0 3
rlabel polysilicon 695 -1059 695 -1059 0 1
rlabel polysilicon 695 -1065 695 -1065 0 3
rlabel polysilicon 702 -1059 702 -1059 0 1
rlabel polysilicon 702 -1065 702 -1065 0 3
rlabel polysilicon 709 -1059 709 -1059 0 1
rlabel polysilicon 709 -1065 709 -1065 0 3
rlabel polysilicon 716 -1059 716 -1059 0 1
rlabel polysilicon 716 -1065 716 -1065 0 3
rlabel polysilicon 723 -1059 723 -1059 0 1
rlabel polysilicon 723 -1065 723 -1065 0 3
rlabel polysilicon 730 -1059 730 -1059 0 1
rlabel polysilicon 730 -1065 730 -1065 0 3
rlabel polysilicon 754 -1065 754 -1065 0 4
rlabel polysilicon 758 -1059 758 -1059 0 1
rlabel polysilicon 758 -1065 758 -1065 0 3
rlabel polysilicon 9 -1126 9 -1126 0 1
rlabel polysilicon 9 -1132 9 -1132 0 3
rlabel polysilicon 16 -1126 16 -1126 0 1
rlabel polysilicon 16 -1132 16 -1132 0 3
rlabel polysilicon 23 -1126 23 -1126 0 1
rlabel polysilicon 26 -1132 26 -1132 0 4
rlabel polysilicon 37 -1126 37 -1126 0 1
rlabel polysilicon 37 -1132 37 -1132 0 3
rlabel polysilicon 44 -1126 44 -1126 0 1
rlabel polysilicon 44 -1132 44 -1132 0 3
rlabel polysilicon 51 -1126 51 -1126 0 1
rlabel polysilicon 51 -1132 51 -1132 0 3
rlabel polysilicon 58 -1126 58 -1126 0 1
rlabel polysilicon 58 -1132 58 -1132 0 3
rlabel polysilicon 65 -1126 65 -1126 0 1
rlabel polysilicon 65 -1132 65 -1132 0 3
rlabel polysilicon 72 -1126 72 -1126 0 1
rlabel polysilicon 72 -1132 72 -1132 0 3
rlabel polysilicon 79 -1126 79 -1126 0 1
rlabel polysilicon 79 -1132 79 -1132 0 3
rlabel polysilicon 86 -1126 86 -1126 0 1
rlabel polysilicon 89 -1126 89 -1126 0 2
rlabel polysilicon 93 -1126 93 -1126 0 1
rlabel polysilicon 93 -1132 93 -1132 0 3
rlabel polysilicon 100 -1126 100 -1126 0 1
rlabel polysilicon 100 -1132 100 -1132 0 3
rlabel polysilicon 107 -1126 107 -1126 0 1
rlabel polysilicon 107 -1132 107 -1132 0 3
rlabel polysilicon 114 -1126 114 -1126 0 1
rlabel polysilicon 117 -1126 117 -1126 0 2
rlabel polysilicon 114 -1132 114 -1132 0 3
rlabel polysilicon 117 -1132 117 -1132 0 4
rlabel polysilicon 121 -1126 121 -1126 0 1
rlabel polysilicon 121 -1132 121 -1132 0 3
rlabel polysilicon 128 -1126 128 -1126 0 1
rlabel polysilicon 128 -1132 128 -1132 0 3
rlabel polysilicon 138 -1126 138 -1126 0 2
rlabel polysilicon 135 -1132 135 -1132 0 3
rlabel polysilicon 138 -1132 138 -1132 0 4
rlabel polysilicon 142 -1126 142 -1126 0 1
rlabel polysilicon 142 -1132 142 -1132 0 3
rlabel polysilicon 149 -1126 149 -1126 0 1
rlabel polysilicon 152 -1132 152 -1132 0 4
rlabel polysilicon 156 -1126 156 -1126 0 1
rlabel polysilicon 156 -1132 156 -1132 0 3
rlabel polysilicon 163 -1126 163 -1126 0 1
rlabel polysilicon 166 -1126 166 -1126 0 2
rlabel polysilicon 163 -1132 163 -1132 0 3
rlabel polysilicon 170 -1126 170 -1126 0 1
rlabel polysilicon 170 -1132 170 -1132 0 3
rlabel polysilicon 177 -1126 177 -1126 0 1
rlabel polysilicon 180 -1126 180 -1126 0 2
rlabel polysilicon 180 -1132 180 -1132 0 4
rlabel polysilicon 184 -1126 184 -1126 0 1
rlabel polysilicon 187 -1126 187 -1126 0 2
rlabel polysilicon 187 -1132 187 -1132 0 4
rlabel polysilicon 191 -1126 191 -1126 0 1
rlabel polysilicon 194 -1126 194 -1126 0 2
rlabel polysilicon 194 -1132 194 -1132 0 4
rlabel polysilicon 198 -1126 198 -1126 0 1
rlabel polysilicon 198 -1132 198 -1132 0 3
rlabel polysilicon 205 -1126 205 -1126 0 1
rlabel polysilicon 208 -1126 208 -1126 0 2
rlabel polysilicon 208 -1132 208 -1132 0 4
rlabel polysilicon 212 -1126 212 -1126 0 1
rlabel polysilicon 212 -1132 212 -1132 0 3
rlabel polysilicon 219 -1126 219 -1126 0 1
rlabel polysilicon 219 -1132 219 -1132 0 3
rlabel polysilicon 226 -1126 226 -1126 0 1
rlabel polysilicon 226 -1132 226 -1132 0 3
rlabel polysilicon 233 -1126 233 -1126 0 1
rlabel polysilicon 233 -1132 233 -1132 0 3
rlabel polysilicon 240 -1126 240 -1126 0 1
rlabel polysilicon 240 -1132 240 -1132 0 3
rlabel polysilicon 247 -1126 247 -1126 0 1
rlabel polysilicon 250 -1126 250 -1126 0 2
rlabel polysilicon 247 -1132 247 -1132 0 3
rlabel polysilicon 250 -1132 250 -1132 0 4
rlabel polysilicon 254 -1126 254 -1126 0 1
rlabel polysilicon 254 -1132 254 -1132 0 3
rlabel polysilicon 261 -1126 261 -1126 0 1
rlabel polysilicon 261 -1132 261 -1132 0 3
rlabel polysilicon 268 -1126 268 -1126 0 1
rlabel polysilicon 268 -1132 268 -1132 0 3
rlabel polysilicon 275 -1126 275 -1126 0 1
rlabel polysilicon 275 -1132 275 -1132 0 3
rlabel polysilicon 282 -1126 282 -1126 0 1
rlabel polysilicon 282 -1132 282 -1132 0 3
rlabel polysilicon 289 -1126 289 -1126 0 1
rlabel polysilicon 292 -1132 292 -1132 0 4
rlabel polysilicon 296 -1126 296 -1126 0 1
rlabel polysilicon 296 -1132 296 -1132 0 3
rlabel polysilicon 303 -1126 303 -1126 0 1
rlabel polysilicon 303 -1132 303 -1132 0 3
rlabel polysilicon 310 -1126 310 -1126 0 1
rlabel polysilicon 310 -1132 310 -1132 0 3
rlabel polysilicon 317 -1126 317 -1126 0 1
rlabel polysilicon 320 -1126 320 -1126 0 2
rlabel polysilicon 317 -1132 317 -1132 0 3
rlabel polysilicon 324 -1126 324 -1126 0 1
rlabel polysilicon 327 -1126 327 -1126 0 2
rlabel polysilicon 324 -1132 324 -1132 0 3
rlabel polysilicon 327 -1132 327 -1132 0 4
rlabel polysilicon 331 -1126 331 -1126 0 1
rlabel polysilicon 331 -1132 331 -1132 0 3
rlabel polysilicon 338 -1126 338 -1126 0 1
rlabel polysilicon 338 -1132 338 -1132 0 3
rlabel polysilicon 345 -1126 345 -1126 0 1
rlabel polysilicon 345 -1132 345 -1132 0 3
rlabel polysilicon 352 -1132 352 -1132 0 3
rlabel polysilicon 355 -1132 355 -1132 0 4
rlabel polysilicon 359 -1126 359 -1126 0 1
rlabel polysilicon 359 -1132 359 -1132 0 3
rlabel polysilicon 366 -1126 366 -1126 0 1
rlabel polysilicon 369 -1126 369 -1126 0 2
rlabel polysilicon 366 -1132 366 -1132 0 3
rlabel polysilicon 369 -1132 369 -1132 0 4
rlabel polysilicon 373 -1126 373 -1126 0 1
rlabel polysilicon 373 -1132 373 -1132 0 3
rlabel polysilicon 380 -1126 380 -1126 0 1
rlabel polysilicon 383 -1126 383 -1126 0 2
rlabel polysilicon 380 -1132 380 -1132 0 3
rlabel polysilicon 387 -1126 387 -1126 0 1
rlabel polysilicon 387 -1132 387 -1132 0 3
rlabel polysilicon 394 -1126 394 -1126 0 1
rlabel polysilicon 394 -1132 394 -1132 0 3
rlabel polysilicon 401 -1126 401 -1126 0 1
rlabel polysilicon 401 -1132 401 -1132 0 3
rlabel polysilicon 408 -1126 408 -1126 0 1
rlabel polysilicon 408 -1132 408 -1132 0 3
rlabel polysilicon 415 -1126 415 -1126 0 1
rlabel polysilicon 415 -1132 415 -1132 0 3
rlabel polysilicon 422 -1126 422 -1126 0 1
rlabel polysilicon 425 -1126 425 -1126 0 2
rlabel polysilicon 425 -1132 425 -1132 0 4
rlabel polysilicon 429 -1126 429 -1126 0 1
rlabel polysilicon 429 -1132 429 -1132 0 3
rlabel polysilicon 432 -1132 432 -1132 0 4
rlabel polysilicon 436 -1126 436 -1126 0 1
rlabel polysilicon 439 -1126 439 -1126 0 2
rlabel polysilicon 443 -1126 443 -1126 0 1
rlabel polysilicon 443 -1132 443 -1132 0 3
rlabel polysilicon 450 -1126 450 -1126 0 1
rlabel polysilicon 450 -1132 450 -1132 0 3
rlabel polysilicon 457 -1126 457 -1126 0 1
rlabel polysilicon 457 -1132 457 -1132 0 3
rlabel polysilicon 464 -1126 464 -1126 0 1
rlabel polysilicon 464 -1132 464 -1132 0 3
rlabel polysilicon 471 -1126 471 -1126 0 1
rlabel polysilicon 474 -1126 474 -1126 0 2
rlabel polysilicon 471 -1132 471 -1132 0 3
rlabel polysilicon 474 -1132 474 -1132 0 4
rlabel polysilicon 478 -1126 478 -1126 0 1
rlabel polysilicon 478 -1132 478 -1132 0 3
rlabel polysilicon 485 -1126 485 -1126 0 1
rlabel polysilicon 485 -1132 485 -1132 0 3
rlabel polysilicon 492 -1126 492 -1126 0 1
rlabel polysilicon 492 -1132 492 -1132 0 3
rlabel polysilicon 499 -1126 499 -1126 0 1
rlabel polysilicon 499 -1132 499 -1132 0 3
rlabel polysilicon 509 -1126 509 -1126 0 2
rlabel polysilicon 509 -1132 509 -1132 0 4
rlabel polysilicon 513 -1126 513 -1126 0 1
rlabel polysilicon 513 -1132 513 -1132 0 3
rlabel polysilicon 520 -1126 520 -1126 0 1
rlabel polysilicon 520 -1132 520 -1132 0 3
rlabel polysilicon 527 -1126 527 -1126 0 1
rlabel polysilicon 527 -1132 527 -1132 0 3
rlabel polysilicon 534 -1126 534 -1126 0 1
rlabel polysilicon 534 -1132 534 -1132 0 3
rlabel polysilicon 541 -1126 541 -1126 0 1
rlabel polysilicon 541 -1132 541 -1132 0 3
rlabel polysilicon 548 -1126 548 -1126 0 1
rlabel polysilicon 548 -1132 548 -1132 0 3
rlabel polysilicon 555 -1126 555 -1126 0 1
rlabel polysilicon 555 -1132 555 -1132 0 3
rlabel polysilicon 562 -1126 562 -1126 0 1
rlabel polysilicon 562 -1132 562 -1132 0 3
rlabel polysilicon 569 -1126 569 -1126 0 1
rlabel polysilicon 569 -1132 569 -1132 0 3
rlabel polysilicon 576 -1126 576 -1126 0 1
rlabel polysilicon 576 -1132 576 -1132 0 3
rlabel polysilicon 583 -1126 583 -1126 0 1
rlabel polysilicon 583 -1132 583 -1132 0 3
rlabel polysilicon 590 -1126 590 -1126 0 1
rlabel polysilicon 590 -1132 590 -1132 0 3
rlabel polysilicon 597 -1126 597 -1126 0 1
rlabel polysilicon 597 -1132 597 -1132 0 3
rlabel polysilicon 604 -1126 604 -1126 0 1
rlabel polysilicon 604 -1132 604 -1132 0 3
rlabel polysilicon 625 -1126 625 -1126 0 1
rlabel polysilicon 625 -1132 625 -1132 0 3
rlabel polysilicon 632 -1126 632 -1126 0 1
rlabel polysilicon 632 -1132 632 -1132 0 3
rlabel polysilicon 639 -1126 639 -1126 0 1
rlabel polysilicon 639 -1132 639 -1132 0 3
rlabel polysilicon 646 -1126 646 -1126 0 1
rlabel polysilicon 646 -1132 646 -1132 0 3
rlabel polysilicon 653 -1126 653 -1126 0 1
rlabel polysilicon 653 -1132 653 -1132 0 3
rlabel polysilicon 660 -1126 660 -1126 0 1
rlabel polysilicon 660 -1132 660 -1132 0 3
rlabel polysilicon 667 -1126 667 -1126 0 1
rlabel polysilicon 667 -1132 667 -1132 0 3
rlabel polysilicon 674 -1126 674 -1126 0 1
rlabel polysilicon 674 -1132 674 -1132 0 3
rlabel polysilicon 681 -1126 681 -1126 0 1
rlabel polysilicon 681 -1132 681 -1132 0 3
rlabel polysilicon 695 -1126 695 -1126 0 1
rlabel polysilicon 695 -1132 695 -1132 0 3
rlabel polysilicon 702 -1126 702 -1126 0 1
rlabel polysilicon 702 -1132 702 -1132 0 3
rlabel polysilicon 709 -1126 709 -1126 0 1
rlabel polysilicon 709 -1132 709 -1132 0 3
rlabel polysilicon 716 -1126 716 -1126 0 1
rlabel polysilicon 716 -1132 716 -1132 0 3
rlabel polysilicon 723 -1126 723 -1126 0 1
rlabel polysilicon 723 -1132 723 -1132 0 3
rlabel polysilicon 730 -1126 730 -1126 0 1
rlabel polysilicon 730 -1132 730 -1132 0 3
rlabel polysilicon 737 -1126 737 -1126 0 1
rlabel polysilicon 740 -1126 740 -1126 0 2
rlabel polysilicon 737 -1132 737 -1132 0 3
rlabel polysilicon 740 -1132 740 -1132 0 4
rlabel polysilicon 747 -1132 747 -1132 0 4
rlabel polysilicon 751 -1126 751 -1126 0 1
rlabel polysilicon 754 -1126 754 -1126 0 2
rlabel polysilicon 751 -1132 751 -1132 0 3
rlabel polysilicon 758 -1126 758 -1126 0 1
rlabel polysilicon 758 -1132 758 -1132 0 3
rlabel polysilicon 779 -1126 779 -1126 0 1
rlabel polysilicon 779 -1132 779 -1132 0 3
rlabel polysilicon 786 -1126 786 -1126 0 1
rlabel polysilicon 786 -1132 786 -1132 0 3
rlabel polysilicon 793 -1126 793 -1126 0 1
rlabel polysilicon 793 -1132 793 -1132 0 3
rlabel polysilicon 814 -1126 814 -1126 0 1
rlabel polysilicon 814 -1132 814 -1132 0 3
rlabel polysilicon 9 -1207 9 -1207 0 1
rlabel polysilicon 9 -1213 9 -1213 0 3
rlabel polysilicon 16 -1207 16 -1207 0 1
rlabel polysilicon 16 -1213 16 -1213 0 3
rlabel polysilicon 23 -1207 23 -1207 0 1
rlabel polysilicon 23 -1213 23 -1213 0 3
rlabel polysilicon 30 -1207 30 -1207 0 1
rlabel polysilicon 33 -1207 33 -1207 0 2
rlabel polysilicon 30 -1213 30 -1213 0 3
rlabel polysilicon 33 -1213 33 -1213 0 4
rlabel polysilicon 40 -1207 40 -1207 0 2
rlabel polysilicon 44 -1207 44 -1207 0 1
rlabel polysilicon 44 -1213 44 -1213 0 3
rlabel polysilicon 51 -1207 51 -1207 0 1
rlabel polysilicon 54 -1207 54 -1207 0 2
rlabel polysilicon 51 -1213 51 -1213 0 3
rlabel polysilicon 54 -1213 54 -1213 0 4
rlabel polysilicon 58 -1207 58 -1207 0 1
rlabel polysilicon 58 -1213 58 -1213 0 3
rlabel polysilicon 65 -1207 65 -1207 0 1
rlabel polysilicon 68 -1207 68 -1207 0 2
rlabel polysilicon 68 -1213 68 -1213 0 4
rlabel polysilicon 72 -1207 72 -1207 0 1
rlabel polysilicon 72 -1213 72 -1213 0 3
rlabel polysilicon 79 -1207 79 -1207 0 1
rlabel polysilicon 79 -1213 79 -1213 0 3
rlabel polysilicon 89 -1213 89 -1213 0 4
rlabel polysilicon 93 -1207 93 -1207 0 1
rlabel polysilicon 93 -1213 93 -1213 0 3
rlabel polysilicon 100 -1207 100 -1207 0 1
rlabel polysilicon 100 -1213 100 -1213 0 3
rlabel polysilicon 107 -1207 107 -1207 0 1
rlabel polysilicon 107 -1213 107 -1213 0 3
rlabel polysilicon 117 -1207 117 -1207 0 2
rlabel polysilicon 114 -1213 114 -1213 0 3
rlabel polysilicon 121 -1207 121 -1207 0 1
rlabel polysilicon 121 -1213 121 -1213 0 3
rlabel polysilicon 128 -1207 128 -1207 0 1
rlabel polysilicon 128 -1213 128 -1213 0 3
rlabel polysilicon 135 -1207 135 -1207 0 1
rlabel polysilicon 135 -1213 135 -1213 0 3
rlabel polysilicon 145 -1207 145 -1207 0 2
rlabel polysilicon 142 -1213 142 -1213 0 3
rlabel polysilicon 145 -1213 145 -1213 0 4
rlabel polysilicon 149 -1207 149 -1207 0 1
rlabel polysilicon 149 -1213 149 -1213 0 3
rlabel polysilicon 156 -1207 156 -1207 0 1
rlabel polysilicon 156 -1213 156 -1213 0 3
rlabel polysilicon 166 -1207 166 -1207 0 2
rlabel polysilicon 170 -1207 170 -1207 0 1
rlabel polysilicon 170 -1213 170 -1213 0 3
rlabel polysilicon 177 -1207 177 -1207 0 1
rlabel polysilicon 177 -1213 177 -1213 0 3
rlabel polysilicon 187 -1207 187 -1207 0 2
rlabel polysilicon 184 -1213 184 -1213 0 3
rlabel polysilicon 191 -1207 191 -1207 0 1
rlabel polysilicon 191 -1213 191 -1213 0 3
rlabel polysilicon 198 -1207 198 -1207 0 1
rlabel polysilicon 198 -1213 198 -1213 0 3
rlabel polysilicon 205 -1207 205 -1207 0 1
rlabel polysilicon 205 -1213 205 -1213 0 3
rlabel polysilicon 212 -1207 212 -1207 0 1
rlabel polysilicon 212 -1213 212 -1213 0 3
rlabel polysilicon 219 -1207 219 -1207 0 1
rlabel polysilicon 219 -1213 219 -1213 0 3
rlabel polysilicon 226 -1207 226 -1207 0 1
rlabel polysilicon 226 -1213 226 -1213 0 3
rlabel polysilicon 236 -1207 236 -1207 0 2
rlabel polysilicon 233 -1213 233 -1213 0 3
rlabel polysilicon 240 -1207 240 -1207 0 1
rlabel polysilicon 240 -1213 240 -1213 0 3
rlabel polysilicon 247 -1207 247 -1207 0 1
rlabel polysilicon 247 -1213 247 -1213 0 3
rlabel polysilicon 257 -1207 257 -1207 0 2
rlabel polysilicon 254 -1213 254 -1213 0 3
rlabel polysilicon 261 -1207 261 -1207 0 1
rlabel polysilicon 261 -1213 261 -1213 0 3
rlabel polysilicon 268 -1207 268 -1207 0 1
rlabel polysilicon 268 -1213 268 -1213 0 3
rlabel polysilicon 275 -1207 275 -1207 0 1
rlabel polysilicon 275 -1213 275 -1213 0 3
rlabel polysilicon 278 -1213 278 -1213 0 4
rlabel polysilicon 282 -1207 282 -1207 0 1
rlabel polysilicon 282 -1213 282 -1213 0 3
rlabel polysilicon 289 -1207 289 -1207 0 1
rlabel polysilicon 289 -1213 289 -1213 0 3
rlabel polysilicon 296 -1207 296 -1207 0 1
rlabel polysilicon 296 -1213 296 -1213 0 3
rlabel polysilicon 303 -1207 303 -1207 0 1
rlabel polysilicon 303 -1213 303 -1213 0 3
rlabel polysilicon 310 -1207 310 -1207 0 1
rlabel polysilicon 310 -1213 310 -1213 0 3
rlabel polysilicon 320 -1207 320 -1207 0 2
rlabel polysilicon 317 -1213 317 -1213 0 3
rlabel polysilicon 324 -1207 324 -1207 0 1
rlabel polysilicon 324 -1213 324 -1213 0 3
rlabel polysilicon 327 -1213 327 -1213 0 4
rlabel polysilicon 331 -1207 331 -1207 0 1
rlabel polysilicon 331 -1213 331 -1213 0 3
rlabel polysilicon 338 -1207 338 -1207 0 1
rlabel polysilicon 341 -1207 341 -1207 0 2
rlabel polysilicon 341 -1213 341 -1213 0 4
rlabel polysilicon 345 -1207 345 -1207 0 1
rlabel polysilicon 348 -1207 348 -1207 0 2
rlabel polysilicon 345 -1213 345 -1213 0 3
rlabel polysilicon 348 -1213 348 -1213 0 4
rlabel polysilicon 352 -1207 352 -1207 0 1
rlabel polysilicon 352 -1213 352 -1213 0 3
rlabel polysilicon 359 -1207 359 -1207 0 1
rlabel polysilicon 359 -1213 359 -1213 0 3
rlabel polysilicon 366 -1207 366 -1207 0 1
rlabel polysilicon 369 -1207 369 -1207 0 2
rlabel polysilicon 366 -1213 366 -1213 0 3
rlabel polysilicon 373 -1207 373 -1207 0 1
rlabel polysilicon 373 -1213 373 -1213 0 3
rlabel polysilicon 380 -1207 380 -1207 0 1
rlabel polysilicon 380 -1213 380 -1213 0 3
rlabel polysilicon 390 -1207 390 -1207 0 2
rlabel polysilicon 390 -1213 390 -1213 0 4
rlabel polysilicon 394 -1207 394 -1207 0 1
rlabel polysilicon 397 -1207 397 -1207 0 2
rlabel polysilicon 397 -1213 397 -1213 0 4
rlabel polysilicon 404 -1207 404 -1207 0 2
rlabel polysilicon 401 -1213 401 -1213 0 3
rlabel polysilicon 404 -1213 404 -1213 0 4
rlabel polysilicon 411 -1207 411 -1207 0 2
rlabel polysilicon 408 -1213 408 -1213 0 3
rlabel polysilicon 411 -1213 411 -1213 0 4
rlabel polysilicon 415 -1207 415 -1207 0 1
rlabel polysilicon 415 -1213 415 -1213 0 3
rlabel polysilicon 422 -1207 422 -1207 0 1
rlabel polysilicon 422 -1213 422 -1213 0 3
rlabel polysilicon 429 -1207 429 -1207 0 1
rlabel polysilicon 429 -1213 429 -1213 0 3
rlabel polysilicon 436 -1207 436 -1207 0 1
rlabel polysilicon 436 -1213 436 -1213 0 3
rlabel polysilicon 443 -1207 443 -1207 0 1
rlabel polysilicon 443 -1213 443 -1213 0 3
rlabel polysilicon 450 -1207 450 -1207 0 1
rlabel polysilicon 450 -1213 450 -1213 0 3
rlabel polysilicon 457 -1207 457 -1207 0 1
rlabel polysilicon 457 -1213 457 -1213 0 3
rlabel polysilicon 467 -1207 467 -1207 0 2
rlabel polysilicon 464 -1213 464 -1213 0 3
rlabel polysilicon 471 -1207 471 -1207 0 1
rlabel polysilicon 474 -1213 474 -1213 0 4
rlabel polysilicon 478 -1207 478 -1207 0 1
rlabel polysilicon 478 -1213 478 -1213 0 3
rlabel polysilicon 481 -1213 481 -1213 0 4
rlabel polysilicon 485 -1207 485 -1207 0 1
rlabel polysilicon 485 -1213 485 -1213 0 3
rlabel polysilicon 492 -1207 492 -1207 0 1
rlabel polysilicon 492 -1213 492 -1213 0 3
rlabel polysilicon 499 -1207 499 -1207 0 1
rlabel polysilicon 499 -1213 499 -1213 0 3
rlabel polysilicon 506 -1207 506 -1207 0 1
rlabel polysilicon 506 -1213 506 -1213 0 3
rlabel polysilicon 513 -1207 513 -1207 0 1
rlabel polysilicon 513 -1213 513 -1213 0 3
rlabel polysilicon 520 -1207 520 -1207 0 1
rlabel polysilicon 520 -1213 520 -1213 0 3
rlabel polysilicon 527 -1207 527 -1207 0 1
rlabel polysilicon 527 -1213 527 -1213 0 3
rlabel polysilicon 534 -1207 534 -1207 0 1
rlabel polysilicon 534 -1213 534 -1213 0 3
rlabel polysilicon 541 -1213 541 -1213 0 3
rlabel polysilicon 548 -1207 548 -1207 0 1
rlabel polysilicon 548 -1213 548 -1213 0 3
rlabel polysilicon 555 -1207 555 -1207 0 1
rlabel polysilicon 555 -1213 555 -1213 0 3
rlabel polysilicon 562 -1207 562 -1207 0 1
rlabel polysilicon 562 -1213 562 -1213 0 3
rlabel polysilicon 569 -1207 569 -1207 0 1
rlabel polysilicon 569 -1213 569 -1213 0 3
rlabel polysilicon 576 -1207 576 -1207 0 1
rlabel polysilicon 576 -1213 576 -1213 0 3
rlabel polysilicon 583 -1207 583 -1207 0 1
rlabel polysilicon 583 -1213 583 -1213 0 3
rlabel polysilicon 593 -1207 593 -1207 0 2
rlabel polysilicon 593 -1213 593 -1213 0 4
rlabel polysilicon 597 -1207 597 -1207 0 1
rlabel polysilicon 597 -1213 597 -1213 0 3
rlabel polysilicon 604 -1207 604 -1207 0 1
rlabel polysilicon 604 -1213 604 -1213 0 3
rlabel polysilicon 611 -1207 611 -1207 0 1
rlabel polysilicon 611 -1213 611 -1213 0 3
rlabel polysilicon 618 -1207 618 -1207 0 1
rlabel polysilicon 618 -1213 618 -1213 0 3
rlabel polysilicon 625 -1207 625 -1207 0 1
rlabel polysilicon 625 -1213 625 -1213 0 3
rlabel polysilicon 632 -1207 632 -1207 0 1
rlabel polysilicon 632 -1213 632 -1213 0 3
rlabel polysilicon 639 -1207 639 -1207 0 1
rlabel polysilicon 639 -1213 639 -1213 0 3
rlabel polysilicon 646 -1207 646 -1207 0 1
rlabel polysilicon 646 -1213 646 -1213 0 3
rlabel polysilicon 653 -1207 653 -1207 0 1
rlabel polysilicon 653 -1213 653 -1213 0 3
rlabel polysilicon 663 -1213 663 -1213 0 4
rlabel polysilicon 667 -1207 667 -1207 0 1
rlabel polysilicon 667 -1213 667 -1213 0 3
rlabel polysilicon 674 -1207 674 -1207 0 1
rlabel polysilicon 674 -1213 674 -1213 0 3
rlabel polysilicon 681 -1207 681 -1207 0 1
rlabel polysilicon 681 -1213 681 -1213 0 3
rlabel polysilicon 688 -1207 688 -1207 0 1
rlabel polysilicon 688 -1213 688 -1213 0 3
rlabel polysilicon 695 -1207 695 -1207 0 1
rlabel polysilicon 695 -1213 695 -1213 0 3
rlabel polysilicon 702 -1207 702 -1207 0 1
rlabel polysilicon 702 -1213 702 -1213 0 3
rlabel polysilicon 709 -1207 709 -1207 0 1
rlabel polysilicon 709 -1213 709 -1213 0 3
rlabel polysilicon 716 -1207 716 -1207 0 1
rlabel polysilicon 716 -1213 716 -1213 0 3
rlabel polysilicon 723 -1207 723 -1207 0 1
rlabel polysilicon 723 -1213 723 -1213 0 3
rlabel polysilicon 730 -1207 730 -1207 0 1
rlabel polysilicon 730 -1213 730 -1213 0 3
rlabel polysilicon 744 -1207 744 -1207 0 1
rlabel polysilicon 744 -1213 744 -1213 0 3
rlabel polysilicon 751 -1207 751 -1207 0 1
rlabel polysilicon 751 -1213 751 -1213 0 3
rlabel polysilicon 758 -1207 758 -1207 0 1
rlabel polysilicon 758 -1213 758 -1213 0 3
rlabel polysilicon 765 -1207 765 -1207 0 1
rlabel polysilicon 765 -1213 765 -1213 0 3
rlabel polysilicon 772 -1207 772 -1207 0 1
rlabel polysilicon 772 -1213 772 -1213 0 3
rlabel polysilicon 779 -1207 779 -1207 0 1
rlabel polysilicon 779 -1213 779 -1213 0 3
rlabel polysilicon 786 -1207 786 -1207 0 1
rlabel polysilicon 786 -1213 786 -1213 0 3
rlabel polysilicon 793 -1207 793 -1207 0 1
rlabel polysilicon 793 -1213 793 -1213 0 3
rlabel polysilicon 800 -1207 800 -1207 0 1
rlabel polysilicon 800 -1213 800 -1213 0 3
rlabel polysilicon 2 -1300 2 -1300 0 1
rlabel polysilicon 2 -1306 2 -1306 0 3
rlabel polysilicon 9 -1300 9 -1300 0 1
rlabel polysilicon 9 -1306 9 -1306 0 3
rlabel polysilicon 16 -1300 16 -1300 0 1
rlabel polysilicon 16 -1306 16 -1306 0 3
rlabel polysilicon 23 -1300 23 -1300 0 1
rlabel polysilicon 23 -1306 23 -1306 0 3
rlabel polysilicon 30 -1300 30 -1300 0 1
rlabel polysilicon 30 -1306 30 -1306 0 3
rlabel polysilicon 37 -1300 37 -1300 0 1
rlabel polysilicon 37 -1306 37 -1306 0 3
rlabel polysilicon 44 -1300 44 -1300 0 1
rlabel polysilicon 44 -1306 44 -1306 0 3
rlabel polysilicon 51 -1300 51 -1300 0 1
rlabel polysilicon 51 -1306 51 -1306 0 3
rlabel polysilicon 58 -1300 58 -1300 0 1
rlabel polysilicon 58 -1306 58 -1306 0 3
rlabel polysilicon 65 -1300 65 -1300 0 1
rlabel polysilicon 65 -1306 65 -1306 0 3
rlabel polysilicon 68 -1306 68 -1306 0 4
rlabel polysilicon 72 -1300 72 -1300 0 1
rlabel polysilicon 75 -1300 75 -1300 0 2
rlabel polysilicon 75 -1306 75 -1306 0 4
rlabel polysilicon 79 -1300 79 -1300 0 1
rlabel polysilicon 79 -1306 79 -1306 0 3
rlabel polysilicon 86 -1300 86 -1300 0 1
rlabel polysilicon 86 -1306 86 -1306 0 3
rlabel polysilicon 93 -1300 93 -1300 0 1
rlabel polysilicon 93 -1306 93 -1306 0 3
rlabel polysilicon 100 -1300 100 -1300 0 1
rlabel polysilicon 100 -1306 100 -1306 0 3
rlabel polysilicon 107 -1300 107 -1300 0 1
rlabel polysilicon 107 -1306 107 -1306 0 3
rlabel polysilicon 114 -1306 114 -1306 0 3
rlabel polysilicon 117 -1306 117 -1306 0 4
rlabel polysilicon 121 -1300 121 -1300 0 1
rlabel polysilicon 121 -1306 121 -1306 0 3
rlabel polysilicon 128 -1300 128 -1300 0 1
rlabel polysilicon 128 -1306 128 -1306 0 3
rlabel polysilicon 135 -1300 135 -1300 0 1
rlabel polysilicon 135 -1306 135 -1306 0 3
rlabel polysilicon 145 -1300 145 -1300 0 2
rlabel polysilicon 142 -1306 142 -1306 0 3
rlabel polysilicon 149 -1300 149 -1300 0 1
rlabel polysilicon 149 -1306 149 -1306 0 3
rlabel polysilicon 156 -1300 156 -1300 0 1
rlabel polysilicon 156 -1306 156 -1306 0 3
rlabel polysilicon 166 -1300 166 -1300 0 2
rlabel polysilicon 163 -1306 163 -1306 0 3
rlabel polysilicon 166 -1306 166 -1306 0 4
rlabel polysilicon 170 -1300 170 -1300 0 1
rlabel polysilicon 170 -1306 170 -1306 0 3
rlabel polysilicon 177 -1300 177 -1300 0 1
rlabel polysilicon 177 -1306 177 -1306 0 3
rlabel polysilicon 184 -1300 184 -1300 0 1
rlabel polysilicon 187 -1300 187 -1300 0 2
rlabel polysilicon 184 -1306 184 -1306 0 3
rlabel polysilicon 187 -1306 187 -1306 0 4
rlabel polysilicon 191 -1300 191 -1300 0 1
rlabel polysilicon 191 -1306 191 -1306 0 3
rlabel polysilicon 198 -1300 198 -1300 0 1
rlabel polysilicon 198 -1306 198 -1306 0 3
rlabel polysilicon 201 -1306 201 -1306 0 4
rlabel polysilicon 205 -1300 205 -1300 0 1
rlabel polysilicon 205 -1306 205 -1306 0 3
rlabel polysilicon 212 -1300 212 -1300 0 1
rlabel polysilicon 212 -1306 212 -1306 0 3
rlabel polysilicon 219 -1300 219 -1300 0 1
rlabel polysilicon 219 -1306 219 -1306 0 3
rlabel polysilicon 229 -1306 229 -1306 0 4
rlabel polysilicon 233 -1300 233 -1300 0 1
rlabel polysilicon 233 -1306 233 -1306 0 3
rlabel polysilicon 240 -1300 240 -1300 0 1
rlabel polysilicon 240 -1306 240 -1306 0 3
rlabel polysilicon 247 -1300 247 -1300 0 1
rlabel polysilicon 247 -1306 247 -1306 0 3
rlabel polysilicon 254 -1300 254 -1300 0 1
rlabel polysilicon 254 -1306 254 -1306 0 3
rlabel polysilicon 261 -1300 261 -1300 0 1
rlabel polysilicon 261 -1306 261 -1306 0 3
rlabel polysilicon 268 -1300 268 -1300 0 1
rlabel polysilicon 268 -1306 268 -1306 0 3
rlabel polysilicon 275 -1300 275 -1300 0 1
rlabel polysilicon 275 -1306 275 -1306 0 3
rlabel polysilicon 282 -1300 282 -1300 0 1
rlabel polysilicon 282 -1306 282 -1306 0 3
rlabel polysilicon 289 -1300 289 -1300 0 1
rlabel polysilicon 289 -1306 289 -1306 0 3
rlabel polysilicon 296 -1300 296 -1300 0 1
rlabel polysilicon 296 -1306 296 -1306 0 3
rlabel polysilicon 303 -1300 303 -1300 0 1
rlabel polysilicon 303 -1306 303 -1306 0 3
rlabel polysilicon 310 -1300 310 -1300 0 1
rlabel polysilicon 313 -1306 313 -1306 0 4
rlabel polysilicon 317 -1300 317 -1300 0 1
rlabel polysilicon 317 -1306 317 -1306 0 3
rlabel polysilicon 324 -1300 324 -1300 0 1
rlabel polysilicon 324 -1306 324 -1306 0 3
rlabel polysilicon 334 -1300 334 -1300 0 2
rlabel polysilicon 334 -1306 334 -1306 0 4
rlabel polysilicon 338 -1300 338 -1300 0 1
rlabel polysilicon 341 -1300 341 -1300 0 2
rlabel polysilicon 345 -1300 345 -1300 0 1
rlabel polysilicon 345 -1306 345 -1306 0 3
rlabel polysilicon 352 -1306 352 -1306 0 3
rlabel polysilicon 355 -1306 355 -1306 0 4
rlabel polysilicon 362 -1300 362 -1300 0 2
rlabel polysilicon 359 -1306 359 -1306 0 3
rlabel polysilicon 362 -1306 362 -1306 0 4
rlabel polysilicon 366 -1306 366 -1306 0 3
rlabel polysilicon 373 -1300 373 -1300 0 1
rlabel polysilicon 373 -1306 373 -1306 0 3
rlabel polysilicon 380 -1300 380 -1300 0 1
rlabel polysilicon 380 -1306 380 -1306 0 3
rlabel polysilicon 387 -1300 387 -1300 0 1
rlabel polysilicon 387 -1306 387 -1306 0 3
rlabel polysilicon 394 -1300 394 -1300 0 1
rlabel polysilicon 394 -1306 394 -1306 0 3
rlabel polysilicon 401 -1300 401 -1300 0 1
rlabel polysilicon 404 -1300 404 -1300 0 2
rlabel polysilicon 401 -1306 401 -1306 0 3
rlabel polysilicon 408 -1300 408 -1300 0 1
rlabel polysilicon 411 -1300 411 -1300 0 2
rlabel polysilicon 408 -1306 408 -1306 0 3
rlabel polysilicon 411 -1306 411 -1306 0 4
rlabel polysilicon 415 -1300 415 -1300 0 1
rlabel polysilicon 415 -1306 415 -1306 0 3
rlabel polysilicon 422 -1300 422 -1300 0 1
rlabel polysilicon 422 -1306 422 -1306 0 3
rlabel polysilicon 425 -1306 425 -1306 0 4
rlabel polysilicon 429 -1300 429 -1300 0 1
rlabel polysilicon 429 -1306 429 -1306 0 3
rlabel polysilicon 436 -1300 436 -1300 0 1
rlabel polysilicon 436 -1306 436 -1306 0 3
rlabel polysilicon 443 -1300 443 -1300 0 1
rlabel polysilicon 443 -1306 443 -1306 0 3
rlabel polysilicon 450 -1300 450 -1300 0 1
rlabel polysilicon 450 -1306 450 -1306 0 3
rlabel polysilicon 457 -1300 457 -1300 0 1
rlabel polysilicon 457 -1306 457 -1306 0 3
rlabel polysilicon 464 -1300 464 -1300 0 1
rlabel polysilicon 464 -1306 464 -1306 0 3
rlabel polysilicon 471 -1300 471 -1300 0 1
rlabel polysilicon 471 -1306 471 -1306 0 3
rlabel polysilicon 478 -1300 478 -1300 0 1
rlabel polysilicon 478 -1306 478 -1306 0 3
rlabel polysilicon 485 -1300 485 -1300 0 1
rlabel polysilicon 485 -1306 485 -1306 0 3
rlabel polysilicon 492 -1300 492 -1300 0 1
rlabel polysilicon 492 -1306 492 -1306 0 3
rlabel polysilicon 499 -1300 499 -1300 0 1
rlabel polysilicon 499 -1306 499 -1306 0 3
rlabel polysilicon 506 -1300 506 -1300 0 1
rlabel polysilicon 506 -1306 506 -1306 0 3
rlabel polysilicon 513 -1300 513 -1300 0 1
rlabel polysilicon 513 -1306 513 -1306 0 3
rlabel polysilicon 520 -1300 520 -1300 0 1
rlabel polysilicon 520 -1306 520 -1306 0 3
rlabel polysilicon 527 -1300 527 -1300 0 1
rlabel polysilicon 527 -1306 527 -1306 0 3
rlabel polysilicon 534 -1300 534 -1300 0 1
rlabel polysilicon 534 -1306 534 -1306 0 3
rlabel polysilicon 537 -1306 537 -1306 0 4
rlabel polysilicon 541 -1300 541 -1300 0 1
rlabel polysilicon 541 -1306 541 -1306 0 3
rlabel polysilicon 548 -1300 548 -1300 0 1
rlabel polysilicon 548 -1306 548 -1306 0 3
rlabel polysilicon 555 -1300 555 -1300 0 1
rlabel polysilicon 555 -1306 555 -1306 0 3
rlabel polysilicon 562 -1300 562 -1300 0 1
rlabel polysilicon 562 -1306 562 -1306 0 3
rlabel polysilicon 572 -1300 572 -1300 0 2
rlabel polysilicon 572 -1306 572 -1306 0 4
rlabel polysilicon 576 -1300 576 -1300 0 1
rlabel polysilicon 576 -1306 576 -1306 0 3
rlabel polysilicon 583 -1300 583 -1300 0 1
rlabel polysilicon 583 -1306 583 -1306 0 3
rlabel polysilicon 590 -1300 590 -1300 0 1
rlabel polysilicon 590 -1306 590 -1306 0 3
rlabel polysilicon 597 -1300 597 -1300 0 1
rlabel polysilicon 597 -1306 597 -1306 0 3
rlabel polysilicon 604 -1300 604 -1300 0 1
rlabel polysilicon 604 -1306 604 -1306 0 3
rlabel polysilicon 611 -1300 611 -1300 0 1
rlabel polysilicon 611 -1306 611 -1306 0 3
rlabel polysilicon 618 -1300 618 -1300 0 1
rlabel polysilicon 618 -1306 618 -1306 0 3
rlabel polysilicon 625 -1300 625 -1300 0 1
rlabel polysilicon 625 -1306 625 -1306 0 3
rlabel polysilicon 632 -1300 632 -1300 0 1
rlabel polysilicon 632 -1306 632 -1306 0 3
rlabel polysilicon 639 -1300 639 -1300 0 1
rlabel polysilicon 639 -1306 639 -1306 0 3
rlabel polysilicon 646 -1300 646 -1300 0 1
rlabel polysilicon 649 -1300 649 -1300 0 2
rlabel polysilicon 653 -1300 653 -1300 0 1
rlabel polysilicon 653 -1306 653 -1306 0 3
rlabel polysilicon 660 -1300 660 -1300 0 1
rlabel polysilicon 660 -1306 660 -1306 0 3
rlabel polysilicon 667 -1300 667 -1300 0 1
rlabel polysilicon 667 -1306 667 -1306 0 3
rlabel polysilicon 674 -1300 674 -1300 0 1
rlabel polysilicon 674 -1306 674 -1306 0 3
rlabel polysilicon 681 -1300 681 -1300 0 1
rlabel polysilicon 681 -1306 681 -1306 0 3
rlabel polysilicon 688 -1300 688 -1300 0 1
rlabel polysilicon 688 -1306 688 -1306 0 3
rlabel polysilicon 695 -1300 695 -1300 0 1
rlabel polysilicon 695 -1306 695 -1306 0 3
rlabel polysilicon 702 -1300 702 -1300 0 1
rlabel polysilicon 702 -1306 702 -1306 0 3
rlabel polysilicon 709 -1300 709 -1300 0 1
rlabel polysilicon 709 -1306 709 -1306 0 3
rlabel polysilicon 716 -1300 716 -1300 0 1
rlabel polysilicon 716 -1306 716 -1306 0 3
rlabel polysilicon 723 -1300 723 -1300 0 1
rlabel polysilicon 723 -1306 723 -1306 0 3
rlabel polysilicon 730 -1300 730 -1300 0 1
rlabel polysilicon 730 -1306 730 -1306 0 3
rlabel polysilicon 737 -1300 737 -1300 0 1
rlabel polysilicon 737 -1306 737 -1306 0 3
rlabel polysilicon 744 -1300 744 -1300 0 1
rlabel polysilicon 744 -1306 744 -1306 0 3
rlabel polysilicon 751 -1300 751 -1300 0 1
rlabel polysilicon 751 -1306 751 -1306 0 3
rlabel polysilicon 758 -1300 758 -1300 0 1
rlabel polysilicon 758 -1306 758 -1306 0 3
rlabel polysilicon 768 -1306 768 -1306 0 4
rlabel polysilicon 772 -1300 772 -1300 0 1
rlabel polysilicon 779 -1300 779 -1300 0 1
rlabel polysilicon 782 -1300 782 -1300 0 2
rlabel polysilicon 782 -1306 782 -1306 0 4
rlabel polysilicon 786 -1300 786 -1300 0 1
rlabel polysilicon 789 -1300 789 -1300 0 2
rlabel polysilicon 9 -1377 9 -1377 0 1
rlabel polysilicon 23 -1377 23 -1377 0 1
rlabel polysilicon 23 -1383 23 -1383 0 3
rlabel polysilicon 30 -1377 30 -1377 0 1
rlabel polysilicon 30 -1383 30 -1383 0 3
rlabel polysilicon 40 -1377 40 -1377 0 2
rlabel polysilicon 44 -1377 44 -1377 0 1
rlabel polysilicon 44 -1383 44 -1383 0 3
rlabel polysilicon 51 -1377 51 -1377 0 1
rlabel polysilicon 51 -1383 51 -1383 0 3
rlabel polysilicon 58 -1377 58 -1377 0 1
rlabel polysilicon 58 -1383 58 -1383 0 3
rlabel polysilicon 65 -1377 65 -1377 0 1
rlabel polysilicon 65 -1383 65 -1383 0 3
rlabel polysilicon 72 -1377 72 -1377 0 1
rlabel polysilicon 75 -1383 75 -1383 0 4
rlabel polysilicon 79 -1377 79 -1377 0 1
rlabel polysilicon 82 -1377 82 -1377 0 2
rlabel polysilicon 79 -1383 79 -1383 0 3
rlabel polysilicon 89 -1383 89 -1383 0 4
rlabel polysilicon 93 -1377 93 -1377 0 1
rlabel polysilicon 93 -1383 93 -1383 0 3
rlabel polysilicon 100 -1377 100 -1377 0 1
rlabel polysilicon 100 -1383 100 -1383 0 3
rlabel polysilicon 107 -1377 107 -1377 0 1
rlabel polysilicon 107 -1383 107 -1383 0 3
rlabel polysilicon 114 -1377 114 -1377 0 1
rlabel polysilicon 117 -1377 117 -1377 0 2
rlabel polysilicon 117 -1383 117 -1383 0 4
rlabel polysilicon 121 -1377 121 -1377 0 1
rlabel polysilicon 121 -1383 121 -1383 0 3
rlabel polysilicon 128 -1377 128 -1377 0 1
rlabel polysilicon 128 -1383 128 -1383 0 3
rlabel polysilicon 135 -1377 135 -1377 0 1
rlabel polysilicon 135 -1383 135 -1383 0 3
rlabel polysilicon 142 -1377 142 -1377 0 1
rlabel polysilicon 145 -1377 145 -1377 0 2
rlabel polysilicon 142 -1383 142 -1383 0 3
rlabel polysilicon 149 -1377 149 -1377 0 1
rlabel polysilicon 149 -1383 149 -1383 0 3
rlabel polysilicon 156 -1377 156 -1377 0 1
rlabel polysilicon 156 -1383 156 -1383 0 3
rlabel polysilicon 163 -1377 163 -1377 0 1
rlabel polysilicon 163 -1383 163 -1383 0 3
rlabel polysilicon 166 -1383 166 -1383 0 4
rlabel polysilicon 170 -1377 170 -1377 0 1
rlabel polysilicon 170 -1383 170 -1383 0 3
rlabel polysilicon 177 -1377 177 -1377 0 1
rlabel polysilicon 180 -1377 180 -1377 0 2
rlabel polysilicon 177 -1383 177 -1383 0 3
rlabel polysilicon 180 -1383 180 -1383 0 4
rlabel polysilicon 184 -1377 184 -1377 0 1
rlabel polysilicon 187 -1377 187 -1377 0 2
rlabel polysilicon 184 -1383 184 -1383 0 3
rlabel polysilicon 191 -1377 191 -1377 0 1
rlabel polysilicon 191 -1383 191 -1383 0 3
rlabel polysilicon 198 -1377 198 -1377 0 1
rlabel polysilicon 198 -1383 198 -1383 0 3
rlabel polysilicon 205 -1377 205 -1377 0 1
rlabel polysilicon 205 -1383 205 -1383 0 3
rlabel polysilicon 212 -1377 212 -1377 0 1
rlabel polysilicon 215 -1377 215 -1377 0 2
rlabel polysilicon 215 -1383 215 -1383 0 4
rlabel polysilicon 219 -1377 219 -1377 0 1
rlabel polysilicon 219 -1383 219 -1383 0 3
rlabel polysilicon 226 -1377 226 -1377 0 1
rlabel polysilicon 226 -1383 226 -1383 0 3
rlabel polysilicon 233 -1377 233 -1377 0 1
rlabel polysilicon 233 -1383 233 -1383 0 3
rlabel polysilicon 240 -1377 240 -1377 0 1
rlabel polysilicon 240 -1383 240 -1383 0 3
rlabel polysilicon 247 -1377 247 -1377 0 1
rlabel polysilicon 247 -1383 247 -1383 0 3
rlabel polysilicon 254 -1377 254 -1377 0 1
rlabel polysilicon 254 -1383 254 -1383 0 3
rlabel polysilicon 261 -1377 261 -1377 0 1
rlabel polysilicon 261 -1383 261 -1383 0 3
rlabel polysilicon 268 -1377 268 -1377 0 1
rlabel polysilicon 268 -1383 268 -1383 0 3
rlabel polysilicon 275 -1377 275 -1377 0 1
rlabel polysilicon 275 -1383 275 -1383 0 3
rlabel polysilicon 278 -1383 278 -1383 0 4
rlabel polysilicon 282 -1377 282 -1377 0 1
rlabel polysilicon 282 -1383 282 -1383 0 3
rlabel polysilicon 289 -1377 289 -1377 0 1
rlabel polysilicon 289 -1383 289 -1383 0 3
rlabel polysilicon 296 -1377 296 -1377 0 1
rlabel polysilicon 296 -1383 296 -1383 0 3
rlabel polysilicon 299 -1383 299 -1383 0 4
rlabel polysilicon 303 -1377 303 -1377 0 1
rlabel polysilicon 303 -1383 303 -1383 0 3
rlabel polysilicon 310 -1377 310 -1377 0 1
rlabel polysilicon 310 -1383 310 -1383 0 3
rlabel polysilicon 317 -1377 317 -1377 0 1
rlabel polysilicon 320 -1377 320 -1377 0 2
rlabel polysilicon 317 -1383 317 -1383 0 3
rlabel polysilicon 324 -1377 324 -1377 0 1
rlabel polysilicon 324 -1383 324 -1383 0 3
rlabel polysilicon 331 -1377 331 -1377 0 1
rlabel polysilicon 334 -1377 334 -1377 0 2
rlabel polysilicon 331 -1383 331 -1383 0 3
rlabel polysilicon 338 -1377 338 -1377 0 1
rlabel polysilicon 338 -1383 338 -1383 0 3
rlabel polysilicon 348 -1377 348 -1377 0 2
rlabel polysilicon 348 -1383 348 -1383 0 4
rlabel polysilicon 352 -1377 352 -1377 0 1
rlabel polysilicon 352 -1383 352 -1383 0 3
rlabel polysilicon 359 -1377 359 -1377 0 1
rlabel polysilicon 359 -1383 359 -1383 0 3
rlabel polysilicon 366 -1377 366 -1377 0 1
rlabel polysilicon 366 -1383 366 -1383 0 3
rlabel polysilicon 373 -1377 373 -1377 0 1
rlabel polysilicon 373 -1383 373 -1383 0 3
rlabel polysilicon 380 -1377 380 -1377 0 1
rlabel polysilicon 380 -1383 380 -1383 0 3
rlabel polysilicon 387 -1377 387 -1377 0 1
rlabel polysilicon 387 -1383 387 -1383 0 3
rlabel polysilicon 394 -1377 394 -1377 0 1
rlabel polysilicon 394 -1383 394 -1383 0 3
rlabel polysilicon 401 -1377 401 -1377 0 1
rlabel polysilicon 404 -1377 404 -1377 0 2
rlabel polysilicon 404 -1383 404 -1383 0 4
rlabel polysilicon 408 -1377 408 -1377 0 1
rlabel polysilicon 408 -1383 408 -1383 0 3
rlabel polysilicon 411 -1383 411 -1383 0 4
rlabel polysilicon 415 -1377 415 -1377 0 1
rlabel polysilicon 415 -1383 415 -1383 0 3
rlabel polysilicon 422 -1377 422 -1377 0 1
rlabel polysilicon 422 -1383 422 -1383 0 3
rlabel polysilicon 429 -1377 429 -1377 0 1
rlabel polysilicon 429 -1383 429 -1383 0 3
rlabel polysilicon 436 -1377 436 -1377 0 1
rlabel polysilicon 436 -1383 436 -1383 0 3
rlabel polysilicon 443 -1377 443 -1377 0 1
rlabel polysilicon 446 -1377 446 -1377 0 2
rlabel polysilicon 443 -1383 443 -1383 0 3
rlabel polysilicon 450 -1377 450 -1377 0 1
rlabel polysilicon 450 -1383 450 -1383 0 3
rlabel polysilicon 457 -1377 457 -1377 0 1
rlabel polysilicon 457 -1383 457 -1383 0 3
rlabel polysilicon 464 -1377 464 -1377 0 1
rlabel polysilicon 464 -1383 464 -1383 0 3
rlabel polysilicon 471 -1377 471 -1377 0 1
rlabel polysilicon 471 -1383 471 -1383 0 3
rlabel polysilicon 478 -1377 478 -1377 0 1
rlabel polysilicon 481 -1377 481 -1377 0 2
rlabel polysilicon 478 -1383 478 -1383 0 3
rlabel polysilicon 485 -1377 485 -1377 0 1
rlabel polysilicon 485 -1383 485 -1383 0 3
rlabel polysilicon 492 -1377 492 -1377 0 1
rlabel polysilicon 492 -1383 492 -1383 0 3
rlabel polysilicon 499 -1377 499 -1377 0 1
rlabel polysilicon 499 -1383 499 -1383 0 3
rlabel polysilicon 506 -1377 506 -1377 0 1
rlabel polysilicon 506 -1383 506 -1383 0 3
rlabel polysilicon 513 -1377 513 -1377 0 1
rlabel polysilicon 516 -1377 516 -1377 0 2
rlabel polysilicon 513 -1383 513 -1383 0 3
rlabel polysilicon 516 -1383 516 -1383 0 4
rlabel polysilicon 520 -1377 520 -1377 0 1
rlabel polysilicon 520 -1383 520 -1383 0 3
rlabel polysilicon 527 -1377 527 -1377 0 1
rlabel polysilicon 527 -1383 527 -1383 0 3
rlabel polysilicon 534 -1377 534 -1377 0 1
rlabel polysilicon 534 -1383 534 -1383 0 3
rlabel polysilicon 541 -1377 541 -1377 0 1
rlabel polysilicon 541 -1383 541 -1383 0 3
rlabel polysilicon 548 -1377 548 -1377 0 1
rlabel polysilicon 548 -1383 548 -1383 0 3
rlabel polysilicon 555 -1377 555 -1377 0 1
rlabel polysilicon 555 -1383 555 -1383 0 3
rlabel polysilicon 562 -1377 562 -1377 0 1
rlabel polysilicon 565 -1377 565 -1377 0 2
rlabel polysilicon 565 -1383 565 -1383 0 4
rlabel polysilicon 572 -1383 572 -1383 0 4
rlabel polysilicon 576 -1377 576 -1377 0 1
rlabel polysilicon 576 -1383 576 -1383 0 3
rlabel polysilicon 583 -1377 583 -1377 0 1
rlabel polysilicon 583 -1383 583 -1383 0 3
rlabel polysilicon 590 -1377 590 -1377 0 1
rlabel polysilicon 590 -1383 590 -1383 0 3
rlabel polysilicon 597 -1377 597 -1377 0 1
rlabel polysilicon 597 -1383 597 -1383 0 3
rlabel polysilicon 604 -1377 604 -1377 0 1
rlabel polysilicon 604 -1383 604 -1383 0 3
rlabel polysilicon 611 -1377 611 -1377 0 1
rlabel polysilicon 611 -1383 611 -1383 0 3
rlabel polysilicon 618 -1377 618 -1377 0 1
rlabel polysilicon 618 -1383 618 -1383 0 3
rlabel polysilicon 632 -1377 632 -1377 0 1
rlabel polysilicon 632 -1383 632 -1383 0 3
rlabel polysilicon 639 -1377 639 -1377 0 1
rlabel polysilicon 639 -1383 639 -1383 0 3
rlabel polysilicon 646 -1377 646 -1377 0 1
rlabel polysilicon 646 -1383 646 -1383 0 3
rlabel polysilicon 653 -1377 653 -1377 0 1
rlabel polysilicon 653 -1383 653 -1383 0 3
rlabel polysilicon 660 -1377 660 -1377 0 1
rlabel polysilicon 660 -1383 660 -1383 0 3
rlabel polysilicon 667 -1377 667 -1377 0 1
rlabel polysilicon 667 -1383 667 -1383 0 3
rlabel polysilicon 674 -1377 674 -1377 0 1
rlabel polysilicon 674 -1383 674 -1383 0 3
rlabel polysilicon 681 -1377 681 -1377 0 1
rlabel polysilicon 681 -1383 681 -1383 0 3
rlabel polysilicon 688 -1377 688 -1377 0 1
rlabel polysilicon 691 -1377 691 -1377 0 2
rlabel polysilicon 688 -1383 688 -1383 0 3
rlabel polysilicon 691 -1383 691 -1383 0 4
rlabel polysilicon 695 -1377 695 -1377 0 1
rlabel polysilicon 695 -1383 695 -1383 0 3
rlabel polysilicon 702 -1377 702 -1377 0 1
rlabel polysilicon 705 -1377 705 -1377 0 2
rlabel polysilicon 705 -1383 705 -1383 0 4
rlabel polysilicon 709 -1377 709 -1377 0 1
rlabel polysilicon 709 -1383 709 -1383 0 3
rlabel polysilicon 716 -1383 716 -1383 0 3
rlabel polysilicon 758 -1377 758 -1377 0 1
rlabel polysilicon 758 -1383 758 -1383 0 3
rlabel polysilicon 779 -1377 779 -1377 0 1
rlabel polysilicon 779 -1383 779 -1383 0 3
rlabel polysilicon 800 -1377 800 -1377 0 1
rlabel polysilicon 800 -1383 800 -1383 0 3
rlabel polysilicon 9 -1446 9 -1446 0 1
rlabel polysilicon 9 -1452 9 -1452 0 3
rlabel polysilicon 16 -1446 16 -1446 0 1
rlabel polysilicon 16 -1452 16 -1452 0 3
rlabel polysilicon 23 -1446 23 -1446 0 1
rlabel polysilicon 23 -1452 23 -1452 0 3
rlabel polysilicon 30 -1446 30 -1446 0 1
rlabel polysilicon 30 -1452 30 -1452 0 3
rlabel polysilicon 37 -1446 37 -1446 0 1
rlabel polysilicon 37 -1452 37 -1452 0 3
rlabel polysilicon 44 -1446 44 -1446 0 1
rlabel polysilicon 44 -1452 44 -1452 0 3
rlabel polysilicon 51 -1446 51 -1446 0 1
rlabel polysilicon 58 -1446 58 -1446 0 1
rlabel polysilicon 58 -1452 58 -1452 0 3
rlabel polysilicon 65 -1446 65 -1446 0 1
rlabel polysilicon 65 -1452 65 -1452 0 3
rlabel polysilicon 75 -1446 75 -1446 0 2
rlabel polysilicon 79 -1446 79 -1446 0 1
rlabel polysilicon 79 -1452 79 -1452 0 3
rlabel polysilicon 86 -1446 86 -1446 0 1
rlabel polysilicon 86 -1452 86 -1452 0 3
rlabel polysilicon 93 -1446 93 -1446 0 1
rlabel polysilicon 93 -1452 93 -1452 0 3
rlabel polysilicon 100 -1446 100 -1446 0 1
rlabel polysilicon 107 -1446 107 -1446 0 1
rlabel polysilicon 107 -1452 107 -1452 0 3
rlabel polysilicon 117 -1446 117 -1446 0 2
rlabel polysilicon 117 -1452 117 -1452 0 4
rlabel polysilicon 121 -1452 121 -1452 0 3
rlabel polysilicon 124 -1452 124 -1452 0 4
rlabel polysilicon 128 -1446 128 -1446 0 1
rlabel polysilicon 128 -1452 128 -1452 0 3
rlabel polysilicon 138 -1446 138 -1446 0 2
rlabel polysilicon 135 -1452 135 -1452 0 3
rlabel polysilicon 138 -1452 138 -1452 0 4
rlabel polysilicon 142 -1446 142 -1446 0 1
rlabel polysilicon 142 -1452 142 -1452 0 3
rlabel polysilicon 149 -1446 149 -1446 0 1
rlabel polysilicon 149 -1452 149 -1452 0 3
rlabel polysilicon 156 -1452 156 -1452 0 3
rlabel polysilicon 159 -1452 159 -1452 0 4
rlabel polysilicon 163 -1446 163 -1446 0 1
rlabel polysilicon 163 -1452 163 -1452 0 3
rlabel polysilicon 170 -1446 170 -1446 0 1
rlabel polysilicon 170 -1452 170 -1452 0 3
rlabel polysilicon 177 -1446 177 -1446 0 1
rlabel polysilicon 177 -1452 177 -1452 0 3
rlabel polysilicon 184 -1452 184 -1452 0 3
rlabel polysilicon 187 -1452 187 -1452 0 4
rlabel polysilicon 191 -1446 191 -1446 0 1
rlabel polysilicon 191 -1452 191 -1452 0 3
rlabel polysilicon 198 -1446 198 -1446 0 1
rlabel polysilicon 198 -1452 198 -1452 0 3
rlabel polysilicon 205 -1446 205 -1446 0 1
rlabel polysilicon 205 -1452 205 -1452 0 3
rlabel polysilicon 212 -1446 212 -1446 0 1
rlabel polysilicon 212 -1452 212 -1452 0 3
rlabel polysilicon 219 -1446 219 -1446 0 1
rlabel polysilicon 219 -1452 219 -1452 0 3
rlabel polysilicon 226 -1446 226 -1446 0 1
rlabel polysilicon 226 -1452 226 -1452 0 3
rlabel polysilicon 233 -1446 233 -1446 0 1
rlabel polysilicon 233 -1452 233 -1452 0 3
rlabel polysilicon 240 -1446 240 -1446 0 1
rlabel polysilicon 240 -1452 240 -1452 0 3
rlabel polysilicon 247 -1446 247 -1446 0 1
rlabel polysilicon 247 -1452 247 -1452 0 3
rlabel polysilicon 254 -1446 254 -1446 0 1
rlabel polysilicon 254 -1452 254 -1452 0 3
rlabel polysilicon 261 -1446 261 -1446 0 1
rlabel polysilicon 261 -1452 261 -1452 0 3
rlabel polysilicon 268 -1446 268 -1446 0 1
rlabel polysilicon 271 -1446 271 -1446 0 2
rlabel polysilicon 271 -1452 271 -1452 0 4
rlabel polysilicon 275 -1446 275 -1446 0 1
rlabel polysilicon 275 -1452 275 -1452 0 3
rlabel polysilicon 282 -1446 282 -1446 0 1
rlabel polysilicon 282 -1452 282 -1452 0 3
rlabel polysilicon 289 -1446 289 -1446 0 1
rlabel polysilicon 289 -1452 289 -1452 0 3
rlabel polysilicon 296 -1446 296 -1446 0 1
rlabel polysilicon 296 -1452 296 -1452 0 3
rlabel polysilicon 303 -1446 303 -1446 0 1
rlabel polysilicon 303 -1452 303 -1452 0 3
rlabel polysilicon 310 -1446 310 -1446 0 1
rlabel polysilicon 310 -1452 310 -1452 0 3
rlabel polysilicon 317 -1446 317 -1446 0 1
rlabel polysilicon 317 -1452 317 -1452 0 3
rlabel polysilicon 324 -1446 324 -1446 0 1
rlabel polysilicon 324 -1452 324 -1452 0 3
rlabel polysilicon 334 -1446 334 -1446 0 2
rlabel polysilicon 331 -1452 331 -1452 0 3
rlabel polysilicon 334 -1452 334 -1452 0 4
rlabel polysilicon 338 -1446 338 -1446 0 1
rlabel polysilicon 338 -1452 338 -1452 0 3
rlabel polysilicon 345 -1446 345 -1446 0 1
rlabel polysilicon 345 -1452 345 -1452 0 3
rlabel polysilicon 352 -1446 352 -1446 0 1
rlabel polysilicon 352 -1452 352 -1452 0 3
rlabel polysilicon 359 -1446 359 -1446 0 1
rlabel polysilicon 359 -1452 359 -1452 0 3
rlabel polysilicon 366 -1446 366 -1446 0 1
rlabel polysilicon 366 -1452 366 -1452 0 3
rlabel polysilicon 373 -1446 373 -1446 0 1
rlabel polysilicon 373 -1452 373 -1452 0 3
rlabel polysilicon 380 -1446 380 -1446 0 1
rlabel polysilicon 383 -1446 383 -1446 0 2
rlabel polysilicon 380 -1452 380 -1452 0 3
rlabel polysilicon 383 -1452 383 -1452 0 4
rlabel polysilicon 387 -1446 387 -1446 0 1
rlabel polysilicon 387 -1452 387 -1452 0 3
rlabel polysilicon 394 -1446 394 -1446 0 1
rlabel polysilicon 397 -1452 397 -1452 0 4
rlabel polysilicon 404 -1446 404 -1446 0 2
rlabel polysilicon 401 -1452 401 -1452 0 3
rlabel polysilicon 404 -1452 404 -1452 0 4
rlabel polysilicon 411 -1446 411 -1446 0 2
rlabel polysilicon 415 -1446 415 -1446 0 1
rlabel polysilicon 415 -1452 415 -1452 0 3
rlabel polysilicon 422 -1446 422 -1446 0 1
rlabel polysilicon 422 -1452 422 -1452 0 3
rlabel polysilicon 429 -1446 429 -1446 0 1
rlabel polysilicon 432 -1446 432 -1446 0 2
rlabel polysilicon 429 -1452 429 -1452 0 3
rlabel polysilicon 432 -1452 432 -1452 0 4
rlabel polysilicon 439 -1446 439 -1446 0 2
rlabel polysilicon 439 -1452 439 -1452 0 4
rlabel polysilicon 443 -1446 443 -1446 0 1
rlabel polysilicon 443 -1452 443 -1452 0 3
rlabel polysilicon 450 -1446 450 -1446 0 1
rlabel polysilicon 450 -1452 450 -1452 0 3
rlabel polysilicon 457 -1446 457 -1446 0 1
rlabel polysilicon 457 -1452 457 -1452 0 3
rlabel polysilicon 464 -1446 464 -1446 0 1
rlabel polysilicon 464 -1452 464 -1452 0 3
rlabel polysilicon 471 -1452 471 -1452 0 3
rlabel polysilicon 474 -1452 474 -1452 0 4
rlabel polysilicon 478 -1446 478 -1446 0 1
rlabel polysilicon 478 -1452 478 -1452 0 3
rlabel polysilicon 485 -1446 485 -1446 0 1
rlabel polysilicon 488 -1446 488 -1446 0 2
rlabel polysilicon 492 -1446 492 -1446 0 1
rlabel polysilicon 492 -1452 492 -1452 0 3
rlabel polysilicon 499 -1446 499 -1446 0 1
rlabel polysilicon 499 -1452 499 -1452 0 3
rlabel polysilicon 506 -1446 506 -1446 0 1
rlabel polysilicon 509 -1446 509 -1446 0 2
rlabel polysilicon 509 -1452 509 -1452 0 4
rlabel polysilicon 513 -1446 513 -1446 0 1
rlabel polysilicon 513 -1452 513 -1452 0 3
rlabel polysilicon 520 -1446 520 -1446 0 1
rlabel polysilicon 520 -1452 520 -1452 0 3
rlabel polysilicon 527 -1446 527 -1446 0 1
rlabel polysilicon 527 -1452 527 -1452 0 3
rlabel polysilicon 534 -1446 534 -1446 0 1
rlabel polysilicon 534 -1452 534 -1452 0 3
rlabel polysilicon 537 -1452 537 -1452 0 4
rlabel polysilicon 541 -1446 541 -1446 0 1
rlabel polysilicon 541 -1452 541 -1452 0 3
rlabel polysilicon 548 -1446 548 -1446 0 1
rlabel polysilicon 551 -1446 551 -1446 0 2
rlabel polysilicon 555 -1446 555 -1446 0 1
rlabel polysilicon 555 -1452 555 -1452 0 3
rlabel polysilicon 562 -1446 562 -1446 0 1
rlabel polysilicon 562 -1452 562 -1452 0 3
rlabel polysilicon 569 -1446 569 -1446 0 1
rlabel polysilicon 569 -1452 569 -1452 0 3
rlabel polysilicon 576 -1446 576 -1446 0 1
rlabel polysilicon 576 -1452 576 -1452 0 3
rlabel polysilicon 583 -1446 583 -1446 0 1
rlabel polysilicon 583 -1452 583 -1452 0 3
rlabel polysilicon 590 -1446 590 -1446 0 1
rlabel polysilicon 590 -1452 590 -1452 0 3
rlabel polysilicon 597 -1446 597 -1446 0 1
rlabel polysilicon 597 -1452 597 -1452 0 3
rlabel polysilicon 604 -1446 604 -1446 0 1
rlabel polysilicon 604 -1452 604 -1452 0 3
rlabel polysilicon 611 -1446 611 -1446 0 1
rlabel polysilicon 611 -1452 611 -1452 0 3
rlabel polysilicon 618 -1446 618 -1446 0 1
rlabel polysilicon 618 -1452 618 -1452 0 3
rlabel polysilicon 625 -1446 625 -1446 0 1
rlabel polysilicon 625 -1452 625 -1452 0 3
rlabel polysilicon 632 -1446 632 -1446 0 1
rlabel polysilicon 632 -1452 632 -1452 0 3
rlabel polysilicon 639 -1446 639 -1446 0 1
rlabel polysilicon 639 -1452 639 -1452 0 3
rlabel polysilicon 646 -1446 646 -1446 0 1
rlabel polysilicon 646 -1452 646 -1452 0 3
rlabel polysilicon 653 -1446 653 -1446 0 1
rlabel polysilicon 653 -1452 653 -1452 0 3
rlabel polysilicon 660 -1446 660 -1446 0 1
rlabel polysilicon 660 -1452 660 -1452 0 3
rlabel polysilicon 667 -1446 667 -1446 0 1
rlabel polysilicon 667 -1452 667 -1452 0 3
rlabel polysilicon 674 -1446 674 -1446 0 1
rlabel polysilicon 674 -1452 674 -1452 0 3
rlabel polysilicon 681 -1446 681 -1446 0 1
rlabel polysilicon 681 -1452 681 -1452 0 3
rlabel polysilicon 688 -1446 688 -1446 0 1
rlabel polysilicon 688 -1452 688 -1452 0 3
rlabel polysilicon 695 -1446 695 -1446 0 1
rlabel polysilicon 695 -1452 695 -1452 0 3
rlabel polysilicon 702 -1446 702 -1446 0 1
rlabel polysilicon 702 -1452 702 -1452 0 3
rlabel polysilicon 709 -1446 709 -1446 0 1
rlabel polysilicon 709 -1452 709 -1452 0 3
rlabel polysilicon 716 -1446 716 -1446 0 1
rlabel polysilicon 716 -1452 716 -1452 0 3
rlabel polysilicon 723 -1446 723 -1446 0 1
rlabel polysilicon 723 -1452 723 -1452 0 3
rlabel polysilicon 730 -1446 730 -1446 0 1
rlabel polysilicon 730 -1452 730 -1452 0 3
rlabel polysilicon 737 -1446 737 -1446 0 1
rlabel polysilicon 737 -1452 737 -1452 0 3
rlabel polysilicon 744 -1446 744 -1446 0 1
rlabel polysilicon 744 -1452 744 -1452 0 3
rlabel polysilicon 751 -1446 751 -1446 0 1
rlabel polysilicon 751 -1452 751 -1452 0 3
rlabel polysilicon 765 -1446 765 -1446 0 1
rlabel polysilicon 768 -1446 768 -1446 0 2
rlabel polysilicon 768 -1452 768 -1452 0 4
rlabel polysilicon 772 -1446 772 -1446 0 1
rlabel polysilicon 772 -1452 772 -1452 0 3
rlabel polysilicon 782 -1446 782 -1446 0 2
rlabel polysilicon 779 -1452 779 -1452 0 3
rlabel polysilicon 786 -1446 786 -1446 0 1
rlabel polysilicon 789 -1446 789 -1446 0 2
rlabel polysilicon 789 -1452 789 -1452 0 4
rlabel polysilicon 796 -1446 796 -1446 0 2
rlabel polysilicon 803 -1446 803 -1446 0 2
rlabel polysilicon 800 -1452 800 -1452 0 3
rlabel polysilicon 807 -1446 807 -1446 0 1
rlabel polysilicon 807 -1452 807 -1452 0 3
rlabel polysilicon 814 -1452 814 -1452 0 3
rlabel polysilicon 817 -1452 817 -1452 0 4
rlabel polysilicon 828 -1446 828 -1446 0 1
rlabel polysilicon 828 -1452 828 -1452 0 3
rlabel polysilicon 835 -1446 835 -1446 0 1
rlabel polysilicon 835 -1452 835 -1452 0 3
rlabel polysilicon 2 -1531 2 -1531 0 3
rlabel polysilicon 9 -1525 9 -1525 0 1
rlabel polysilicon 9 -1531 9 -1531 0 3
rlabel polysilicon 16 -1525 16 -1525 0 1
rlabel polysilicon 16 -1531 16 -1531 0 3
rlabel polysilicon 23 -1525 23 -1525 0 1
rlabel polysilicon 23 -1531 23 -1531 0 3
rlabel polysilicon 30 -1525 30 -1525 0 1
rlabel polysilicon 30 -1531 30 -1531 0 3
rlabel polysilicon 37 -1525 37 -1525 0 1
rlabel polysilicon 37 -1531 37 -1531 0 3
rlabel polysilicon 44 -1525 44 -1525 0 1
rlabel polysilicon 44 -1531 44 -1531 0 3
rlabel polysilicon 54 -1525 54 -1525 0 2
rlabel polysilicon 51 -1531 51 -1531 0 3
rlabel polysilicon 58 -1525 58 -1525 0 1
rlabel polysilicon 58 -1531 58 -1531 0 3
rlabel polysilicon 65 -1525 65 -1525 0 1
rlabel polysilicon 65 -1531 65 -1531 0 3
rlabel polysilicon 72 -1525 72 -1525 0 1
rlabel polysilicon 79 -1525 79 -1525 0 1
rlabel polysilicon 79 -1531 79 -1531 0 3
rlabel polysilicon 86 -1525 86 -1525 0 1
rlabel polysilicon 86 -1531 86 -1531 0 3
rlabel polysilicon 96 -1525 96 -1525 0 2
rlabel polysilicon 96 -1531 96 -1531 0 4
rlabel polysilicon 100 -1531 100 -1531 0 3
rlabel polysilicon 107 -1525 107 -1525 0 1
rlabel polysilicon 107 -1531 107 -1531 0 3
rlabel polysilicon 114 -1525 114 -1525 0 1
rlabel polysilicon 114 -1531 114 -1531 0 3
rlabel polysilicon 121 -1525 121 -1525 0 1
rlabel polysilicon 121 -1531 121 -1531 0 3
rlabel polysilicon 128 -1525 128 -1525 0 1
rlabel polysilicon 128 -1531 128 -1531 0 3
rlabel polysilicon 138 -1525 138 -1525 0 2
rlabel polysilicon 138 -1531 138 -1531 0 4
rlabel polysilicon 142 -1525 142 -1525 0 1
rlabel polysilicon 142 -1531 142 -1531 0 3
rlabel polysilicon 149 -1525 149 -1525 0 1
rlabel polysilicon 149 -1531 149 -1531 0 3
rlabel polysilicon 156 -1525 156 -1525 0 1
rlabel polysilicon 156 -1531 156 -1531 0 3
rlabel polysilicon 166 -1525 166 -1525 0 2
rlabel polysilicon 170 -1525 170 -1525 0 1
rlabel polysilicon 170 -1531 170 -1531 0 3
rlabel polysilicon 177 -1525 177 -1525 0 1
rlabel polysilicon 180 -1525 180 -1525 0 2
rlabel polysilicon 177 -1531 177 -1531 0 3
rlabel polysilicon 184 -1531 184 -1531 0 3
rlabel polysilicon 187 -1531 187 -1531 0 4
rlabel polysilicon 191 -1525 191 -1525 0 1
rlabel polysilicon 191 -1531 191 -1531 0 3
rlabel polysilicon 198 -1525 198 -1525 0 1
rlabel polysilicon 198 -1531 198 -1531 0 3
rlabel polysilicon 205 -1531 205 -1531 0 3
rlabel polysilicon 208 -1531 208 -1531 0 4
rlabel polysilicon 212 -1525 212 -1525 0 1
rlabel polysilicon 212 -1531 212 -1531 0 3
rlabel polysilicon 219 -1525 219 -1525 0 1
rlabel polysilicon 219 -1531 219 -1531 0 3
rlabel polysilicon 226 -1525 226 -1525 0 1
rlabel polysilicon 226 -1531 226 -1531 0 3
rlabel polysilicon 233 -1525 233 -1525 0 1
rlabel polysilicon 240 -1525 240 -1525 0 1
rlabel polysilicon 247 -1525 247 -1525 0 1
rlabel polysilicon 250 -1525 250 -1525 0 2
rlabel polysilicon 247 -1531 247 -1531 0 3
rlabel polysilicon 250 -1531 250 -1531 0 4
rlabel polysilicon 257 -1525 257 -1525 0 2
rlabel polysilicon 257 -1531 257 -1531 0 4
rlabel polysilicon 261 -1525 261 -1525 0 1
rlabel polysilicon 261 -1531 261 -1531 0 3
rlabel polysilicon 268 -1525 268 -1525 0 1
rlabel polysilicon 275 -1525 275 -1525 0 1
rlabel polysilicon 275 -1531 275 -1531 0 3
rlabel polysilicon 282 -1525 282 -1525 0 1
rlabel polysilicon 282 -1531 282 -1531 0 3
rlabel polysilicon 289 -1525 289 -1525 0 1
rlabel polysilicon 289 -1531 289 -1531 0 3
rlabel polysilicon 296 -1525 296 -1525 0 1
rlabel polysilicon 296 -1531 296 -1531 0 3
rlabel polysilicon 306 -1525 306 -1525 0 2
rlabel polysilicon 303 -1531 303 -1531 0 3
rlabel polysilicon 306 -1531 306 -1531 0 4
rlabel polysilicon 310 -1525 310 -1525 0 1
rlabel polysilicon 310 -1531 310 -1531 0 3
rlabel polysilicon 317 -1525 317 -1525 0 1
rlabel polysilicon 317 -1531 317 -1531 0 3
rlabel polysilicon 324 -1525 324 -1525 0 1
rlabel polysilicon 324 -1531 324 -1531 0 3
rlabel polysilicon 331 -1525 331 -1525 0 1
rlabel polysilicon 331 -1531 331 -1531 0 3
rlabel polysilicon 334 -1531 334 -1531 0 4
rlabel polysilicon 338 -1525 338 -1525 0 1
rlabel polysilicon 341 -1525 341 -1525 0 2
rlabel polysilicon 338 -1531 338 -1531 0 3
rlabel polysilicon 341 -1531 341 -1531 0 4
rlabel polysilicon 345 -1525 345 -1525 0 1
rlabel polysilicon 345 -1531 345 -1531 0 3
rlabel polysilicon 352 -1525 352 -1525 0 1
rlabel polysilicon 352 -1531 352 -1531 0 3
rlabel polysilicon 359 -1525 359 -1525 0 1
rlabel polysilicon 362 -1525 362 -1525 0 2
rlabel polysilicon 362 -1531 362 -1531 0 4
rlabel polysilicon 366 -1525 366 -1525 0 1
rlabel polysilicon 369 -1525 369 -1525 0 2
rlabel polysilicon 373 -1525 373 -1525 0 1
rlabel polysilicon 373 -1531 373 -1531 0 3
rlabel polysilicon 380 -1525 380 -1525 0 1
rlabel polysilicon 383 -1525 383 -1525 0 2
rlabel polysilicon 380 -1531 380 -1531 0 3
rlabel polysilicon 387 -1525 387 -1525 0 1
rlabel polysilicon 390 -1525 390 -1525 0 2
rlabel polysilicon 387 -1531 387 -1531 0 3
rlabel polysilicon 394 -1525 394 -1525 0 1
rlabel polysilicon 394 -1531 394 -1531 0 3
rlabel polysilicon 401 -1525 401 -1525 0 1
rlabel polysilicon 401 -1531 401 -1531 0 3
rlabel polysilicon 408 -1525 408 -1525 0 1
rlabel polysilicon 408 -1531 408 -1531 0 3
rlabel polysilicon 415 -1525 415 -1525 0 1
rlabel polysilicon 418 -1525 418 -1525 0 2
rlabel polysilicon 415 -1531 415 -1531 0 3
rlabel polysilicon 418 -1531 418 -1531 0 4
rlabel polysilicon 422 -1525 422 -1525 0 1
rlabel polysilicon 422 -1531 422 -1531 0 3
rlabel polysilicon 429 -1525 429 -1525 0 1
rlabel polysilicon 429 -1531 429 -1531 0 3
rlabel polysilicon 436 -1525 436 -1525 0 1
rlabel polysilicon 439 -1525 439 -1525 0 2
rlabel polysilicon 439 -1531 439 -1531 0 4
rlabel polysilicon 443 -1525 443 -1525 0 1
rlabel polysilicon 443 -1531 443 -1531 0 3
rlabel polysilicon 450 -1525 450 -1525 0 1
rlabel polysilicon 450 -1531 450 -1531 0 3
rlabel polysilicon 457 -1525 457 -1525 0 1
rlabel polysilicon 457 -1531 457 -1531 0 3
rlabel polysilicon 464 -1525 464 -1525 0 1
rlabel polysilicon 464 -1531 464 -1531 0 3
rlabel polysilicon 471 -1525 471 -1525 0 1
rlabel polysilicon 471 -1531 471 -1531 0 3
rlabel polysilicon 478 -1525 478 -1525 0 1
rlabel polysilicon 478 -1531 478 -1531 0 3
rlabel polysilicon 485 -1525 485 -1525 0 1
rlabel polysilicon 485 -1531 485 -1531 0 3
rlabel polysilicon 492 -1525 492 -1525 0 1
rlabel polysilicon 492 -1531 492 -1531 0 3
rlabel polysilicon 499 -1525 499 -1525 0 1
rlabel polysilicon 499 -1531 499 -1531 0 3
rlabel polysilicon 506 -1525 506 -1525 0 1
rlabel polysilicon 506 -1531 506 -1531 0 3
rlabel polysilicon 513 -1525 513 -1525 0 1
rlabel polysilicon 513 -1531 513 -1531 0 3
rlabel polysilicon 520 -1525 520 -1525 0 1
rlabel polysilicon 523 -1525 523 -1525 0 2
rlabel polysilicon 527 -1525 527 -1525 0 1
rlabel polysilicon 527 -1531 527 -1531 0 3
rlabel polysilicon 534 -1525 534 -1525 0 1
rlabel polysilicon 537 -1525 537 -1525 0 2
rlabel polysilicon 534 -1531 534 -1531 0 3
rlabel polysilicon 541 -1525 541 -1525 0 1
rlabel polysilicon 541 -1531 541 -1531 0 3
rlabel polysilicon 548 -1525 548 -1525 0 1
rlabel polysilicon 548 -1531 548 -1531 0 3
rlabel polysilicon 555 -1525 555 -1525 0 1
rlabel polysilicon 555 -1531 555 -1531 0 3
rlabel polysilicon 562 -1525 562 -1525 0 1
rlabel polysilicon 562 -1531 562 -1531 0 3
rlabel polysilicon 569 -1525 569 -1525 0 1
rlabel polysilicon 569 -1531 569 -1531 0 3
rlabel polysilicon 576 -1525 576 -1525 0 1
rlabel polysilicon 576 -1531 576 -1531 0 3
rlabel polysilicon 583 -1525 583 -1525 0 1
rlabel polysilicon 583 -1531 583 -1531 0 3
rlabel polysilicon 590 -1525 590 -1525 0 1
rlabel polysilicon 590 -1531 590 -1531 0 3
rlabel polysilicon 597 -1525 597 -1525 0 1
rlabel polysilicon 597 -1531 597 -1531 0 3
rlabel polysilicon 600 -1531 600 -1531 0 4
rlabel polysilicon 604 -1525 604 -1525 0 1
rlabel polysilicon 604 -1531 604 -1531 0 3
rlabel polysilicon 611 -1525 611 -1525 0 1
rlabel polysilicon 611 -1531 611 -1531 0 3
rlabel polysilicon 618 -1525 618 -1525 0 1
rlabel polysilicon 625 -1525 625 -1525 0 1
rlabel polysilicon 625 -1531 625 -1531 0 3
rlabel polysilicon 632 -1525 632 -1525 0 1
rlabel polysilicon 632 -1531 632 -1531 0 3
rlabel polysilicon 639 -1525 639 -1525 0 1
rlabel polysilicon 639 -1531 639 -1531 0 3
rlabel polysilicon 646 -1525 646 -1525 0 1
rlabel polysilicon 646 -1531 646 -1531 0 3
rlabel polysilicon 653 -1525 653 -1525 0 1
rlabel polysilicon 653 -1531 653 -1531 0 3
rlabel polysilicon 660 -1525 660 -1525 0 1
rlabel polysilicon 660 -1531 660 -1531 0 3
rlabel polysilicon 667 -1525 667 -1525 0 1
rlabel polysilicon 667 -1531 667 -1531 0 3
rlabel polysilicon 674 -1525 674 -1525 0 1
rlabel polysilicon 674 -1531 674 -1531 0 3
rlabel polysilicon 681 -1525 681 -1525 0 1
rlabel polysilicon 681 -1531 681 -1531 0 3
rlabel polysilicon 688 -1525 688 -1525 0 1
rlabel polysilicon 688 -1531 688 -1531 0 3
rlabel polysilicon 695 -1525 695 -1525 0 1
rlabel polysilicon 695 -1531 695 -1531 0 3
rlabel polysilicon 702 -1525 702 -1525 0 1
rlabel polysilicon 702 -1531 702 -1531 0 3
rlabel polysilicon 709 -1525 709 -1525 0 1
rlabel polysilicon 709 -1531 709 -1531 0 3
rlabel polysilicon 716 -1525 716 -1525 0 1
rlabel polysilicon 716 -1531 716 -1531 0 3
rlabel polysilicon 723 -1525 723 -1525 0 1
rlabel polysilicon 723 -1531 723 -1531 0 3
rlabel polysilicon 730 -1525 730 -1525 0 1
rlabel polysilicon 730 -1531 730 -1531 0 3
rlabel polysilicon 737 -1525 737 -1525 0 1
rlabel polysilicon 737 -1531 737 -1531 0 3
rlabel polysilicon 744 -1525 744 -1525 0 1
rlabel polysilicon 744 -1531 744 -1531 0 3
rlabel polysilicon 751 -1525 751 -1525 0 1
rlabel polysilicon 751 -1531 751 -1531 0 3
rlabel polysilicon 5 -1610 5 -1610 0 4
rlabel polysilicon 12 -1604 12 -1604 0 2
rlabel polysilicon 16 -1604 16 -1604 0 1
rlabel polysilicon 16 -1610 16 -1610 0 3
rlabel polysilicon 23 -1604 23 -1604 0 1
rlabel polysilicon 23 -1610 23 -1610 0 3
rlabel polysilicon 30 -1604 30 -1604 0 1
rlabel polysilicon 30 -1610 30 -1610 0 3
rlabel polysilicon 37 -1604 37 -1604 0 1
rlabel polysilicon 37 -1610 37 -1610 0 3
rlabel polysilicon 44 -1604 44 -1604 0 1
rlabel polysilicon 47 -1610 47 -1610 0 4
rlabel polysilicon 51 -1604 51 -1604 0 1
rlabel polysilicon 51 -1610 51 -1610 0 3
rlabel polysilicon 58 -1604 58 -1604 0 1
rlabel polysilicon 58 -1610 58 -1610 0 3
rlabel polysilicon 65 -1604 65 -1604 0 1
rlabel polysilicon 65 -1610 65 -1610 0 3
rlabel polysilicon 72 -1604 72 -1604 0 1
rlabel polysilicon 72 -1610 72 -1610 0 3
rlabel polysilicon 82 -1604 82 -1604 0 2
rlabel polysilicon 82 -1610 82 -1610 0 4
rlabel polysilicon 89 -1604 89 -1604 0 2
rlabel polysilicon 86 -1610 86 -1610 0 3
rlabel polysilicon 89 -1610 89 -1610 0 4
rlabel polysilicon 93 -1604 93 -1604 0 1
rlabel polysilicon 93 -1610 93 -1610 0 3
rlabel polysilicon 103 -1604 103 -1604 0 2
rlabel polysilicon 107 -1604 107 -1604 0 1
rlabel polysilicon 107 -1610 107 -1610 0 3
rlabel polysilicon 114 -1604 114 -1604 0 1
rlabel polysilicon 117 -1604 117 -1604 0 2
rlabel polysilicon 114 -1610 114 -1610 0 3
rlabel polysilicon 121 -1604 121 -1604 0 1
rlabel polysilicon 121 -1610 121 -1610 0 3
rlabel polysilicon 128 -1604 128 -1604 0 1
rlabel polysilicon 128 -1610 128 -1610 0 3
rlabel polysilicon 138 -1604 138 -1604 0 2
rlabel polysilicon 135 -1610 135 -1610 0 3
rlabel polysilicon 138 -1610 138 -1610 0 4
rlabel polysilicon 142 -1610 142 -1610 0 3
rlabel polysilicon 152 -1604 152 -1604 0 2
rlabel polysilicon 152 -1610 152 -1610 0 4
rlabel polysilicon 156 -1604 156 -1604 0 1
rlabel polysilicon 156 -1610 156 -1610 0 3
rlabel polysilicon 163 -1604 163 -1604 0 1
rlabel polysilicon 163 -1610 163 -1610 0 3
rlabel polysilicon 170 -1604 170 -1604 0 1
rlabel polysilicon 170 -1610 170 -1610 0 3
rlabel polysilicon 177 -1604 177 -1604 0 1
rlabel polysilicon 177 -1610 177 -1610 0 3
rlabel polysilicon 184 -1604 184 -1604 0 1
rlabel polysilicon 184 -1610 184 -1610 0 3
rlabel polysilicon 191 -1604 191 -1604 0 1
rlabel polysilicon 191 -1610 191 -1610 0 3
rlabel polysilicon 194 -1610 194 -1610 0 4
rlabel polysilicon 198 -1604 198 -1604 0 1
rlabel polysilicon 198 -1610 198 -1610 0 3
rlabel polysilicon 205 -1604 205 -1604 0 1
rlabel polysilicon 205 -1610 205 -1610 0 3
rlabel polysilicon 212 -1604 212 -1604 0 1
rlabel polysilicon 212 -1610 212 -1610 0 3
rlabel polysilicon 219 -1604 219 -1604 0 1
rlabel polysilicon 219 -1610 219 -1610 0 3
rlabel polysilicon 226 -1604 226 -1604 0 1
rlabel polysilicon 226 -1610 226 -1610 0 3
rlabel polysilicon 233 -1604 233 -1604 0 1
rlabel polysilicon 236 -1604 236 -1604 0 2
rlabel polysilicon 233 -1610 233 -1610 0 3
rlabel polysilicon 240 -1604 240 -1604 0 1
rlabel polysilicon 240 -1610 240 -1610 0 3
rlabel polysilicon 247 -1604 247 -1604 0 1
rlabel polysilicon 247 -1610 247 -1610 0 3
rlabel polysilicon 254 -1604 254 -1604 0 1
rlabel polysilicon 254 -1610 254 -1610 0 3
rlabel polysilicon 261 -1604 261 -1604 0 1
rlabel polysilicon 261 -1610 261 -1610 0 3
rlabel polysilicon 268 -1604 268 -1604 0 1
rlabel polysilicon 268 -1610 268 -1610 0 3
rlabel polysilicon 275 -1604 275 -1604 0 1
rlabel polysilicon 278 -1604 278 -1604 0 2
rlabel polysilicon 275 -1610 275 -1610 0 3
rlabel polysilicon 278 -1610 278 -1610 0 4
rlabel polysilicon 282 -1604 282 -1604 0 1
rlabel polysilicon 282 -1610 282 -1610 0 3
rlabel polysilicon 289 -1604 289 -1604 0 1
rlabel polysilicon 289 -1610 289 -1610 0 3
rlabel polysilicon 296 -1604 296 -1604 0 1
rlabel polysilicon 296 -1610 296 -1610 0 3
rlabel polysilicon 303 -1604 303 -1604 0 1
rlabel polysilicon 306 -1604 306 -1604 0 2
rlabel polysilicon 306 -1610 306 -1610 0 4
rlabel polysilicon 310 -1604 310 -1604 0 1
rlabel polysilicon 313 -1604 313 -1604 0 2
rlabel polysilicon 320 -1604 320 -1604 0 2
rlabel polysilicon 317 -1610 317 -1610 0 3
rlabel polysilicon 320 -1610 320 -1610 0 4
rlabel polysilicon 324 -1604 324 -1604 0 1
rlabel polysilicon 324 -1610 324 -1610 0 3
rlabel polysilicon 331 -1604 331 -1604 0 1
rlabel polysilicon 331 -1610 331 -1610 0 3
rlabel polysilicon 341 -1604 341 -1604 0 2
rlabel polysilicon 338 -1610 338 -1610 0 3
rlabel polysilicon 345 -1604 345 -1604 0 1
rlabel polysilicon 345 -1610 345 -1610 0 3
rlabel polysilicon 352 -1604 352 -1604 0 1
rlabel polysilicon 352 -1610 352 -1610 0 3
rlabel polysilicon 362 -1604 362 -1604 0 2
rlabel polysilicon 359 -1610 359 -1610 0 3
rlabel polysilicon 362 -1610 362 -1610 0 4
rlabel polysilicon 366 -1604 366 -1604 0 1
rlabel polysilicon 373 -1604 373 -1604 0 1
rlabel polysilicon 373 -1610 373 -1610 0 3
rlabel polysilicon 380 -1604 380 -1604 0 1
rlabel polysilicon 380 -1610 380 -1610 0 3
rlabel polysilicon 387 -1604 387 -1604 0 1
rlabel polysilicon 387 -1610 387 -1610 0 3
rlabel polysilicon 394 -1604 394 -1604 0 1
rlabel polysilicon 394 -1610 394 -1610 0 3
rlabel polysilicon 401 -1604 401 -1604 0 1
rlabel polysilicon 401 -1610 401 -1610 0 3
rlabel polysilicon 408 -1604 408 -1604 0 1
rlabel polysilicon 411 -1604 411 -1604 0 2
rlabel polysilicon 408 -1610 408 -1610 0 3
rlabel polysilicon 411 -1610 411 -1610 0 4
rlabel polysilicon 415 -1604 415 -1604 0 1
rlabel polysilicon 415 -1610 415 -1610 0 3
rlabel polysilicon 422 -1604 422 -1604 0 1
rlabel polysilicon 422 -1610 422 -1610 0 3
rlabel polysilicon 429 -1604 429 -1604 0 1
rlabel polysilicon 429 -1610 429 -1610 0 3
rlabel polysilicon 436 -1604 436 -1604 0 1
rlabel polysilicon 439 -1610 439 -1610 0 4
rlabel polysilicon 443 -1604 443 -1604 0 1
rlabel polysilicon 443 -1610 443 -1610 0 3
rlabel polysilicon 446 -1610 446 -1610 0 4
rlabel polysilicon 450 -1604 450 -1604 0 1
rlabel polysilicon 450 -1610 450 -1610 0 3
rlabel polysilicon 457 -1604 457 -1604 0 1
rlabel polysilicon 457 -1610 457 -1610 0 3
rlabel polysilicon 464 -1604 464 -1604 0 1
rlabel polysilicon 464 -1610 464 -1610 0 3
rlabel polysilicon 471 -1604 471 -1604 0 1
rlabel polysilicon 471 -1610 471 -1610 0 3
rlabel polysilicon 478 -1604 478 -1604 0 1
rlabel polysilicon 478 -1610 478 -1610 0 3
rlabel polysilicon 485 -1604 485 -1604 0 1
rlabel polysilicon 488 -1604 488 -1604 0 2
rlabel polysilicon 492 -1604 492 -1604 0 1
rlabel polysilicon 492 -1610 492 -1610 0 3
rlabel polysilicon 499 -1604 499 -1604 0 1
rlabel polysilicon 499 -1610 499 -1610 0 3
rlabel polysilicon 506 -1604 506 -1604 0 1
rlabel polysilicon 506 -1610 506 -1610 0 3
rlabel polysilicon 513 -1604 513 -1604 0 1
rlabel polysilicon 513 -1610 513 -1610 0 3
rlabel polysilicon 520 -1604 520 -1604 0 1
rlabel polysilicon 520 -1610 520 -1610 0 3
rlabel polysilicon 527 -1604 527 -1604 0 1
rlabel polysilicon 527 -1610 527 -1610 0 3
rlabel polysilicon 534 -1604 534 -1604 0 1
rlabel polysilicon 534 -1610 534 -1610 0 3
rlabel polysilicon 541 -1604 541 -1604 0 1
rlabel polysilicon 541 -1610 541 -1610 0 3
rlabel polysilicon 548 -1604 548 -1604 0 1
rlabel polysilicon 548 -1610 548 -1610 0 3
rlabel polysilicon 555 -1610 555 -1610 0 3
rlabel polysilicon 558 -1610 558 -1610 0 4
rlabel polysilicon 562 -1604 562 -1604 0 1
rlabel polysilicon 562 -1610 562 -1610 0 3
rlabel polysilicon 569 -1604 569 -1604 0 1
rlabel polysilicon 569 -1610 569 -1610 0 3
rlabel polysilicon 576 -1604 576 -1604 0 1
rlabel polysilicon 576 -1610 576 -1610 0 3
rlabel polysilicon 583 -1604 583 -1604 0 1
rlabel polysilicon 583 -1610 583 -1610 0 3
rlabel polysilicon 590 -1604 590 -1604 0 1
rlabel polysilicon 590 -1610 590 -1610 0 3
rlabel polysilicon 597 -1604 597 -1604 0 1
rlabel polysilicon 597 -1610 597 -1610 0 3
rlabel polysilicon 604 -1604 604 -1604 0 1
rlabel polysilicon 604 -1610 604 -1610 0 3
rlabel polysilicon 611 -1604 611 -1604 0 1
rlabel polysilicon 611 -1610 611 -1610 0 3
rlabel polysilicon 618 -1604 618 -1604 0 1
rlabel polysilicon 618 -1610 618 -1610 0 3
rlabel polysilicon 625 -1604 625 -1604 0 1
rlabel polysilicon 625 -1610 625 -1610 0 3
rlabel polysilicon 632 -1604 632 -1604 0 1
rlabel polysilicon 632 -1610 632 -1610 0 3
rlabel polysilicon 639 -1604 639 -1604 0 1
rlabel polysilicon 639 -1610 639 -1610 0 3
rlabel polysilicon 646 -1604 646 -1604 0 1
rlabel polysilicon 646 -1610 646 -1610 0 3
rlabel polysilicon 653 -1604 653 -1604 0 1
rlabel polysilicon 653 -1610 653 -1610 0 3
rlabel polysilicon 660 -1604 660 -1604 0 1
rlabel polysilicon 660 -1610 660 -1610 0 3
rlabel polysilicon 667 -1604 667 -1604 0 1
rlabel polysilicon 667 -1610 667 -1610 0 3
rlabel polysilicon 674 -1604 674 -1604 0 1
rlabel polysilicon 674 -1610 674 -1610 0 3
rlabel polysilicon 681 -1604 681 -1604 0 1
rlabel polysilicon 681 -1610 681 -1610 0 3
rlabel polysilicon 9 -1673 9 -1673 0 1
rlabel polysilicon 9 -1679 9 -1679 0 3
rlabel polysilicon 16 -1673 16 -1673 0 1
rlabel polysilicon 16 -1679 16 -1679 0 3
rlabel polysilicon 23 -1673 23 -1673 0 1
rlabel polysilicon 23 -1679 23 -1679 0 3
rlabel polysilicon 30 -1673 30 -1673 0 1
rlabel polysilicon 37 -1673 37 -1673 0 1
rlabel polysilicon 37 -1679 37 -1679 0 3
rlabel polysilicon 47 -1679 47 -1679 0 4
rlabel polysilicon 51 -1673 51 -1673 0 1
rlabel polysilicon 58 -1673 58 -1673 0 1
rlabel polysilicon 58 -1679 58 -1679 0 3
rlabel polysilicon 65 -1673 65 -1673 0 1
rlabel polysilicon 65 -1679 65 -1679 0 3
rlabel polysilicon 72 -1673 72 -1673 0 1
rlabel polysilicon 72 -1679 72 -1679 0 3
rlabel polysilicon 79 -1673 79 -1673 0 1
rlabel polysilicon 79 -1679 79 -1679 0 3
rlabel polysilicon 86 -1673 86 -1673 0 1
rlabel polysilicon 86 -1679 86 -1679 0 3
rlabel polysilicon 93 -1673 93 -1673 0 1
rlabel polysilicon 93 -1679 93 -1679 0 3
rlabel polysilicon 100 -1673 100 -1673 0 1
rlabel polysilicon 110 -1673 110 -1673 0 2
rlabel polysilicon 107 -1679 107 -1679 0 3
rlabel polysilicon 114 -1673 114 -1673 0 1
rlabel polysilicon 117 -1673 117 -1673 0 2
rlabel polysilicon 114 -1679 114 -1679 0 3
rlabel polysilicon 121 -1673 121 -1673 0 1
rlabel polysilicon 121 -1679 121 -1679 0 3
rlabel polysilicon 128 -1673 128 -1673 0 1
rlabel polysilicon 128 -1679 128 -1679 0 3
rlabel polysilicon 135 -1673 135 -1673 0 1
rlabel polysilicon 135 -1679 135 -1679 0 3
rlabel polysilicon 142 -1679 142 -1679 0 3
rlabel polysilicon 145 -1679 145 -1679 0 4
rlabel polysilicon 149 -1673 149 -1673 0 1
rlabel polysilicon 149 -1679 149 -1679 0 3
rlabel polysilicon 156 -1673 156 -1673 0 1
rlabel polysilicon 156 -1679 156 -1679 0 3
rlabel polysilicon 163 -1673 163 -1673 0 1
rlabel polysilicon 163 -1679 163 -1679 0 3
rlabel polysilicon 170 -1673 170 -1673 0 1
rlabel polysilicon 173 -1673 173 -1673 0 2
rlabel polysilicon 173 -1679 173 -1679 0 4
rlabel polysilicon 177 -1673 177 -1673 0 1
rlabel polysilicon 177 -1679 177 -1679 0 3
rlabel polysilicon 187 -1673 187 -1673 0 2
rlabel polysilicon 187 -1679 187 -1679 0 4
rlabel polysilicon 191 -1673 191 -1673 0 1
rlabel polysilicon 198 -1673 198 -1673 0 1
rlabel polysilicon 198 -1679 198 -1679 0 3
rlabel polysilicon 205 -1673 205 -1673 0 1
rlabel polysilicon 205 -1679 205 -1679 0 3
rlabel polysilicon 212 -1673 212 -1673 0 1
rlabel polysilicon 212 -1679 212 -1679 0 3
rlabel polysilicon 219 -1673 219 -1673 0 1
rlabel polysilicon 219 -1679 219 -1679 0 3
rlabel polysilicon 226 -1673 226 -1673 0 1
rlabel polysilicon 226 -1679 226 -1679 0 3
rlabel polysilicon 233 -1673 233 -1673 0 1
rlabel polysilicon 233 -1679 233 -1679 0 3
rlabel polysilicon 236 -1679 236 -1679 0 4
rlabel polysilicon 243 -1679 243 -1679 0 4
rlabel polysilicon 247 -1673 247 -1673 0 1
rlabel polysilicon 247 -1679 247 -1679 0 3
rlabel polysilicon 254 -1673 254 -1673 0 1
rlabel polysilicon 254 -1679 254 -1679 0 3
rlabel polysilicon 261 -1679 261 -1679 0 3
rlabel polysilicon 264 -1679 264 -1679 0 4
rlabel polysilicon 268 -1673 268 -1673 0 1
rlabel polysilicon 268 -1679 268 -1679 0 3
rlabel polysilicon 275 -1673 275 -1673 0 1
rlabel polysilicon 275 -1679 275 -1679 0 3
rlabel polysilicon 282 -1673 282 -1673 0 1
rlabel polysilicon 282 -1679 282 -1679 0 3
rlabel polysilicon 289 -1673 289 -1673 0 1
rlabel polysilicon 292 -1673 292 -1673 0 2
rlabel polysilicon 289 -1679 289 -1679 0 3
rlabel polysilicon 292 -1679 292 -1679 0 4
rlabel polysilicon 296 -1673 296 -1673 0 1
rlabel polysilicon 299 -1673 299 -1673 0 2
rlabel polysilicon 296 -1679 296 -1679 0 3
rlabel polysilicon 306 -1679 306 -1679 0 4
rlabel polysilicon 310 -1673 310 -1673 0 1
rlabel polysilicon 310 -1679 310 -1679 0 3
rlabel polysilicon 317 -1673 317 -1673 0 1
rlabel polysilicon 317 -1679 317 -1679 0 3
rlabel polysilicon 324 -1673 324 -1673 0 1
rlabel polysilicon 324 -1679 324 -1679 0 3
rlabel polysilicon 331 -1679 331 -1679 0 3
rlabel polysilicon 334 -1679 334 -1679 0 4
rlabel polysilicon 338 -1673 338 -1673 0 1
rlabel polysilicon 345 -1673 345 -1673 0 1
rlabel polysilicon 345 -1679 345 -1679 0 3
rlabel polysilicon 352 -1679 352 -1679 0 3
rlabel polysilicon 355 -1679 355 -1679 0 4
rlabel polysilicon 359 -1673 359 -1673 0 1
rlabel polysilicon 359 -1679 359 -1679 0 3
rlabel polysilicon 362 -1679 362 -1679 0 4
rlabel polysilicon 366 -1673 366 -1673 0 1
rlabel polysilicon 369 -1673 369 -1673 0 2
rlabel polysilicon 376 -1673 376 -1673 0 2
rlabel polysilicon 373 -1679 373 -1679 0 3
rlabel polysilicon 380 -1673 380 -1673 0 1
rlabel polysilicon 380 -1679 380 -1679 0 3
rlabel polysilicon 387 -1673 387 -1673 0 1
rlabel polysilicon 390 -1679 390 -1679 0 4
rlabel polysilicon 394 -1673 394 -1673 0 1
rlabel polysilicon 394 -1679 394 -1679 0 3
rlabel polysilicon 401 -1673 401 -1673 0 1
rlabel polysilicon 401 -1679 401 -1679 0 3
rlabel polysilicon 408 -1673 408 -1673 0 1
rlabel polysilicon 408 -1679 408 -1679 0 3
rlabel polysilicon 415 -1673 415 -1673 0 1
rlabel polysilicon 415 -1679 415 -1679 0 3
rlabel polysilicon 422 -1673 422 -1673 0 1
rlabel polysilicon 422 -1679 422 -1679 0 3
rlabel polysilicon 429 -1673 429 -1673 0 1
rlabel polysilicon 429 -1679 429 -1679 0 3
rlabel polysilicon 436 -1673 436 -1673 0 1
rlabel polysilicon 436 -1679 436 -1679 0 3
rlabel polysilicon 443 -1673 443 -1673 0 1
rlabel polysilicon 443 -1679 443 -1679 0 3
rlabel polysilicon 450 -1673 450 -1673 0 1
rlabel polysilicon 450 -1679 450 -1679 0 3
rlabel polysilicon 457 -1673 457 -1673 0 1
rlabel polysilicon 457 -1679 457 -1679 0 3
rlabel polysilicon 464 -1673 464 -1673 0 1
rlabel polysilicon 464 -1679 464 -1679 0 3
rlabel polysilicon 471 -1673 471 -1673 0 1
rlabel polysilicon 471 -1679 471 -1679 0 3
rlabel polysilicon 478 -1673 478 -1673 0 1
rlabel polysilicon 478 -1679 478 -1679 0 3
rlabel polysilicon 485 -1673 485 -1673 0 1
rlabel polysilicon 485 -1679 485 -1679 0 3
rlabel polysilicon 492 -1673 492 -1673 0 1
rlabel polysilicon 492 -1679 492 -1679 0 3
rlabel polysilicon 499 -1673 499 -1673 0 1
rlabel polysilicon 499 -1679 499 -1679 0 3
rlabel polysilicon 506 -1673 506 -1673 0 1
rlabel polysilicon 506 -1679 506 -1679 0 3
rlabel polysilicon 513 -1673 513 -1673 0 1
rlabel polysilicon 513 -1679 513 -1679 0 3
rlabel polysilicon 520 -1673 520 -1673 0 1
rlabel polysilicon 520 -1679 520 -1679 0 3
rlabel polysilicon 527 -1673 527 -1673 0 1
rlabel polysilicon 527 -1679 527 -1679 0 3
rlabel polysilicon 534 -1673 534 -1673 0 1
rlabel polysilicon 534 -1679 534 -1679 0 3
rlabel polysilicon 541 -1673 541 -1673 0 1
rlabel polysilicon 541 -1679 541 -1679 0 3
rlabel polysilicon 548 -1673 548 -1673 0 1
rlabel polysilicon 548 -1679 548 -1679 0 3
rlabel polysilicon 555 -1673 555 -1673 0 1
rlabel polysilicon 555 -1679 555 -1679 0 3
rlabel polysilicon 562 -1673 562 -1673 0 1
rlabel polysilicon 562 -1679 562 -1679 0 3
rlabel polysilicon 569 -1673 569 -1673 0 1
rlabel polysilicon 569 -1679 569 -1679 0 3
rlabel polysilicon 576 -1673 576 -1673 0 1
rlabel polysilicon 576 -1679 576 -1679 0 3
rlabel polysilicon 583 -1673 583 -1673 0 1
rlabel polysilicon 583 -1679 583 -1679 0 3
rlabel polysilicon 590 -1673 590 -1673 0 1
rlabel polysilicon 590 -1679 590 -1679 0 3
rlabel polysilicon 597 -1673 597 -1673 0 1
rlabel polysilicon 597 -1679 597 -1679 0 3
rlabel polysilicon 611 -1673 611 -1673 0 1
rlabel polysilicon 611 -1679 611 -1679 0 3
rlabel polysilicon 618 -1679 618 -1679 0 3
rlabel polysilicon 621 -1679 621 -1679 0 4
rlabel polysilicon 649 -1673 649 -1673 0 2
rlabel polysilicon 649 -1679 649 -1679 0 4
rlabel polysilicon 660 -1673 660 -1673 0 1
rlabel polysilicon 660 -1679 660 -1679 0 3
rlabel polysilicon 677 -1673 677 -1673 0 2
rlabel polysilicon 681 -1673 681 -1673 0 1
rlabel polysilicon 681 -1679 681 -1679 0 3
rlabel polysilicon 9 -1730 9 -1730 0 1
rlabel polysilicon 9 -1736 9 -1736 0 3
rlabel polysilicon 16 -1730 16 -1730 0 1
rlabel polysilicon 16 -1736 16 -1736 0 3
rlabel polysilicon 23 -1730 23 -1730 0 1
rlabel polysilicon 23 -1736 23 -1736 0 3
rlabel polysilicon 30 -1730 30 -1730 0 1
rlabel polysilicon 40 -1730 40 -1730 0 2
rlabel polysilicon 44 -1730 44 -1730 0 1
rlabel polysilicon 44 -1736 44 -1736 0 3
rlabel polysilicon 51 -1730 51 -1730 0 1
rlabel polysilicon 51 -1736 51 -1736 0 3
rlabel polysilicon 58 -1730 58 -1730 0 1
rlabel polysilicon 58 -1736 58 -1736 0 3
rlabel polysilicon 65 -1730 65 -1730 0 1
rlabel polysilicon 65 -1736 65 -1736 0 3
rlabel polysilicon 72 -1730 72 -1730 0 1
rlabel polysilicon 72 -1736 72 -1736 0 3
rlabel polysilicon 79 -1730 79 -1730 0 1
rlabel polysilicon 79 -1736 79 -1736 0 3
rlabel polysilicon 86 -1730 86 -1730 0 1
rlabel polysilicon 86 -1736 86 -1736 0 3
rlabel polysilicon 93 -1736 93 -1736 0 3
rlabel polysilicon 103 -1736 103 -1736 0 4
rlabel polysilicon 107 -1730 107 -1730 0 1
rlabel polysilicon 107 -1736 107 -1736 0 3
rlabel polysilicon 114 -1730 114 -1730 0 1
rlabel polysilicon 114 -1736 114 -1736 0 3
rlabel polysilicon 121 -1730 121 -1730 0 1
rlabel polysilicon 124 -1730 124 -1730 0 2
rlabel polysilicon 128 -1730 128 -1730 0 1
rlabel polysilicon 131 -1730 131 -1730 0 2
rlabel polysilicon 135 -1730 135 -1730 0 1
rlabel polysilicon 135 -1736 135 -1736 0 3
rlabel polysilicon 142 -1730 142 -1730 0 1
rlabel polysilicon 145 -1736 145 -1736 0 4
rlabel polysilicon 152 -1736 152 -1736 0 4
rlabel polysilicon 159 -1730 159 -1730 0 2
rlabel polysilicon 159 -1736 159 -1736 0 4
rlabel polysilicon 163 -1730 163 -1730 0 1
rlabel polysilicon 163 -1736 163 -1736 0 3
rlabel polysilicon 170 -1730 170 -1730 0 1
rlabel polysilicon 170 -1736 170 -1736 0 3
rlabel polysilicon 177 -1736 177 -1736 0 3
rlabel polysilicon 184 -1730 184 -1730 0 1
rlabel polysilicon 187 -1730 187 -1730 0 2
rlabel polysilicon 191 -1730 191 -1730 0 1
rlabel polysilicon 191 -1736 191 -1736 0 3
rlabel polysilicon 198 -1730 198 -1730 0 1
rlabel polysilicon 198 -1736 198 -1736 0 3
rlabel polysilicon 208 -1736 208 -1736 0 4
rlabel polysilicon 212 -1730 212 -1730 0 1
rlabel polysilicon 212 -1736 212 -1736 0 3
rlabel polysilicon 219 -1730 219 -1730 0 1
rlabel polysilicon 219 -1736 219 -1736 0 3
rlabel polysilicon 226 -1730 226 -1730 0 1
rlabel polysilicon 226 -1736 226 -1736 0 3
rlabel polysilicon 233 -1730 233 -1730 0 1
rlabel polysilicon 233 -1736 233 -1736 0 3
rlabel polysilicon 240 -1730 240 -1730 0 1
rlabel polysilicon 243 -1736 243 -1736 0 4
rlabel polysilicon 247 -1730 247 -1730 0 1
rlabel polysilicon 250 -1730 250 -1730 0 2
rlabel polysilicon 250 -1736 250 -1736 0 4
rlabel polysilicon 257 -1730 257 -1730 0 2
rlabel polysilicon 257 -1736 257 -1736 0 4
rlabel polysilicon 261 -1730 261 -1730 0 1
rlabel polysilicon 261 -1736 261 -1736 0 3
rlabel polysilicon 268 -1730 268 -1730 0 1
rlabel polysilicon 271 -1730 271 -1730 0 2
rlabel polysilicon 268 -1736 268 -1736 0 3
rlabel polysilicon 275 -1730 275 -1730 0 1
rlabel polysilicon 275 -1736 275 -1736 0 3
rlabel polysilicon 282 -1730 282 -1730 0 1
rlabel polysilicon 282 -1736 282 -1736 0 3
rlabel polysilicon 289 -1730 289 -1730 0 1
rlabel polysilicon 292 -1736 292 -1736 0 4
rlabel polysilicon 296 -1730 296 -1730 0 1
rlabel polysilicon 296 -1736 296 -1736 0 3
rlabel polysilicon 303 -1730 303 -1730 0 1
rlabel polysilicon 303 -1736 303 -1736 0 3
rlabel polysilicon 310 -1730 310 -1730 0 1
rlabel polysilicon 313 -1730 313 -1730 0 2
rlabel polysilicon 310 -1736 310 -1736 0 3
rlabel polysilicon 317 -1730 317 -1730 0 1
rlabel polysilicon 320 -1730 320 -1730 0 2
rlabel polysilicon 324 -1730 324 -1730 0 1
rlabel polysilicon 324 -1736 324 -1736 0 3
rlabel polysilicon 331 -1730 331 -1730 0 1
rlabel polysilicon 331 -1736 331 -1736 0 3
rlabel polysilicon 338 -1730 338 -1730 0 1
rlabel polysilicon 345 -1730 345 -1730 0 1
rlabel polysilicon 345 -1736 345 -1736 0 3
rlabel polysilicon 352 -1736 352 -1736 0 3
rlabel polysilicon 355 -1736 355 -1736 0 4
rlabel polysilicon 359 -1730 359 -1730 0 1
rlabel polysilicon 362 -1736 362 -1736 0 4
rlabel polysilicon 366 -1730 366 -1730 0 1
rlabel polysilicon 366 -1736 366 -1736 0 3
rlabel polysilicon 373 -1730 373 -1730 0 1
rlabel polysilicon 376 -1730 376 -1730 0 2
rlabel polysilicon 380 -1730 380 -1730 0 1
rlabel polysilicon 380 -1736 380 -1736 0 3
rlabel polysilicon 394 -1730 394 -1730 0 1
rlabel polysilicon 394 -1736 394 -1736 0 3
rlabel polysilicon 401 -1730 401 -1730 0 1
rlabel polysilicon 401 -1736 401 -1736 0 3
rlabel polysilicon 408 -1730 408 -1730 0 1
rlabel polysilicon 408 -1736 408 -1736 0 3
rlabel polysilicon 415 -1730 415 -1730 0 1
rlabel polysilicon 415 -1736 415 -1736 0 3
rlabel polysilicon 422 -1730 422 -1730 0 1
rlabel polysilicon 422 -1736 422 -1736 0 3
rlabel polysilicon 429 -1730 429 -1730 0 1
rlabel polysilicon 429 -1736 429 -1736 0 3
rlabel polysilicon 436 -1730 436 -1730 0 1
rlabel polysilicon 436 -1736 436 -1736 0 3
rlabel polysilicon 446 -1730 446 -1730 0 2
rlabel polysilicon 457 -1730 457 -1730 0 1
rlabel polysilicon 460 -1736 460 -1736 0 4
rlabel polysilicon 464 -1730 464 -1730 0 1
rlabel polysilicon 464 -1736 464 -1736 0 3
rlabel polysilicon 471 -1730 471 -1730 0 1
rlabel polysilicon 471 -1736 471 -1736 0 3
rlabel polysilicon 478 -1730 478 -1730 0 1
rlabel polysilicon 478 -1736 478 -1736 0 3
rlabel polysilicon 485 -1730 485 -1730 0 1
rlabel polysilicon 485 -1736 485 -1736 0 3
rlabel polysilicon 492 -1730 492 -1730 0 1
rlabel polysilicon 492 -1736 492 -1736 0 3
rlabel polysilicon 499 -1730 499 -1730 0 1
rlabel polysilicon 499 -1736 499 -1736 0 3
rlabel polysilicon 520 -1730 520 -1730 0 1
rlabel polysilicon 520 -1736 520 -1736 0 3
rlabel polysilicon 527 -1730 527 -1730 0 1
rlabel polysilicon 527 -1736 527 -1736 0 3
rlabel polysilicon 555 -1730 555 -1730 0 1
rlabel polysilicon 555 -1736 555 -1736 0 3
rlabel polysilicon 579 -1730 579 -1730 0 2
rlabel polysilicon 618 -1730 618 -1730 0 1
rlabel polysilicon 618 -1736 618 -1736 0 3
rlabel polysilicon 653 -1730 653 -1730 0 1
rlabel polysilicon 653 -1736 653 -1736 0 3
rlabel polysilicon 670 -1736 670 -1736 0 4
rlabel polysilicon 674 -1730 674 -1730 0 1
rlabel polysilicon 674 -1736 674 -1736 0 3
rlabel polysilicon 37 -1771 37 -1771 0 1
rlabel polysilicon 37 -1777 37 -1777 0 3
rlabel polysilicon 51 -1771 51 -1771 0 1
rlabel polysilicon 51 -1777 51 -1777 0 3
rlabel polysilicon 61 -1777 61 -1777 0 4
rlabel polysilicon 65 -1771 65 -1771 0 1
rlabel polysilicon 65 -1777 65 -1777 0 3
rlabel polysilicon 72 -1771 72 -1771 0 1
rlabel polysilicon 72 -1777 72 -1777 0 3
rlabel polysilicon 86 -1771 86 -1771 0 1
rlabel polysilicon 86 -1777 86 -1777 0 3
rlabel polysilicon 93 -1771 93 -1771 0 1
rlabel polysilicon 93 -1777 93 -1777 0 3
rlabel polysilicon 103 -1777 103 -1777 0 4
rlabel polysilicon 107 -1771 107 -1771 0 1
rlabel polysilicon 117 -1771 117 -1771 0 2
rlabel polysilicon 117 -1777 117 -1777 0 4
rlabel polysilicon 121 -1771 121 -1771 0 1
rlabel polysilicon 124 -1771 124 -1771 0 2
rlabel polysilicon 128 -1771 128 -1771 0 1
rlabel polysilicon 128 -1777 128 -1777 0 3
rlabel polysilicon 135 -1771 135 -1771 0 1
rlabel polysilicon 135 -1777 135 -1777 0 3
rlabel polysilicon 142 -1771 142 -1771 0 1
rlabel polysilicon 142 -1777 142 -1777 0 3
rlabel polysilicon 152 -1771 152 -1771 0 2
rlabel polysilicon 156 -1771 156 -1771 0 1
rlabel polysilicon 159 -1771 159 -1771 0 2
rlabel polysilicon 156 -1777 156 -1777 0 3
rlabel polysilicon 159 -1777 159 -1777 0 4
rlabel polysilicon 163 -1771 163 -1771 0 1
rlabel polysilicon 163 -1777 163 -1777 0 3
rlabel polysilicon 173 -1771 173 -1771 0 2
rlabel polysilicon 177 -1777 177 -1777 0 3
rlabel polysilicon 184 -1777 184 -1777 0 3
rlabel polysilicon 191 -1771 191 -1771 0 1
rlabel polysilicon 191 -1777 191 -1777 0 3
rlabel polysilicon 198 -1771 198 -1771 0 1
rlabel polysilicon 198 -1777 198 -1777 0 3
rlabel polysilicon 205 -1771 205 -1771 0 1
rlabel polysilicon 212 -1777 212 -1777 0 3
rlabel polysilicon 219 -1771 219 -1771 0 1
rlabel polysilicon 219 -1777 219 -1777 0 3
rlabel polysilicon 226 -1771 226 -1771 0 1
rlabel polysilicon 226 -1777 226 -1777 0 3
rlabel polysilicon 233 -1771 233 -1771 0 1
rlabel polysilicon 233 -1777 233 -1777 0 3
rlabel polysilicon 240 -1771 240 -1771 0 1
rlabel polysilicon 240 -1777 240 -1777 0 3
rlabel polysilicon 254 -1771 254 -1771 0 1
rlabel polysilicon 261 -1771 261 -1771 0 1
rlabel polysilicon 261 -1777 261 -1777 0 3
rlabel polysilicon 268 -1771 268 -1771 0 1
rlabel polysilicon 268 -1777 268 -1777 0 3
rlabel polysilicon 275 -1771 275 -1771 0 1
rlabel polysilicon 289 -1771 289 -1771 0 1
rlabel polysilicon 289 -1777 289 -1777 0 3
rlabel polysilicon 296 -1771 296 -1771 0 1
rlabel polysilicon 296 -1777 296 -1777 0 3
rlabel polysilicon 310 -1771 310 -1771 0 1
rlabel polysilicon 310 -1777 310 -1777 0 3
rlabel polysilicon 317 -1771 317 -1771 0 1
rlabel polysilicon 317 -1777 317 -1777 0 3
rlabel polysilicon 324 -1771 324 -1771 0 1
rlabel polysilicon 324 -1777 324 -1777 0 3
rlabel polysilicon 334 -1771 334 -1771 0 2
rlabel polysilicon 334 -1777 334 -1777 0 4
rlabel polysilicon 338 -1771 338 -1771 0 1
rlabel polysilicon 338 -1777 338 -1777 0 3
rlabel polysilicon 345 -1771 345 -1771 0 1
rlabel polysilicon 345 -1777 345 -1777 0 3
rlabel polysilicon 352 -1771 352 -1771 0 1
rlabel polysilicon 352 -1777 352 -1777 0 3
rlabel polysilicon 366 -1771 366 -1771 0 1
rlabel polysilicon 366 -1777 366 -1777 0 3
rlabel polysilicon 383 -1777 383 -1777 0 4
rlabel polysilicon 404 -1771 404 -1771 0 2
rlabel polysilicon 418 -1771 418 -1771 0 2
rlabel polysilicon 418 -1777 418 -1777 0 4
rlabel polysilicon 422 -1771 422 -1771 0 1
rlabel polysilicon 422 -1777 422 -1777 0 3
rlabel polysilicon 429 -1771 429 -1771 0 1
rlabel polysilicon 429 -1777 429 -1777 0 3
rlabel polysilicon 453 -1771 453 -1771 0 2
rlabel polysilicon 460 -1771 460 -1771 0 2
rlabel polysilicon 464 -1771 464 -1771 0 1
rlabel polysilicon 464 -1777 464 -1777 0 3
rlabel polysilicon 471 -1771 471 -1771 0 1
rlabel polysilicon 471 -1777 471 -1777 0 3
rlabel polysilicon 478 -1771 478 -1771 0 1
rlabel polysilicon 478 -1777 478 -1777 0 3
rlabel polysilicon 488 -1771 488 -1771 0 2
rlabel polysilicon 485 -1777 485 -1777 0 3
rlabel polysilicon 502 -1777 502 -1777 0 4
rlabel polysilicon 513 -1771 513 -1771 0 1
rlabel polysilicon 513 -1777 513 -1777 0 3
rlabel polysilicon 520 -1771 520 -1771 0 1
rlabel polysilicon 520 -1777 520 -1777 0 3
rlabel polysilicon 527 -1771 527 -1771 0 1
rlabel polysilicon 527 -1777 527 -1777 0 3
rlabel polysilicon 534 -1771 534 -1771 0 1
rlabel polysilicon 534 -1777 534 -1777 0 3
rlabel polysilicon 541 -1777 541 -1777 0 3
rlabel polysilicon 548 -1771 548 -1771 0 1
rlabel polysilicon 548 -1777 548 -1777 0 3
rlabel polysilicon 562 -1777 562 -1777 0 3
rlabel polysilicon 614 -1777 614 -1777 0 4
rlabel polysilicon 618 -1771 618 -1771 0 1
rlabel polysilicon 618 -1777 618 -1777 0 3
rlabel polysilicon 632 -1771 632 -1771 0 1
rlabel polysilicon 632 -1777 632 -1777 0 3
rlabel polysilicon 51 -1800 51 -1800 0 1
rlabel polysilicon 51 -1806 51 -1806 0 3
rlabel polysilicon 61 -1806 61 -1806 0 4
rlabel polysilicon 89 -1800 89 -1800 0 2
rlabel polysilicon 103 -1800 103 -1800 0 2
rlabel polysilicon 110 -1800 110 -1800 0 2
rlabel polysilicon 117 -1800 117 -1800 0 2
rlabel polysilicon 124 -1800 124 -1800 0 2
rlabel polysilicon 131 -1800 131 -1800 0 2
rlabel polysilicon 135 -1800 135 -1800 0 1
rlabel polysilicon 138 -1800 138 -1800 0 2
rlabel polysilicon 142 -1800 142 -1800 0 1
rlabel polysilicon 145 -1806 145 -1806 0 4
rlabel polysilicon 149 -1800 149 -1800 0 1
rlabel polysilicon 149 -1806 149 -1806 0 3
rlabel polysilicon 156 -1800 156 -1800 0 1
rlabel polysilicon 156 -1806 156 -1806 0 3
rlabel polysilicon 173 -1800 173 -1800 0 2
rlabel polysilicon 177 -1806 177 -1806 0 3
rlabel polysilicon 180 -1806 180 -1806 0 4
rlabel polysilicon 184 -1806 184 -1806 0 3
rlabel polysilicon 205 -1800 205 -1800 0 1
rlabel polysilicon 205 -1806 205 -1806 0 3
rlabel polysilicon 233 -1800 233 -1800 0 1
rlabel polysilicon 233 -1806 233 -1806 0 3
rlabel polysilicon 247 -1800 247 -1800 0 1
rlabel polysilicon 250 -1800 250 -1800 0 2
rlabel polysilicon 254 -1800 254 -1800 0 1
rlabel polysilicon 261 -1800 261 -1800 0 1
rlabel polysilicon 264 -1800 264 -1800 0 2
rlabel polysilicon 261 -1806 261 -1806 0 3
rlabel polysilicon 271 -1806 271 -1806 0 4
rlabel polysilicon 310 -1800 310 -1800 0 1
rlabel polysilicon 352 -1800 352 -1800 0 1
rlabel polysilicon 352 -1806 352 -1806 0 3
rlabel polysilicon 373 -1800 373 -1800 0 1
rlabel polysilicon 387 -1800 387 -1800 0 1
rlabel polysilicon 411 -1800 411 -1800 0 2
rlabel polysilicon 418 -1800 418 -1800 0 2
rlabel polysilicon 418 -1806 418 -1806 0 4
rlabel polysilicon 467 -1800 467 -1800 0 2
rlabel polysilicon 471 -1800 471 -1800 0 1
rlabel polysilicon 471 -1806 471 -1806 0 3
rlabel polysilicon 478 -1806 478 -1806 0 3
rlabel polysilicon 499 -1800 499 -1800 0 1
rlabel polysilicon 520 -1800 520 -1800 0 1
rlabel polysilicon 520 -1806 520 -1806 0 3
rlabel polysilicon 527 -1806 527 -1806 0 3
rlabel polysilicon 639 -1800 639 -1800 0 1
rlabel metal2 58 1 58 1 0 net=1703
rlabel metal2 114 1 114 1 0 net=3055
rlabel metal2 152 1 152 1 0 net=885
rlabel metal2 177 1 177 1 0 net=1567
rlabel metal2 257 1 257 1 0 net=1747
rlabel metal2 124 -1 124 -1 0 net=3327
rlabel metal2 128 -3 128 -3 0 net=1663
rlabel metal2 156 -3 156 -3 0 net=1731
rlabel metal2 184 -3 184 -3 0 net=2739
rlabel metal2 198 -3 198 -3 0 net=3895
rlabel metal2 205 -5 205 -5 0 net=3755
rlabel metal2 44 -16 44 -16 0 net=591
rlabel metal2 72 -16 72 -16 0 net=1705
rlabel metal2 103 -16 103 -16 0 net=2749
rlabel metal2 285 -16 285 -16 0 net=4033
rlabel metal2 79 -18 79 -18 0 net=797
rlabel metal2 205 -18 205 -18 0 net=3757
rlabel metal2 338 -18 338 -18 0 net=3859
rlabel metal2 114 -20 114 -20 0 net=3056
rlabel metal2 177 -20 177 -20 0 net=3896
rlabel metal2 205 -20 205 -20 0 net=3901
rlabel metal2 124 -22 124 -22 0 net=1568
rlabel metal2 222 -22 222 -22 0 net=3328
rlabel metal2 247 -22 247 -22 0 net=1861
rlabel metal2 128 -24 128 -24 0 net=1665
rlabel metal2 149 -24 149 -24 0 net=2707
rlabel metal2 184 -24 184 -24 0 net=2741
rlabel metal2 240 -24 240 -24 0 net=1749
rlabel metal2 271 -24 271 -24 0 net=3961
rlabel metal2 93 -26 93 -26 0 net=2801
rlabel metal2 163 -26 163 -26 0 net=1733
rlabel metal2 212 -26 212 -26 0 net=1685
rlabel metal2 254 -26 254 -26 0 net=1867
rlabel metal2 289 -26 289 -26 0 net=3333
rlabel metal2 313 -26 313 -26 0 net=4027
rlabel metal2 170 -28 170 -28 0 net=887
rlabel metal2 226 -28 226 -28 0 net=3627
rlabel metal2 142 -30 142 -30 0 net=2529
rlabel metal2 163 -32 163 -32 0 net=1297
rlabel metal2 16 -43 16 -43 0 net=1751
rlabel metal2 254 -43 254 -43 0 net=1868
rlabel metal2 345 -43 345 -43 0 net=4035
rlabel metal2 23 -45 23 -45 0 net=1545
rlabel metal2 128 -45 128 -45 0 net=1773
rlabel metal2 163 -45 163 -45 0 net=1299
rlabel metal2 191 -45 191 -45 0 net=798
rlabel metal2 233 -45 233 -45 0 net=2531
rlabel metal2 317 -45 317 -45 0 net=3759
rlabel metal2 387 -45 387 -45 0 net=3861
rlabel metal2 44 -47 44 -47 0 net=1787
rlabel metal2 65 -47 65 -47 0 net=3169
rlabel metal2 114 -47 114 -47 0 net=2101
rlabel metal2 135 -47 135 -47 0 net=1667
rlabel metal2 156 -47 156 -47 0 net=1471
rlabel metal2 205 -47 205 -47 0 net=2742
rlabel metal2 247 -47 247 -47 0 net=1863
rlabel metal2 275 -47 275 -47 0 net=2751
rlabel metal2 338 -47 338 -47 0 net=4029
rlabel metal2 51 -49 51 -49 0 net=3513
rlabel metal2 352 -49 352 -49 0 net=3963
rlabel metal2 404 -49 404 -49 0 net=3977
rlabel metal2 61 -51 61 -51 0 net=223
rlabel metal2 208 -51 208 -51 0 net=3628
rlabel metal2 268 -51 268 -51 0 net=1973
rlabel metal2 282 -51 282 -51 0 net=2623
rlabel metal2 324 -51 324 -51 0 net=3903
rlabel metal2 72 -53 72 -53 0 net=1706
rlabel metal2 170 -53 170 -53 0 net=1025
rlabel metal2 184 -53 184 -53 0 net=889
rlabel metal2 296 -53 296 -53 0 net=3335
rlabel metal2 373 -53 373 -53 0 net=3535
rlabel metal2 82 -55 82 -55 0 net=943
rlabel metal2 184 -55 184 -55 0 net=1647
rlabel metal2 299 -55 299 -55 0 net=3127
rlabel metal2 86 -57 86 -57 0 net=2708
rlabel metal2 212 -57 212 -57 0 net=1687
rlabel metal2 93 -59 93 -59 0 net=2803
rlabel metal2 93 -61 93 -61 0 net=3573
rlabel metal2 100 -63 100 -63 0 net=2815
rlabel metal2 177 -63 177 -63 0 net=1734
rlabel metal2 212 -63 212 -63 0 net=1255
rlabel metal2 198 -65 198 -65 0 net=1925
rlabel metal2 261 -67 261 -67 0 net=671
rlabel metal2 23 -78 23 -78 0 net=1546
rlabel metal2 205 -78 205 -78 0 net=3841
rlabel metal2 37 -80 37 -80 0 net=2245
rlabel metal2 233 -80 233 -80 0 net=1688
rlabel metal2 250 -80 250 -80 0 net=3747
rlabel metal2 44 -82 44 -82 0 net=1789
rlabel metal2 303 -82 303 -82 0 net=3315
rlabel metal2 397 -82 397 -82 0 net=3605
rlabel metal2 58 -84 58 -84 0 net=1473
rlabel metal2 170 -84 170 -84 0 net=1027
rlabel metal2 208 -84 208 -84 0 net=1648
rlabel metal2 254 -84 254 -84 0 net=1865
rlabel metal2 275 -84 275 -84 0 net=1975
rlabel metal2 373 -84 373 -84 0 net=3537
rlabel metal2 436 -84 436 -84 0 net=4037
rlabel metal2 65 -86 65 -86 0 net=3170
rlabel metal2 156 -86 156 -86 0 net=1521
rlabel metal2 254 -86 254 -86 0 net=2624
rlabel metal2 345 -86 345 -86 0 net=3515
rlabel metal2 72 -88 72 -88 0 net=342
rlabel metal2 121 -88 121 -88 0 net=2103
rlabel metal2 222 -88 222 -88 0 net=2177
rlabel metal2 338 -88 338 -88 0 net=2651
rlabel metal2 380 -88 380 -88 0 net=3761
rlabel metal2 79 -90 79 -90 0 net=2187
rlabel metal2 275 -90 275 -90 0 net=2533
rlabel metal2 387 -90 387 -90 0 net=3905
rlabel metal2 16 -92 16 -92 0 net=1753
rlabel metal2 285 -92 285 -92 0 net=3609
rlabel metal2 86 -94 86 -94 0 net=2817
rlabel metal2 107 -94 107 -94 0 net=1257
rlabel metal2 292 -94 292 -94 0 net=4030
rlabel metal2 93 -96 93 -96 0 net=3575
rlabel metal2 93 -98 93 -98 0 net=3121
rlabel metal2 310 -98 310 -98 0 net=1927
rlabel metal2 380 -98 380 -98 0 net=3527
rlabel metal2 128 -100 128 -100 0 net=1774
rlabel metal2 212 -100 212 -100 0 net=1175
rlabel metal2 401 -100 401 -100 0 net=3965
rlabel metal2 128 -102 128 -102 0 net=2109
rlabel metal2 359 -102 359 -102 0 net=3337
rlabel metal2 408 -102 408 -102 0 net=3863
rlabel metal2 135 -104 135 -104 0 net=945
rlabel metal2 324 -104 324 -104 0 net=2805
rlabel metal2 366 -104 366 -104 0 net=3129
rlabel metal2 415 -104 415 -104 0 net=3979
rlabel metal2 149 -106 149 -106 0 net=3311
rlabel metal2 149 -108 149 -108 0 net=1301
rlabel metal2 173 -108 173 -108 0 net=1926
rlabel metal2 331 -108 331 -108 0 net=2753
rlabel metal2 373 -108 373 -108 0 net=3563
rlabel metal2 121 -110 121 -110 0 net=3405
rlabel metal2 331 -110 331 -110 0 net=4209
rlabel metal2 177 -112 177 -112 0 net=1365
rlabel metal2 187 -114 187 -114 0 net=890
rlabel metal2 142 -116 142 -116 0 net=1669
rlabel metal2 142 -118 142 -118 0 net=1859
rlabel metal2 163 -120 163 -120 0 net=747
rlabel metal2 12 -131 12 -131 0 net=2163
rlabel metal2 75 -131 75 -131 0 net=3842
rlabel metal2 520 -131 520 -131 0 net=4211
rlabel metal2 51 -133 51 -133 0 net=667
rlabel metal2 180 -133 180 -133 0 net=2806
rlabel metal2 373 -133 373 -133 0 net=3011
rlabel metal2 383 -133 383 -133 0 net=3748
rlabel metal2 471 -133 471 -133 0 net=3763
rlabel metal2 58 -135 58 -135 0 net=1474
rlabel metal2 296 -135 296 -135 0 net=1791
rlabel metal2 334 -135 334 -135 0 net=3576
rlabel metal2 457 -135 457 -135 0 net=3607
rlabel metal2 58 -137 58 -137 0 net=1537
rlabel metal2 250 -137 250 -137 0 net=1866
rlabel metal2 282 -137 282 -137 0 net=3338
rlabel metal2 415 -137 415 -137 0 net=3565
rlabel metal2 65 -139 65 -139 0 net=1417
rlabel metal2 65 -139 65 -139 0 net=1417
rlabel metal2 79 -139 79 -139 0 net=2189
rlabel metal2 422 -139 422 -139 0 net=3529
rlabel metal2 478 -139 478 -139 0 net=3981
rlabel metal2 79 -141 79 -141 0 net=1689
rlabel metal2 121 -141 121 -141 0 net=3407
rlabel metal2 44 -143 44 -143 0 net=1991
rlabel metal2 128 -143 128 -143 0 net=2111
rlabel metal2 390 -143 390 -143 0 net=4189
rlabel metal2 44 -145 44 -145 0 net=1833
rlabel metal2 240 -145 240 -145 0 net=2534
rlabel metal2 282 -145 282 -145 0 net=3201
rlabel metal2 513 -145 513 -145 0 net=4039
rlabel metal2 89 -147 89 -147 0 net=2104
rlabel metal2 247 -147 247 -147 0 net=1523
rlabel metal2 292 -147 292 -147 0 net=3013
rlabel metal2 499 -147 499 -147 0 net=3967
rlabel metal2 93 -149 93 -149 0 net=3123
rlabel metal2 485 -149 485 -149 0 net=3865
rlabel metal2 93 -151 93 -151 0 net=843
rlabel metal2 296 -151 296 -151 0 net=1633
rlabel metal2 327 -151 327 -151 0 net=3651
rlabel metal2 100 -153 100 -153 0 net=3555
rlabel metal2 100 -155 100 -155 0 net=1303
rlabel metal2 152 -155 152 -155 0 net=3425
rlabel metal2 128 -157 128 -157 0 net=2247
rlabel metal2 261 -157 261 -157 0 net=1755
rlabel metal2 422 -157 422 -157 0 net=3099
rlabel metal2 107 -159 107 -159 0 net=1259
rlabel metal2 303 -159 303 -159 0 net=1977
rlabel metal2 373 -159 373 -159 0 net=3611
rlabel metal2 107 -161 107 -161 0 net=1215
rlabel metal2 163 -161 163 -161 0 net=749
rlabel metal2 163 -161 163 -161 0 net=749
rlabel metal2 170 -161 170 -161 0 net=2871
rlabel metal2 117 -163 117 -163 0 net=879
rlabel metal2 226 -163 226 -163 0 net=1671
rlabel metal2 341 -163 341 -163 0 net=3617
rlabel metal2 135 -165 135 -165 0 net=3659
rlabel metal2 138 -167 138 -167 0 net=1860
rlabel metal2 149 -167 149 -167 0 net=3045
rlabel metal2 142 -169 142 -169 0 net=305
rlabel metal2 352 -169 352 -169 0 net=3906
rlabel metal2 156 -171 156 -171 0 net=863
rlabel metal2 191 -171 191 -171 0 net=947
rlabel metal2 170 -173 170 -173 0 net=1367
rlabel metal2 289 -173 289 -173 0 net=3139
rlabel metal2 177 -175 177 -175 0 net=2015
rlabel metal2 180 -177 180 -177 0 net=1211
rlabel metal2 387 -177 387 -177 0 net=3313
rlabel metal2 191 -179 191 -179 0 net=1963
rlabel metal2 324 -179 324 -179 0 net=1809
rlabel metal2 394 -179 394 -179 0 net=3317
rlabel metal2 198 -181 198 -181 0 net=3187
rlabel metal2 205 -183 205 -183 0 net=1029
rlabel metal2 317 -183 317 -183 0 net=2179
rlabel metal2 408 -183 408 -183 0 net=3131
rlabel metal2 135 -185 135 -185 0 net=2489
rlabel metal2 408 -185 408 -185 0 net=3577
rlabel metal2 212 -187 212 -187 0 net=1177
rlabel metal2 429 -187 429 -187 0 net=3539
rlabel metal2 366 -189 366 -189 0 net=2755
rlabel metal2 436 -189 436 -189 0 net=3517
rlabel metal2 86 -191 86 -191 0 net=2819
rlabel metal2 345 -193 345 -193 0 net=2653
rlabel metal2 310 -195 310 -195 0 net=1929
rlabel metal2 16 -206 16 -206 0 net=576
rlabel metal2 16 -206 16 -206 0 net=576
rlabel metal2 30 -206 30 -206 0 net=2689
rlabel metal2 30 -206 30 -206 0 net=2689
rlabel metal2 33 -206 33 -206 0 net=2016
rlabel metal2 597 -206 597 -206 0 net=3619
rlabel metal2 51 -208 51 -208 0 net=1543
rlabel metal2 215 -208 215 -208 0 net=3652
rlabel metal2 65 -210 65 -210 0 net=1418
rlabel metal2 205 -210 205 -210 0 net=1213
rlabel metal2 243 -210 243 -210 0 net=3314
rlabel metal2 520 -210 520 -210 0 net=4041
rlabel metal2 79 -212 79 -212 0 net=1690
rlabel metal2 310 -212 310 -212 0 net=1811
rlabel metal2 338 -212 338 -212 0 net=3188
rlabel metal2 44 -214 44 -214 0 net=1835
rlabel metal2 366 -214 366 -214 0 net=2655
rlabel metal2 411 -214 411 -214 0 net=3202
rlabel metal2 513 -214 513 -214 0 net=3409
rlabel metal2 590 -214 590 -214 0 net=3969
rlabel metal2 89 -216 89 -216 0 net=2783
rlabel metal2 464 -216 464 -216 0 net=3047
rlabel metal2 527 -216 527 -216 0 net=3519
rlabel metal2 597 -216 597 -216 0 net=3983
rlabel metal2 100 -218 100 -218 0 net=1304
rlabel metal2 187 -218 187 -218 0 net=1030
rlabel metal2 254 -218 254 -218 0 net=1930
rlabel metal2 373 -218 373 -218 0 net=3613
rlabel metal2 625 -218 625 -218 0 net=4191
rlabel metal2 103 -220 103 -220 0 net=517
rlabel metal2 198 -220 198 -220 0 net=3014
rlabel metal2 464 -220 464 -220 0 net=3133
rlabel metal2 492 -220 492 -220 0 net=3141
rlabel metal2 492 -220 492 -220 0 net=3141
rlabel metal2 632 -220 632 -220 0 net=4213
rlabel metal2 72 -222 72 -222 0 net=2165
rlabel metal2 208 -222 208 -222 0 net=3426
rlabel metal2 72 -224 72 -224 0 net=1023
rlabel metal2 114 -224 114 -224 0 net=2105
rlabel metal2 219 -224 219 -224 0 net=881
rlabel metal2 247 -224 247 -224 0 net=2833
rlabel metal2 478 -224 478 -224 0 net=3125
rlabel metal2 478 -224 478 -224 0 net=3125
rlabel metal2 485 -224 485 -224 0 net=3557
rlabel metal2 58 -226 58 -226 0 net=1539
rlabel metal2 257 -226 257 -226 0 net=1978
rlabel metal2 373 -226 373 -226 0 net=2191
rlabel metal2 499 -226 499 -226 0 net=3867
rlabel metal2 58 -228 58 -228 0 net=3329
rlabel metal2 534 -228 534 -228 0 net=3541
rlabel metal2 114 -230 114 -230 0 net=1965
rlabel metal2 257 -230 257 -230 0 net=3578
rlabel metal2 121 -232 121 -232 0 net=1993
rlabel metal2 359 -232 359 -232 0 net=2113
rlabel metal2 387 -232 387 -232 0 net=3608
rlabel metal2 121 -234 121 -234 0 net=3935
rlabel metal2 124 -236 124 -236 0 net=1672
rlabel metal2 313 -236 313 -236 0 net=2872
rlabel metal2 65 -238 65 -238 0 net=1869
rlabel metal2 317 -238 317 -238 0 net=2491
rlabel metal2 548 -238 548 -238 0 net=3765
rlabel metal2 128 -240 128 -240 0 net=2249
rlabel metal2 387 -240 387 -240 0 net=2757
rlabel metal2 576 -240 576 -240 0 net=3849
rlabel metal2 128 -242 128 -242 0 net=1083
rlabel metal2 268 -242 268 -242 0 net=3660
rlabel metal2 135 -244 135 -244 0 net=948
rlabel metal2 429 -244 429 -244 0 net=3101
rlabel metal2 100 -246 100 -246 0 net=789
rlabel metal2 142 -246 142 -246 0 net=750
rlabel metal2 170 -246 170 -246 0 net=1369
rlabel metal2 268 -246 268 -246 0 net=3203
rlabel metal2 93 -248 93 -248 0 net=845
rlabel metal2 191 -248 191 -248 0 net=875
rlabel metal2 275 -248 275 -248 0 net=1525
rlabel metal2 292 -248 292 -248 0 net=2180
rlabel metal2 443 -248 443 -248 0 net=3531
rlabel metal2 89 -250 89 -250 0 net=2251
rlabel metal2 436 -250 436 -250 0 net=2821
rlabel metal2 93 -252 93 -252 0 net=1635
rlabel metal2 299 -252 299 -252 0 net=1792
rlabel metal2 334 -252 334 -252 0 net=4065
rlabel metal2 107 -254 107 -254 0 net=1217
rlabel metal2 282 -254 282 -254 0 net=3566
rlabel metal2 107 -256 107 -256 0 net=865
rlabel metal2 180 -256 180 -256 0 net=4109
rlabel metal2 142 -258 142 -258 0 net=1265
rlabel metal2 320 -258 320 -258 0 net=3012
rlabel metal2 149 -260 149 -260 0 net=1179
rlabel metal2 285 -260 285 -260 0 net=3031
rlabel metal2 23 -262 23 -262 0 net=2203
rlabel metal2 285 -262 285 -262 0 net=1756
rlabel metal2 425 -262 425 -262 0 net=2763
rlabel metal2 152 -264 152 -264 0 net=1260
rlabel metal2 282 -264 282 -264 0 net=2709
rlabel metal2 261 -266 261 -266 0 net=1339
rlabel metal2 331 -266 331 -266 0 net=3318
rlabel metal2 338 -268 338 -268 0 net=837
rlabel metal2 44 -279 44 -279 0 net=140
rlabel metal2 58 -279 58 -279 0 net=1370
rlabel metal2 219 -279 219 -279 0 net=1541
rlabel metal2 219 -279 219 -279 0 net=1541
rlabel metal2 226 -279 226 -279 0 net=883
rlabel metal2 226 -279 226 -279 0 net=883
rlabel metal2 247 -279 247 -279 0 net=1995
rlabel metal2 355 -279 355 -279 0 net=2758
rlabel metal2 390 -279 390 -279 0 net=3126
rlabel metal2 506 -279 506 -279 0 net=3331
rlabel metal2 667 -279 667 -279 0 net=3621
rlabel metal2 58 -281 58 -281 0 net=2051
rlabel metal2 261 -281 261 -281 0 net=1341
rlabel metal2 282 -281 282 -281 0 net=1812
rlabel metal2 317 -281 317 -281 0 net=3339
rlabel metal2 72 -283 72 -283 0 net=1024
rlabel metal2 187 -283 187 -283 0 net=1237
rlabel metal2 282 -283 282 -283 0 net=839
rlabel metal2 341 -283 341 -283 0 net=3048
rlabel metal2 555 -283 555 -283 0 net=3355
rlabel metal2 72 -285 72 -285 0 net=4110
rlabel metal2 583 -285 583 -285 0 net=3937
rlabel metal2 89 -287 89 -287 0 net=2853
rlabel metal2 513 -287 513 -287 0 net=3411
rlabel metal2 89 -289 89 -289 0 net=3558
rlabel metal2 527 -289 527 -289 0 net=3521
rlabel metal2 590 -289 590 -289 0 net=3971
rlabel metal2 100 -291 100 -291 0 net=3975
rlabel metal2 107 -293 107 -293 0 net=867
rlabel metal2 285 -293 285 -293 0 net=2883
rlabel metal2 492 -293 492 -293 0 net=3143
rlabel metal2 534 -293 534 -293 0 net=3543
rlabel metal2 604 -293 604 -293 0 net=4043
rlabel metal2 16 -295 16 -295 0 net=3713
rlabel metal2 107 -297 107 -297 0 net=1085
rlabel metal2 145 -297 145 -297 0 net=118
rlabel metal2 163 -297 163 -297 0 net=1219
rlabel metal2 289 -297 289 -297 0 net=1527
rlabel metal2 289 -297 289 -297 0 net=1527
rlabel metal2 296 -297 296 -297 0 net=4192
rlabel metal2 54 -299 54 -299 0 net=3907
rlabel metal2 65 -301 65 -301 0 net=1871
rlabel metal2 299 -301 299 -301 0 net=2037
rlabel metal2 362 -301 362 -301 0 net=3061
rlabel metal2 541 -301 541 -301 0 net=3615
rlabel metal2 114 -303 114 -303 0 net=1967
rlabel metal2 149 -303 149 -303 0 net=1180
rlabel metal2 306 -303 306 -303 0 net=4214
rlabel metal2 114 -305 114 -305 0 net=2979
rlabel metal2 320 -305 320 -305 0 net=3102
rlabel metal2 450 -305 450 -305 0 net=3033
rlabel metal2 541 -305 541 -305 0 net=3869
rlabel metal2 30 -307 30 -307 0 net=2691
rlabel metal2 436 -307 436 -307 0 net=2765
rlabel metal2 464 -307 464 -307 0 net=3135
rlabel metal2 562 -307 562 -307 0 net=4067
rlabel metal2 30 -309 30 -309 0 net=616
rlabel metal2 121 -309 121 -309 0 net=183
rlabel metal2 401 -309 401 -309 0 net=2493
rlabel metal2 401 -309 401 -309 0 net=2493
rlabel metal2 415 -309 415 -309 0 net=2711
rlabel metal2 443 -309 443 -309 0 net=2823
rlabel metal2 499 -309 499 -309 0 net=3205
rlabel metal2 576 -309 576 -309 0 net=3851
rlabel metal2 23 -311 23 -311 0 net=803
rlabel metal2 142 -311 142 -311 0 net=1267
rlabel metal2 320 -311 320 -311 0 net=3919
rlabel metal2 159 -313 159 -313 0 net=2250
rlabel metal2 408 -313 408 -313 0 net=2657
rlabel metal2 471 -313 471 -313 0 net=3533
rlabel metal2 65 -315 65 -315 0 net=2443
rlabel metal2 415 -315 415 -315 0 net=2785
rlabel metal2 457 -315 457 -315 0 net=2835
rlabel metal2 79 -317 79 -317 0 net=2797
rlabel metal2 51 -319 51 -319 0 net=1544
rlabel metal2 142 -319 142 -319 0 net=2263
rlabel metal2 394 -319 394 -319 0 net=2253
rlabel metal2 37 -321 37 -321 0 net=2373
rlabel metal2 170 -321 170 -321 0 net=847
rlabel metal2 191 -321 191 -321 0 net=876
rlabel metal2 352 -321 352 -321 0 net=2521
rlabel metal2 135 -323 135 -323 0 net=791
rlabel metal2 191 -323 191 -323 0 net=2167
rlabel metal2 201 -323 201 -323 0 net=180
rlabel metal2 324 -323 324 -323 0 net=1837
rlabel metal2 366 -323 366 -323 0 net=2193
rlabel metal2 135 -325 135 -325 0 net=2204
rlabel metal2 313 -325 313 -325 0 net=2685
rlabel metal2 184 -327 184 -327 0 net=2107
rlabel metal2 324 -327 324 -327 0 net=3021
rlabel metal2 149 -329 149 -329 0 net=959
rlabel metal2 205 -329 205 -329 0 net=1214
rlabel metal2 369 -329 369 -329 0 net=3766
rlabel metal2 93 -331 93 -331 0 net=1637
rlabel metal2 233 -331 233 -331 0 net=2115
rlabel metal2 548 -331 548 -331 0 net=3985
rlabel metal2 93 -333 93 -333 0 net=981
rlabel metal2 9 -344 9 -344 0 net=3340
rlabel metal2 709 -344 709 -344 0 net=3623
rlabel metal2 12 -346 12 -346 0 net=513
rlabel metal2 68 -346 68 -346 0 net=3332
rlabel metal2 23 -348 23 -348 0 net=1969
rlabel metal2 142 -348 142 -348 0 net=2108
rlabel metal2 313 -348 313 -348 0 net=2194
rlabel metal2 436 -348 436 -348 0 net=2713
rlabel metal2 436 -348 436 -348 0 net=2713
rlabel metal2 467 -348 467 -348 0 net=3908
rlabel metal2 30 -350 30 -350 0 net=170
rlabel metal2 89 -350 89 -350 0 net=3034
rlabel metal2 548 -350 548 -350 0 net=3987
rlabel metal2 37 -352 37 -352 0 net=2374
rlabel metal2 51 -352 51 -352 0 net=1781
rlabel metal2 506 -352 506 -352 0 net=3207
rlabel metal2 555 -352 555 -352 0 net=3357
rlabel metal2 555 -352 555 -352 0 net=3357
rlabel metal2 597 -352 597 -352 0 net=3921
rlabel metal2 37 -354 37 -354 0 net=2825
rlabel metal2 471 -354 471 -354 0 net=2837
rlabel metal2 44 -356 44 -356 0 net=2039
rlabel metal2 338 -356 338 -356 0 net=2658
rlabel metal2 450 -356 450 -356 0 net=2767
rlabel metal2 72 -358 72 -358 0 net=1609
rlabel metal2 117 -358 117 -358 0 net=2168
rlabel metal2 198 -358 198 -358 0 net=1997
rlabel metal2 275 -358 275 -358 0 net=1343
rlabel metal2 275 -358 275 -358 0 net=1343
rlabel metal2 282 -358 282 -358 0 net=840
rlabel metal2 390 -358 390 -358 0 net=3221
rlabel metal2 75 -360 75 -360 0 net=2444
rlabel metal2 411 -360 411 -360 0 net=4049
rlabel metal2 79 -362 79 -362 0 net=2729
rlabel metal2 163 -362 163 -362 0 net=868
rlabel metal2 226 -362 226 -362 0 net=884
rlabel metal2 355 -362 355 -362 0 net=3976
rlabel metal2 86 -364 86 -364 0 net=1951
rlabel metal2 107 -364 107 -364 0 net=1087
rlabel metal2 177 -364 177 -364 0 net=849
rlabel metal2 219 -364 219 -364 0 net=1542
rlabel metal2 233 -364 233 -364 0 net=2117
rlabel metal2 390 -364 390 -364 0 net=2786
rlabel metal2 443 -364 443 -364 0 net=2885
rlabel metal2 590 -364 590 -364 0 net=3616
rlabel metal2 86 -366 86 -366 0 net=983
rlabel metal2 110 -366 110 -366 0 net=1919
rlabel metal2 233 -366 233 -366 0 net=1269
rlabel metal2 282 -366 282 -366 0 net=675
rlabel metal2 359 -366 359 -366 0 net=3544
rlabel metal2 590 -366 590 -366 0 net=3853
rlabel metal2 58 -368 58 -368 0 net=2053
rlabel metal2 394 -368 394 -368 0 net=2523
rlabel metal2 450 -368 450 -368 0 net=2855
rlabel metal2 485 -368 485 -368 0 net=3063
rlabel metal2 583 -368 583 -368 0 net=3671
rlabel metal2 58 -370 58 -370 0 net=903
rlabel metal2 201 -370 201 -370 0 net=1638
rlabel metal2 247 -370 247 -370 0 net=1221
rlabel metal2 268 -370 268 -370 0 net=1431
rlabel metal2 317 -370 317 -370 0 net=2265
rlabel metal2 457 -370 457 -370 0 net=2799
rlabel metal2 121 -372 121 -372 0 net=805
rlabel metal2 254 -372 254 -372 0 net=2353
rlabel metal2 457 -372 457 -372 0 net=3137
rlabel metal2 121 -374 121 -374 0 net=2254
rlabel metal2 492 -374 492 -374 0 net=3247
rlabel metal2 128 -376 128 -376 0 net=793
rlabel metal2 187 -376 187 -376 0 net=2153
rlabel metal2 296 -376 296 -376 0 net=1873
rlabel metal2 324 -376 324 -376 0 net=3412
rlabel metal2 114 -378 114 -378 0 net=2981
rlabel metal2 303 -378 303 -378 0 net=1839
rlabel metal2 352 -378 352 -378 0 net=3155
rlabel metal2 135 -380 135 -380 0 net=2061
rlabel metal2 334 -380 334 -380 0 net=2271
rlabel metal2 422 -380 422 -380 0 net=3145
rlabel metal2 135 -382 135 -382 0 net=1529
rlabel metal2 345 -382 345 -382 0 net=2687
rlabel metal2 380 -382 380 -382 0 net=3972
rlabel metal2 142 -384 142 -384 0 net=961
rlabel metal2 170 -384 170 -384 0 net=1239
rlabel metal2 289 -384 289 -384 0 net=2693
rlabel metal2 492 -384 492 -384 0 net=3939
rlabel metal2 93 -386 93 -386 0 net=1877
rlabel metal2 261 -386 261 -386 0 net=813
rlabel metal2 495 -386 495 -386 0 net=3483
rlabel metal2 562 -386 562 -386 0 net=4069
rlabel metal2 355 -388 355 -388 0 net=3925
rlabel metal2 373 -390 373 -390 0 net=3534
rlabel metal2 604 -390 604 -390 0 net=3715
rlabel metal2 541 -392 541 -392 0 net=3871
rlabel metal2 604 -392 604 -392 0 net=4045
rlabel metal2 243 -394 243 -394 0 net=3349
rlabel metal2 562 -394 562 -394 0 net=3523
rlabel metal2 324 -396 324 -396 0 net=3369
rlabel metal2 401 -398 401 -398 0 net=2495
rlabel metal2 401 -400 401 -400 0 net=3023
rlabel metal2 9 -411 9 -411 0 net=3275
rlabel metal2 100 -411 100 -411 0 net=1952
rlabel metal2 198 -411 198 -411 0 net=1998
rlabel metal2 268 -411 268 -411 0 net=1432
rlabel metal2 383 -411 383 -411 0 net=3484
rlabel metal2 562 -411 562 -411 0 net=3525
rlabel metal2 656 -411 656 -411 0 net=2838
rlabel metal2 716 -411 716 -411 0 net=3625
rlabel metal2 16 -413 16 -413 0 net=2731
rlabel metal2 93 -413 93 -413 0 net=3146
rlabel metal2 425 -413 425 -413 0 net=3872
rlabel metal2 597 -413 597 -413 0 net=3923
rlabel metal2 23 -415 23 -415 0 net=1970
rlabel metal2 114 -415 114 -415 0 net=1241
rlabel metal2 180 -415 180 -415 0 net=3716
rlabel metal2 30 -417 30 -417 0 net=2043
rlabel metal2 121 -417 121 -417 0 net=3345
rlabel metal2 583 -417 583 -417 0 net=3673
rlabel metal2 37 -419 37 -419 0 net=2826
rlabel metal2 156 -419 156 -419 0 net=809
rlabel metal2 247 -419 247 -419 0 net=1223
rlabel metal2 275 -419 275 -419 0 net=1345
rlabel metal2 275 -419 275 -419 0 net=1345
rlabel metal2 282 -419 282 -419 0 net=3156
rlabel metal2 534 -419 534 -419 0 net=3223
rlabel metal2 569 -419 569 -419 0 net=3371
rlabel metal2 37 -421 37 -421 0 net=1783
rlabel metal2 58 -421 58 -421 0 net=904
rlabel metal2 373 -421 373 -421 0 net=1795
rlabel metal2 432 -421 432 -421 0 net=2743
rlabel metal2 513 -421 513 -421 0 net=3249
rlabel metal2 604 -421 604 -421 0 net=4047
rlabel metal2 44 -423 44 -423 0 net=2041
rlabel metal2 100 -423 100 -423 0 net=743
rlabel metal2 135 -423 135 -423 0 net=1531
rlabel metal2 303 -423 303 -423 0 net=1841
rlabel metal2 387 -423 387 -423 0 net=344
rlabel metal2 464 -423 464 -423 0 net=3443
rlabel metal2 611 -423 611 -423 0 net=3927
rlabel metal2 44 -425 44 -425 0 net=963
rlabel metal2 163 -425 163 -425 0 net=1089
rlabel metal2 390 -425 390 -425 0 net=3988
rlabel metal2 625 -425 625 -425 0 net=4051
rlabel metal2 58 -427 58 -427 0 net=795
rlabel metal2 135 -427 135 -427 0 net=2155
rlabel metal2 219 -427 219 -427 0 net=1921
rlabel metal2 233 -427 233 -427 0 net=1271
rlabel metal2 296 -427 296 -427 0 net=2982
rlabel metal2 390 -427 390 -427 0 net=3003
rlabel metal2 541 -427 541 -427 0 net=3351
rlabel metal2 65 -429 65 -429 0 net=995
rlabel metal2 149 -429 149 -429 0 net=1879
rlabel metal2 212 -429 212 -429 0 net=851
rlabel metal2 313 -429 313 -429 0 net=2463
rlabel metal2 481 -429 481 -429 0 net=3493
rlabel metal2 68 -431 68 -431 0 net=3157
rlabel metal2 555 -431 555 -431 0 net=3359
rlabel metal2 72 -433 72 -433 0 net=1610
rlabel metal2 149 -433 149 -433 0 net=833
rlabel metal2 324 -433 324 -433 0 net=2055
rlabel metal2 401 -433 401 -433 0 net=3025
rlabel metal2 72 -435 72 -435 0 net=154
rlabel metal2 408 -435 408 -435 0 net=4070
rlabel metal2 86 -437 86 -437 0 net=985
rlabel metal2 327 -437 327 -437 0 net=2800
rlabel metal2 590 -437 590 -437 0 net=3855
rlabel metal2 86 -439 86 -439 0 net=2355
rlabel metal2 331 -439 331 -439 0 net=2181
rlabel metal2 450 -439 450 -439 0 net=2857
rlabel metal2 170 -441 170 -441 0 net=1445
rlabel metal2 345 -441 345 -441 0 net=2688
rlabel metal2 411 -441 411 -441 0 net=3427
rlabel metal2 177 -443 177 -443 0 net=2063
rlabel metal2 254 -443 254 -443 0 net=2267
rlabel metal2 359 -443 359 -443 0 net=608
rlabel metal2 436 -443 436 -443 0 net=2715
rlabel metal2 128 -445 128 -445 0 net=1419
rlabel metal2 184 -445 184 -445 0 net=2694
rlabel metal2 310 -445 310 -445 0 net=1875
rlabel metal2 366 -445 366 -445 0 net=2119
rlabel metal2 436 -445 436 -445 0 net=3485
rlabel metal2 184 -447 184 -447 0 net=2017
rlabel metal2 229 -447 229 -447 0 net=1623
rlabel metal2 439 -447 439 -447 0 net=139
rlabel metal2 191 -449 191 -449 0 net=807
rlabel metal2 443 -449 443 -449 0 net=2887
rlabel metal2 51 -451 51 -451 0 net=1651
rlabel metal2 198 -451 198 -451 0 net=815
rlabel metal2 289 -451 289 -451 0 net=2273
rlabel metal2 492 -451 492 -451 0 net=3941
rlabel metal2 166 -453 166 -453 0 net=2009
rlabel metal2 394 -453 394 -453 0 net=3138
rlabel metal2 485 -453 485 -453 0 net=3065
rlabel metal2 502 -453 502 -453 0 net=3365
rlabel metal2 341 -455 341 -455 0 net=2365
rlabel metal2 506 -455 506 -455 0 net=3209
rlabel metal2 366 -457 366 -457 0 net=2671
rlabel metal2 471 -459 471 -459 0 net=2769
rlabel metal2 471 -461 471 -461 0 net=2497
rlabel metal2 478 -463 478 -463 0 net=3661
rlabel metal2 415 -465 415 -465 0 net=2525
rlabel metal2 58 -476 58 -476 0 net=796
rlabel metal2 177 -476 177 -476 0 net=3360
rlabel metal2 639 -476 639 -476 0 net=3675
rlabel metal2 716 -476 716 -476 0 net=3626
rlabel metal2 75 -478 75 -478 0 net=4147
rlabel metal2 23 -480 23 -480 0 net=1915
rlabel metal2 79 -480 79 -480 0 net=4245
rlabel metal2 79 -482 79 -482 0 net=2157
rlabel metal2 145 -482 145 -482 0 net=3942
rlabel metal2 723 -482 723 -482 0 net=3373
rlabel metal2 93 -484 93 -484 0 net=2042
rlabel metal2 152 -484 152 -484 0 net=1880
rlabel metal2 219 -484 219 -484 0 net=2019
rlabel metal2 243 -484 243 -484 0 net=1876
rlabel metal2 359 -484 359 -484 0 net=2793
rlabel metal2 646 -484 646 -484 0 net=3857
rlabel metal2 37 -486 37 -486 0 net=1785
rlabel metal2 121 -486 121 -486 0 net=744
rlabel metal2 198 -486 198 -486 0 net=817
rlabel metal2 198 -486 198 -486 0 net=817
rlabel metal2 219 -486 219 -486 0 net=2269
rlabel metal2 275 -486 275 -486 0 net=1347
rlabel metal2 275 -486 275 -486 0 net=1347
rlabel metal2 289 -486 289 -486 0 net=2275
rlabel metal2 555 -486 555 -486 0 net=3211
rlabel metal2 674 -486 674 -486 0 net=4053
rlabel metal2 121 -488 121 -488 0 net=1224
rlabel metal2 289 -488 289 -488 0 net=2183
rlabel metal2 345 -488 345 -488 0 net=1797
rlabel metal2 383 -488 383 -488 0 net=2129
rlabel metal2 422 -488 422 -488 0 net=3301
rlabel metal2 51 -490 51 -490 0 net=1653
rlabel metal2 352 -490 352 -490 0 net=1843
rlabel metal2 366 -490 366 -490 0 net=2716
rlabel metal2 555 -490 555 -490 0 net=3429
rlabel metal2 597 -490 597 -490 0 net=3445
rlabel metal2 16 -492 16 -492 0 net=2733
rlabel metal2 30 -494 30 -494 0 net=2044
rlabel metal2 124 -494 124 -494 0 net=3773
rlabel metal2 128 -496 128 -496 0 net=1421
rlabel metal2 390 -496 390 -496 0 net=3366
rlabel metal2 107 -498 107 -498 0 net=997
rlabel metal2 135 -498 135 -498 0 net=1159
rlabel metal2 44 -500 44 -500 0 net=965
rlabel metal2 149 -500 149 -500 0 net=835
rlabel metal2 394 -500 394 -500 0 net=4193
rlabel metal2 44 -502 44 -502 0 net=1243
rlabel metal2 156 -502 156 -502 0 net=811
rlabel metal2 156 -502 156 -502 0 net=811
rlabel metal2 180 -502 180 -502 0 net=2064
rlabel metal2 247 -502 247 -502 0 net=987
rlabel metal2 247 -502 247 -502 0 net=987
rlabel metal2 408 -502 408 -502 0 net=2255
rlabel metal2 439 -502 439 -502 0 net=3924
rlabel metal2 61 -504 61 -504 0 net=915
rlabel metal2 187 -504 187 -504 0 net=1090
rlabel metal2 401 -504 401 -504 0 net=2121
rlabel metal2 411 -504 411 -504 0 net=2526
rlabel metal2 513 -504 513 -504 0 net=2859
rlabel metal2 562 -504 562 -504 0 net=3225
rlabel metal2 625 -504 625 -504 0 net=3487
rlabel metal2 65 -506 65 -506 0 net=3273
rlabel metal2 170 -508 170 -508 0 net=3175
rlabel metal2 576 -508 576 -508 0 net=3347
rlabel metal2 170 -510 170 -510 0 net=1273
rlabel metal2 303 -510 303 -510 0 net=1447
rlabel metal2 429 -510 429 -510 0 net=3526
rlabel metal2 191 -512 191 -512 0 net=1829
rlabel metal2 324 -512 324 -512 0 net=2057
rlabel metal2 432 -512 432 -512 0 net=2957
rlabel metal2 142 -514 142 -514 0 net=1457
rlabel metal2 317 -514 317 -514 0 net=1625
rlabel metal2 432 -514 432 -514 0 net=3662
rlabel metal2 212 -516 212 -516 0 net=808
rlabel metal2 303 -516 303 -516 0 net=4059
rlabel metal2 226 -518 226 -518 0 net=1922
rlabel metal2 397 -518 397 -518 0 net=3379
rlabel metal2 226 -520 226 -520 0 net=853
rlabel metal2 240 -520 240 -520 0 net=1533
rlabel metal2 443 -520 443 -520 0 net=4048
rlabel metal2 233 -522 233 -522 0 net=1813
rlabel metal2 387 -522 387 -522 0 net=3639
rlabel metal2 240 -524 240 -524 0 net=1885
rlabel metal2 443 -524 443 -524 0 net=3928
rlabel metal2 261 -526 261 -526 0 net=2011
rlabel metal2 478 -526 478 -526 0 net=3005
rlabel metal2 534 -526 534 -526 0 net=3027
rlabel metal2 583 -526 583 -526 0 net=3353
rlabel metal2 282 -528 282 -528 0 net=979
rlabel metal2 453 -528 453 -528 0 net=2791
rlabel metal2 632 -528 632 -528 0 net=3495
rlabel metal2 9 -530 9 -530 0 net=3277
rlabel metal2 492 -532 492 -532 0 net=3067
rlabel metal2 446 -534 446 -534 0 net=2589
rlabel metal2 506 -534 506 -534 0 net=2771
rlabel metal2 261 -536 261 -536 0 net=1137
rlabel metal2 513 -536 513 -536 0 net=3159
rlabel metal2 320 -538 320 -538 0 net=2695
rlabel metal2 520 -538 520 -538 0 net=2889
rlabel metal2 499 -540 499 -540 0 net=2745
rlabel metal2 541 -540 541 -540 0 net=3251
rlabel metal2 464 -542 464 -542 0 net=2465
rlabel metal2 457 -544 457 -544 0 net=2367
rlabel metal2 485 -544 485 -544 0 net=2673
rlabel metal2 86 -546 86 -546 0 net=2357
rlabel metal2 471 -546 471 -546 0 net=2499
rlabel metal2 68 -548 68 -548 0 net=2435
rlabel metal2 26 -550 26 -550 0 net=99
rlabel metal2 86 -550 86 -550 0 net=891
rlabel metal2 16 -561 16 -561 0 net=2123
rlabel metal2 418 -561 418 -561 0 net=3858
rlabel metal2 779 -561 779 -561 0 net=3375
rlabel metal2 23 -563 23 -563 0 net=1916
rlabel metal2 58 -563 58 -563 0 net=1161
rlabel metal2 156 -563 156 -563 0 net=812
rlabel metal2 187 -563 187 -563 0 net=980
rlabel metal2 306 -563 306 -563 0 net=1626
rlabel metal2 355 -563 355 -563 0 net=2746
rlabel metal2 541 -563 541 -563 0 net=3253
rlabel metal2 562 -563 562 -563 0 net=3177
rlabel metal2 562 -563 562 -563 0 net=3177
rlabel metal2 23 -565 23 -565 0 net=1999
rlabel metal2 128 -565 128 -565 0 net=999
rlabel metal2 166 -565 166 -565 0 net=2890
rlabel metal2 30 -567 30 -567 0 net=271
rlabel metal2 100 -567 100 -567 0 net=1971
rlabel metal2 177 -567 177 -567 0 net=753
rlabel metal2 205 -567 205 -567 0 net=836
rlabel metal2 219 -567 219 -567 0 net=2270
rlabel metal2 366 -567 366 -567 0 net=2674
rlabel metal2 541 -567 541 -567 0 net=3029
rlabel metal2 33 -569 33 -569 0 net=548
rlabel metal2 61 -569 61 -569 0 net=3274
rlabel metal2 40 -571 40 -571 0 net=6
rlabel metal2 40 -571 40 -571 0 net=6
rlabel metal2 44 -571 44 -571 0 net=1244
rlabel metal2 191 -571 191 -571 0 net=1831
rlabel metal2 369 -571 369 -571 0 net=3915
rlabel metal2 47 -573 47 -573 0 net=3354
rlabel metal2 51 -575 51 -575 0 net=967
rlabel metal2 394 -575 394 -575 0 net=3348
rlabel metal2 65 -577 65 -577 0 net=382
rlabel metal2 411 -577 411 -577 0 net=2779
rlabel metal2 625 -577 625 -577 0 net=3497
rlabel metal2 65 -579 65 -579 0 net=1815
rlabel metal2 394 -579 394 -579 0 net=4194
rlabel metal2 72 -581 72 -581 0 net=2734
rlabel metal2 646 -581 646 -581 0 net=3775
rlabel metal2 72 -583 72 -583 0 net=2839
rlabel metal2 191 -583 191 -583 0 net=819
rlabel metal2 212 -583 212 -583 0 net=4229
rlabel metal2 107 -585 107 -585 0 net=966
rlabel metal2 212 -585 212 -585 0 net=2059
rlabel metal2 425 -585 425 -585 0 net=2792
rlabel metal2 590 -585 590 -585 0 net=3303
rlabel metal2 688 -585 688 -585 0 net=4061
rlabel metal2 114 -587 114 -587 0 net=917
rlabel metal2 219 -587 219 -587 0 net=1459
rlabel metal2 338 -587 338 -587 0 net=1448
rlabel metal2 401 -587 401 -587 0 net=2131
rlabel metal2 429 -587 429 -587 0 net=2466
rlabel metal2 597 -587 597 -587 0 net=2959
rlabel metal2 730 -587 730 -587 0 net=4247
rlabel metal2 226 -589 226 -589 0 net=855
rlabel metal2 569 -589 569 -589 0 net=3213
rlabel metal2 226 -591 226 -591 0 net=1139
rlabel metal2 275 -591 275 -591 0 net=1348
rlabel metal2 282 -591 282 -591 0 net=1535
rlabel metal2 310 -591 310 -591 0 net=2277
rlabel metal2 471 -591 471 -591 0 net=2437
rlabel metal2 233 -593 233 -593 0 net=1613
rlabel metal2 331 -593 331 -593 0 net=1654
rlabel metal2 429 -593 429 -593 0 net=2369
rlabel metal2 471 -593 471 -593 0 net=2591
rlabel metal2 604 -593 604 -593 0 net=3447
rlabel metal2 163 -595 163 -595 0 net=38
rlabel metal2 233 -597 233 -597 0 net=2021
rlabel metal2 261 -597 261 -597 0 net=2013
rlabel metal2 432 -597 432 -597 0 net=3676
rlabel metal2 142 -599 142 -599 0 net=4077
rlabel metal2 184 -601 184 -601 0 net=1091
rlabel metal2 275 -601 275 -601 0 net=3813
rlabel metal2 236 -603 236 -603 0 net=4148
rlabel metal2 240 -605 240 -605 0 net=988
rlabel metal2 289 -605 289 -605 0 net=2185
rlabel metal2 331 -605 331 -605 0 net=1887
rlabel metal2 387 -605 387 -605 0 net=3380
rlabel metal2 79 -607 79 -607 0 net=2159
rlabel metal2 247 -607 247 -607 0 net=1423
rlabel metal2 303 -607 303 -607 0 net=2089
rlabel metal2 390 -607 390 -607 0 net=3873
rlabel metal2 79 -609 79 -609 0 net=1275
rlabel metal2 198 -609 198 -609 0 net=2621
rlabel metal2 303 -609 303 -609 0 net=1799
rlabel metal2 348 -609 348 -609 0 net=2509
rlabel metal2 86 -611 86 -611 0 net=893
rlabel metal2 268 -611 268 -611 0 net=1691
rlabel metal2 338 -611 338 -611 0 net=2359
rlabel metal2 464 -611 464 -611 0 net=3431
rlabel metal2 86 -613 86 -613 0 net=3677
rlabel metal2 320 -613 320 -613 0 net=3507
rlabel metal2 478 -613 478 -613 0 net=3007
rlabel metal2 555 -613 555 -613 0 net=4055
rlabel metal2 93 -615 93 -615 0 net=1786
rlabel metal2 352 -615 352 -615 0 net=2794
rlabel metal2 93 -617 93 -617 0 net=2911
rlabel metal2 383 -617 383 -617 0 net=3601
rlabel metal2 443 -619 443 -619 0 net=3226
rlabel metal2 446 -621 446 -621 0 net=3640
rlabel metal2 446 -623 446 -623 0 net=3721
rlabel metal2 450 -625 450 -625 0 net=2861
rlabel metal2 485 -627 485 -627 0 net=2501
rlabel metal2 485 -629 485 -629 0 net=2697
rlabel metal2 513 -629 513 -629 0 net=3161
rlabel metal2 478 -631 478 -631 0 net=2473
rlabel metal2 516 -631 516 -631 0 net=4155
rlabel metal2 506 -633 506 -633 0 net=2773
rlabel metal2 548 -633 548 -633 0 net=3069
rlabel metal2 380 -635 380 -635 0 net=3959
rlabel metal2 583 -635 583 -635 0 net=3279
rlabel metal2 359 -637 359 -637 0 net=1845
rlabel metal2 632 -637 632 -637 0 net=3489
rlabel metal2 359 -639 359 -639 0 net=2257
rlabel metal2 75 -641 75 -641 0 net=2393
rlabel metal2 425 -643 425 -643 0 net=3943
rlabel metal2 58 -654 58 -654 0 net=1162
rlabel metal2 100 -654 100 -654 0 net=1972
rlabel metal2 117 -654 117 -654 0 net=1000
rlabel metal2 166 -654 166 -654 0 net=754
rlabel metal2 184 -654 184 -654 0 net=2160
rlabel metal2 254 -654 254 -654 0 net=1093
rlabel metal2 348 -654 348 -654 0 net=2862
rlabel metal2 474 -654 474 -654 0 net=3973
rlabel metal2 807 -654 807 -654 0 net=3377
rlabel metal2 9 -656 9 -656 0 net=2891
rlabel metal2 117 -656 117 -656 0 net=2622
rlabel metal2 212 -656 212 -656 0 net=2060
rlabel metal2 261 -656 261 -656 0 net=2014
rlabel metal2 282 -656 282 -656 0 net=1536
rlabel metal2 352 -656 352 -656 0 net=2045
rlabel metal2 418 -656 418 -656 0 net=2445
rlabel metal2 555 -656 555 -656 0 net=4057
rlabel metal2 16 -658 16 -658 0 net=2125
rlabel metal2 366 -658 366 -658 0 net=3008
rlabel metal2 597 -658 597 -658 0 net=2510
rlabel metal2 16 -660 16 -660 0 net=2841
rlabel metal2 86 -660 86 -660 0 net=3678
rlabel metal2 124 -660 124 -660 0 net=151
rlabel metal2 443 -660 443 -660 0 net=2807
rlabel metal2 660 -660 660 -660 0 net=2961
rlabel metal2 709 -660 709 -660 0 net=4079
rlabel metal2 51 -662 51 -662 0 net=969
rlabel metal2 107 -662 107 -662 0 net=3280
rlabel metal2 646 -662 646 -662 0 net=3777
rlabel metal2 716 -662 716 -662 0 net=4157
rlabel metal2 58 -664 58 -664 0 net=4215
rlabel metal2 65 -666 65 -666 0 net=1817
rlabel metal2 152 -666 152 -666 0 net=338
rlabel metal2 261 -666 261 -666 0 net=1491
rlabel metal2 380 -666 380 -666 0 net=1847
rlabel metal2 408 -666 408 -666 0 net=2502
rlabel metal2 667 -666 667 -666 0 net=3875
rlabel metal2 730 -666 730 -666 0 net=4249
rlabel metal2 23 -668 23 -668 0 net=2000
rlabel metal2 86 -668 86 -668 0 net=2279
rlabel metal2 411 -668 411 -668 0 net=4217
rlabel metal2 23 -670 23 -670 0 net=1597
rlabel metal2 303 -670 303 -670 0 net=1801
rlabel metal2 422 -670 422 -670 0 net=3162
rlabel metal2 30 -672 30 -672 0 net=1043
rlabel metal2 429 -672 429 -672 0 net=2371
rlabel metal2 590 -672 590 -672 0 net=3305
rlabel metal2 618 -672 618 -672 0 net=3603
rlabel metal2 37 -674 37 -674 0 net=1451
rlabel metal2 443 -674 443 -674 0 net=2475
rlabel metal2 548 -674 548 -674 0 net=3071
rlabel metal2 604 -674 604 -674 0 net=3449
rlabel metal2 653 -674 653 -674 0 net=3815
rlabel metal2 674 -674 674 -674 0 net=3917
rlabel metal2 44 -676 44 -676 0 net=3441
rlabel metal2 681 -676 681 -676 0 net=3945
rlabel metal2 44 -678 44 -678 0 net=949
rlabel metal2 107 -678 107 -678 0 net=989
rlabel metal2 177 -678 177 -678 0 net=2133
rlabel metal2 439 -678 439 -678 0 net=3361
rlabel metal2 576 -678 576 -678 0 net=3255
rlabel metal2 681 -678 681 -678 0 net=4231
rlabel metal2 79 -680 79 -680 0 net=1277
rlabel metal2 310 -680 310 -680 0 net=2361
rlabel metal2 394 -680 394 -680 0 net=2083
rlabel metal2 457 -680 457 -680 0 net=3509
rlabel metal2 688 -680 688 -680 0 net=4063
rlabel metal2 79 -682 79 -682 0 net=1003
rlabel metal2 397 -682 397 -682 0 net=2999
rlabel metal2 632 -682 632 -682 0 net=3491
rlabel metal2 121 -684 121 -684 0 net=3960
rlabel metal2 625 -684 625 -684 0 net=3499
rlabel metal2 639 -684 639 -684 0 net=3723
rlabel metal2 128 -686 128 -686 0 net=1693
rlabel metal2 282 -686 282 -686 0 net=1117
rlabel metal2 467 -686 467 -686 0 net=2341
rlabel metal2 499 -686 499 -686 0 net=2781
rlabel metal2 131 -688 131 -688 0 net=3030
rlabel metal2 569 -688 569 -688 0 net=3215
rlabel metal2 135 -690 135 -690 0 net=919
rlabel metal2 219 -690 219 -690 0 net=1461
rlabel metal2 359 -690 359 -690 0 net=2259
rlabel metal2 471 -690 471 -690 0 net=2593
rlabel metal2 124 -692 124 -692 0 net=2237
rlabel metal2 226 -692 226 -692 0 net=1141
rlabel metal2 292 -692 292 -692 0 net=3115
rlabel metal2 110 -694 110 -694 0 net=721
rlabel metal2 236 -694 236 -694 0 net=3887
rlabel metal2 135 -696 135 -696 0 net=1099
rlabel metal2 156 -696 156 -696 0 net=1832
rlabel metal2 331 -696 331 -696 0 net=1889
rlabel metal2 436 -696 436 -696 0 net=2395
rlabel metal2 506 -696 506 -696 0 net=2775
rlabel metal2 142 -698 142 -698 0 net=2698
rlabel metal2 506 -698 506 -698 0 net=2439
rlabel metal2 47 -700 47 -700 0 net=1759
rlabel metal2 163 -700 163 -700 0 net=3178
rlabel metal2 166 -702 166 -702 0 net=2827
rlabel metal2 184 -704 184 -704 0 net=1111
rlabel metal2 296 -704 296 -704 0 net=1615
rlabel metal2 369 -704 369 -704 0 net=4071
rlabel metal2 173 -706 173 -706 0 net=1021
rlabel metal2 317 -706 317 -706 0 net=1383
rlabel metal2 191 -708 191 -708 0 net=821
rlabel metal2 191 -708 191 -708 0 net=821
rlabel metal2 198 -708 198 -708 0 net=1425
rlabel metal2 324 -708 324 -708 0 net=2186
rlabel metal2 446 -708 446 -708 0 net=1325
rlabel metal2 205 -710 205 -710 0 net=2913
rlabel metal2 170 -712 170 -712 0 net=895
rlabel metal2 233 -712 233 -712 0 net=2023
rlabel metal2 324 -712 324 -712 0 net=2091
rlabel metal2 233 -714 233 -714 0 net=856
rlabel metal2 240 -716 240 -716 0 net=3843
rlabel metal2 247 -718 247 -718 0 net=1247
rlabel metal2 464 -718 464 -718 0 net=3433
rlabel metal2 331 -720 331 -720 0 net=2535
rlabel metal2 334 -722 334 -722 0 net=2943
rlabel metal2 373 -724 373 -724 0 net=2291
rlabel metal2 9 -735 9 -735 0 net=2893
rlabel metal2 9 -735 9 -735 0 net=2893
rlabel metal2 40 -735 40 -735 0 net=1261
rlabel metal2 124 -735 124 -735 0 net=3844
rlabel metal2 817 -735 817 -735 0 net=3378
rlabel metal2 44 -737 44 -737 0 net=950
rlabel metal2 72 -737 72 -737 0 net=920
rlabel metal2 236 -737 236 -737 0 net=463
rlabel metal2 467 -737 467 -737 0 net=4158
rlabel metal2 47 -739 47 -739 0 net=311
rlabel metal2 72 -739 72 -739 0 net=690
rlabel metal2 324 -739 324 -739 0 net=2093
rlabel metal2 474 -739 474 -739 0 net=4064
rlabel metal2 51 -741 51 -741 0 net=2914
rlabel metal2 597 -741 597 -741 0 net=3501
rlabel metal2 639 -741 639 -741 0 net=2782
rlabel metal2 58 -743 58 -743 0 net=3442
rlabel metal2 681 -743 681 -743 0 net=4233
rlabel metal2 58 -745 58 -745 0 net=1463
rlabel metal2 341 -745 341 -745 0 net=4218
rlabel metal2 75 -747 75 -747 0 net=3217
rlabel metal2 660 -747 660 -747 0 net=2963
rlabel metal2 96 -749 96 -749 0 net=3239
rlabel metal2 100 -751 100 -751 0 net=971
rlabel metal2 100 -751 100 -751 0 net=971
rlabel metal2 117 -751 117 -751 0 net=3604
rlabel metal2 142 -753 142 -753 0 net=1761
rlabel metal2 240 -753 240 -753 0 net=584
rlabel metal2 79 -755 79 -755 0 net=1005
rlabel metal2 254 -755 254 -755 0 net=1143
rlabel metal2 289 -755 289 -755 0 net=3974
rlabel metal2 86 -757 86 -757 0 net=2280
rlabel metal2 282 -757 282 -757 0 net=1119
rlabel metal2 292 -757 292 -757 0 net=1326
rlabel metal2 506 -757 506 -757 0 net=2441
rlabel metal2 86 -759 86 -759 0 net=1059
rlabel metal2 275 -759 275 -759 0 net=2025
rlabel metal2 310 -759 310 -759 0 net=2363
rlabel metal2 583 -759 583 -759 0 net=3725
rlabel metal2 37 -761 37 -761 0 net=1453
rlabel metal2 324 -761 324 -761 0 net=1095
rlabel metal2 348 -761 348 -761 0 net=4253
rlabel metal2 37 -763 37 -763 0 net=4216
rlabel metal2 107 -765 107 -765 0 net=991
rlabel metal2 331 -765 331 -765 0 net=2126
rlabel metal2 366 -765 366 -765 0 net=2931
rlabel metal2 107 -767 107 -767 0 net=1381
rlabel metal2 548 -767 548 -767 0 net=3363
rlabel metal2 82 -769 82 -769 0 net=2637
rlabel metal2 590 -769 590 -769 0 net=3073
rlabel metal2 135 -771 135 -771 0 net=1101
rlabel metal2 296 -771 296 -771 0 net=1022
rlabel metal2 352 -771 352 -771 0 net=677
rlabel metal2 394 -771 394 -771 0 net=2372
rlabel metal2 600 -771 600 -771 0 net=3918
rlabel metal2 135 -773 135 -773 0 net=785
rlabel metal2 387 -773 387 -773 0 net=1849
rlabel metal2 408 -773 408 -773 0 net=2476
rlabel metal2 450 -773 450 -773 0 net=3116
rlabel metal2 709 -773 709 -773 0 net=3877
rlabel metal2 142 -775 142 -775 0 net=1113
rlabel metal2 191 -775 191 -775 0 net=823
rlabel metal2 191 -775 191 -775 0 net=823
rlabel metal2 226 -775 226 -775 0 net=722
rlabel metal2 408 -775 408 -775 0 net=2047
rlabel metal2 429 -775 429 -775 0 net=3434
rlabel metal2 611 -775 611 -775 0 net=3307
rlabel metal2 611 -775 611 -775 0 net=3307
rlabel metal2 632 -775 632 -775 0 net=3817
rlabel metal2 159 -777 159 -777 0 net=4058
rlabel metal2 163 -779 163 -779 0 net=1891
rlabel metal2 411 -779 411 -779 0 net=3216
rlabel metal2 639 -779 639 -779 0 net=4073
rlabel metal2 170 -781 170 -781 0 net=897
rlabel metal2 296 -781 296 -781 0 net=1305
rlabel metal2 446 -781 446 -781 0 net=3267
rlabel metal2 198 -783 198 -783 0 net=1427
rlabel metal2 380 -783 380 -783 0 net=1803
rlabel metal2 436 -783 436 -783 0 net=3492
rlabel metal2 16 -785 16 -785 0 net=2843
rlabel metal2 198 -787 198 -787 0 net=2293
rlabel metal2 380 -787 380 -787 0 net=3888
rlabel metal2 205 -789 205 -789 0 net=1249
rlabel metal2 359 -789 359 -789 0 net=1617
rlabel metal2 404 -789 404 -789 0 net=3059
rlabel metal2 23 -791 23 -791 0 net=1599
rlabel metal2 338 -791 338 -791 0 net=801
rlabel metal2 436 -791 436 -791 0 net=3829
rlabel metal2 23 -793 23 -793 0 net=1611
rlabel metal2 457 -793 457 -793 0 net=2261
rlabel metal2 492 -793 492 -793 0 net=2777
rlabel metal2 604 -793 604 -793 0 net=3257
rlabel metal2 93 -795 93 -795 0 net=1707
rlabel metal2 422 -795 422 -795 0 net=2085
rlabel metal2 471 -795 471 -795 0 net=2447
rlabel metal2 520 -795 520 -795 0 net=3001
rlabel metal2 625 -795 625 -795 0 net=3779
rlabel metal2 93 -797 93 -797 0 net=1492
rlabel metal2 453 -797 453 -797 0 net=4175
rlabel metal2 534 -797 534 -797 0 net=2595
rlabel metal2 562 -797 562 -797 0 net=2829
rlabel metal2 618 -797 618 -797 0 net=3451
rlabel metal2 16 -799 16 -799 0 net=2787
rlabel metal2 569 -799 569 -799 0 net=2945
rlabel metal2 646 -799 646 -799 0 net=3511
rlabel metal2 149 -801 149 -801 0 net=1819
rlabel metal2 499 -801 499 -801 0 net=2397
rlabel metal2 114 -803 114 -803 0 net=1547
rlabel metal2 261 -803 261 -803 0 net=755
rlabel metal2 478 -803 478 -803 0 net=2343
rlabel metal2 527 -803 527 -803 0 net=2537
rlabel metal2 555 -803 555 -803 0 net=2809
rlabel metal2 646 -803 646 -803 0 net=3107
rlabel metal2 177 -805 177 -805 0 net=2135
rlabel metal2 555 -805 555 -805 0 net=4080
rlabel metal2 128 -807 128 -807 0 net=1695
rlabel metal2 219 -807 219 -807 0 net=2239
rlabel metal2 758 -807 758 -807 0 net=4251
rlabel metal2 30 -809 30 -809 0 net=1045
rlabel metal2 219 -809 219 -809 0 net=1385
rlabel metal2 716 -809 716 -809 0 net=3947
rlabel metal2 30 -811 30 -811 0 net=1193
rlabel metal2 271 -811 271 -811 0 net=2987
rlabel metal2 303 -813 303 -813 0 net=1279
rlabel metal2 390 -813 390 -813 0 net=3629
rlabel metal2 9 -824 9 -824 0 net=2894
rlabel metal2 96 -824 96 -824 0 net=1006
rlabel metal2 303 -824 303 -824 0 net=2398
rlabel metal2 23 -826 23 -826 0 net=1612
rlabel metal2 54 -826 54 -826 0 net=435
rlabel metal2 369 -826 369 -826 0 net=3512
rlabel metal2 37 -828 37 -828 0 net=2844
rlabel metal2 37 -830 37 -830 0 net=174
rlabel metal2 331 -830 331 -830 0 net=3830
rlabel metal2 26 -832 26 -832 0 net=3381
rlabel metal2 348 -832 348 -832 0 net=2136
rlabel metal2 530 -832 530 -832 0 net=4234
rlabel metal2 51 -834 51 -834 0 net=1762
rlabel metal2 352 -834 352 -834 0 net=2442
rlabel metal2 58 -836 58 -836 0 net=1465
rlabel metal2 359 -836 359 -836 0 net=802
rlabel metal2 390 -836 390 -836 0 net=3074
rlabel metal2 58 -838 58 -838 0 net=825
rlabel metal2 212 -838 212 -838 0 net=1145
rlabel metal2 373 -838 373 -838 0 net=1618
rlabel metal2 404 -838 404 -838 0 net=2810
rlabel metal2 590 -838 590 -838 0 net=3364
rlabel metal2 709 -838 709 -838 0 net=3949
rlabel metal2 30 -840 30 -840 0 net=1195
rlabel metal2 257 -840 257 -840 0 net=2549
rlabel metal2 380 -840 380 -840 0 net=2831
rlabel metal2 625 -840 625 -840 0 net=3781
rlabel metal2 625 -840 625 -840 0 net=3781
rlabel metal2 632 -840 632 -840 0 net=3819
rlabel metal2 681 -840 681 -840 0 net=2965
rlabel metal2 30 -842 30 -842 0 net=973
rlabel metal2 128 -842 128 -842 0 net=1047
rlabel metal2 187 -842 187 -842 0 net=2026
rlabel metal2 306 -842 306 -842 0 net=2487
rlabel metal2 65 -844 65 -844 0 net=3218
rlabel metal2 65 -846 65 -846 0 net=933
rlabel metal2 72 -846 72 -846 0 net=1382
rlabel metal2 114 -846 114 -846 0 net=1549
rlabel metal2 145 -846 145 -846 0 net=3060
rlabel metal2 16 -848 16 -848 0 net=1509
rlabel metal2 149 -848 149 -848 0 net=1280
rlabel metal2 324 -848 324 -848 0 net=1097
rlabel metal2 394 -848 394 -848 0 net=1850
rlabel metal2 411 -848 411 -848 0 net=2932
rlabel metal2 716 -848 716 -848 0 net=3631
rlabel metal2 44 -850 44 -850 0 net=1923
rlabel metal2 44 -852 44 -852 0 net=1601
rlabel metal2 310 -852 310 -852 0 net=1455
rlabel metal2 338 -852 338 -852 0 net=3219
rlabel metal2 611 -852 611 -852 0 net=3309
rlabel metal2 72 -854 72 -854 0 net=2295
rlabel metal2 219 -854 219 -854 0 net=1387
rlabel metal2 394 -854 394 -854 0 net=2049
rlabel metal2 422 -854 422 -854 0 net=1821
rlabel metal2 82 -856 82 -856 0 net=2364
rlabel metal2 537 -856 537 -856 0 net=3452
rlabel metal2 86 -858 86 -858 0 net=1061
rlabel metal2 226 -858 226 -858 0 net=1429
rlabel metal2 422 -858 422 -858 0 net=2789
rlabel metal2 569 -858 569 -858 0 net=3259
rlabel metal2 86 -860 86 -860 0 net=1263
rlabel metal2 149 -860 149 -860 0 net=757
rlabel metal2 429 -860 429 -860 0 net=2262
rlabel metal2 555 -860 555 -860 0 net=4254
rlabel metal2 93 -862 93 -862 0 net=1115
rlabel metal2 152 -862 152 -862 0 net=1102
rlabel metal2 299 -862 299 -862 0 net=2735
rlabel metal2 436 -862 436 -862 0 net=3002
rlabel metal2 555 -862 555 -862 0 net=2989
rlabel metal2 632 -862 632 -862 0 net=4075
rlabel metal2 667 -862 667 -862 0 net=3879
rlabel metal2 107 -864 107 -864 0 net=2851
rlabel metal2 436 -864 436 -864 0 net=2241
rlabel metal2 485 -864 485 -864 0 net=2639
rlabel metal2 562 -864 562 -864 0 net=3241
rlabel metal2 121 -866 121 -866 0 net=899
rlabel metal2 173 -866 173 -866 0 net=1306
rlabel metal2 306 -866 306 -866 0 net=4195
rlabel metal2 513 -866 513 -866 0 net=4177
rlabel metal2 142 -868 142 -868 0 net=1775
rlabel metal2 275 -868 275 -868 0 net=419
rlabel metal2 450 -868 450 -868 0 net=3689
rlabel metal2 156 -870 156 -870 0 net=1709
rlabel metal2 163 -870 163 -870 0 net=1893
rlabel metal2 345 -870 345 -870 0 net=4111
rlabel metal2 156 -872 156 -872 0 net=1251
rlabel metal2 345 -872 345 -872 0 net=1805
rlabel metal2 443 -872 443 -872 0 net=2345
rlabel metal2 513 -872 513 -872 0 net=2947
rlabel metal2 117 -874 117 -874 0 net=4235
rlabel metal2 453 -874 453 -874 0 net=2778
rlabel metal2 597 -874 597 -874 0 net=3503
rlabel metal2 635 -874 635 -874 0 net=1
rlabel metal2 163 -876 163 -876 0 net=775
rlabel metal2 453 -876 453 -876 0 net=4252
rlabel metal2 170 -878 170 -878 0 net=74
rlabel metal2 457 -878 457 -878 0 net=2087
rlabel metal2 135 -880 135 -880 0 net=787
rlabel metal2 471 -880 471 -880 0 net=2449
rlabel metal2 471 -880 471 -880 0 net=2449
rlabel metal2 492 -880 492 -880 0 net=2597
rlabel metal2 135 -882 135 -882 0 net=2469
rlabel metal2 268 -882 268 -882 0 net=1121
rlabel metal2 541 -882 541 -882 0 net=3109
rlabel metal2 79 -884 79 -884 0 net=1897
rlabel metal2 583 -884 583 -884 0 net=3727
rlabel metal2 177 -886 177 -886 0 net=1697
rlabel metal2 583 -886 583 -886 0 net=3269
rlabel metal2 177 -888 177 -888 0 net=992
rlabel metal2 674 -888 674 -888 0 net=4123
rlabel metal2 180 -890 180 -890 0 net=1679
rlabel metal2 233 -892 233 -892 0 net=1157
rlabel metal2 366 -894 366 -894 0 net=2095
rlabel metal2 464 -896 464 -896 0 net=2539
rlabel metal2 534 -898 534 -898 0 net=4159
rlabel metal2 2 -909 2 -909 0 net=1979
rlabel metal2 103 -909 103 -909 0 net=1158
rlabel metal2 240 -909 240 -909 0 net=1466
rlabel metal2 317 -909 317 -909 0 net=1895
rlabel metal2 317 -909 317 -909 0 net=1895
rlabel metal2 338 -909 338 -909 0 net=1699
rlabel metal2 359 -909 359 -909 0 net=42
rlabel metal2 548 -909 548 -909 0 net=3243
rlabel metal2 576 -909 576 -909 0 net=3220
rlabel metal2 607 -909 607 -909 0 net=3310
rlabel metal2 695 -909 695 -909 0 net=2966
rlabel metal2 23 -911 23 -911 0 net=2088
rlabel metal2 509 -911 509 -911 0 net=4076
rlabel metal2 737 -911 737 -911 0 net=3633
rlabel metal2 26 -913 26 -913 0 net=1983
rlabel metal2 205 -913 205 -913 0 net=1710
rlabel metal2 257 -913 257 -913 0 net=3199
rlabel metal2 30 -915 30 -915 0 net=974
rlabel metal2 205 -915 205 -915 0 net=1361
rlabel metal2 404 -915 404 -915 0 net=3728
rlabel metal2 30 -917 30 -917 0 net=1309
rlabel metal2 212 -917 212 -917 0 net=1146
rlabel metal2 296 -917 296 -917 0 net=1389
rlabel metal2 383 -917 383 -917 0 net=2050
rlabel metal2 408 -917 408 -917 0 net=4219
rlabel metal2 618 -917 618 -917 0 net=3691
rlabel metal2 37 -919 37 -919 0 net=1181
rlabel metal2 54 -919 54 -919 0 net=2488
rlabel metal2 40 -921 40 -921 0 net=1924
rlabel metal2 65 -923 65 -923 0 net=934
rlabel metal2 156 -923 156 -923 0 net=1253
rlabel metal2 229 -923 229 -923 0 net=3413
rlabel metal2 597 -923 597 -923 0 net=4161
rlabel metal2 65 -925 65 -925 0 net=2990
rlabel metal2 576 -925 576 -925 0 net=3505
rlabel metal2 621 -925 621 -925 0 net=3950
rlabel metal2 72 -927 72 -927 0 net=2297
rlabel metal2 275 -927 275 -927 0 net=4171
rlabel metal2 72 -929 72 -929 0 net=2097
rlabel metal2 387 -929 387 -929 0 net=1098
rlabel metal2 478 -929 478 -929 0 net=4197
rlabel metal2 79 -931 79 -931 0 net=1898
rlabel metal2 219 -931 219 -931 0 net=1777
rlabel metal2 394 -931 394 -931 0 net=4178
rlabel metal2 688 -931 688 -931 0 net=4149
rlabel metal2 61 -933 61 -933 0 net=1519
rlabel metal2 86 -933 86 -933 0 net=1264
rlabel metal2 275 -933 275 -933 0 net=1807
rlabel metal2 362 -933 362 -933 0 net=4081
rlabel metal2 93 -935 93 -935 0 net=1116
rlabel metal2 156 -935 156 -935 0 net=777
rlabel metal2 226 -935 226 -935 0 net=2471
rlabel metal2 415 -935 415 -935 0 net=4237
rlabel metal2 93 -937 93 -937 0 net=1063
rlabel metal2 233 -937 233 -937 0 net=2553
rlabel metal2 303 -937 303 -937 0 net=1477
rlabel metal2 436 -937 436 -937 0 net=2243
rlabel metal2 436 -937 436 -937 0 net=2243
rlabel metal2 450 -937 450 -937 0 net=2451
rlabel metal2 478 -937 478 -937 0 net=3075
rlabel metal2 534 -937 534 -937 0 net=3261
rlabel metal2 625 -937 625 -937 0 net=3783
rlabel metal2 44 -939 44 -939 0 net=1603
rlabel metal2 240 -939 240 -939 0 net=1123
rlabel metal2 278 -939 278 -939 0 net=1456
rlabel metal2 499 -939 499 -939 0 net=3669
rlabel metal2 44 -941 44 -941 0 net=3009
rlabel metal2 625 -941 625 -941 0 net=3821
rlabel metal2 107 -943 107 -943 0 net=2852
rlabel metal2 513 -943 513 -943 0 net=2949
rlabel metal2 555 -943 555 -943 0 net=4125
rlabel metal2 107 -945 107 -945 0 net=1769
rlabel metal2 513 -945 513 -945 0 net=3271
rlabel metal2 114 -947 114 -947 0 net=1551
rlabel metal2 135 -947 135 -947 0 net=2557
rlabel metal2 520 -947 520 -947 0 net=4113
rlabel metal2 16 -949 16 -949 0 net=1511
rlabel metal2 163 -949 163 -949 0 net=1293
rlabel metal2 261 -949 261 -949 0 net=1681
rlabel metal2 520 -949 520 -949 0 net=3111
rlabel metal2 562 -949 562 -949 0 net=3281
rlabel metal2 16 -951 16 -951 0 net=1197
rlabel metal2 261 -951 261 -951 0 net=1225
rlabel metal2 100 -953 100 -953 0 net=1569
rlabel metal2 149 -953 149 -953 0 net=759
rlabel metal2 282 -953 282 -953 0 net=2599
rlabel metal2 117 -955 117 -955 0 net=1430
rlabel metal2 285 -955 285 -955 0 net=2790
rlabel metal2 485 -955 485 -955 0 net=2641
rlabel metal2 121 -957 121 -957 0 net=901
rlabel metal2 310 -957 310 -957 0 net=1822
rlabel metal2 58 -959 58 -959 0 net=827
rlabel metal2 142 -959 142 -959 0 net=2231
rlabel metal2 653 -959 653 -959 0 net=3881
rlabel metal2 9 -961 9 -961 0 net=369
rlabel metal2 149 -961 149 -961 0 net=2215
rlabel metal2 180 -963 180 -963 0 net=788
rlabel metal2 324 -965 324 -965 0 net=869
rlabel metal2 313 -967 313 -967 0 net=2873
rlabel metal2 331 -969 331 -969 0 net=3383
rlabel metal2 51 -971 51 -971 0 net=1619
rlabel metal2 373 -971 373 -971 0 net=2551
rlabel metal2 184 -973 184 -973 0 net=1049
rlabel metal2 401 -973 401 -973 0 net=4091
rlabel metal2 184 -975 184 -975 0 net=3653
rlabel metal2 401 -975 401 -975 0 net=2205
rlabel metal2 457 -975 457 -975 0 net=2541
rlabel metal2 429 -977 429 -977 0 net=2737
rlabel metal2 429 -979 429 -979 0 net=2347
rlabel metal2 380 -981 380 -981 0 net=2832
rlabel metal2 9 -992 9 -992 0 net=630
rlabel metal2 187 -992 187 -992 0 net=2298
rlabel metal2 275 -992 275 -992 0 net=1808
rlabel metal2 404 -992 404 -992 0 net=2244
rlabel metal2 443 -992 443 -992 0 net=2453
rlabel metal2 464 -992 464 -992 0 net=2738
rlabel metal2 499 -992 499 -992 0 net=2875
rlabel metal2 520 -992 520 -992 0 net=3113
rlabel metal2 527 -992 527 -992 0 net=2951
rlabel metal2 751 -992 751 -992 0 net=3635
rlabel metal2 26 -994 26 -994 0 net=2235
rlabel metal2 79 -994 79 -994 0 net=1520
rlabel metal2 89 -994 89 -994 0 net=4220
rlabel metal2 618 -994 618 -994 0 net=3693
rlabel metal2 639 -994 639 -994 0 net=3785
rlabel metal2 639 -994 639 -994 0 net=3785
rlabel metal2 653 -994 653 -994 0 net=3883
rlabel metal2 653 -994 653 -994 0 net=3883
rlabel metal2 716 -994 716 -994 0 net=4239
rlabel metal2 30 -996 30 -996 0 net=1310
rlabel metal2 425 -996 425 -996 0 net=3079
rlabel metal2 548 -996 548 -996 0 net=3245
rlabel metal2 548 -996 548 -996 0 net=3245
rlabel metal2 604 -996 604 -996 0 net=662
rlabel metal2 625 -996 625 -996 0 net=3823
rlabel metal2 709 -996 709 -996 0 net=4199
rlabel metal2 37 -998 37 -998 0 net=1182
rlabel metal2 149 -998 149 -998 0 net=410
rlabel metal2 436 -998 436 -998 0 net=2543
rlabel metal2 464 -998 464 -998 0 net=2643
rlabel metal2 502 -998 502 -998 0 net=3506
rlabel metal2 695 -998 695 -998 0 net=4163
rlabel metal2 37 -1000 37 -1000 0 net=2099
rlabel metal2 79 -1000 79 -1000 0 net=2349
rlabel metal2 457 -1000 457 -1000 0 net=2559
rlabel metal2 478 -1000 478 -1000 0 net=3077
rlabel metal2 520 -1000 520 -1000 0 net=3283
rlabel metal2 695 -1000 695 -1000 0 net=4173
rlabel metal2 44 -1002 44 -1002 0 net=3200
rlabel metal2 688 -1002 688 -1002 0 net=4151
rlabel metal2 47 -1004 47 -1004 0 net=1604
rlabel metal2 205 -1004 205 -1004 0 net=1362
rlabel metal2 485 -1004 485 -1004 0 net=2759
rlabel metal2 674 -1004 674 -1004 0 net=4115
rlabel metal2 54 -1006 54 -1006 0 net=3010
rlabel metal2 660 -1006 660 -1006 0 net=4083
rlabel metal2 58 -1008 58 -1008 0 net=2217
rlabel metal2 488 -1008 488 -1008 0 net=3771
rlabel metal2 660 -1008 660 -1008 0 net=4093
rlabel metal2 68 -1010 68 -1010 0 net=2477
rlabel metal2 569 -1010 569 -1010 0 net=3385
rlabel metal2 86 -1012 86 -1012 0 net=1621
rlabel metal2 352 -1012 352 -1012 0 net=1771
rlabel metal2 555 -1012 555 -1012 0 net=4127
rlabel metal2 93 -1014 93 -1014 0 net=1064
rlabel metal2 191 -1014 191 -1014 0 net=761
rlabel metal2 205 -1014 205 -1014 0 net=1683
rlabel metal2 366 -1014 366 -1014 0 net=1779
rlabel metal2 2 -1016 2 -1016 0 net=1981
rlabel metal2 366 -1016 366 -1016 0 net=3641
rlabel metal2 383 -1016 383 -1016 0 net=2723
rlabel metal2 534 -1016 534 -1016 0 net=3263
rlabel metal2 93 -1018 93 -1018 0 net=1571
rlabel metal2 107 -1018 107 -1018 0 net=3670
rlabel metal2 16 -1020 16 -1020 0 net=1199
rlabel metal2 114 -1020 114 -1020 0 net=1553
rlabel metal2 292 -1020 292 -1020 0 net=4201
rlabel metal2 16 -1022 16 -1022 0 net=1985
rlabel metal2 180 -1022 180 -1022 0 net=1050
rlabel metal2 394 -1022 394 -1022 0 net=2552
rlabel metal2 100 -1024 100 -1024 0 net=1254
rlabel metal2 219 -1024 219 -1024 0 net=902
rlabel metal2 240 -1024 240 -1024 0 net=1124
rlabel metal2 317 -1024 317 -1024 0 net=1896
rlabel metal2 373 -1024 373 -1024 0 net=3272
rlabel metal2 534 -1024 534 -1024 0 net=3415
rlabel metal2 23 -1026 23 -1026 0 net=3567
rlabel metal2 75 -1028 75 -1028 0 net=1481
rlabel metal2 247 -1028 247 -1028 0 net=1227
rlabel metal2 268 -1028 268 -1028 0 net=3655
rlabel metal2 117 -1030 117 -1030 0 net=2319
rlabel metal2 226 -1030 226 -1030 0 net=871
rlabel metal2 331 -1030 331 -1030 0 net=3421
rlabel metal2 142 -1032 142 -1032 0 net=2207
rlabel metal2 156 -1034 156 -1034 0 net=778
rlabel metal2 177 -1034 177 -1034 0 net=3227
rlabel metal2 128 -1036 128 -1036 0 net=1513
rlabel metal2 212 -1036 212 -1036 0 net=1721
rlabel metal2 317 -1036 317 -1036 0 net=1700
rlabel metal2 401 -1036 401 -1036 0 net=4005
rlabel metal2 103 -1038 103 -1038 0 net=1131
rlabel metal2 135 -1038 135 -1038 0 net=745
rlabel metal2 163 -1038 163 -1038 0 net=1295
rlabel metal2 250 -1038 250 -1038 0 net=3801
rlabel metal2 121 -1040 121 -1040 0 net=829
rlabel metal2 254 -1040 254 -1040 0 net=2233
rlabel metal2 30 -1042 30 -1042 0 net=2633
rlabel metal2 135 -1042 135 -1042 0 net=935
rlabel metal2 261 -1042 261 -1042 0 net=1391
rlabel metal2 306 -1042 306 -1042 0 net=1957
rlabel metal2 422 -1042 422 -1042 0 net=2967
rlabel metal2 233 -1044 233 -1044 0 net=2555
rlabel metal2 310 -1044 310 -1044 0 net=3729
rlabel metal2 233 -1046 233 -1046 0 net=1191
rlabel metal2 268 -1048 268 -1048 0 net=2417
rlabel metal2 275 -1050 275 -1050 0 net=1479
rlabel metal2 320 -1050 320 -1050 0 net=2472
rlabel metal2 282 -1052 282 -1052 0 net=2600
rlabel metal2 303 -1054 303 -1054 0 net=2865
rlabel metal2 324 -1056 324 -1056 0 net=2717
rlabel metal2 387 -1056 387 -1056 0 net=2429
rlabel metal2 16 -1067 16 -1067 0 net=1987
rlabel metal2 362 -1067 362 -1067 0 net=4174
rlabel metal2 702 -1067 702 -1067 0 net=4153
rlabel metal2 702 -1067 702 -1067 0 net=4153
rlabel metal2 730 -1067 730 -1067 0 net=2952
rlabel metal2 751 -1067 751 -1067 0 net=653
rlabel metal2 758 -1067 758 -1067 0 net=3637
rlabel metal2 758 -1067 758 -1067 0 net=3637
rlabel metal2 16 -1069 16 -1069 0 net=1393
rlabel metal2 268 -1069 268 -1069 0 net=1555
rlabel metal2 306 -1069 306 -1069 0 net=4128
rlabel metal2 754 -1069 754 -1069 0 net=3479
rlabel metal2 26 -1071 26 -1071 0 net=1622
rlabel metal2 89 -1071 89 -1071 0 net=670
rlabel metal2 177 -1071 177 -1071 0 net=1515
rlabel metal2 310 -1071 310 -1071 0 net=1982
rlabel metal2 369 -1071 369 -1071 0 net=3246
rlabel metal2 597 -1071 597 -1071 0 net=4203
rlabel metal2 9 -1073 9 -1073 0 net=694
rlabel metal2 93 -1073 93 -1073 0 net=1573
rlabel metal2 93 -1073 93 -1073 0 net=1573
rlabel metal2 107 -1073 107 -1073 0 net=1200
rlabel metal2 310 -1073 310 -1073 0 net=2719
rlabel metal2 327 -1073 327 -1073 0 net=2507
rlabel metal2 383 -1073 383 -1073 0 net=3078
rlabel metal2 509 -1073 509 -1073 0 net=4031
rlabel metal2 9 -1075 9 -1075 0 net=2635
rlabel metal2 156 -1075 156 -1075 0 net=746
rlabel metal2 205 -1075 205 -1075 0 net=1684
rlabel metal2 394 -1075 394 -1075 0 net=3645
rlabel metal2 464 -1075 464 -1075 0 net=2645
rlabel metal2 30 -1077 30 -1077 0 net=1772
rlabel metal2 474 -1077 474 -1077 0 net=3772
rlabel metal2 604 -1077 604 -1077 0 net=3884
rlabel metal2 660 -1077 660 -1077 0 net=4095
rlabel metal2 37 -1079 37 -1079 0 net=2100
rlabel metal2 156 -1079 156 -1079 0 net=735
rlabel metal2 170 -1079 170 -1079 0 net=1673
rlabel metal2 331 -1079 331 -1079 0 net=3423
rlabel metal2 632 -1079 632 -1079 0 net=3825
rlabel metal2 667 -1079 667 -1079 0 net=4007
rlabel metal2 44 -1081 44 -1081 0 net=2321
rlabel metal2 226 -1081 226 -1081 0 net=873
rlabel metal2 226 -1081 226 -1081 0 net=873
rlabel metal2 247 -1081 247 -1081 0 net=1228
rlabel metal2 418 -1081 418 -1081 0 net=4240
rlabel metal2 47 -1083 47 -1083 0 net=2236
rlabel metal2 72 -1083 72 -1083 0 net=1077
rlabel metal2 138 -1083 138 -1083 0 net=1780
rlabel metal2 625 -1083 625 -1083 0 net=3731
rlabel metal2 709 -1083 709 -1083 0 net=4165
rlabel metal2 23 -1085 23 -1085 0 net=1823
rlabel metal2 100 -1085 100 -1085 0 net=2513
rlabel metal2 198 -1085 198 -1085 0 net=763
rlabel metal2 250 -1085 250 -1085 0 net=1480
rlabel metal2 345 -1085 345 -1085 0 net=2301
rlabel metal2 450 -1085 450 -1085 0 net=3035
rlabel metal2 632 -1085 632 -1085 0 net=4085
rlabel metal2 688 -1085 688 -1085 0 net=4117
rlabel metal2 58 -1087 58 -1087 0 net=2219
rlabel metal2 114 -1087 114 -1087 0 net=1296
rlabel metal2 208 -1087 208 -1087 0 net=2234
rlabel metal2 275 -1087 275 -1087 0 net=1959
rlabel metal2 380 -1087 380 -1087 0 net=3643
rlabel metal2 639 -1087 639 -1087 0 net=3787
rlabel metal2 58 -1089 58 -1089 0 net=2209
rlabel metal2 163 -1089 163 -1089 0 net=831
rlabel metal2 380 -1089 380 -1089 0 net=144
rlabel metal2 114 -1091 114 -1091 0 net=1722
rlabel metal2 387 -1091 387 -1091 0 net=2431
rlabel metal2 425 -1091 425 -1091 0 net=4200
rlabel metal2 79 -1093 79 -1093 0 net=2351
rlabel metal2 397 -1093 397 -1093 0 net=3403
rlabel metal2 611 -1093 611 -1093 0 net=3657
rlabel metal2 646 -1093 646 -1093 0 net=3803
rlabel metal2 117 -1095 117 -1095 0 net=2556
rlabel metal2 401 -1095 401 -1095 0 net=2419
rlabel metal2 436 -1095 436 -1095 0 net=2545
rlabel metal2 457 -1095 457 -1095 0 net=2561
rlabel metal2 471 -1095 471 -1095 0 net=4129
rlabel metal2 51 -1097 51 -1097 0 net=2747
rlabel metal2 499 -1097 499 -1097 0 net=2877
rlabel metal2 51 -1099 51 -1099 0 net=2601
rlabel metal2 212 -1099 212 -1099 0 net=751
rlabel metal2 436 -1099 436 -1099 0 net=3114
rlabel metal2 618 -1099 618 -1099 0 net=3695
rlabel metal2 37 -1101 37 -1101 0 net=1001
rlabel metal2 513 -1101 513 -1101 0 net=2969
rlabel metal2 562 -1101 562 -1101 0 net=3387
rlabel metal2 103 -1103 103 -1103 0 net=2905
rlabel metal2 520 -1103 520 -1103 0 net=3285
rlabel metal2 520 -1103 520 -1103 0 net=3285
rlabel metal2 534 -1103 534 -1103 0 net=3417
rlabel metal2 121 -1105 121 -1105 0 net=723
rlabel metal2 527 -1105 527 -1105 0 net=3081
rlabel metal2 541 -1105 541 -1105 0 net=3229
rlabel metal2 541 -1105 541 -1105 0 net=3229
rlabel metal2 128 -1107 128 -1107 0 net=1133
rlabel metal2 163 -1107 163 -1107 0 net=2478
rlabel metal2 527 -1107 527 -1107 0 net=3265
rlabel metal2 128 -1109 128 -1109 0 net=937
rlabel metal2 177 -1109 177 -1109 0 net=75
rlabel metal2 289 -1109 289 -1109 0 net=3367
rlabel metal2 79 -1111 79 -1111 0 net=733
rlabel metal2 180 -1111 180 -1111 0 net=669
rlabel metal2 429 -1111 429 -1111 0 net=2725
rlabel metal2 555 -1111 555 -1111 0 net=3569
rlabel metal2 184 -1113 184 -1113 0 net=1147
rlabel metal2 240 -1113 240 -1113 0 net=1483
rlabel metal2 366 -1113 366 -1113 0 net=3437
rlabel metal2 184 -1115 184 -1115 0 net=1192
rlabel metal2 240 -1115 240 -1115 0 net=927
rlabel metal2 282 -1115 282 -1115 0 net=1711
rlabel metal2 366 -1115 366 -1115 0 net=2991
rlabel metal2 191 -1117 191 -1117 0 net=1493
rlabel metal2 429 -1117 429 -1117 0 net=2454
rlabel metal2 194 -1119 194 -1119 0 net=1321
rlabel metal2 443 -1119 443 -1119 0 net=2867
rlabel metal2 233 -1121 233 -1121 0 net=2573
rlabel metal2 485 -1121 485 -1121 0 net=2761
rlabel metal2 320 -1123 320 -1123 0 net=3455
rlabel metal2 9 -1134 9 -1134 0 net=2636
rlabel metal2 348 -1134 348 -1134 0 net=2479
rlabel metal2 509 -1134 509 -1134 0 net=4154
rlabel metal2 716 -1134 716 -1134 0 net=4131
rlabel metal2 793 -1134 793 -1134 0 net=3481
rlabel metal2 9 -1136 9 -1136 0 net=1039
rlabel metal2 310 -1136 310 -1136 0 net=2720
rlabel metal2 355 -1136 355 -1136 0 net=2508
rlabel metal2 422 -1136 422 -1136 0 net=1403
rlabel metal2 646 -1136 646 -1136 0 net=3697
rlabel metal2 740 -1136 740 -1136 0 net=2127
rlabel metal2 23 -1138 23 -1138 0 net=1713
rlabel metal2 366 -1138 366 -1138 0 net=2970
rlabel metal2 555 -1138 555 -1138 0 net=3571
rlabel metal2 26 -1140 26 -1140 0 net=3658
rlabel metal2 744 -1140 744 -1140 0 net=4009
rlabel metal2 30 -1142 30 -1142 0 net=3424
rlabel metal2 723 -1142 723 -1142 0 net=4167
rlabel metal2 37 -1144 37 -1144 0 net=1002
rlabel metal2 194 -1144 194 -1144 0 net=832
rlabel metal2 341 -1144 341 -1144 0 net=3663
rlabel metal2 674 -1144 674 -1144 0 net=3805
rlabel metal2 751 -1144 751 -1144 0 net=3638
rlabel metal2 44 -1146 44 -1146 0 net=2322
rlabel metal2 373 -1146 373 -1146 0 net=2993
rlabel metal2 520 -1146 520 -1146 0 net=3287
rlabel metal2 44 -1148 44 -1148 0 net=1353
rlabel metal2 432 -1148 432 -1148 0 net=3797
rlabel metal2 54 -1150 54 -1150 0 net=2748
rlabel metal2 467 -1150 467 -1150 0 net=2762
rlabel metal2 534 -1150 534 -1150 0 net=3083
rlabel metal2 632 -1150 632 -1150 0 net=4087
rlabel metal2 72 -1152 72 -1152 0 net=1078
rlabel metal2 254 -1152 254 -1152 0 net=1323
rlabel metal2 324 -1152 324 -1152 0 net=236
rlabel metal2 394 -1152 394 -1152 0 net=3647
rlabel metal2 695 -1152 695 -1152 0 net=4097
rlabel metal2 79 -1154 79 -1154 0 net=734
rlabel metal2 331 -1154 331 -1154 0 net=1371
rlabel metal2 397 -1154 397 -1154 0 net=3929
rlabel metal2 562 -1154 562 -1154 0 net=3389
rlabel metal2 79 -1156 79 -1156 0 net=1135
rlabel metal2 145 -1156 145 -1156 0 net=259
rlabel metal2 212 -1156 212 -1156 0 net=752
rlabel metal2 247 -1156 247 -1156 0 net=1735
rlabel metal2 275 -1156 275 -1156 0 net=1961
rlabel metal2 443 -1156 443 -1156 0 net=2869
rlabel metal2 569 -1156 569 -1156 0 net=3368
rlabel metal2 16 -1158 16 -1158 0 net=1394
rlabel metal2 292 -1158 292 -1158 0 net=1007
rlabel metal2 401 -1158 401 -1158 0 net=2421
rlabel metal2 541 -1158 541 -1158 0 net=3231
rlabel metal2 16 -1160 16 -1160 0 net=993
rlabel metal2 166 -1160 166 -1160 0 net=247
rlabel metal2 187 -1160 187 -1160 0 net=2143
rlabel metal2 474 -1160 474 -1160 0 net=3266
rlabel metal2 548 -1160 548 -1160 0 net=2647
rlabel metal2 100 -1162 100 -1162 0 net=2515
rlabel metal2 569 -1162 569 -1162 0 net=2879
rlabel metal2 93 -1164 93 -1164 0 net=1575
rlabel metal2 107 -1164 107 -1164 0 net=2221
rlabel metal2 107 -1164 107 -1164 0 net=2221
rlabel metal2 114 -1164 114 -1164 0 net=4032
rlabel metal2 730 -1164 730 -1164 0 net=4205
rlabel metal2 93 -1166 93 -1166 0 net=1281
rlabel metal2 408 -1166 408 -1166 0 net=2575
rlabel metal2 576 -1166 576 -1166 0 net=3419
rlabel metal2 653 -1166 653 -1166 0 net=3827
rlabel metal2 117 -1168 117 -1168 0 net=2313
rlabel metal2 352 -1168 352 -1168 0 net=3717
rlabel metal2 117 -1170 117 -1170 0 net=921
rlabel metal2 198 -1170 198 -1170 0 net=1149
rlabel metal2 296 -1170 296 -1170 0 net=1485
rlabel metal2 359 -1170 359 -1170 0 net=1989
rlabel metal2 450 -1170 450 -1170 0 net=2547
rlabel metal2 590 -1170 590 -1170 0 net=3439
rlabel metal2 121 -1172 121 -1172 0 net=725
rlabel metal2 152 -1172 152 -1172 0 net=3404
rlabel metal2 625 -1172 625 -1172 0 net=3037
rlabel metal2 121 -1174 121 -1174 0 net=939
rlabel metal2 135 -1174 135 -1174 0 net=2925
rlabel metal2 625 -1174 625 -1174 0 net=3789
rlabel metal2 51 -1176 51 -1176 0 net=2603
rlabel metal2 138 -1176 138 -1176 0 net=267
rlabel metal2 429 -1176 429 -1176 0 net=1943
rlabel metal2 485 -1176 485 -1176 0 net=3457
rlabel metal2 33 -1178 33 -1178 0 net=1793
rlabel metal2 499 -1178 499 -1178 0 net=2907
rlabel metal2 51 -1180 51 -1180 0 net=29
rlabel metal2 58 -1182 58 -1182 0 net=2211
rlabel metal2 156 -1182 156 -1182 0 net=737
rlabel metal2 156 -1182 156 -1182 0 net=737
rlabel metal2 170 -1182 170 -1182 0 net=1675
rlabel metal2 170 -1182 170 -1182 0 net=1675
rlabel metal2 177 -1182 177 -1182 0 net=1035
rlabel metal2 415 -1182 415 -1182 0 net=2433
rlabel metal2 58 -1184 58 -1184 0 net=1899
rlabel metal2 198 -1184 198 -1184 0 net=1517
rlabel metal2 296 -1184 296 -1184 0 net=1187
rlabel metal2 450 -1184 450 -1184 0 net=2727
rlabel metal2 65 -1186 65 -1186 0 net=1825
rlabel metal2 464 -1186 464 -1186 0 net=2563
rlabel metal2 65 -1188 65 -1188 0 net=841
rlabel metal2 205 -1188 205 -1188 0 net=857
rlabel metal2 471 -1188 471 -1188 0 net=3644
rlabel metal2 212 -1190 212 -1190 0 net=929
rlabel metal2 250 -1190 250 -1190 0 net=3049
rlabel metal2 226 -1192 226 -1192 0 net=874
rlabel metal2 240 -1192 240 -1192 0 net=1327
rlabel metal2 219 -1194 219 -1194 0 net=765
rlabel metal2 261 -1194 261 -1194 0 net=1557
rlabel metal2 303 -1194 303 -1194 0 net=1495
rlabel metal2 369 -1194 369 -1194 0 net=2352
rlabel metal2 40 -1196 40 -1196 0 net=1079
rlabel metal2 268 -1196 268 -1196 0 net=1467
rlabel metal2 303 -1198 303 -1198 0 net=2303
rlabel metal2 345 -1200 345 -1200 0 net=3732
rlabel metal2 667 -1202 667 -1202 0 net=4119
rlabel metal2 478 -1204 478 -1204 0 net=3793
rlabel metal2 2 -1215 2 -1215 0 net=2213
rlabel metal2 149 -1215 149 -1215 0 net=727
rlabel metal2 149 -1215 149 -1215 0 net=727
rlabel metal2 156 -1215 156 -1215 0 net=739
rlabel metal2 156 -1215 156 -1215 0 net=739
rlabel metal2 184 -1215 184 -1215 0 net=1518
rlabel metal2 254 -1215 254 -1215 0 net=1324
rlabel metal2 317 -1215 317 -1215 0 net=1990
rlabel metal2 471 -1215 471 -1215 0 net=2481
rlabel metal2 541 -1215 541 -1215 0 net=3440
rlabel metal2 649 -1215 649 -1215 0 net=4206
rlabel metal2 789 -1215 789 -1215 0 net=3482
rlabel metal2 9 -1217 9 -1217 0 net=1040
rlabel metal2 362 -1217 362 -1217 0 net=3664
rlabel metal2 660 -1217 660 -1217 0 net=2701
rlabel metal2 9 -1219 9 -1219 0 net=1337
rlabel metal2 33 -1219 33 -1219 0 net=182
rlabel metal2 667 -1219 667 -1219 0 net=4121
rlabel metal2 16 -1221 16 -1221 0 net=994
rlabel metal2 100 -1221 100 -1221 0 net=1577
rlabel metal2 100 -1221 100 -1221 0 net=1577
rlabel metal2 128 -1221 128 -1221 0 net=2605
rlabel metal2 397 -1221 397 -1221 0 net=2548
rlabel metal2 593 -1221 593 -1221 0 net=3828
rlabel metal2 16 -1223 16 -1223 0 net=2001
rlabel metal2 198 -1223 198 -1223 0 net=1008
rlabel metal2 387 -1223 387 -1223 0 net=2577
rlabel metal2 681 -1223 681 -1223 0 net=3039
rlabel metal2 30 -1225 30 -1225 0 net=2699
rlabel metal2 254 -1225 254 -1225 0 net=1163
rlabel metal2 345 -1225 345 -1225 0 net=1794
rlabel metal2 506 -1225 506 -1225 0 net=3085
rlabel metal2 37 -1227 37 -1227 0 net=1469
rlabel metal2 278 -1227 278 -1227 0 net=4139
rlabel metal2 23 -1229 23 -1229 0 net=1715
rlabel metal2 282 -1229 282 -1229 0 net=2315
rlabel metal2 366 -1229 366 -1229 0 net=2434
rlabel metal2 520 -1229 520 -1229 0 net=2909
rlabel metal2 23 -1231 23 -1231 0 net=1081
rlabel metal2 247 -1231 247 -1231 0 net=1737
rlabel metal2 555 -1231 555 -1231 0 net=3931
rlabel metal2 51 -1233 51 -1233 0 net=1900
rlabel metal2 68 -1233 68 -1233 0 net=842
rlabel metal2 75 -1233 75 -1233 0 net=1962
rlabel metal2 443 -1233 443 -1233 0 net=2423
rlabel metal2 555 -1233 555 -1233 0 net=3459
rlabel metal2 51 -1235 51 -1235 0 net=941
rlabel metal2 128 -1235 128 -1235 0 net=1763
rlabel metal2 373 -1235 373 -1235 0 net=2995
rlabel metal2 576 -1235 576 -1235 0 net=3051
rlabel metal2 653 -1235 653 -1235 0 net=3699
rlabel metal2 54 -1237 54 -1237 0 net=3057
rlabel metal2 688 -1237 688 -1237 0 net=4099
rlabel metal2 58 -1239 58 -1239 0 net=1329
rlabel metal2 247 -1239 247 -1239 0 net=1151
rlabel metal2 317 -1239 317 -1239 0 net=1405
rlabel metal2 464 -1239 464 -1239 0 net=3193
rlabel metal2 758 -1239 758 -1239 0 net=4169
rlabel metal2 79 -1241 79 -1241 0 net=1136
rlabel metal2 145 -1241 145 -1241 0 net=922
rlabel metal2 212 -1241 212 -1241 0 net=931
rlabel metal2 240 -1241 240 -1241 0 net=1487
rlabel metal2 373 -1241 373 -1241 0 net=1945
rlabel metal2 464 -1241 464 -1241 0 net=2517
rlabel metal2 79 -1243 79 -1243 0 net=1373
rlabel metal2 334 -1243 334 -1243 0 net=3687
rlabel metal2 86 -1245 86 -1245 0 net=1497
rlabel metal2 390 -1245 390 -1245 0 net=3390
rlabel metal2 93 -1247 93 -1247 0 net=1283
rlabel metal2 135 -1247 135 -1247 0 net=859
rlabel metal2 212 -1247 212 -1247 0 net=1827
rlabel metal2 422 -1247 422 -1247 0 net=2728
rlabel metal2 478 -1247 478 -1247 0 net=4088
rlabel metal2 93 -1249 93 -1249 0 net=1037
rlabel metal2 184 -1249 184 -1249 0 net=2527
rlabel metal2 450 -1249 450 -1249 0 net=3897
rlabel metal2 44 -1251 44 -1251 0 net=1355
rlabel metal2 191 -1251 191 -1251 0 net=2305
rlabel metal2 324 -1251 324 -1251 0 net=3806
rlabel metal2 44 -1253 44 -1253 0 net=1449
rlabel metal2 107 -1253 107 -1253 0 net=2223
rlabel metal2 324 -1253 324 -1253 0 net=2145
rlabel metal2 478 -1253 478 -1253 0 net=2565
rlabel metal2 632 -1253 632 -1253 0 net=3679
rlabel metal2 107 -1255 107 -1255 0 net=1677
rlabel metal2 205 -1255 205 -1255 0 net=767
rlabel metal2 282 -1255 282 -1255 0 net=3401
rlabel metal2 401 -1255 401 -1255 0 net=2648
rlabel metal2 723 -1255 723 -1255 0 net=4011
rlabel metal2 65 -1257 65 -1257 0 net=1395
rlabel metal2 341 -1257 341 -1257 0 net=2870
rlabel metal2 744 -1257 744 -1257 0 net=4133
rlabel metal2 114 -1259 114 -1259 0 net=4145
rlabel metal2 772 -1259 772 -1259 0 net=2128
rlabel metal2 166 -1261 166 -1261 0 net=2281
rlabel metal2 401 -1261 401 -1261 0 net=3572
rlabel metal2 310 -1263 310 -1263 0 net=2863
rlabel metal2 404 -1265 404 -1265 0 net=3321
rlabel metal2 404 -1267 404 -1267 0 net=159
rlabel metal2 548 -1267 548 -1267 0 net=3233
rlabel metal2 411 -1269 411 -1269 0 net=3420
rlabel metal2 411 -1271 411 -1271 0 net=3288
rlabel metal2 429 -1273 429 -1273 0 net=2927
rlabel metal2 639 -1273 639 -1273 0 net=3719
rlabel metal2 702 -1273 702 -1273 0 net=3799
rlabel metal2 457 -1275 457 -1275 0 net=2895
rlabel metal2 513 -1275 513 -1275 0 net=2583
rlabel metal2 646 -1275 646 -1275 0 net=3993
rlabel metal2 474 -1277 474 -1277 0 net=2675
rlabel metal2 695 -1277 695 -1277 0 net=3795
rlabel metal2 303 -1279 303 -1279 0 net=4107
rlabel metal2 481 -1281 481 -1281 0 net=470
rlabel metal2 527 -1283 527 -1283 0 net=3649
rlabel metal2 569 -1285 569 -1285 0 net=2881
rlabel metal2 625 -1285 625 -1285 0 net=3791
rlabel metal2 275 -1287 275 -1287 0 net=3341
rlabel metal2 233 -1289 233 -1289 0 net=1307
rlabel metal2 233 -1291 233 -1291 0 net=1559
rlabel metal2 261 -1293 261 -1293 0 net=1189
rlabel metal2 296 -1295 296 -1295 0 net=1363
rlabel metal2 408 -1297 408 -1297 0 net=2455
rlabel metal2 2 -1308 2 -1308 0 net=2214
rlabel metal2 355 -1308 355 -1308 0 net=4146
rlabel metal2 782 -1308 782 -1308 0 net=3889
rlabel metal2 9 -1310 9 -1310 0 net=1338
rlabel metal2 191 -1310 191 -1310 0 net=2306
rlabel metal2 359 -1310 359 -1310 0 net=1738
rlabel metal2 516 -1310 516 -1310 0 net=3792
rlabel metal2 709 -1310 709 -1310 0 net=4108
rlabel metal2 9 -1312 9 -1312 0 net=20
rlabel metal2 362 -1312 362 -1312 0 net=2864
rlabel metal2 565 -1312 565 -1312 0 net=341
rlabel metal2 730 -1312 730 -1312 0 net=3041
rlabel metal2 30 -1314 30 -1314 0 net=2700
rlabel metal2 40 -1314 40 -1314 0 net=1450
rlabel metal2 65 -1314 65 -1314 0 net=3650
rlabel metal2 537 -1314 537 -1314 0 net=4122
rlabel metal2 30 -1316 30 -1316 0 net=1765
rlabel metal2 149 -1316 149 -1316 0 net=728
rlabel metal2 198 -1316 198 -1316 0 net=495
rlabel metal2 404 -1316 404 -1316 0 net=3058
rlabel metal2 527 -1316 527 -1316 0 net=3461
rlabel metal2 562 -1316 562 -1316 0 net=3796
rlabel metal2 44 -1318 44 -1318 0 net=2519
rlabel metal2 492 -1318 492 -1318 0 net=2677
rlabel metal2 590 -1318 590 -1318 0 net=4141
rlabel metal2 51 -1320 51 -1320 0 net=942
rlabel metal2 198 -1320 198 -1320 0 net=769
rlabel metal2 215 -1320 215 -1320 0 net=2171
rlabel metal2 408 -1320 408 -1320 0 net=3800
rlabel metal2 51 -1322 51 -1322 0 net=1033
rlabel metal2 149 -1322 149 -1322 0 net=741
rlabel metal2 163 -1322 163 -1322 0 net=2224
rlabel metal2 296 -1322 296 -1322 0 net=1364
rlabel metal2 457 -1322 457 -1322 0 net=2910
rlabel metal2 534 -1322 534 -1322 0 net=3587
rlabel metal2 632 -1322 632 -1322 0 net=3681
rlabel metal2 632 -1322 632 -1322 0 net=3681
rlabel metal2 639 -1322 639 -1322 0 net=3720
rlabel metal2 702 -1322 702 -1322 0 net=4012
rlabel metal2 68 -1324 68 -1324 0 net=1038
rlabel metal2 100 -1324 100 -1324 0 net=1579
rlabel metal2 100 -1324 100 -1324 0 net=1579
rlabel metal2 114 -1324 114 -1324 0 net=560
rlabel metal2 219 -1324 219 -1324 0 net=932
rlabel metal2 268 -1324 268 -1324 0 net=1717
rlabel metal2 310 -1324 310 -1324 0 net=2607
rlabel metal2 429 -1324 429 -1324 0 net=2929
rlabel metal2 541 -1324 541 -1324 0 net=2997
rlabel metal2 572 -1324 572 -1324 0 net=4170
rlabel metal2 58 -1326 58 -1326 0 net=1331
rlabel metal2 226 -1326 226 -1326 0 net=1153
rlabel metal2 275 -1326 275 -1326 0 net=1308
rlabel metal2 457 -1326 457 -1326 0 net=2567
rlabel metal2 485 -1326 485 -1326 0 net=2897
rlabel metal2 541 -1326 541 -1326 0 net=3235
rlabel metal2 576 -1326 576 -1326 0 net=3053
rlabel metal2 639 -1326 639 -1326 0 net=3701
rlabel metal2 688 -1326 688 -1326 0 net=4101
rlabel metal2 744 -1326 744 -1326 0 net=4135
rlabel metal2 23 -1328 23 -1328 0 net=1082
rlabel metal2 296 -1328 296 -1328 0 net=3189
rlabel metal2 653 -1328 653 -1328 0 net=3899
rlabel metal2 23 -1330 23 -1330 0 net=2457
rlabel metal2 425 -1330 425 -1330 0 net=4185
rlabel metal2 65 -1332 65 -1332 0 net=1183
rlabel metal2 114 -1332 114 -1332 0 net=3402
rlabel metal2 345 -1332 345 -1332 0 net=2317
rlabel metal2 471 -1332 471 -1332 0 net=2483
rlabel metal2 506 -1332 506 -1332 0 net=3087
rlabel metal2 72 -1334 72 -1334 0 net=3989
rlabel metal2 75 -1336 75 -1336 0 net=2311
rlabel metal2 506 -1336 506 -1336 0 net=2585
rlabel metal2 82 -1338 82 -1338 0 net=1678
rlabel metal2 117 -1338 117 -1338 0 net=2933
rlabel metal2 107 -1340 107 -1340 0 net=1433
rlabel metal2 191 -1340 191 -1340 0 net=1125
rlabel metal2 117 -1342 117 -1342 0 net=657
rlabel metal2 156 -1342 156 -1342 0 net=1397
rlabel metal2 177 -1342 177 -1342 0 net=1357
rlabel metal2 268 -1342 268 -1342 0 net=1639
rlabel metal2 16 -1344 16 -1344 0 net=2003
rlabel metal2 184 -1344 184 -1344 0 net=1953
rlabel metal2 352 -1344 352 -1344 0 net=1947
rlabel metal2 380 -1344 380 -1344 0 net=2283
rlabel metal2 464 -1344 464 -1344 0 net=2385
rlabel metal2 37 -1346 37 -1346 0 net=1470
rlabel metal2 163 -1346 163 -1346 0 net=2528
rlabel metal2 58 -1348 58 -1348 0 net=2195
rlabel metal2 233 -1348 233 -1348 0 net=1561
rlabel metal2 366 -1348 366 -1348 0 net=2375
rlabel metal2 86 -1350 86 -1350 0 net=1499
rlabel metal2 373 -1350 373 -1350 0 net=1901
rlabel metal2 121 -1352 121 -1352 0 net=1285
rlabel metal2 135 -1352 135 -1352 0 net=861
rlabel metal2 380 -1352 380 -1352 0 net=3195
rlabel metal2 121 -1354 121 -1354 0 net=1165
rlabel metal2 387 -1354 387 -1354 0 net=2579
rlabel metal2 597 -1354 597 -1354 0 net=3323
rlabel metal2 135 -1356 135 -1356 0 net=2139
rlabel metal2 387 -1356 387 -1356 0 net=2169
rlabel metal2 422 -1356 422 -1356 0 net=2399
rlabel metal2 443 -1356 443 -1356 0 net=2425
rlabel metal2 611 -1356 611 -1356 0 net=3343
rlabel metal2 166 -1358 166 -1358 0 net=453
rlabel metal2 254 -1360 254 -1360 0 net=1407
rlabel metal2 401 -1360 401 -1360 0 net=4013
rlabel metal2 212 -1362 212 -1362 0 net=1828
rlabel metal2 443 -1362 443 -1362 0 net=2882
rlabel metal2 261 -1364 261 -1364 0 net=1190
rlabel metal2 618 -1364 618 -1364 0 net=2703
rlabel metal2 79 -1366 79 -1366 0 net=1375
rlabel metal2 303 -1366 303 -1366 0 net=2299
rlabel metal2 660 -1366 660 -1366 0 net=3933
rlabel metal2 79 -1368 79 -1368 0 net=3688
rlabel metal2 681 -1368 681 -1368 0 net=3995
rlabel metal2 303 -1370 303 -1370 0 net=2147
rlabel metal2 331 -1370 331 -1370 0 net=3463
rlabel metal2 240 -1372 240 -1372 0 net=1489
rlabel metal2 240 -1374 240 -1374 0 net=2227
rlabel metal2 9 -1385 9 -1385 0 net=4207
rlabel metal2 149 -1385 149 -1385 0 net=742
rlabel metal2 170 -1385 170 -1385 0 net=2005
rlabel metal2 271 -1385 271 -1385 0 net=1490
rlabel metal2 338 -1385 338 -1385 0 net=1955
rlabel metal2 383 -1385 383 -1385 0 net=3749
rlabel metal2 758 -1385 758 -1385 0 net=4136
rlabel metal2 786 -1385 786 -1385 0 net=4137
rlabel metal2 16 -1387 16 -1387 0 net=3319
rlabel metal2 275 -1387 275 -1387 0 net=3196
rlabel metal2 411 -1387 411 -1387 0 net=3741
rlabel metal2 779 -1387 779 -1387 0 net=3043
rlabel metal2 37 -1389 37 -1389 0 net=2141
rlabel metal2 149 -1389 149 -1389 0 net=923
rlabel metal2 296 -1389 296 -1389 0 net=2312
rlabel metal2 443 -1389 443 -1389 0 net=3900
rlabel metal2 674 -1389 674 -1389 0 net=4015
rlabel metal2 789 -1389 789 -1389 0 net=3890
rlabel metal2 44 -1391 44 -1391 0 net=2520
rlabel metal2 247 -1391 247 -1391 0 net=1359
rlabel metal2 310 -1391 310 -1391 0 net=2608
rlabel metal2 338 -1391 338 -1391 0 net=1659
rlabel metal2 443 -1391 443 -1391 0 net=2071
rlabel metal2 534 -1391 534 -1391 0 net=2930
rlabel metal2 695 -1391 695 -1391 0 net=4103
rlabel metal2 796 -1391 796 -1391 0 net=692
rlabel metal2 44 -1393 44 -1393 0 net=1435
rlabel metal2 121 -1393 121 -1393 0 net=1167
rlabel metal2 156 -1393 156 -1393 0 net=1399
rlabel metal2 177 -1393 177 -1393 0 net=2300
rlabel metal2 457 -1393 457 -1393 0 net=2569
rlabel metal2 51 -1395 51 -1395 0 net=1034
rlabel metal2 163 -1395 163 -1395 0 net=1103
rlabel metal2 226 -1395 226 -1395 0 net=1155
rlabel metal2 324 -1395 324 -1395 0 net=1949
rlabel metal2 394 -1395 394 -1395 0 net=2285
rlabel metal2 450 -1395 450 -1395 0 net=2427
rlabel metal2 464 -1395 464 -1395 0 net=2387
rlabel metal2 464 -1395 464 -1395 0 net=2387
rlabel metal2 478 -1395 478 -1395 0 net=3054
rlabel metal2 590 -1395 590 -1395 0 net=3589
rlabel metal2 709 -1395 709 -1395 0 net=4143
rlabel metal2 51 -1397 51 -1397 0 net=2170
rlabel metal2 394 -1397 394 -1397 0 net=2318
rlabel metal2 488 -1397 488 -1397 0 net=3462
rlabel metal2 551 -1397 551 -1397 0 net=3934
rlabel metal2 674 -1397 674 -1397 0 net=3997
rlabel metal2 58 -1399 58 -1399 0 net=2197
rlabel metal2 75 -1399 75 -1399 0 net=269
rlabel metal2 226 -1399 226 -1399 0 net=1937
rlabel metal2 404 -1399 404 -1399 0 net=3705
rlabel metal2 58 -1401 58 -1401 0 net=1185
rlabel metal2 75 -1401 75 -1401 0 net=862
rlabel metal2 254 -1401 254 -1401 0 net=1409
rlabel metal2 303 -1401 303 -1401 0 net=2149
rlabel metal2 404 -1401 404 -1401 0 net=3579
rlabel metal2 79 -1403 79 -1403 0 net=1065
rlabel metal2 205 -1403 205 -1403 0 net=1627
rlabel metal2 348 -1403 348 -1403 0 net=3831
rlabel metal2 555 -1403 555 -1403 0 net=2998
rlabel metal2 79 -1405 79 -1405 0 net=1287
rlabel metal2 261 -1405 261 -1405 0 net=1377
rlabel metal2 317 -1405 317 -1405 0 net=3733
rlabel metal2 86 -1407 86 -1407 0 net=1581
rlabel metal2 117 -1407 117 -1407 0 net=2335
rlabel metal2 506 -1407 506 -1407 0 net=2587
rlabel metal2 639 -1407 639 -1407 0 net=3703
rlabel metal2 89 -1409 89 -1409 0 net=1313
rlabel metal2 261 -1409 261 -1409 0 net=1641
rlabel metal2 282 -1409 282 -1409 0 net=1563
rlabel metal2 352 -1409 352 -1409 0 net=2323
rlabel metal2 520 -1409 520 -1409 0 net=2899
rlabel metal2 618 -1409 618 -1409 0 net=2705
rlabel metal2 93 -1411 93 -1411 0 net=3344
rlabel metal2 646 -1411 646 -1411 0 net=3991
rlabel metal2 30 -1413 30 -1413 0 net=1767
rlabel metal2 100 -1413 100 -1413 0 net=2228
rlabel metal2 359 -1413 359 -1413 0 net=2173
rlabel metal2 506 -1413 506 -1413 0 net=3197
rlabel metal2 23 -1415 23 -1415 0 net=2459
rlabel metal2 107 -1415 107 -1415 0 net=907
rlabel metal2 128 -1415 128 -1415 0 net=771
rlabel metal2 219 -1415 219 -1415 0 net=1333
rlabel metal2 359 -1415 359 -1415 0 net=1903
rlabel metal2 411 -1415 411 -1415 0 net=2307
rlabel metal2 432 -1415 432 -1415 0 net=4179
rlabel metal2 562 -1415 562 -1415 0 net=3683
rlabel metal2 23 -1417 23 -1417 0 net=2581
rlabel metal2 492 -1417 492 -1417 0 net=2679
rlabel metal2 198 -1419 198 -1419 0 net=1719
rlabel metal2 366 -1419 366 -1419 0 net=2377
rlabel metal2 513 -1419 513 -1419 0 net=3163
rlabel metal2 219 -1421 219 -1421 0 net=1009
rlabel metal2 439 -1421 439 -1421 0 net=2405
rlabel metal2 520 -1421 520 -1421 0 net=2609
rlabel metal2 233 -1423 233 -1423 0 net=1501
rlabel metal2 334 -1423 334 -1423 0 net=1655
rlabel metal2 527 -1423 527 -1423 0 net=3089
rlabel metal2 565 -1423 565 -1423 0 net=3545
rlabel metal2 191 -1425 191 -1425 0 net=1127
rlabel metal2 240 -1425 240 -1425 0 net=1073
rlabel metal2 268 -1425 268 -1425 0 net=1739
rlabel metal2 541 -1425 541 -1425 0 net=3237
rlabel metal2 191 -1427 191 -1427 0 net=975
rlabel metal2 541 -1429 541 -1429 0 net=3289
rlabel metal2 548 -1431 548 -1431 0 net=3435
rlabel metal2 572 -1433 572 -1433 0 net=4186
rlabel metal2 576 -1435 576 -1435 0 net=3191
rlabel metal2 576 -1435 576 -1435 0 net=3191
rlabel metal2 583 -1435 583 -1435 0 net=3465
rlabel metal2 667 -1435 667 -1435 0 net=3547
rlabel metal2 485 -1437 485 -1437 0 net=2485
rlabel metal2 485 -1439 485 -1439 0 net=2915
rlabel metal2 597 -1439 597 -1439 0 net=3325
rlabel metal2 499 -1441 499 -1441 0 net=2935
rlabel metal2 436 -1443 436 -1443 0 net=2401
rlabel metal2 9 -1454 9 -1454 0 net=4208
rlabel metal2 128 -1454 128 -1454 0 net=773
rlabel metal2 681 -1454 681 -1454 0 net=3436
rlabel metal2 800 -1454 800 -1454 0 net=712
rlabel metal2 817 -1454 817 -1454 0 net=4138
rlabel metal2 9 -1456 9 -1456 0 net=1051
rlabel metal2 16 -1458 16 -1458 0 net=3320
rlabel metal2 439 -1458 439 -1458 0 net=2680
rlabel metal2 681 -1458 681 -1458 0 net=3743
rlabel metal2 768 -1458 768 -1458 0 net=3044
rlabel metal2 16 -1460 16 -1460 0 net=1941
rlabel metal2 474 -1460 474 -1460 0 net=4144
rlabel metal2 23 -1462 23 -1462 0 net=2582
rlabel metal2 156 -1462 156 -1462 0 net=3992
rlabel metal2 737 -1462 737 -1462 0 net=4105
rlabel metal2 23 -1464 23 -1464 0 net=1105
rlabel metal2 198 -1464 198 -1464 0 net=1720
rlabel metal2 394 -1464 394 -1464 0 net=2287
rlabel metal2 429 -1464 429 -1464 0 net=2486
rlabel metal2 632 -1464 632 -1464 0 net=3549
rlabel metal2 674 -1464 674 -1464 0 net=3999
rlabel metal2 30 -1466 30 -1466 0 net=2460
rlabel metal2 250 -1466 250 -1466 0 net=475
rlabel metal2 422 -1466 422 -1466 0 net=2379
rlabel metal2 509 -1466 509 -1466 0 net=3704
rlabel metal2 30 -1468 30 -1468 0 net=2503
rlabel metal2 257 -1468 257 -1468 0 net=3198
rlabel metal2 667 -1468 667 -1468 0 net=3735
rlabel metal2 37 -1470 37 -1470 0 net=2142
rlabel metal2 268 -1470 268 -1470 0 net=1360
rlabel metal2 303 -1470 303 -1470 0 net=1379
rlabel metal2 523 -1470 523 -1470 0 net=2588
rlabel metal2 688 -1470 688 -1470 0 net=3751
rlabel metal2 44 -1472 44 -1472 0 net=1436
rlabel metal2 128 -1472 128 -1472 0 net=1169
rlabel metal2 159 -1472 159 -1472 0 net=1723
rlabel metal2 432 -1472 432 -1472 0 net=3238
rlabel metal2 54 -1474 54 -1474 0 net=3909
rlabel metal2 58 -1476 58 -1476 0 net=1186
rlabel metal2 79 -1476 79 -1476 0 net=1289
rlabel metal2 114 -1476 114 -1476 0 net=1589
rlabel metal2 142 -1476 142 -1476 0 net=1067
rlabel metal2 296 -1476 296 -1476 0 net=1229
rlabel metal2 383 -1476 383 -1476 0 net=3117
rlabel metal2 37 -1478 37 -1478 0 net=1907
rlabel metal2 401 -1478 401 -1478 0 net=2428
rlabel metal2 527 -1478 527 -1478 0 net=3091
rlabel metal2 44 -1480 44 -1480 0 net=3171
rlabel metal2 212 -1480 212 -1480 0 net=2007
rlabel metal2 464 -1480 464 -1480 0 net=2389
rlabel metal2 534 -1480 534 -1480 0 net=3833
rlabel metal2 541 -1480 541 -1480 0 net=3291
rlabel metal2 58 -1482 58 -1482 0 net=1583
rlabel metal2 135 -1482 135 -1482 0 net=1201
rlabel metal2 212 -1482 212 -1482 0 net=1851
rlabel metal2 306 -1482 306 -1482 0 net=4016
rlabel metal2 65 -1484 65 -1484 0 net=2198
rlabel metal2 331 -1484 331 -1484 0 net=1956
rlabel metal2 352 -1484 352 -1484 0 net=2325
rlabel metal2 513 -1484 513 -1484 0 net=2407
rlabel metal2 555 -1484 555 -1484 0 net=4181
rlabel metal2 65 -1486 65 -1486 0 net=925
rlabel metal2 289 -1486 289 -1486 0 net=1503
rlabel metal2 359 -1486 359 -1486 0 net=1905
rlabel metal2 439 -1486 439 -1486 0 net=3326
rlabel metal2 79 -1488 79 -1488 0 net=1041
rlabel metal2 149 -1488 149 -1488 0 net=1011
rlabel metal2 289 -1488 289 -1488 0 net=1741
rlabel metal2 390 -1488 390 -1488 0 net=2027
rlabel metal2 478 -1488 478 -1488 0 net=2337
rlabel metal2 534 -1488 534 -1488 0 net=3165
rlabel metal2 646 -1488 646 -1488 0 net=2571
rlabel metal2 86 -1490 86 -1490 0 net=1411
rlabel metal2 317 -1490 317 -1490 0 net=1565
rlabel metal2 366 -1490 366 -1490 0 net=1657
rlabel metal2 555 -1490 555 -1490 0 net=3467
rlabel metal2 597 -1490 597 -1490 0 net=2937
rlabel metal2 170 -1492 170 -1492 0 net=1401
rlabel metal2 233 -1492 233 -1492 0 net=1129
rlabel metal2 282 -1492 282 -1492 0 net=1335
rlabel metal2 331 -1492 331 -1492 0 net=3192
rlabel metal2 597 -1492 597 -1492 0 net=4017
rlabel metal2 93 -1494 93 -1494 0 net=1768
rlabel metal2 191 -1494 191 -1494 0 net=977
rlabel metal2 387 -1494 387 -1494 0 net=2151
rlabel metal2 562 -1494 562 -1494 0 net=3685
rlabel metal2 121 -1496 121 -1496 0 net=729
rlabel metal2 233 -1496 233 -1496 0 net=227
rlabel metal2 310 -1496 310 -1496 0 net=1156
rlabel metal2 397 -1496 397 -1496 0 net=2659
rlabel metal2 618 -1496 618 -1496 0 net=2706
rlabel metal2 107 -1498 107 -1498 0 net=909
rlabel metal2 247 -1498 247 -1498 0 net=1315
rlabel metal2 334 -1498 334 -1498 0 net=3546
rlabel metal2 107 -1500 107 -1500 0 net=1593
rlabel metal2 198 -1500 198 -1500 0 net=951
rlabel metal2 261 -1500 261 -1500 0 net=1643
rlabel metal2 338 -1500 338 -1500 0 net=1661
rlabel metal2 450 -1500 450 -1500 0 net=2175
rlabel metal2 653 -1500 653 -1500 0 net=3581
rlabel metal2 240 -1502 240 -1502 0 net=1075
rlabel metal2 324 -1502 324 -1502 0 net=1950
rlabel metal2 341 -1502 341 -1502 0 net=2681
rlabel metal2 660 -1502 660 -1502 0 net=3591
rlabel metal2 240 -1504 240 -1504 0 net=394
rlabel metal2 450 -1504 450 -1504 0 net=2403
rlabel metal2 520 -1504 520 -1504 0 net=2611
rlabel metal2 324 -1506 324 -1506 0 net=2073
rlabel metal2 485 -1506 485 -1506 0 net=3393
rlabel metal2 537 -1506 537 -1506 0 net=1
rlabel metal2 226 -1508 226 -1508 0 net=1939
rlabel metal2 205 -1510 205 -1510 0 net=1629
rlabel metal2 362 -1510 362 -1510 0 net=3769
rlabel metal2 366 -1512 366 -1512 0 net=3706
rlabel metal2 380 -1514 380 -1514 0 net=3845
rlabel metal2 415 -1516 415 -1516 0 net=2309
rlabel metal2 415 -1518 415 -1518 0 net=2900
rlabel metal2 569 -1520 569 -1520 0 net=2917
rlabel metal2 359 -1522 359 -1522 0 net=2649
rlabel metal2 12 -1533 12 -1533 0 net=1942
rlabel metal2 51 -1533 51 -1533 0 net=230
rlabel metal2 208 -1533 208 -1533 0 net=1076
rlabel metal2 303 -1533 303 -1533 0 net=1336
rlabel metal2 331 -1533 331 -1533 0 net=265
rlabel metal2 488 -1533 488 -1533 0 net=4182
rlabel metal2 16 -1535 16 -1535 0 net=1853
rlabel metal2 226 -1535 226 -1535 0 net=1631
rlabel metal2 226 -1535 226 -1535 0 net=1631
rlabel metal2 240 -1535 240 -1535 0 net=2075
rlabel metal2 338 -1535 338 -1535 0 net=1380
rlabel metal2 520 -1535 520 -1535 0 net=3093
rlabel metal2 618 -1535 618 -1535 0 net=3737
rlabel metal2 2 -1537 2 -1537 0 net=1649
rlabel metal2 341 -1537 341 -1537 0 net=3951
rlabel metal2 23 -1539 23 -1539 0 net=1107
rlabel metal2 212 -1539 212 -1539 0 net=1743
rlabel metal2 303 -1539 303 -1539 0 net=2176
rlabel metal2 23 -1541 23 -1541 0 net=1505
rlabel metal2 362 -1541 362 -1541 0 net=1940
rlabel metal2 471 -1541 471 -1541 0 net=3770
rlabel metal2 44 -1543 44 -1543 0 net=3173
rlabel metal2 341 -1543 341 -1543 0 net=2310
rlabel metal2 597 -1543 597 -1543 0 net=4106
rlabel metal2 44 -1545 44 -1545 0 net=2650
rlabel metal2 604 -1545 604 -1545 0 net=3583
rlabel metal2 51 -1547 51 -1547 0 net=1171
rlabel metal2 138 -1547 138 -1547 0 net=2152
rlabel metal2 499 -1547 499 -1547 0 net=2939
rlabel metal2 58 -1549 58 -1549 0 net=1584
rlabel metal2 103 -1549 103 -1549 0 net=730
rlabel metal2 233 -1549 233 -1549 0 net=2811
rlabel metal2 569 -1549 569 -1549 0 net=3551
rlabel metal2 653 -1549 653 -1549 0 net=3847
rlabel metal2 58 -1551 58 -1551 0 net=2845
rlabel metal2 184 -1551 184 -1551 0 net=1130
rlabel metal2 278 -1551 278 -1551 0 net=2137
rlabel metal2 632 -1551 632 -1551 0 net=3753
rlabel metal2 72 -1553 72 -1553 0 net=1291
rlabel metal2 117 -1553 117 -1553 0 net=910
rlabel metal2 128 -1553 128 -1553 0 net=779
rlabel metal2 345 -1553 345 -1553 0 net=2409
rlabel metal2 79 -1555 79 -1555 0 net=1042
rlabel metal2 93 -1555 93 -1555 0 net=1591
rlabel metal2 121 -1555 121 -1555 0 net=1231
rlabel metal2 306 -1555 306 -1555 0 net=2008
rlabel metal2 82 -1557 82 -1557 0 net=1605
rlabel metal2 257 -1557 257 -1557 0 net=774
rlabel metal2 86 -1559 86 -1559 0 net=1413
rlabel metal2 289 -1559 289 -1559 0 net=1725
rlabel metal2 415 -1559 415 -1559 0 net=2572
rlabel metal2 65 -1561 65 -1561 0 net=926
rlabel metal2 415 -1561 415 -1561 0 net=2381
rlabel metal2 443 -1561 443 -1561 0 net=3166
rlabel metal2 548 -1561 548 -1561 0 net=3807
rlabel metal2 646 -1561 646 -1561 0 net=3835
rlabel metal2 30 -1563 30 -1563 0 net=2505
rlabel metal2 138 -1563 138 -1563 0 net=1402
rlabel metal2 247 -1563 247 -1563 0 net=1662
rlabel metal2 422 -1563 422 -1563 0 net=2327
rlabel metal2 534 -1563 534 -1563 0 net=3119
rlabel metal2 30 -1565 30 -1565 0 net=2682
rlabel metal2 611 -1565 611 -1565 0 net=3593
rlabel metal2 149 -1567 149 -1567 0 net=1013
rlabel metal2 170 -1567 170 -1567 0 net=1585
rlabel metal2 247 -1567 247 -1567 0 net=1645
rlabel metal2 296 -1567 296 -1567 0 net=2339
rlabel metal2 555 -1567 555 -1567 0 net=3469
rlabel metal2 660 -1567 660 -1567 0 net=3911
rlabel metal2 152 -1569 152 -1569 0 net=1566
rlabel metal2 362 -1569 362 -1569 0 net=3147
rlabel metal2 37 -1571 37 -1571 0 net=1909
rlabel metal2 366 -1571 366 -1571 0 net=1658
rlabel metal2 37 -1573 37 -1573 0 net=1595
rlabel metal2 184 -1573 184 -1573 0 net=953
rlabel metal2 219 -1573 219 -1573 0 net=3167
rlabel metal2 9 -1575 9 -1575 0 net=1053
rlabel metal2 177 -1575 177 -1575 0 net=2721
rlabel metal2 250 -1575 250 -1575 0 net=978
rlabel metal2 380 -1575 380 -1575 0 net=2404
rlabel metal2 457 -1575 457 -1575 0 net=2661
rlabel metal2 114 -1577 114 -1577 0 net=2199
rlabel metal2 387 -1577 387 -1577 0 net=3686
rlabel metal2 156 -1579 156 -1579 0 net=1203
rlabel metal2 187 -1579 187 -1579 0 net=526
rlabel metal2 261 -1579 261 -1579 0 net=1317
rlabel metal2 313 -1579 313 -1579 0 net=1906
rlabel metal2 439 -1579 439 -1579 0 net=2971
rlabel metal2 674 -1579 674 -1579 0 net=4001
rlabel metal2 142 -1581 142 -1581 0 net=1069
rlabel metal2 275 -1581 275 -1581 0 net=3559
rlabel metal2 394 -1581 394 -1581 0 net=2289
rlabel metal2 394 -1581 394 -1581 0 net=2289
rlabel metal2 401 -1581 401 -1581 0 net=2391
rlabel metal2 282 -1583 282 -1583 0 net=2683
rlabel metal2 334 -1583 334 -1583 0 net=3015
rlabel metal2 306 -1585 306 -1585 0 net=3103
rlabel metal2 418 -1587 418 -1587 0 net=2625
rlabel metal2 485 -1587 485 -1587 0 net=3395
rlabel metal2 387 -1589 387 -1589 0 net=2225
rlabel metal2 492 -1589 492 -1589 0 net=2919
rlabel metal2 411 -1591 411 -1591 0 net=3391
rlabel metal2 429 -1593 429 -1593 0 net=2029
rlabel metal2 464 -1595 464 -1595 0 net=2613
rlabel metal2 562 -1597 562 -1597 0 net=3293
rlabel metal2 625 -1599 625 -1599 0 net=3745
rlabel metal2 681 -1601 681 -1601 0 net=4019
rlabel metal2 5 -1612 5 -1612 0 net=1650
rlabel metal2 359 -1612 359 -1612 0 net=219
rlabel metal2 485 -1612 485 -1612 0 net=3095
rlabel metal2 558 -1612 558 -1612 0 net=3836
rlabel metal2 9 -1614 9 -1614 0 net=1071
rlabel metal2 163 -1614 163 -1614 0 net=1015
rlabel metal2 163 -1614 163 -1614 0 net=1015
rlabel metal2 187 -1614 187 -1614 0 net=2722
rlabel metal2 226 -1614 226 -1614 0 net=1632
rlabel metal2 317 -1614 317 -1614 0 net=2940
rlabel metal2 520 -1614 520 -1614 0 net=3397
rlabel metal2 625 -1614 625 -1614 0 net=3746
rlabel metal2 23 -1616 23 -1616 0 net=1507
rlabel metal2 82 -1616 82 -1616 0 net=3168
rlabel metal2 23 -1618 23 -1618 0 net=799
rlabel metal2 114 -1618 114 -1618 0 net=709
rlabel metal2 359 -1618 359 -1618 0 net=3120
rlabel metal2 30 -1620 30 -1620 0 net=2795
rlabel metal2 362 -1620 362 -1620 0 net=2290
rlabel metal2 401 -1620 401 -1620 0 net=2392
rlabel metal2 411 -1620 411 -1620 0 net=3754
rlabel metal2 30 -1622 30 -1622 0 net=661
rlabel metal2 233 -1622 233 -1622 0 net=1646
rlabel metal2 254 -1622 254 -1622 0 net=1607
rlabel metal2 366 -1622 366 -1622 0 net=2614
rlabel metal2 478 -1622 478 -1622 0 net=2813
rlabel metal2 534 -1622 534 -1622 0 net=3585
rlabel metal2 16 -1624 16 -1624 0 net=1855
rlabel metal2 16 -1626 16 -1626 0 net=905
rlabel metal2 152 -1626 152 -1626 0 net=2615
rlabel metal2 268 -1626 268 -1626 0 net=1415
rlabel metal2 373 -1626 373 -1626 0 net=3561
rlabel metal2 37 -1628 37 -1628 0 net=1596
rlabel metal2 128 -1628 128 -1628 0 net=781
rlabel metal2 170 -1628 170 -1628 0 net=1587
rlabel metal2 240 -1628 240 -1628 0 net=2077
rlabel metal2 376 -1628 376 -1628 0 net=2226
rlabel metal2 394 -1628 394 -1628 0 net=2973
rlabel metal2 37 -1630 37 -1630 0 net=1745
rlabel metal2 380 -1630 380 -1630 0 net=2201
rlabel metal2 506 -1630 506 -1630 0 net=3595
rlabel metal2 65 -1632 65 -1632 0 net=2506
rlabel metal2 292 -1632 292 -1632 0 net=4221
rlabel metal2 58 -1634 58 -1634 0 net=2847
rlabel metal2 72 -1634 72 -1634 0 net=1292
rlabel metal2 173 -1634 173 -1634 0 net=1701
rlabel metal2 205 -1634 205 -1634 0 net=1109
rlabel metal2 275 -1634 275 -1634 0 net=1911
rlabel metal2 380 -1634 380 -1634 0 net=2031
rlabel metal2 436 -1634 436 -1634 0 net=2663
rlabel metal2 58 -1636 58 -1636 0 net=877
rlabel metal2 205 -1636 205 -1636 0 net=1437
rlabel metal2 401 -1636 401 -1636 0 net=2329
rlabel metal2 429 -1636 429 -1636 0 net=2627
rlabel metal2 457 -1636 457 -1636 0 net=3179
rlabel metal2 47 -1638 47 -1638 0 net=109
rlabel metal2 212 -1638 212 -1638 0 net=1744
rlabel metal2 296 -1638 296 -1638 0 net=2340
rlabel metal2 408 -1638 408 -1638 0 net=3913
rlabel metal2 51 -1640 51 -1640 0 net=1173
rlabel metal2 439 -1640 439 -1640 0 net=3392
rlabel metal2 660 -1640 660 -1640 0 net=4003
rlabel metal2 51 -1642 51 -1642 0 net=674
rlabel metal2 443 -1642 443 -1642 0 net=2138
rlabel metal2 86 -1644 86 -1644 0 net=1881
rlabel metal2 184 -1644 184 -1644 0 net=955
rlabel metal2 296 -1644 296 -1644 0 net=4187
rlabel metal2 597 -1644 597 -1644 0 net=4021
rlabel metal2 72 -1646 72 -1646 0 net=1311
rlabel metal2 89 -1646 89 -1646 0 net=3848
rlabel metal2 677 -1646 677 -1646 0 net=4241
rlabel metal2 93 -1648 93 -1648 0 net=1592
rlabel metal2 128 -1648 128 -1648 0 net=1205
rlabel metal2 194 -1648 194 -1648 0 net=1917
rlabel metal2 93 -1650 93 -1650 0 net=1233
rlabel metal2 135 -1650 135 -1650 0 net=1931
rlabel metal2 212 -1650 212 -1650 0 net=1319
rlabel metal2 331 -1650 331 -1650 0 net=3174
rlabel metal2 443 -1650 443 -1650 0 net=3017
rlabel metal2 107 -1652 107 -1652 0 net=1055
rlabel metal2 446 -1652 446 -1652 0 net=3707
rlabel metal2 114 -1654 114 -1654 0 net=433
rlabel metal2 450 -1654 450 -1654 0 net=3149
rlabel metal2 121 -1656 121 -1656 0 net=1727
rlabel metal2 320 -1656 320 -1656 0 net=3767
rlabel metal2 282 -1658 282 -1658 0 net=2684
rlabel metal2 513 -1658 513 -1658 0 net=3295
rlabel metal2 282 -1660 282 -1660 0 net=2383
rlabel metal2 548 -1660 548 -1660 0 net=3809
rlabel metal2 345 -1662 345 -1662 0 net=2411
rlabel metal2 548 -1662 548 -1662 0 net=3553
rlabel metal2 345 -1664 345 -1664 0 net=2921
rlabel metal2 569 -1664 569 -1664 0 net=3739
rlabel metal2 492 -1666 492 -1666 0 net=3105
rlabel metal2 527 -1668 527 -1668 0 net=3471
rlabel metal2 583 -1670 583 -1670 0 net=3953
rlabel metal2 16 -1681 16 -1681 0 net=906
rlabel metal2 107 -1681 107 -1681 0 net=40
rlabel metal2 170 -1681 170 -1681 0 net=1933
rlabel metal2 187 -1681 187 -1681 0 net=1174
rlabel metal2 446 -1681 446 -1681 0 net=3106
rlabel metal2 506 -1681 506 -1681 0 net=3597
rlabel metal2 674 -1681 674 -1681 0 net=4243
rlabel metal2 16 -1683 16 -1683 0 net=1235
rlabel metal2 145 -1683 145 -1683 0 net=702
rlabel metal2 306 -1683 306 -1683 0 net=2202
rlabel metal2 534 -1683 534 -1683 0 net=3586
rlabel metal2 649 -1683 649 -1683 0 net=4004
rlabel metal2 23 -1685 23 -1685 0 net=800
rlabel metal2 156 -1685 156 -1685 0 net=783
rlabel metal2 212 -1685 212 -1685 0 net=1320
rlabel metal2 264 -1685 264 -1685 0 net=1856
rlabel metal2 471 -1685 471 -1685 0 net=3297
rlabel metal2 548 -1685 548 -1685 0 net=3554
rlabel metal2 23 -1687 23 -1687 0 net=2923
rlabel metal2 352 -1687 352 -1687 0 net=1918
rlabel metal2 30 -1689 30 -1689 0 net=1588
rlabel metal2 243 -1689 243 -1689 0 net=2796
rlabel metal2 331 -1689 331 -1689 0 net=3768
rlabel metal2 569 -1689 569 -1689 0 net=3740
rlabel metal2 37 -1691 37 -1691 0 net=1746
rlabel metal2 317 -1691 317 -1691 0 net=1608
rlabel metal2 376 -1691 376 -1691 0 net=2814
rlabel metal2 597 -1691 597 -1691 0 net=4023
rlabel metal2 9 -1693 9 -1693 0 net=1072
rlabel metal2 320 -1693 320 -1693 0 net=3914
rlabel metal2 499 -1693 499 -1693 0 net=3473
rlabel metal2 9 -1695 9 -1695 0 net=1207
rlabel metal2 173 -1695 173 -1695 0 net=491
rlabel metal2 338 -1695 338 -1695 0 net=4188
rlabel metal2 40 -1697 40 -1697 0 net=1702
rlabel metal2 212 -1697 212 -1697 0 net=1913
rlabel metal2 282 -1697 282 -1697 0 net=2384
rlabel metal2 390 -1697 390 -1697 0 net=3018
rlabel metal2 527 -1697 527 -1697 0 net=4223
rlabel metal2 44 -1699 44 -1699 0 net=1757
rlabel metal2 187 -1699 187 -1699 0 net=250
rlabel metal2 247 -1699 247 -1699 0 net=1110
rlabel metal2 292 -1699 292 -1699 0 net=2941
rlabel metal2 310 -1699 310 -1699 0 net=1416
rlabel metal2 408 -1699 408 -1699 0 net=2665
rlabel metal2 47 -1701 47 -1701 0 net=878
rlabel metal2 65 -1701 65 -1701 0 net=2849
rlabel metal2 271 -1701 271 -1701 0 net=3891
rlabel metal2 51 -1703 51 -1703 0 net=2161
rlabel metal2 275 -1703 275 -1703 0 net=2975
rlabel metal2 436 -1703 436 -1703 0 net=3151
rlabel metal2 58 -1705 58 -1705 0 net=3399
rlabel metal2 65 -1707 65 -1707 0 net=2467
rlabel metal2 198 -1707 198 -1707 0 net=1031
rlabel metal2 247 -1707 247 -1707 0 net=164
rlabel metal2 380 -1707 380 -1707 0 net=2033
rlabel metal2 520 -1707 520 -1707 0 net=3811
rlabel metal2 72 -1709 72 -1709 0 net=1312
rlabel metal2 219 -1709 219 -1709 0 net=957
rlabel metal2 250 -1709 250 -1709 0 net=4089
rlabel metal2 72 -1711 72 -1711 0 net=1439
rlabel metal2 254 -1711 254 -1711 0 net=2617
rlabel metal2 331 -1711 331 -1711 0 net=2413
rlabel metal2 79 -1713 79 -1713 0 net=1508
rlabel metal2 310 -1713 310 -1713 0 net=3562
rlabel metal2 79 -1715 79 -1715 0 net=2079
rlabel metal2 282 -1715 282 -1715 0 net=2629
rlabel metal2 86 -1717 86 -1717 0 net=1475
rlabel metal2 121 -1717 121 -1717 0 net=1729
rlabel metal2 240 -1717 240 -1717 0 net=3665
rlabel metal2 107 -1719 107 -1719 0 net=1349
rlabel metal2 149 -1719 149 -1719 0 net=1883
rlabel metal2 268 -1719 268 -1719 0 net=2667
rlabel metal2 373 -1719 373 -1719 0 net=3019
rlabel metal2 429 -1719 429 -1719 0 net=3097
rlabel metal2 114 -1721 114 -1721 0 net=1057
rlabel metal2 345 -1721 345 -1721 0 net=2331
rlabel metal2 485 -1721 485 -1721 0 net=3709
rlabel metal2 121 -1723 121 -1723 0 net=2901
rlabel metal2 401 -1723 401 -1723 0 net=3181
rlabel metal2 555 -1723 555 -1723 0 net=3955
rlabel metal2 135 -1725 135 -1725 0 net=1017
rlabel metal2 303 -1725 303 -1725 0 net=2065
rlabel metal2 163 -1727 163 -1727 0 net=2953
rlabel metal2 362 -1727 362 -1727 0 net=2983
rlabel metal2 16 -1738 16 -1738 0 net=1236
rlabel metal2 156 -1738 156 -1738 0 net=2511
rlabel metal2 254 -1738 254 -1738 0 net=11
rlabel metal2 261 -1738 261 -1738 0 net=2850
rlabel metal2 418 -1738 418 -1738 0 net=3885
rlabel metal2 548 -1738 548 -1738 0 net=3957
rlabel metal2 618 -1738 618 -1738 0 net=4025
rlabel metal2 618 -1738 618 -1738 0 net=4025
rlabel metal2 632 -1738 632 -1738 0 net=3599
rlabel metal2 670 -1738 670 -1738 0 net=4244
rlabel metal2 23 -1740 23 -1740 0 net=2924
rlabel metal2 422 -1740 422 -1740 0 net=3020
rlabel metal2 460 -1740 460 -1740 0 net=3812
rlabel metal2 37 -1742 37 -1742 0 net=1351
rlabel metal2 114 -1742 114 -1742 0 net=1058
rlabel metal2 208 -1742 208 -1742 0 net=2942
rlabel metal2 331 -1742 331 -1742 0 net=2415
rlabel metal2 408 -1742 408 -1742 0 net=2666
rlabel metal2 471 -1742 471 -1742 0 net=3299
rlabel metal2 44 -1744 44 -1744 0 net=1758
rlabel metal2 334 -1744 334 -1744 0 net=4090
rlabel metal2 51 -1746 51 -1746 0 net=2162
rlabel metal2 296 -1746 296 -1746 0 net=2669
rlabel metal2 422 -1746 422 -1746 0 net=3667
rlabel metal2 51 -1748 51 -1748 0 net=1019
rlabel metal2 145 -1748 145 -1748 0 net=1884
rlabel metal2 226 -1748 226 -1748 0 net=958
rlabel metal2 282 -1748 282 -1748 0 net=2631
rlabel metal2 338 -1748 338 -1748 0 net=3183
rlabel metal2 429 -1748 429 -1748 0 net=3098
rlabel metal2 58 -1750 58 -1750 0 net=3400
rlabel metal2 429 -1750 429 -1750 0 net=3893
rlabel metal2 471 -1750 471 -1750 0 net=4225
rlabel metal2 65 -1752 65 -1752 0 net=2468
rlabel metal2 117 -1752 117 -1752 0 net=593
rlabel metal2 212 -1752 212 -1752 0 net=1914
rlabel metal2 289 -1752 289 -1752 0 net=2619
rlabel metal2 345 -1752 345 -1752 0 net=2333
rlabel metal2 394 -1752 394 -1752 0 net=2035
rlabel metal2 478 -1752 478 -1752 0 net=3711
rlabel metal2 499 -1752 499 -1752 0 net=3475
rlabel metal2 72 -1754 72 -1754 0 net=1441
rlabel metal2 152 -1754 152 -1754 0 net=784
rlabel metal2 219 -1754 219 -1754 0 net=2067
rlabel metal2 310 -1754 310 -1754 0 net=4183
rlabel metal2 436 -1754 436 -1754 0 net=3153
rlabel metal2 72 -1756 72 -1756 0 net=2081
rlabel metal2 86 -1756 86 -1756 0 net=1476
rlabel metal2 124 -1756 124 -1756 0 net=731
rlabel metal2 159 -1756 159 -1756 0 net=2229
rlabel metal2 268 -1756 268 -1756 0 net=2903
rlabel metal2 65 -1758 65 -1758 0 net=2461
rlabel metal2 163 -1758 163 -1758 0 net=2955
rlabel metal2 275 -1758 275 -1758 0 net=2977
rlabel metal2 86 -1760 86 -1760 0 net=1857
rlabel metal2 128 -1760 128 -1760 0 net=911
rlabel metal2 324 -1760 324 -1760 0 net=2985
rlabel metal2 93 -1762 93 -1762 0 net=1245
rlabel metal2 163 -1762 163 -1762 0 net=3837
rlabel metal2 173 -1764 173 -1764 0 net=1032
rlabel metal2 233 -1764 233 -1764 0 net=1730
rlabel metal2 9 -1766 9 -1766 0 net=1209
rlabel metal2 170 -1768 170 -1768 0 net=1935
rlabel metal2 51 -1779 51 -1779 0 net=1020
rlabel metal2 198 -1779 198 -1779 0 net=1210
rlabel metal2 254 -1779 254 -1779 0 net=2620
rlabel metal2 317 -1779 317 -1779 0 net=2632
rlabel metal2 387 -1779 387 -1779 0 net=3894
rlabel metal2 464 -1779 464 -1779 0 net=2036
rlabel metal2 499 -1779 499 -1779 0 net=3886
rlabel metal2 541 -1779 541 -1779 0 net=3958
rlabel metal2 614 -1779 614 -1779 0 net=3600
rlabel metal2 51 -1781 51 -1781 0 net=3453
rlabel metal2 72 -1781 72 -1781 0 net=2082
rlabel metal2 345 -1781 345 -1781 0 net=2978
rlabel metal2 467 -1781 467 -1781 0 net=3154
rlabel metal2 618 -1781 618 -1781 0 net=4026
rlabel metal2 86 -1783 86 -1783 0 net=1858
rlabel metal2 110 -1783 110 -1783 0 net=87
rlabel metal2 247 -1783 247 -1783 0 net=2986
rlabel metal2 352 -1783 352 -1783 0 net=2416
rlabel metal2 471 -1783 471 -1783 0 net=4227
rlabel metal2 471 -1783 471 -1783 0 net=4227
rlabel metal2 478 -1783 478 -1783 0 net=3712
rlabel metal2 513 -1783 513 -1783 0 net=3300
rlabel metal2 93 -1785 93 -1785 0 net=1246
rlabel metal2 117 -1785 117 -1785 0 net=912
rlabel metal2 135 -1785 135 -1785 0 net=1443
rlabel metal2 156 -1785 156 -1785 0 net=2956
rlabel metal2 264 -1785 264 -1785 0 net=4184
rlabel metal2 338 -1785 338 -1785 0 net=3185
rlabel metal2 366 -1785 366 -1785 0 net=2334
rlabel metal2 520 -1785 520 -1785 0 net=3477
rlabel metal2 65 -1787 65 -1787 0 net=2462
rlabel metal2 124 -1787 124 -1787 0 net=2512
rlabel metal2 296 -1787 296 -1787 0 net=2670
rlabel metal2 373 -1787 373 -1787 0 net=3668
rlabel metal2 89 -1789 89 -1789 0 net=202
rlabel metal2 138 -1789 138 -1789 0 net=913
rlabel metal2 163 -1789 163 -1789 0 net=2904
rlabel metal2 142 -1791 142 -1791 0 net=732
rlabel metal2 173 -1791 173 -1791 0 net=2230
rlabel metal2 205 -1791 205 -1791 0 net=2069
rlabel metal2 37 -1793 37 -1793 0 net=1352
rlabel metal2 177 -1793 177 -1793 0 net=1936
rlabel metal2 233 -1795 233 -1795 0 net=3839
rlabel metal2 131 -1797 131 -1797 0 net=27
rlabel metal2 51 -1808 51 -1808 0 net=3454
rlabel metal2 145 -1808 145 -1808 0 net=2070
rlabel metal2 233 -1808 233 -1808 0 net=3840
rlabel metal2 352 -1808 352 -1808 0 net=3186
rlabel metal2 471 -1808 471 -1808 0 net=4228
rlabel metal2 520 -1808 520 -1808 0 net=3478
rlabel metal2 149 -1810 149 -1810 0 net=1444
rlabel metal2 156 -1812 156 -1812 0 net=914
rlabel metal2 180 -1812 180 -1812 0 net=335
<< end >>
