magic
tech scmos
timestamp 1555071772 
<< pdiffusion >>
rect 1 -8 7 -2
rect 8 -8 14 -2
rect 15 -8 21 -2
rect 22 -8 28 -2
rect 29 -8 35 -2
rect 36 -8 42 -2
rect 43 -8 49 -2
rect 50 -8 56 -2
rect 57 -8 63 -2
rect 134 -8 137 -2
rect 141 -8 147 -2
rect 148 -8 154 -2
rect 155 -8 161 -2
rect 183 -8 189 -2
rect 190 -8 196 -2
rect 211 -8 214 -2
rect 218 -8 224 -2
rect 253 -8 259 -2
rect 1 -23 7 -17
rect 8 -23 14 -17
rect 15 -23 21 -17
rect 22 -23 28 -17
rect 29 -23 35 -17
rect 36 -23 42 -17
rect 43 -23 49 -17
rect 50 -23 56 -17
rect 141 -23 147 -17
rect 148 -23 151 -17
rect 155 -23 158 -17
rect 162 -23 168 -17
rect 169 -23 175 -17
rect 176 -23 182 -17
rect 183 -23 186 -17
rect 190 -23 196 -17
rect 197 -23 200 -17
rect 204 -23 210 -17
rect 211 -23 214 -17
rect 218 -23 224 -17
rect 239 -23 245 -17
rect 253 -23 256 -17
rect 260 -23 266 -17
rect 267 -23 273 -17
rect 309 -23 315 -17
rect 1 -42 7 -36
rect 8 -42 14 -36
rect 15 -42 21 -36
rect 22 -42 28 -36
rect 29 -42 35 -36
rect 36 -42 42 -36
rect 43 -42 49 -36
rect 50 -42 56 -36
rect 99 -42 105 -36
rect 141 -42 147 -36
rect 148 -42 151 -36
rect 162 -42 165 -36
rect 169 -42 175 -36
rect 176 -42 182 -36
rect 183 -42 189 -36
rect 190 -42 193 -36
rect 197 -42 203 -36
rect 204 -42 210 -36
rect 211 -42 214 -36
rect 218 -42 221 -36
rect 225 -42 231 -36
rect 232 -42 238 -36
rect 239 -42 242 -36
rect 246 -42 249 -36
rect 253 -42 256 -36
rect 260 -42 263 -36
rect 267 -42 273 -36
rect 309 -42 312 -36
rect 337 -42 343 -36
rect 344 -42 347 -36
rect 358 -42 364 -36
rect 1 -65 7 -59
rect 8 -65 14 -59
rect 15 -65 21 -59
rect 22 -65 28 -59
rect 29 -65 35 -59
rect 36 -65 42 -59
rect 50 -65 56 -59
rect 71 -65 74 -59
rect 92 -65 98 -59
rect 99 -65 102 -59
rect 134 -65 140 -59
rect 141 -65 144 -59
rect 148 -65 154 -59
rect 155 -65 161 -59
rect 162 -65 165 -59
rect 169 -65 172 -59
rect 176 -65 182 -59
rect 183 -65 189 -59
rect 190 -65 196 -59
rect 197 -65 203 -59
rect 204 -65 207 -59
rect 211 -65 214 -59
rect 218 -65 221 -59
rect 225 -65 231 -59
rect 232 -65 235 -59
rect 239 -65 245 -59
rect 246 -65 249 -59
rect 253 -65 256 -59
rect 260 -65 263 -59
rect 267 -65 270 -59
rect 274 -65 280 -59
rect 281 -65 287 -59
rect 288 -65 291 -59
rect 295 -65 298 -59
rect 309 -65 312 -59
rect 316 -65 322 -59
rect 337 -65 340 -59
rect 344 -65 350 -59
rect 351 -65 354 -59
rect 365 -65 368 -59
rect 1 -96 7 -90
rect 8 -96 14 -90
rect 15 -96 21 -90
rect 22 -96 28 -90
rect 29 -96 35 -90
rect 50 -96 56 -90
rect 57 -96 60 -90
rect 64 -96 67 -90
rect 71 -96 74 -90
rect 78 -96 81 -90
rect 85 -96 91 -90
rect 92 -96 95 -90
rect 99 -96 105 -90
rect 106 -96 109 -90
rect 113 -96 116 -90
rect 120 -96 123 -90
rect 127 -96 130 -90
rect 134 -96 140 -90
rect 141 -96 147 -90
rect 148 -96 151 -90
rect 155 -96 158 -90
rect 162 -96 165 -90
rect 169 -96 175 -90
rect 176 -96 182 -90
rect 183 -96 189 -90
rect 190 -96 196 -90
rect 197 -96 203 -90
rect 204 -96 210 -90
rect 211 -96 214 -90
rect 218 -96 221 -90
rect 225 -96 231 -90
rect 232 -96 238 -90
rect 239 -96 245 -90
rect 246 -96 252 -90
rect 253 -96 259 -90
rect 260 -96 263 -90
rect 267 -96 270 -90
rect 274 -96 277 -90
rect 281 -96 284 -90
rect 288 -96 291 -90
rect 295 -96 298 -90
rect 302 -96 305 -90
rect 309 -96 312 -90
rect 316 -96 319 -90
rect 323 -96 326 -90
rect 330 -96 333 -90
rect 337 -96 340 -90
rect 344 -96 347 -90
rect 351 -96 354 -90
rect 365 -96 368 -90
rect 372 -96 378 -90
rect 1 -139 7 -133
rect 8 -139 14 -133
rect 15 -139 21 -133
rect 22 -139 28 -133
rect 85 -139 88 -133
rect 92 -139 95 -133
rect 99 -139 102 -133
rect 106 -139 109 -133
rect 113 -139 119 -133
rect 120 -139 126 -133
rect 127 -139 130 -133
rect 134 -139 137 -133
rect 141 -139 147 -133
rect 148 -139 151 -133
rect 155 -139 161 -133
rect 162 -139 165 -133
rect 169 -139 175 -133
rect 176 -139 182 -133
rect 183 -139 186 -133
rect 190 -139 196 -133
rect 197 -139 200 -133
rect 204 -139 210 -133
rect 211 -139 214 -133
rect 218 -139 221 -133
rect 225 -139 231 -133
rect 232 -139 238 -133
rect 239 -139 242 -133
rect 246 -139 252 -133
rect 253 -139 256 -133
rect 260 -139 266 -133
rect 267 -139 273 -133
rect 274 -139 277 -133
rect 281 -139 287 -133
rect 288 -139 294 -133
rect 295 -139 298 -133
rect 302 -139 305 -133
rect 309 -139 315 -133
rect 316 -139 319 -133
rect 323 -139 326 -133
rect 330 -139 333 -133
rect 337 -139 343 -133
rect 344 -139 347 -133
rect 351 -139 357 -133
rect 365 -139 368 -133
rect 379 -139 382 -133
rect 393 -139 396 -133
rect 400 -139 403 -133
rect 1 -174 7 -168
rect 8 -174 14 -168
rect 15 -174 21 -168
rect 64 -174 67 -168
rect 71 -174 74 -168
rect 78 -174 84 -168
rect 85 -174 88 -168
rect 92 -174 95 -168
rect 99 -174 102 -168
rect 106 -174 109 -168
rect 113 -174 119 -168
rect 120 -174 123 -168
rect 127 -174 133 -168
rect 134 -174 140 -168
rect 141 -174 147 -168
rect 148 -174 154 -168
rect 155 -174 158 -168
rect 162 -174 168 -168
rect 169 -174 172 -168
rect 176 -174 182 -168
rect 183 -174 186 -168
rect 190 -174 193 -168
rect 197 -174 203 -168
rect 204 -174 210 -168
rect 211 -174 214 -168
rect 218 -174 224 -168
rect 225 -174 231 -168
rect 232 -174 235 -168
rect 239 -174 245 -168
rect 246 -174 252 -168
rect 253 -174 256 -168
rect 260 -174 263 -168
rect 267 -174 270 -168
rect 274 -174 277 -168
rect 281 -174 287 -168
rect 288 -174 291 -168
rect 295 -174 298 -168
rect 302 -174 305 -168
rect 309 -174 315 -168
rect 316 -174 322 -168
rect 323 -174 326 -168
rect 330 -174 333 -168
rect 337 -174 343 -168
rect 344 -174 347 -168
rect 351 -174 354 -168
rect 358 -174 361 -168
rect 365 -174 368 -168
rect 372 -174 378 -168
rect 379 -174 382 -168
rect 386 -174 392 -168
rect 393 -174 396 -168
rect 400 -174 403 -168
rect 407 -174 410 -168
rect 414 -174 417 -168
rect 421 -174 424 -168
rect 428 -174 434 -168
rect 435 -174 441 -168
rect 1 -213 7 -207
rect 8 -213 14 -207
rect 22 -213 25 -207
rect 29 -213 32 -207
rect 36 -213 39 -207
rect 43 -213 46 -207
rect 50 -213 53 -207
rect 57 -213 63 -207
rect 64 -213 70 -207
rect 71 -213 77 -207
rect 78 -213 81 -207
rect 85 -213 91 -207
rect 92 -213 98 -207
rect 99 -213 102 -207
rect 106 -213 109 -207
rect 113 -213 116 -207
rect 120 -213 123 -207
rect 127 -213 130 -207
rect 134 -213 140 -207
rect 141 -213 147 -207
rect 148 -213 154 -207
rect 155 -213 161 -207
rect 162 -213 165 -207
rect 169 -213 172 -207
rect 176 -213 179 -207
rect 183 -213 186 -207
rect 190 -213 196 -207
rect 197 -213 203 -207
rect 204 -213 210 -207
rect 211 -213 217 -207
rect 218 -213 221 -207
rect 225 -213 228 -207
rect 232 -213 238 -207
rect 239 -213 245 -207
rect 246 -213 249 -207
rect 253 -213 256 -207
rect 260 -213 263 -207
rect 267 -213 273 -207
rect 274 -213 277 -207
rect 281 -213 287 -207
rect 288 -213 291 -207
rect 295 -213 301 -207
rect 302 -213 305 -207
rect 309 -213 312 -207
rect 316 -213 319 -207
rect 323 -213 329 -207
rect 330 -213 333 -207
rect 337 -213 343 -207
rect 344 -213 347 -207
rect 351 -213 354 -207
rect 358 -213 361 -207
rect 365 -213 368 -207
rect 372 -213 378 -207
rect 379 -213 382 -207
rect 386 -213 389 -207
rect 393 -213 396 -207
rect 400 -213 403 -207
rect 407 -213 413 -207
rect 414 -213 417 -207
rect 421 -213 424 -207
rect 428 -213 431 -207
rect 435 -213 438 -207
rect 442 -213 445 -207
rect 449 -213 452 -207
rect 456 -213 459 -207
rect 463 -213 466 -207
rect 540 -213 546 -207
rect 1 -260 7 -254
rect 36 -260 39 -254
rect 43 -260 46 -254
rect 50 -260 53 -254
rect 57 -260 60 -254
rect 64 -260 67 -254
rect 71 -260 77 -254
rect 78 -260 81 -254
rect 85 -260 88 -254
rect 92 -260 95 -254
rect 99 -260 102 -254
rect 106 -260 112 -254
rect 113 -260 119 -254
rect 120 -260 126 -254
rect 127 -260 133 -254
rect 134 -260 137 -254
rect 141 -260 147 -254
rect 148 -260 154 -254
rect 155 -260 158 -254
rect 162 -260 168 -254
rect 169 -260 175 -254
rect 176 -260 182 -254
rect 183 -260 186 -254
rect 190 -260 193 -254
rect 197 -260 203 -254
rect 204 -260 210 -254
rect 211 -260 214 -254
rect 218 -260 221 -254
rect 225 -260 231 -254
rect 232 -260 238 -254
rect 239 -260 245 -254
rect 246 -260 249 -254
rect 253 -260 256 -254
rect 260 -260 263 -254
rect 267 -260 270 -254
rect 274 -260 277 -254
rect 281 -260 287 -254
rect 288 -260 291 -254
rect 295 -260 298 -254
rect 302 -260 308 -254
rect 309 -260 312 -254
rect 316 -260 319 -254
rect 323 -260 329 -254
rect 330 -260 336 -254
rect 337 -260 343 -254
rect 344 -260 350 -254
rect 351 -260 357 -254
rect 358 -260 361 -254
rect 365 -260 368 -254
rect 372 -260 375 -254
rect 379 -260 382 -254
rect 386 -260 389 -254
rect 393 -260 396 -254
rect 400 -260 403 -254
rect 407 -260 410 -254
rect 414 -260 417 -254
rect 421 -260 424 -254
rect 428 -260 431 -254
rect 435 -260 438 -254
rect 442 -260 445 -254
rect 449 -260 452 -254
rect 456 -260 459 -254
rect 463 -260 466 -254
rect 470 -260 473 -254
rect 477 -260 480 -254
rect 484 -260 487 -254
rect 491 -260 494 -254
rect 498 -260 501 -254
rect 505 -260 508 -254
rect 512 -260 515 -254
rect 519 -260 522 -254
rect 526 -260 532 -254
rect 533 -260 539 -254
rect 540 -260 543 -254
rect 1 -307 7 -301
rect 36 -307 39 -301
rect 43 -307 49 -301
rect 50 -307 53 -301
rect 57 -307 63 -301
rect 64 -307 67 -301
rect 71 -307 74 -301
rect 78 -307 84 -301
rect 85 -307 91 -301
rect 92 -307 98 -301
rect 99 -307 102 -301
rect 106 -307 109 -301
rect 113 -307 119 -301
rect 120 -307 123 -301
rect 127 -307 133 -301
rect 134 -307 137 -301
rect 141 -307 144 -301
rect 148 -307 151 -301
rect 155 -307 158 -301
rect 162 -307 165 -301
rect 169 -307 172 -301
rect 176 -307 179 -301
rect 183 -307 186 -301
rect 190 -307 196 -301
rect 197 -307 200 -301
rect 204 -307 207 -301
rect 211 -307 214 -301
rect 218 -307 221 -301
rect 225 -307 228 -301
rect 232 -307 235 -301
rect 239 -307 242 -301
rect 246 -307 252 -301
rect 253 -307 256 -301
rect 260 -307 263 -301
rect 267 -307 273 -301
rect 274 -307 277 -301
rect 281 -307 287 -301
rect 288 -307 291 -301
rect 295 -307 298 -301
rect 302 -307 308 -301
rect 309 -307 312 -301
rect 316 -307 322 -301
rect 323 -307 326 -301
rect 330 -307 336 -301
rect 337 -307 343 -301
rect 344 -307 350 -301
rect 351 -307 354 -301
rect 358 -307 364 -301
rect 365 -307 371 -301
rect 372 -307 375 -301
rect 379 -307 385 -301
rect 386 -307 389 -301
rect 393 -307 396 -301
rect 400 -307 403 -301
rect 407 -307 410 -301
rect 414 -307 417 -301
rect 421 -307 424 -301
rect 428 -307 431 -301
rect 435 -307 438 -301
rect 442 -307 445 -301
rect 449 -307 452 -301
rect 456 -307 459 -301
rect 463 -307 469 -301
rect 470 -307 473 -301
rect 477 -307 480 -301
rect 484 -307 487 -301
rect 491 -307 494 -301
rect 498 -307 501 -301
rect 505 -307 508 -301
rect 512 -307 515 -301
rect 519 -307 522 -301
rect 526 -307 529 -301
rect 533 -307 536 -301
rect 540 -307 546 -301
rect 547 -307 550 -301
rect 554 -307 560 -301
rect 561 -307 567 -301
rect 568 -307 574 -301
rect 575 -307 578 -301
rect 8 -368 11 -362
rect 15 -368 18 -362
rect 22 -368 25 -362
rect 29 -368 32 -362
rect 36 -368 42 -362
rect 43 -368 46 -362
rect 50 -368 53 -362
rect 57 -368 63 -362
rect 64 -368 67 -362
rect 71 -368 74 -362
rect 78 -368 81 -362
rect 85 -368 88 -362
rect 92 -368 95 -362
rect 99 -368 105 -362
rect 106 -368 112 -362
rect 113 -368 116 -362
rect 120 -368 126 -362
rect 127 -368 133 -362
rect 134 -368 140 -362
rect 141 -368 144 -362
rect 148 -368 154 -362
rect 155 -368 161 -362
rect 162 -368 165 -362
rect 169 -368 172 -362
rect 176 -368 182 -362
rect 183 -368 186 -362
rect 190 -368 196 -362
rect 197 -368 200 -362
rect 204 -368 210 -362
rect 211 -368 214 -362
rect 218 -368 221 -362
rect 225 -368 228 -362
rect 232 -368 235 -362
rect 239 -368 245 -362
rect 246 -368 249 -362
rect 253 -368 256 -362
rect 260 -368 263 -362
rect 267 -368 273 -362
rect 274 -368 277 -362
rect 281 -368 287 -362
rect 288 -368 294 -362
rect 295 -368 301 -362
rect 302 -368 305 -362
rect 309 -368 315 -362
rect 316 -368 319 -362
rect 323 -368 329 -362
rect 330 -368 336 -362
rect 337 -368 343 -362
rect 344 -368 350 -362
rect 351 -368 357 -362
rect 358 -368 361 -362
rect 365 -368 371 -362
rect 372 -368 375 -362
rect 379 -368 385 -362
rect 386 -368 389 -362
rect 393 -368 396 -362
rect 400 -368 403 -362
rect 407 -368 410 -362
rect 414 -368 417 -362
rect 421 -368 424 -362
rect 428 -368 431 -362
rect 435 -368 438 -362
rect 442 -368 445 -362
rect 449 -368 452 -362
rect 456 -368 459 -362
rect 463 -368 466 -362
rect 470 -368 473 -362
rect 477 -368 480 -362
rect 484 -368 487 -362
rect 491 -368 494 -362
rect 498 -368 501 -362
rect 505 -368 508 -362
rect 512 -368 515 -362
rect 519 -368 522 -362
rect 526 -368 529 -362
rect 533 -368 536 -362
rect 540 -368 543 -362
rect 547 -368 550 -362
rect 554 -368 560 -362
rect 561 -368 564 -362
rect 568 -368 571 -362
rect 575 -368 578 -362
rect 1 -423 4 -417
rect 8 -423 14 -417
rect 15 -423 21 -417
rect 22 -423 25 -417
rect 29 -423 35 -417
rect 36 -423 39 -417
rect 43 -423 46 -417
rect 50 -423 53 -417
rect 57 -423 60 -417
rect 64 -423 70 -417
rect 71 -423 74 -417
rect 78 -423 81 -417
rect 85 -423 91 -417
rect 92 -423 98 -417
rect 99 -423 105 -417
rect 106 -423 109 -417
rect 113 -423 116 -417
rect 120 -423 123 -417
rect 127 -423 133 -417
rect 134 -423 140 -417
rect 141 -423 144 -417
rect 148 -423 154 -417
rect 155 -423 161 -417
rect 162 -423 165 -417
rect 169 -423 172 -417
rect 176 -423 179 -417
rect 183 -423 186 -417
rect 190 -423 193 -417
rect 197 -423 203 -417
rect 204 -423 210 -417
rect 211 -423 214 -417
rect 218 -423 221 -417
rect 225 -423 228 -417
rect 232 -423 235 -417
rect 239 -423 245 -417
rect 246 -423 252 -417
rect 253 -423 259 -417
rect 260 -423 263 -417
rect 267 -423 273 -417
rect 274 -423 280 -417
rect 281 -423 284 -417
rect 288 -423 294 -417
rect 295 -423 298 -417
rect 302 -423 308 -417
rect 309 -423 312 -417
rect 316 -423 322 -417
rect 323 -423 329 -417
rect 330 -423 333 -417
rect 337 -423 340 -417
rect 344 -423 350 -417
rect 351 -423 354 -417
rect 358 -423 364 -417
rect 365 -423 368 -417
rect 372 -423 375 -417
rect 379 -423 385 -417
rect 386 -423 392 -417
rect 393 -423 396 -417
rect 400 -423 403 -417
rect 407 -423 413 -417
rect 414 -423 417 -417
rect 421 -423 424 -417
rect 428 -423 431 -417
rect 435 -423 438 -417
rect 442 -423 445 -417
rect 449 -423 452 -417
rect 456 -423 459 -417
rect 463 -423 466 -417
rect 470 -423 473 -417
rect 477 -423 480 -417
rect 484 -423 487 -417
rect 491 -423 494 -417
rect 498 -423 501 -417
rect 505 -423 508 -417
rect 512 -423 515 -417
rect 519 -423 525 -417
rect 526 -423 529 -417
rect 533 -423 536 -417
rect 540 -423 543 -417
rect 547 -423 550 -417
rect 554 -423 557 -417
rect 561 -423 564 -417
rect 568 -423 571 -417
rect 575 -423 578 -417
rect 582 -423 585 -417
rect 610 -423 613 -417
rect 1 -500 4 -494
rect 8 -500 11 -494
rect 15 -500 18 -494
rect 22 -500 25 -494
rect 29 -500 32 -494
rect 36 -500 42 -494
rect 43 -500 49 -494
rect 50 -500 53 -494
rect 57 -500 60 -494
rect 64 -500 70 -494
rect 71 -500 74 -494
rect 78 -500 81 -494
rect 85 -500 88 -494
rect 92 -500 95 -494
rect 99 -500 102 -494
rect 106 -500 109 -494
rect 113 -500 119 -494
rect 120 -500 126 -494
rect 127 -500 133 -494
rect 134 -500 140 -494
rect 141 -500 147 -494
rect 148 -500 151 -494
rect 155 -500 158 -494
rect 162 -500 165 -494
rect 169 -500 175 -494
rect 176 -500 179 -494
rect 183 -500 189 -494
rect 190 -500 196 -494
rect 197 -500 203 -494
rect 204 -500 210 -494
rect 211 -500 214 -494
rect 218 -500 221 -494
rect 225 -500 228 -494
rect 232 -500 238 -494
rect 239 -500 245 -494
rect 246 -500 249 -494
rect 253 -500 256 -494
rect 260 -500 266 -494
rect 267 -500 270 -494
rect 274 -500 277 -494
rect 281 -500 284 -494
rect 288 -500 291 -494
rect 295 -500 298 -494
rect 302 -500 308 -494
rect 309 -500 315 -494
rect 316 -500 319 -494
rect 323 -500 329 -494
rect 330 -500 336 -494
rect 337 -500 340 -494
rect 344 -500 347 -494
rect 351 -500 357 -494
rect 358 -500 364 -494
rect 365 -500 368 -494
rect 372 -500 375 -494
rect 379 -500 382 -494
rect 386 -500 389 -494
rect 393 -500 399 -494
rect 400 -500 403 -494
rect 407 -500 410 -494
rect 414 -500 417 -494
rect 421 -500 427 -494
rect 428 -500 431 -494
rect 435 -500 438 -494
rect 442 -500 445 -494
rect 449 -500 452 -494
rect 456 -500 459 -494
rect 463 -500 466 -494
rect 470 -500 473 -494
rect 477 -500 480 -494
rect 484 -500 487 -494
rect 491 -500 497 -494
rect 498 -500 501 -494
rect 505 -500 508 -494
rect 512 -500 515 -494
rect 519 -500 522 -494
rect 526 -500 529 -494
rect 533 -500 536 -494
rect 540 -500 543 -494
rect 547 -500 550 -494
rect 554 -500 557 -494
rect 561 -500 564 -494
rect 568 -500 571 -494
rect 575 -500 578 -494
rect 582 -500 585 -494
rect 589 -500 592 -494
rect 596 -500 599 -494
rect 603 -500 606 -494
rect 610 -500 613 -494
rect 617 -500 623 -494
rect 624 -500 627 -494
rect 631 -500 637 -494
rect 638 -500 641 -494
rect 645 -500 648 -494
rect 652 -500 658 -494
rect 659 -500 665 -494
rect 666 -500 669 -494
rect 673 -500 676 -494
rect 15 -565 18 -559
rect 22 -565 25 -559
rect 29 -565 32 -559
rect 36 -565 39 -559
rect 43 -565 49 -559
rect 50 -565 53 -559
rect 57 -565 63 -559
rect 64 -565 67 -559
rect 71 -565 77 -559
rect 78 -565 84 -559
rect 85 -565 88 -559
rect 92 -565 95 -559
rect 99 -565 102 -559
rect 106 -565 109 -559
rect 113 -565 116 -559
rect 120 -565 123 -559
rect 127 -565 133 -559
rect 134 -565 137 -559
rect 141 -565 147 -559
rect 148 -565 154 -559
rect 155 -565 161 -559
rect 162 -565 165 -559
rect 169 -565 175 -559
rect 176 -565 179 -559
rect 183 -565 186 -559
rect 190 -565 196 -559
rect 197 -565 200 -559
rect 204 -565 210 -559
rect 211 -565 214 -559
rect 218 -565 221 -559
rect 225 -565 228 -559
rect 232 -565 235 -559
rect 239 -565 242 -559
rect 246 -565 249 -559
rect 253 -565 256 -559
rect 260 -565 266 -559
rect 267 -565 273 -559
rect 274 -565 280 -559
rect 281 -565 284 -559
rect 288 -565 291 -559
rect 295 -565 298 -559
rect 302 -565 305 -559
rect 309 -565 312 -559
rect 316 -565 319 -559
rect 323 -565 326 -559
rect 330 -565 336 -559
rect 337 -565 340 -559
rect 344 -565 350 -559
rect 351 -565 357 -559
rect 358 -565 361 -559
rect 365 -565 371 -559
rect 372 -565 375 -559
rect 379 -565 385 -559
rect 386 -565 392 -559
rect 393 -565 399 -559
rect 400 -565 406 -559
rect 407 -565 413 -559
rect 414 -565 417 -559
rect 421 -565 424 -559
rect 428 -565 431 -559
rect 435 -565 438 -559
rect 442 -565 445 -559
rect 449 -565 452 -559
rect 456 -565 459 -559
rect 463 -565 466 -559
rect 470 -565 473 -559
rect 477 -565 480 -559
rect 484 -565 490 -559
rect 491 -565 494 -559
rect 498 -565 501 -559
rect 505 -565 508 -559
rect 512 -565 515 -559
rect 519 -565 522 -559
rect 526 -565 529 -559
rect 533 -565 536 -559
rect 540 -565 543 -559
rect 547 -565 550 -559
rect 554 -565 557 -559
rect 561 -565 564 -559
rect 568 -565 571 -559
rect 575 -565 578 -559
rect 582 -565 585 -559
rect 589 -565 592 -559
rect 596 -565 599 -559
rect 603 -565 606 -559
rect 610 -565 616 -559
rect 617 -565 623 -559
rect 624 -565 630 -559
rect 631 -565 634 -559
rect 638 -565 644 -559
rect 645 -565 648 -559
rect 652 -565 655 -559
rect 1 -620 4 -614
rect 8 -620 11 -614
rect 15 -620 18 -614
rect 22 -620 25 -614
rect 29 -620 32 -614
rect 36 -620 39 -614
rect 43 -620 46 -614
rect 50 -620 53 -614
rect 57 -620 63 -614
rect 64 -620 70 -614
rect 71 -620 74 -614
rect 78 -620 81 -614
rect 85 -620 88 -614
rect 92 -620 95 -614
rect 99 -620 105 -614
rect 106 -620 109 -614
rect 113 -620 116 -614
rect 120 -620 126 -614
rect 127 -620 133 -614
rect 134 -620 137 -614
rect 141 -620 144 -614
rect 148 -620 154 -614
rect 155 -620 158 -614
rect 162 -620 168 -614
rect 169 -620 172 -614
rect 176 -620 182 -614
rect 183 -620 189 -614
rect 190 -620 196 -614
rect 197 -620 203 -614
rect 204 -620 210 -614
rect 211 -620 214 -614
rect 218 -620 221 -614
rect 225 -620 231 -614
rect 232 -620 235 -614
rect 239 -620 242 -614
rect 246 -620 249 -614
rect 253 -620 259 -614
rect 260 -620 263 -614
rect 267 -620 270 -614
rect 274 -620 280 -614
rect 281 -620 284 -614
rect 288 -620 291 -614
rect 295 -620 298 -614
rect 302 -620 305 -614
rect 309 -620 315 -614
rect 316 -620 319 -614
rect 323 -620 329 -614
rect 330 -620 336 -614
rect 337 -620 340 -614
rect 344 -620 350 -614
rect 351 -620 357 -614
rect 358 -620 364 -614
rect 365 -620 368 -614
rect 372 -620 375 -614
rect 379 -620 382 -614
rect 386 -620 389 -614
rect 393 -620 396 -614
rect 400 -620 406 -614
rect 407 -620 410 -614
rect 414 -620 417 -614
rect 421 -620 424 -614
rect 428 -620 431 -614
rect 435 -620 438 -614
rect 442 -620 445 -614
rect 449 -620 452 -614
rect 456 -620 462 -614
rect 463 -620 466 -614
rect 470 -620 473 -614
rect 477 -620 483 -614
rect 484 -620 487 -614
rect 491 -620 494 -614
rect 498 -620 501 -614
rect 505 -620 508 -614
rect 512 -620 515 -614
rect 519 -620 522 -614
rect 526 -620 532 -614
rect 533 -620 536 -614
rect 540 -620 546 -614
rect 547 -620 550 -614
rect 554 -620 557 -614
rect 561 -620 567 -614
rect 568 -620 571 -614
rect 575 -620 578 -614
rect 582 -620 585 -614
rect 589 -620 592 -614
rect 596 -620 599 -614
rect 603 -620 606 -614
rect 610 -620 613 -614
rect 617 -620 620 -614
rect 624 -620 630 -614
rect 631 -620 634 -614
rect 652 -620 655 -614
rect 1 -685 4 -679
rect 8 -685 11 -679
rect 15 -685 18 -679
rect 22 -685 28 -679
rect 29 -685 32 -679
rect 36 -685 39 -679
rect 43 -685 46 -679
rect 50 -685 56 -679
rect 57 -685 60 -679
rect 64 -685 67 -679
rect 71 -685 74 -679
rect 78 -685 81 -679
rect 85 -685 88 -679
rect 92 -685 98 -679
rect 99 -685 102 -679
rect 106 -685 109 -679
rect 113 -685 119 -679
rect 120 -685 126 -679
rect 127 -685 133 -679
rect 134 -685 140 -679
rect 141 -685 144 -679
rect 148 -685 154 -679
rect 155 -685 158 -679
rect 162 -685 165 -679
rect 169 -685 175 -679
rect 176 -685 182 -679
rect 183 -685 189 -679
rect 190 -685 193 -679
rect 197 -685 203 -679
rect 204 -685 210 -679
rect 211 -685 214 -679
rect 218 -685 224 -679
rect 225 -685 228 -679
rect 232 -685 235 -679
rect 239 -685 242 -679
rect 246 -685 249 -679
rect 253 -685 259 -679
rect 260 -685 263 -679
rect 267 -685 270 -679
rect 274 -685 280 -679
rect 281 -685 287 -679
rect 288 -685 294 -679
rect 295 -685 298 -679
rect 302 -685 305 -679
rect 309 -685 315 -679
rect 316 -685 319 -679
rect 323 -685 326 -679
rect 330 -685 336 -679
rect 337 -685 340 -679
rect 344 -685 347 -679
rect 351 -685 354 -679
rect 358 -685 361 -679
rect 365 -685 371 -679
rect 372 -685 378 -679
rect 379 -685 382 -679
rect 386 -685 389 -679
rect 393 -685 399 -679
rect 400 -685 406 -679
rect 407 -685 410 -679
rect 414 -685 417 -679
rect 421 -685 427 -679
rect 428 -685 434 -679
rect 435 -685 438 -679
rect 442 -685 445 -679
rect 449 -685 452 -679
rect 456 -685 459 -679
rect 463 -685 466 -679
rect 470 -685 473 -679
rect 477 -685 480 -679
rect 484 -685 487 -679
rect 491 -685 494 -679
rect 498 -685 501 -679
rect 505 -685 508 -679
rect 512 -685 515 -679
rect 519 -685 522 -679
rect 526 -685 529 -679
rect 533 -685 536 -679
rect 540 -685 543 -679
rect 547 -685 550 -679
rect 554 -685 560 -679
rect 561 -685 567 -679
rect 631 -685 634 -679
rect 638 -685 644 -679
rect 652 -685 655 -679
rect 1 -752 4 -746
rect 8 -752 14 -746
rect 15 -752 21 -746
rect 22 -752 28 -746
rect 29 -752 32 -746
rect 36 -752 39 -746
rect 43 -752 49 -746
rect 50 -752 53 -746
rect 57 -752 63 -746
rect 64 -752 67 -746
rect 71 -752 74 -746
rect 78 -752 84 -746
rect 85 -752 88 -746
rect 92 -752 95 -746
rect 99 -752 105 -746
rect 106 -752 109 -746
rect 113 -752 119 -746
rect 120 -752 123 -746
rect 127 -752 130 -746
rect 134 -752 137 -746
rect 141 -752 147 -746
rect 148 -752 154 -746
rect 155 -752 158 -746
rect 162 -752 168 -746
rect 169 -752 172 -746
rect 176 -752 179 -746
rect 183 -752 189 -746
rect 190 -752 196 -746
rect 197 -752 203 -746
rect 204 -752 210 -746
rect 211 -752 214 -746
rect 218 -752 221 -746
rect 225 -752 231 -746
rect 232 -752 235 -746
rect 239 -752 242 -746
rect 246 -752 249 -746
rect 253 -752 256 -746
rect 260 -752 266 -746
rect 267 -752 273 -746
rect 274 -752 280 -746
rect 281 -752 287 -746
rect 288 -752 291 -746
rect 295 -752 298 -746
rect 302 -752 308 -746
rect 309 -752 312 -746
rect 316 -752 319 -746
rect 323 -752 326 -746
rect 330 -752 333 -746
rect 337 -752 343 -746
rect 344 -752 347 -746
rect 351 -752 357 -746
rect 358 -752 364 -746
rect 365 -752 368 -746
rect 372 -752 378 -746
rect 379 -752 385 -746
rect 386 -752 389 -746
rect 393 -752 396 -746
rect 400 -752 403 -746
rect 407 -752 413 -746
rect 414 -752 417 -746
rect 421 -752 424 -746
rect 428 -752 431 -746
rect 435 -752 438 -746
rect 442 -752 445 -746
rect 449 -752 452 -746
rect 456 -752 459 -746
rect 463 -752 466 -746
rect 470 -752 476 -746
rect 477 -752 480 -746
rect 484 -752 487 -746
rect 491 -752 494 -746
rect 498 -752 501 -746
rect 505 -752 508 -746
rect 512 -752 515 -746
rect 519 -752 522 -746
rect 526 -752 529 -746
rect 533 -752 536 -746
rect 540 -752 543 -746
rect 547 -752 550 -746
rect 554 -752 557 -746
rect 561 -752 564 -746
rect 568 -752 571 -746
rect 575 -752 578 -746
rect 582 -752 585 -746
rect 589 -752 592 -746
rect 596 -752 599 -746
rect 603 -752 606 -746
rect 610 -752 613 -746
rect 617 -752 620 -746
rect 624 -752 627 -746
rect 631 -752 634 -746
rect 638 -752 641 -746
rect 645 -752 648 -746
rect 652 -752 658 -746
rect 659 -752 665 -746
rect 22 -825 25 -819
rect 29 -825 32 -819
rect 36 -825 42 -819
rect 43 -825 46 -819
rect 50 -825 56 -819
rect 57 -825 60 -819
rect 64 -825 67 -819
rect 71 -825 74 -819
rect 78 -825 84 -819
rect 85 -825 91 -819
rect 92 -825 98 -819
rect 99 -825 102 -819
rect 106 -825 109 -819
rect 113 -825 116 -819
rect 120 -825 123 -819
rect 127 -825 133 -819
rect 134 -825 140 -819
rect 141 -825 147 -819
rect 148 -825 154 -819
rect 155 -825 158 -819
rect 162 -825 165 -819
rect 169 -825 172 -819
rect 176 -825 179 -819
rect 183 -825 186 -819
rect 190 -825 193 -819
rect 197 -825 200 -819
rect 204 -825 207 -819
rect 211 -825 214 -819
rect 218 -825 221 -819
rect 225 -825 228 -819
rect 232 -825 235 -819
rect 239 -825 245 -819
rect 246 -825 249 -819
rect 253 -825 256 -819
rect 260 -825 263 -819
rect 267 -825 270 -819
rect 274 -825 280 -819
rect 281 -825 287 -819
rect 288 -825 291 -819
rect 295 -825 301 -819
rect 302 -825 305 -819
rect 309 -825 315 -819
rect 316 -825 322 -819
rect 323 -825 329 -819
rect 330 -825 336 -819
rect 337 -825 343 -819
rect 344 -825 347 -819
rect 351 -825 357 -819
rect 358 -825 361 -819
rect 365 -825 368 -819
rect 372 -825 378 -819
rect 379 -825 382 -819
rect 386 -825 392 -819
rect 393 -825 396 -819
rect 400 -825 406 -819
rect 407 -825 410 -819
rect 414 -825 417 -819
rect 421 -825 424 -819
rect 428 -825 431 -819
rect 435 -825 438 -819
rect 442 -825 445 -819
rect 449 -825 452 -819
rect 456 -825 459 -819
rect 463 -825 466 -819
rect 470 -825 473 -819
rect 477 -825 483 -819
rect 484 -825 487 -819
rect 491 -825 494 -819
rect 498 -825 501 -819
rect 505 -825 508 -819
rect 512 -825 518 -819
rect 519 -825 522 -819
rect 526 -825 529 -819
rect 533 -825 539 -819
rect 540 -825 543 -819
rect 547 -825 550 -819
rect 554 -825 560 -819
rect 561 -825 564 -819
rect 568 -825 574 -819
rect 575 -825 578 -819
rect 582 -825 585 -819
rect 589 -825 592 -819
rect 596 -825 602 -819
rect 603 -825 606 -819
rect 617 -825 620 -819
rect 1 -868 4 -862
rect 8 -868 11 -862
rect 15 -868 18 -862
rect 22 -868 25 -862
rect 29 -868 35 -862
rect 36 -868 42 -862
rect 43 -868 49 -862
rect 50 -868 53 -862
rect 57 -868 63 -862
rect 64 -868 67 -862
rect 71 -868 74 -862
rect 78 -868 84 -862
rect 85 -868 88 -862
rect 92 -868 95 -862
rect 99 -868 102 -862
rect 106 -868 109 -862
rect 113 -868 116 -862
rect 120 -868 123 -862
rect 127 -868 130 -862
rect 134 -868 140 -862
rect 141 -868 147 -862
rect 148 -868 151 -862
rect 155 -868 158 -862
rect 162 -868 168 -862
rect 169 -868 175 -862
rect 176 -868 182 -862
rect 183 -868 186 -862
rect 190 -868 196 -862
rect 197 -868 203 -862
rect 204 -868 210 -862
rect 211 -868 217 -862
rect 218 -868 224 -862
rect 225 -868 231 -862
rect 232 -868 235 -862
rect 239 -868 242 -862
rect 246 -868 249 -862
rect 253 -868 256 -862
rect 260 -868 266 -862
rect 267 -868 270 -862
rect 274 -868 277 -862
rect 281 -868 284 -862
rect 288 -868 294 -862
rect 295 -868 298 -862
rect 302 -868 305 -862
rect 309 -868 312 -862
rect 316 -868 322 -862
rect 323 -868 326 -862
rect 330 -868 333 -862
rect 337 -868 340 -862
rect 344 -868 350 -862
rect 351 -868 354 -862
rect 358 -868 361 -862
rect 365 -868 368 -862
rect 372 -868 378 -862
rect 379 -868 385 -862
rect 386 -868 389 -862
rect 393 -868 396 -862
rect 400 -868 403 -862
rect 407 -868 410 -862
rect 414 -868 417 -862
rect 421 -868 427 -862
rect 428 -868 431 -862
rect 435 -868 438 -862
rect 442 -868 445 -862
rect 449 -868 455 -862
rect 456 -868 459 -862
rect 463 -868 466 -862
rect 470 -868 473 -862
rect 477 -868 480 -862
rect 484 -868 487 -862
rect 491 -868 494 -862
rect 498 -868 501 -862
rect 505 -868 508 -862
rect 512 -868 518 -862
rect 519 -868 522 -862
rect 526 -868 532 -862
rect 533 -868 539 -862
rect 540 -868 546 -862
rect 547 -868 553 -862
rect 554 -868 557 -862
rect 561 -868 564 -862
rect 1 -923 4 -917
rect 8 -923 14 -917
rect 15 -923 18 -917
rect 22 -923 25 -917
rect 29 -923 35 -917
rect 36 -923 42 -917
rect 43 -923 49 -917
rect 50 -923 56 -917
rect 57 -923 63 -917
rect 64 -923 70 -917
rect 71 -923 77 -917
rect 78 -923 81 -917
rect 85 -923 88 -917
rect 92 -923 98 -917
rect 99 -923 105 -917
rect 106 -923 112 -917
rect 113 -923 116 -917
rect 120 -923 126 -917
rect 127 -923 133 -917
rect 134 -923 137 -917
rect 141 -923 144 -917
rect 148 -923 154 -917
rect 155 -923 158 -917
rect 162 -923 165 -917
rect 169 -923 175 -917
rect 176 -923 182 -917
rect 183 -923 189 -917
rect 190 -923 196 -917
rect 197 -923 203 -917
rect 204 -923 210 -917
rect 211 -923 214 -917
rect 218 -923 221 -917
rect 225 -923 231 -917
rect 232 -923 235 -917
rect 239 -923 245 -917
rect 246 -923 249 -917
rect 253 -923 256 -917
rect 260 -923 263 -917
rect 267 -923 270 -917
rect 274 -923 277 -917
rect 281 -923 284 -917
rect 288 -923 294 -917
rect 295 -923 301 -917
rect 302 -923 308 -917
rect 309 -923 315 -917
rect 316 -923 319 -917
rect 323 -923 326 -917
rect 330 -923 333 -917
rect 337 -923 340 -917
rect 344 -923 347 -917
rect 351 -923 354 -917
rect 358 -923 364 -917
rect 365 -923 368 -917
rect 372 -923 375 -917
rect 379 -923 382 -917
rect 386 -923 389 -917
rect 393 -923 396 -917
rect 400 -923 403 -917
rect 407 -923 410 -917
rect 414 -923 417 -917
rect 421 -923 424 -917
rect 428 -923 431 -917
rect 435 -923 438 -917
rect 442 -923 448 -917
rect 449 -923 452 -917
rect 456 -923 459 -917
rect 463 -923 466 -917
rect 470 -923 476 -917
rect 477 -923 480 -917
rect 484 -923 487 -917
rect 491 -923 494 -917
rect 498 -923 501 -917
rect 505 -923 508 -917
rect 512 -923 515 -917
rect 519 -923 522 -917
rect 526 -923 532 -917
rect 533 -923 536 -917
rect 540 -923 543 -917
rect 547 -923 550 -917
rect 22 -976 25 -970
rect 29 -976 32 -970
rect 36 -976 42 -970
rect 43 -976 49 -970
rect 50 -976 56 -970
rect 57 -976 60 -970
rect 64 -976 70 -970
rect 71 -976 74 -970
rect 78 -976 81 -970
rect 85 -976 88 -970
rect 92 -976 95 -970
rect 99 -976 102 -970
rect 106 -976 112 -970
rect 113 -976 119 -970
rect 120 -976 123 -970
rect 127 -976 133 -970
rect 134 -976 137 -970
rect 141 -976 147 -970
rect 148 -976 154 -970
rect 155 -976 158 -970
rect 162 -976 168 -970
rect 169 -976 172 -970
rect 176 -976 179 -970
rect 183 -976 189 -970
rect 190 -976 193 -970
rect 197 -976 203 -970
rect 204 -976 210 -970
rect 211 -976 214 -970
rect 218 -976 221 -970
rect 225 -976 231 -970
rect 232 -976 238 -970
rect 239 -976 242 -970
rect 246 -976 249 -970
rect 253 -976 256 -970
rect 260 -976 266 -970
rect 267 -976 270 -970
rect 274 -976 280 -970
rect 281 -976 287 -970
rect 288 -976 291 -970
rect 295 -976 301 -970
rect 302 -976 305 -970
rect 309 -976 312 -970
rect 316 -976 322 -970
rect 323 -976 326 -970
rect 330 -976 333 -970
rect 337 -976 340 -970
rect 344 -976 347 -970
rect 351 -976 357 -970
rect 358 -976 361 -970
rect 365 -976 368 -970
rect 372 -976 375 -970
rect 379 -976 385 -970
rect 386 -976 389 -970
rect 393 -976 396 -970
rect 400 -976 403 -970
rect 407 -976 413 -970
rect 414 -976 417 -970
rect 421 -976 427 -970
rect 428 -976 431 -970
rect 435 -976 438 -970
rect 442 -976 445 -970
rect 449 -976 452 -970
rect 456 -976 459 -970
rect 463 -976 469 -970
rect 470 -976 473 -970
rect 477 -976 483 -970
rect 484 -976 490 -970
rect 491 -976 494 -970
rect 498 -976 501 -970
rect 505 -976 511 -970
rect 519 -976 522 -970
rect 15 -1017 18 -1011
rect 22 -1017 28 -1011
rect 29 -1017 32 -1011
rect 36 -1017 39 -1011
rect 43 -1017 49 -1011
rect 50 -1017 53 -1011
rect 57 -1017 60 -1011
rect 64 -1017 70 -1011
rect 71 -1017 74 -1011
rect 78 -1017 81 -1011
rect 85 -1017 91 -1011
rect 92 -1017 98 -1011
rect 99 -1017 102 -1011
rect 106 -1017 109 -1011
rect 113 -1017 119 -1011
rect 120 -1017 123 -1011
rect 127 -1017 133 -1011
rect 134 -1017 137 -1011
rect 141 -1017 144 -1011
rect 148 -1017 151 -1011
rect 155 -1017 158 -1011
rect 162 -1017 165 -1011
rect 169 -1017 175 -1011
rect 176 -1017 179 -1011
rect 183 -1017 189 -1011
rect 190 -1017 196 -1011
rect 197 -1017 203 -1011
rect 204 -1017 210 -1011
rect 211 -1017 214 -1011
rect 218 -1017 221 -1011
rect 225 -1017 231 -1011
rect 232 -1017 238 -1011
rect 239 -1017 242 -1011
rect 246 -1017 249 -1011
rect 253 -1017 256 -1011
rect 260 -1017 263 -1011
rect 267 -1017 273 -1011
rect 274 -1017 280 -1011
rect 281 -1017 287 -1011
rect 288 -1017 294 -1011
rect 295 -1017 301 -1011
rect 302 -1017 305 -1011
rect 309 -1017 312 -1011
rect 316 -1017 319 -1011
rect 323 -1017 329 -1011
rect 330 -1017 333 -1011
rect 337 -1017 340 -1011
rect 344 -1017 347 -1011
rect 351 -1017 354 -1011
rect 358 -1017 361 -1011
rect 365 -1017 371 -1011
rect 372 -1017 375 -1011
rect 379 -1017 382 -1011
rect 386 -1017 392 -1011
rect 393 -1017 396 -1011
rect 400 -1017 403 -1011
rect 407 -1017 410 -1011
rect 414 -1017 417 -1011
rect 421 -1017 424 -1011
rect 428 -1017 434 -1011
rect 435 -1017 438 -1011
rect 442 -1017 448 -1011
rect 449 -1017 455 -1011
rect 456 -1017 459 -1011
rect 463 -1017 466 -1011
rect 470 -1017 473 -1011
rect 477 -1017 480 -1011
rect 519 -1017 525 -1011
rect 526 -1017 529 -1011
rect 64 -1054 67 -1048
rect 71 -1054 74 -1048
rect 78 -1054 84 -1048
rect 85 -1054 91 -1048
rect 92 -1054 95 -1048
rect 99 -1054 105 -1048
rect 106 -1054 109 -1048
rect 113 -1054 119 -1048
rect 120 -1054 123 -1048
rect 127 -1054 130 -1048
rect 134 -1054 137 -1048
rect 141 -1054 147 -1048
rect 148 -1054 154 -1048
rect 155 -1054 161 -1048
rect 162 -1054 168 -1048
rect 169 -1054 172 -1048
rect 176 -1054 179 -1048
rect 183 -1054 186 -1048
rect 190 -1054 193 -1048
rect 197 -1054 203 -1048
rect 204 -1054 210 -1048
rect 211 -1054 217 -1048
rect 218 -1054 221 -1048
rect 225 -1054 231 -1048
rect 232 -1054 238 -1048
rect 239 -1054 242 -1048
rect 246 -1054 252 -1048
rect 253 -1054 259 -1048
rect 260 -1054 263 -1048
rect 267 -1054 270 -1048
rect 274 -1054 277 -1048
rect 281 -1054 284 -1048
rect 288 -1054 294 -1048
rect 295 -1054 298 -1048
rect 302 -1054 305 -1048
rect 309 -1054 312 -1048
rect 316 -1054 319 -1048
rect 323 -1054 326 -1048
rect 330 -1054 336 -1048
rect 337 -1054 340 -1048
rect 344 -1054 347 -1048
rect 351 -1054 357 -1048
rect 358 -1054 361 -1048
rect 365 -1054 368 -1048
rect 372 -1054 375 -1048
rect 379 -1054 382 -1048
rect 386 -1054 389 -1048
rect 393 -1054 396 -1048
rect 400 -1054 403 -1048
rect 407 -1054 410 -1048
rect 414 -1054 417 -1048
rect 421 -1054 427 -1048
rect 428 -1054 434 -1048
rect 442 -1054 448 -1048
rect 449 -1054 455 -1048
rect 456 -1054 459 -1048
rect 477 -1054 480 -1048
rect 512 -1054 518 -1048
rect 519 -1054 525 -1048
rect 526 -1054 529 -1048
rect 50 -1099 53 -1093
rect 57 -1099 63 -1093
rect 64 -1099 67 -1093
rect 71 -1099 77 -1093
rect 78 -1099 84 -1093
rect 85 -1099 91 -1093
rect 92 -1099 95 -1093
rect 99 -1099 102 -1093
rect 106 -1099 112 -1093
rect 113 -1099 116 -1093
rect 120 -1099 123 -1093
rect 127 -1099 133 -1093
rect 134 -1099 140 -1093
rect 141 -1099 144 -1093
rect 148 -1099 151 -1093
rect 155 -1099 158 -1093
rect 162 -1099 165 -1093
rect 169 -1099 172 -1093
rect 176 -1099 182 -1093
rect 183 -1099 189 -1093
rect 190 -1099 196 -1093
rect 197 -1099 200 -1093
rect 204 -1099 207 -1093
rect 211 -1099 214 -1093
rect 218 -1099 224 -1093
rect 225 -1099 228 -1093
rect 232 -1099 238 -1093
rect 239 -1099 242 -1093
rect 246 -1099 249 -1093
rect 253 -1099 256 -1093
rect 260 -1099 263 -1093
rect 267 -1099 270 -1093
rect 274 -1099 277 -1093
rect 281 -1099 284 -1093
rect 288 -1099 294 -1093
rect 295 -1099 301 -1093
rect 302 -1099 308 -1093
rect 309 -1099 312 -1093
rect 316 -1099 322 -1093
rect 323 -1099 326 -1093
rect 330 -1099 333 -1093
rect 337 -1099 340 -1093
rect 344 -1099 347 -1093
rect 351 -1099 354 -1093
rect 358 -1099 361 -1093
rect 365 -1099 368 -1093
rect 372 -1099 378 -1093
rect 379 -1099 382 -1093
rect 386 -1099 392 -1093
rect 393 -1099 396 -1093
rect 400 -1099 403 -1093
rect 407 -1099 410 -1093
rect 414 -1099 420 -1093
rect 421 -1099 424 -1093
rect 428 -1099 431 -1093
rect 435 -1099 441 -1093
rect 456 -1099 462 -1093
rect 463 -1099 466 -1093
rect 477 -1099 480 -1093
rect 29 -1136 32 -1130
rect 36 -1136 39 -1130
rect 43 -1136 46 -1130
rect 50 -1136 56 -1130
rect 57 -1136 60 -1130
rect 64 -1136 67 -1130
rect 71 -1136 77 -1130
rect 78 -1136 84 -1130
rect 85 -1136 91 -1130
rect 92 -1136 98 -1130
rect 99 -1136 102 -1130
rect 106 -1136 109 -1130
rect 113 -1136 119 -1130
rect 120 -1136 123 -1130
rect 127 -1136 133 -1130
rect 134 -1136 137 -1130
rect 141 -1136 144 -1130
rect 148 -1136 151 -1130
rect 155 -1136 161 -1130
rect 162 -1136 165 -1130
rect 169 -1136 175 -1130
rect 176 -1136 179 -1130
rect 183 -1136 186 -1130
rect 190 -1136 196 -1130
rect 197 -1136 203 -1130
rect 204 -1136 210 -1130
rect 211 -1136 214 -1130
rect 218 -1136 221 -1130
rect 225 -1136 231 -1130
rect 232 -1136 235 -1130
rect 239 -1136 242 -1130
rect 246 -1136 249 -1130
rect 253 -1136 259 -1130
rect 260 -1136 266 -1130
rect 267 -1136 270 -1130
rect 274 -1136 280 -1130
rect 281 -1136 284 -1130
rect 288 -1136 291 -1130
rect 295 -1136 298 -1130
rect 302 -1136 308 -1130
rect 309 -1136 312 -1130
rect 316 -1136 322 -1130
rect 323 -1136 329 -1130
rect 330 -1136 333 -1130
rect 337 -1136 340 -1130
rect 344 -1136 347 -1130
rect 351 -1136 354 -1130
rect 358 -1136 364 -1130
rect 365 -1136 371 -1130
rect 372 -1136 375 -1130
rect 379 -1136 382 -1130
rect 386 -1136 389 -1130
rect 393 -1136 396 -1130
rect 400 -1136 403 -1130
rect 407 -1136 410 -1130
rect 414 -1136 417 -1130
rect 421 -1136 424 -1130
rect 428 -1136 431 -1130
rect 435 -1136 438 -1130
rect 442 -1136 445 -1130
rect 477 -1136 480 -1130
rect 484 -1136 490 -1130
rect 50 -1179 56 -1173
rect 57 -1179 63 -1173
rect 71 -1179 74 -1173
rect 78 -1179 84 -1173
rect 85 -1179 88 -1173
rect 92 -1179 98 -1173
rect 99 -1179 102 -1173
rect 106 -1179 109 -1173
rect 113 -1179 119 -1173
rect 120 -1179 126 -1173
rect 127 -1179 130 -1173
rect 134 -1179 137 -1173
rect 141 -1179 147 -1173
rect 148 -1179 151 -1173
rect 155 -1179 158 -1173
rect 162 -1179 168 -1173
rect 169 -1179 175 -1173
rect 176 -1179 179 -1173
rect 183 -1179 186 -1173
rect 190 -1179 193 -1173
rect 197 -1179 203 -1173
rect 204 -1179 210 -1173
rect 211 -1179 214 -1173
rect 218 -1179 221 -1173
rect 225 -1179 228 -1173
rect 232 -1179 235 -1173
rect 239 -1179 245 -1173
rect 246 -1179 252 -1173
rect 253 -1179 259 -1173
rect 260 -1179 266 -1173
rect 267 -1179 270 -1173
rect 274 -1179 277 -1173
rect 281 -1179 284 -1173
rect 288 -1179 291 -1173
rect 295 -1179 301 -1173
rect 302 -1179 308 -1173
rect 309 -1179 312 -1173
rect 316 -1179 319 -1173
rect 323 -1179 326 -1173
rect 330 -1179 333 -1173
rect 337 -1179 340 -1173
rect 344 -1179 347 -1173
rect 351 -1179 354 -1173
rect 358 -1179 361 -1173
rect 365 -1179 368 -1173
rect 372 -1179 378 -1173
rect 379 -1179 382 -1173
rect 386 -1179 389 -1173
rect 393 -1179 399 -1173
rect 400 -1179 403 -1173
rect 407 -1179 413 -1173
rect 64 -1210 67 -1204
rect 71 -1210 74 -1204
rect 78 -1210 81 -1204
rect 85 -1210 91 -1204
rect 92 -1210 95 -1204
rect 99 -1210 102 -1204
rect 106 -1210 112 -1204
rect 113 -1210 116 -1204
rect 120 -1210 123 -1204
rect 127 -1210 133 -1204
rect 134 -1210 140 -1204
rect 141 -1210 144 -1204
rect 148 -1210 154 -1204
rect 155 -1210 161 -1204
rect 162 -1210 165 -1204
rect 169 -1210 175 -1204
rect 176 -1210 182 -1204
rect 183 -1210 189 -1204
rect 190 -1210 196 -1204
rect 197 -1210 200 -1204
rect 204 -1210 210 -1204
rect 211 -1210 214 -1204
rect 218 -1210 221 -1204
rect 225 -1210 231 -1204
rect 232 -1210 235 -1204
rect 239 -1210 245 -1204
rect 246 -1210 249 -1204
rect 253 -1210 256 -1204
rect 260 -1210 266 -1204
rect 267 -1210 270 -1204
rect 274 -1210 277 -1204
rect 281 -1210 284 -1204
rect 288 -1210 294 -1204
rect 295 -1210 298 -1204
rect 302 -1210 308 -1204
rect 309 -1210 312 -1204
rect 316 -1210 322 -1204
rect 323 -1210 329 -1204
rect 330 -1210 333 -1204
rect 337 -1210 340 -1204
rect 344 -1210 347 -1204
rect 351 -1210 354 -1204
rect 358 -1210 361 -1204
rect 365 -1210 368 -1204
rect 372 -1210 375 -1204
rect 379 -1210 385 -1204
rect 386 -1210 389 -1204
rect 393 -1210 396 -1204
rect 92 -1239 95 -1233
rect 99 -1239 105 -1233
rect 106 -1239 112 -1233
rect 113 -1239 116 -1233
rect 120 -1239 126 -1233
rect 127 -1239 130 -1233
rect 134 -1239 137 -1233
rect 141 -1239 144 -1233
rect 148 -1239 154 -1233
rect 155 -1239 158 -1233
rect 162 -1239 165 -1233
rect 169 -1239 175 -1233
rect 176 -1239 182 -1233
rect 183 -1239 189 -1233
rect 190 -1239 196 -1233
rect 197 -1239 203 -1233
rect 204 -1239 207 -1233
rect 211 -1239 214 -1233
rect 218 -1239 224 -1233
rect 225 -1239 228 -1233
rect 232 -1239 235 -1233
rect 239 -1239 242 -1233
rect 246 -1239 249 -1233
rect 253 -1239 259 -1233
rect 260 -1239 266 -1233
rect 267 -1239 273 -1233
rect 274 -1239 277 -1233
rect 281 -1239 284 -1233
rect 288 -1239 291 -1233
rect 295 -1239 301 -1233
rect 302 -1239 308 -1233
rect 309 -1239 312 -1233
rect 316 -1239 319 -1233
rect 323 -1239 326 -1233
rect 330 -1239 333 -1233
rect 344 -1239 350 -1233
rect 351 -1239 354 -1233
rect 379 -1239 382 -1233
rect 1 -1260 7 -1254
rect 71 -1260 77 -1254
rect 78 -1260 84 -1254
rect 85 -1260 88 -1254
rect 99 -1260 102 -1254
rect 106 -1260 109 -1254
rect 113 -1260 119 -1254
rect 120 -1260 126 -1254
rect 127 -1260 133 -1254
rect 134 -1260 137 -1254
rect 141 -1260 147 -1254
rect 148 -1260 154 -1254
rect 155 -1260 161 -1254
rect 162 -1260 168 -1254
rect 169 -1260 175 -1254
rect 176 -1260 179 -1254
rect 183 -1260 189 -1254
rect 190 -1260 193 -1254
rect 197 -1260 203 -1254
rect 204 -1260 207 -1254
rect 211 -1260 217 -1254
rect 218 -1260 221 -1254
rect 225 -1260 231 -1254
rect 232 -1260 235 -1254
rect 239 -1260 242 -1254
rect 246 -1260 252 -1254
rect 253 -1260 256 -1254
rect 260 -1260 263 -1254
rect 267 -1260 270 -1254
rect 274 -1260 280 -1254
rect 281 -1260 287 -1254
rect 288 -1260 294 -1254
rect 295 -1260 298 -1254
rect 302 -1260 305 -1254
rect 316 -1260 322 -1254
rect 323 -1260 326 -1254
rect 379 -1260 382 -1254
rect 1 -1275 7 -1269
rect 85 -1275 91 -1269
rect 92 -1275 98 -1269
rect 106 -1275 109 -1269
rect 113 -1275 119 -1269
rect 120 -1275 123 -1269
rect 127 -1275 133 -1269
rect 134 -1275 137 -1269
rect 141 -1275 147 -1269
rect 148 -1275 151 -1269
rect 155 -1275 161 -1269
rect 162 -1275 168 -1269
rect 169 -1275 175 -1269
rect 183 -1275 189 -1269
rect 204 -1275 210 -1269
rect 211 -1275 217 -1269
rect 218 -1275 224 -1269
rect 225 -1275 228 -1269
rect 232 -1275 238 -1269
rect 239 -1275 245 -1269
rect 267 -1275 273 -1269
rect 274 -1275 277 -1269
rect 281 -1275 287 -1269
rect 295 -1275 301 -1269
rect 302 -1275 305 -1269
rect 379 -1275 385 -1269
rect 386 -1275 389 -1269
<< polysilicon >>
rect 135 -3 136 -1
rect 135 -9 136 -7
rect 142 -3 143 -1
rect 145 -3 146 -1
rect 142 -9 143 -7
rect 149 -9 150 -7
rect 152 -9 153 -7
rect 156 -3 157 -1
rect 184 -3 185 -1
rect 184 -9 185 -7
rect 194 -3 195 -1
rect 212 -3 213 -1
rect 212 -9 213 -7
rect 219 -3 220 -1
rect 254 -9 255 -7
rect 257 -9 258 -7
rect 142 -18 143 -16
rect 149 -18 150 -16
rect 149 -24 150 -22
rect 156 -18 157 -16
rect 156 -24 157 -22
rect 163 -24 164 -22
rect 166 -24 167 -22
rect 173 -24 174 -22
rect 177 -18 178 -16
rect 180 -18 181 -16
rect 177 -24 178 -22
rect 184 -18 185 -16
rect 184 -24 185 -22
rect 191 -18 192 -16
rect 198 -18 199 -16
rect 198 -24 199 -22
rect 205 -18 206 -16
rect 208 -18 209 -16
rect 205 -24 206 -22
rect 212 -18 213 -16
rect 212 -24 213 -22
rect 222 -18 223 -16
rect 243 -24 244 -22
rect 254 -18 255 -16
rect 254 -24 255 -22
rect 261 -18 262 -16
rect 268 -24 269 -22
rect 310 -24 311 -22
rect 54 -43 55 -41
rect 100 -43 101 -41
rect 145 -37 146 -35
rect 149 -37 150 -35
rect 149 -43 150 -41
rect 163 -37 164 -35
rect 163 -43 164 -41
rect 170 -37 171 -35
rect 177 -43 178 -41
rect 187 -37 188 -35
rect 187 -43 188 -41
rect 191 -37 192 -35
rect 191 -43 192 -41
rect 201 -37 202 -35
rect 198 -43 199 -41
rect 208 -37 209 -35
rect 208 -43 209 -41
rect 212 -37 213 -35
rect 212 -43 213 -41
rect 219 -37 220 -35
rect 219 -43 220 -41
rect 229 -37 230 -35
rect 233 -37 234 -35
rect 233 -43 234 -41
rect 236 -43 237 -41
rect 240 -37 241 -35
rect 240 -43 241 -41
rect 247 -37 248 -35
rect 247 -43 248 -41
rect 254 -37 255 -35
rect 254 -43 255 -41
rect 261 -37 262 -35
rect 261 -43 262 -41
rect 271 -37 272 -35
rect 268 -43 269 -41
rect 310 -37 311 -35
rect 310 -43 311 -41
rect 341 -37 342 -35
rect 338 -43 339 -41
rect 345 -37 346 -35
rect 345 -43 346 -41
rect 359 -43 360 -41
rect 362 -43 363 -41
rect 26 -66 27 -64
rect 51 -60 52 -58
rect 72 -60 73 -58
rect 72 -66 73 -64
rect 96 -60 97 -58
rect 93 -66 94 -64
rect 96 -66 97 -64
rect 100 -60 101 -58
rect 100 -66 101 -64
rect 138 -60 139 -58
rect 142 -60 143 -58
rect 142 -66 143 -64
rect 149 -66 150 -64
rect 156 -60 157 -58
rect 163 -60 164 -58
rect 163 -66 164 -64
rect 170 -60 171 -58
rect 170 -66 171 -64
rect 177 -60 178 -58
rect 187 -60 188 -58
rect 187 -66 188 -64
rect 191 -60 192 -58
rect 194 -60 195 -58
rect 198 -60 199 -58
rect 201 -60 202 -58
rect 201 -66 202 -64
rect 205 -60 206 -58
rect 205 -66 206 -64
rect 212 -60 213 -58
rect 212 -66 213 -64
rect 219 -60 220 -58
rect 219 -66 220 -64
rect 226 -60 227 -58
rect 226 -66 227 -64
rect 229 -66 230 -64
rect 233 -60 234 -58
rect 233 -66 234 -64
rect 240 -60 241 -58
rect 243 -60 244 -58
rect 240 -66 241 -64
rect 247 -60 248 -58
rect 247 -66 248 -64
rect 254 -60 255 -58
rect 254 -66 255 -64
rect 261 -60 262 -58
rect 261 -66 262 -64
rect 268 -60 269 -58
rect 268 -66 269 -64
rect 275 -60 276 -58
rect 278 -66 279 -64
rect 282 -60 283 -58
rect 282 -66 283 -64
rect 289 -60 290 -58
rect 289 -66 290 -64
rect 296 -60 297 -58
rect 296 -66 297 -64
rect 310 -60 311 -58
rect 310 -66 311 -64
rect 317 -66 318 -64
rect 320 -66 321 -64
rect 338 -60 339 -58
rect 338 -66 339 -64
rect 345 -60 346 -58
rect 348 -66 349 -64
rect 352 -60 353 -58
rect 352 -66 353 -64
rect 366 -60 367 -58
rect 366 -66 367 -64
rect 26 -91 27 -89
rect 51 -91 52 -89
rect 58 -91 59 -89
rect 58 -97 59 -95
rect 65 -91 66 -89
rect 65 -97 66 -95
rect 72 -91 73 -89
rect 72 -97 73 -95
rect 79 -91 80 -89
rect 79 -97 80 -95
rect 86 -91 87 -89
rect 93 -91 94 -89
rect 93 -97 94 -95
rect 103 -91 104 -89
rect 103 -97 104 -95
rect 107 -91 108 -89
rect 107 -97 108 -95
rect 114 -91 115 -89
rect 114 -97 115 -95
rect 121 -91 122 -89
rect 121 -97 122 -95
rect 128 -91 129 -89
rect 128 -97 129 -95
rect 135 -91 136 -89
rect 138 -91 139 -89
rect 145 -91 146 -89
rect 142 -97 143 -95
rect 145 -97 146 -95
rect 149 -91 150 -89
rect 149 -97 150 -95
rect 156 -91 157 -89
rect 156 -97 157 -95
rect 163 -91 164 -89
rect 163 -97 164 -95
rect 170 -97 171 -95
rect 173 -97 174 -95
rect 177 -97 178 -95
rect 180 -97 181 -95
rect 187 -91 188 -89
rect 187 -97 188 -95
rect 191 -91 192 -89
rect 194 -91 195 -89
rect 191 -97 192 -95
rect 194 -97 195 -95
rect 198 -91 199 -89
rect 201 -97 202 -95
rect 205 -91 206 -89
rect 208 -91 209 -89
rect 205 -97 206 -95
rect 208 -97 209 -95
rect 212 -91 213 -89
rect 212 -97 213 -95
rect 219 -91 220 -89
rect 219 -97 220 -95
rect 226 -91 227 -89
rect 226 -97 227 -95
rect 236 -91 237 -89
rect 236 -97 237 -95
rect 243 -91 244 -89
rect 240 -97 241 -95
rect 243 -97 244 -95
rect 250 -91 251 -89
rect 247 -97 248 -95
rect 250 -97 251 -95
rect 254 -91 255 -89
rect 257 -91 258 -89
rect 254 -97 255 -95
rect 257 -97 258 -95
rect 261 -91 262 -89
rect 261 -97 262 -95
rect 268 -91 269 -89
rect 268 -97 269 -95
rect 275 -91 276 -89
rect 275 -97 276 -95
rect 282 -91 283 -89
rect 282 -97 283 -95
rect 289 -91 290 -89
rect 289 -97 290 -95
rect 296 -91 297 -89
rect 296 -97 297 -95
rect 303 -91 304 -89
rect 303 -97 304 -95
rect 310 -91 311 -89
rect 310 -97 311 -95
rect 317 -91 318 -89
rect 317 -97 318 -95
rect 324 -91 325 -89
rect 324 -97 325 -95
rect 331 -91 332 -89
rect 331 -97 332 -95
rect 338 -91 339 -89
rect 338 -97 339 -95
rect 345 -91 346 -89
rect 345 -97 346 -95
rect 352 -91 353 -89
rect 352 -97 353 -95
rect 366 -91 367 -89
rect 366 -97 367 -95
rect 376 -91 377 -89
rect 373 -97 374 -95
rect 376 -97 377 -95
rect 86 -134 87 -132
rect 86 -140 87 -138
rect 93 -134 94 -132
rect 93 -140 94 -138
rect 100 -134 101 -132
rect 100 -140 101 -138
rect 107 -134 108 -132
rect 107 -140 108 -138
rect 117 -140 118 -138
rect 121 -134 122 -132
rect 124 -140 125 -138
rect 128 -134 129 -132
rect 128 -140 129 -138
rect 135 -134 136 -132
rect 135 -140 136 -138
rect 142 -134 143 -132
rect 145 -134 146 -132
rect 142 -140 143 -138
rect 149 -134 150 -132
rect 149 -140 150 -138
rect 156 -134 157 -132
rect 163 -134 164 -132
rect 163 -140 164 -138
rect 170 -134 171 -132
rect 170 -140 171 -138
rect 173 -140 174 -138
rect 180 -134 181 -132
rect 184 -134 185 -132
rect 184 -140 185 -138
rect 191 -134 192 -132
rect 194 -134 195 -132
rect 198 -134 199 -132
rect 198 -140 199 -138
rect 205 -134 206 -132
rect 208 -134 209 -132
rect 205 -140 206 -138
rect 212 -134 213 -132
rect 212 -140 213 -138
rect 219 -134 220 -132
rect 219 -140 220 -138
rect 226 -134 227 -132
rect 229 -140 230 -138
rect 236 -134 237 -132
rect 236 -140 237 -138
rect 240 -134 241 -132
rect 240 -140 241 -138
rect 250 -134 251 -132
rect 247 -140 248 -138
rect 254 -134 255 -132
rect 254 -140 255 -138
rect 261 -134 262 -132
rect 264 -134 265 -132
rect 264 -140 265 -138
rect 271 -134 272 -132
rect 275 -134 276 -132
rect 275 -140 276 -138
rect 282 -140 283 -138
rect 289 -134 290 -132
rect 289 -140 290 -138
rect 296 -134 297 -132
rect 296 -140 297 -138
rect 303 -134 304 -132
rect 303 -140 304 -138
rect 310 -134 311 -132
rect 310 -140 311 -138
rect 317 -134 318 -132
rect 317 -140 318 -138
rect 324 -134 325 -132
rect 324 -140 325 -138
rect 331 -134 332 -132
rect 331 -140 332 -138
rect 338 -134 339 -132
rect 341 -140 342 -138
rect 345 -134 346 -132
rect 345 -140 346 -138
rect 355 -140 356 -138
rect 366 -134 367 -132
rect 366 -140 367 -138
rect 380 -134 381 -132
rect 380 -140 381 -138
rect 394 -134 395 -132
rect 394 -140 395 -138
rect 401 -134 402 -132
rect 401 -140 402 -138
rect 65 -169 66 -167
rect 65 -175 66 -173
rect 72 -169 73 -167
rect 72 -175 73 -173
rect 79 -175 80 -173
rect 82 -175 83 -173
rect 86 -169 87 -167
rect 86 -175 87 -173
rect 93 -169 94 -167
rect 93 -175 94 -173
rect 100 -169 101 -167
rect 100 -175 101 -173
rect 107 -169 108 -167
rect 107 -175 108 -173
rect 117 -169 118 -167
rect 114 -175 115 -173
rect 121 -169 122 -167
rect 121 -175 122 -173
rect 128 -169 129 -167
rect 131 -175 132 -173
rect 135 -169 136 -167
rect 135 -175 136 -173
rect 138 -175 139 -173
rect 142 -169 143 -167
rect 142 -175 143 -173
rect 145 -175 146 -173
rect 149 -169 150 -167
rect 152 -169 153 -167
rect 156 -169 157 -167
rect 156 -175 157 -173
rect 163 -169 164 -167
rect 163 -175 164 -173
rect 170 -169 171 -167
rect 170 -175 171 -173
rect 177 -169 178 -167
rect 180 -175 181 -173
rect 184 -169 185 -167
rect 184 -175 185 -173
rect 191 -169 192 -167
rect 191 -175 192 -173
rect 198 -169 199 -167
rect 198 -175 199 -173
rect 201 -175 202 -173
rect 205 -169 206 -167
rect 205 -175 206 -173
rect 212 -169 213 -167
rect 212 -175 213 -173
rect 219 -175 220 -173
rect 222 -175 223 -173
rect 226 -169 227 -167
rect 229 -169 230 -167
rect 233 -169 234 -167
rect 233 -175 234 -173
rect 243 -169 244 -167
rect 240 -175 241 -173
rect 243 -175 244 -173
rect 247 -169 248 -167
rect 247 -175 248 -173
rect 254 -169 255 -167
rect 254 -175 255 -173
rect 261 -169 262 -167
rect 261 -175 262 -173
rect 268 -169 269 -167
rect 268 -175 269 -173
rect 275 -169 276 -167
rect 275 -175 276 -173
rect 285 -169 286 -167
rect 285 -175 286 -173
rect 289 -169 290 -167
rect 289 -175 290 -173
rect 296 -169 297 -167
rect 296 -175 297 -173
rect 303 -169 304 -167
rect 303 -175 304 -173
rect 313 -175 314 -173
rect 317 -169 318 -167
rect 317 -175 318 -173
rect 320 -175 321 -173
rect 324 -169 325 -167
rect 324 -175 325 -173
rect 331 -169 332 -167
rect 331 -175 332 -173
rect 341 -169 342 -167
rect 341 -175 342 -173
rect 345 -169 346 -167
rect 345 -175 346 -173
rect 352 -169 353 -167
rect 352 -175 353 -173
rect 359 -169 360 -167
rect 359 -175 360 -173
rect 366 -169 367 -167
rect 366 -175 367 -173
rect 373 -169 374 -167
rect 380 -169 381 -167
rect 380 -175 381 -173
rect 387 -169 388 -167
rect 387 -175 388 -173
rect 394 -169 395 -167
rect 394 -175 395 -173
rect 401 -169 402 -167
rect 401 -175 402 -173
rect 408 -169 409 -167
rect 408 -175 409 -173
rect 415 -169 416 -167
rect 415 -175 416 -173
rect 422 -169 423 -167
rect 422 -175 423 -173
rect 429 -169 430 -167
rect 432 -175 433 -173
rect 439 -175 440 -173
rect 23 -208 24 -206
rect 23 -214 24 -212
rect 30 -208 31 -206
rect 30 -214 31 -212
rect 37 -208 38 -206
rect 37 -214 38 -212
rect 44 -208 45 -206
rect 44 -214 45 -212
rect 51 -208 52 -206
rect 51 -214 52 -212
rect 58 -214 59 -212
rect 65 -208 66 -206
rect 68 -208 69 -206
rect 65 -214 66 -212
rect 72 -208 73 -206
rect 79 -208 80 -206
rect 79 -214 80 -212
rect 86 -208 87 -206
rect 89 -214 90 -212
rect 96 -208 97 -206
rect 93 -214 94 -212
rect 100 -208 101 -206
rect 100 -214 101 -212
rect 107 -208 108 -206
rect 107 -214 108 -212
rect 114 -208 115 -206
rect 114 -214 115 -212
rect 121 -208 122 -206
rect 121 -214 122 -212
rect 128 -208 129 -206
rect 128 -214 129 -212
rect 135 -208 136 -206
rect 135 -214 136 -212
rect 138 -214 139 -212
rect 142 -208 143 -206
rect 145 -208 146 -206
rect 142 -214 143 -212
rect 145 -214 146 -212
rect 149 -208 150 -206
rect 152 -208 153 -206
rect 156 -208 157 -206
rect 159 -208 160 -206
rect 159 -214 160 -212
rect 163 -208 164 -206
rect 163 -214 164 -212
rect 170 -208 171 -206
rect 170 -214 171 -212
rect 177 -208 178 -206
rect 177 -214 178 -212
rect 184 -208 185 -206
rect 184 -214 185 -212
rect 191 -208 192 -206
rect 194 -208 195 -206
rect 191 -214 192 -212
rect 198 -208 199 -206
rect 201 -214 202 -212
rect 205 -208 206 -206
rect 205 -214 206 -212
rect 208 -214 209 -212
rect 215 -208 216 -206
rect 215 -214 216 -212
rect 219 -208 220 -206
rect 219 -214 220 -212
rect 226 -208 227 -206
rect 226 -214 227 -212
rect 233 -208 234 -206
rect 236 -208 237 -206
rect 236 -214 237 -212
rect 243 -208 244 -206
rect 240 -214 241 -212
rect 243 -214 244 -212
rect 247 -208 248 -206
rect 247 -214 248 -212
rect 254 -208 255 -206
rect 254 -214 255 -212
rect 261 -208 262 -206
rect 261 -214 262 -212
rect 268 -208 269 -206
rect 271 -208 272 -206
rect 268 -214 269 -212
rect 271 -214 272 -212
rect 275 -208 276 -206
rect 275 -214 276 -212
rect 285 -208 286 -206
rect 282 -214 283 -212
rect 289 -208 290 -206
rect 289 -214 290 -212
rect 296 -208 297 -206
rect 299 -214 300 -212
rect 303 -208 304 -206
rect 303 -214 304 -212
rect 310 -208 311 -206
rect 310 -214 311 -212
rect 317 -208 318 -206
rect 317 -214 318 -212
rect 324 -208 325 -206
rect 331 -208 332 -206
rect 331 -214 332 -212
rect 341 -208 342 -206
rect 338 -214 339 -212
rect 345 -208 346 -206
rect 345 -214 346 -212
rect 352 -208 353 -206
rect 352 -214 353 -212
rect 359 -208 360 -206
rect 359 -214 360 -212
rect 366 -208 367 -206
rect 366 -214 367 -212
rect 373 -208 374 -206
rect 380 -208 381 -206
rect 380 -214 381 -212
rect 387 -208 388 -206
rect 387 -214 388 -212
rect 394 -208 395 -206
rect 394 -214 395 -212
rect 401 -208 402 -206
rect 401 -214 402 -212
rect 411 -208 412 -206
rect 408 -214 409 -212
rect 415 -208 416 -206
rect 415 -214 416 -212
rect 422 -208 423 -206
rect 422 -214 423 -212
rect 429 -208 430 -206
rect 429 -214 430 -212
rect 436 -208 437 -206
rect 436 -214 437 -212
rect 443 -208 444 -206
rect 443 -214 444 -212
rect 450 -208 451 -206
rect 450 -214 451 -212
rect 457 -208 458 -206
rect 457 -214 458 -212
rect 464 -208 465 -206
rect 464 -214 465 -212
rect 544 -214 545 -212
rect 37 -255 38 -253
rect 37 -261 38 -259
rect 44 -255 45 -253
rect 44 -261 45 -259
rect 51 -255 52 -253
rect 51 -261 52 -259
rect 58 -255 59 -253
rect 58 -261 59 -259
rect 65 -255 66 -253
rect 65 -261 66 -259
rect 72 -255 73 -253
rect 72 -261 73 -259
rect 75 -261 76 -259
rect 79 -255 80 -253
rect 79 -261 80 -259
rect 86 -255 87 -253
rect 86 -261 87 -259
rect 93 -255 94 -253
rect 93 -261 94 -259
rect 100 -255 101 -253
rect 100 -261 101 -259
rect 110 -255 111 -253
rect 107 -261 108 -259
rect 114 -261 115 -259
rect 117 -261 118 -259
rect 121 -255 122 -253
rect 124 -255 125 -253
rect 128 -261 129 -259
rect 131 -261 132 -259
rect 135 -255 136 -253
rect 135 -261 136 -259
rect 142 -255 143 -253
rect 145 -261 146 -259
rect 149 -255 150 -253
rect 152 -255 153 -253
rect 149 -261 150 -259
rect 152 -261 153 -259
rect 156 -255 157 -253
rect 156 -261 157 -259
rect 163 -255 164 -253
rect 166 -255 167 -253
rect 166 -261 167 -259
rect 170 -255 171 -253
rect 173 -261 174 -259
rect 177 -255 178 -253
rect 180 -255 181 -253
rect 177 -261 178 -259
rect 184 -255 185 -253
rect 184 -261 185 -259
rect 191 -255 192 -253
rect 191 -261 192 -259
rect 198 -255 199 -253
rect 201 -255 202 -253
rect 205 -255 206 -253
rect 208 -255 209 -253
rect 205 -261 206 -259
rect 208 -261 209 -259
rect 212 -255 213 -253
rect 212 -261 213 -259
rect 219 -255 220 -253
rect 219 -261 220 -259
rect 226 -255 227 -253
rect 229 -255 230 -253
rect 226 -261 227 -259
rect 229 -261 230 -259
rect 233 -255 234 -253
rect 240 -255 241 -253
rect 243 -255 244 -253
rect 243 -261 244 -259
rect 247 -255 248 -253
rect 247 -261 248 -259
rect 254 -255 255 -253
rect 254 -261 255 -259
rect 261 -255 262 -253
rect 261 -261 262 -259
rect 268 -255 269 -253
rect 268 -261 269 -259
rect 275 -255 276 -253
rect 275 -261 276 -259
rect 282 -255 283 -253
rect 285 -255 286 -253
rect 282 -261 283 -259
rect 289 -255 290 -253
rect 289 -261 290 -259
rect 296 -255 297 -253
rect 296 -261 297 -259
rect 306 -255 307 -253
rect 303 -261 304 -259
rect 310 -255 311 -253
rect 310 -261 311 -259
rect 317 -255 318 -253
rect 317 -261 318 -259
rect 324 -255 325 -253
rect 327 -255 328 -253
rect 331 -255 332 -253
rect 331 -261 332 -259
rect 334 -261 335 -259
rect 338 -255 339 -253
rect 341 -255 342 -253
rect 338 -261 339 -259
rect 348 -255 349 -253
rect 345 -261 346 -259
rect 348 -261 349 -259
rect 355 -255 356 -253
rect 352 -261 353 -259
rect 359 -255 360 -253
rect 359 -261 360 -259
rect 366 -255 367 -253
rect 366 -261 367 -259
rect 373 -255 374 -253
rect 373 -261 374 -259
rect 380 -255 381 -253
rect 380 -261 381 -259
rect 387 -255 388 -253
rect 387 -261 388 -259
rect 394 -255 395 -253
rect 394 -261 395 -259
rect 401 -255 402 -253
rect 401 -261 402 -259
rect 408 -255 409 -253
rect 408 -261 409 -259
rect 415 -255 416 -253
rect 415 -261 416 -259
rect 422 -255 423 -253
rect 422 -261 423 -259
rect 429 -255 430 -253
rect 429 -261 430 -259
rect 436 -255 437 -253
rect 436 -261 437 -259
rect 443 -255 444 -253
rect 443 -261 444 -259
rect 450 -255 451 -253
rect 450 -261 451 -259
rect 457 -255 458 -253
rect 457 -261 458 -259
rect 464 -255 465 -253
rect 464 -261 465 -259
rect 471 -255 472 -253
rect 471 -261 472 -259
rect 478 -255 479 -253
rect 478 -261 479 -259
rect 485 -255 486 -253
rect 485 -261 486 -259
rect 492 -255 493 -253
rect 492 -261 493 -259
rect 499 -255 500 -253
rect 499 -261 500 -259
rect 506 -255 507 -253
rect 506 -261 507 -259
rect 513 -255 514 -253
rect 513 -261 514 -259
rect 520 -255 521 -253
rect 520 -261 521 -259
rect 527 -261 528 -259
rect 534 -255 535 -253
rect 537 -255 538 -253
rect 534 -261 535 -259
rect 541 -255 542 -253
rect 541 -261 542 -259
rect 37 -302 38 -300
rect 37 -308 38 -306
rect 44 -308 45 -306
rect 51 -302 52 -300
rect 51 -308 52 -306
rect 61 -308 62 -306
rect 65 -302 66 -300
rect 65 -308 66 -306
rect 72 -302 73 -300
rect 72 -308 73 -306
rect 79 -302 80 -300
rect 86 -302 87 -300
rect 86 -308 87 -306
rect 96 -302 97 -300
rect 96 -308 97 -306
rect 100 -302 101 -300
rect 100 -308 101 -306
rect 107 -302 108 -300
rect 107 -308 108 -306
rect 114 -302 115 -300
rect 117 -302 118 -300
rect 114 -308 115 -306
rect 121 -302 122 -300
rect 121 -308 122 -306
rect 128 -302 129 -300
rect 131 -308 132 -306
rect 135 -302 136 -300
rect 135 -308 136 -306
rect 142 -302 143 -300
rect 142 -308 143 -306
rect 149 -302 150 -300
rect 149 -308 150 -306
rect 156 -302 157 -300
rect 156 -308 157 -306
rect 163 -302 164 -300
rect 163 -308 164 -306
rect 170 -302 171 -300
rect 170 -308 171 -306
rect 177 -302 178 -300
rect 177 -308 178 -306
rect 184 -302 185 -300
rect 184 -308 185 -306
rect 191 -302 192 -300
rect 191 -308 192 -306
rect 194 -308 195 -306
rect 198 -302 199 -300
rect 198 -308 199 -306
rect 205 -302 206 -300
rect 205 -308 206 -306
rect 212 -302 213 -300
rect 212 -308 213 -306
rect 219 -302 220 -300
rect 219 -308 220 -306
rect 226 -302 227 -300
rect 226 -308 227 -306
rect 233 -302 234 -300
rect 233 -308 234 -306
rect 240 -302 241 -300
rect 240 -308 241 -306
rect 247 -302 248 -300
rect 247 -308 248 -306
rect 250 -308 251 -306
rect 254 -302 255 -300
rect 254 -308 255 -306
rect 261 -302 262 -300
rect 261 -308 262 -306
rect 268 -302 269 -300
rect 268 -308 269 -306
rect 271 -308 272 -306
rect 275 -302 276 -300
rect 275 -308 276 -306
rect 285 -302 286 -300
rect 282 -308 283 -306
rect 285 -308 286 -306
rect 289 -302 290 -300
rect 289 -308 290 -306
rect 296 -302 297 -300
rect 296 -308 297 -306
rect 303 -302 304 -300
rect 306 -302 307 -300
rect 303 -308 304 -306
rect 310 -302 311 -300
rect 310 -308 311 -306
rect 317 -302 318 -300
rect 320 -302 321 -300
rect 317 -308 318 -306
rect 324 -302 325 -300
rect 324 -308 325 -306
rect 334 -302 335 -300
rect 334 -308 335 -306
rect 338 -308 339 -306
rect 345 -308 346 -306
rect 348 -308 349 -306
rect 352 -302 353 -300
rect 352 -308 353 -306
rect 362 -302 363 -300
rect 366 -302 367 -300
rect 366 -308 367 -306
rect 373 -302 374 -300
rect 373 -308 374 -306
rect 383 -302 384 -300
rect 383 -308 384 -306
rect 387 -302 388 -300
rect 387 -308 388 -306
rect 394 -302 395 -300
rect 394 -308 395 -306
rect 401 -302 402 -300
rect 401 -308 402 -306
rect 408 -302 409 -300
rect 408 -308 409 -306
rect 415 -302 416 -300
rect 415 -308 416 -306
rect 422 -302 423 -300
rect 422 -308 423 -306
rect 429 -302 430 -300
rect 429 -308 430 -306
rect 436 -302 437 -300
rect 436 -308 437 -306
rect 443 -302 444 -300
rect 443 -308 444 -306
rect 450 -302 451 -300
rect 450 -308 451 -306
rect 457 -302 458 -300
rect 457 -308 458 -306
rect 464 -308 465 -306
rect 471 -302 472 -300
rect 471 -308 472 -306
rect 478 -302 479 -300
rect 478 -308 479 -306
rect 485 -302 486 -300
rect 485 -308 486 -306
rect 492 -302 493 -300
rect 492 -308 493 -306
rect 499 -302 500 -300
rect 499 -308 500 -306
rect 506 -302 507 -300
rect 506 -308 507 -306
rect 513 -302 514 -300
rect 513 -308 514 -306
rect 520 -302 521 -300
rect 520 -308 521 -306
rect 527 -302 528 -300
rect 527 -308 528 -306
rect 534 -302 535 -300
rect 534 -308 535 -306
rect 541 -302 542 -300
rect 541 -308 542 -306
rect 544 -308 545 -306
rect 548 -302 549 -300
rect 548 -308 549 -306
rect 555 -302 556 -300
rect 562 -302 563 -300
rect 569 -308 570 -306
rect 576 -302 577 -300
rect 576 -308 577 -306
rect 9 -363 10 -361
rect 9 -369 10 -367
rect 16 -363 17 -361
rect 16 -369 17 -367
rect 23 -363 24 -361
rect 23 -369 24 -367
rect 30 -363 31 -361
rect 30 -369 31 -367
rect 37 -369 38 -367
rect 44 -363 45 -361
rect 44 -369 45 -367
rect 51 -363 52 -361
rect 51 -369 52 -367
rect 61 -363 62 -361
rect 58 -369 59 -367
rect 61 -369 62 -367
rect 65 -363 66 -361
rect 65 -369 66 -367
rect 72 -363 73 -361
rect 72 -369 73 -367
rect 79 -363 80 -361
rect 79 -369 80 -367
rect 86 -363 87 -361
rect 86 -369 87 -367
rect 93 -363 94 -361
rect 93 -369 94 -367
rect 103 -363 104 -361
rect 103 -369 104 -367
rect 107 -369 108 -367
rect 114 -363 115 -361
rect 114 -369 115 -367
rect 121 -363 122 -361
rect 124 -369 125 -367
rect 128 -369 129 -367
rect 131 -369 132 -367
rect 138 -363 139 -361
rect 135 -369 136 -367
rect 138 -369 139 -367
rect 142 -363 143 -361
rect 142 -369 143 -367
rect 149 -363 150 -361
rect 149 -369 150 -367
rect 152 -369 153 -367
rect 156 -363 157 -361
rect 156 -369 157 -367
rect 163 -363 164 -361
rect 163 -369 164 -367
rect 170 -363 171 -361
rect 170 -369 171 -367
rect 180 -363 181 -361
rect 177 -369 178 -367
rect 184 -363 185 -361
rect 184 -369 185 -367
rect 194 -363 195 -361
rect 191 -369 192 -367
rect 198 -363 199 -361
rect 198 -369 199 -367
rect 205 -363 206 -361
rect 208 -363 209 -361
rect 208 -369 209 -367
rect 212 -363 213 -361
rect 212 -369 213 -367
rect 219 -363 220 -361
rect 219 -369 220 -367
rect 226 -363 227 -361
rect 226 -369 227 -367
rect 233 -363 234 -361
rect 233 -369 234 -367
rect 240 -363 241 -361
rect 243 -369 244 -367
rect 247 -363 248 -361
rect 247 -369 248 -367
rect 254 -363 255 -361
rect 254 -369 255 -367
rect 261 -363 262 -361
rect 261 -369 262 -367
rect 268 -363 269 -361
rect 271 -369 272 -367
rect 275 -363 276 -361
rect 275 -369 276 -367
rect 282 -363 283 -361
rect 285 -363 286 -361
rect 285 -369 286 -367
rect 289 -363 290 -361
rect 292 -363 293 -361
rect 296 -363 297 -361
rect 299 -363 300 -361
rect 296 -369 297 -367
rect 299 -369 300 -367
rect 303 -363 304 -361
rect 303 -369 304 -367
rect 310 -363 311 -361
rect 313 -363 314 -361
rect 313 -369 314 -367
rect 317 -363 318 -361
rect 317 -369 318 -367
rect 324 -369 325 -367
rect 327 -369 328 -367
rect 331 -363 332 -361
rect 334 -363 335 -361
rect 338 -363 339 -361
rect 341 -363 342 -361
rect 345 -363 346 -361
rect 348 -363 349 -361
rect 345 -369 346 -367
rect 348 -369 349 -367
rect 352 -363 353 -361
rect 355 -363 356 -361
rect 355 -369 356 -367
rect 359 -363 360 -361
rect 359 -369 360 -367
rect 366 -369 367 -367
rect 373 -363 374 -361
rect 373 -369 374 -367
rect 380 -363 381 -361
rect 380 -369 381 -367
rect 387 -363 388 -361
rect 387 -369 388 -367
rect 394 -363 395 -361
rect 394 -369 395 -367
rect 401 -363 402 -361
rect 401 -369 402 -367
rect 408 -363 409 -361
rect 408 -369 409 -367
rect 415 -363 416 -361
rect 415 -369 416 -367
rect 422 -363 423 -361
rect 422 -369 423 -367
rect 429 -363 430 -361
rect 429 -369 430 -367
rect 436 -363 437 -361
rect 436 -369 437 -367
rect 443 -363 444 -361
rect 443 -369 444 -367
rect 450 -363 451 -361
rect 450 -369 451 -367
rect 457 -363 458 -361
rect 457 -369 458 -367
rect 464 -363 465 -361
rect 464 -369 465 -367
rect 471 -363 472 -361
rect 471 -369 472 -367
rect 478 -363 479 -361
rect 478 -369 479 -367
rect 485 -363 486 -361
rect 485 -369 486 -367
rect 492 -363 493 -361
rect 492 -369 493 -367
rect 499 -363 500 -361
rect 499 -369 500 -367
rect 506 -363 507 -361
rect 506 -369 507 -367
rect 513 -363 514 -361
rect 513 -369 514 -367
rect 520 -363 521 -361
rect 520 -369 521 -367
rect 527 -363 528 -361
rect 527 -369 528 -367
rect 534 -363 535 -361
rect 534 -369 535 -367
rect 541 -363 542 -361
rect 541 -369 542 -367
rect 548 -363 549 -361
rect 548 -369 549 -367
rect 555 -363 556 -361
rect 558 -369 559 -367
rect 562 -363 563 -361
rect 562 -369 563 -367
rect 569 -363 570 -361
rect 569 -369 570 -367
rect 576 -363 577 -361
rect 576 -369 577 -367
rect 2 -418 3 -416
rect 2 -424 3 -422
rect 9 -418 10 -416
rect 19 -424 20 -422
rect 23 -418 24 -416
rect 23 -424 24 -422
rect 33 -418 34 -416
rect 37 -418 38 -416
rect 37 -424 38 -422
rect 44 -418 45 -416
rect 44 -424 45 -422
rect 51 -418 52 -416
rect 51 -424 52 -422
rect 58 -418 59 -416
rect 58 -424 59 -422
rect 68 -418 69 -416
rect 72 -418 73 -416
rect 72 -424 73 -422
rect 79 -418 80 -416
rect 79 -424 80 -422
rect 86 -424 87 -422
rect 96 -418 97 -416
rect 93 -424 94 -422
rect 96 -424 97 -422
rect 100 -418 101 -416
rect 107 -418 108 -416
rect 107 -424 108 -422
rect 114 -418 115 -416
rect 114 -424 115 -422
rect 121 -418 122 -416
rect 121 -424 122 -422
rect 131 -424 132 -422
rect 138 -418 139 -416
rect 135 -424 136 -422
rect 138 -424 139 -422
rect 142 -418 143 -416
rect 142 -424 143 -422
rect 149 -418 150 -416
rect 152 -418 153 -416
rect 156 -418 157 -416
rect 156 -424 157 -422
rect 159 -424 160 -422
rect 163 -418 164 -416
rect 163 -424 164 -422
rect 170 -418 171 -416
rect 170 -424 171 -422
rect 177 -418 178 -416
rect 177 -424 178 -422
rect 184 -418 185 -416
rect 184 -424 185 -422
rect 191 -418 192 -416
rect 191 -424 192 -422
rect 201 -418 202 -416
rect 198 -424 199 -422
rect 205 -418 206 -416
rect 205 -424 206 -422
rect 208 -424 209 -422
rect 212 -418 213 -416
rect 212 -424 213 -422
rect 219 -418 220 -416
rect 219 -424 220 -422
rect 226 -418 227 -416
rect 226 -424 227 -422
rect 233 -418 234 -416
rect 233 -424 234 -422
rect 243 -418 244 -416
rect 240 -424 241 -422
rect 243 -424 244 -422
rect 247 -418 248 -416
rect 250 -418 251 -416
rect 250 -424 251 -422
rect 254 -424 255 -422
rect 257 -424 258 -422
rect 261 -418 262 -416
rect 261 -424 262 -422
rect 268 -418 269 -416
rect 268 -424 269 -422
rect 271 -424 272 -422
rect 275 -418 276 -416
rect 275 -424 276 -422
rect 278 -424 279 -422
rect 282 -418 283 -416
rect 282 -424 283 -422
rect 289 -424 290 -422
rect 296 -418 297 -416
rect 296 -424 297 -422
rect 306 -418 307 -416
rect 310 -418 311 -416
rect 310 -424 311 -422
rect 320 -418 321 -416
rect 317 -424 318 -422
rect 320 -424 321 -422
rect 327 -418 328 -416
rect 324 -424 325 -422
rect 327 -424 328 -422
rect 331 -418 332 -416
rect 331 -424 332 -422
rect 338 -418 339 -416
rect 338 -424 339 -422
rect 348 -418 349 -416
rect 348 -424 349 -422
rect 352 -418 353 -416
rect 352 -424 353 -422
rect 359 -424 360 -422
rect 362 -424 363 -422
rect 366 -418 367 -416
rect 366 -424 367 -422
rect 373 -418 374 -416
rect 373 -424 374 -422
rect 380 -418 381 -416
rect 383 -418 384 -416
rect 380 -424 381 -422
rect 383 -424 384 -422
rect 387 -418 388 -416
rect 390 -418 391 -416
rect 394 -418 395 -416
rect 394 -424 395 -422
rect 401 -418 402 -416
rect 401 -424 402 -422
rect 408 -418 409 -416
rect 411 -418 412 -416
rect 415 -418 416 -416
rect 415 -424 416 -422
rect 422 -418 423 -416
rect 422 -424 423 -422
rect 429 -418 430 -416
rect 429 -424 430 -422
rect 436 -418 437 -416
rect 436 -424 437 -422
rect 443 -418 444 -416
rect 443 -424 444 -422
rect 450 -418 451 -416
rect 450 -424 451 -422
rect 457 -418 458 -416
rect 457 -424 458 -422
rect 464 -418 465 -416
rect 464 -424 465 -422
rect 471 -418 472 -416
rect 471 -424 472 -422
rect 478 -418 479 -416
rect 478 -424 479 -422
rect 485 -418 486 -416
rect 485 -424 486 -422
rect 492 -418 493 -416
rect 492 -424 493 -422
rect 499 -418 500 -416
rect 499 -424 500 -422
rect 506 -418 507 -416
rect 506 -424 507 -422
rect 513 -418 514 -416
rect 513 -424 514 -422
rect 523 -418 524 -416
rect 527 -418 528 -416
rect 527 -424 528 -422
rect 534 -418 535 -416
rect 534 -424 535 -422
rect 541 -418 542 -416
rect 541 -424 542 -422
rect 548 -418 549 -416
rect 548 -424 549 -422
rect 555 -418 556 -416
rect 555 -424 556 -422
rect 562 -418 563 -416
rect 562 -424 563 -422
rect 569 -418 570 -416
rect 569 -424 570 -422
rect 576 -418 577 -416
rect 576 -424 577 -422
rect 583 -418 584 -416
rect 583 -424 584 -422
rect 611 -418 612 -416
rect 611 -424 612 -422
rect 2 -495 3 -493
rect 2 -501 3 -499
rect 9 -495 10 -493
rect 9 -501 10 -499
rect 16 -495 17 -493
rect 16 -501 17 -499
rect 23 -495 24 -493
rect 23 -501 24 -499
rect 30 -495 31 -493
rect 30 -501 31 -499
rect 37 -495 38 -493
rect 40 -495 41 -493
rect 44 -495 45 -493
rect 47 -495 48 -493
rect 47 -501 48 -499
rect 51 -495 52 -493
rect 51 -501 52 -499
rect 58 -495 59 -493
rect 58 -501 59 -499
rect 68 -495 69 -493
rect 72 -495 73 -493
rect 72 -501 73 -499
rect 79 -495 80 -493
rect 79 -501 80 -499
rect 86 -495 87 -493
rect 86 -501 87 -499
rect 93 -495 94 -493
rect 93 -501 94 -499
rect 100 -495 101 -493
rect 100 -501 101 -499
rect 107 -495 108 -493
rect 107 -501 108 -499
rect 114 -495 115 -493
rect 117 -495 118 -493
rect 124 -495 125 -493
rect 124 -501 125 -499
rect 128 -495 129 -493
rect 131 -495 132 -493
rect 128 -501 129 -499
rect 131 -501 132 -499
rect 135 -495 136 -493
rect 138 -495 139 -493
rect 142 -495 143 -493
rect 145 -495 146 -493
rect 142 -501 143 -499
rect 149 -495 150 -493
rect 149 -501 150 -499
rect 156 -495 157 -493
rect 156 -501 157 -499
rect 163 -495 164 -493
rect 163 -501 164 -499
rect 170 -495 171 -493
rect 173 -495 174 -493
rect 170 -501 171 -499
rect 177 -495 178 -493
rect 177 -501 178 -499
rect 187 -495 188 -493
rect 191 -495 192 -493
rect 191 -501 192 -499
rect 201 -495 202 -493
rect 198 -501 199 -499
rect 205 -501 206 -499
rect 208 -501 209 -499
rect 212 -495 213 -493
rect 212 -501 213 -499
rect 219 -495 220 -493
rect 219 -501 220 -499
rect 226 -495 227 -493
rect 226 -501 227 -499
rect 233 -495 234 -493
rect 236 -501 237 -499
rect 243 -495 244 -493
rect 240 -501 241 -499
rect 247 -495 248 -493
rect 247 -501 248 -499
rect 254 -495 255 -493
rect 254 -501 255 -499
rect 264 -495 265 -493
rect 268 -495 269 -493
rect 268 -501 269 -499
rect 275 -495 276 -493
rect 275 -501 276 -499
rect 282 -495 283 -493
rect 282 -501 283 -499
rect 289 -495 290 -493
rect 289 -501 290 -499
rect 296 -495 297 -493
rect 296 -501 297 -499
rect 303 -495 304 -493
rect 303 -501 304 -499
rect 306 -501 307 -499
rect 310 -495 311 -493
rect 313 -495 314 -493
rect 310 -501 311 -499
rect 313 -501 314 -499
rect 317 -495 318 -493
rect 317 -501 318 -499
rect 324 -495 325 -493
rect 327 -495 328 -493
rect 324 -501 325 -499
rect 331 -495 332 -493
rect 334 -495 335 -493
rect 331 -501 332 -499
rect 334 -501 335 -499
rect 338 -495 339 -493
rect 338 -501 339 -499
rect 345 -495 346 -493
rect 345 -501 346 -499
rect 352 -495 353 -493
rect 355 -495 356 -493
rect 355 -501 356 -499
rect 362 -495 363 -493
rect 362 -501 363 -499
rect 366 -495 367 -493
rect 366 -501 367 -499
rect 373 -495 374 -493
rect 373 -501 374 -499
rect 380 -495 381 -493
rect 380 -501 381 -499
rect 387 -495 388 -493
rect 387 -501 388 -499
rect 394 -495 395 -493
rect 397 -495 398 -493
rect 397 -501 398 -499
rect 401 -495 402 -493
rect 401 -501 402 -499
rect 408 -495 409 -493
rect 408 -501 409 -499
rect 415 -495 416 -493
rect 415 -501 416 -499
rect 422 -495 423 -493
rect 425 -501 426 -499
rect 429 -495 430 -493
rect 429 -501 430 -499
rect 436 -495 437 -493
rect 436 -501 437 -499
rect 443 -495 444 -493
rect 443 -501 444 -499
rect 450 -495 451 -493
rect 450 -501 451 -499
rect 457 -495 458 -493
rect 457 -501 458 -499
rect 464 -495 465 -493
rect 464 -501 465 -499
rect 471 -495 472 -493
rect 471 -501 472 -499
rect 478 -495 479 -493
rect 478 -501 479 -499
rect 485 -495 486 -493
rect 485 -501 486 -499
rect 492 -501 493 -499
rect 495 -501 496 -499
rect 499 -495 500 -493
rect 499 -501 500 -499
rect 506 -495 507 -493
rect 506 -501 507 -499
rect 513 -495 514 -493
rect 513 -501 514 -499
rect 520 -495 521 -493
rect 520 -501 521 -499
rect 527 -495 528 -493
rect 527 -501 528 -499
rect 534 -495 535 -493
rect 534 -501 535 -499
rect 541 -495 542 -493
rect 541 -501 542 -499
rect 548 -495 549 -493
rect 548 -501 549 -499
rect 555 -495 556 -493
rect 555 -501 556 -499
rect 562 -495 563 -493
rect 562 -501 563 -499
rect 569 -495 570 -493
rect 569 -501 570 -499
rect 576 -495 577 -493
rect 576 -501 577 -499
rect 583 -495 584 -493
rect 583 -501 584 -499
rect 590 -495 591 -493
rect 590 -501 591 -499
rect 597 -495 598 -493
rect 597 -501 598 -499
rect 604 -495 605 -493
rect 604 -501 605 -499
rect 611 -495 612 -493
rect 611 -501 612 -499
rect 621 -495 622 -493
rect 618 -501 619 -499
rect 621 -501 622 -499
rect 625 -495 626 -493
rect 625 -501 626 -499
rect 635 -495 636 -493
rect 632 -501 633 -499
rect 635 -501 636 -499
rect 639 -495 640 -493
rect 639 -501 640 -499
rect 646 -495 647 -493
rect 646 -501 647 -499
rect 653 -501 654 -499
rect 663 -495 664 -493
rect 667 -495 668 -493
rect 667 -501 668 -499
rect 674 -495 675 -493
rect 674 -501 675 -499
rect 16 -560 17 -558
rect 16 -566 17 -564
rect 23 -560 24 -558
rect 23 -566 24 -564
rect 30 -560 31 -558
rect 30 -566 31 -564
rect 37 -560 38 -558
rect 37 -566 38 -564
rect 44 -566 45 -564
rect 51 -560 52 -558
rect 51 -566 52 -564
rect 61 -560 62 -558
rect 58 -566 59 -564
rect 65 -560 66 -558
rect 65 -566 66 -564
rect 75 -560 76 -558
rect 72 -566 73 -564
rect 79 -566 80 -564
rect 82 -566 83 -564
rect 86 -560 87 -558
rect 86 -566 87 -564
rect 93 -560 94 -558
rect 93 -566 94 -564
rect 100 -560 101 -558
rect 100 -566 101 -564
rect 107 -560 108 -558
rect 107 -566 108 -564
rect 114 -560 115 -558
rect 114 -566 115 -564
rect 121 -560 122 -558
rect 121 -566 122 -564
rect 131 -560 132 -558
rect 135 -560 136 -558
rect 135 -566 136 -564
rect 145 -560 146 -558
rect 142 -566 143 -564
rect 149 -560 150 -558
rect 152 -560 153 -558
rect 149 -566 150 -564
rect 152 -566 153 -564
rect 156 -560 157 -558
rect 156 -566 157 -564
rect 163 -560 164 -558
rect 163 -566 164 -564
rect 170 -560 171 -558
rect 173 -560 174 -558
rect 170 -566 171 -564
rect 177 -560 178 -558
rect 177 -566 178 -564
rect 184 -560 185 -558
rect 184 -566 185 -564
rect 191 -560 192 -558
rect 191 -566 192 -564
rect 194 -566 195 -564
rect 198 -560 199 -558
rect 198 -566 199 -564
rect 205 -560 206 -558
rect 208 -560 209 -558
rect 205 -566 206 -564
rect 212 -560 213 -558
rect 212 -566 213 -564
rect 219 -560 220 -558
rect 219 -566 220 -564
rect 226 -560 227 -558
rect 226 -566 227 -564
rect 233 -560 234 -558
rect 233 -566 234 -564
rect 240 -560 241 -558
rect 240 -566 241 -564
rect 247 -560 248 -558
rect 247 -566 248 -564
rect 254 -560 255 -558
rect 254 -566 255 -564
rect 264 -560 265 -558
rect 261 -566 262 -564
rect 264 -566 265 -564
rect 268 -560 269 -558
rect 271 -560 272 -558
rect 268 -566 269 -564
rect 271 -566 272 -564
rect 275 -560 276 -558
rect 278 -560 279 -558
rect 282 -560 283 -558
rect 282 -566 283 -564
rect 289 -560 290 -558
rect 289 -566 290 -564
rect 296 -560 297 -558
rect 296 -566 297 -564
rect 303 -560 304 -558
rect 303 -566 304 -564
rect 310 -560 311 -558
rect 310 -566 311 -564
rect 317 -560 318 -558
rect 317 -566 318 -564
rect 324 -560 325 -558
rect 324 -566 325 -564
rect 334 -560 335 -558
rect 334 -566 335 -564
rect 338 -560 339 -558
rect 338 -566 339 -564
rect 348 -560 349 -558
rect 348 -566 349 -564
rect 352 -560 353 -558
rect 352 -566 353 -564
rect 355 -566 356 -564
rect 359 -560 360 -558
rect 359 -566 360 -564
rect 366 -560 367 -558
rect 369 -560 370 -558
rect 369 -566 370 -564
rect 373 -560 374 -558
rect 373 -566 374 -564
rect 380 -560 381 -558
rect 383 -560 384 -558
rect 383 -566 384 -564
rect 390 -560 391 -558
rect 387 -566 388 -564
rect 394 -560 395 -558
rect 397 -560 398 -558
rect 394 -566 395 -564
rect 401 -566 402 -564
rect 404 -566 405 -564
rect 411 -560 412 -558
rect 408 -566 409 -564
rect 411 -566 412 -564
rect 415 -560 416 -558
rect 415 -566 416 -564
rect 422 -560 423 -558
rect 422 -566 423 -564
rect 429 -560 430 -558
rect 429 -566 430 -564
rect 436 -560 437 -558
rect 436 -566 437 -564
rect 443 -560 444 -558
rect 443 -566 444 -564
rect 450 -560 451 -558
rect 450 -566 451 -564
rect 457 -560 458 -558
rect 457 -566 458 -564
rect 464 -560 465 -558
rect 464 -566 465 -564
rect 471 -560 472 -558
rect 471 -566 472 -564
rect 478 -560 479 -558
rect 478 -566 479 -564
rect 485 -560 486 -558
rect 485 -566 486 -564
rect 492 -560 493 -558
rect 492 -566 493 -564
rect 499 -560 500 -558
rect 499 -566 500 -564
rect 506 -560 507 -558
rect 506 -566 507 -564
rect 513 -560 514 -558
rect 513 -566 514 -564
rect 520 -560 521 -558
rect 520 -566 521 -564
rect 527 -560 528 -558
rect 527 -566 528 -564
rect 534 -560 535 -558
rect 534 -566 535 -564
rect 541 -560 542 -558
rect 541 -566 542 -564
rect 548 -560 549 -558
rect 548 -566 549 -564
rect 555 -560 556 -558
rect 555 -566 556 -564
rect 562 -560 563 -558
rect 562 -566 563 -564
rect 569 -560 570 -558
rect 569 -566 570 -564
rect 576 -560 577 -558
rect 576 -566 577 -564
rect 583 -560 584 -558
rect 583 -566 584 -564
rect 590 -560 591 -558
rect 590 -566 591 -564
rect 597 -560 598 -558
rect 597 -566 598 -564
rect 604 -560 605 -558
rect 604 -566 605 -564
rect 611 -560 612 -558
rect 614 -560 615 -558
rect 618 -560 619 -558
rect 618 -566 619 -564
rect 621 -566 622 -564
rect 625 -560 626 -558
rect 628 -560 629 -558
rect 628 -566 629 -564
rect 632 -560 633 -558
rect 632 -566 633 -564
rect 639 -560 640 -558
rect 642 -560 643 -558
rect 642 -566 643 -564
rect 646 -560 647 -558
rect 646 -566 647 -564
rect 653 -560 654 -558
rect 653 -566 654 -564
rect 2 -615 3 -613
rect 2 -621 3 -619
rect 9 -615 10 -613
rect 9 -621 10 -619
rect 16 -615 17 -613
rect 16 -621 17 -619
rect 23 -615 24 -613
rect 23 -621 24 -619
rect 30 -615 31 -613
rect 30 -621 31 -619
rect 37 -615 38 -613
rect 37 -621 38 -619
rect 44 -615 45 -613
rect 44 -621 45 -619
rect 51 -615 52 -613
rect 51 -621 52 -619
rect 61 -615 62 -613
rect 61 -621 62 -619
rect 68 -615 69 -613
rect 65 -621 66 -619
rect 68 -621 69 -619
rect 72 -615 73 -613
rect 72 -621 73 -619
rect 79 -615 80 -613
rect 79 -621 80 -619
rect 86 -615 87 -613
rect 86 -621 87 -619
rect 93 -615 94 -613
rect 93 -621 94 -619
rect 100 -615 101 -613
rect 103 -615 104 -613
rect 103 -621 104 -619
rect 107 -615 108 -613
rect 107 -621 108 -619
rect 114 -615 115 -613
rect 114 -621 115 -619
rect 121 -615 122 -613
rect 124 -615 125 -613
rect 121 -621 122 -619
rect 128 -615 129 -613
rect 128 -621 129 -619
rect 131 -621 132 -619
rect 135 -615 136 -613
rect 135 -621 136 -619
rect 142 -615 143 -613
rect 142 -621 143 -619
rect 152 -615 153 -613
rect 152 -621 153 -619
rect 156 -615 157 -613
rect 156 -621 157 -619
rect 163 -615 164 -613
rect 163 -621 164 -619
rect 170 -615 171 -613
rect 170 -621 171 -619
rect 177 -615 178 -613
rect 180 -615 181 -613
rect 177 -621 178 -619
rect 180 -621 181 -619
rect 184 -615 185 -613
rect 184 -621 185 -619
rect 191 -615 192 -613
rect 194 -621 195 -619
rect 198 -615 199 -613
rect 201 -615 202 -613
rect 198 -621 199 -619
rect 201 -621 202 -619
rect 205 -615 206 -613
rect 208 -615 209 -613
rect 205 -621 206 -619
rect 208 -621 209 -619
rect 212 -615 213 -613
rect 212 -621 213 -619
rect 219 -615 220 -613
rect 219 -621 220 -619
rect 226 -615 227 -613
rect 229 -615 230 -613
rect 226 -621 227 -619
rect 229 -621 230 -619
rect 233 -615 234 -613
rect 233 -621 234 -619
rect 240 -615 241 -613
rect 240 -621 241 -619
rect 247 -615 248 -613
rect 247 -621 248 -619
rect 257 -615 258 -613
rect 257 -621 258 -619
rect 261 -615 262 -613
rect 261 -621 262 -619
rect 268 -615 269 -613
rect 268 -621 269 -619
rect 278 -615 279 -613
rect 278 -621 279 -619
rect 282 -615 283 -613
rect 282 -621 283 -619
rect 289 -615 290 -613
rect 289 -621 290 -619
rect 296 -615 297 -613
rect 296 -621 297 -619
rect 303 -615 304 -613
rect 303 -621 304 -619
rect 310 -615 311 -613
rect 310 -621 311 -619
rect 313 -621 314 -619
rect 317 -615 318 -613
rect 317 -621 318 -619
rect 324 -615 325 -613
rect 324 -621 325 -619
rect 327 -621 328 -619
rect 331 -615 332 -613
rect 334 -621 335 -619
rect 338 -615 339 -613
rect 338 -621 339 -619
rect 345 -615 346 -613
rect 348 -615 349 -613
rect 345 -621 346 -619
rect 348 -621 349 -619
rect 352 -615 353 -613
rect 355 -621 356 -619
rect 359 -615 360 -613
rect 362 -615 363 -613
rect 362 -621 363 -619
rect 366 -615 367 -613
rect 366 -621 367 -619
rect 373 -615 374 -613
rect 373 -621 374 -619
rect 380 -615 381 -613
rect 380 -621 381 -619
rect 387 -615 388 -613
rect 387 -621 388 -619
rect 394 -615 395 -613
rect 394 -621 395 -619
rect 401 -615 402 -613
rect 404 -621 405 -619
rect 408 -615 409 -613
rect 408 -621 409 -619
rect 415 -615 416 -613
rect 415 -621 416 -619
rect 422 -615 423 -613
rect 422 -621 423 -619
rect 429 -615 430 -613
rect 429 -621 430 -619
rect 436 -615 437 -613
rect 436 -621 437 -619
rect 443 -615 444 -613
rect 443 -621 444 -619
rect 450 -615 451 -613
rect 450 -621 451 -619
rect 457 -621 458 -619
rect 460 -621 461 -619
rect 464 -615 465 -613
rect 464 -621 465 -619
rect 471 -615 472 -613
rect 471 -621 472 -619
rect 478 -615 479 -613
rect 485 -615 486 -613
rect 485 -621 486 -619
rect 492 -615 493 -613
rect 492 -621 493 -619
rect 499 -615 500 -613
rect 499 -621 500 -619
rect 506 -615 507 -613
rect 506 -621 507 -619
rect 513 -615 514 -613
rect 513 -621 514 -619
rect 520 -615 521 -613
rect 520 -621 521 -619
rect 527 -621 528 -619
rect 534 -615 535 -613
rect 534 -621 535 -619
rect 544 -615 545 -613
rect 548 -615 549 -613
rect 548 -621 549 -619
rect 555 -615 556 -613
rect 555 -621 556 -619
rect 565 -615 566 -613
rect 569 -615 570 -613
rect 569 -621 570 -619
rect 576 -615 577 -613
rect 576 -621 577 -619
rect 583 -615 584 -613
rect 583 -621 584 -619
rect 590 -615 591 -613
rect 590 -621 591 -619
rect 597 -615 598 -613
rect 597 -621 598 -619
rect 604 -615 605 -613
rect 604 -621 605 -619
rect 611 -615 612 -613
rect 611 -621 612 -619
rect 618 -615 619 -613
rect 618 -621 619 -619
rect 625 -615 626 -613
rect 625 -621 626 -619
rect 632 -615 633 -613
rect 632 -621 633 -619
rect 653 -615 654 -613
rect 653 -621 654 -619
rect 2 -680 3 -678
rect 2 -686 3 -684
rect 9 -680 10 -678
rect 9 -686 10 -684
rect 16 -680 17 -678
rect 16 -686 17 -684
rect 23 -680 24 -678
rect 30 -680 31 -678
rect 30 -686 31 -684
rect 37 -680 38 -678
rect 37 -686 38 -684
rect 44 -680 45 -678
rect 44 -686 45 -684
rect 51 -680 52 -678
rect 54 -686 55 -684
rect 58 -680 59 -678
rect 58 -686 59 -684
rect 65 -680 66 -678
rect 65 -686 66 -684
rect 72 -680 73 -678
rect 72 -686 73 -684
rect 79 -680 80 -678
rect 79 -686 80 -684
rect 86 -680 87 -678
rect 86 -686 87 -684
rect 96 -680 97 -678
rect 96 -686 97 -684
rect 100 -680 101 -678
rect 100 -686 101 -684
rect 107 -680 108 -678
rect 107 -686 108 -684
rect 114 -686 115 -684
rect 117 -686 118 -684
rect 121 -680 122 -678
rect 121 -686 122 -684
rect 128 -680 129 -678
rect 131 -680 132 -678
rect 128 -686 129 -684
rect 135 -680 136 -678
rect 138 -680 139 -678
rect 142 -680 143 -678
rect 142 -686 143 -684
rect 149 -680 150 -678
rect 152 -680 153 -678
rect 149 -686 150 -684
rect 156 -680 157 -678
rect 156 -686 157 -684
rect 163 -680 164 -678
rect 163 -686 164 -684
rect 170 -680 171 -678
rect 173 -680 174 -678
rect 173 -686 174 -684
rect 177 -680 178 -678
rect 177 -686 178 -684
rect 180 -686 181 -684
rect 184 -680 185 -678
rect 187 -686 188 -684
rect 191 -680 192 -678
rect 191 -686 192 -684
rect 201 -680 202 -678
rect 198 -686 199 -684
rect 201 -686 202 -684
rect 205 -680 206 -678
rect 208 -680 209 -678
rect 205 -686 206 -684
rect 212 -680 213 -678
rect 212 -686 213 -684
rect 219 -680 220 -678
rect 222 -680 223 -678
rect 219 -686 220 -684
rect 226 -680 227 -678
rect 226 -686 227 -684
rect 233 -680 234 -678
rect 233 -686 234 -684
rect 240 -680 241 -678
rect 240 -686 241 -684
rect 247 -680 248 -678
rect 247 -686 248 -684
rect 257 -680 258 -678
rect 254 -686 255 -684
rect 257 -686 258 -684
rect 261 -680 262 -678
rect 261 -686 262 -684
rect 268 -680 269 -678
rect 268 -686 269 -684
rect 275 -680 276 -678
rect 278 -680 279 -678
rect 275 -686 276 -684
rect 278 -686 279 -684
rect 285 -686 286 -684
rect 289 -680 290 -678
rect 292 -686 293 -684
rect 296 -680 297 -678
rect 296 -686 297 -684
rect 303 -680 304 -678
rect 303 -686 304 -684
rect 310 -680 311 -678
rect 313 -680 314 -678
rect 310 -686 311 -684
rect 313 -686 314 -684
rect 317 -680 318 -678
rect 317 -686 318 -684
rect 324 -680 325 -678
rect 324 -686 325 -684
rect 331 -680 332 -678
rect 334 -680 335 -678
rect 331 -686 332 -684
rect 338 -680 339 -678
rect 338 -686 339 -684
rect 345 -680 346 -678
rect 345 -686 346 -684
rect 352 -680 353 -678
rect 352 -686 353 -684
rect 359 -680 360 -678
rect 359 -686 360 -684
rect 369 -680 370 -678
rect 366 -686 367 -684
rect 369 -686 370 -684
rect 373 -680 374 -678
rect 376 -686 377 -684
rect 380 -680 381 -678
rect 380 -686 381 -684
rect 387 -680 388 -678
rect 387 -686 388 -684
rect 394 -680 395 -678
rect 397 -680 398 -678
rect 397 -686 398 -684
rect 401 -680 402 -678
rect 404 -680 405 -678
rect 404 -686 405 -684
rect 408 -680 409 -678
rect 408 -686 409 -684
rect 415 -680 416 -678
rect 415 -686 416 -684
rect 422 -680 423 -678
rect 425 -686 426 -684
rect 429 -680 430 -678
rect 432 -686 433 -684
rect 436 -680 437 -678
rect 436 -686 437 -684
rect 443 -680 444 -678
rect 443 -686 444 -684
rect 450 -680 451 -678
rect 450 -686 451 -684
rect 457 -680 458 -678
rect 457 -686 458 -684
rect 464 -680 465 -678
rect 464 -686 465 -684
rect 471 -680 472 -678
rect 471 -686 472 -684
rect 478 -680 479 -678
rect 478 -686 479 -684
rect 485 -680 486 -678
rect 485 -686 486 -684
rect 492 -680 493 -678
rect 492 -686 493 -684
rect 499 -680 500 -678
rect 499 -686 500 -684
rect 506 -680 507 -678
rect 506 -686 507 -684
rect 513 -680 514 -678
rect 513 -686 514 -684
rect 520 -680 521 -678
rect 520 -686 521 -684
rect 527 -680 528 -678
rect 527 -686 528 -684
rect 534 -680 535 -678
rect 534 -686 535 -684
rect 541 -680 542 -678
rect 541 -686 542 -684
rect 548 -680 549 -678
rect 548 -686 549 -684
rect 555 -680 556 -678
rect 558 -680 559 -678
rect 562 -680 563 -678
rect 565 -680 566 -678
rect 562 -686 563 -684
rect 632 -680 633 -678
rect 632 -686 633 -684
rect 639 -680 640 -678
rect 639 -686 640 -684
rect 653 -680 654 -678
rect 653 -686 654 -684
rect 2 -747 3 -745
rect 2 -753 3 -751
rect 12 -747 13 -745
rect 16 -747 17 -745
rect 23 -753 24 -751
rect 30 -747 31 -745
rect 30 -753 31 -751
rect 37 -747 38 -745
rect 37 -753 38 -751
rect 47 -747 48 -745
rect 51 -747 52 -745
rect 51 -753 52 -751
rect 58 -753 59 -751
rect 61 -753 62 -751
rect 65 -747 66 -745
rect 65 -753 66 -751
rect 72 -747 73 -745
rect 72 -753 73 -751
rect 82 -747 83 -745
rect 82 -753 83 -751
rect 86 -747 87 -745
rect 86 -753 87 -751
rect 93 -747 94 -745
rect 93 -753 94 -751
rect 100 -753 101 -751
rect 103 -753 104 -751
rect 107 -747 108 -745
rect 107 -753 108 -751
rect 114 -747 115 -745
rect 117 -747 118 -745
rect 114 -753 115 -751
rect 117 -753 118 -751
rect 121 -747 122 -745
rect 121 -753 122 -751
rect 128 -747 129 -745
rect 128 -753 129 -751
rect 135 -747 136 -745
rect 135 -753 136 -751
rect 145 -747 146 -745
rect 142 -753 143 -751
rect 145 -753 146 -751
rect 149 -747 150 -745
rect 149 -753 150 -751
rect 152 -753 153 -751
rect 156 -747 157 -745
rect 156 -753 157 -751
rect 166 -747 167 -745
rect 163 -753 164 -751
rect 170 -747 171 -745
rect 170 -753 171 -751
rect 177 -747 178 -745
rect 177 -753 178 -751
rect 184 -747 185 -745
rect 187 -747 188 -745
rect 187 -753 188 -751
rect 191 -747 192 -745
rect 194 -747 195 -745
rect 198 -747 199 -745
rect 198 -753 199 -751
rect 205 -753 206 -751
rect 208 -753 209 -751
rect 212 -747 213 -745
rect 212 -753 213 -751
rect 219 -747 220 -745
rect 219 -753 220 -751
rect 226 -747 227 -745
rect 229 -747 230 -745
rect 229 -753 230 -751
rect 233 -747 234 -745
rect 233 -753 234 -751
rect 240 -747 241 -745
rect 240 -753 241 -751
rect 247 -747 248 -745
rect 247 -753 248 -751
rect 254 -747 255 -745
rect 254 -753 255 -751
rect 261 -747 262 -745
rect 261 -753 262 -751
rect 268 -747 269 -745
rect 271 -747 272 -745
rect 268 -753 269 -751
rect 275 -747 276 -745
rect 278 -747 279 -745
rect 275 -753 276 -751
rect 278 -753 279 -751
rect 282 -747 283 -745
rect 285 -747 286 -745
rect 289 -747 290 -745
rect 289 -753 290 -751
rect 296 -747 297 -745
rect 296 -753 297 -751
rect 306 -747 307 -745
rect 310 -747 311 -745
rect 310 -753 311 -751
rect 317 -747 318 -745
rect 317 -753 318 -751
rect 324 -747 325 -745
rect 324 -753 325 -751
rect 331 -747 332 -745
rect 331 -753 332 -751
rect 338 -747 339 -745
rect 341 -747 342 -745
rect 341 -753 342 -751
rect 345 -747 346 -745
rect 345 -753 346 -751
rect 352 -747 353 -745
rect 355 -747 356 -745
rect 359 -747 360 -745
rect 362 -747 363 -745
rect 359 -753 360 -751
rect 362 -753 363 -751
rect 366 -747 367 -745
rect 366 -753 367 -751
rect 373 -747 374 -745
rect 376 -747 377 -745
rect 373 -753 374 -751
rect 376 -753 377 -751
rect 380 -753 381 -751
rect 387 -747 388 -745
rect 387 -753 388 -751
rect 394 -747 395 -745
rect 394 -753 395 -751
rect 401 -747 402 -745
rect 401 -753 402 -751
rect 408 -753 409 -751
rect 411 -753 412 -751
rect 415 -747 416 -745
rect 415 -753 416 -751
rect 422 -747 423 -745
rect 422 -753 423 -751
rect 429 -747 430 -745
rect 429 -753 430 -751
rect 436 -747 437 -745
rect 436 -753 437 -751
rect 443 -747 444 -745
rect 443 -753 444 -751
rect 450 -747 451 -745
rect 450 -753 451 -751
rect 457 -747 458 -745
rect 457 -753 458 -751
rect 464 -747 465 -745
rect 464 -753 465 -751
rect 471 -753 472 -751
rect 474 -753 475 -751
rect 478 -747 479 -745
rect 478 -753 479 -751
rect 485 -747 486 -745
rect 485 -753 486 -751
rect 492 -747 493 -745
rect 492 -753 493 -751
rect 499 -747 500 -745
rect 499 -753 500 -751
rect 506 -747 507 -745
rect 506 -753 507 -751
rect 513 -747 514 -745
rect 513 -753 514 -751
rect 520 -747 521 -745
rect 520 -753 521 -751
rect 527 -747 528 -745
rect 527 -753 528 -751
rect 534 -747 535 -745
rect 534 -753 535 -751
rect 541 -747 542 -745
rect 541 -753 542 -751
rect 548 -747 549 -745
rect 548 -753 549 -751
rect 555 -747 556 -745
rect 555 -753 556 -751
rect 562 -747 563 -745
rect 562 -753 563 -751
rect 569 -747 570 -745
rect 569 -753 570 -751
rect 576 -747 577 -745
rect 576 -753 577 -751
rect 583 -747 584 -745
rect 583 -753 584 -751
rect 590 -747 591 -745
rect 590 -753 591 -751
rect 597 -747 598 -745
rect 597 -753 598 -751
rect 604 -747 605 -745
rect 604 -753 605 -751
rect 611 -747 612 -745
rect 611 -753 612 -751
rect 618 -747 619 -745
rect 618 -753 619 -751
rect 625 -747 626 -745
rect 625 -753 626 -751
rect 632 -747 633 -745
rect 632 -753 633 -751
rect 639 -747 640 -745
rect 639 -753 640 -751
rect 646 -747 647 -745
rect 646 -753 647 -751
rect 653 -747 654 -745
rect 656 -747 657 -745
rect 653 -753 654 -751
rect 663 -747 664 -745
rect 660 -753 661 -751
rect 23 -820 24 -818
rect 23 -826 24 -824
rect 30 -820 31 -818
rect 30 -826 31 -824
rect 40 -826 41 -824
rect 44 -820 45 -818
rect 44 -826 45 -824
rect 54 -820 55 -818
rect 51 -826 52 -824
rect 54 -826 55 -824
rect 58 -820 59 -818
rect 58 -826 59 -824
rect 65 -820 66 -818
rect 65 -826 66 -824
rect 72 -820 73 -818
rect 72 -826 73 -824
rect 79 -820 80 -818
rect 82 -820 83 -818
rect 82 -826 83 -824
rect 86 -826 87 -824
rect 89 -826 90 -824
rect 96 -820 97 -818
rect 93 -826 94 -824
rect 96 -826 97 -824
rect 100 -820 101 -818
rect 100 -826 101 -824
rect 107 -820 108 -818
rect 107 -826 108 -824
rect 114 -820 115 -818
rect 114 -826 115 -824
rect 121 -820 122 -818
rect 121 -826 122 -824
rect 128 -826 129 -824
rect 135 -826 136 -824
rect 145 -826 146 -824
rect 149 -820 150 -818
rect 152 -820 153 -818
rect 152 -826 153 -824
rect 156 -820 157 -818
rect 156 -826 157 -824
rect 163 -820 164 -818
rect 163 -826 164 -824
rect 170 -820 171 -818
rect 170 -826 171 -824
rect 177 -820 178 -818
rect 177 -826 178 -824
rect 184 -820 185 -818
rect 184 -826 185 -824
rect 191 -820 192 -818
rect 191 -826 192 -824
rect 198 -820 199 -818
rect 198 -826 199 -824
rect 205 -820 206 -818
rect 205 -826 206 -824
rect 212 -820 213 -818
rect 212 -826 213 -824
rect 219 -820 220 -818
rect 219 -826 220 -824
rect 226 -820 227 -818
rect 226 -826 227 -824
rect 233 -820 234 -818
rect 233 -826 234 -824
rect 243 -820 244 -818
rect 247 -820 248 -818
rect 247 -826 248 -824
rect 254 -820 255 -818
rect 254 -826 255 -824
rect 261 -820 262 -818
rect 261 -826 262 -824
rect 268 -820 269 -818
rect 268 -826 269 -824
rect 275 -820 276 -818
rect 278 -820 279 -818
rect 275 -826 276 -824
rect 278 -826 279 -824
rect 282 -820 283 -818
rect 285 -820 286 -818
rect 285 -826 286 -824
rect 289 -820 290 -818
rect 289 -826 290 -824
rect 299 -820 300 -818
rect 296 -826 297 -824
rect 303 -820 304 -818
rect 303 -826 304 -824
rect 310 -820 311 -818
rect 313 -820 314 -818
rect 320 -820 321 -818
rect 317 -826 318 -824
rect 320 -826 321 -824
rect 327 -820 328 -818
rect 331 -820 332 -818
rect 331 -826 332 -824
rect 334 -826 335 -824
rect 338 -820 339 -818
rect 341 -820 342 -818
rect 338 -826 339 -824
rect 345 -820 346 -818
rect 345 -826 346 -824
rect 352 -820 353 -818
rect 355 -826 356 -824
rect 359 -820 360 -818
rect 359 -826 360 -824
rect 366 -820 367 -818
rect 366 -826 367 -824
rect 373 -820 374 -818
rect 376 -820 377 -818
rect 373 -826 374 -824
rect 376 -826 377 -824
rect 380 -820 381 -818
rect 380 -826 381 -824
rect 387 -820 388 -818
rect 390 -820 391 -818
rect 394 -820 395 -818
rect 394 -826 395 -824
rect 401 -826 402 -824
rect 404 -826 405 -824
rect 408 -820 409 -818
rect 408 -826 409 -824
rect 415 -820 416 -818
rect 415 -826 416 -824
rect 422 -820 423 -818
rect 422 -826 423 -824
rect 429 -820 430 -818
rect 429 -826 430 -824
rect 436 -820 437 -818
rect 436 -826 437 -824
rect 443 -820 444 -818
rect 443 -826 444 -824
rect 450 -820 451 -818
rect 450 -826 451 -824
rect 457 -820 458 -818
rect 457 -826 458 -824
rect 464 -820 465 -818
rect 464 -826 465 -824
rect 471 -820 472 -818
rect 471 -826 472 -824
rect 478 -826 479 -824
rect 485 -820 486 -818
rect 485 -826 486 -824
rect 492 -820 493 -818
rect 492 -826 493 -824
rect 499 -820 500 -818
rect 499 -826 500 -824
rect 506 -820 507 -818
rect 506 -826 507 -824
rect 513 -820 514 -818
rect 520 -820 521 -818
rect 520 -826 521 -824
rect 527 -820 528 -818
rect 527 -826 528 -824
rect 537 -820 538 -818
rect 541 -820 542 -818
rect 541 -826 542 -824
rect 548 -820 549 -818
rect 548 -826 549 -824
rect 555 -820 556 -818
rect 558 -820 559 -818
rect 562 -820 563 -818
rect 562 -826 563 -824
rect 569 -820 570 -818
rect 572 -826 573 -824
rect 576 -820 577 -818
rect 576 -826 577 -824
rect 583 -820 584 -818
rect 583 -826 584 -824
rect 590 -820 591 -818
rect 590 -826 591 -824
rect 597 -820 598 -818
rect 604 -820 605 -818
rect 604 -826 605 -824
rect 618 -820 619 -818
rect 618 -826 619 -824
rect 2 -863 3 -861
rect 2 -869 3 -867
rect 9 -863 10 -861
rect 9 -869 10 -867
rect 16 -863 17 -861
rect 16 -869 17 -867
rect 23 -863 24 -861
rect 23 -869 24 -867
rect 33 -863 34 -861
rect 30 -869 31 -867
rect 37 -863 38 -861
rect 37 -869 38 -867
rect 40 -869 41 -867
rect 44 -869 45 -867
rect 47 -869 48 -867
rect 51 -863 52 -861
rect 51 -869 52 -867
rect 61 -863 62 -861
rect 61 -869 62 -867
rect 65 -863 66 -861
rect 65 -869 66 -867
rect 72 -863 73 -861
rect 72 -869 73 -867
rect 79 -869 80 -867
rect 86 -863 87 -861
rect 86 -869 87 -867
rect 93 -863 94 -861
rect 93 -869 94 -867
rect 100 -863 101 -861
rect 100 -869 101 -867
rect 107 -863 108 -861
rect 107 -869 108 -867
rect 114 -863 115 -861
rect 114 -869 115 -867
rect 121 -863 122 -861
rect 121 -869 122 -867
rect 128 -863 129 -861
rect 128 -869 129 -867
rect 135 -863 136 -861
rect 135 -869 136 -867
rect 142 -863 143 -861
rect 149 -863 150 -861
rect 149 -869 150 -867
rect 156 -863 157 -861
rect 156 -869 157 -867
rect 163 -863 164 -861
rect 163 -869 164 -867
rect 170 -863 171 -861
rect 173 -863 174 -861
rect 173 -869 174 -867
rect 180 -863 181 -861
rect 184 -863 185 -861
rect 184 -869 185 -867
rect 191 -863 192 -861
rect 194 -863 195 -861
rect 191 -869 192 -867
rect 198 -863 199 -861
rect 201 -863 202 -861
rect 205 -863 206 -861
rect 205 -869 206 -867
rect 208 -869 209 -867
rect 215 -863 216 -861
rect 222 -863 223 -861
rect 219 -869 220 -867
rect 222 -869 223 -867
rect 226 -863 227 -861
rect 229 -863 230 -861
rect 226 -869 227 -867
rect 233 -863 234 -861
rect 233 -869 234 -867
rect 240 -863 241 -861
rect 240 -869 241 -867
rect 247 -863 248 -861
rect 247 -869 248 -867
rect 254 -863 255 -861
rect 254 -869 255 -867
rect 261 -863 262 -861
rect 268 -863 269 -861
rect 268 -869 269 -867
rect 275 -863 276 -861
rect 275 -869 276 -867
rect 282 -863 283 -861
rect 282 -869 283 -867
rect 289 -863 290 -861
rect 292 -863 293 -861
rect 289 -869 290 -867
rect 292 -869 293 -867
rect 296 -863 297 -861
rect 296 -869 297 -867
rect 303 -863 304 -861
rect 303 -869 304 -867
rect 310 -863 311 -861
rect 310 -869 311 -867
rect 317 -863 318 -861
rect 320 -863 321 -861
rect 320 -869 321 -867
rect 324 -863 325 -861
rect 324 -869 325 -867
rect 331 -863 332 -861
rect 331 -869 332 -867
rect 338 -863 339 -861
rect 338 -869 339 -867
rect 345 -863 346 -861
rect 348 -863 349 -861
rect 348 -869 349 -867
rect 352 -863 353 -861
rect 352 -869 353 -867
rect 359 -863 360 -861
rect 359 -869 360 -867
rect 366 -863 367 -861
rect 366 -869 367 -867
rect 373 -863 374 -861
rect 373 -869 374 -867
rect 376 -869 377 -867
rect 380 -863 381 -861
rect 380 -869 381 -867
rect 387 -863 388 -861
rect 387 -869 388 -867
rect 394 -863 395 -861
rect 394 -869 395 -867
rect 401 -863 402 -861
rect 401 -869 402 -867
rect 408 -863 409 -861
rect 408 -869 409 -867
rect 415 -863 416 -861
rect 415 -869 416 -867
rect 425 -863 426 -861
rect 425 -869 426 -867
rect 429 -863 430 -861
rect 429 -869 430 -867
rect 436 -863 437 -861
rect 436 -869 437 -867
rect 443 -863 444 -861
rect 443 -869 444 -867
rect 450 -869 451 -867
rect 453 -869 454 -867
rect 457 -863 458 -861
rect 457 -869 458 -867
rect 464 -863 465 -861
rect 464 -869 465 -867
rect 471 -863 472 -861
rect 471 -869 472 -867
rect 478 -863 479 -861
rect 478 -869 479 -867
rect 485 -863 486 -861
rect 485 -869 486 -867
rect 492 -863 493 -861
rect 492 -869 493 -867
rect 499 -863 500 -861
rect 499 -869 500 -867
rect 506 -863 507 -861
rect 506 -869 507 -867
rect 513 -863 514 -861
rect 516 -863 517 -861
rect 513 -869 514 -867
rect 516 -869 517 -867
rect 520 -863 521 -861
rect 520 -869 521 -867
rect 527 -863 528 -861
rect 527 -869 528 -867
rect 534 -863 535 -861
rect 537 -869 538 -867
rect 544 -869 545 -867
rect 548 -863 549 -861
rect 548 -869 549 -867
rect 555 -863 556 -861
rect 555 -869 556 -867
rect 562 -863 563 -861
rect 562 -869 563 -867
rect 2 -918 3 -916
rect 2 -924 3 -922
rect 9 -924 10 -922
rect 16 -918 17 -916
rect 16 -924 17 -922
rect 23 -918 24 -916
rect 23 -924 24 -922
rect 30 -924 31 -922
rect 37 -918 38 -916
rect 44 -918 45 -916
rect 54 -918 55 -916
rect 58 -924 59 -922
rect 65 -918 66 -916
rect 68 -918 69 -916
rect 72 -924 73 -922
rect 79 -918 80 -916
rect 79 -924 80 -922
rect 86 -918 87 -916
rect 86 -924 87 -922
rect 96 -918 97 -916
rect 93 -924 94 -922
rect 96 -924 97 -922
rect 100 -918 101 -916
rect 103 -918 104 -916
rect 100 -924 101 -922
rect 110 -924 111 -922
rect 114 -918 115 -916
rect 114 -924 115 -922
rect 121 -918 122 -916
rect 124 -918 125 -916
rect 124 -924 125 -922
rect 131 -918 132 -916
rect 128 -924 129 -922
rect 135 -918 136 -916
rect 135 -924 136 -922
rect 142 -918 143 -916
rect 142 -924 143 -922
rect 149 -918 150 -916
rect 152 -918 153 -916
rect 152 -924 153 -922
rect 156 -918 157 -916
rect 156 -924 157 -922
rect 163 -918 164 -916
rect 163 -924 164 -922
rect 173 -918 174 -916
rect 170 -924 171 -922
rect 173 -924 174 -922
rect 177 -918 178 -916
rect 177 -924 178 -922
rect 184 -918 185 -916
rect 184 -924 185 -922
rect 187 -924 188 -922
rect 191 -918 192 -916
rect 194 -918 195 -916
rect 194 -924 195 -922
rect 198 -918 199 -916
rect 201 -918 202 -916
rect 198 -924 199 -922
rect 208 -918 209 -916
rect 208 -924 209 -922
rect 212 -918 213 -916
rect 212 -924 213 -922
rect 219 -918 220 -916
rect 219 -924 220 -922
rect 229 -918 230 -916
rect 233 -918 234 -916
rect 233 -924 234 -922
rect 240 -918 241 -916
rect 243 -918 244 -916
rect 240 -924 241 -922
rect 243 -924 244 -922
rect 247 -918 248 -916
rect 247 -924 248 -922
rect 254 -918 255 -916
rect 254 -924 255 -922
rect 261 -918 262 -916
rect 261 -924 262 -922
rect 268 -918 269 -916
rect 268 -924 269 -922
rect 275 -918 276 -916
rect 275 -924 276 -922
rect 282 -918 283 -916
rect 282 -924 283 -922
rect 289 -918 290 -916
rect 292 -918 293 -916
rect 289 -924 290 -922
rect 299 -918 300 -916
rect 306 -918 307 -916
rect 303 -924 304 -922
rect 306 -924 307 -922
rect 313 -918 314 -916
rect 310 -924 311 -922
rect 317 -918 318 -916
rect 317 -924 318 -922
rect 324 -918 325 -916
rect 324 -924 325 -922
rect 331 -918 332 -916
rect 331 -924 332 -922
rect 338 -918 339 -916
rect 338 -924 339 -922
rect 345 -918 346 -916
rect 345 -924 346 -922
rect 352 -918 353 -916
rect 352 -924 353 -922
rect 359 -924 360 -922
rect 362 -924 363 -922
rect 366 -918 367 -916
rect 366 -924 367 -922
rect 373 -918 374 -916
rect 373 -924 374 -922
rect 380 -918 381 -916
rect 380 -924 381 -922
rect 387 -918 388 -916
rect 387 -924 388 -922
rect 394 -918 395 -916
rect 394 -924 395 -922
rect 401 -918 402 -916
rect 401 -924 402 -922
rect 408 -918 409 -916
rect 408 -924 409 -922
rect 415 -918 416 -916
rect 415 -924 416 -922
rect 422 -918 423 -916
rect 422 -924 423 -922
rect 429 -918 430 -916
rect 429 -924 430 -922
rect 436 -918 437 -916
rect 436 -924 437 -922
rect 446 -918 447 -916
rect 450 -918 451 -916
rect 450 -924 451 -922
rect 457 -918 458 -916
rect 457 -924 458 -922
rect 464 -918 465 -916
rect 464 -924 465 -922
rect 471 -918 472 -916
rect 474 -924 475 -922
rect 478 -918 479 -916
rect 478 -924 479 -922
rect 485 -918 486 -916
rect 485 -924 486 -922
rect 492 -918 493 -916
rect 492 -924 493 -922
rect 499 -918 500 -916
rect 499 -924 500 -922
rect 506 -918 507 -916
rect 506 -924 507 -922
rect 513 -918 514 -916
rect 513 -924 514 -922
rect 520 -918 521 -916
rect 520 -924 521 -922
rect 527 -918 528 -916
rect 530 -918 531 -916
rect 530 -924 531 -922
rect 534 -918 535 -916
rect 534 -924 535 -922
rect 541 -918 542 -916
rect 541 -924 542 -922
rect 548 -918 549 -916
rect 548 -924 549 -922
rect 23 -971 24 -969
rect 23 -977 24 -975
rect 30 -971 31 -969
rect 30 -977 31 -975
rect 37 -971 38 -969
rect 37 -977 38 -975
rect 44 -971 45 -969
rect 54 -971 55 -969
rect 58 -971 59 -969
rect 58 -977 59 -975
rect 65 -971 66 -969
rect 68 -971 69 -969
rect 65 -977 66 -975
rect 68 -977 69 -975
rect 72 -971 73 -969
rect 72 -977 73 -975
rect 79 -971 80 -969
rect 79 -977 80 -975
rect 86 -971 87 -969
rect 86 -977 87 -975
rect 93 -971 94 -969
rect 93 -977 94 -975
rect 100 -971 101 -969
rect 100 -977 101 -975
rect 110 -971 111 -969
rect 107 -977 108 -975
rect 110 -977 111 -975
rect 114 -971 115 -969
rect 117 -971 118 -969
rect 117 -977 118 -975
rect 121 -971 122 -969
rect 121 -977 122 -975
rect 128 -977 129 -975
rect 131 -977 132 -975
rect 135 -971 136 -969
rect 135 -977 136 -975
rect 142 -971 143 -969
rect 145 -971 146 -969
rect 142 -977 143 -975
rect 149 -971 150 -969
rect 152 -971 153 -969
rect 156 -971 157 -969
rect 156 -977 157 -975
rect 166 -971 167 -969
rect 170 -971 171 -969
rect 170 -977 171 -975
rect 177 -971 178 -969
rect 177 -977 178 -975
rect 184 -971 185 -969
rect 187 -971 188 -969
rect 184 -977 185 -975
rect 191 -971 192 -969
rect 191 -977 192 -975
rect 198 -971 199 -969
rect 201 -971 202 -969
rect 198 -977 199 -975
rect 201 -977 202 -975
rect 205 -971 206 -969
rect 208 -971 209 -969
rect 208 -977 209 -975
rect 212 -971 213 -969
rect 212 -977 213 -975
rect 219 -971 220 -969
rect 219 -977 220 -975
rect 226 -971 227 -969
rect 229 -977 230 -975
rect 233 -971 234 -969
rect 240 -971 241 -969
rect 240 -977 241 -975
rect 247 -971 248 -969
rect 247 -977 248 -975
rect 254 -971 255 -969
rect 254 -977 255 -975
rect 261 -971 262 -969
rect 264 -971 265 -969
rect 261 -977 262 -975
rect 264 -977 265 -975
rect 268 -971 269 -969
rect 268 -977 269 -975
rect 275 -971 276 -969
rect 275 -977 276 -975
rect 278 -977 279 -975
rect 282 -971 283 -969
rect 285 -971 286 -969
rect 289 -971 290 -969
rect 289 -977 290 -975
rect 296 -971 297 -969
rect 299 -971 300 -969
rect 299 -977 300 -975
rect 303 -971 304 -969
rect 303 -977 304 -975
rect 310 -971 311 -969
rect 310 -977 311 -975
rect 320 -971 321 -969
rect 320 -977 321 -975
rect 324 -971 325 -969
rect 324 -977 325 -975
rect 331 -971 332 -969
rect 331 -977 332 -975
rect 338 -971 339 -969
rect 338 -977 339 -975
rect 345 -971 346 -969
rect 345 -977 346 -975
rect 352 -971 353 -969
rect 352 -977 353 -975
rect 359 -971 360 -969
rect 359 -977 360 -975
rect 366 -971 367 -969
rect 366 -977 367 -975
rect 373 -971 374 -969
rect 373 -977 374 -975
rect 383 -971 384 -969
rect 380 -977 381 -975
rect 387 -971 388 -969
rect 387 -977 388 -975
rect 394 -971 395 -969
rect 394 -977 395 -975
rect 401 -971 402 -969
rect 401 -977 402 -975
rect 411 -971 412 -969
rect 411 -977 412 -975
rect 415 -971 416 -969
rect 415 -977 416 -975
rect 422 -977 423 -975
rect 429 -971 430 -969
rect 429 -977 430 -975
rect 436 -971 437 -969
rect 436 -977 437 -975
rect 443 -971 444 -969
rect 443 -977 444 -975
rect 450 -971 451 -969
rect 450 -977 451 -975
rect 457 -971 458 -969
rect 457 -977 458 -975
rect 464 -971 465 -969
rect 467 -971 468 -969
rect 464 -977 465 -975
rect 471 -971 472 -969
rect 471 -977 472 -975
rect 478 -971 479 -969
rect 481 -971 482 -969
rect 478 -977 479 -975
rect 485 -971 486 -969
rect 485 -977 486 -975
rect 492 -971 493 -969
rect 492 -977 493 -975
rect 499 -971 500 -969
rect 499 -977 500 -975
rect 506 -971 507 -969
rect 509 -971 510 -969
rect 509 -977 510 -975
rect 520 -971 521 -969
rect 520 -977 521 -975
rect 16 -1012 17 -1010
rect 16 -1018 17 -1016
rect 26 -1012 27 -1010
rect 30 -1012 31 -1010
rect 30 -1018 31 -1016
rect 37 -1012 38 -1010
rect 37 -1018 38 -1016
rect 47 -1018 48 -1016
rect 51 -1012 52 -1010
rect 51 -1018 52 -1016
rect 58 -1012 59 -1010
rect 58 -1018 59 -1016
rect 65 -1012 66 -1010
rect 68 -1012 69 -1010
rect 72 -1012 73 -1010
rect 72 -1018 73 -1016
rect 79 -1012 80 -1010
rect 79 -1018 80 -1016
rect 86 -1018 87 -1016
rect 89 -1018 90 -1016
rect 96 -1012 97 -1010
rect 96 -1018 97 -1016
rect 100 -1012 101 -1010
rect 100 -1018 101 -1016
rect 107 -1012 108 -1010
rect 107 -1018 108 -1016
rect 114 -1012 115 -1010
rect 117 -1012 118 -1010
rect 114 -1018 115 -1016
rect 117 -1018 118 -1016
rect 121 -1012 122 -1010
rect 121 -1018 122 -1016
rect 128 -1012 129 -1010
rect 131 -1012 132 -1010
rect 135 -1012 136 -1010
rect 135 -1018 136 -1016
rect 142 -1012 143 -1010
rect 142 -1018 143 -1016
rect 149 -1012 150 -1010
rect 149 -1018 150 -1016
rect 156 -1012 157 -1010
rect 156 -1018 157 -1016
rect 163 -1012 164 -1010
rect 163 -1018 164 -1016
rect 170 -1012 171 -1010
rect 173 -1012 174 -1010
rect 177 -1012 178 -1010
rect 177 -1018 178 -1016
rect 187 -1012 188 -1010
rect 184 -1018 185 -1016
rect 187 -1018 188 -1016
rect 191 -1012 192 -1010
rect 194 -1018 195 -1016
rect 198 -1012 199 -1010
rect 201 -1012 202 -1010
rect 201 -1018 202 -1016
rect 205 -1012 206 -1010
rect 208 -1012 209 -1010
rect 208 -1018 209 -1016
rect 212 -1012 213 -1010
rect 212 -1018 213 -1016
rect 219 -1012 220 -1010
rect 219 -1018 220 -1016
rect 226 -1012 227 -1010
rect 229 -1012 230 -1010
rect 226 -1018 227 -1016
rect 229 -1018 230 -1016
rect 233 -1012 234 -1010
rect 236 -1012 237 -1010
rect 233 -1018 234 -1016
rect 240 -1012 241 -1010
rect 240 -1018 241 -1016
rect 247 -1012 248 -1010
rect 247 -1018 248 -1016
rect 254 -1012 255 -1010
rect 254 -1018 255 -1016
rect 261 -1012 262 -1010
rect 261 -1018 262 -1016
rect 271 -1012 272 -1010
rect 268 -1018 269 -1016
rect 275 -1018 276 -1016
rect 278 -1018 279 -1016
rect 282 -1012 283 -1010
rect 285 -1018 286 -1016
rect 289 -1012 290 -1010
rect 292 -1012 293 -1010
rect 292 -1018 293 -1016
rect 296 -1012 297 -1010
rect 299 -1012 300 -1010
rect 303 -1012 304 -1010
rect 303 -1018 304 -1016
rect 310 -1012 311 -1010
rect 310 -1018 311 -1016
rect 317 -1012 318 -1010
rect 317 -1018 318 -1016
rect 324 -1012 325 -1010
rect 324 -1018 325 -1016
rect 327 -1018 328 -1016
rect 331 -1012 332 -1010
rect 331 -1018 332 -1016
rect 338 -1012 339 -1010
rect 338 -1018 339 -1016
rect 345 -1012 346 -1010
rect 345 -1018 346 -1016
rect 352 -1012 353 -1010
rect 352 -1018 353 -1016
rect 359 -1012 360 -1010
rect 359 -1018 360 -1016
rect 366 -1012 367 -1010
rect 369 -1018 370 -1016
rect 373 -1012 374 -1010
rect 373 -1018 374 -1016
rect 380 -1012 381 -1010
rect 380 -1018 381 -1016
rect 387 -1012 388 -1010
rect 390 -1012 391 -1010
rect 387 -1018 388 -1016
rect 394 -1012 395 -1010
rect 394 -1018 395 -1016
rect 401 -1012 402 -1010
rect 401 -1018 402 -1016
rect 408 -1012 409 -1010
rect 408 -1018 409 -1016
rect 415 -1012 416 -1010
rect 415 -1018 416 -1016
rect 422 -1012 423 -1010
rect 422 -1018 423 -1016
rect 429 -1012 430 -1010
rect 432 -1012 433 -1010
rect 436 -1012 437 -1010
rect 436 -1018 437 -1016
rect 443 -1012 444 -1010
rect 446 -1012 447 -1010
rect 443 -1018 444 -1016
rect 453 -1018 454 -1016
rect 457 -1012 458 -1010
rect 457 -1018 458 -1016
rect 464 -1012 465 -1010
rect 464 -1018 465 -1016
rect 471 -1012 472 -1010
rect 471 -1018 472 -1016
rect 478 -1012 479 -1010
rect 478 -1018 479 -1016
rect 520 -1018 521 -1016
rect 523 -1018 524 -1016
rect 527 -1012 528 -1010
rect 527 -1018 528 -1016
rect 65 -1049 66 -1047
rect 65 -1055 66 -1053
rect 72 -1049 73 -1047
rect 72 -1055 73 -1053
rect 79 -1055 80 -1053
rect 86 -1049 87 -1047
rect 89 -1055 90 -1053
rect 93 -1049 94 -1047
rect 93 -1055 94 -1053
rect 103 -1049 104 -1047
rect 103 -1055 104 -1053
rect 107 -1049 108 -1047
rect 107 -1055 108 -1053
rect 114 -1049 115 -1047
rect 117 -1049 118 -1047
rect 114 -1055 115 -1053
rect 117 -1055 118 -1053
rect 121 -1049 122 -1047
rect 121 -1055 122 -1053
rect 128 -1049 129 -1047
rect 128 -1055 129 -1053
rect 135 -1049 136 -1047
rect 135 -1055 136 -1053
rect 142 -1055 143 -1053
rect 145 -1055 146 -1053
rect 149 -1049 150 -1047
rect 149 -1055 150 -1053
rect 152 -1055 153 -1053
rect 159 -1055 160 -1053
rect 166 -1049 167 -1047
rect 163 -1055 164 -1053
rect 170 -1049 171 -1047
rect 177 -1049 178 -1047
rect 177 -1055 178 -1053
rect 184 -1049 185 -1047
rect 184 -1055 185 -1053
rect 191 -1049 192 -1047
rect 191 -1055 192 -1053
rect 201 -1049 202 -1047
rect 201 -1055 202 -1053
rect 205 -1049 206 -1047
rect 208 -1049 209 -1047
rect 205 -1055 206 -1053
rect 208 -1055 209 -1053
rect 212 -1049 213 -1047
rect 215 -1049 216 -1047
rect 212 -1055 213 -1053
rect 215 -1055 216 -1053
rect 219 -1049 220 -1047
rect 219 -1055 220 -1053
rect 226 -1049 227 -1047
rect 229 -1049 230 -1047
rect 236 -1049 237 -1047
rect 236 -1055 237 -1053
rect 240 -1049 241 -1047
rect 240 -1055 241 -1053
rect 247 -1049 248 -1047
rect 250 -1049 251 -1047
rect 247 -1055 248 -1053
rect 250 -1055 251 -1053
rect 254 -1049 255 -1047
rect 254 -1055 255 -1053
rect 261 -1049 262 -1047
rect 261 -1055 262 -1053
rect 268 -1049 269 -1047
rect 268 -1055 269 -1053
rect 275 -1049 276 -1047
rect 275 -1055 276 -1053
rect 282 -1049 283 -1047
rect 282 -1055 283 -1053
rect 289 -1049 290 -1047
rect 292 -1049 293 -1047
rect 289 -1055 290 -1053
rect 292 -1055 293 -1053
rect 296 -1049 297 -1047
rect 296 -1055 297 -1053
rect 303 -1049 304 -1047
rect 303 -1055 304 -1053
rect 310 -1049 311 -1047
rect 310 -1055 311 -1053
rect 317 -1049 318 -1047
rect 317 -1055 318 -1053
rect 324 -1049 325 -1047
rect 324 -1055 325 -1053
rect 334 -1049 335 -1047
rect 334 -1055 335 -1053
rect 338 -1049 339 -1047
rect 338 -1055 339 -1053
rect 345 -1049 346 -1047
rect 345 -1055 346 -1053
rect 355 -1049 356 -1047
rect 359 -1049 360 -1047
rect 359 -1055 360 -1053
rect 362 -1055 363 -1053
rect 366 -1049 367 -1047
rect 366 -1055 367 -1053
rect 373 -1049 374 -1047
rect 373 -1055 374 -1053
rect 380 -1049 381 -1047
rect 380 -1055 381 -1053
rect 387 -1049 388 -1047
rect 387 -1055 388 -1053
rect 394 -1049 395 -1047
rect 394 -1055 395 -1053
rect 401 -1049 402 -1047
rect 401 -1055 402 -1053
rect 408 -1049 409 -1047
rect 408 -1055 409 -1053
rect 415 -1049 416 -1047
rect 415 -1055 416 -1053
rect 422 -1049 423 -1047
rect 429 -1049 430 -1047
rect 429 -1055 430 -1053
rect 443 -1049 444 -1047
rect 450 -1049 451 -1047
rect 453 -1049 454 -1047
rect 457 -1049 458 -1047
rect 457 -1055 458 -1053
rect 478 -1049 479 -1047
rect 478 -1055 479 -1053
rect 516 -1049 517 -1047
rect 523 -1049 524 -1047
rect 520 -1055 521 -1053
rect 527 -1049 528 -1047
rect 527 -1055 528 -1053
rect 51 -1094 52 -1092
rect 51 -1100 52 -1098
rect 61 -1094 62 -1092
rect 65 -1094 66 -1092
rect 65 -1100 66 -1098
rect 75 -1094 76 -1092
rect 72 -1100 73 -1098
rect 79 -1100 80 -1098
rect 89 -1100 90 -1098
rect 93 -1094 94 -1092
rect 93 -1100 94 -1098
rect 100 -1094 101 -1092
rect 100 -1100 101 -1098
rect 107 -1094 108 -1092
rect 110 -1094 111 -1092
rect 107 -1100 108 -1098
rect 110 -1100 111 -1098
rect 114 -1094 115 -1092
rect 114 -1100 115 -1098
rect 121 -1094 122 -1092
rect 121 -1100 122 -1098
rect 131 -1094 132 -1092
rect 135 -1094 136 -1092
rect 135 -1100 136 -1098
rect 138 -1100 139 -1098
rect 142 -1094 143 -1092
rect 142 -1100 143 -1098
rect 149 -1094 150 -1092
rect 149 -1100 150 -1098
rect 156 -1094 157 -1092
rect 156 -1100 157 -1098
rect 163 -1094 164 -1092
rect 163 -1100 164 -1098
rect 170 -1100 171 -1098
rect 177 -1094 178 -1092
rect 180 -1094 181 -1092
rect 180 -1100 181 -1098
rect 184 -1100 185 -1098
rect 187 -1100 188 -1098
rect 191 -1100 192 -1098
rect 198 -1094 199 -1092
rect 198 -1100 199 -1098
rect 205 -1094 206 -1092
rect 205 -1100 206 -1098
rect 212 -1094 213 -1092
rect 212 -1100 213 -1098
rect 219 -1094 220 -1092
rect 222 -1094 223 -1092
rect 222 -1100 223 -1098
rect 226 -1094 227 -1092
rect 226 -1100 227 -1098
rect 233 -1094 234 -1092
rect 236 -1094 237 -1092
rect 236 -1100 237 -1098
rect 240 -1094 241 -1092
rect 240 -1100 241 -1098
rect 247 -1094 248 -1092
rect 247 -1100 248 -1098
rect 254 -1094 255 -1092
rect 254 -1100 255 -1098
rect 261 -1094 262 -1092
rect 261 -1100 262 -1098
rect 268 -1094 269 -1092
rect 268 -1100 269 -1098
rect 275 -1094 276 -1092
rect 275 -1100 276 -1098
rect 282 -1094 283 -1092
rect 282 -1100 283 -1098
rect 289 -1094 290 -1092
rect 299 -1094 300 -1092
rect 296 -1100 297 -1098
rect 299 -1100 300 -1098
rect 306 -1094 307 -1092
rect 303 -1100 304 -1098
rect 306 -1100 307 -1098
rect 310 -1094 311 -1092
rect 310 -1100 311 -1098
rect 317 -1094 318 -1092
rect 320 -1094 321 -1092
rect 320 -1100 321 -1098
rect 324 -1094 325 -1092
rect 324 -1100 325 -1098
rect 331 -1094 332 -1092
rect 331 -1100 332 -1098
rect 338 -1094 339 -1092
rect 338 -1100 339 -1098
rect 345 -1094 346 -1092
rect 345 -1100 346 -1098
rect 352 -1094 353 -1092
rect 352 -1100 353 -1098
rect 359 -1094 360 -1092
rect 362 -1094 363 -1092
rect 359 -1100 360 -1098
rect 366 -1094 367 -1092
rect 366 -1100 367 -1098
rect 373 -1094 374 -1092
rect 373 -1100 374 -1098
rect 376 -1100 377 -1098
rect 380 -1094 381 -1092
rect 380 -1100 381 -1098
rect 387 -1094 388 -1092
rect 390 -1094 391 -1092
rect 387 -1100 388 -1098
rect 394 -1094 395 -1092
rect 394 -1100 395 -1098
rect 401 -1094 402 -1092
rect 401 -1100 402 -1098
rect 408 -1094 409 -1092
rect 408 -1100 409 -1098
rect 415 -1100 416 -1098
rect 418 -1100 419 -1098
rect 422 -1094 423 -1092
rect 422 -1100 423 -1098
rect 429 -1094 430 -1092
rect 429 -1100 430 -1098
rect 436 -1094 437 -1092
rect 460 -1100 461 -1098
rect 464 -1094 465 -1092
rect 464 -1100 465 -1098
rect 478 -1094 479 -1092
rect 478 -1100 479 -1098
rect 30 -1131 31 -1129
rect 30 -1137 31 -1135
rect 37 -1131 38 -1129
rect 37 -1137 38 -1135
rect 44 -1131 45 -1129
rect 44 -1137 45 -1135
rect 54 -1131 55 -1129
rect 58 -1131 59 -1129
rect 58 -1137 59 -1135
rect 65 -1131 66 -1129
rect 65 -1137 66 -1135
rect 75 -1131 76 -1129
rect 75 -1137 76 -1135
rect 79 -1131 80 -1129
rect 82 -1131 83 -1129
rect 79 -1137 80 -1135
rect 86 -1131 87 -1129
rect 89 -1137 90 -1135
rect 96 -1137 97 -1135
rect 100 -1131 101 -1129
rect 100 -1137 101 -1135
rect 107 -1131 108 -1129
rect 107 -1137 108 -1135
rect 114 -1131 115 -1129
rect 117 -1137 118 -1135
rect 121 -1131 122 -1129
rect 121 -1137 122 -1135
rect 131 -1131 132 -1129
rect 128 -1137 129 -1135
rect 135 -1131 136 -1129
rect 135 -1137 136 -1135
rect 142 -1131 143 -1129
rect 142 -1137 143 -1135
rect 149 -1131 150 -1129
rect 149 -1137 150 -1135
rect 159 -1131 160 -1129
rect 159 -1137 160 -1135
rect 163 -1131 164 -1129
rect 163 -1137 164 -1135
rect 170 -1131 171 -1129
rect 170 -1137 171 -1135
rect 177 -1131 178 -1129
rect 177 -1137 178 -1135
rect 184 -1131 185 -1129
rect 184 -1137 185 -1135
rect 191 -1131 192 -1129
rect 194 -1131 195 -1129
rect 191 -1137 192 -1135
rect 198 -1137 199 -1135
rect 201 -1137 202 -1135
rect 205 -1131 206 -1129
rect 208 -1131 209 -1129
rect 205 -1137 206 -1135
rect 208 -1137 209 -1135
rect 212 -1131 213 -1129
rect 212 -1137 213 -1135
rect 219 -1131 220 -1129
rect 219 -1137 220 -1135
rect 226 -1131 227 -1129
rect 226 -1137 227 -1135
rect 229 -1137 230 -1135
rect 233 -1131 234 -1129
rect 233 -1137 234 -1135
rect 240 -1131 241 -1129
rect 240 -1137 241 -1135
rect 247 -1131 248 -1129
rect 247 -1137 248 -1135
rect 254 -1131 255 -1129
rect 254 -1137 255 -1135
rect 261 -1131 262 -1129
rect 264 -1131 265 -1129
rect 261 -1137 262 -1135
rect 264 -1137 265 -1135
rect 268 -1131 269 -1129
rect 268 -1137 269 -1135
rect 275 -1131 276 -1129
rect 278 -1131 279 -1129
rect 275 -1137 276 -1135
rect 278 -1137 279 -1135
rect 282 -1131 283 -1129
rect 282 -1137 283 -1135
rect 289 -1131 290 -1129
rect 289 -1137 290 -1135
rect 296 -1131 297 -1129
rect 296 -1137 297 -1135
rect 303 -1137 304 -1135
rect 306 -1137 307 -1135
rect 310 -1131 311 -1129
rect 310 -1137 311 -1135
rect 317 -1131 318 -1129
rect 320 -1131 321 -1129
rect 327 -1137 328 -1135
rect 331 -1131 332 -1129
rect 331 -1137 332 -1135
rect 338 -1131 339 -1129
rect 338 -1137 339 -1135
rect 345 -1131 346 -1129
rect 345 -1137 346 -1135
rect 352 -1131 353 -1129
rect 352 -1137 353 -1135
rect 359 -1131 360 -1129
rect 362 -1131 363 -1129
rect 369 -1131 370 -1129
rect 369 -1137 370 -1135
rect 373 -1131 374 -1129
rect 373 -1137 374 -1135
rect 380 -1131 381 -1129
rect 380 -1137 381 -1135
rect 387 -1131 388 -1129
rect 387 -1137 388 -1135
rect 394 -1131 395 -1129
rect 394 -1137 395 -1135
rect 401 -1131 402 -1129
rect 401 -1137 402 -1135
rect 408 -1131 409 -1129
rect 408 -1137 409 -1135
rect 415 -1131 416 -1129
rect 415 -1137 416 -1135
rect 422 -1131 423 -1129
rect 422 -1137 423 -1135
rect 429 -1131 430 -1129
rect 429 -1137 430 -1135
rect 436 -1131 437 -1129
rect 436 -1137 437 -1135
rect 443 -1131 444 -1129
rect 443 -1137 444 -1135
rect 478 -1131 479 -1129
rect 478 -1137 479 -1135
rect 485 -1137 486 -1135
rect 54 -1174 55 -1172
rect 61 -1180 62 -1178
rect 72 -1174 73 -1172
rect 72 -1180 73 -1178
rect 82 -1174 83 -1172
rect 86 -1174 87 -1172
rect 86 -1180 87 -1178
rect 93 -1174 94 -1172
rect 100 -1174 101 -1172
rect 100 -1180 101 -1178
rect 107 -1174 108 -1172
rect 107 -1180 108 -1178
rect 114 -1174 115 -1172
rect 117 -1174 118 -1172
rect 114 -1180 115 -1178
rect 121 -1174 122 -1172
rect 124 -1174 125 -1172
rect 121 -1180 122 -1178
rect 124 -1180 125 -1178
rect 128 -1174 129 -1172
rect 128 -1180 129 -1178
rect 135 -1174 136 -1172
rect 135 -1180 136 -1178
rect 145 -1174 146 -1172
rect 149 -1174 150 -1172
rect 149 -1180 150 -1178
rect 156 -1174 157 -1172
rect 156 -1180 157 -1178
rect 163 -1174 164 -1172
rect 166 -1174 167 -1172
rect 170 -1174 171 -1172
rect 173 -1174 174 -1172
rect 170 -1180 171 -1178
rect 177 -1174 178 -1172
rect 177 -1180 178 -1178
rect 184 -1174 185 -1172
rect 184 -1180 185 -1178
rect 191 -1174 192 -1172
rect 191 -1180 192 -1178
rect 198 -1174 199 -1172
rect 198 -1180 199 -1178
rect 201 -1180 202 -1178
rect 205 -1174 206 -1172
rect 208 -1174 209 -1172
rect 205 -1180 206 -1178
rect 208 -1180 209 -1178
rect 212 -1174 213 -1172
rect 212 -1180 213 -1178
rect 219 -1174 220 -1172
rect 219 -1180 220 -1178
rect 226 -1174 227 -1172
rect 226 -1180 227 -1178
rect 233 -1174 234 -1172
rect 233 -1180 234 -1178
rect 240 -1174 241 -1172
rect 243 -1174 244 -1172
rect 240 -1180 241 -1178
rect 250 -1174 251 -1172
rect 247 -1180 248 -1178
rect 250 -1180 251 -1178
rect 254 -1174 255 -1172
rect 257 -1180 258 -1178
rect 261 -1174 262 -1172
rect 264 -1174 265 -1172
rect 261 -1180 262 -1178
rect 268 -1174 269 -1172
rect 268 -1180 269 -1178
rect 275 -1174 276 -1172
rect 275 -1180 276 -1178
rect 282 -1174 283 -1172
rect 282 -1180 283 -1178
rect 289 -1174 290 -1172
rect 289 -1180 290 -1178
rect 299 -1174 300 -1172
rect 296 -1180 297 -1178
rect 306 -1174 307 -1172
rect 303 -1180 304 -1178
rect 310 -1174 311 -1172
rect 310 -1180 311 -1178
rect 317 -1174 318 -1172
rect 317 -1180 318 -1178
rect 324 -1174 325 -1172
rect 324 -1180 325 -1178
rect 331 -1174 332 -1172
rect 331 -1180 332 -1178
rect 338 -1174 339 -1172
rect 338 -1180 339 -1178
rect 345 -1174 346 -1172
rect 345 -1180 346 -1178
rect 352 -1174 353 -1172
rect 352 -1180 353 -1178
rect 359 -1174 360 -1172
rect 359 -1180 360 -1178
rect 366 -1174 367 -1172
rect 366 -1180 367 -1178
rect 376 -1174 377 -1172
rect 376 -1180 377 -1178
rect 380 -1174 381 -1172
rect 380 -1180 381 -1178
rect 387 -1174 388 -1172
rect 387 -1180 388 -1178
rect 397 -1174 398 -1172
rect 401 -1174 402 -1172
rect 401 -1180 402 -1178
rect 408 -1174 409 -1172
rect 65 -1205 66 -1203
rect 65 -1211 66 -1209
rect 72 -1205 73 -1203
rect 72 -1211 73 -1209
rect 79 -1205 80 -1203
rect 79 -1211 80 -1209
rect 89 -1211 90 -1209
rect 93 -1205 94 -1203
rect 93 -1211 94 -1209
rect 100 -1205 101 -1203
rect 100 -1211 101 -1209
rect 107 -1205 108 -1203
rect 107 -1211 108 -1209
rect 114 -1205 115 -1203
rect 114 -1211 115 -1209
rect 121 -1205 122 -1203
rect 121 -1211 122 -1209
rect 131 -1205 132 -1203
rect 128 -1211 129 -1209
rect 138 -1205 139 -1203
rect 138 -1211 139 -1209
rect 142 -1205 143 -1203
rect 142 -1211 143 -1209
rect 149 -1211 150 -1209
rect 156 -1205 157 -1203
rect 159 -1211 160 -1209
rect 163 -1205 164 -1203
rect 163 -1211 164 -1209
rect 170 -1205 171 -1203
rect 173 -1205 174 -1203
rect 177 -1211 178 -1209
rect 180 -1211 181 -1209
rect 184 -1205 185 -1203
rect 187 -1211 188 -1209
rect 191 -1205 192 -1203
rect 194 -1205 195 -1203
rect 191 -1211 192 -1209
rect 198 -1205 199 -1203
rect 198 -1211 199 -1209
rect 208 -1205 209 -1203
rect 212 -1205 213 -1203
rect 212 -1211 213 -1209
rect 219 -1205 220 -1203
rect 219 -1211 220 -1209
rect 229 -1211 230 -1209
rect 233 -1205 234 -1203
rect 233 -1211 234 -1209
rect 240 -1205 241 -1203
rect 240 -1211 241 -1209
rect 243 -1211 244 -1209
rect 247 -1205 248 -1203
rect 247 -1211 248 -1209
rect 254 -1205 255 -1203
rect 254 -1211 255 -1209
rect 261 -1211 262 -1209
rect 264 -1211 265 -1209
rect 268 -1205 269 -1203
rect 268 -1211 269 -1209
rect 275 -1205 276 -1203
rect 275 -1211 276 -1209
rect 282 -1205 283 -1203
rect 282 -1211 283 -1209
rect 292 -1205 293 -1203
rect 292 -1211 293 -1209
rect 296 -1205 297 -1203
rect 296 -1211 297 -1209
rect 303 -1211 304 -1209
rect 310 -1205 311 -1203
rect 310 -1211 311 -1209
rect 317 -1211 318 -1209
rect 324 -1205 325 -1203
rect 331 -1205 332 -1203
rect 331 -1211 332 -1209
rect 338 -1205 339 -1203
rect 338 -1211 339 -1209
rect 345 -1205 346 -1203
rect 345 -1211 346 -1209
rect 352 -1205 353 -1203
rect 352 -1211 353 -1209
rect 359 -1205 360 -1203
rect 359 -1211 360 -1209
rect 366 -1205 367 -1203
rect 366 -1211 367 -1209
rect 373 -1205 374 -1203
rect 373 -1211 374 -1209
rect 380 -1205 381 -1203
rect 383 -1205 384 -1203
rect 383 -1211 384 -1209
rect 387 -1205 388 -1203
rect 387 -1211 388 -1209
rect 394 -1205 395 -1203
rect 394 -1211 395 -1209
rect 93 -1234 94 -1232
rect 93 -1240 94 -1238
rect 100 -1240 101 -1238
rect 110 -1240 111 -1238
rect 114 -1234 115 -1232
rect 114 -1240 115 -1238
rect 121 -1234 122 -1232
rect 128 -1234 129 -1232
rect 128 -1240 129 -1238
rect 135 -1234 136 -1232
rect 135 -1240 136 -1238
rect 142 -1234 143 -1232
rect 142 -1240 143 -1238
rect 152 -1234 153 -1232
rect 152 -1240 153 -1238
rect 156 -1234 157 -1232
rect 156 -1240 157 -1238
rect 163 -1234 164 -1232
rect 163 -1240 164 -1238
rect 170 -1234 171 -1232
rect 180 -1234 181 -1232
rect 180 -1240 181 -1238
rect 184 -1234 185 -1232
rect 187 -1240 188 -1238
rect 194 -1234 195 -1232
rect 191 -1240 192 -1238
rect 201 -1240 202 -1238
rect 205 -1234 206 -1232
rect 205 -1240 206 -1238
rect 212 -1234 213 -1232
rect 212 -1240 213 -1238
rect 219 -1240 220 -1238
rect 226 -1234 227 -1232
rect 226 -1240 227 -1238
rect 233 -1234 234 -1232
rect 233 -1240 234 -1238
rect 240 -1234 241 -1232
rect 240 -1240 241 -1238
rect 247 -1234 248 -1232
rect 247 -1240 248 -1238
rect 254 -1234 255 -1232
rect 261 -1234 262 -1232
rect 261 -1240 262 -1238
rect 268 -1234 269 -1232
rect 275 -1234 276 -1232
rect 275 -1240 276 -1238
rect 282 -1234 283 -1232
rect 282 -1240 283 -1238
rect 289 -1234 290 -1232
rect 289 -1240 290 -1238
rect 296 -1234 297 -1232
rect 299 -1240 300 -1238
rect 306 -1240 307 -1238
rect 310 -1234 311 -1232
rect 310 -1240 311 -1238
rect 317 -1234 318 -1232
rect 317 -1240 318 -1238
rect 324 -1234 325 -1232
rect 324 -1240 325 -1238
rect 331 -1234 332 -1232
rect 331 -1240 332 -1238
rect 348 -1240 349 -1238
rect 352 -1234 353 -1232
rect 352 -1240 353 -1238
rect 380 -1234 381 -1232
rect 380 -1240 381 -1238
rect 5 -1261 6 -1259
rect 75 -1261 76 -1259
rect 82 -1255 83 -1253
rect 79 -1261 80 -1259
rect 86 -1255 87 -1253
rect 86 -1261 87 -1259
rect 100 -1255 101 -1253
rect 100 -1261 101 -1259
rect 107 -1255 108 -1253
rect 107 -1261 108 -1259
rect 117 -1255 118 -1253
rect 114 -1261 115 -1259
rect 121 -1255 122 -1253
rect 121 -1261 122 -1259
rect 128 -1255 129 -1253
rect 128 -1261 129 -1259
rect 135 -1255 136 -1253
rect 135 -1261 136 -1259
rect 145 -1261 146 -1259
rect 149 -1255 150 -1253
rect 149 -1261 150 -1259
rect 156 -1255 157 -1253
rect 163 -1261 164 -1259
rect 166 -1261 167 -1259
rect 173 -1255 174 -1253
rect 173 -1261 174 -1259
rect 177 -1255 178 -1253
rect 177 -1261 178 -1259
rect 184 -1261 185 -1259
rect 191 -1255 192 -1253
rect 191 -1261 192 -1259
rect 198 -1255 199 -1253
rect 205 -1255 206 -1253
rect 205 -1261 206 -1259
rect 215 -1255 216 -1253
rect 219 -1255 220 -1253
rect 219 -1261 220 -1259
rect 226 -1255 227 -1253
rect 233 -1255 234 -1253
rect 233 -1261 234 -1259
rect 240 -1255 241 -1253
rect 240 -1261 241 -1259
rect 247 -1255 248 -1253
rect 254 -1255 255 -1253
rect 254 -1261 255 -1259
rect 261 -1255 262 -1253
rect 261 -1261 262 -1259
rect 268 -1255 269 -1253
rect 268 -1261 269 -1259
rect 278 -1255 279 -1253
rect 275 -1261 276 -1259
rect 278 -1261 279 -1259
rect 285 -1255 286 -1253
rect 289 -1255 290 -1253
rect 296 -1255 297 -1253
rect 296 -1261 297 -1259
rect 303 -1255 304 -1253
rect 303 -1261 304 -1259
rect 320 -1255 321 -1253
rect 320 -1261 321 -1259
rect 324 -1255 325 -1253
rect 324 -1261 325 -1259
rect 380 -1255 381 -1253
rect 380 -1261 381 -1259
rect 5 -1270 6 -1268
rect 86 -1270 87 -1268
rect 86 -1276 87 -1274
rect 96 -1276 97 -1274
rect 107 -1270 108 -1268
rect 107 -1276 108 -1274
rect 117 -1270 118 -1268
rect 117 -1276 118 -1274
rect 121 -1270 122 -1268
rect 121 -1276 122 -1274
rect 128 -1276 129 -1274
rect 135 -1270 136 -1268
rect 135 -1276 136 -1274
rect 145 -1276 146 -1274
rect 149 -1270 150 -1268
rect 149 -1276 150 -1274
rect 156 -1276 157 -1274
rect 159 -1276 160 -1274
rect 166 -1276 167 -1274
rect 170 -1270 171 -1268
rect 184 -1270 185 -1268
rect 205 -1270 206 -1268
rect 215 -1270 216 -1268
rect 219 -1276 220 -1274
rect 226 -1270 227 -1268
rect 226 -1276 227 -1274
rect 233 -1270 234 -1268
rect 240 -1270 241 -1268
rect 271 -1270 272 -1268
rect 275 -1270 276 -1268
rect 275 -1276 276 -1274
rect 282 -1276 283 -1274
rect 299 -1276 300 -1274
rect 303 -1270 304 -1268
rect 303 -1276 304 -1274
rect 383 -1276 384 -1274
rect 387 -1270 388 -1268
rect 387 -1276 388 -1274
<< metal1 >>
rect 135 0 143 1
rect 145 0 157 1
rect 184 0 195 1
rect 212 0 220 1
rect 135 -11 150 -10
rect 156 -11 181 -10
rect 191 -11 199 -10
rect 208 -11 213 -10
rect 257 -11 262 -10
rect 149 -13 153 -12
rect 177 -13 185 -12
rect 212 -13 223 -12
rect 184 -15 206 -14
rect 149 -26 167 -25
rect 170 -26 185 -25
rect 187 -26 192 -25
rect 198 -26 220 -25
rect 229 -26 262 -25
rect 268 -26 272 -25
rect 341 -26 346 -25
rect 145 -28 150 -27
rect 156 -28 174 -27
rect 177 -28 209 -27
rect 243 -28 248 -27
rect 201 -30 213 -29
rect 205 -32 241 -31
rect 212 -34 234 -33
rect 51 -45 55 -44
rect 72 -45 97 -44
rect 138 -45 150 -44
rect 156 -45 199 -44
rect 201 -45 220 -44
rect 236 -45 248 -44
rect 282 -45 290 -44
rect 345 -45 353 -44
rect 359 -45 367 -44
rect 142 -47 199 -46
rect 208 -47 213 -46
rect 240 -47 244 -46
rect 247 -47 262 -46
rect 345 -47 363 -46
rect 163 -49 188 -48
rect 191 -49 206 -48
rect 240 -49 297 -48
rect 170 -51 276 -50
rect 177 -53 192 -52
rect 194 -53 220 -52
rect 261 -53 269 -52
rect 163 -55 178 -54
rect 187 -55 213 -54
rect 254 -55 269 -54
rect 226 -57 255 -56
rect 51 -68 73 -67
rect 79 -68 143 -67
rect 149 -68 188 -67
rect 194 -68 213 -67
rect 219 -68 276 -67
rect 282 -68 377 -67
rect 58 -70 146 -69
rect 149 -70 244 -69
rect 247 -70 304 -69
rect 310 -70 318 -69
rect 320 -70 332 -69
rect 338 -70 349 -69
rect 65 -72 171 -71
rect 198 -72 283 -71
rect 289 -72 311 -71
rect 345 -72 353 -71
rect 72 -74 87 -73
rect 93 -74 139 -73
rect 156 -74 188 -73
rect 201 -74 255 -73
rect 257 -74 325 -73
rect 93 -76 227 -75
rect 229 -76 318 -75
rect 96 -78 101 -77
rect 103 -78 115 -77
rect 121 -78 251 -77
rect 254 -78 269 -77
rect 278 -78 353 -77
rect 107 -80 136 -79
rect 205 -80 220 -79
rect 226 -80 290 -79
rect 296 -80 339 -79
rect 128 -82 192 -81
rect 205 -82 269 -81
rect 212 -84 237 -83
rect 261 -84 297 -83
rect 208 -86 262 -85
rect 233 -88 241 -87
rect 58 -99 171 -98
rect 173 -99 262 -98
rect 352 -99 381 -98
rect 65 -101 181 -100
rect 184 -101 213 -100
rect 236 -101 283 -100
rect 366 -101 374 -100
rect 376 -101 402 -100
rect 72 -103 104 -102
rect 107 -103 202 -102
rect 205 -103 220 -102
rect 243 -103 339 -102
rect 100 -105 115 -104
rect 135 -105 181 -104
rect 187 -105 304 -104
rect 324 -105 367 -104
rect 107 -107 122 -106
rect 145 -107 195 -106
rect 198 -107 272 -106
rect 338 -107 395 -106
rect 86 -109 122 -108
rect 142 -109 146 -108
rect 149 -109 227 -108
rect 236 -109 325 -108
rect 79 -111 143 -110
rect 149 -111 157 -110
rect 163 -111 213 -110
rect 247 -111 297 -110
rect 93 -113 157 -112
rect 163 -113 241 -112
rect 250 -113 297 -112
rect 93 -115 129 -114
rect 177 -115 227 -114
rect 254 -115 318 -114
rect 128 -117 171 -116
rect 191 -117 311 -116
rect 317 -117 332 -116
rect 191 -119 276 -118
rect 310 -119 332 -118
rect 194 -121 241 -120
rect 254 -121 265 -120
rect 205 -123 276 -122
rect 208 -125 262 -124
rect 208 -127 269 -126
rect 219 -129 251 -128
rect 257 -129 290 -128
rect 289 -131 304 -130
rect 65 -142 185 -141
rect 191 -142 342 -141
rect 380 -142 409 -141
rect 93 -144 125 -143
rect 142 -144 157 -143
rect 170 -144 241 -143
rect 243 -144 416 -143
rect 93 -146 118 -145
rect 121 -146 150 -145
rect 163 -146 171 -145
rect 184 -146 237 -145
rect 264 -146 353 -145
rect 380 -146 388 -145
rect 401 -146 430 -145
rect 72 -148 150 -147
rect 152 -148 164 -147
rect 205 -148 213 -147
rect 226 -148 262 -147
rect 289 -148 423 -147
rect 86 -150 118 -149
rect 177 -150 213 -149
rect 233 -150 255 -149
rect 289 -150 297 -149
rect 310 -150 318 -149
rect 331 -150 360 -149
rect 394 -150 402 -149
rect 86 -152 129 -151
rect 229 -152 255 -151
rect 285 -152 297 -151
rect 317 -152 374 -151
rect 107 -154 174 -153
rect 331 -154 356 -153
rect 366 -154 395 -153
rect 107 -156 136 -155
rect 142 -156 230 -155
rect 324 -156 367 -155
rect 100 -158 136 -157
rect 219 -158 325 -157
rect 341 -158 346 -157
rect 100 -160 199 -159
rect 303 -160 346 -159
rect 128 -162 206 -161
rect 247 -162 304 -161
rect 198 -164 269 -163
rect 247 -166 283 -165
rect 23 -177 69 -176
rect 72 -177 202 -176
rect 205 -177 209 -176
rect 219 -177 304 -176
rect 313 -177 353 -176
rect 387 -177 409 -176
rect 411 -177 437 -176
rect 37 -179 244 -178
rect 285 -179 332 -178
rect 341 -179 458 -178
rect 44 -181 80 -180
rect 82 -181 132 -180
rect 149 -181 157 -180
rect 170 -181 181 -180
rect 191 -181 220 -180
rect 236 -181 272 -180
rect 296 -181 311 -180
rect 317 -181 465 -180
rect 51 -183 108 -182
rect 128 -183 195 -182
rect 198 -183 234 -182
rect 240 -183 290 -182
rect 303 -183 325 -182
rect 352 -183 367 -182
rect 380 -183 388 -182
rect 394 -183 430 -182
rect 65 -185 227 -184
rect 243 -185 381 -184
rect 401 -185 440 -184
rect 72 -187 80 -186
rect 86 -187 153 -186
rect 156 -187 223 -186
rect 247 -187 332 -186
rect 359 -187 402 -186
rect 415 -187 444 -186
rect 65 -189 87 -188
rect 93 -189 143 -188
rect 177 -189 216 -188
rect 268 -189 342 -188
rect 373 -189 395 -188
rect 415 -189 433 -188
rect 100 -191 234 -190
rect 275 -191 318 -190
rect 320 -191 367 -190
rect 422 -191 451 -190
rect 96 -193 101 -192
rect 107 -193 164 -192
rect 191 -193 248 -192
rect 268 -193 423 -192
rect 121 -195 143 -194
rect 159 -195 276 -194
rect 285 -195 290 -194
rect 324 -195 360 -194
rect 121 -197 136 -196
rect 138 -197 171 -196
rect 198 -197 213 -196
rect 135 -199 146 -198
rect 163 -199 297 -198
rect 30 -201 146 -200
rect 205 -201 346 -200
rect 254 -203 346 -202
rect 208 -205 255 -204
rect 23 -216 73 -215
rect 100 -216 111 -215
rect 152 -216 451 -215
rect 457 -216 500 -215
rect 541 -216 545 -215
rect 30 -218 206 -217
rect 215 -218 349 -217
rect 408 -218 479 -217
rect 485 -218 538 -217
rect 37 -220 125 -219
rect 156 -220 178 -219
rect 184 -220 213 -219
rect 226 -220 269 -219
rect 271 -220 402 -219
rect 436 -220 472 -219
rect 37 -222 146 -221
rect 149 -222 185 -221
rect 191 -222 304 -221
rect 317 -222 342 -221
rect 345 -222 507 -221
rect 44 -224 59 -223
rect 65 -224 80 -223
rect 100 -224 115 -223
rect 142 -224 178 -223
rect 229 -224 388 -223
rect 429 -224 437 -223
rect 450 -224 535 -223
rect 44 -226 94 -225
rect 107 -226 244 -225
rect 261 -226 297 -225
rect 299 -226 367 -225
rect 464 -226 514 -225
rect 51 -228 139 -227
rect 159 -228 234 -227
rect 236 -228 269 -227
rect 275 -228 325 -227
rect 327 -228 409 -227
rect 443 -228 465 -227
rect 58 -230 227 -229
rect 240 -230 255 -229
rect 275 -230 332 -229
rect 338 -230 521 -229
rect 65 -232 129 -231
rect 163 -232 202 -231
rect 205 -232 262 -231
rect 285 -232 374 -231
rect 51 -234 202 -233
rect 219 -234 255 -233
rect 306 -234 388 -233
rect 79 -236 136 -235
rect 142 -236 220 -235
rect 310 -236 318 -235
rect 331 -236 493 -235
rect 86 -238 164 -237
rect 166 -238 192 -237
rect 198 -238 241 -237
rect 289 -238 311 -237
rect 338 -238 458 -237
rect 93 -240 122 -239
rect 135 -240 181 -239
rect 352 -240 402 -239
rect 89 -242 122 -241
rect 170 -242 209 -241
rect 355 -242 430 -241
rect 170 -244 290 -243
rect 366 -244 395 -243
rect 208 -246 360 -245
rect 394 -246 416 -245
rect 243 -248 360 -247
rect 282 -250 416 -249
rect 282 -252 444 -251
rect 37 -263 230 -262
rect 240 -263 269 -262
rect 282 -263 402 -262
rect 443 -263 556 -262
rect 562 -263 577 -262
rect 37 -265 108 -264
rect 142 -265 213 -264
rect 285 -265 297 -264
rect 303 -265 318 -264
rect 320 -265 507 -264
rect 527 -265 535 -264
rect 44 -267 118 -266
rect 152 -267 234 -266
rect 296 -267 423 -266
rect 464 -267 507 -266
rect 65 -269 132 -268
rect 163 -269 220 -268
rect 306 -269 521 -268
rect 65 -271 115 -270
rect 145 -271 220 -270
rect 324 -271 381 -270
rect 383 -271 549 -270
rect 75 -273 150 -272
rect 170 -273 192 -272
rect 198 -273 290 -272
rect 331 -273 367 -272
rect 408 -273 528 -272
rect 86 -275 129 -274
rect 149 -275 227 -274
rect 289 -275 388 -274
rect 408 -275 416 -274
rect 422 -275 430 -274
rect 499 -275 535 -274
rect 86 -277 115 -276
rect 173 -277 213 -276
rect 226 -277 262 -276
rect 334 -277 479 -276
rect 520 -277 542 -276
rect 79 -279 262 -278
rect 338 -279 388 -278
rect 394 -279 500 -278
rect 93 -281 129 -280
rect 191 -281 269 -280
rect 345 -281 514 -280
rect 96 -283 118 -282
rect 208 -283 276 -282
rect 317 -283 514 -282
rect 100 -285 122 -284
rect 275 -285 360 -284
rect 362 -285 367 -284
rect 415 -285 451 -284
rect 471 -285 479 -284
rect 51 -287 101 -286
rect 107 -287 136 -286
rect 243 -287 451 -286
rect 457 -287 472 -286
rect 51 -289 73 -288
rect 135 -289 167 -288
rect 205 -289 458 -288
rect 72 -291 178 -290
rect 184 -291 206 -290
rect 348 -291 395 -290
rect 429 -291 437 -290
rect 443 -291 542 -290
rect 58 -293 185 -292
rect 303 -293 437 -292
rect 177 -295 248 -294
rect 352 -295 402 -294
rect 247 -297 255 -296
rect 334 -297 353 -296
rect 79 -299 255 -298
rect 9 -310 87 -309
rect 93 -310 150 -309
rect 177 -310 304 -309
rect 334 -310 346 -309
rect 366 -310 479 -309
rect 520 -310 545 -309
rect 548 -310 563 -309
rect 16 -312 276 -311
rect 285 -312 311 -311
rect 334 -312 577 -311
rect 23 -314 97 -313
rect 100 -314 314 -313
rect 338 -314 458 -313
rect 464 -314 493 -313
rect 527 -314 549 -313
rect 30 -316 45 -315
rect 51 -316 62 -315
rect 65 -316 248 -315
rect 250 -316 458 -315
rect 471 -316 556 -315
rect 37 -318 209 -317
rect 240 -318 269 -317
rect 285 -318 577 -317
rect 44 -320 234 -319
rect 240 -320 423 -319
rect 429 -320 528 -319
rect 51 -322 136 -321
rect 180 -322 276 -321
rect 296 -322 430 -321
rect 450 -322 570 -321
rect 61 -324 139 -323
rect 184 -324 248 -323
rect 254 -324 356 -323
rect 373 -324 423 -323
rect 471 -324 514 -323
rect 65 -326 73 -325
rect 79 -326 199 -325
rect 226 -326 255 -325
rect 268 -326 325 -325
rect 348 -326 521 -325
rect 72 -328 143 -327
rect 184 -328 206 -327
rect 219 -328 227 -327
rect 282 -328 570 -327
rect 86 -330 171 -329
rect 194 -330 213 -329
rect 219 -330 262 -329
rect 299 -330 514 -329
rect 103 -332 234 -331
rect 261 -332 297 -331
rect 310 -332 451 -331
rect 107 -334 132 -333
rect 142 -334 339 -333
rect 348 -334 542 -333
rect 114 -336 409 -335
rect 534 -336 542 -335
rect 114 -338 122 -337
rect 149 -338 171 -337
rect 194 -338 304 -337
rect 317 -338 493 -337
rect 121 -340 192 -339
rect 198 -340 283 -339
rect 317 -340 332 -339
rect 345 -340 535 -339
rect 163 -342 213 -341
rect 352 -342 409 -341
rect 156 -344 164 -343
rect 352 -344 479 -343
rect 156 -346 360 -345
rect 373 -346 402 -345
rect 380 -348 507 -347
rect 383 -350 500 -349
rect 387 -352 465 -351
rect 341 -354 388 -353
rect 394 -354 507 -353
rect 271 -356 395 -355
rect 401 -356 416 -355
rect 443 -356 500 -355
rect 292 -358 416 -357
rect 436 -358 444 -357
rect 205 -360 437 -359
rect 2 -371 192 -370
rect 201 -371 332 -370
rect 345 -371 423 -370
rect 513 -371 584 -370
rect 9 -373 136 -372
rect 156 -373 164 -372
rect 184 -373 339 -372
rect 348 -373 395 -372
rect 422 -373 479 -372
rect 534 -373 612 -372
rect 16 -375 251 -374
rect 254 -375 286 -374
rect 296 -375 500 -374
rect 555 -375 577 -374
rect 23 -377 150 -376
rect 156 -377 307 -376
rect 313 -377 472 -376
rect 23 -379 34 -378
rect 37 -379 62 -378
rect 65 -379 178 -378
rect 219 -379 328 -378
rect 352 -379 524 -378
rect 30 -381 59 -380
rect 68 -381 178 -380
rect 226 -381 283 -380
rect 296 -381 318 -380
rect 355 -381 549 -380
rect 37 -383 125 -382
rect 149 -383 164 -382
rect 170 -383 185 -382
rect 299 -383 409 -382
rect 443 -383 500 -382
rect 44 -385 272 -384
rect 303 -385 311 -384
rect 366 -385 465 -384
rect 471 -385 521 -384
rect 44 -387 108 -386
rect 121 -387 262 -386
rect 268 -387 367 -386
rect 380 -387 549 -386
rect 51 -389 220 -388
rect 233 -389 262 -388
rect 320 -389 465 -388
rect 51 -391 104 -390
rect 107 -391 115 -390
rect 170 -391 213 -390
rect 233 -391 276 -390
rect 380 -391 528 -390
rect 58 -393 206 -392
rect 212 -393 328 -392
rect 390 -393 577 -392
rect 72 -395 153 -394
rect 191 -395 276 -394
rect 394 -395 402 -394
rect 408 -395 416 -394
rect 443 -395 493 -394
rect 527 -395 570 -394
rect 72 -397 97 -396
rect 100 -397 227 -396
rect 373 -397 402 -396
rect 415 -397 507 -396
rect 558 -397 570 -396
rect 79 -399 209 -398
rect 348 -399 374 -398
rect 387 -399 493 -398
rect 79 -401 143 -400
rect 152 -401 430 -400
rect 450 -401 535 -400
rect 86 -403 244 -402
rect 383 -403 451 -402
rect 457 -403 479 -402
rect 93 -405 132 -404
rect 138 -405 388 -404
rect 411 -405 507 -404
rect 9 -407 139 -406
rect 142 -407 199 -406
rect 243 -407 248 -406
rect 429 -407 542 -406
rect 114 -409 129 -408
rect 247 -409 514 -408
rect 541 -409 563 -408
rect 359 -411 563 -410
rect 436 -413 458 -412
rect 324 -415 437 -414
rect 2 -426 157 -425
rect 198 -426 220 -425
rect 240 -426 521 -425
rect 576 -426 598 -425
rect 611 -426 640 -425
rect 663 -426 675 -425
rect 2 -428 52 -427
rect 79 -428 188 -427
rect 208 -428 353 -427
rect 355 -428 395 -427
rect 464 -428 626 -427
rect 635 -428 668 -427
rect 9 -430 73 -429
rect 79 -430 178 -429
rect 257 -430 339 -429
rect 348 -430 472 -429
rect 506 -430 591 -429
rect 16 -432 115 -431
rect 128 -432 160 -431
rect 170 -432 220 -431
rect 271 -432 283 -431
rect 310 -432 384 -431
rect 422 -432 507 -431
rect 513 -432 577 -431
rect 583 -432 605 -431
rect 19 -434 248 -433
rect 275 -434 290 -433
rect 313 -434 416 -433
rect 436 -434 584 -433
rect 30 -436 41 -435
rect 44 -436 206 -435
rect 226 -436 416 -435
rect 492 -436 514 -435
rect 527 -436 612 -435
rect 44 -438 622 -437
rect 47 -440 213 -439
rect 233 -440 290 -439
rect 317 -440 549 -439
rect 51 -442 360 -441
rect 362 -442 556 -441
rect 68 -444 339 -443
rect 373 -444 388 -443
rect 401 -444 437 -443
rect 457 -444 549 -443
rect 72 -446 262 -445
rect 275 -446 398 -445
rect 478 -446 556 -445
rect 86 -448 174 -447
rect 177 -448 192 -447
rect 278 -448 297 -447
rect 303 -448 458 -447
rect 499 -448 528 -447
rect 86 -450 244 -449
rect 282 -450 363 -449
rect 380 -450 430 -449
rect 93 -452 465 -451
rect 93 -454 115 -453
rect 121 -454 213 -453
rect 243 -454 374 -453
rect 429 -454 563 -453
rect 96 -456 118 -455
rect 138 -456 251 -455
rect 296 -456 395 -455
rect 534 -456 563 -455
rect 100 -458 185 -457
rect 191 -458 346 -457
rect 145 -460 227 -459
rect 254 -460 535 -459
rect 149 -462 164 -461
rect 170 -462 402 -461
rect 58 -464 164 -463
rect 254 -464 265 -463
rect 310 -464 479 -463
rect 58 -466 132 -465
rect 156 -466 234 -465
rect 317 -466 353 -465
rect 37 -468 132 -467
rect 320 -468 367 -467
rect 23 -470 38 -469
rect 201 -470 367 -469
rect 23 -472 143 -471
rect 324 -472 472 -471
rect 135 -474 143 -473
rect 324 -474 500 -473
rect 107 -476 136 -475
rect 327 -476 444 -475
rect 107 -478 139 -477
rect 327 -478 647 -477
rect 124 -480 444 -479
rect 331 -482 409 -481
rect 331 -484 542 -483
rect 334 -486 381 -485
rect 450 -486 542 -485
rect 450 -488 570 -487
rect 485 -490 570 -489
rect 422 -492 486 -491
rect 2 -503 48 -502
rect 51 -503 125 -502
rect 128 -503 213 -502
rect 236 -503 458 -502
rect 492 -503 563 -502
rect 597 -503 629 -502
rect 635 -503 675 -502
rect 9 -505 174 -504
rect 205 -505 416 -504
rect 422 -505 465 -504
rect 492 -505 570 -504
rect 597 -505 647 -504
rect 16 -507 192 -506
rect 208 -507 220 -506
rect 240 -507 444 -506
rect 464 -507 549 -506
rect 604 -507 615 -506
rect 618 -507 668 -506
rect 16 -509 76 -508
rect 79 -509 265 -508
rect 289 -509 307 -508
rect 310 -509 416 -508
rect 513 -509 605 -508
rect 639 -509 647 -508
rect 23 -511 199 -510
rect 212 -511 335 -510
rect 345 -511 549 -510
rect 576 -511 619 -510
rect 23 -513 31 -512
rect 37 -513 395 -512
rect 397 -513 528 -512
rect 30 -515 73 -514
rect 86 -515 153 -514
rect 170 -515 507 -514
rect 513 -515 556 -514
rect 51 -517 332 -516
rect 334 -517 570 -516
rect 58 -519 209 -518
rect 303 -519 500 -518
rect 527 -519 654 -518
rect 86 -521 283 -520
rect 310 -521 367 -520
rect 369 -521 500 -520
rect 555 -521 591 -520
rect 621 -521 654 -520
rect 93 -523 115 -522
rect 131 -523 563 -522
rect 590 -523 626 -522
rect 93 -525 279 -524
rect 282 -525 353 -524
rect 355 -525 479 -524
rect 495 -525 507 -524
rect 625 -525 643 -524
rect 100 -527 185 -526
rect 191 -527 227 -526
rect 275 -527 304 -526
rect 324 -527 430 -526
rect 478 -527 535 -526
rect 100 -529 164 -528
rect 170 -529 220 -528
rect 226 -529 269 -528
rect 275 -529 472 -528
rect 485 -529 535 -528
rect 107 -531 290 -530
rect 324 -531 391 -530
rect 397 -531 612 -530
rect 107 -533 150 -532
rect 163 -533 612 -532
rect 65 -535 150 -534
rect 177 -535 241 -534
rect 348 -535 444 -534
rect 457 -535 486 -534
rect 61 -537 178 -536
rect 198 -537 255 -536
rect 362 -537 451 -536
rect 121 -539 132 -538
rect 135 -539 157 -538
rect 205 -539 472 -538
rect 142 -541 234 -540
rect 254 -541 314 -540
rect 366 -541 409 -540
rect 429 -541 521 -540
rect 145 -543 633 -542
rect 156 -545 360 -544
rect 373 -545 412 -544
rect 436 -545 451 -544
rect 520 -545 584 -544
rect 632 -545 640 -544
rect 271 -547 584 -546
rect 338 -549 437 -548
rect 296 -551 339 -550
rect 373 -551 402 -550
rect 296 -553 318 -552
rect 380 -553 426 -552
rect 247 -555 318 -554
rect 380 -555 577 -554
rect 247 -557 269 -556
rect 383 -557 388 -556
rect 2 -568 94 -567
rect 100 -568 143 -567
rect 156 -568 241 -567
rect 254 -568 356 -567
rect 369 -568 465 -567
rect 485 -568 556 -567
rect 576 -568 612 -567
rect 618 -568 629 -567
rect 642 -568 654 -567
rect 9 -570 101 -569
rect 114 -570 150 -569
rect 170 -570 213 -569
rect 233 -570 269 -569
rect 271 -570 318 -569
rect 352 -570 591 -569
rect 646 -570 654 -569
rect 16 -572 104 -571
rect 114 -572 136 -571
rect 142 -572 206 -571
rect 208 -572 230 -571
rect 261 -572 405 -571
rect 408 -572 605 -571
rect 16 -574 311 -573
rect 331 -574 591 -573
rect 23 -576 80 -575
rect 82 -576 94 -575
rect 135 -576 258 -575
rect 268 -576 325 -575
rect 373 -576 577 -575
rect 583 -576 619 -575
rect 23 -578 192 -577
rect 194 -578 227 -577
rect 278 -578 318 -577
rect 324 -578 451 -577
rect 464 -578 472 -577
rect 544 -578 598 -577
rect 30 -580 381 -579
rect 383 -580 412 -579
rect 429 -580 433 -579
rect 450 -580 626 -579
rect 30 -582 73 -581
rect 79 -582 164 -581
rect 170 -582 185 -581
rect 198 -582 202 -581
rect 205 -582 409 -581
rect 429 -582 479 -581
rect 506 -582 598 -581
rect 51 -584 234 -583
rect 303 -584 335 -583
rect 387 -584 521 -583
rect 565 -584 605 -583
rect 51 -586 122 -585
rect 152 -586 164 -585
rect 177 -586 262 -585
rect 296 -586 304 -585
rect 310 -586 437 -585
rect 443 -586 479 -585
rect 506 -586 549 -585
rect 569 -586 584 -585
rect 61 -588 241 -587
rect 264 -588 437 -587
rect 471 -588 500 -587
rect 520 -588 535 -587
rect 548 -588 563 -587
rect 65 -590 297 -589
rect 345 -590 500 -589
rect 527 -590 570 -589
rect 68 -592 129 -591
rect 152 -592 339 -591
rect 394 -592 486 -591
rect 534 -592 542 -591
rect 72 -594 220 -593
rect 226 -594 283 -593
rect 338 -594 363 -593
rect 401 -594 514 -593
rect 58 -596 220 -595
rect 247 -596 395 -595
rect 401 -596 493 -595
rect 86 -598 349 -597
rect 432 -598 444 -597
rect 457 -598 514 -597
rect 86 -600 192 -599
rect 198 -600 556 -599
rect 107 -602 185 -601
rect 212 -602 353 -601
rect 492 -602 622 -601
rect 37 -604 108 -603
rect 121 -604 374 -603
rect 37 -606 45 -605
rect 156 -606 178 -605
rect 180 -606 248 -605
rect 282 -606 416 -605
rect 44 -608 125 -607
rect 348 -608 367 -607
rect 415 -608 423 -607
rect 359 -610 423 -609
rect 359 -612 388 -611
rect 2 -623 129 -622
rect 131 -623 209 -622
rect 212 -623 335 -622
rect 345 -623 570 -622
rect 625 -623 640 -622
rect 2 -625 94 -624
rect 100 -625 153 -624
rect 173 -625 584 -624
rect 9 -627 206 -626
rect 208 -627 605 -626
rect 9 -629 69 -628
rect 103 -629 195 -628
rect 201 -629 262 -628
rect 296 -629 328 -628
rect 334 -629 563 -628
rect 565 -629 591 -628
rect 16 -631 279 -630
rect 289 -631 297 -630
rect 313 -631 430 -630
rect 443 -631 479 -630
rect 513 -631 542 -630
rect 16 -633 132 -632
rect 184 -633 360 -632
rect 362 -633 598 -632
rect 23 -635 178 -634
rect 219 -635 332 -634
rect 348 -635 577 -634
rect 23 -637 97 -636
rect 107 -637 111 -636
rect 114 -637 139 -636
rect 170 -637 185 -636
rect 219 -637 402 -636
rect 443 -637 493 -636
rect 520 -637 559 -636
rect 30 -639 153 -638
rect 177 -639 381 -638
rect 429 -639 493 -638
rect 520 -639 549 -638
rect 30 -641 279 -640
rect 324 -641 549 -640
rect 37 -643 66 -642
rect 107 -643 164 -642
rect 222 -643 318 -642
rect 324 -643 405 -642
rect 460 -643 612 -642
rect 37 -645 143 -644
rect 226 -645 388 -644
rect 527 -645 619 -644
rect 44 -647 199 -646
rect 226 -647 248 -646
rect 257 -647 465 -646
rect 44 -649 206 -648
rect 240 -649 290 -648
rect 303 -649 318 -648
rect 338 -649 381 -648
rect 387 -649 395 -648
rect 436 -649 528 -648
rect 51 -651 202 -650
rect 247 -651 458 -650
rect 51 -653 262 -652
rect 275 -653 339 -652
rect 345 -653 405 -652
rect 408 -653 437 -652
rect 58 -655 171 -654
rect 282 -655 304 -654
rect 310 -655 465 -654
rect 61 -657 556 -656
rect 65 -659 230 -658
rect 268 -659 311 -658
rect 313 -659 458 -658
rect 513 -659 556 -658
rect 72 -661 269 -660
rect 352 -661 374 -660
rect 408 -661 451 -660
rect 72 -663 129 -662
rect 135 -663 143 -662
rect 180 -663 451 -662
rect 79 -665 241 -664
rect 355 -665 423 -664
rect 79 -667 136 -666
rect 191 -667 374 -666
rect 422 -667 535 -666
rect 110 -669 164 -668
rect 366 -669 398 -668
rect 506 -669 535 -668
rect 121 -671 234 -670
rect 369 -671 472 -670
rect 485 -671 507 -670
rect 86 -673 234 -672
rect 257 -673 472 -672
rect 86 -675 150 -674
rect 394 -675 486 -674
rect 121 -677 213 -676
rect 2 -688 206 -687
rect 219 -688 286 -687
rect 289 -688 307 -687
rect 313 -688 416 -687
rect 422 -688 426 -687
rect 429 -688 451 -687
rect 457 -688 612 -687
rect 632 -688 640 -687
rect 2 -690 59 -689
rect 96 -690 174 -689
rect 177 -690 255 -689
rect 278 -690 297 -689
rect 331 -690 458 -689
rect 478 -690 584 -689
rect 9 -692 122 -691
rect 135 -692 157 -691
rect 170 -692 192 -691
rect 194 -692 227 -691
rect 229 -692 591 -691
rect 12 -694 395 -693
rect 397 -694 549 -693
rect 562 -694 664 -693
rect 16 -696 118 -695
rect 121 -696 181 -695
rect 187 -696 563 -695
rect 16 -698 94 -697
rect 114 -698 577 -697
rect 30 -700 129 -699
rect 156 -700 213 -699
rect 219 -700 262 -699
rect 271 -700 332 -699
rect 338 -700 598 -699
rect 30 -702 108 -701
rect 114 -702 479 -701
rect 485 -702 570 -701
rect 37 -704 258 -703
rect 278 -704 402 -703
rect 404 -704 556 -703
rect 37 -706 87 -705
rect 117 -706 297 -705
rect 341 -706 444 -705
rect 464 -706 549 -705
rect 44 -708 48 -707
rect 51 -708 262 -707
rect 345 -708 416 -707
rect 432 -708 507 -707
rect 520 -708 619 -707
rect 54 -710 241 -709
rect 247 -710 286 -709
rect 292 -710 507 -709
rect 527 -710 626 -709
rect 82 -712 213 -711
rect 226 -712 472 -711
rect 492 -712 605 -711
rect 86 -714 143 -713
rect 145 -714 528 -713
rect 100 -716 248 -715
rect 254 -716 374 -715
rect 376 -716 542 -715
rect 128 -718 185 -717
rect 198 -718 325 -717
rect 345 -718 367 -717
rect 376 -718 647 -717
rect 107 -720 199 -719
rect 233 -720 370 -719
rect 380 -720 633 -719
rect 149 -722 339 -721
rect 355 -722 451 -721
rect 499 -722 521 -721
rect 72 -724 500 -723
rect 72 -726 80 -725
rect 149 -726 311 -725
rect 359 -726 486 -725
rect 163 -728 241 -727
rect 268 -728 325 -727
rect 359 -728 535 -727
rect 166 -730 444 -729
rect 513 -730 535 -729
rect 177 -732 202 -731
rect 268 -732 640 -731
rect 191 -734 234 -733
rect 275 -734 542 -733
rect 187 -736 276 -735
rect 303 -736 493 -735
rect 310 -738 353 -737
rect 366 -738 657 -737
rect 352 -740 388 -739
rect 408 -740 465 -739
rect 282 -742 388 -741
rect 436 -742 514 -741
rect 362 -744 437 -743
rect 2 -755 164 -754
rect 184 -755 255 -754
rect 261 -755 363 -754
rect 373 -755 437 -754
rect 471 -755 626 -754
rect 23 -757 388 -756
rect 471 -757 542 -756
rect 558 -757 647 -756
rect 23 -759 101 -758
rect 114 -759 241 -758
rect 243 -759 297 -758
rect 299 -759 598 -758
rect 30 -761 104 -760
rect 114 -761 136 -760
rect 142 -761 605 -760
rect 30 -763 108 -762
rect 117 -763 255 -762
rect 261 -763 346 -762
rect 376 -763 584 -762
rect 597 -763 605 -762
rect 37 -765 150 -764
rect 152 -765 164 -764
rect 187 -765 395 -764
rect 474 -765 556 -764
rect 583 -765 612 -764
rect 54 -767 353 -766
rect 376 -767 619 -766
rect 61 -769 640 -768
rect 65 -771 230 -770
rect 268 -771 318 -770
rect 327 -771 416 -770
rect 443 -771 556 -770
rect 618 -771 661 -770
rect 65 -773 157 -772
rect 191 -773 339 -772
rect 345 -773 360 -772
rect 380 -773 514 -772
rect 541 -773 591 -772
rect 79 -775 549 -774
rect 82 -777 493 -776
rect 44 -779 83 -778
rect 86 -779 206 -778
rect 208 -779 577 -778
rect 96 -781 101 -780
rect 107 -781 122 -780
rect 145 -781 171 -780
rect 198 -781 479 -780
rect 93 -783 122 -782
rect 149 -783 206 -782
rect 219 -783 227 -782
rect 268 -783 311 -782
rect 331 -783 514 -782
rect 156 -785 178 -784
rect 219 -785 654 -784
rect 58 -787 178 -786
rect 275 -787 325 -786
rect 359 -787 367 -786
rect 373 -787 591 -786
rect 58 -789 73 -788
rect 170 -789 283 -788
rect 285 -789 500 -788
rect 72 -791 129 -790
rect 275 -791 633 -790
rect 278 -793 465 -792
rect 499 -793 521 -792
rect 198 -795 279 -794
rect 289 -795 409 -794
rect 411 -795 549 -794
rect 212 -797 409 -796
rect 415 -797 528 -796
rect 152 -799 213 -798
rect 233 -799 290 -798
rect 303 -799 332 -798
rect 380 -799 430 -798
rect 443 -799 535 -798
rect 51 -801 234 -800
rect 310 -801 507 -800
rect 527 -801 563 -800
rect 320 -803 367 -802
rect 387 -803 521 -802
rect 562 -803 570 -802
rect 341 -805 507 -804
rect 341 -807 437 -806
rect 450 -807 577 -806
rect 390 -809 493 -808
rect 394 -811 402 -810
rect 422 -811 430 -810
rect 450 -811 486 -810
rect 313 -813 423 -812
rect 457 -813 486 -812
rect 457 -815 538 -814
rect 464 -817 570 -816
rect 9 -828 34 -827
rect 40 -828 97 -827
rect 107 -828 136 -827
rect 149 -828 230 -827
rect 233 -828 374 -827
rect 387 -828 409 -827
rect 425 -828 493 -827
rect 513 -828 563 -827
rect 572 -828 619 -827
rect 16 -830 38 -829
rect 54 -830 472 -829
rect 478 -830 542 -829
rect 555 -830 591 -829
rect 30 -832 94 -831
rect 107 -832 185 -831
rect 194 -832 213 -831
rect 222 -832 286 -831
rect 292 -832 493 -831
rect 534 -832 584 -831
rect 58 -834 87 -833
rect 89 -834 101 -833
rect 114 -834 146 -833
rect 170 -834 325 -833
rect 334 -834 549 -833
rect 562 -834 577 -833
rect 23 -836 171 -835
rect 180 -836 241 -835
rect 247 -836 251 -835
rect 268 -836 318 -835
rect 320 -836 437 -835
rect 478 -836 507 -835
rect 548 -836 605 -835
rect 23 -838 45 -837
rect 51 -838 101 -837
rect 114 -838 199 -837
rect 226 -838 276 -837
rect 303 -838 374 -837
rect 401 -838 451 -837
rect 499 -838 507 -837
rect 51 -840 62 -839
rect 65 -840 202 -839
rect 247 -840 290 -839
rect 317 -840 500 -839
rect 65 -842 164 -841
rect 173 -842 269 -841
rect 320 -842 409 -841
rect 422 -842 472 -841
rect 72 -844 129 -843
rect 135 -844 216 -843
rect 250 -844 290 -843
rect 338 -844 381 -843
rect 404 -844 521 -843
rect 72 -846 83 -845
rect 86 -846 220 -845
rect 254 -846 339 -845
rect 345 -846 517 -845
rect 93 -848 143 -847
rect 163 -848 283 -847
rect 348 -848 458 -847
rect 121 -850 153 -849
rect 177 -850 276 -849
rect 352 -850 360 -849
rect 376 -850 402 -849
rect 436 -850 444 -849
rect 121 -852 157 -851
rect 184 -852 192 -851
rect 198 -852 311 -851
rect 331 -852 444 -851
rect 2 -854 192 -853
rect 205 -854 255 -853
rect 261 -854 304 -853
rect 345 -854 360 -853
rect 128 -856 279 -855
rect 296 -856 332 -855
rect 355 -856 528 -855
rect 156 -858 206 -857
rect 226 -858 458 -857
rect 520 -858 528 -857
rect 233 -860 262 -859
rect 296 -860 381 -859
rect 2 -871 136 -870
rect 152 -871 388 -870
rect 425 -871 500 -870
rect 516 -871 545 -870
rect 2 -873 115 -872
rect 121 -873 174 -872
rect 205 -873 234 -872
rect 247 -873 321 -872
rect 345 -873 402 -872
rect 443 -873 549 -872
rect 9 -875 45 -874
rect 47 -875 104 -874
rect 135 -875 150 -874
rect 156 -875 234 -874
rect 240 -875 248 -874
rect 261 -875 297 -874
rect 299 -875 388 -874
rect 401 -875 451 -874
rect 453 -875 486 -874
rect 520 -875 535 -874
rect 537 -875 542 -874
rect 548 -875 556 -874
rect 16 -877 31 -876
rect 44 -877 52 -876
rect 54 -877 125 -876
rect 142 -877 241 -876
rect 268 -877 500 -876
rect 520 -877 531 -876
rect 16 -879 41 -878
rect 61 -879 73 -878
rect 79 -879 129 -878
rect 173 -879 374 -878
rect 376 -879 465 -878
rect 485 -879 507 -878
rect 527 -879 563 -878
rect 23 -881 38 -880
rect 65 -881 164 -880
rect 191 -881 465 -880
rect 478 -881 507 -880
rect 23 -883 132 -882
rect 163 -883 185 -882
rect 208 -883 339 -882
rect 348 -883 353 -882
rect 380 -883 437 -882
rect 68 -885 87 -884
rect 93 -885 202 -884
rect 212 -885 276 -884
rect 282 -885 374 -884
rect 422 -885 528 -884
rect 79 -887 178 -886
rect 194 -887 339 -886
rect 352 -887 367 -886
rect 86 -889 108 -888
rect 121 -889 185 -888
rect 198 -889 381 -888
rect 96 -891 150 -890
rect 219 -891 269 -890
rect 275 -891 290 -890
rect 292 -891 416 -890
rect 100 -893 157 -892
rect 191 -893 220 -892
rect 222 -893 367 -892
rect 415 -893 430 -892
rect 100 -895 115 -894
rect 226 -895 325 -894
rect 331 -895 437 -894
rect 37 -897 332 -896
rect 408 -897 430 -896
rect 229 -899 255 -898
rect 282 -899 514 -898
rect 208 -901 514 -900
rect 243 -903 479 -902
rect 254 -905 290 -904
rect 292 -905 472 -904
rect 303 -907 314 -906
rect 317 -907 360 -906
rect 394 -907 409 -906
rect 65 -909 395 -908
rect 306 -911 447 -910
rect 310 -913 451 -912
rect 324 -915 472 -914
rect 9 -926 395 -925
rect 429 -926 444 -925
rect 450 -926 472 -925
rect 474 -926 486 -925
rect 506 -926 510 -925
rect 530 -926 549 -925
rect 16 -928 31 -927
rect 37 -928 171 -927
rect 173 -928 482 -927
rect 485 -928 521 -927
rect 23 -930 73 -929
rect 79 -930 146 -929
rect 149 -930 332 -929
rect 359 -930 479 -929
rect 506 -930 521 -929
rect 23 -932 118 -931
rect 163 -932 199 -931
rect 201 -932 388 -931
rect 415 -932 430 -931
rect 450 -932 493 -931
rect 44 -934 125 -933
rect 184 -934 248 -933
rect 264 -934 437 -933
rect 478 -934 542 -933
rect 54 -936 199 -935
rect 208 -936 213 -935
rect 226 -936 423 -935
rect 436 -936 500 -935
rect 58 -938 87 -937
rect 93 -938 241 -937
rect 268 -938 272 -937
rect 285 -938 384 -937
rect 387 -938 402 -937
rect 499 -938 535 -937
rect 58 -940 143 -939
rect 177 -940 241 -939
rect 268 -940 325 -939
rect 345 -940 416 -939
rect 2 -942 143 -941
rect 152 -942 178 -941
rect 187 -942 213 -941
rect 233 -942 248 -941
rect 271 -942 325 -941
rect 338 -942 346 -941
rect 359 -942 367 -941
rect 373 -942 402 -941
rect 30 -944 234 -943
rect 243 -944 367 -943
rect 373 -944 468 -943
rect 72 -946 255 -945
rect 299 -946 318 -945
rect 320 -946 395 -945
rect 79 -948 111 -947
rect 114 -948 122 -947
rect 187 -948 465 -947
rect 68 -950 465 -949
rect 86 -952 311 -951
rect 338 -952 412 -951
rect 93 -954 185 -953
rect 191 -954 206 -953
rect 208 -954 514 -953
rect 96 -956 290 -955
rect 303 -956 332 -955
rect 362 -956 409 -955
rect 100 -958 157 -957
rect 194 -958 220 -957
rect 254 -958 262 -957
rect 282 -958 304 -957
rect 306 -958 353 -957
rect 100 -960 153 -959
rect 170 -960 262 -959
rect 289 -960 297 -959
rect 310 -960 381 -959
rect 110 -962 115 -961
rect 128 -962 283 -961
rect 352 -962 493 -961
rect 135 -964 157 -963
rect 219 -964 276 -963
rect 65 -966 276 -965
rect 135 -968 167 -967
rect 16 -979 80 -978
rect 107 -979 188 -978
rect 219 -979 276 -978
rect 292 -979 325 -978
rect 331 -979 486 -978
rect 520 -979 528 -978
rect 23 -981 265 -980
rect 320 -981 402 -980
rect 408 -981 433 -980
rect 464 -981 500 -980
rect 26 -983 38 -982
rect 51 -983 136 -982
rect 156 -983 209 -982
rect 261 -983 346 -982
rect 352 -983 472 -982
rect 30 -985 230 -984
rect 271 -985 353 -984
rect 380 -985 444 -984
rect 446 -985 465 -984
rect 471 -985 493 -984
rect 37 -987 132 -986
rect 135 -987 192 -986
rect 208 -987 300 -986
rect 303 -987 346 -986
rect 411 -987 430 -986
rect 58 -989 129 -988
rect 131 -989 213 -988
rect 229 -989 255 -988
rect 278 -989 402 -988
rect 422 -989 458 -988
rect 58 -991 101 -990
rect 107 -991 122 -990
rect 128 -991 199 -990
rect 212 -991 290 -990
rect 296 -991 381 -990
rect 390 -991 423 -990
rect 429 -991 510 -990
rect 65 -993 115 -992
rect 121 -993 185 -992
rect 191 -993 262 -992
rect 299 -993 311 -992
rect 324 -993 416 -992
rect 443 -993 458 -992
rect 65 -995 118 -994
rect 156 -995 171 -994
rect 173 -995 202 -994
rect 233 -995 290 -994
rect 303 -995 339 -994
rect 394 -995 416 -994
rect 68 -997 94 -996
rect 100 -997 118 -996
rect 149 -997 171 -996
rect 177 -997 227 -996
rect 240 -997 311 -996
rect 338 -997 374 -996
rect 394 -997 437 -996
rect 30 -999 69 -998
rect 72 -999 220 -998
rect 236 -999 241 -998
rect 366 -999 374 -998
rect 436 -999 451 -998
rect 72 -1001 87 -1000
rect 110 -1001 360 -1000
rect 79 -1003 97 -1002
rect 163 -1003 206 -1002
rect 317 -1003 367 -1002
rect 177 -1005 283 -1004
rect 359 -1005 388 -1004
rect 198 -1007 332 -1006
rect 201 -1009 255 -1008
rect 268 -1009 388 -1008
rect 30 -1020 48 -1019
rect 51 -1020 202 -1019
rect 208 -1020 220 -1019
rect 247 -1020 269 -1019
rect 278 -1020 339 -1019
rect 355 -1020 381 -1019
rect 436 -1020 444 -1019
rect 453 -1020 472 -1019
rect 523 -1020 528 -1019
rect 58 -1022 97 -1021
rect 114 -1022 237 -1021
rect 240 -1022 269 -1021
rect 289 -1022 395 -1021
rect 443 -1022 451 -1021
rect 453 -1022 465 -1021
rect 516 -1022 524 -1021
rect 16 -1024 115 -1023
rect 121 -1024 195 -1023
rect 205 -1024 241 -1023
rect 247 -1024 283 -1023
rect 296 -1024 304 -1023
rect 324 -1024 335 -1023
rect 359 -1024 367 -1023
rect 369 -1024 402 -1023
rect 520 -1024 528 -1023
rect 65 -1026 80 -1025
rect 86 -1026 104 -1025
rect 107 -1026 122 -1025
rect 142 -1026 167 -1025
rect 177 -1026 220 -1025
rect 229 -1026 395 -1025
rect 72 -1028 129 -1027
rect 135 -1028 178 -1027
rect 184 -1028 202 -1027
rect 208 -1028 213 -1027
rect 215 -1028 304 -1027
rect 324 -1028 328 -1027
rect 380 -1028 409 -1027
rect 72 -1030 90 -1029
rect 93 -1030 101 -1029
rect 107 -1030 293 -1029
rect 387 -1030 409 -1029
rect 86 -1032 118 -1031
rect 135 -1032 150 -1031
rect 156 -1032 192 -1031
rect 212 -1032 360 -1031
rect 37 -1034 150 -1033
rect 163 -1034 185 -1033
rect 187 -1034 255 -1033
rect 261 -1034 339 -1033
rect 117 -1036 227 -1035
rect 233 -1036 293 -1035
rect 331 -1036 388 -1035
rect 170 -1038 230 -1037
rect 250 -1038 346 -1037
rect 226 -1040 374 -1039
rect 261 -1042 276 -1041
rect 285 -1042 402 -1041
rect 275 -1044 318 -1043
rect 345 -1044 353 -1043
rect 373 -1044 430 -1043
rect 254 -1046 318 -1045
rect 51 -1057 118 -1056
rect 128 -1057 181 -1056
rect 201 -1057 304 -1056
rect 320 -1057 381 -1056
rect 429 -1057 437 -1056
rect 457 -1057 465 -1056
rect 520 -1057 528 -1056
rect 61 -1059 90 -1058
rect 93 -1059 104 -1058
rect 107 -1059 255 -1058
rect 334 -1059 374 -1058
rect 408 -1059 430 -1058
rect 65 -1061 80 -1060
rect 93 -1061 150 -1060
rect 152 -1061 262 -1060
rect 359 -1061 363 -1060
rect 373 -1061 381 -1060
rect 408 -1061 416 -1060
rect 65 -1063 132 -1062
rect 135 -1063 160 -1062
rect 163 -1063 167 -1062
rect 177 -1063 209 -1062
rect 212 -1063 276 -1062
rect 359 -1063 367 -1062
rect 72 -1065 111 -1064
rect 135 -1065 300 -1064
rect 366 -1065 402 -1064
rect 75 -1067 108 -1066
rect 145 -1067 216 -1066
rect 219 -1067 223 -1066
rect 226 -1067 248 -1066
rect 250 -1067 388 -1066
rect 394 -1067 402 -1066
rect 100 -1069 143 -1068
rect 149 -1069 234 -1068
rect 236 -1069 423 -1068
rect 156 -1071 206 -1070
rect 219 -1071 332 -1070
rect 163 -1073 171 -1072
rect 177 -1073 199 -1072
rect 236 -1073 353 -1072
rect 184 -1075 213 -1074
rect 247 -1075 293 -1074
rect 306 -1075 388 -1074
rect 191 -1077 206 -1076
rect 254 -1077 269 -1076
rect 275 -1077 318 -1076
rect 362 -1077 395 -1076
rect 142 -1079 318 -1078
rect 261 -1081 290 -1080
rect 268 -1083 283 -1082
rect 289 -1083 339 -1082
rect 282 -1085 391 -1084
rect 324 -1087 339 -1086
rect 310 -1089 325 -1088
rect 296 -1091 311 -1090
rect 30 -1102 94 -1101
rect 100 -1102 111 -1101
rect 114 -1102 223 -1101
rect 226 -1102 444 -1101
rect 460 -1102 465 -1101
rect 37 -1104 237 -1103
rect 254 -1104 300 -1103
rect 306 -1104 346 -1103
rect 352 -1104 419 -1103
rect 422 -1104 437 -1103
rect 51 -1106 90 -1105
rect 100 -1106 115 -1105
rect 121 -1106 139 -1105
rect 142 -1106 178 -1105
rect 184 -1106 248 -1105
rect 254 -1106 353 -1105
rect 359 -1106 374 -1105
rect 387 -1106 409 -1105
rect 415 -1106 430 -1105
rect 54 -1108 59 -1107
rect 65 -1108 188 -1107
rect 219 -1108 304 -1107
rect 317 -1108 339 -1107
rect 345 -1108 360 -1107
rect 362 -1108 367 -1107
rect 380 -1108 409 -1107
rect 65 -1110 157 -1109
rect 163 -1110 192 -1109
rect 226 -1110 241 -1109
rect 247 -1110 269 -1109
rect 320 -1110 374 -1109
rect 394 -1110 423 -1109
rect 72 -1112 80 -1111
rect 82 -1112 87 -1111
rect 121 -1112 136 -1111
rect 142 -1112 150 -1111
rect 159 -1112 164 -1111
rect 170 -1112 185 -1111
rect 191 -1112 209 -1111
rect 233 -1112 377 -1111
rect 401 -1112 430 -1111
rect 44 -1114 80 -1113
rect 107 -1114 136 -1113
rect 170 -1114 213 -1113
rect 268 -1114 283 -1113
rect 289 -1114 321 -1113
rect 324 -1114 381 -1113
rect 75 -1116 108 -1115
rect 131 -1116 150 -1115
rect 198 -1116 213 -1115
rect 278 -1116 395 -1115
rect 205 -1118 241 -1117
rect 282 -1118 311 -1117
rect 331 -1118 416 -1117
rect 194 -1120 311 -1119
rect 338 -1120 370 -1119
rect 205 -1122 388 -1121
rect 261 -1124 332 -1123
rect 180 -1126 262 -1125
rect 296 -1126 402 -1125
rect 264 -1128 297 -1127
rect 30 -1139 97 -1138
rect 107 -1139 129 -1138
rect 149 -1139 199 -1138
rect 205 -1139 241 -1138
rect 250 -1139 269 -1138
rect 275 -1139 381 -1138
rect 397 -1139 437 -1138
rect 478 -1139 486 -1138
rect 37 -1141 171 -1140
rect 184 -1141 199 -1140
rect 229 -1141 276 -1140
rect 296 -1141 325 -1140
rect 327 -1141 402 -1140
rect 44 -1143 55 -1142
rect 58 -1143 73 -1142
rect 75 -1143 83 -1142
rect 86 -1143 244 -1142
rect 254 -1143 444 -1142
rect 65 -1145 160 -1144
rect 163 -1145 174 -1144
rect 184 -1145 206 -1144
rect 261 -1145 283 -1144
rect 299 -1145 416 -1144
rect 79 -1147 101 -1146
rect 107 -1147 122 -1146
rect 128 -1147 304 -1146
rect 306 -1147 430 -1146
rect 89 -1149 115 -1148
rect 117 -1149 167 -1148
rect 201 -1149 283 -1148
rect 306 -1149 360 -1148
rect 369 -1149 409 -1148
rect 93 -1151 209 -1150
rect 261 -1151 374 -1150
rect 376 -1151 423 -1150
rect 100 -1153 125 -1152
rect 149 -1153 192 -1152
rect 208 -1153 395 -1152
rect 401 -1153 409 -1152
rect 117 -1155 227 -1154
rect 268 -1155 290 -1154
rect 310 -1155 381 -1154
rect 121 -1157 136 -1156
rect 156 -1157 171 -1156
rect 191 -1157 220 -1156
rect 278 -1157 311 -1156
rect 317 -1157 332 -1156
rect 338 -1157 367 -1156
rect 135 -1159 146 -1158
rect 163 -1159 290 -1158
rect 212 -1161 227 -1160
rect 240 -1161 339 -1160
rect 142 -1163 213 -1162
rect 219 -1163 234 -1162
rect 264 -1163 332 -1162
rect 233 -1165 248 -1164
rect 264 -1165 388 -1164
rect 352 -1167 388 -1166
rect 345 -1169 353 -1168
rect 254 -1171 346 -1170
rect 61 -1182 73 -1181
rect 79 -1182 136 -1181
rect 163 -1182 185 -1181
rect 198 -1182 206 -1181
rect 208 -1182 213 -1181
rect 240 -1182 283 -1181
rect 292 -1182 402 -1181
rect 72 -1184 115 -1183
rect 121 -1184 150 -1183
rect 177 -1184 209 -1183
rect 212 -1184 241 -1183
rect 247 -1184 269 -1183
rect 303 -1184 381 -1183
rect 86 -1186 171 -1185
rect 173 -1186 248 -1185
rect 250 -1186 374 -1185
rect 376 -1186 395 -1185
rect 65 -1188 171 -1187
rect 184 -1188 227 -1187
rect 254 -1188 346 -1187
rect 366 -1188 381 -1187
rect 93 -1190 125 -1189
rect 128 -1190 199 -1189
rect 201 -1190 269 -1189
rect 324 -1190 328 -1189
rect 366 -1190 388 -1189
rect 107 -1192 132 -1191
rect 194 -1192 283 -1191
rect 324 -1192 339 -1191
rect 383 -1192 388 -1191
rect 100 -1194 108 -1193
rect 114 -1194 157 -1193
rect 233 -1194 346 -1193
rect 100 -1196 262 -1195
rect 338 -1196 353 -1195
rect 121 -1198 220 -1197
rect 233 -1198 297 -1197
rect 327 -1198 353 -1197
rect 142 -1200 157 -1199
rect 191 -1200 220 -1199
rect 257 -1200 276 -1199
rect 296 -1200 311 -1199
rect 138 -1202 192 -1201
rect 275 -1202 290 -1201
rect 310 -1202 318 -1201
rect 65 -1213 192 -1212
rect 194 -1213 248 -1212
rect 261 -1213 290 -1212
rect 292 -1213 353 -1212
rect 380 -1213 388 -1212
rect 72 -1215 90 -1214
rect 114 -1215 157 -1214
rect 170 -1215 248 -1214
rect 261 -1215 374 -1214
rect 383 -1215 395 -1214
rect 79 -1217 139 -1216
rect 149 -1217 220 -1216
rect 240 -1217 360 -1216
rect 107 -1219 115 -1218
rect 121 -1219 244 -1218
rect 264 -1219 346 -1218
rect 352 -1219 367 -1218
rect 121 -1221 181 -1220
rect 184 -1221 227 -1220
rect 275 -1221 318 -1220
rect 324 -1221 332 -1220
rect 128 -1223 160 -1222
rect 177 -1223 255 -1222
rect 268 -1223 318 -1222
rect 331 -1223 339 -1222
rect 100 -1225 129 -1224
rect 135 -1225 188 -1224
rect 205 -1225 213 -1224
rect 233 -1225 269 -1224
rect 303 -1225 311 -1224
rect 142 -1227 181 -1226
rect 198 -1227 234 -1226
rect 240 -1227 255 -1226
rect 282 -1227 311 -1226
rect 142 -1229 153 -1228
rect 212 -1229 230 -1228
rect 282 -1229 297 -1228
rect 275 -1231 297 -1230
rect 82 -1242 87 -1241
rect 93 -1242 101 -1241
rect 107 -1242 118 -1241
rect 128 -1242 153 -1241
rect 156 -1242 202 -1241
rect 212 -1242 220 -1241
rect 233 -1242 262 -1241
rect 275 -1242 297 -1241
rect 299 -1242 311 -1241
rect 317 -1242 321 -1241
rect 348 -1242 353 -1241
rect 100 -1244 122 -1243
rect 128 -1244 143 -1243
rect 156 -1244 227 -1243
rect 240 -1244 262 -1243
rect 282 -1244 304 -1243
rect 306 -1244 325 -1243
rect 110 -1246 115 -1245
rect 135 -1246 174 -1245
rect 177 -1246 192 -1245
rect 198 -1246 220 -1245
rect 226 -1246 234 -1245
rect 254 -1246 279 -1245
rect 285 -1246 290 -1245
rect 324 -1246 332 -1245
rect 135 -1248 150 -1247
rect 163 -1248 188 -1247
rect 191 -1248 206 -1247
rect 268 -1248 290 -1247
rect 180 -1250 248 -1249
rect 205 -1252 216 -1251
rect 240 -1252 248 -1251
rect 75 -1263 80 -1262
rect 100 -1263 129 -1262
rect 135 -1263 167 -1262
rect 170 -1263 174 -1262
rect 205 -1263 227 -1262
rect 254 -1263 272 -1262
rect 275 -1263 297 -1262
rect 320 -1263 325 -1262
rect 380 -1263 388 -1262
rect 114 -1265 122 -1264
rect 135 -1265 146 -1264
rect 163 -1265 178 -1264
rect 191 -1265 206 -1264
rect 215 -1265 220 -1264
rect 261 -1265 279 -1264
rect 117 -1267 122 -1266
rect 268 -1267 276 -1266
rect 86 -1278 97 -1277
rect 107 -1278 118 -1277
rect 121 -1278 129 -1277
rect 135 -1278 146 -1277
rect 149 -1278 160 -1277
rect 219 -1278 227 -1277
rect 275 -1278 283 -1277
rect 299 -1278 304 -1277
rect 383 -1278 388 -1277
rect 156 -1280 167 -1279
<< m2contact >>
rect 135 0 136 1
rect 142 0 143 1
rect 145 0 146 1
rect 156 0 157 1
rect 184 0 185 1
rect 194 0 195 1
rect 212 0 213 1
rect 219 0 220 1
rect 135 -11 136 -10
rect 149 -11 150 -10
rect 156 -11 157 -10
rect 180 -11 181 -10
rect 191 -11 192 -10
rect 198 -11 199 -10
rect 208 -11 209 -10
rect 212 -11 213 -10
rect 257 -11 258 -10
rect 261 -11 262 -10
rect 149 -13 150 -12
rect 152 -13 153 -12
rect 177 -13 178 -12
rect 184 -13 185 -12
rect 212 -13 213 -12
rect 222 -13 223 -12
rect 184 -15 185 -14
rect 205 -15 206 -14
rect 149 -26 150 -25
rect 166 -26 167 -25
rect 170 -26 171 -25
rect 184 -26 185 -25
rect 187 -26 188 -25
rect 191 -26 192 -25
rect 198 -26 199 -25
rect 219 -26 220 -25
rect 229 -26 230 -25
rect 261 -26 262 -25
rect 268 -26 269 -25
rect 271 -26 272 -25
rect 341 -26 342 -25
rect 345 -26 346 -25
rect 145 -28 146 -27
rect 149 -28 150 -27
rect 156 -28 157 -27
rect 173 -28 174 -27
rect 177 -28 178 -27
rect 208 -28 209 -27
rect 243 -28 244 -27
rect 247 -28 248 -27
rect 201 -30 202 -29
rect 212 -30 213 -29
rect 205 -32 206 -31
rect 240 -32 241 -31
rect 212 -34 213 -33
rect 233 -34 234 -33
rect 51 -45 52 -44
rect 54 -45 55 -44
rect 72 -45 73 -44
rect 96 -45 97 -44
rect 138 -45 139 -44
rect 149 -45 150 -44
rect 156 -45 157 -44
rect 198 -45 199 -44
rect 201 -45 202 -44
rect 219 -45 220 -44
rect 236 -45 237 -44
rect 247 -45 248 -44
rect 282 -45 283 -44
rect 289 -45 290 -44
rect 345 -45 346 -44
rect 352 -45 353 -44
rect 359 -45 360 -44
rect 366 -45 367 -44
rect 142 -47 143 -46
rect 198 -47 199 -46
rect 208 -47 209 -46
rect 212 -47 213 -46
rect 240 -47 241 -46
rect 243 -47 244 -46
rect 247 -47 248 -46
rect 261 -47 262 -46
rect 345 -47 346 -46
rect 362 -47 363 -46
rect 163 -49 164 -48
rect 187 -49 188 -48
rect 191 -49 192 -48
rect 205 -49 206 -48
rect 240 -49 241 -48
rect 296 -49 297 -48
rect 170 -51 171 -50
rect 275 -51 276 -50
rect 177 -53 178 -52
rect 191 -53 192 -52
rect 194 -53 195 -52
rect 219 -53 220 -52
rect 261 -53 262 -52
rect 268 -53 269 -52
rect 163 -55 164 -54
rect 177 -55 178 -54
rect 187 -55 188 -54
rect 212 -55 213 -54
rect 254 -55 255 -54
rect 268 -55 269 -54
rect 226 -57 227 -56
rect 254 -57 255 -56
rect 51 -68 52 -67
rect 72 -68 73 -67
rect 79 -68 80 -67
rect 142 -68 143 -67
rect 149 -68 150 -67
rect 187 -68 188 -67
rect 194 -68 195 -67
rect 212 -68 213 -67
rect 219 -68 220 -67
rect 275 -68 276 -67
rect 282 -68 283 -67
rect 376 -68 377 -67
rect 58 -70 59 -69
rect 145 -70 146 -69
rect 149 -70 150 -69
rect 243 -70 244 -69
rect 247 -70 248 -69
rect 303 -70 304 -69
rect 310 -70 311 -69
rect 317 -70 318 -69
rect 320 -70 321 -69
rect 331 -70 332 -69
rect 338 -70 339 -69
rect 348 -70 349 -69
rect 65 -72 66 -71
rect 170 -72 171 -71
rect 198 -72 199 -71
rect 282 -72 283 -71
rect 289 -72 290 -71
rect 310 -72 311 -71
rect 345 -72 346 -71
rect 352 -72 353 -71
rect 72 -74 73 -73
rect 86 -74 87 -73
rect 93 -74 94 -73
rect 138 -74 139 -73
rect 156 -74 157 -73
rect 187 -74 188 -73
rect 201 -74 202 -73
rect 254 -74 255 -73
rect 257 -74 258 -73
rect 324 -74 325 -73
rect 93 -76 94 -75
rect 226 -76 227 -75
rect 229 -76 230 -75
rect 317 -76 318 -75
rect 96 -78 97 -77
rect 100 -78 101 -77
rect 103 -78 104 -77
rect 114 -78 115 -77
rect 121 -78 122 -77
rect 250 -78 251 -77
rect 254 -78 255 -77
rect 268 -78 269 -77
rect 278 -78 279 -77
rect 352 -78 353 -77
rect 107 -80 108 -79
rect 135 -80 136 -79
rect 205 -80 206 -79
rect 219 -80 220 -79
rect 226 -80 227 -79
rect 289 -80 290 -79
rect 296 -80 297 -79
rect 338 -80 339 -79
rect 128 -82 129 -81
rect 191 -82 192 -81
rect 205 -82 206 -81
rect 268 -82 269 -81
rect 212 -84 213 -83
rect 236 -84 237 -83
rect 261 -84 262 -83
rect 296 -84 297 -83
rect 208 -86 209 -85
rect 261 -86 262 -85
rect 233 -88 234 -87
rect 240 -88 241 -87
rect 58 -99 59 -98
rect 170 -99 171 -98
rect 173 -99 174 -98
rect 261 -99 262 -98
rect 352 -99 353 -98
rect 380 -99 381 -98
rect 65 -101 66 -100
rect 180 -101 181 -100
rect 184 -101 185 -100
rect 212 -101 213 -100
rect 236 -101 237 -100
rect 282 -101 283 -100
rect 366 -101 367 -100
rect 373 -101 374 -100
rect 376 -101 377 -100
rect 401 -101 402 -100
rect 72 -103 73 -102
rect 103 -103 104 -102
rect 107 -103 108 -102
rect 201 -103 202 -102
rect 205 -103 206 -102
rect 219 -103 220 -102
rect 243 -103 244 -102
rect 338 -103 339 -102
rect 100 -105 101 -104
rect 114 -105 115 -104
rect 135 -105 136 -104
rect 180 -105 181 -104
rect 187 -105 188 -104
rect 303 -105 304 -104
rect 324 -105 325 -104
rect 366 -105 367 -104
rect 107 -107 108 -106
rect 121 -107 122 -106
rect 145 -107 146 -106
rect 194 -107 195 -106
rect 198 -107 199 -106
rect 271 -107 272 -106
rect 338 -107 339 -106
rect 394 -107 395 -106
rect 86 -109 87 -108
rect 121 -109 122 -108
rect 142 -109 143 -108
rect 145 -109 146 -108
rect 149 -109 150 -108
rect 226 -109 227 -108
rect 236 -109 237 -108
rect 324 -109 325 -108
rect 79 -111 80 -110
rect 142 -111 143 -110
rect 149 -111 150 -110
rect 156 -111 157 -110
rect 163 -111 164 -110
rect 212 -111 213 -110
rect 247 -111 248 -110
rect 296 -111 297 -110
rect 93 -113 94 -112
rect 156 -113 157 -112
rect 163 -113 164 -112
rect 240 -113 241 -112
rect 250 -113 251 -112
rect 296 -113 297 -112
rect 93 -115 94 -114
rect 128 -115 129 -114
rect 177 -115 178 -114
rect 226 -115 227 -114
rect 254 -115 255 -114
rect 317 -115 318 -114
rect 128 -117 129 -116
rect 170 -117 171 -116
rect 191 -117 192 -116
rect 310 -117 311 -116
rect 317 -117 318 -116
rect 331 -117 332 -116
rect 191 -119 192 -118
rect 275 -119 276 -118
rect 310 -119 311 -118
rect 331 -119 332 -118
rect 194 -121 195 -120
rect 240 -121 241 -120
rect 254 -121 255 -120
rect 264 -121 265 -120
rect 205 -123 206 -122
rect 275 -123 276 -122
rect 208 -125 209 -124
rect 261 -125 262 -124
rect 208 -127 209 -126
rect 268 -127 269 -126
rect 219 -129 220 -128
rect 250 -129 251 -128
rect 257 -129 258 -128
rect 289 -129 290 -128
rect 289 -131 290 -130
rect 303 -131 304 -130
rect 65 -142 66 -141
rect 184 -142 185 -141
rect 191 -142 192 -141
rect 341 -142 342 -141
rect 380 -142 381 -141
rect 408 -142 409 -141
rect 93 -144 94 -143
rect 124 -144 125 -143
rect 142 -144 143 -143
rect 156 -144 157 -143
rect 170 -144 171 -143
rect 240 -144 241 -143
rect 243 -144 244 -143
rect 415 -144 416 -143
rect 93 -146 94 -145
rect 117 -146 118 -145
rect 121 -146 122 -145
rect 149 -146 150 -145
rect 163 -146 164 -145
rect 170 -146 171 -145
rect 184 -146 185 -145
rect 236 -146 237 -145
rect 264 -146 265 -145
rect 352 -146 353 -145
rect 380 -146 381 -145
rect 387 -146 388 -145
rect 401 -146 402 -145
rect 429 -146 430 -145
rect 72 -148 73 -147
rect 149 -148 150 -147
rect 152 -148 153 -147
rect 163 -148 164 -147
rect 205 -148 206 -147
rect 212 -148 213 -147
rect 226 -148 227 -147
rect 261 -148 262 -147
rect 289 -148 290 -147
rect 422 -148 423 -147
rect 86 -150 87 -149
rect 117 -150 118 -149
rect 177 -150 178 -149
rect 212 -150 213 -149
rect 233 -150 234 -149
rect 254 -150 255 -149
rect 289 -150 290 -149
rect 296 -150 297 -149
rect 310 -150 311 -149
rect 317 -150 318 -149
rect 331 -150 332 -149
rect 359 -150 360 -149
rect 394 -150 395 -149
rect 401 -150 402 -149
rect 86 -152 87 -151
rect 128 -152 129 -151
rect 229 -152 230 -151
rect 254 -152 255 -151
rect 285 -152 286 -151
rect 296 -152 297 -151
rect 317 -152 318 -151
rect 373 -152 374 -151
rect 107 -154 108 -153
rect 173 -154 174 -153
rect 331 -154 332 -153
rect 355 -154 356 -153
rect 366 -154 367 -153
rect 394 -154 395 -153
rect 107 -156 108 -155
rect 135 -156 136 -155
rect 142 -156 143 -155
rect 229 -156 230 -155
rect 324 -156 325 -155
rect 366 -156 367 -155
rect 100 -158 101 -157
rect 135 -158 136 -157
rect 219 -158 220 -157
rect 324 -158 325 -157
rect 341 -158 342 -157
rect 345 -158 346 -157
rect 100 -160 101 -159
rect 198 -160 199 -159
rect 303 -160 304 -159
rect 345 -160 346 -159
rect 128 -162 129 -161
rect 205 -162 206 -161
rect 247 -162 248 -161
rect 303 -162 304 -161
rect 198 -164 199 -163
rect 268 -164 269 -163
rect 247 -166 248 -165
rect 282 -166 283 -165
rect 23 -177 24 -176
rect 68 -177 69 -176
rect 72 -177 73 -176
rect 201 -177 202 -176
rect 205 -177 206 -176
rect 208 -177 209 -176
rect 219 -177 220 -176
rect 303 -177 304 -176
rect 313 -177 314 -176
rect 352 -177 353 -176
rect 387 -177 388 -176
rect 408 -177 409 -176
rect 411 -177 412 -176
rect 436 -177 437 -176
rect 37 -179 38 -178
rect 243 -179 244 -178
rect 285 -179 286 -178
rect 331 -179 332 -178
rect 341 -179 342 -178
rect 457 -179 458 -178
rect 44 -181 45 -180
rect 79 -181 80 -180
rect 82 -181 83 -180
rect 131 -181 132 -180
rect 149 -181 150 -180
rect 156 -181 157 -180
rect 170 -181 171 -180
rect 180 -181 181 -180
rect 191 -181 192 -180
rect 219 -181 220 -180
rect 236 -181 237 -180
rect 271 -181 272 -180
rect 296 -181 297 -180
rect 310 -181 311 -180
rect 317 -181 318 -180
rect 464 -181 465 -180
rect 51 -183 52 -182
rect 107 -183 108 -182
rect 128 -183 129 -182
rect 194 -183 195 -182
rect 198 -183 199 -182
rect 233 -183 234 -182
rect 240 -183 241 -182
rect 289 -183 290 -182
rect 303 -183 304 -182
rect 324 -183 325 -182
rect 352 -183 353 -182
rect 366 -183 367 -182
rect 380 -183 381 -182
rect 387 -183 388 -182
rect 394 -183 395 -182
rect 429 -183 430 -182
rect 65 -185 66 -184
rect 226 -185 227 -184
rect 243 -185 244 -184
rect 380 -185 381 -184
rect 401 -185 402 -184
rect 439 -185 440 -184
rect 72 -187 73 -186
rect 79 -187 80 -186
rect 86 -187 87 -186
rect 152 -187 153 -186
rect 156 -187 157 -186
rect 222 -187 223 -186
rect 247 -187 248 -186
rect 331 -187 332 -186
rect 359 -187 360 -186
rect 401 -187 402 -186
rect 415 -187 416 -186
rect 443 -187 444 -186
rect 65 -189 66 -188
rect 86 -189 87 -188
rect 93 -189 94 -188
rect 142 -189 143 -188
rect 177 -189 178 -188
rect 215 -189 216 -188
rect 268 -189 269 -188
rect 341 -189 342 -188
rect 373 -189 374 -188
rect 394 -189 395 -188
rect 415 -189 416 -188
rect 432 -189 433 -188
rect 100 -191 101 -190
rect 233 -191 234 -190
rect 275 -191 276 -190
rect 317 -191 318 -190
rect 320 -191 321 -190
rect 366 -191 367 -190
rect 422 -191 423 -190
rect 450 -191 451 -190
rect 96 -193 97 -192
rect 100 -193 101 -192
rect 107 -193 108 -192
rect 163 -193 164 -192
rect 191 -193 192 -192
rect 247 -193 248 -192
rect 268 -193 269 -192
rect 422 -193 423 -192
rect 121 -195 122 -194
rect 142 -195 143 -194
rect 159 -195 160 -194
rect 275 -195 276 -194
rect 285 -195 286 -194
rect 289 -195 290 -194
rect 324 -195 325 -194
rect 359 -195 360 -194
rect 121 -197 122 -196
rect 135 -197 136 -196
rect 138 -197 139 -196
rect 170 -197 171 -196
rect 198 -197 199 -196
rect 212 -197 213 -196
rect 135 -199 136 -198
rect 145 -199 146 -198
rect 163 -199 164 -198
rect 296 -199 297 -198
rect 30 -201 31 -200
rect 145 -201 146 -200
rect 205 -201 206 -200
rect 345 -201 346 -200
rect 254 -203 255 -202
rect 345 -203 346 -202
rect 208 -205 209 -204
rect 254 -205 255 -204
rect 23 -216 24 -215
rect 72 -216 73 -215
rect 100 -216 101 -215
rect 110 -216 111 -215
rect 152 -216 153 -215
rect 450 -216 451 -215
rect 457 -216 458 -215
rect 499 -216 500 -215
rect 541 -216 542 -215
rect 544 -216 545 -215
rect 30 -218 31 -217
rect 205 -218 206 -217
rect 215 -218 216 -217
rect 348 -218 349 -217
rect 408 -218 409 -217
rect 478 -218 479 -217
rect 485 -218 486 -217
rect 537 -218 538 -217
rect 37 -220 38 -219
rect 124 -220 125 -219
rect 156 -220 157 -219
rect 177 -220 178 -219
rect 184 -220 185 -219
rect 212 -220 213 -219
rect 226 -220 227 -219
rect 268 -220 269 -219
rect 271 -220 272 -219
rect 401 -220 402 -219
rect 436 -220 437 -219
rect 471 -220 472 -219
rect 37 -222 38 -221
rect 145 -222 146 -221
rect 149 -222 150 -221
rect 184 -222 185 -221
rect 191 -222 192 -221
rect 303 -222 304 -221
rect 317 -222 318 -221
rect 341 -222 342 -221
rect 345 -222 346 -221
rect 506 -222 507 -221
rect 44 -224 45 -223
rect 58 -224 59 -223
rect 65 -224 66 -223
rect 79 -224 80 -223
rect 100 -224 101 -223
rect 114 -224 115 -223
rect 142 -224 143 -223
rect 177 -224 178 -223
rect 229 -224 230 -223
rect 387 -224 388 -223
rect 429 -224 430 -223
rect 436 -224 437 -223
rect 450 -224 451 -223
rect 534 -224 535 -223
rect 44 -226 45 -225
rect 93 -226 94 -225
rect 107 -226 108 -225
rect 243 -226 244 -225
rect 261 -226 262 -225
rect 296 -226 297 -225
rect 299 -226 300 -225
rect 366 -226 367 -225
rect 464 -226 465 -225
rect 513 -226 514 -225
rect 51 -228 52 -227
rect 138 -228 139 -227
rect 159 -228 160 -227
rect 233 -228 234 -227
rect 236 -228 237 -227
rect 268 -228 269 -227
rect 275 -228 276 -227
rect 324 -228 325 -227
rect 327 -228 328 -227
rect 408 -228 409 -227
rect 443 -228 444 -227
rect 464 -228 465 -227
rect 58 -230 59 -229
rect 226 -230 227 -229
rect 240 -230 241 -229
rect 254 -230 255 -229
rect 275 -230 276 -229
rect 331 -230 332 -229
rect 338 -230 339 -229
rect 520 -230 521 -229
rect 65 -232 66 -231
rect 128 -232 129 -231
rect 163 -232 164 -231
rect 201 -232 202 -231
rect 205 -232 206 -231
rect 261 -232 262 -231
rect 285 -232 286 -231
rect 373 -232 374 -231
rect 51 -234 52 -233
rect 201 -234 202 -233
rect 219 -234 220 -233
rect 254 -234 255 -233
rect 306 -234 307 -233
rect 387 -234 388 -233
rect 79 -236 80 -235
rect 135 -236 136 -235
rect 142 -236 143 -235
rect 219 -236 220 -235
rect 310 -236 311 -235
rect 317 -236 318 -235
rect 331 -236 332 -235
rect 492 -236 493 -235
rect 86 -238 87 -237
rect 163 -238 164 -237
rect 166 -238 167 -237
rect 191 -238 192 -237
rect 198 -238 199 -237
rect 240 -238 241 -237
rect 289 -238 290 -237
rect 310 -238 311 -237
rect 338 -238 339 -237
rect 457 -238 458 -237
rect 93 -240 94 -239
rect 121 -240 122 -239
rect 135 -240 136 -239
rect 180 -240 181 -239
rect 352 -240 353 -239
rect 401 -240 402 -239
rect 89 -242 90 -241
rect 121 -242 122 -241
rect 170 -242 171 -241
rect 208 -242 209 -241
rect 355 -242 356 -241
rect 429 -242 430 -241
rect 170 -244 171 -243
rect 289 -244 290 -243
rect 366 -244 367 -243
rect 394 -244 395 -243
rect 208 -246 209 -245
rect 359 -246 360 -245
rect 394 -246 395 -245
rect 415 -246 416 -245
rect 243 -248 244 -247
rect 359 -248 360 -247
rect 282 -250 283 -249
rect 415 -250 416 -249
rect 282 -252 283 -251
rect 443 -252 444 -251
rect 37 -263 38 -262
rect 229 -263 230 -262
rect 240 -263 241 -262
rect 268 -263 269 -262
rect 282 -263 283 -262
rect 401 -263 402 -262
rect 443 -263 444 -262
rect 555 -263 556 -262
rect 562 -263 563 -262
rect 576 -263 577 -262
rect 37 -265 38 -264
rect 107 -265 108 -264
rect 142 -265 143 -264
rect 212 -265 213 -264
rect 285 -265 286 -264
rect 296 -265 297 -264
rect 303 -265 304 -264
rect 317 -265 318 -264
rect 320 -265 321 -264
rect 506 -265 507 -264
rect 527 -265 528 -264
rect 534 -265 535 -264
rect 44 -267 45 -266
rect 117 -267 118 -266
rect 152 -267 153 -266
rect 233 -267 234 -266
rect 296 -267 297 -266
rect 422 -267 423 -266
rect 464 -267 465 -266
rect 506 -267 507 -266
rect 65 -269 66 -268
rect 131 -269 132 -268
rect 163 -269 164 -268
rect 219 -269 220 -268
rect 306 -269 307 -268
rect 520 -269 521 -268
rect 65 -271 66 -270
rect 114 -271 115 -270
rect 145 -271 146 -270
rect 219 -271 220 -270
rect 324 -271 325 -270
rect 380 -271 381 -270
rect 383 -271 384 -270
rect 548 -271 549 -270
rect 75 -273 76 -272
rect 149 -273 150 -272
rect 170 -273 171 -272
rect 191 -273 192 -272
rect 198 -273 199 -272
rect 289 -273 290 -272
rect 331 -273 332 -272
rect 366 -273 367 -272
rect 408 -273 409 -272
rect 527 -273 528 -272
rect 86 -275 87 -274
rect 128 -275 129 -274
rect 149 -275 150 -274
rect 226 -275 227 -274
rect 289 -275 290 -274
rect 387 -275 388 -274
rect 408 -275 409 -274
rect 415 -275 416 -274
rect 422 -275 423 -274
rect 429 -275 430 -274
rect 499 -275 500 -274
rect 534 -275 535 -274
rect 86 -277 87 -276
rect 114 -277 115 -276
rect 173 -277 174 -276
rect 212 -277 213 -276
rect 226 -277 227 -276
rect 261 -277 262 -276
rect 334 -277 335 -276
rect 478 -277 479 -276
rect 520 -277 521 -276
rect 541 -277 542 -276
rect 79 -279 80 -278
rect 261 -279 262 -278
rect 338 -279 339 -278
rect 387 -279 388 -278
rect 394 -279 395 -278
rect 499 -279 500 -278
rect 93 -281 94 -280
rect 128 -281 129 -280
rect 191 -281 192 -280
rect 268 -281 269 -280
rect 345 -281 346 -280
rect 513 -281 514 -280
rect 96 -283 97 -282
rect 117 -283 118 -282
rect 208 -283 209 -282
rect 275 -283 276 -282
rect 317 -283 318 -282
rect 513 -283 514 -282
rect 100 -285 101 -284
rect 121 -285 122 -284
rect 275 -285 276 -284
rect 359 -285 360 -284
rect 362 -285 363 -284
rect 366 -285 367 -284
rect 415 -285 416 -284
rect 450 -285 451 -284
rect 471 -285 472 -284
rect 478 -285 479 -284
rect 51 -287 52 -286
rect 100 -287 101 -286
rect 107 -287 108 -286
rect 135 -287 136 -286
rect 243 -287 244 -286
rect 450 -287 451 -286
rect 457 -287 458 -286
rect 471 -287 472 -286
rect 51 -289 52 -288
rect 72 -289 73 -288
rect 135 -289 136 -288
rect 166 -289 167 -288
rect 205 -289 206 -288
rect 457 -289 458 -288
rect 72 -291 73 -290
rect 177 -291 178 -290
rect 184 -291 185 -290
rect 205 -291 206 -290
rect 348 -291 349 -290
rect 394 -291 395 -290
rect 429 -291 430 -290
rect 436 -291 437 -290
rect 443 -291 444 -290
rect 541 -291 542 -290
rect 58 -293 59 -292
rect 184 -293 185 -292
rect 303 -293 304 -292
rect 436 -293 437 -292
rect 177 -295 178 -294
rect 247 -295 248 -294
rect 352 -295 353 -294
rect 401 -295 402 -294
rect 247 -297 248 -296
rect 254 -297 255 -296
rect 334 -297 335 -296
rect 352 -297 353 -296
rect 79 -299 80 -298
rect 254 -299 255 -298
rect 9 -310 10 -309
rect 86 -310 87 -309
rect 93 -310 94 -309
rect 149 -310 150 -309
rect 177 -310 178 -309
rect 303 -310 304 -309
rect 334 -310 335 -309
rect 345 -310 346 -309
rect 366 -310 367 -309
rect 478 -310 479 -309
rect 520 -310 521 -309
rect 544 -310 545 -309
rect 548 -310 549 -309
rect 562 -310 563 -309
rect 16 -312 17 -311
rect 275 -312 276 -311
rect 285 -312 286 -311
rect 310 -312 311 -311
rect 334 -312 335 -311
rect 576 -312 577 -311
rect 23 -314 24 -313
rect 96 -314 97 -313
rect 100 -314 101 -313
rect 313 -314 314 -313
rect 338 -314 339 -313
rect 457 -314 458 -313
rect 464 -314 465 -313
rect 492 -314 493 -313
rect 527 -314 528 -313
rect 548 -314 549 -313
rect 30 -316 31 -315
rect 44 -316 45 -315
rect 51 -316 52 -315
rect 61 -316 62 -315
rect 65 -316 66 -315
rect 247 -316 248 -315
rect 250 -316 251 -315
rect 457 -316 458 -315
rect 471 -316 472 -315
rect 555 -316 556 -315
rect 37 -318 38 -317
rect 208 -318 209 -317
rect 240 -318 241 -317
rect 268 -318 269 -317
rect 285 -318 286 -317
rect 576 -318 577 -317
rect 44 -320 45 -319
rect 233 -320 234 -319
rect 240 -320 241 -319
rect 422 -320 423 -319
rect 429 -320 430 -319
rect 527 -320 528 -319
rect 51 -322 52 -321
rect 135 -322 136 -321
rect 180 -322 181 -321
rect 275 -322 276 -321
rect 296 -322 297 -321
rect 429 -322 430 -321
rect 450 -322 451 -321
rect 569 -322 570 -321
rect 61 -324 62 -323
rect 138 -324 139 -323
rect 184 -324 185 -323
rect 247 -324 248 -323
rect 254 -324 255 -323
rect 355 -324 356 -323
rect 373 -324 374 -323
rect 422 -324 423 -323
rect 471 -324 472 -323
rect 513 -324 514 -323
rect 65 -326 66 -325
rect 72 -326 73 -325
rect 79 -326 80 -325
rect 198 -326 199 -325
rect 226 -326 227 -325
rect 254 -326 255 -325
rect 268 -326 269 -325
rect 324 -326 325 -325
rect 348 -326 349 -325
rect 520 -326 521 -325
rect 72 -328 73 -327
rect 142 -328 143 -327
rect 184 -328 185 -327
rect 205 -328 206 -327
rect 219 -328 220 -327
rect 226 -328 227 -327
rect 282 -328 283 -327
rect 569 -328 570 -327
rect 86 -330 87 -329
rect 170 -330 171 -329
rect 194 -330 195 -329
rect 212 -330 213 -329
rect 219 -330 220 -329
rect 261 -330 262 -329
rect 299 -330 300 -329
rect 513 -330 514 -329
rect 103 -332 104 -331
rect 233 -332 234 -331
rect 261 -332 262 -331
rect 296 -332 297 -331
rect 310 -332 311 -331
rect 450 -332 451 -331
rect 107 -334 108 -333
rect 131 -334 132 -333
rect 142 -334 143 -333
rect 338 -334 339 -333
rect 348 -334 349 -333
rect 541 -334 542 -333
rect 114 -336 115 -335
rect 408 -336 409 -335
rect 534 -336 535 -335
rect 541 -336 542 -335
rect 114 -338 115 -337
rect 121 -338 122 -337
rect 149 -338 150 -337
rect 170 -338 171 -337
rect 194 -338 195 -337
rect 303 -338 304 -337
rect 317 -338 318 -337
rect 492 -338 493 -337
rect 121 -340 122 -339
rect 191 -340 192 -339
rect 198 -340 199 -339
rect 282 -340 283 -339
rect 317 -340 318 -339
rect 331 -340 332 -339
rect 345 -340 346 -339
rect 534 -340 535 -339
rect 163 -342 164 -341
rect 212 -342 213 -341
rect 352 -342 353 -341
rect 408 -342 409 -341
rect 156 -344 157 -343
rect 163 -344 164 -343
rect 352 -344 353 -343
rect 478 -344 479 -343
rect 156 -346 157 -345
rect 359 -346 360 -345
rect 373 -346 374 -345
rect 401 -346 402 -345
rect 380 -348 381 -347
rect 506 -348 507 -347
rect 383 -350 384 -349
rect 499 -350 500 -349
rect 387 -352 388 -351
rect 464 -352 465 -351
rect 341 -354 342 -353
rect 387 -354 388 -353
rect 394 -354 395 -353
rect 506 -354 507 -353
rect 271 -356 272 -355
rect 394 -356 395 -355
rect 401 -356 402 -355
rect 415 -356 416 -355
rect 443 -356 444 -355
rect 499 -356 500 -355
rect 292 -358 293 -357
rect 415 -358 416 -357
rect 436 -358 437 -357
rect 443 -358 444 -357
rect 205 -360 206 -359
rect 436 -360 437 -359
rect 2 -371 3 -370
rect 191 -371 192 -370
rect 201 -371 202 -370
rect 331 -371 332 -370
rect 345 -371 346 -370
rect 422 -371 423 -370
rect 513 -371 514 -370
rect 583 -371 584 -370
rect 9 -373 10 -372
rect 135 -373 136 -372
rect 156 -373 157 -372
rect 163 -373 164 -372
rect 184 -373 185 -372
rect 338 -373 339 -372
rect 348 -373 349 -372
rect 394 -373 395 -372
rect 422 -373 423 -372
rect 478 -373 479 -372
rect 534 -373 535 -372
rect 611 -373 612 -372
rect 16 -375 17 -374
rect 250 -375 251 -374
rect 254 -375 255 -374
rect 285 -375 286 -374
rect 296 -375 297 -374
rect 499 -375 500 -374
rect 555 -375 556 -374
rect 576 -375 577 -374
rect 23 -377 24 -376
rect 149 -377 150 -376
rect 156 -377 157 -376
rect 306 -377 307 -376
rect 313 -377 314 -376
rect 471 -377 472 -376
rect 23 -379 24 -378
rect 33 -379 34 -378
rect 37 -379 38 -378
rect 61 -379 62 -378
rect 65 -379 66 -378
rect 177 -379 178 -378
rect 219 -379 220 -378
rect 327 -379 328 -378
rect 352 -379 353 -378
rect 523 -379 524 -378
rect 30 -381 31 -380
rect 58 -381 59 -380
rect 68 -381 69 -380
rect 177 -381 178 -380
rect 226 -381 227 -380
rect 282 -381 283 -380
rect 296 -381 297 -380
rect 317 -381 318 -380
rect 355 -381 356 -380
rect 548 -381 549 -380
rect 37 -383 38 -382
rect 124 -383 125 -382
rect 149 -383 150 -382
rect 163 -383 164 -382
rect 170 -383 171 -382
rect 184 -383 185 -382
rect 299 -383 300 -382
rect 408 -383 409 -382
rect 443 -383 444 -382
rect 499 -383 500 -382
rect 44 -385 45 -384
rect 271 -385 272 -384
rect 303 -385 304 -384
rect 310 -385 311 -384
rect 366 -385 367 -384
rect 464 -385 465 -384
rect 471 -385 472 -384
rect 520 -385 521 -384
rect 44 -387 45 -386
rect 107 -387 108 -386
rect 121 -387 122 -386
rect 261 -387 262 -386
rect 268 -387 269 -386
rect 366 -387 367 -386
rect 380 -387 381 -386
rect 548 -387 549 -386
rect 51 -389 52 -388
rect 219 -389 220 -388
rect 233 -389 234 -388
rect 261 -389 262 -388
rect 320 -389 321 -388
rect 464 -389 465 -388
rect 51 -391 52 -390
rect 103 -391 104 -390
rect 107 -391 108 -390
rect 114 -391 115 -390
rect 170 -391 171 -390
rect 212 -391 213 -390
rect 233 -391 234 -390
rect 275 -391 276 -390
rect 380 -391 381 -390
rect 527 -391 528 -390
rect 58 -393 59 -392
rect 205 -393 206 -392
rect 212 -393 213 -392
rect 327 -393 328 -392
rect 390 -393 391 -392
rect 576 -393 577 -392
rect 72 -395 73 -394
rect 152 -395 153 -394
rect 191 -395 192 -394
rect 275 -395 276 -394
rect 394 -395 395 -394
rect 401 -395 402 -394
rect 408 -395 409 -394
rect 415 -395 416 -394
rect 443 -395 444 -394
rect 492 -395 493 -394
rect 527 -395 528 -394
rect 569 -395 570 -394
rect 72 -397 73 -396
rect 96 -397 97 -396
rect 100 -397 101 -396
rect 226 -397 227 -396
rect 373 -397 374 -396
rect 401 -397 402 -396
rect 415 -397 416 -396
rect 506 -397 507 -396
rect 558 -397 559 -396
rect 569 -397 570 -396
rect 79 -399 80 -398
rect 208 -399 209 -398
rect 348 -399 349 -398
rect 373 -399 374 -398
rect 387 -399 388 -398
rect 492 -399 493 -398
rect 79 -401 80 -400
rect 142 -401 143 -400
rect 152 -401 153 -400
rect 429 -401 430 -400
rect 450 -401 451 -400
rect 534 -401 535 -400
rect 86 -403 87 -402
rect 243 -403 244 -402
rect 383 -403 384 -402
rect 450 -403 451 -402
rect 457 -403 458 -402
rect 478 -403 479 -402
rect 93 -405 94 -404
rect 131 -405 132 -404
rect 138 -405 139 -404
rect 387 -405 388 -404
rect 411 -405 412 -404
rect 506 -405 507 -404
rect 9 -407 10 -406
rect 138 -407 139 -406
rect 142 -407 143 -406
rect 198 -407 199 -406
rect 243 -407 244 -406
rect 247 -407 248 -406
rect 429 -407 430 -406
rect 541 -407 542 -406
rect 114 -409 115 -408
rect 128 -409 129 -408
rect 247 -409 248 -408
rect 513 -409 514 -408
rect 541 -409 542 -408
rect 562 -409 563 -408
rect 359 -411 360 -410
rect 562 -411 563 -410
rect 436 -413 437 -412
rect 457 -413 458 -412
rect 324 -415 325 -414
rect 436 -415 437 -414
rect 2 -426 3 -425
rect 156 -426 157 -425
rect 198 -426 199 -425
rect 219 -426 220 -425
rect 240 -426 241 -425
rect 520 -426 521 -425
rect 576 -426 577 -425
rect 597 -426 598 -425
rect 611 -426 612 -425
rect 639 -426 640 -425
rect 663 -426 664 -425
rect 674 -426 675 -425
rect 2 -428 3 -427
rect 51 -428 52 -427
rect 79 -428 80 -427
rect 187 -428 188 -427
rect 208 -428 209 -427
rect 352 -428 353 -427
rect 355 -428 356 -427
rect 394 -428 395 -427
rect 464 -428 465 -427
rect 625 -428 626 -427
rect 635 -428 636 -427
rect 667 -428 668 -427
rect 9 -430 10 -429
rect 72 -430 73 -429
rect 79 -430 80 -429
rect 177 -430 178 -429
rect 257 -430 258 -429
rect 338 -430 339 -429
rect 348 -430 349 -429
rect 471 -430 472 -429
rect 506 -430 507 -429
rect 590 -430 591 -429
rect 16 -432 17 -431
rect 114 -432 115 -431
rect 128 -432 129 -431
rect 159 -432 160 -431
rect 170 -432 171 -431
rect 219 -432 220 -431
rect 271 -432 272 -431
rect 282 -432 283 -431
rect 310 -432 311 -431
rect 383 -432 384 -431
rect 422 -432 423 -431
rect 506 -432 507 -431
rect 513 -432 514 -431
rect 576 -432 577 -431
rect 583 -432 584 -431
rect 604 -432 605 -431
rect 19 -434 20 -433
rect 247 -434 248 -433
rect 275 -434 276 -433
rect 289 -434 290 -433
rect 313 -434 314 -433
rect 415 -434 416 -433
rect 436 -434 437 -433
rect 583 -434 584 -433
rect 30 -436 31 -435
rect 40 -436 41 -435
rect 44 -436 45 -435
rect 205 -436 206 -435
rect 226 -436 227 -435
rect 415 -436 416 -435
rect 492 -436 493 -435
rect 513 -436 514 -435
rect 527 -436 528 -435
rect 611 -436 612 -435
rect 44 -438 45 -437
rect 621 -438 622 -437
rect 47 -440 48 -439
rect 212 -440 213 -439
rect 233 -440 234 -439
rect 289 -440 290 -439
rect 317 -440 318 -439
rect 548 -440 549 -439
rect 51 -442 52 -441
rect 359 -442 360 -441
rect 362 -442 363 -441
rect 555 -442 556 -441
rect 68 -444 69 -443
rect 338 -444 339 -443
rect 373 -444 374 -443
rect 387 -444 388 -443
rect 401 -444 402 -443
rect 436 -444 437 -443
rect 457 -444 458 -443
rect 548 -444 549 -443
rect 72 -446 73 -445
rect 261 -446 262 -445
rect 275 -446 276 -445
rect 397 -446 398 -445
rect 478 -446 479 -445
rect 555 -446 556 -445
rect 86 -448 87 -447
rect 173 -448 174 -447
rect 177 -448 178 -447
rect 191 -448 192 -447
rect 278 -448 279 -447
rect 296 -448 297 -447
rect 303 -448 304 -447
rect 457 -448 458 -447
rect 499 -448 500 -447
rect 527 -448 528 -447
rect 86 -450 87 -449
rect 243 -450 244 -449
rect 282 -450 283 -449
rect 362 -450 363 -449
rect 380 -450 381 -449
rect 429 -450 430 -449
rect 93 -452 94 -451
rect 464 -452 465 -451
rect 93 -454 94 -453
rect 114 -454 115 -453
rect 121 -454 122 -453
rect 212 -454 213 -453
rect 243 -454 244 -453
rect 373 -454 374 -453
rect 429 -454 430 -453
rect 562 -454 563 -453
rect 96 -456 97 -455
rect 117 -456 118 -455
rect 138 -456 139 -455
rect 250 -456 251 -455
rect 296 -456 297 -455
rect 394 -456 395 -455
rect 534 -456 535 -455
rect 562 -456 563 -455
rect 100 -458 101 -457
rect 184 -458 185 -457
rect 191 -458 192 -457
rect 345 -458 346 -457
rect 145 -460 146 -459
rect 226 -460 227 -459
rect 254 -460 255 -459
rect 534 -460 535 -459
rect 149 -462 150 -461
rect 163 -462 164 -461
rect 170 -462 171 -461
rect 401 -462 402 -461
rect 58 -464 59 -463
rect 163 -464 164 -463
rect 254 -464 255 -463
rect 264 -464 265 -463
rect 310 -464 311 -463
rect 478 -464 479 -463
rect 58 -466 59 -465
rect 131 -466 132 -465
rect 156 -466 157 -465
rect 233 -466 234 -465
rect 317 -466 318 -465
rect 352 -466 353 -465
rect 37 -468 38 -467
rect 131 -468 132 -467
rect 320 -468 321 -467
rect 366 -468 367 -467
rect 23 -470 24 -469
rect 37 -470 38 -469
rect 201 -470 202 -469
rect 366 -470 367 -469
rect 23 -472 24 -471
rect 142 -472 143 -471
rect 324 -472 325 -471
rect 471 -472 472 -471
rect 135 -474 136 -473
rect 142 -474 143 -473
rect 324 -474 325 -473
rect 499 -474 500 -473
rect 107 -476 108 -475
rect 135 -476 136 -475
rect 327 -476 328 -475
rect 443 -476 444 -475
rect 107 -478 108 -477
rect 138 -478 139 -477
rect 327 -478 328 -477
rect 646 -478 647 -477
rect 124 -480 125 -479
rect 443 -480 444 -479
rect 331 -482 332 -481
rect 408 -482 409 -481
rect 331 -484 332 -483
rect 541 -484 542 -483
rect 334 -486 335 -485
rect 380 -486 381 -485
rect 450 -486 451 -485
rect 541 -486 542 -485
rect 450 -488 451 -487
rect 569 -488 570 -487
rect 485 -490 486 -489
rect 569 -490 570 -489
rect 422 -492 423 -491
rect 485 -492 486 -491
rect 2 -503 3 -502
rect 47 -503 48 -502
rect 51 -503 52 -502
rect 124 -503 125 -502
rect 128 -503 129 -502
rect 212 -503 213 -502
rect 236 -503 237 -502
rect 457 -503 458 -502
rect 492 -503 493 -502
rect 562 -503 563 -502
rect 597 -503 598 -502
rect 628 -503 629 -502
rect 635 -503 636 -502
rect 674 -503 675 -502
rect 9 -505 10 -504
rect 173 -505 174 -504
rect 205 -505 206 -504
rect 415 -505 416 -504
rect 422 -505 423 -504
rect 464 -505 465 -504
rect 492 -505 493 -504
rect 569 -505 570 -504
rect 597 -505 598 -504
rect 646 -505 647 -504
rect 16 -507 17 -506
rect 191 -507 192 -506
rect 208 -507 209 -506
rect 219 -507 220 -506
rect 240 -507 241 -506
rect 443 -507 444 -506
rect 464 -507 465 -506
rect 548 -507 549 -506
rect 604 -507 605 -506
rect 614 -507 615 -506
rect 618 -507 619 -506
rect 667 -507 668 -506
rect 16 -509 17 -508
rect 75 -509 76 -508
rect 79 -509 80 -508
rect 264 -509 265 -508
rect 289 -509 290 -508
rect 306 -509 307 -508
rect 310 -509 311 -508
rect 415 -509 416 -508
rect 513 -509 514 -508
rect 604 -509 605 -508
rect 639 -509 640 -508
rect 646 -509 647 -508
rect 23 -511 24 -510
rect 198 -511 199 -510
rect 212 -511 213 -510
rect 334 -511 335 -510
rect 345 -511 346 -510
rect 548 -511 549 -510
rect 576 -511 577 -510
rect 618 -511 619 -510
rect 23 -513 24 -512
rect 30 -513 31 -512
rect 37 -513 38 -512
rect 394 -513 395 -512
rect 397 -513 398 -512
rect 527 -513 528 -512
rect 30 -515 31 -514
rect 72 -515 73 -514
rect 86 -515 87 -514
rect 152 -515 153 -514
rect 170 -515 171 -514
rect 506 -515 507 -514
rect 513 -515 514 -514
rect 555 -515 556 -514
rect 51 -517 52 -516
rect 331 -517 332 -516
rect 334 -517 335 -516
rect 569 -517 570 -516
rect 58 -519 59 -518
rect 208 -519 209 -518
rect 303 -519 304 -518
rect 499 -519 500 -518
rect 527 -519 528 -518
rect 653 -519 654 -518
rect 86 -521 87 -520
rect 282 -521 283 -520
rect 310 -521 311 -520
rect 366 -521 367 -520
rect 369 -521 370 -520
rect 499 -521 500 -520
rect 555 -521 556 -520
rect 590 -521 591 -520
rect 621 -521 622 -520
rect 653 -521 654 -520
rect 93 -523 94 -522
rect 114 -523 115 -522
rect 131 -523 132 -522
rect 562 -523 563 -522
rect 590 -523 591 -522
rect 625 -523 626 -522
rect 93 -525 94 -524
rect 278 -525 279 -524
rect 282 -525 283 -524
rect 352 -525 353 -524
rect 355 -525 356 -524
rect 478 -525 479 -524
rect 495 -525 496 -524
rect 506 -525 507 -524
rect 625 -525 626 -524
rect 642 -525 643 -524
rect 100 -527 101 -526
rect 184 -527 185 -526
rect 191 -527 192 -526
rect 226 -527 227 -526
rect 275 -527 276 -526
rect 303 -527 304 -526
rect 324 -527 325 -526
rect 429 -527 430 -526
rect 478 -527 479 -526
rect 534 -527 535 -526
rect 100 -529 101 -528
rect 163 -529 164 -528
rect 170 -529 171 -528
rect 219 -529 220 -528
rect 226 -529 227 -528
rect 268 -529 269 -528
rect 275 -529 276 -528
rect 471 -529 472 -528
rect 485 -529 486 -528
rect 534 -529 535 -528
rect 107 -531 108 -530
rect 289 -531 290 -530
rect 324 -531 325 -530
rect 390 -531 391 -530
rect 397 -531 398 -530
rect 611 -531 612 -530
rect 107 -533 108 -532
rect 149 -533 150 -532
rect 163 -533 164 -532
rect 611 -533 612 -532
rect 65 -535 66 -534
rect 149 -535 150 -534
rect 177 -535 178 -534
rect 240 -535 241 -534
rect 348 -535 349 -534
rect 443 -535 444 -534
rect 457 -535 458 -534
rect 485 -535 486 -534
rect 61 -537 62 -536
rect 177 -537 178 -536
rect 198 -537 199 -536
rect 254 -537 255 -536
rect 362 -537 363 -536
rect 450 -537 451 -536
rect 121 -539 122 -538
rect 131 -539 132 -538
rect 135 -539 136 -538
rect 156 -539 157 -538
rect 205 -539 206 -538
rect 471 -539 472 -538
rect 142 -541 143 -540
rect 233 -541 234 -540
rect 254 -541 255 -540
rect 313 -541 314 -540
rect 366 -541 367 -540
rect 408 -541 409 -540
rect 429 -541 430 -540
rect 520 -541 521 -540
rect 145 -543 146 -542
rect 632 -543 633 -542
rect 156 -545 157 -544
rect 359 -545 360 -544
rect 373 -545 374 -544
rect 411 -545 412 -544
rect 436 -545 437 -544
rect 450 -545 451 -544
rect 520 -545 521 -544
rect 583 -545 584 -544
rect 632 -545 633 -544
rect 639 -545 640 -544
rect 271 -547 272 -546
rect 583 -547 584 -546
rect 338 -549 339 -548
rect 436 -549 437 -548
rect 296 -551 297 -550
rect 338 -551 339 -550
rect 373 -551 374 -550
rect 401 -551 402 -550
rect 296 -553 297 -552
rect 317 -553 318 -552
rect 380 -553 381 -552
rect 425 -553 426 -552
rect 247 -555 248 -554
rect 317 -555 318 -554
rect 380 -555 381 -554
rect 576 -555 577 -554
rect 247 -557 248 -556
rect 268 -557 269 -556
rect 383 -557 384 -556
rect 387 -557 388 -556
rect 2 -568 3 -567
rect 93 -568 94 -567
rect 100 -568 101 -567
rect 142 -568 143 -567
rect 156 -568 157 -567
rect 240 -568 241 -567
rect 254 -568 255 -567
rect 355 -568 356 -567
rect 369 -568 370 -567
rect 464 -568 465 -567
rect 485 -568 486 -567
rect 555 -568 556 -567
rect 576 -568 577 -567
rect 611 -568 612 -567
rect 618 -568 619 -567
rect 628 -568 629 -567
rect 642 -568 643 -567
rect 653 -568 654 -567
rect 9 -570 10 -569
rect 100 -570 101 -569
rect 114 -570 115 -569
rect 149 -570 150 -569
rect 170 -570 171 -569
rect 212 -570 213 -569
rect 233 -570 234 -569
rect 268 -570 269 -569
rect 271 -570 272 -569
rect 317 -570 318 -569
rect 352 -570 353 -569
rect 590 -570 591 -569
rect 646 -570 647 -569
rect 653 -570 654 -569
rect 16 -572 17 -571
rect 103 -572 104 -571
rect 114 -572 115 -571
rect 135 -572 136 -571
rect 142 -572 143 -571
rect 205 -572 206 -571
rect 208 -572 209 -571
rect 229 -572 230 -571
rect 261 -572 262 -571
rect 404 -572 405 -571
rect 408 -572 409 -571
rect 604 -572 605 -571
rect 16 -574 17 -573
rect 310 -574 311 -573
rect 331 -574 332 -573
rect 590 -574 591 -573
rect 23 -576 24 -575
rect 79 -576 80 -575
rect 82 -576 83 -575
rect 93 -576 94 -575
rect 135 -576 136 -575
rect 257 -576 258 -575
rect 268 -576 269 -575
rect 324 -576 325 -575
rect 373 -576 374 -575
rect 576 -576 577 -575
rect 583 -576 584 -575
rect 618 -576 619 -575
rect 23 -578 24 -577
rect 191 -578 192 -577
rect 194 -578 195 -577
rect 226 -578 227 -577
rect 278 -578 279 -577
rect 317 -578 318 -577
rect 324 -578 325 -577
rect 450 -578 451 -577
rect 464 -578 465 -577
rect 471 -578 472 -577
rect 544 -578 545 -577
rect 597 -578 598 -577
rect 30 -580 31 -579
rect 380 -580 381 -579
rect 383 -580 384 -579
rect 411 -580 412 -579
rect 429 -580 430 -579
rect 432 -580 433 -579
rect 450 -580 451 -579
rect 625 -580 626 -579
rect 30 -582 31 -581
rect 72 -582 73 -581
rect 79 -582 80 -581
rect 163 -582 164 -581
rect 170 -582 171 -581
rect 184 -582 185 -581
rect 198 -582 199 -581
rect 201 -582 202 -581
rect 205 -582 206 -581
rect 408 -582 409 -581
rect 429 -582 430 -581
rect 478 -582 479 -581
rect 506 -582 507 -581
rect 597 -582 598 -581
rect 51 -584 52 -583
rect 233 -584 234 -583
rect 303 -584 304 -583
rect 334 -584 335 -583
rect 387 -584 388 -583
rect 520 -584 521 -583
rect 565 -584 566 -583
rect 604 -584 605 -583
rect 51 -586 52 -585
rect 121 -586 122 -585
rect 152 -586 153 -585
rect 163 -586 164 -585
rect 177 -586 178 -585
rect 261 -586 262 -585
rect 296 -586 297 -585
rect 303 -586 304 -585
rect 310 -586 311 -585
rect 436 -586 437 -585
rect 443 -586 444 -585
rect 478 -586 479 -585
rect 506 -586 507 -585
rect 548 -586 549 -585
rect 569 -586 570 -585
rect 583 -586 584 -585
rect 61 -588 62 -587
rect 240 -588 241 -587
rect 264 -588 265 -587
rect 436 -588 437 -587
rect 471 -588 472 -587
rect 499 -588 500 -587
rect 520 -588 521 -587
rect 534 -588 535 -587
rect 548 -588 549 -587
rect 562 -588 563 -587
rect 65 -590 66 -589
rect 296 -590 297 -589
rect 345 -590 346 -589
rect 499 -590 500 -589
rect 527 -590 528 -589
rect 569 -590 570 -589
rect 68 -592 69 -591
rect 128 -592 129 -591
rect 152 -592 153 -591
rect 338 -592 339 -591
rect 394 -592 395 -591
rect 485 -592 486 -591
rect 534 -592 535 -591
rect 541 -592 542 -591
rect 72 -594 73 -593
rect 219 -594 220 -593
rect 226 -594 227 -593
rect 282 -594 283 -593
rect 338 -594 339 -593
rect 362 -594 363 -593
rect 401 -594 402 -593
rect 513 -594 514 -593
rect 58 -596 59 -595
rect 219 -596 220 -595
rect 247 -596 248 -595
rect 394 -596 395 -595
rect 401 -596 402 -595
rect 492 -596 493 -595
rect 86 -598 87 -597
rect 348 -598 349 -597
rect 432 -598 433 -597
rect 443 -598 444 -597
rect 457 -598 458 -597
rect 513 -598 514 -597
rect 86 -600 87 -599
rect 191 -600 192 -599
rect 198 -600 199 -599
rect 555 -600 556 -599
rect 107 -602 108 -601
rect 184 -602 185 -601
rect 212 -602 213 -601
rect 352 -602 353 -601
rect 492 -602 493 -601
rect 621 -602 622 -601
rect 37 -604 38 -603
rect 107 -604 108 -603
rect 121 -604 122 -603
rect 373 -604 374 -603
rect 37 -606 38 -605
rect 44 -606 45 -605
rect 156 -606 157 -605
rect 177 -606 178 -605
rect 180 -606 181 -605
rect 247 -606 248 -605
rect 282 -606 283 -605
rect 415 -606 416 -605
rect 44 -608 45 -607
rect 124 -608 125 -607
rect 348 -608 349 -607
rect 366 -608 367 -607
rect 415 -608 416 -607
rect 422 -608 423 -607
rect 359 -610 360 -609
rect 422 -610 423 -609
rect 359 -612 360 -611
rect 387 -612 388 -611
rect 2 -623 3 -622
rect 128 -623 129 -622
rect 131 -623 132 -622
rect 208 -623 209 -622
rect 212 -623 213 -622
rect 334 -623 335 -622
rect 345 -623 346 -622
rect 569 -623 570 -622
rect 625 -623 626 -622
rect 639 -623 640 -622
rect 2 -625 3 -624
rect 93 -625 94 -624
rect 100 -625 101 -624
rect 152 -625 153 -624
rect 173 -625 174 -624
rect 583 -625 584 -624
rect 9 -627 10 -626
rect 205 -627 206 -626
rect 208 -627 209 -626
rect 604 -627 605 -626
rect 9 -629 10 -628
rect 68 -629 69 -628
rect 103 -629 104 -628
rect 194 -629 195 -628
rect 201 -629 202 -628
rect 261 -629 262 -628
rect 296 -629 297 -628
rect 327 -629 328 -628
rect 334 -629 335 -628
rect 562 -629 563 -628
rect 565 -629 566 -628
rect 590 -629 591 -628
rect 16 -631 17 -630
rect 278 -631 279 -630
rect 289 -631 290 -630
rect 296 -631 297 -630
rect 313 -631 314 -630
rect 429 -631 430 -630
rect 443 -631 444 -630
rect 478 -631 479 -630
rect 513 -631 514 -630
rect 541 -631 542 -630
rect 16 -633 17 -632
rect 131 -633 132 -632
rect 184 -633 185 -632
rect 359 -633 360 -632
rect 362 -633 363 -632
rect 597 -633 598 -632
rect 23 -635 24 -634
rect 177 -635 178 -634
rect 219 -635 220 -634
rect 331 -635 332 -634
rect 348 -635 349 -634
rect 576 -635 577 -634
rect 23 -637 24 -636
rect 96 -637 97 -636
rect 107 -637 108 -636
rect 110 -637 111 -636
rect 114 -637 115 -636
rect 138 -637 139 -636
rect 170 -637 171 -636
rect 184 -637 185 -636
rect 219 -637 220 -636
rect 401 -637 402 -636
rect 443 -637 444 -636
rect 492 -637 493 -636
rect 520 -637 521 -636
rect 558 -637 559 -636
rect 30 -639 31 -638
rect 152 -639 153 -638
rect 177 -639 178 -638
rect 380 -639 381 -638
rect 429 -639 430 -638
rect 492 -639 493 -638
rect 520 -639 521 -638
rect 548 -639 549 -638
rect 30 -641 31 -640
rect 278 -641 279 -640
rect 324 -641 325 -640
rect 548 -641 549 -640
rect 37 -643 38 -642
rect 65 -643 66 -642
rect 107 -643 108 -642
rect 163 -643 164 -642
rect 222 -643 223 -642
rect 317 -643 318 -642
rect 324 -643 325 -642
rect 404 -643 405 -642
rect 460 -643 461 -642
rect 611 -643 612 -642
rect 37 -645 38 -644
rect 142 -645 143 -644
rect 226 -645 227 -644
rect 387 -645 388 -644
rect 527 -645 528 -644
rect 618 -645 619 -644
rect 44 -647 45 -646
rect 198 -647 199 -646
rect 226 -647 227 -646
rect 247 -647 248 -646
rect 257 -647 258 -646
rect 464 -647 465 -646
rect 44 -649 45 -648
rect 205 -649 206 -648
rect 240 -649 241 -648
rect 289 -649 290 -648
rect 303 -649 304 -648
rect 317 -649 318 -648
rect 338 -649 339 -648
rect 380 -649 381 -648
rect 387 -649 388 -648
rect 394 -649 395 -648
rect 436 -649 437 -648
rect 527 -649 528 -648
rect 51 -651 52 -650
rect 201 -651 202 -650
rect 247 -651 248 -650
rect 457 -651 458 -650
rect 51 -653 52 -652
rect 261 -653 262 -652
rect 275 -653 276 -652
rect 338 -653 339 -652
rect 345 -653 346 -652
rect 404 -653 405 -652
rect 408 -653 409 -652
rect 436 -653 437 -652
rect 58 -655 59 -654
rect 170 -655 171 -654
rect 282 -655 283 -654
rect 303 -655 304 -654
rect 310 -655 311 -654
rect 464 -655 465 -654
rect 61 -657 62 -656
rect 555 -657 556 -656
rect 65 -659 66 -658
rect 229 -659 230 -658
rect 268 -659 269 -658
rect 310 -659 311 -658
rect 313 -659 314 -658
rect 457 -659 458 -658
rect 513 -659 514 -658
rect 555 -659 556 -658
rect 72 -661 73 -660
rect 268 -661 269 -660
rect 352 -661 353 -660
rect 373 -661 374 -660
rect 408 -661 409 -660
rect 450 -661 451 -660
rect 72 -663 73 -662
rect 128 -663 129 -662
rect 135 -663 136 -662
rect 142 -663 143 -662
rect 180 -663 181 -662
rect 450 -663 451 -662
rect 79 -665 80 -664
rect 240 -665 241 -664
rect 355 -665 356 -664
rect 422 -665 423 -664
rect 79 -667 80 -666
rect 135 -667 136 -666
rect 191 -667 192 -666
rect 373 -667 374 -666
rect 422 -667 423 -666
rect 534 -667 535 -666
rect 110 -669 111 -668
rect 163 -669 164 -668
rect 366 -669 367 -668
rect 397 -669 398 -668
rect 506 -669 507 -668
rect 534 -669 535 -668
rect 121 -671 122 -670
rect 233 -671 234 -670
rect 369 -671 370 -670
rect 471 -671 472 -670
rect 485 -671 486 -670
rect 506 -671 507 -670
rect 86 -673 87 -672
rect 233 -673 234 -672
rect 257 -673 258 -672
rect 471 -673 472 -672
rect 86 -675 87 -674
rect 149 -675 150 -674
rect 394 -675 395 -674
rect 485 -675 486 -674
rect 121 -677 122 -676
rect 212 -677 213 -676
rect 2 -688 3 -687
rect 205 -688 206 -687
rect 219 -688 220 -687
rect 285 -688 286 -687
rect 289 -688 290 -687
rect 306 -688 307 -687
rect 313 -688 314 -687
rect 415 -688 416 -687
rect 422 -688 423 -687
rect 425 -688 426 -687
rect 429 -688 430 -687
rect 450 -688 451 -687
rect 457 -688 458 -687
rect 611 -688 612 -687
rect 632 -688 633 -687
rect 639 -688 640 -687
rect 2 -690 3 -689
rect 58 -690 59 -689
rect 96 -690 97 -689
rect 173 -690 174 -689
rect 177 -690 178 -689
rect 254 -690 255 -689
rect 278 -690 279 -689
rect 296 -690 297 -689
rect 331 -690 332 -689
rect 457 -690 458 -689
rect 478 -690 479 -689
rect 583 -690 584 -689
rect 9 -692 10 -691
rect 121 -692 122 -691
rect 135 -692 136 -691
rect 156 -692 157 -691
rect 170 -692 171 -691
rect 191 -692 192 -691
rect 194 -692 195 -691
rect 226 -692 227 -691
rect 229 -692 230 -691
rect 590 -692 591 -691
rect 12 -694 13 -693
rect 394 -694 395 -693
rect 397 -694 398 -693
rect 548 -694 549 -693
rect 562 -694 563 -693
rect 663 -694 664 -693
rect 16 -696 17 -695
rect 117 -696 118 -695
rect 121 -696 122 -695
rect 180 -696 181 -695
rect 187 -696 188 -695
rect 562 -696 563 -695
rect 16 -698 17 -697
rect 93 -698 94 -697
rect 114 -698 115 -697
rect 576 -698 577 -697
rect 30 -700 31 -699
rect 128 -700 129 -699
rect 156 -700 157 -699
rect 212 -700 213 -699
rect 219 -700 220 -699
rect 261 -700 262 -699
rect 271 -700 272 -699
rect 331 -700 332 -699
rect 338 -700 339 -699
rect 597 -700 598 -699
rect 30 -702 31 -701
rect 107 -702 108 -701
rect 114 -702 115 -701
rect 478 -702 479 -701
rect 485 -702 486 -701
rect 569 -702 570 -701
rect 37 -704 38 -703
rect 257 -704 258 -703
rect 278 -704 279 -703
rect 401 -704 402 -703
rect 404 -704 405 -703
rect 555 -704 556 -703
rect 37 -706 38 -705
rect 86 -706 87 -705
rect 117 -706 118 -705
rect 296 -706 297 -705
rect 341 -706 342 -705
rect 443 -706 444 -705
rect 464 -706 465 -705
rect 548 -706 549 -705
rect 44 -708 45 -707
rect 47 -708 48 -707
rect 51 -708 52 -707
rect 261 -708 262 -707
rect 345 -708 346 -707
rect 415 -708 416 -707
rect 432 -708 433 -707
rect 506 -708 507 -707
rect 520 -708 521 -707
rect 618 -708 619 -707
rect 54 -710 55 -709
rect 240 -710 241 -709
rect 247 -710 248 -709
rect 285 -710 286 -709
rect 292 -710 293 -709
rect 506 -710 507 -709
rect 527 -710 528 -709
rect 625 -710 626 -709
rect 82 -712 83 -711
rect 212 -712 213 -711
rect 226 -712 227 -711
rect 471 -712 472 -711
rect 492 -712 493 -711
rect 604 -712 605 -711
rect 86 -714 87 -713
rect 142 -714 143 -713
rect 145 -714 146 -713
rect 527 -714 528 -713
rect 100 -716 101 -715
rect 247 -716 248 -715
rect 254 -716 255 -715
rect 373 -716 374 -715
rect 376 -716 377 -715
rect 541 -716 542 -715
rect 128 -718 129 -717
rect 184 -718 185 -717
rect 198 -718 199 -717
rect 324 -718 325 -717
rect 345 -718 346 -717
rect 366 -718 367 -717
rect 376 -718 377 -717
rect 646 -718 647 -717
rect 107 -720 108 -719
rect 198 -720 199 -719
rect 233 -720 234 -719
rect 369 -720 370 -719
rect 380 -720 381 -719
rect 632 -720 633 -719
rect 149 -722 150 -721
rect 338 -722 339 -721
rect 355 -722 356 -721
rect 450 -722 451 -721
rect 499 -722 500 -721
rect 520 -722 521 -721
rect 72 -724 73 -723
rect 499 -724 500 -723
rect 72 -726 73 -725
rect 79 -726 80 -725
rect 149 -726 150 -725
rect 310 -726 311 -725
rect 359 -726 360 -725
rect 485 -726 486 -725
rect 163 -728 164 -727
rect 240 -728 241 -727
rect 268 -728 269 -727
rect 324 -728 325 -727
rect 359 -728 360 -727
rect 534 -728 535 -727
rect 166 -730 167 -729
rect 443 -730 444 -729
rect 513 -730 514 -729
rect 534 -730 535 -729
rect 177 -732 178 -731
rect 201 -732 202 -731
rect 268 -732 269 -731
rect 639 -732 640 -731
rect 191 -734 192 -733
rect 233 -734 234 -733
rect 275 -734 276 -733
rect 541 -734 542 -733
rect 187 -736 188 -735
rect 275 -736 276 -735
rect 303 -736 304 -735
rect 492 -736 493 -735
rect 310 -738 311 -737
rect 352 -738 353 -737
rect 366 -738 367 -737
rect 656 -738 657 -737
rect 352 -740 353 -739
rect 387 -740 388 -739
rect 408 -740 409 -739
rect 464 -740 465 -739
rect 282 -742 283 -741
rect 387 -742 388 -741
rect 436 -742 437 -741
rect 513 -742 514 -741
rect 362 -744 363 -743
rect 436 -744 437 -743
rect 2 -755 3 -754
rect 163 -755 164 -754
rect 184 -755 185 -754
rect 254 -755 255 -754
rect 261 -755 262 -754
rect 362 -755 363 -754
rect 373 -755 374 -754
rect 436 -755 437 -754
rect 471 -755 472 -754
rect 625 -755 626 -754
rect 23 -757 24 -756
rect 387 -757 388 -756
rect 471 -757 472 -756
rect 541 -757 542 -756
rect 558 -757 559 -756
rect 646 -757 647 -756
rect 23 -759 24 -758
rect 100 -759 101 -758
rect 114 -759 115 -758
rect 240 -759 241 -758
rect 243 -759 244 -758
rect 296 -759 297 -758
rect 299 -759 300 -758
rect 597 -759 598 -758
rect 30 -761 31 -760
rect 103 -761 104 -760
rect 114 -761 115 -760
rect 135 -761 136 -760
rect 142 -761 143 -760
rect 604 -761 605 -760
rect 30 -763 31 -762
rect 107 -763 108 -762
rect 117 -763 118 -762
rect 254 -763 255 -762
rect 261 -763 262 -762
rect 345 -763 346 -762
rect 376 -763 377 -762
rect 583 -763 584 -762
rect 597 -763 598 -762
rect 604 -763 605 -762
rect 37 -765 38 -764
rect 149 -765 150 -764
rect 152 -765 153 -764
rect 163 -765 164 -764
rect 187 -765 188 -764
rect 394 -765 395 -764
rect 474 -765 475 -764
rect 555 -765 556 -764
rect 583 -765 584 -764
rect 611 -765 612 -764
rect 54 -767 55 -766
rect 352 -767 353 -766
rect 376 -767 377 -766
rect 618 -767 619 -766
rect 61 -769 62 -768
rect 639 -769 640 -768
rect 65 -771 66 -770
rect 229 -771 230 -770
rect 268 -771 269 -770
rect 317 -771 318 -770
rect 327 -771 328 -770
rect 415 -771 416 -770
rect 443 -771 444 -770
rect 555 -771 556 -770
rect 618 -771 619 -770
rect 660 -771 661 -770
rect 65 -773 66 -772
rect 156 -773 157 -772
rect 191 -773 192 -772
rect 338 -773 339 -772
rect 345 -773 346 -772
rect 359 -773 360 -772
rect 380 -773 381 -772
rect 513 -773 514 -772
rect 541 -773 542 -772
rect 590 -773 591 -772
rect 79 -775 80 -774
rect 548 -775 549 -774
rect 82 -777 83 -776
rect 492 -777 493 -776
rect 44 -779 45 -778
rect 82 -779 83 -778
rect 86 -779 87 -778
rect 205 -779 206 -778
rect 208 -779 209 -778
rect 576 -779 577 -778
rect 96 -781 97 -780
rect 100 -781 101 -780
rect 107 -781 108 -780
rect 121 -781 122 -780
rect 145 -781 146 -780
rect 170 -781 171 -780
rect 198 -781 199 -780
rect 478 -781 479 -780
rect 93 -783 94 -782
rect 121 -783 122 -782
rect 149 -783 150 -782
rect 205 -783 206 -782
rect 219 -783 220 -782
rect 226 -783 227 -782
rect 268 -783 269 -782
rect 310 -783 311 -782
rect 331 -783 332 -782
rect 513 -783 514 -782
rect 156 -785 157 -784
rect 177 -785 178 -784
rect 219 -785 220 -784
rect 653 -785 654 -784
rect 58 -787 59 -786
rect 177 -787 178 -786
rect 275 -787 276 -786
rect 324 -787 325 -786
rect 359 -787 360 -786
rect 366 -787 367 -786
rect 373 -787 374 -786
rect 590 -787 591 -786
rect 58 -789 59 -788
rect 72 -789 73 -788
rect 170 -789 171 -788
rect 282 -789 283 -788
rect 285 -789 286 -788
rect 499 -789 500 -788
rect 72 -791 73 -790
rect 128 -791 129 -790
rect 275 -791 276 -790
rect 632 -791 633 -790
rect 278 -793 279 -792
rect 464 -793 465 -792
rect 499 -793 500 -792
rect 520 -793 521 -792
rect 198 -795 199 -794
rect 278 -795 279 -794
rect 289 -795 290 -794
rect 408 -795 409 -794
rect 411 -795 412 -794
rect 548 -795 549 -794
rect 212 -797 213 -796
rect 408 -797 409 -796
rect 415 -797 416 -796
rect 527 -797 528 -796
rect 152 -799 153 -798
rect 212 -799 213 -798
rect 233 -799 234 -798
rect 289 -799 290 -798
rect 303 -799 304 -798
rect 331 -799 332 -798
rect 380 -799 381 -798
rect 429 -799 430 -798
rect 443 -799 444 -798
rect 534 -799 535 -798
rect 51 -801 52 -800
rect 233 -801 234 -800
rect 310 -801 311 -800
rect 506 -801 507 -800
rect 527 -801 528 -800
rect 562 -801 563 -800
rect 320 -803 321 -802
rect 366 -803 367 -802
rect 387 -803 388 -802
rect 520 -803 521 -802
rect 562 -803 563 -802
rect 569 -803 570 -802
rect 341 -805 342 -804
rect 506 -805 507 -804
rect 341 -807 342 -806
rect 436 -807 437 -806
rect 450 -807 451 -806
rect 576 -807 577 -806
rect 390 -809 391 -808
rect 492 -809 493 -808
rect 394 -811 395 -810
rect 401 -811 402 -810
rect 422 -811 423 -810
rect 429 -811 430 -810
rect 450 -811 451 -810
rect 485 -811 486 -810
rect 313 -813 314 -812
rect 422 -813 423 -812
rect 457 -813 458 -812
rect 485 -813 486 -812
rect 457 -815 458 -814
rect 537 -815 538 -814
rect 464 -817 465 -816
rect 569 -817 570 -816
rect 9 -828 10 -827
rect 33 -828 34 -827
rect 40 -828 41 -827
rect 96 -828 97 -827
rect 107 -828 108 -827
rect 135 -828 136 -827
rect 149 -828 150 -827
rect 229 -828 230 -827
rect 233 -828 234 -827
rect 373 -828 374 -827
rect 387 -828 388 -827
rect 408 -828 409 -827
rect 425 -828 426 -827
rect 492 -828 493 -827
rect 513 -828 514 -827
rect 562 -828 563 -827
rect 572 -828 573 -827
rect 618 -828 619 -827
rect 16 -830 17 -829
rect 37 -830 38 -829
rect 54 -830 55 -829
rect 471 -830 472 -829
rect 478 -830 479 -829
rect 541 -830 542 -829
rect 555 -830 556 -829
rect 590 -830 591 -829
rect 30 -832 31 -831
rect 93 -832 94 -831
rect 107 -832 108 -831
rect 184 -832 185 -831
rect 194 -832 195 -831
rect 212 -832 213 -831
rect 222 -832 223 -831
rect 285 -832 286 -831
rect 292 -832 293 -831
rect 492 -832 493 -831
rect 534 -832 535 -831
rect 583 -832 584 -831
rect 58 -834 59 -833
rect 86 -834 87 -833
rect 89 -834 90 -833
rect 100 -834 101 -833
rect 114 -834 115 -833
rect 145 -834 146 -833
rect 170 -834 171 -833
rect 324 -834 325 -833
rect 334 -834 335 -833
rect 548 -834 549 -833
rect 562 -834 563 -833
rect 576 -834 577 -833
rect 23 -836 24 -835
rect 170 -836 171 -835
rect 180 -836 181 -835
rect 240 -836 241 -835
rect 247 -836 248 -835
rect 250 -836 251 -835
rect 268 -836 269 -835
rect 317 -836 318 -835
rect 320 -836 321 -835
rect 436 -836 437 -835
rect 478 -836 479 -835
rect 506 -836 507 -835
rect 548 -836 549 -835
rect 604 -836 605 -835
rect 23 -838 24 -837
rect 44 -838 45 -837
rect 51 -838 52 -837
rect 100 -838 101 -837
rect 114 -838 115 -837
rect 198 -838 199 -837
rect 226 -838 227 -837
rect 275 -838 276 -837
rect 303 -838 304 -837
rect 373 -838 374 -837
rect 401 -838 402 -837
rect 450 -838 451 -837
rect 499 -838 500 -837
rect 506 -838 507 -837
rect 51 -840 52 -839
rect 61 -840 62 -839
rect 65 -840 66 -839
rect 201 -840 202 -839
rect 247 -840 248 -839
rect 289 -840 290 -839
rect 317 -840 318 -839
rect 499 -840 500 -839
rect 65 -842 66 -841
rect 163 -842 164 -841
rect 173 -842 174 -841
rect 268 -842 269 -841
rect 320 -842 321 -841
rect 408 -842 409 -841
rect 422 -842 423 -841
rect 471 -842 472 -841
rect 72 -844 73 -843
rect 128 -844 129 -843
rect 135 -844 136 -843
rect 215 -844 216 -843
rect 250 -844 251 -843
rect 289 -844 290 -843
rect 338 -844 339 -843
rect 380 -844 381 -843
rect 404 -844 405 -843
rect 520 -844 521 -843
rect 72 -846 73 -845
rect 82 -846 83 -845
rect 86 -846 87 -845
rect 219 -846 220 -845
rect 254 -846 255 -845
rect 338 -846 339 -845
rect 345 -846 346 -845
rect 516 -846 517 -845
rect 93 -848 94 -847
rect 142 -848 143 -847
rect 163 -848 164 -847
rect 282 -848 283 -847
rect 348 -848 349 -847
rect 457 -848 458 -847
rect 121 -850 122 -849
rect 152 -850 153 -849
rect 177 -850 178 -849
rect 275 -850 276 -849
rect 352 -850 353 -849
rect 359 -850 360 -849
rect 376 -850 377 -849
rect 401 -850 402 -849
rect 436 -850 437 -849
rect 443 -850 444 -849
rect 121 -852 122 -851
rect 156 -852 157 -851
rect 184 -852 185 -851
rect 191 -852 192 -851
rect 198 -852 199 -851
rect 310 -852 311 -851
rect 331 -852 332 -851
rect 443 -852 444 -851
rect 2 -854 3 -853
rect 191 -854 192 -853
rect 205 -854 206 -853
rect 254 -854 255 -853
rect 261 -854 262 -853
rect 303 -854 304 -853
rect 345 -854 346 -853
rect 359 -854 360 -853
rect 128 -856 129 -855
rect 278 -856 279 -855
rect 296 -856 297 -855
rect 331 -856 332 -855
rect 355 -856 356 -855
rect 527 -856 528 -855
rect 156 -858 157 -857
rect 205 -858 206 -857
rect 226 -858 227 -857
rect 457 -858 458 -857
rect 520 -858 521 -857
rect 527 -858 528 -857
rect 233 -860 234 -859
rect 261 -860 262 -859
rect 296 -860 297 -859
rect 380 -860 381 -859
rect 2 -871 3 -870
rect 135 -871 136 -870
rect 152 -871 153 -870
rect 387 -871 388 -870
rect 425 -871 426 -870
rect 499 -871 500 -870
rect 516 -871 517 -870
rect 544 -871 545 -870
rect 2 -873 3 -872
rect 114 -873 115 -872
rect 121 -873 122 -872
rect 173 -873 174 -872
rect 205 -873 206 -872
rect 233 -873 234 -872
rect 247 -873 248 -872
rect 320 -873 321 -872
rect 345 -873 346 -872
rect 401 -873 402 -872
rect 443 -873 444 -872
rect 548 -873 549 -872
rect 9 -875 10 -874
rect 44 -875 45 -874
rect 47 -875 48 -874
rect 103 -875 104 -874
rect 135 -875 136 -874
rect 149 -875 150 -874
rect 156 -875 157 -874
rect 233 -875 234 -874
rect 240 -875 241 -874
rect 247 -875 248 -874
rect 261 -875 262 -874
rect 296 -875 297 -874
rect 299 -875 300 -874
rect 387 -875 388 -874
rect 401 -875 402 -874
rect 450 -875 451 -874
rect 453 -875 454 -874
rect 485 -875 486 -874
rect 520 -875 521 -874
rect 534 -875 535 -874
rect 537 -875 538 -874
rect 541 -875 542 -874
rect 548 -875 549 -874
rect 555 -875 556 -874
rect 16 -877 17 -876
rect 30 -877 31 -876
rect 44 -877 45 -876
rect 51 -877 52 -876
rect 54 -877 55 -876
rect 124 -877 125 -876
rect 142 -877 143 -876
rect 240 -877 241 -876
rect 268 -877 269 -876
rect 499 -877 500 -876
rect 520 -877 521 -876
rect 530 -877 531 -876
rect 16 -879 17 -878
rect 40 -879 41 -878
rect 61 -879 62 -878
rect 72 -879 73 -878
rect 79 -879 80 -878
rect 128 -879 129 -878
rect 173 -879 174 -878
rect 373 -879 374 -878
rect 376 -879 377 -878
rect 464 -879 465 -878
rect 485 -879 486 -878
rect 506 -879 507 -878
rect 527 -879 528 -878
rect 562 -879 563 -878
rect 23 -881 24 -880
rect 37 -881 38 -880
rect 65 -881 66 -880
rect 163 -881 164 -880
rect 191 -881 192 -880
rect 464 -881 465 -880
rect 478 -881 479 -880
rect 506 -881 507 -880
rect 23 -883 24 -882
rect 131 -883 132 -882
rect 163 -883 164 -882
rect 184 -883 185 -882
rect 208 -883 209 -882
rect 338 -883 339 -882
rect 348 -883 349 -882
rect 352 -883 353 -882
rect 380 -883 381 -882
rect 436 -883 437 -882
rect 68 -885 69 -884
rect 86 -885 87 -884
rect 93 -885 94 -884
rect 201 -885 202 -884
rect 212 -885 213 -884
rect 275 -885 276 -884
rect 282 -885 283 -884
rect 373 -885 374 -884
rect 422 -885 423 -884
rect 527 -885 528 -884
rect 79 -887 80 -886
rect 177 -887 178 -886
rect 194 -887 195 -886
rect 338 -887 339 -886
rect 352 -887 353 -886
rect 366 -887 367 -886
rect 86 -889 87 -888
rect 107 -889 108 -888
rect 121 -889 122 -888
rect 184 -889 185 -888
rect 198 -889 199 -888
rect 380 -889 381 -888
rect 96 -891 97 -890
rect 149 -891 150 -890
rect 219 -891 220 -890
rect 268 -891 269 -890
rect 275 -891 276 -890
rect 289 -891 290 -890
rect 292 -891 293 -890
rect 415 -891 416 -890
rect 100 -893 101 -892
rect 156 -893 157 -892
rect 191 -893 192 -892
rect 219 -893 220 -892
rect 222 -893 223 -892
rect 366 -893 367 -892
rect 415 -893 416 -892
rect 429 -893 430 -892
rect 100 -895 101 -894
rect 114 -895 115 -894
rect 226 -895 227 -894
rect 324 -895 325 -894
rect 331 -895 332 -894
rect 436 -895 437 -894
rect 37 -897 38 -896
rect 331 -897 332 -896
rect 408 -897 409 -896
rect 429 -897 430 -896
rect 229 -899 230 -898
rect 254 -899 255 -898
rect 282 -899 283 -898
rect 513 -899 514 -898
rect 208 -901 209 -900
rect 513 -901 514 -900
rect 243 -903 244 -902
rect 478 -903 479 -902
rect 254 -905 255 -904
rect 289 -905 290 -904
rect 292 -905 293 -904
rect 471 -905 472 -904
rect 303 -907 304 -906
rect 313 -907 314 -906
rect 317 -907 318 -906
rect 359 -907 360 -906
rect 394 -907 395 -906
rect 408 -907 409 -906
rect 65 -909 66 -908
rect 394 -909 395 -908
rect 306 -911 307 -910
rect 446 -911 447 -910
rect 310 -913 311 -912
rect 450 -913 451 -912
rect 324 -915 325 -914
rect 471 -915 472 -914
rect 9 -926 10 -925
rect 394 -926 395 -925
rect 429 -926 430 -925
rect 443 -926 444 -925
rect 450 -926 451 -925
rect 471 -926 472 -925
rect 474 -926 475 -925
rect 485 -926 486 -925
rect 506 -926 507 -925
rect 509 -926 510 -925
rect 530 -926 531 -925
rect 548 -926 549 -925
rect 16 -928 17 -927
rect 30 -928 31 -927
rect 37 -928 38 -927
rect 170 -928 171 -927
rect 173 -928 174 -927
rect 481 -928 482 -927
rect 485 -928 486 -927
rect 520 -928 521 -927
rect 23 -930 24 -929
rect 72 -930 73 -929
rect 79 -930 80 -929
rect 145 -930 146 -929
rect 149 -930 150 -929
rect 331 -930 332 -929
rect 359 -930 360 -929
rect 478 -930 479 -929
rect 506 -930 507 -929
rect 520 -930 521 -929
rect 23 -932 24 -931
rect 117 -932 118 -931
rect 163 -932 164 -931
rect 198 -932 199 -931
rect 201 -932 202 -931
rect 387 -932 388 -931
rect 415 -932 416 -931
rect 429 -932 430 -931
rect 450 -932 451 -931
rect 492 -932 493 -931
rect 44 -934 45 -933
rect 124 -934 125 -933
rect 184 -934 185 -933
rect 247 -934 248 -933
rect 264 -934 265 -933
rect 436 -934 437 -933
rect 478 -934 479 -933
rect 541 -934 542 -933
rect 54 -936 55 -935
rect 198 -936 199 -935
rect 208 -936 209 -935
rect 212 -936 213 -935
rect 226 -936 227 -935
rect 422 -936 423 -935
rect 436 -936 437 -935
rect 499 -936 500 -935
rect 58 -938 59 -937
rect 86 -938 87 -937
rect 93 -938 94 -937
rect 240 -938 241 -937
rect 268 -938 269 -937
rect 271 -938 272 -937
rect 285 -938 286 -937
rect 383 -938 384 -937
rect 387 -938 388 -937
rect 401 -938 402 -937
rect 499 -938 500 -937
rect 534 -938 535 -937
rect 58 -940 59 -939
rect 142 -940 143 -939
rect 177 -940 178 -939
rect 240 -940 241 -939
rect 268 -940 269 -939
rect 324 -940 325 -939
rect 345 -940 346 -939
rect 415 -940 416 -939
rect 2 -942 3 -941
rect 142 -942 143 -941
rect 152 -942 153 -941
rect 177 -942 178 -941
rect 187 -942 188 -941
rect 212 -942 213 -941
rect 233 -942 234 -941
rect 247 -942 248 -941
rect 271 -942 272 -941
rect 324 -942 325 -941
rect 338 -942 339 -941
rect 345 -942 346 -941
rect 359 -942 360 -941
rect 366 -942 367 -941
rect 373 -942 374 -941
rect 401 -942 402 -941
rect 30 -944 31 -943
rect 233 -944 234 -943
rect 243 -944 244 -943
rect 366 -944 367 -943
rect 373 -944 374 -943
rect 467 -944 468 -943
rect 72 -946 73 -945
rect 254 -946 255 -945
rect 299 -946 300 -945
rect 317 -946 318 -945
rect 320 -946 321 -945
rect 394 -946 395 -945
rect 79 -948 80 -947
rect 110 -948 111 -947
rect 114 -948 115 -947
rect 121 -948 122 -947
rect 187 -948 188 -947
rect 464 -948 465 -947
rect 68 -950 69 -949
rect 464 -950 465 -949
rect 86 -952 87 -951
rect 310 -952 311 -951
rect 338 -952 339 -951
rect 411 -952 412 -951
rect 93 -954 94 -953
rect 184 -954 185 -953
rect 191 -954 192 -953
rect 205 -954 206 -953
rect 208 -954 209 -953
rect 513 -954 514 -953
rect 96 -956 97 -955
rect 289 -956 290 -955
rect 303 -956 304 -955
rect 331 -956 332 -955
rect 362 -956 363 -955
rect 408 -956 409 -955
rect 100 -958 101 -957
rect 156 -958 157 -957
rect 194 -958 195 -957
rect 219 -958 220 -957
rect 254 -958 255 -957
rect 261 -958 262 -957
rect 282 -958 283 -957
rect 303 -958 304 -957
rect 306 -958 307 -957
rect 352 -958 353 -957
rect 100 -960 101 -959
rect 152 -960 153 -959
rect 170 -960 171 -959
rect 261 -960 262 -959
rect 289 -960 290 -959
rect 296 -960 297 -959
rect 310 -960 311 -959
rect 380 -960 381 -959
rect 110 -962 111 -961
rect 114 -962 115 -961
rect 128 -962 129 -961
rect 282 -962 283 -961
rect 352 -962 353 -961
rect 492 -962 493 -961
rect 135 -964 136 -963
rect 156 -964 157 -963
rect 219 -964 220 -963
rect 275 -964 276 -963
rect 65 -966 66 -965
rect 275 -966 276 -965
rect 135 -968 136 -967
rect 166 -968 167 -967
rect 16 -979 17 -978
rect 79 -979 80 -978
rect 107 -979 108 -978
rect 187 -979 188 -978
rect 219 -979 220 -978
rect 275 -979 276 -978
rect 292 -979 293 -978
rect 324 -979 325 -978
rect 331 -979 332 -978
rect 485 -979 486 -978
rect 520 -979 521 -978
rect 527 -979 528 -978
rect 23 -981 24 -980
rect 264 -981 265 -980
rect 320 -981 321 -980
rect 401 -981 402 -980
rect 408 -981 409 -980
rect 432 -981 433 -980
rect 464 -981 465 -980
rect 499 -981 500 -980
rect 26 -983 27 -982
rect 37 -983 38 -982
rect 51 -983 52 -982
rect 135 -983 136 -982
rect 156 -983 157 -982
rect 208 -983 209 -982
rect 261 -983 262 -982
rect 345 -983 346 -982
rect 352 -983 353 -982
rect 471 -983 472 -982
rect 30 -985 31 -984
rect 229 -985 230 -984
rect 271 -985 272 -984
rect 352 -985 353 -984
rect 380 -985 381 -984
rect 443 -985 444 -984
rect 446 -985 447 -984
rect 464 -985 465 -984
rect 471 -985 472 -984
rect 492 -985 493 -984
rect 37 -987 38 -986
rect 131 -987 132 -986
rect 135 -987 136 -986
rect 191 -987 192 -986
rect 208 -987 209 -986
rect 299 -987 300 -986
rect 303 -987 304 -986
rect 345 -987 346 -986
rect 411 -987 412 -986
rect 429 -987 430 -986
rect 58 -989 59 -988
rect 128 -989 129 -988
rect 131 -989 132 -988
rect 212 -989 213 -988
rect 229 -989 230 -988
rect 254 -989 255 -988
rect 278 -989 279 -988
rect 401 -989 402 -988
rect 422 -989 423 -988
rect 457 -989 458 -988
rect 58 -991 59 -990
rect 100 -991 101 -990
rect 107 -991 108 -990
rect 121 -991 122 -990
rect 128 -991 129 -990
rect 198 -991 199 -990
rect 212 -991 213 -990
rect 289 -991 290 -990
rect 296 -991 297 -990
rect 380 -991 381 -990
rect 390 -991 391 -990
rect 422 -991 423 -990
rect 429 -991 430 -990
rect 509 -991 510 -990
rect 65 -993 66 -992
rect 114 -993 115 -992
rect 121 -993 122 -992
rect 184 -993 185 -992
rect 191 -993 192 -992
rect 261 -993 262 -992
rect 299 -993 300 -992
rect 310 -993 311 -992
rect 324 -993 325 -992
rect 415 -993 416 -992
rect 443 -993 444 -992
rect 457 -993 458 -992
rect 65 -995 66 -994
rect 117 -995 118 -994
rect 156 -995 157 -994
rect 170 -995 171 -994
rect 173 -995 174 -994
rect 201 -995 202 -994
rect 233 -995 234 -994
rect 289 -995 290 -994
rect 303 -995 304 -994
rect 338 -995 339 -994
rect 394 -995 395 -994
rect 415 -995 416 -994
rect 68 -997 69 -996
rect 93 -997 94 -996
rect 100 -997 101 -996
rect 117 -997 118 -996
rect 149 -997 150 -996
rect 170 -997 171 -996
rect 177 -997 178 -996
rect 226 -997 227 -996
rect 240 -997 241 -996
rect 310 -997 311 -996
rect 338 -997 339 -996
rect 373 -997 374 -996
rect 394 -997 395 -996
rect 436 -997 437 -996
rect 30 -999 31 -998
rect 68 -999 69 -998
rect 72 -999 73 -998
rect 219 -999 220 -998
rect 236 -999 237 -998
rect 240 -999 241 -998
rect 366 -999 367 -998
rect 373 -999 374 -998
rect 436 -999 437 -998
rect 450 -999 451 -998
rect 72 -1001 73 -1000
rect 86 -1001 87 -1000
rect 110 -1001 111 -1000
rect 359 -1001 360 -1000
rect 79 -1003 80 -1002
rect 96 -1003 97 -1002
rect 163 -1003 164 -1002
rect 205 -1003 206 -1002
rect 317 -1003 318 -1002
rect 366 -1003 367 -1002
rect 177 -1005 178 -1004
rect 282 -1005 283 -1004
rect 359 -1005 360 -1004
rect 387 -1005 388 -1004
rect 198 -1007 199 -1006
rect 331 -1007 332 -1006
rect 201 -1009 202 -1008
rect 254 -1009 255 -1008
rect 268 -1009 269 -1008
rect 387 -1009 388 -1008
rect 30 -1020 31 -1019
rect 47 -1020 48 -1019
rect 51 -1020 52 -1019
rect 201 -1020 202 -1019
rect 208 -1020 209 -1019
rect 219 -1020 220 -1019
rect 247 -1020 248 -1019
rect 268 -1020 269 -1019
rect 278 -1020 279 -1019
rect 338 -1020 339 -1019
rect 355 -1020 356 -1019
rect 380 -1020 381 -1019
rect 436 -1020 437 -1019
rect 443 -1020 444 -1019
rect 453 -1020 454 -1019
rect 471 -1020 472 -1019
rect 523 -1020 524 -1019
rect 527 -1020 528 -1019
rect 58 -1022 59 -1021
rect 96 -1022 97 -1021
rect 114 -1022 115 -1021
rect 236 -1022 237 -1021
rect 240 -1022 241 -1021
rect 268 -1022 269 -1021
rect 289 -1022 290 -1021
rect 394 -1022 395 -1021
rect 443 -1022 444 -1021
rect 450 -1022 451 -1021
rect 453 -1022 454 -1021
rect 464 -1022 465 -1021
rect 516 -1022 517 -1021
rect 523 -1022 524 -1021
rect 16 -1024 17 -1023
rect 114 -1024 115 -1023
rect 121 -1024 122 -1023
rect 194 -1024 195 -1023
rect 205 -1024 206 -1023
rect 240 -1024 241 -1023
rect 247 -1024 248 -1023
rect 282 -1024 283 -1023
rect 296 -1024 297 -1023
rect 303 -1024 304 -1023
rect 324 -1024 325 -1023
rect 334 -1024 335 -1023
rect 359 -1024 360 -1023
rect 366 -1024 367 -1023
rect 369 -1024 370 -1023
rect 401 -1024 402 -1023
rect 520 -1024 521 -1023
rect 527 -1024 528 -1023
rect 65 -1026 66 -1025
rect 79 -1026 80 -1025
rect 86 -1026 87 -1025
rect 103 -1026 104 -1025
rect 107 -1026 108 -1025
rect 121 -1026 122 -1025
rect 142 -1026 143 -1025
rect 166 -1026 167 -1025
rect 177 -1026 178 -1025
rect 219 -1026 220 -1025
rect 229 -1026 230 -1025
rect 394 -1026 395 -1025
rect 72 -1028 73 -1027
rect 128 -1028 129 -1027
rect 135 -1028 136 -1027
rect 177 -1028 178 -1027
rect 184 -1028 185 -1027
rect 201 -1028 202 -1027
rect 208 -1028 209 -1027
rect 212 -1028 213 -1027
rect 215 -1028 216 -1027
rect 303 -1028 304 -1027
rect 324 -1028 325 -1027
rect 327 -1028 328 -1027
rect 380 -1028 381 -1027
rect 408 -1028 409 -1027
rect 72 -1030 73 -1029
rect 89 -1030 90 -1029
rect 93 -1030 94 -1029
rect 100 -1030 101 -1029
rect 107 -1030 108 -1029
rect 292 -1030 293 -1029
rect 387 -1030 388 -1029
rect 408 -1030 409 -1029
rect 86 -1032 87 -1031
rect 117 -1032 118 -1031
rect 135 -1032 136 -1031
rect 149 -1032 150 -1031
rect 156 -1032 157 -1031
rect 191 -1032 192 -1031
rect 212 -1032 213 -1031
rect 359 -1032 360 -1031
rect 37 -1034 38 -1033
rect 149 -1034 150 -1033
rect 163 -1034 164 -1033
rect 184 -1034 185 -1033
rect 187 -1034 188 -1033
rect 254 -1034 255 -1033
rect 261 -1034 262 -1033
rect 338 -1034 339 -1033
rect 117 -1036 118 -1035
rect 226 -1036 227 -1035
rect 233 -1036 234 -1035
rect 292 -1036 293 -1035
rect 331 -1036 332 -1035
rect 387 -1036 388 -1035
rect 170 -1038 171 -1037
rect 229 -1038 230 -1037
rect 250 -1038 251 -1037
rect 345 -1038 346 -1037
rect 226 -1040 227 -1039
rect 373 -1040 374 -1039
rect 261 -1042 262 -1041
rect 275 -1042 276 -1041
rect 285 -1042 286 -1041
rect 401 -1042 402 -1041
rect 275 -1044 276 -1043
rect 317 -1044 318 -1043
rect 345 -1044 346 -1043
rect 352 -1044 353 -1043
rect 373 -1044 374 -1043
rect 429 -1044 430 -1043
rect 254 -1046 255 -1045
rect 317 -1046 318 -1045
rect 51 -1057 52 -1056
rect 117 -1057 118 -1056
rect 128 -1057 129 -1056
rect 180 -1057 181 -1056
rect 201 -1057 202 -1056
rect 303 -1057 304 -1056
rect 320 -1057 321 -1056
rect 380 -1057 381 -1056
rect 429 -1057 430 -1056
rect 436 -1057 437 -1056
rect 457 -1057 458 -1056
rect 464 -1057 465 -1056
rect 520 -1057 521 -1056
rect 527 -1057 528 -1056
rect 61 -1059 62 -1058
rect 89 -1059 90 -1058
rect 93 -1059 94 -1058
rect 103 -1059 104 -1058
rect 107 -1059 108 -1058
rect 254 -1059 255 -1058
rect 334 -1059 335 -1058
rect 373 -1059 374 -1058
rect 408 -1059 409 -1058
rect 429 -1059 430 -1058
rect 65 -1061 66 -1060
rect 79 -1061 80 -1060
rect 93 -1061 94 -1060
rect 149 -1061 150 -1060
rect 152 -1061 153 -1060
rect 261 -1061 262 -1060
rect 359 -1061 360 -1060
rect 362 -1061 363 -1060
rect 373 -1061 374 -1060
rect 380 -1061 381 -1060
rect 408 -1061 409 -1060
rect 415 -1061 416 -1060
rect 65 -1063 66 -1062
rect 131 -1063 132 -1062
rect 135 -1063 136 -1062
rect 159 -1063 160 -1062
rect 163 -1063 164 -1062
rect 166 -1063 167 -1062
rect 177 -1063 178 -1062
rect 208 -1063 209 -1062
rect 212 -1063 213 -1062
rect 275 -1063 276 -1062
rect 359 -1063 360 -1062
rect 366 -1063 367 -1062
rect 72 -1065 73 -1064
rect 110 -1065 111 -1064
rect 135 -1065 136 -1064
rect 299 -1065 300 -1064
rect 366 -1065 367 -1064
rect 401 -1065 402 -1064
rect 75 -1067 76 -1066
rect 107 -1067 108 -1066
rect 145 -1067 146 -1066
rect 215 -1067 216 -1066
rect 219 -1067 220 -1066
rect 222 -1067 223 -1066
rect 226 -1067 227 -1066
rect 247 -1067 248 -1066
rect 250 -1067 251 -1066
rect 387 -1067 388 -1066
rect 394 -1067 395 -1066
rect 401 -1067 402 -1066
rect 100 -1069 101 -1068
rect 142 -1069 143 -1068
rect 149 -1069 150 -1068
rect 233 -1069 234 -1068
rect 236 -1069 237 -1068
rect 422 -1069 423 -1068
rect 156 -1071 157 -1070
rect 205 -1071 206 -1070
rect 219 -1071 220 -1070
rect 331 -1071 332 -1070
rect 163 -1073 164 -1072
rect 170 -1073 171 -1072
rect 177 -1073 178 -1072
rect 198 -1073 199 -1072
rect 236 -1073 237 -1072
rect 352 -1073 353 -1072
rect 184 -1075 185 -1074
rect 212 -1075 213 -1074
rect 247 -1075 248 -1074
rect 292 -1075 293 -1074
rect 306 -1075 307 -1074
rect 387 -1075 388 -1074
rect 191 -1077 192 -1076
rect 205 -1077 206 -1076
rect 254 -1077 255 -1076
rect 268 -1077 269 -1076
rect 275 -1077 276 -1076
rect 317 -1077 318 -1076
rect 362 -1077 363 -1076
rect 394 -1077 395 -1076
rect 142 -1079 143 -1078
rect 317 -1079 318 -1078
rect 261 -1081 262 -1080
rect 289 -1081 290 -1080
rect 268 -1083 269 -1082
rect 282 -1083 283 -1082
rect 289 -1083 290 -1082
rect 338 -1083 339 -1082
rect 282 -1085 283 -1084
rect 390 -1085 391 -1084
rect 324 -1087 325 -1086
rect 338 -1087 339 -1086
rect 310 -1089 311 -1088
rect 324 -1089 325 -1088
rect 296 -1091 297 -1090
rect 310 -1091 311 -1090
rect 30 -1102 31 -1101
rect 93 -1102 94 -1101
rect 100 -1102 101 -1101
rect 110 -1102 111 -1101
rect 114 -1102 115 -1101
rect 222 -1102 223 -1101
rect 226 -1102 227 -1101
rect 443 -1102 444 -1101
rect 460 -1102 461 -1101
rect 464 -1102 465 -1101
rect 37 -1104 38 -1103
rect 236 -1104 237 -1103
rect 254 -1104 255 -1103
rect 299 -1104 300 -1103
rect 306 -1104 307 -1103
rect 345 -1104 346 -1103
rect 352 -1104 353 -1103
rect 418 -1104 419 -1103
rect 422 -1104 423 -1103
rect 436 -1104 437 -1103
rect 51 -1106 52 -1105
rect 89 -1106 90 -1105
rect 100 -1106 101 -1105
rect 114 -1106 115 -1105
rect 121 -1106 122 -1105
rect 138 -1106 139 -1105
rect 142 -1106 143 -1105
rect 177 -1106 178 -1105
rect 184 -1106 185 -1105
rect 247 -1106 248 -1105
rect 254 -1106 255 -1105
rect 352 -1106 353 -1105
rect 359 -1106 360 -1105
rect 373 -1106 374 -1105
rect 387 -1106 388 -1105
rect 408 -1106 409 -1105
rect 415 -1106 416 -1105
rect 429 -1106 430 -1105
rect 54 -1108 55 -1107
rect 58 -1108 59 -1107
rect 65 -1108 66 -1107
rect 187 -1108 188 -1107
rect 219 -1108 220 -1107
rect 303 -1108 304 -1107
rect 317 -1108 318 -1107
rect 338 -1108 339 -1107
rect 345 -1108 346 -1107
rect 359 -1108 360 -1107
rect 362 -1108 363 -1107
rect 366 -1108 367 -1107
rect 380 -1108 381 -1107
rect 408 -1108 409 -1107
rect 65 -1110 66 -1109
rect 156 -1110 157 -1109
rect 163 -1110 164 -1109
rect 191 -1110 192 -1109
rect 226 -1110 227 -1109
rect 240 -1110 241 -1109
rect 247 -1110 248 -1109
rect 268 -1110 269 -1109
rect 320 -1110 321 -1109
rect 373 -1110 374 -1109
rect 394 -1110 395 -1109
rect 422 -1110 423 -1109
rect 72 -1112 73 -1111
rect 79 -1112 80 -1111
rect 82 -1112 83 -1111
rect 86 -1112 87 -1111
rect 121 -1112 122 -1111
rect 135 -1112 136 -1111
rect 142 -1112 143 -1111
rect 149 -1112 150 -1111
rect 159 -1112 160 -1111
rect 163 -1112 164 -1111
rect 170 -1112 171 -1111
rect 184 -1112 185 -1111
rect 191 -1112 192 -1111
rect 208 -1112 209 -1111
rect 233 -1112 234 -1111
rect 376 -1112 377 -1111
rect 401 -1112 402 -1111
rect 429 -1112 430 -1111
rect 44 -1114 45 -1113
rect 79 -1114 80 -1113
rect 107 -1114 108 -1113
rect 135 -1114 136 -1113
rect 170 -1114 171 -1113
rect 212 -1114 213 -1113
rect 268 -1114 269 -1113
rect 282 -1114 283 -1113
rect 289 -1114 290 -1113
rect 320 -1114 321 -1113
rect 324 -1114 325 -1113
rect 380 -1114 381 -1113
rect 75 -1116 76 -1115
rect 107 -1116 108 -1115
rect 131 -1116 132 -1115
rect 149 -1116 150 -1115
rect 198 -1116 199 -1115
rect 212 -1116 213 -1115
rect 278 -1116 279 -1115
rect 394 -1116 395 -1115
rect 205 -1118 206 -1117
rect 240 -1118 241 -1117
rect 282 -1118 283 -1117
rect 310 -1118 311 -1117
rect 331 -1118 332 -1117
rect 415 -1118 416 -1117
rect 194 -1120 195 -1119
rect 310 -1120 311 -1119
rect 338 -1120 339 -1119
rect 369 -1120 370 -1119
rect 205 -1122 206 -1121
rect 387 -1122 388 -1121
rect 261 -1124 262 -1123
rect 331 -1124 332 -1123
rect 180 -1126 181 -1125
rect 261 -1126 262 -1125
rect 296 -1126 297 -1125
rect 401 -1126 402 -1125
rect 264 -1128 265 -1127
rect 296 -1128 297 -1127
rect 30 -1139 31 -1138
rect 96 -1139 97 -1138
rect 107 -1139 108 -1138
rect 128 -1139 129 -1138
rect 149 -1139 150 -1138
rect 198 -1139 199 -1138
rect 205 -1139 206 -1138
rect 240 -1139 241 -1138
rect 250 -1139 251 -1138
rect 268 -1139 269 -1138
rect 275 -1139 276 -1138
rect 380 -1139 381 -1138
rect 397 -1139 398 -1138
rect 436 -1139 437 -1138
rect 478 -1139 479 -1138
rect 485 -1139 486 -1138
rect 37 -1141 38 -1140
rect 170 -1141 171 -1140
rect 184 -1141 185 -1140
rect 198 -1141 199 -1140
rect 229 -1141 230 -1140
rect 275 -1141 276 -1140
rect 296 -1141 297 -1140
rect 324 -1141 325 -1140
rect 327 -1141 328 -1140
rect 401 -1141 402 -1140
rect 44 -1143 45 -1142
rect 54 -1143 55 -1142
rect 58 -1143 59 -1142
rect 72 -1143 73 -1142
rect 75 -1143 76 -1142
rect 82 -1143 83 -1142
rect 86 -1143 87 -1142
rect 243 -1143 244 -1142
rect 254 -1143 255 -1142
rect 443 -1143 444 -1142
rect 65 -1145 66 -1144
rect 159 -1145 160 -1144
rect 163 -1145 164 -1144
rect 173 -1145 174 -1144
rect 184 -1145 185 -1144
rect 205 -1145 206 -1144
rect 261 -1145 262 -1144
rect 282 -1145 283 -1144
rect 299 -1145 300 -1144
rect 415 -1145 416 -1144
rect 79 -1147 80 -1146
rect 100 -1147 101 -1146
rect 107 -1147 108 -1146
rect 121 -1147 122 -1146
rect 128 -1147 129 -1146
rect 303 -1147 304 -1146
rect 306 -1147 307 -1146
rect 429 -1147 430 -1146
rect 89 -1149 90 -1148
rect 114 -1149 115 -1148
rect 117 -1149 118 -1148
rect 166 -1149 167 -1148
rect 201 -1149 202 -1148
rect 282 -1149 283 -1148
rect 306 -1149 307 -1148
rect 359 -1149 360 -1148
rect 369 -1149 370 -1148
rect 408 -1149 409 -1148
rect 93 -1151 94 -1150
rect 208 -1151 209 -1150
rect 261 -1151 262 -1150
rect 373 -1151 374 -1150
rect 376 -1151 377 -1150
rect 422 -1151 423 -1150
rect 100 -1153 101 -1152
rect 124 -1153 125 -1152
rect 149 -1153 150 -1152
rect 191 -1153 192 -1152
rect 208 -1153 209 -1152
rect 394 -1153 395 -1152
rect 401 -1153 402 -1152
rect 408 -1153 409 -1152
rect 117 -1155 118 -1154
rect 226 -1155 227 -1154
rect 268 -1155 269 -1154
rect 289 -1155 290 -1154
rect 310 -1155 311 -1154
rect 380 -1155 381 -1154
rect 121 -1157 122 -1156
rect 135 -1157 136 -1156
rect 156 -1157 157 -1156
rect 170 -1157 171 -1156
rect 191 -1157 192 -1156
rect 219 -1157 220 -1156
rect 278 -1157 279 -1156
rect 310 -1157 311 -1156
rect 317 -1157 318 -1156
rect 331 -1157 332 -1156
rect 338 -1157 339 -1156
rect 366 -1157 367 -1156
rect 135 -1159 136 -1158
rect 145 -1159 146 -1158
rect 163 -1159 164 -1158
rect 289 -1159 290 -1158
rect 212 -1161 213 -1160
rect 226 -1161 227 -1160
rect 240 -1161 241 -1160
rect 338 -1161 339 -1160
rect 142 -1163 143 -1162
rect 212 -1163 213 -1162
rect 219 -1163 220 -1162
rect 233 -1163 234 -1162
rect 264 -1163 265 -1162
rect 331 -1163 332 -1162
rect 233 -1165 234 -1164
rect 247 -1165 248 -1164
rect 264 -1165 265 -1164
rect 387 -1165 388 -1164
rect 352 -1167 353 -1166
rect 387 -1167 388 -1166
rect 345 -1169 346 -1168
rect 352 -1169 353 -1168
rect 254 -1171 255 -1170
rect 345 -1171 346 -1170
rect 61 -1182 62 -1181
rect 72 -1182 73 -1181
rect 79 -1182 80 -1181
rect 135 -1182 136 -1181
rect 163 -1182 164 -1181
rect 184 -1182 185 -1181
rect 198 -1182 199 -1181
rect 205 -1182 206 -1181
rect 208 -1182 209 -1181
rect 212 -1182 213 -1181
rect 240 -1182 241 -1181
rect 282 -1182 283 -1181
rect 292 -1182 293 -1181
rect 401 -1182 402 -1181
rect 72 -1184 73 -1183
rect 114 -1184 115 -1183
rect 121 -1184 122 -1183
rect 149 -1184 150 -1183
rect 177 -1184 178 -1183
rect 208 -1184 209 -1183
rect 212 -1184 213 -1183
rect 240 -1184 241 -1183
rect 247 -1184 248 -1183
rect 268 -1184 269 -1183
rect 303 -1184 304 -1183
rect 380 -1184 381 -1183
rect 86 -1186 87 -1185
rect 170 -1186 171 -1185
rect 173 -1186 174 -1185
rect 247 -1186 248 -1185
rect 250 -1186 251 -1185
rect 373 -1186 374 -1185
rect 376 -1186 377 -1185
rect 394 -1186 395 -1185
rect 65 -1188 66 -1187
rect 170 -1188 171 -1187
rect 184 -1188 185 -1187
rect 226 -1188 227 -1187
rect 254 -1188 255 -1187
rect 345 -1188 346 -1187
rect 366 -1188 367 -1187
rect 380 -1188 381 -1187
rect 93 -1190 94 -1189
rect 124 -1190 125 -1189
rect 128 -1190 129 -1189
rect 198 -1190 199 -1189
rect 201 -1190 202 -1189
rect 268 -1190 269 -1189
rect 324 -1190 325 -1189
rect 327 -1190 328 -1189
rect 366 -1190 367 -1189
rect 387 -1190 388 -1189
rect 107 -1192 108 -1191
rect 131 -1192 132 -1191
rect 194 -1192 195 -1191
rect 282 -1192 283 -1191
rect 324 -1192 325 -1191
rect 338 -1192 339 -1191
rect 383 -1192 384 -1191
rect 387 -1192 388 -1191
rect 100 -1194 101 -1193
rect 107 -1194 108 -1193
rect 114 -1194 115 -1193
rect 156 -1194 157 -1193
rect 233 -1194 234 -1193
rect 345 -1194 346 -1193
rect 100 -1196 101 -1195
rect 261 -1196 262 -1195
rect 338 -1196 339 -1195
rect 352 -1196 353 -1195
rect 121 -1198 122 -1197
rect 219 -1198 220 -1197
rect 233 -1198 234 -1197
rect 296 -1198 297 -1197
rect 327 -1198 328 -1197
rect 352 -1198 353 -1197
rect 142 -1200 143 -1199
rect 156 -1200 157 -1199
rect 191 -1200 192 -1199
rect 219 -1200 220 -1199
rect 257 -1200 258 -1199
rect 275 -1200 276 -1199
rect 296 -1200 297 -1199
rect 310 -1200 311 -1199
rect 138 -1202 139 -1201
rect 191 -1202 192 -1201
rect 275 -1202 276 -1201
rect 289 -1202 290 -1201
rect 310 -1202 311 -1201
rect 317 -1202 318 -1201
rect 65 -1213 66 -1212
rect 191 -1213 192 -1212
rect 194 -1213 195 -1212
rect 247 -1213 248 -1212
rect 261 -1213 262 -1212
rect 289 -1213 290 -1212
rect 292 -1213 293 -1212
rect 352 -1213 353 -1212
rect 380 -1213 381 -1212
rect 387 -1213 388 -1212
rect 72 -1215 73 -1214
rect 89 -1215 90 -1214
rect 114 -1215 115 -1214
rect 156 -1215 157 -1214
rect 170 -1215 171 -1214
rect 247 -1215 248 -1214
rect 261 -1215 262 -1214
rect 373 -1215 374 -1214
rect 383 -1215 384 -1214
rect 394 -1215 395 -1214
rect 79 -1217 80 -1216
rect 138 -1217 139 -1216
rect 149 -1217 150 -1216
rect 219 -1217 220 -1216
rect 240 -1217 241 -1216
rect 359 -1217 360 -1216
rect 107 -1219 108 -1218
rect 114 -1219 115 -1218
rect 121 -1219 122 -1218
rect 243 -1219 244 -1218
rect 264 -1219 265 -1218
rect 345 -1219 346 -1218
rect 352 -1219 353 -1218
rect 366 -1219 367 -1218
rect 121 -1221 122 -1220
rect 180 -1221 181 -1220
rect 184 -1221 185 -1220
rect 226 -1221 227 -1220
rect 275 -1221 276 -1220
rect 317 -1221 318 -1220
rect 324 -1221 325 -1220
rect 331 -1221 332 -1220
rect 128 -1223 129 -1222
rect 159 -1223 160 -1222
rect 177 -1223 178 -1222
rect 254 -1223 255 -1222
rect 268 -1223 269 -1222
rect 317 -1223 318 -1222
rect 331 -1223 332 -1222
rect 338 -1223 339 -1222
rect 100 -1225 101 -1224
rect 128 -1225 129 -1224
rect 135 -1225 136 -1224
rect 187 -1225 188 -1224
rect 205 -1225 206 -1224
rect 212 -1225 213 -1224
rect 233 -1225 234 -1224
rect 268 -1225 269 -1224
rect 303 -1225 304 -1224
rect 310 -1225 311 -1224
rect 142 -1227 143 -1226
rect 180 -1227 181 -1226
rect 198 -1227 199 -1226
rect 233 -1227 234 -1226
rect 240 -1227 241 -1226
rect 254 -1227 255 -1226
rect 282 -1227 283 -1226
rect 310 -1227 311 -1226
rect 142 -1229 143 -1228
rect 152 -1229 153 -1228
rect 212 -1229 213 -1228
rect 229 -1229 230 -1228
rect 282 -1229 283 -1228
rect 296 -1229 297 -1228
rect 275 -1231 276 -1230
rect 296 -1231 297 -1230
rect 82 -1242 83 -1241
rect 86 -1242 87 -1241
rect 93 -1242 94 -1241
rect 100 -1242 101 -1241
rect 107 -1242 108 -1241
rect 117 -1242 118 -1241
rect 128 -1242 129 -1241
rect 152 -1242 153 -1241
rect 156 -1242 157 -1241
rect 201 -1242 202 -1241
rect 212 -1242 213 -1241
rect 219 -1242 220 -1241
rect 233 -1242 234 -1241
rect 261 -1242 262 -1241
rect 275 -1242 276 -1241
rect 296 -1242 297 -1241
rect 299 -1242 300 -1241
rect 310 -1242 311 -1241
rect 317 -1242 318 -1241
rect 320 -1242 321 -1241
rect 348 -1242 349 -1241
rect 352 -1242 353 -1241
rect 100 -1244 101 -1243
rect 121 -1244 122 -1243
rect 128 -1244 129 -1243
rect 142 -1244 143 -1243
rect 156 -1244 157 -1243
rect 226 -1244 227 -1243
rect 240 -1244 241 -1243
rect 261 -1244 262 -1243
rect 282 -1244 283 -1243
rect 303 -1244 304 -1243
rect 306 -1244 307 -1243
rect 324 -1244 325 -1243
rect 110 -1246 111 -1245
rect 114 -1246 115 -1245
rect 135 -1246 136 -1245
rect 173 -1246 174 -1245
rect 177 -1246 178 -1245
rect 191 -1246 192 -1245
rect 198 -1246 199 -1245
rect 219 -1246 220 -1245
rect 226 -1246 227 -1245
rect 233 -1246 234 -1245
rect 254 -1246 255 -1245
rect 278 -1246 279 -1245
rect 285 -1246 286 -1245
rect 289 -1246 290 -1245
rect 324 -1246 325 -1245
rect 331 -1246 332 -1245
rect 135 -1248 136 -1247
rect 149 -1248 150 -1247
rect 163 -1248 164 -1247
rect 187 -1248 188 -1247
rect 191 -1248 192 -1247
rect 205 -1248 206 -1247
rect 268 -1248 269 -1247
rect 289 -1248 290 -1247
rect 180 -1250 181 -1249
rect 247 -1250 248 -1249
rect 205 -1252 206 -1251
rect 215 -1252 216 -1251
rect 240 -1252 241 -1251
rect 247 -1252 248 -1251
rect 75 -1263 76 -1262
rect 79 -1263 80 -1262
rect 100 -1263 101 -1262
rect 128 -1263 129 -1262
rect 135 -1263 136 -1262
rect 166 -1263 167 -1262
rect 170 -1263 171 -1262
rect 173 -1263 174 -1262
rect 205 -1263 206 -1262
rect 226 -1263 227 -1262
rect 254 -1263 255 -1262
rect 271 -1263 272 -1262
rect 275 -1263 276 -1262
rect 296 -1263 297 -1262
rect 320 -1263 321 -1262
rect 324 -1263 325 -1262
rect 380 -1263 381 -1262
rect 387 -1263 388 -1262
rect 114 -1265 115 -1264
rect 121 -1265 122 -1264
rect 135 -1265 136 -1264
rect 145 -1265 146 -1264
rect 163 -1265 164 -1264
rect 177 -1265 178 -1264
rect 191 -1265 192 -1264
rect 205 -1265 206 -1264
rect 215 -1265 216 -1264
rect 219 -1265 220 -1264
rect 261 -1265 262 -1264
rect 278 -1265 279 -1264
rect 117 -1267 118 -1266
rect 121 -1267 122 -1266
rect 268 -1267 269 -1266
rect 275 -1267 276 -1266
rect 86 -1278 87 -1277
rect 96 -1278 97 -1277
rect 107 -1278 108 -1277
rect 117 -1278 118 -1277
rect 121 -1278 122 -1277
rect 128 -1278 129 -1277
rect 135 -1278 136 -1277
rect 145 -1278 146 -1277
rect 149 -1278 150 -1277
rect 159 -1278 160 -1277
rect 219 -1278 220 -1277
rect 226 -1278 227 -1277
rect 275 -1278 276 -1277
rect 282 -1278 283 -1277
rect 299 -1278 300 -1277
rect 303 -1278 304 -1277
rect 383 -1278 384 -1277
rect 387 -1278 388 -1277
rect 156 -1280 157 -1279
rect 166 -1280 167 -1279
<< metal2 >>
rect 135 -1 136 1
rect 142 -1 143 1
rect 145 -1 146 1
rect 156 -1 157 1
rect 184 -1 185 1
rect 194 -1 195 1
rect 212 -1 213 1
rect 219 -1 220 1
rect 135 -11 136 -9
rect 149 -11 150 -9
rect 156 -16 157 -10
rect 180 -16 181 -10
rect 191 -16 192 -10
rect 198 -16 199 -10
rect 208 -16 209 -10
rect 212 -11 213 -9
rect 254 -11 255 -9
rect 254 -16 255 -10
rect 254 -11 255 -9
rect 254 -16 255 -10
rect 257 -11 258 -9
rect 261 -16 262 -10
rect 142 -13 143 -9
rect 142 -16 143 -12
rect 142 -13 143 -9
rect 142 -16 143 -12
rect 149 -16 150 -12
rect 152 -13 153 -9
rect 177 -16 178 -12
rect 184 -13 185 -9
rect 212 -16 213 -12
rect 222 -16 223 -12
rect 184 -16 185 -14
rect 205 -16 206 -14
rect 149 -26 150 -24
rect 166 -26 167 -24
rect 170 -35 171 -25
rect 184 -26 185 -24
rect 187 -35 188 -25
rect 191 -35 192 -25
rect 198 -26 199 -24
rect 219 -35 220 -25
rect 229 -35 230 -25
rect 261 -35 262 -25
rect 268 -26 269 -24
rect 271 -35 272 -25
rect 310 -26 311 -24
rect 310 -35 311 -25
rect 310 -26 311 -24
rect 310 -35 311 -25
rect 341 -35 342 -25
rect 345 -35 346 -25
rect 145 -35 146 -27
rect 149 -35 150 -27
rect 156 -28 157 -24
rect 173 -28 174 -24
rect 177 -28 178 -24
rect 208 -35 209 -27
rect 243 -28 244 -24
rect 247 -35 248 -27
rect 254 -28 255 -24
rect 254 -35 255 -27
rect 254 -28 255 -24
rect 254 -35 255 -27
rect 163 -30 164 -24
rect 163 -35 164 -29
rect 163 -30 164 -24
rect 163 -35 164 -29
rect 201 -35 202 -29
rect 212 -30 213 -24
rect 205 -32 206 -24
rect 240 -35 241 -31
rect 212 -35 213 -33
rect 233 -35 234 -33
rect 51 -58 52 -44
rect 54 -45 55 -43
rect 72 -58 73 -44
rect 96 -58 97 -44
rect 100 -45 101 -43
rect 100 -58 101 -44
rect 100 -45 101 -43
rect 100 -58 101 -44
rect 138 -58 139 -44
rect 149 -45 150 -43
rect 156 -58 157 -44
rect 198 -45 199 -43
rect 201 -58 202 -44
rect 219 -45 220 -43
rect 233 -45 234 -43
rect 233 -58 234 -44
rect 233 -45 234 -43
rect 233 -58 234 -44
rect 236 -45 237 -43
rect 247 -45 248 -43
rect 282 -58 283 -44
rect 289 -58 290 -44
rect 310 -45 311 -43
rect 310 -58 311 -44
rect 310 -45 311 -43
rect 310 -58 311 -44
rect 338 -45 339 -43
rect 338 -58 339 -44
rect 338 -45 339 -43
rect 338 -58 339 -44
rect 345 -45 346 -43
rect 352 -58 353 -44
rect 359 -45 360 -43
rect 366 -58 367 -44
rect 142 -58 143 -46
rect 198 -58 199 -46
rect 208 -47 209 -43
rect 212 -47 213 -43
rect 240 -47 241 -43
rect 243 -58 244 -46
rect 247 -58 248 -46
rect 261 -47 262 -43
rect 345 -58 346 -46
rect 362 -47 363 -43
rect 163 -49 164 -43
rect 187 -49 188 -43
rect 191 -49 192 -43
rect 205 -58 206 -48
rect 240 -58 241 -48
rect 296 -58 297 -48
rect 170 -58 171 -50
rect 275 -58 276 -50
rect 177 -53 178 -43
rect 191 -58 192 -52
rect 194 -58 195 -52
rect 219 -58 220 -52
rect 261 -58 262 -52
rect 268 -53 269 -43
rect 163 -58 164 -54
rect 177 -58 178 -54
rect 187 -58 188 -54
rect 212 -58 213 -54
rect 254 -55 255 -43
rect 268 -58 269 -54
rect 226 -58 227 -56
rect 254 -58 255 -56
rect 26 -68 27 -66
rect 26 -89 27 -67
rect 26 -68 27 -66
rect 26 -89 27 -67
rect 51 -89 52 -67
rect 72 -68 73 -66
rect 79 -89 80 -67
rect 142 -68 143 -66
rect 149 -68 150 -66
rect 187 -68 188 -66
rect 194 -89 195 -67
rect 212 -68 213 -66
rect 219 -68 220 -66
rect 275 -89 276 -67
rect 282 -68 283 -66
rect 376 -89 377 -67
rect 58 -89 59 -69
rect 145 -89 146 -69
rect 149 -89 150 -69
rect 243 -89 244 -69
rect 247 -70 248 -66
rect 303 -89 304 -69
rect 310 -70 311 -66
rect 317 -70 318 -66
rect 320 -70 321 -66
rect 331 -89 332 -69
rect 338 -70 339 -66
rect 348 -70 349 -66
rect 366 -70 367 -66
rect 366 -89 367 -69
rect 366 -70 367 -66
rect 366 -89 367 -69
rect 65 -89 66 -71
rect 170 -72 171 -66
rect 198 -89 199 -71
rect 282 -89 283 -71
rect 289 -72 290 -66
rect 310 -89 311 -71
rect 345 -89 346 -71
rect 352 -72 353 -66
rect 72 -89 73 -73
rect 86 -89 87 -73
rect 93 -74 94 -66
rect 138 -89 139 -73
rect 156 -89 157 -73
rect 187 -89 188 -73
rect 201 -74 202 -66
rect 254 -74 255 -66
rect 257 -89 258 -73
rect 324 -89 325 -73
rect 93 -89 94 -75
rect 226 -76 227 -66
rect 229 -76 230 -66
rect 317 -89 318 -75
rect 96 -78 97 -66
rect 100 -78 101 -66
rect 103 -89 104 -77
rect 114 -89 115 -77
rect 121 -89 122 -77
rect 250 -89 251 -77
rect 254 -89 255 -77
rect 268 -78 269 -66
rect 278 -78 279 -66
rect 352 -89 353 -77
rect 107 -89 108 -79
rect 135 -89 136 -79
rect 163 -80 164 -66
rect 163 -89 164 -79
rect 163 -80 164 -66
rect 163 -89 164 -79
rect 205 -80 206 -66
rect 219 -89 220 -79
rect 226 -89 227 -79
rect 289 -89 290 -79
rect 296 -80 297 -66
rect 338 -89 339 -79
rect 128 -89 129 -81
rect 191 -89 192 -81
rect 205 -89 206 -81
rect 268 -89 269 -81
rect 212 -89 213 -83
rect 236 -89 237 -83
rect 261 -84 262 -66
rect 296 -89 297 -83
rect 208 -89 209 -85
rect 261 -89 262 -85
rect 233 -88 234 -66
rect 240 -88 241 -66
rect 58 -99 59 -97
rect 170 -99 171 -97
rect 173 -99 174 -97
rect 261 -99 262 -97
rect 345 -99 346 -97
rect 345 -132 346 -98
rect 345 -99 346 -97
rect 345 -132 346 -98
rect 352 -99 353 -97
rect 380 -132 381 -98
rect 65 -101 66 -97
rect 180 -101 181 -97
rect 184 -132 185 -100
rect 212 -101 213 -97
rect 236 -101 237 -97
rect 282 -101 283 -97
rect 366 -101 367 -97
rect 373 -101 374 -97
rect 376 -101 377 -97
rect 401 -132 402 -100
rect 72 -103 73 -97
rect 103 -103 104 -97
rect 107 -103 108 -97
rect 201 -103 202 -97
rect 205 -103 206 -97
rect 219 -103 220 -97
rect 243 -103 244 -97
rect 338 -103 339 -97
rect 100 -132 101 -104
rect 114 -105 115 -97
rect 135 -132 136 -104
rect 180 -132 181 -104
rect 187 -105 188 -97
rect 303 -105 304 -97
rect 324 -105 325 -97
rect 366 -132 367 -104
rect 107 -132 108 -106
rect 121 -107 122 -97
rect 145 -107 146 -97
rect 194 -107 195 -97
rect 198 -132 199 -106
rect 271 -132 272 -106
rect 338 -132 339 -106
rect 394 -132 395 -106
rect 86 -132 87 -108
rect 121 -132 122 -108
rect 142 -109 143 -97
rect 145 -132 146 -108
rect 149 -109 150 -97
rect 226 -109 227 -97
rect 236 -132 237 -108
rect 324 -132 325 -108
rect 79 -111 80 -97
rect 142 -132 143 -110
rect 149 -132 150 -110
rect 156 -111 157 -97
rect 163 -111 164 -97
rect 212 -132 213 -110
rect 247 -111 248 -97
rect 296 -111 297 -97
rect 93 -113 94 -97
rect 156 -132 157 -112
rect 163 -132 164 -112
rect 240 -113 241 -97
rect 250 -113 251 -97
rect 296 -132 297 -112
rect 93 -132 94 -114
rect 128 -115 129 -97
rect 177 -115 178 -97
rect 226 -132 227 -114
rect 254 -115 255 -97
rect 317 -115 318 -97
rect 128 -132 129 -116
rect 170 -132 171 -116
rect 191 -117 192 -97
rect 310 -117 311 -97
rect 317 -132 318 -116
rect 331 -117 332 -97
rect 191 -132 192 -118
rect 275 -119 276 -97
rect 310 -132 311 -118
rect 331 -132 332 -118
rect 194 -132 195 -120
rect 240 -132 241 -120
rect 254 -132 255 -120
rect 264 -132 265 -120
rect 205 -132 206 -122
rect 275 -132 276 -122
rect 208 -125 209 -97
rect 261 -132 262 -124
rect 208 -132 209 -126
rect 268 -127 269 -97
rect 219 -132 220 -128
rect 250 -132 251 -128
rect 257 -129 258 -97
rect 289 -129 290 -97
rect 289 -132 290 -130
rect 303 -132 304 -130
rect 65 -167 66 -141
rect 184 -142 185 -140
rect 191 -167 192 -141
rect 341 -142 342 -140
rect 380 -142 381 -140
rect 408 -167 409 -141
rect 93 -144 94 -140
rect 124 -144 125 -140
rect 142 -144 143 -140
rect 156 -167 157 -143
rect 170 -144 171 -140
rect 240 -144 241 -140
rect 243 -167 244 -143
rect 415 -167 416 -143
rect 93 -167 94 -145
rect 117 -146 118 -140
rect 121 -167 122 -145
rect 149 -146 150 -140
rect 163 -146 164 -140
rect 170 -167 171 -145
rect 184 -167 185 -145
rect 236 -146 237 -140
rect 264 -146 265 -140
rect 352 -167 353 -145
rect 380 -167 381 -145
rect 387 -167 388 -145
rect 401 -146 402 -140
rect 429 -167 430 -145
rect 72 -167 73 -147
rect 149 -167 150 -147
rect 152 -167 153 -147
rect 163 -167 164 -147
rect 205 -148 206 -140
rect 212 -148 213 -140
rect 226 -167 227 -147
rect 261 -167 262 -147
rect 275 -148 276 -140
rect 275 -167 276 -147
rect 275 -148 276 -140
rect 275 -167 276 -147
rect 289 -148 290 -140
rect 422 -167 423 -147
rect 86 -150 87 -140
rect 117 -167 118 -149
rect 177 -167 178 -149
rect 212 -167 213 -149
rect 233 -167 234 -149
rect 254 -150 255 -140
rect 289 -167 290 -149
rect 296 -150 297 -140
rect 310 -150 311 -140
rect 317 -150 318 -140
rect 331 -150 332 -140
rect 359 -167 360 -149
rect 394 -150 395 -140
rect 401 -167 402 -149
rect 86 -167 87 -151
rect 128 -152 129 -140
rect 229 -152 230 -140
rect 254 -167 255 -151
rect 285 -167 286 -151
rect 296 -167 297 -151
rect 317 -167 318 -151
rect 373 -167 374 -151
rect 107 -154 108 -140
rect 173 -154 174 -140
rect 331 -167 332 -153
rect 355 -154 356 -140
rect 366 -154 367 -140
rect 394 -167 395 -153
rect 107 -167 108 -155
rect 135 -156 136 -140
rect 142 -167 143 -155
rect 229 -167 230 -155
rect 324 -156 325 -140
rect 366 -167 367 -155
rect 100 -158 101 -140
rect 135 -167 136 -157
rect 219 -158 220 -140
rect 324 -167 325 -157
rect 341 -167 342 -157
rect 345 -158 346 -140
rect 100 -167 101 -159
rect 198 -160 199 -140
rect 303 -160 304 -140
rect 345 -167 346 -159
rect 128 -167 129 -161
rect 205 -167 206 -161
rect 247 -162 248 -140
rect 303 -167 304 -161
rect 198 -167 199 -163
rect 268 -167 269 -163
rect 247 -167 248 -165
rect 282 -166 283 -140
rect 23 -206 24 -176
rect 68 -206 69 -176
rect 72 -177 73 -175
rect 201 -177 202 -175
rect 205 -177 206 -175
rect 208 -205 209 -176
rect 219 -177 220 -175
rect 303 -177 304 -175
rect 313 -177 314 -175
rect 352 -177 353 -175
rect 387 -177 388 -175
rect 408 -177 409 -175
rect 411 -206 412 -176
rect 436 -206 437 -176
rect 37 -206 38 -178
rect 243 -179 244 -175
rect 261 -179 262 -175
rect 261 -206 262 -178
rect 261 -179 262 -175
rect 261 -206 262 -178
rect 285 -179 286 -175
rect 331 -179 332 -175
rect 341 -179 342 -175
rect 457 -206 458 -178
rect 44 -206 45 -180
rect 79 -181 80 -175
rect 82 -181 83 -175
rect 131 -181 132 -175
rect 149 -206 150 -180
rect 156 -181 157 -175
rect 170 -181 171 -175
rect 180 -181 181 -175
rect 184 -181 185 -175
rect 184 -206 185 -180
rect 184 -181 185 -175
rect 184 -206 185 -180
rect 191 -181 192 -175
rect 219 -206 220 -180
rect 236 -206 237 -180
rect 271 -206 272 -180
rect 296 -181 297 -175
rect 310 -206 311 -180
rect 317 -181 318 -175
rect 464 -206 465 -180
rect 51 -206 52 -182
rect 107 -183 108 -175
rect 114 -183 115 -175
rect 114 -206 115 -182
rect 114 -183 115 -175
rect 114 -206 115 -182
rect 128 -206 129 -182
rect 194 -206 195 -182
rect 198 -183 199 -175
rect 233 -183 234 -175
rect 240 -183 241 -175
rect 289 -183 290 -175
rect 303 -206 304 -182
rect 324 -183 325 -175
rect 352 -206 353 -182
rect 366 -183 367 -175
rect 380 -183 381 -175
rect 387 -206 388 -182
rect 394 -183 395 -175
rect 429 -206 430 -182
rect 65 -185 66 -175
rect 226 -206 227 -184
rect 243 -206 244 -184
rect 380 -206 381 -184
rect 401 -185 402 -175
rect 439 -185 440 -175
rect 72 -206 73 -186
rect 79 -206 80 -186
rect 86 -187 87 -175
rect 152 -206 153 -186
rect 156 -206 157 -186
rect 222 -187 223 -175
rect 247 -187 248 -175
rect 331 -206 332 -186
rect 359 -187 360 -175
rect 401 -206 402 -186
rect 415 -187 416 -175
rect 443 -206 444 -186
rect 65 -206 66 -188
rect 86 -206 87 -188
rect 93 -189 94 -175
rect 142 -189 143 -175
rect 177 -206 178 -188
rect 215 -206 216 -188
rect 268 -189 269 -175
rect 341 -206 342 -188
rect 373 -206 374 -188
rect 394 -206 395 -188
rect 415 -206 416 -188
rect 432 -189 433 -175
rect 100 -191 101 -175
rect 233 -206 234 -190
rect 275 -191 276 -175
rect 317 -206 318 -190
rect 320 -191 321 -175
rect 366 -206 367 -190
rect 422 -191 423 -175
rect 450 -206 451 -190
rect 96 -206 97 -192
rect 100 -206 101 -192
rect 107 -206 108 -192
rect 163 -193 164 -175
rect 191 -206 192 -192
rect 247 -206 248 -192
rect 268 -206 269 -192
rect 422 -206 423 -192
rect 121 -195 122 -175
rect 142 -206 143 -194
rect 159 -206 160 -194
rect 275 -206 276 -194
rect 285 -206 286 -194
rect 289 -206 290 -194
rect 324 -206 325 -194
rect 359 -206 360 -194
rect 121 -206 122 -196
rect 135 -197 136 -175
rect 138 -197 139 -175
rect 170 -206 171 -196
rect 198 -206 199 -196
rect 212 -197 213 -175
rect 135 -206 136 -198
rect 145 -199 146 -175
rect 163 -206 164 -198
rect 296 -206 297 -198
rect 30 -206 31 -200
rect 145 -206 146 -200
rect 205 -206 206 -200
rect 345 -201 346 -175
rect 254 -203 255 -175
rect 345 -206 346 -202
rect 254 -206 255 -204
rect 23 -216 24 -214
rect 72 -253 73 -215
rect 100 -216 101 -214
rect 110 -253 111 -215
rect 152 -253 153 -215
rect 450 -216 451 -214
rect 457 -216 458 -214
rect 499 -253 500 -215
rect 541 -253 542 -215
rect 544 -216 545 -214
rect 30 -218 31 -214
rect 205 -218 206 -214
rect 215 -218 216 -214
rect 348 -253 349 -217
rect 380 -218 381 -214
rect 380 -253 381 -217
rect 380 -218 381 -214
rect 380 -253 381 -217
rect 408 -218 409 -214
rect 478 -253 479 -217
rect 485 -253 486 -217
rect 537 -253 538 -217
rect 37 -220 38 -214
rect 124 -253 125 -219
rect 156 -253 157 -219
rect 177 -220 178 -214
rect 184 -220 185 -214
rect 212 -253 213 -219
rect 226 -220 227 -214
rect 268 -220 269 -214
rect 271 -220 272 -214
rect 401 -220 402 -214
rect 422 -220 423 -214
rect 422 -253 423 -219
rect 422 -220 423 -214
rect 422 -253 423 -219
rect 436 -220 437 -214
rect 471 -253 472 -219
rect 37 -253 38 -221
rect 145 -222 146 -214
rect 149 -253 150 -221
rect 184 -253 185 -221
rect 191 -222 192 -214
rect 303 -222 304 -214
rect 317 -222 318 -214
rect 341 -253 342 -221
rect 345 -222 346 -214
rect 506 -253 507 -221
rect 44 -224 45 -214
rect 58 -224 59 -214
rect 65 -224 66 -214
rect 79 -224 80 -214
rect 100 -253 101 -223
rect 114 -224 115 -214
rect 142 -224 143 -214
rect 177 -253 178 -223
rect 229 -253 230 -223
rect 387 -224 388 -214
rect 429 -224 430 -214
rect 436 -253 437 -223
rect 450 -253 451 -223
rect 534 -253 535 -223
rect 44 -253 45 -225
rect 93 -226 94 -214
rect 107 -226 108 -214
rect 243 -226 244 -214
rect 247 -226 248 -214
rect 247 -253 248 -225
rect 247 -226 248 -214
rect 247 -253 248 -225
rect 261 -226 262 -214
rect 296 -253 297 -225
rect 299 -226 300 -214
rect 366 -226 367 -214
rect 464 -226 465 -214
rect 513 -253 514 -225
rect 51 -228 52 -214
rect 138 -228 139 -214
rect 159 -228 160 -214
rect 233 -253 234 -227
rect 236 -228 237 -214
rect 268 -253 269 -227
rect 275 -228 276 -214
rect 324 -253 325 -227
rect 327 -253 328 -227
rect 408 -253 409 -227
rect 443 -228 444 -214
rect 464 -253 465 -227
rect 58 -253 59 -229
rect 226 -253 227 -229
rect 240 -230 241 -214
rect 254 -230 255 -214
rect 275 -253 276 -229
rect 331 -230 332 -214
rect 338 -230 339 -214
rect 520 -253 521 -229
rect 65 -253 66 -231
rect 128 -232 129 -214
rect 163 -232 164 -214
rect 201 -232 202 -214
rect 205 -253 206 -231
rect 261 -253 262 -231
rect 285 -253 286 -231
rect 373 -253 374 -231
rect 51 -253 52 -233
rect 201 -253 202 -233
rect 219 -234 220 -214
rect 254 -253 255 -233
rect 306 -253 307 -233
rect 387 -253 388 -233
rect 79 -253 80 -235
rect 135 -236 136 -214
rect 142 -253 143 -235
rect 219 -253 220 -235
rect 310 -236 311 -214
rect 317 -253 318 -235
rect 331 -253 332 -235
rect 492 -253 493 -235
rect 86 -253 87 -237
rect 163 -253 164 -237
rect 166 -253 167 -237
rect 191 -253 192 -237
rect 198 -253 199 -237
rect 240 -253 241 -237
rect 289 -238 290 -214
rect 310 -253 311 -237
rect 338 -253 339 -237
rect 457 -253 458 -237
rect 93 -253 94 -239
rect 121 -240 122 -214
rect 135 -253 136 -239
rect 180 -253 181 -239
rect 352 -240 353 -214
rect 401 -253 402 -239
rect 89 -242 90 -214
rect 121 -253 122 -241
rect 170 -242 171 -214
rect 208 -242 209 -214
rect 355 -253 356 -241
rect 429 -253 430 -241
rect 170 -253 171 -243
rect 289 -253 290 -243
rect 366 -253 367 -243
rect 394 -244 395 -214
rect 208 -253 209 -245
rect 359 -246 360 -214
rect 394 -253 395 -245
rect 415 -246 416 -214
rect 243 -253 244 -247
rect 359 -253 360 -247
rect 282 -250 283 -214
rect 415 -253 416 -249
rect 282 -253 283 -251
rect 443 -253 444 -251
rect 37 -263 38 -261
rect 229 -263 230 -261
rect 240 -300 241 -262
rect 268 -263 269 -261
rect 282 -263 283 -261
rect 401 -263 402 -261
rect 443 -263 444 -261
rect 555 -300 556 -262
rect 562 -300 563 -262
rect 576 -300 577 -262
rect 37 -300 38 -264
rect 107 -265 108 -261
rect 142 -300 143 -264
rect 212 -265 213 -261
rect 285 -300 286 -264
rect 296 -265 297 -261
rect 303 -265 304 -261
rect 317 -265 318 -261
rect 320 -300 321 -264
rect 506 -265 507 -261
rect 527 -265 528 -261
rect 534 -265 535 -261
rect 44 -267 45 -261
rect 117 -267 118 -261
rect 152 -267 153 -261
rect 233 -300 234 -266
rect 296 -300 297 -266
rect 422 -267 423 -261
rect 464 -267 465 -261
rect 506 -300 507 -266
rect 65 -269 66 -261
rect 131 -269 132 -261
rect 156 -269 157 -261
rect 156 -300 157 -268
rect 156 -269 157 -261
rect 156 -300 157 -268
rect 163 -300 164 -268
rect 219 -269 220 -261
rect 306 -300 307 -268
rect 520 -269 521 -261
rect 65 -300 66 -270
rect 114 -271 115 -261
rect 145 -271 146 -261
rect 219 -300 220 -270
rect 310 -271 311 -261
rect 310 -300 311 -270
rect 310 -271 311 -261
rect 310 -300 311 -270
rect 324 -300 325 -270
rect 380 -271 381 -261
rect 383 -300 384 -270
rect 548 -300 549 -270
rect 75 -273 76 -261
rect 149 -273 150 -261
rect 170 -300 171 -272
rect 191 -273 192 -261
rect 198 -300 199 -272
rect 289 -273 290 -261
rect 331 -273 332 -261
rect 366 -273 367 -261
rect 373 -273 374 -261
rect 373 -300 374 -272
rect 373 -273 374 -261
rect 373 -300 374 -272
rect 408 -273 409 -261
rect 527 -300 528 -272
rect 86 -275 87 -261
rect 128 -275 129 -261
rect 149 -300 150 -274
rect 226 -275 227 -261
rect 289 -300 290 -274
rect 387 -275 388 -261
rect 408 -300 409 -274
rect 415 -275 416 -261
rect 422 -300 423 -274
rect 429 -275 430 -261
rect 485 -275 486 -261
rect 485 -300 486 -274
rect 485 -275 486 -261
rect 485 -300 486 -274
rect 492 -275 493 -261
rect 492 -300 493 -274
rect 492 -275 493 -261
rect 492 -300 493 -274
rect 499 -275 500 -261
rect 534 -300 535 -274
rect 86 -300 87 -276
rect 114 -300 115 -276
rect 173 -277 174 -261
rect 212 -300 213 -276
rect 226 -300 227 -276
rect 261 -277 262 -261
rect 334 -277 335 -261
rect 478 -277 479 -261
rect 520 -300 521 -276
rect 541 -277 542 -261
rect 79 -279 80 -261
rect 261 -300 262 -278
rect 338 -279 339 -261
rect 387 -300 388 -278
rect 394 -279 395 -261
rect 499 -300 500 -278
rect 93 -281 94 -261
rect 128 -300 129 -280
rect 191 -300 192 -280
rect 268 -300 269 -280
rect 345 -281 346 -261
rect 513 -281 514 -261
rect 96 -300 97 -282
rect 117 -300 118 -282
rect 208 -283 209 -261
rect 275 -283 276 -261
rect 317 -300 318 -282
rect 513 -300 514 -282
rect 100 -285 101 -261
rect 121 -300 122 -284
rect 275 -300 276 -284
rect 359 -285 360 -261
rect 362 -300 363 -284
rect 366 -300 367 -284
rect 415 -300 416 -284
rect 450 -285 451 -261
rect 471 -285 472 -261
rect 478 -300 479 -284
rect 51 -287 52 -261
rect 100 -300 101 -286
rect 107 -300 108 -286
rect 135 -287 136 -261
rect 243 -287 244 -261
rect 450 -300 451 -286
rect 457 -287 458 -261
rect 471 -300 472 -286
rect 51 -300 52 -288
rect 72 -289 73 -261
rect 135 -300 136 -288
rect 166 -289 167 -261
rect 205 -289 206 -261
rect 457 -300 458 -288
rect 72 -300 73 -290
rect 177 -291 178 -261
rect 184 -291 185 -261
rect 205 -300 206 -290
rect 348 -291 349 -261
rect 394 -300 395 -290
rect 429 -300 430 -290
rect 436 -291 437 -261
rect 443 -300 444 -290
rect 541 -300 542 -290
rect 58 -293 59 -261
rect 184 -300 185 -292
rect 303 -300 304 -292
rect 436 -300 437 -292
rect 177 -300 178 -294
rect 247 -295 248 -261
rect 352 -295 353 -261
rect 401 -300 402 -294
rect 247 -300 248 -296
rect 254 -297 255 -261
rect 334 -300 335 -296
rect 352 -300 353 -296
rect 79 -300 80 -298
rect 254 -300 255 -298
rect 9 -361 10 -309
rect 86 -310 87 -308
rect 93 -361 94 -309
rect 149 -310 150 -308
rect 177 -310 178 -308
rect 303 -310 304 -308
rect 334 -310 335 -308
rect 345 -310 346 -308
rect 366 -310 367 -308
rect 478 -310 479 -308
rect 485 -310 486 -308
rect 485 -361 486 -309
rect 485 -310 486 -308
rect 485 -361 486 -309
rect 520 -310 521 -308
rect 544 -310 545 -308
rect 548 -310 549 -308
rect 562 -361 563 -309
rect 16 -361 17 -311
rect 275 -312 276 -308
rect 285 -312 286 -308
rect 310 -312 311 -308
rect 334 -361 335 -311
rect 576 -312 577 -308
rect 23 -361 24 -313
rect 96 -314 97 -308
rect 100 -314 101 -308
rect 313 -361 314 -313
rect 338 -314 339 -308
rect 457 -314 458 -308
rect 464 -314 465 -308
rect 492 -314 493 -308
rect 527 -314 528 -308
rect 548 -361 549 -313
rect 30 -361 31 -315
rect 44 -316 45 -308
rect 51 -316 52 -308
rect 61 -316 62 -308
rect 65 -316 66 -308
rect 247 -316 248 -308
rect 250 -316 251 -308
rect 457 -361 458 -315
rect 471 -316 472 -308
rect 555 -361 556 -315
rect 37 -318 38 -308
rect 208 -361 209 -317
rect 240 -318 241 -308
rect 268 -318 269 -308
rect 285 -361 286 -317
rect 576 -361 577 -317
rect 44 -361 45 -319
rect 233 -320 234 -308
rect 240 -361 241 -319
rect 422 -320 423 -308
rect 429 -320 430 -308
rect 527 -361 528 -319
rect 51 -361 52 -321
rect 135 -322 136 -308
rect 180 -361 181 -321
rect 275 -361 276 -321
rect 289 -322 290 -308
rect 289 -361 290 -321
rect 289 -322 290 -308
rect 289 -361 290 -321
rect 296 -322 297 -308
rect 429 -361 430 -321
rect 450 -322 451 -308
rect 569 -322 570 -308
rect 61 -361 62 -323
rect 138 -361 139 -323
rect 184 -324 185 -308
rect 247 -361 248 -323
rect 254 -324 255 -308
rect 355 -361 356 -323
rect 373 -324 374 -308
rect 422 -361 423 -323
rect 471 -361 472 -323
rect 513 -324 514 -308
rect 65 -361 66 -325
rect 72 -326 73 -308
rect 79 -361 80 -325
rect 198 -326 199 -308
rect 226 -326 227 -308
rect 254 -361 255 -325
rect 268 -361 269 -325
rect 324 -326 325 -308
rect 348 -326 349 -308
rect 520 -361 521 -325
rect 72 -361 73 -327
rect 142 -328 143 -308
rect 184 -361 185 -327
rect 205 -328 206 -308
rect 219 -328 220 -308
rect 226 -361 227 -327
rect 282 -328 283 -308
rect 569 -361 570 -327
rect 86 -361 87 -329
rect 170 -330 171 -308
rect 194 -330 195 -308
rect 212 -330 213 -308
rect 219 -361 220 -329
rect 261 -330 262 -308
rect 299 -361 300 -329
rect 513 -361 514 -329
rect 103 -361 104 -331
rect 233 -361 234 -331
rect 261 -361 262 -331
rect 296 -361 297 -331
rect 310 -361 311 -331
rect 450 -361 451 -331
rect 107 -334 108 -308
rect 131 -334 132 -308
rect 142 -361 143 -333
rect 338 -361 339 -333
rect 348 -361 349 -333
rect 541 -334 542 -308
rect 114 -336 115 -308
rect 408 -336 409 -308
rect 534 -336 535 -308
rect 541 -361 542 -335
rect 114 -361 115 -337
rect 121 -338 122 -308
rect 149 -361 150 -337
rect 170 -361 171 -337
rect 194 -361 195 -337
rect 303 -361 304 -337
rect 317 -338 318 -308
rect 492 -361 493 -337
rect 121 -361 122 -339
rect 191 -340 192 -308
rect 198 -361 199 -339
rect 282 -361 283 -339
rect 317 -361 318 -339
rect 331 -361 332 -339
rect 345 -361 346 -339
rect 534 -361 535 -339
rect 163 -342 164 -308
rect 212 -361 213 -341
rect 352 -342 353 -308
rect 408 -361 409 -341
rect 156 -344 157 -308
rect 163 -361 164 -343
rect 352 -361 353 -343
rect 478 -361 479 -343
rect 156 -361 157 -345
rect 359 -361 360 -345
rect 373 -361 374 -345
rect 401 -346 402 -308
rect 380 -361 381 -347
rect 506 -348 507 -308
rect 383 -350 384 -308
rect 499 -350 500 -308
rect 387 -352 388 -308
rect 464 -361 465 -351
rect 341 -361 342 -353
rect 387 -361 388 -353
rect 394 -354 395 -308
rect 506 -361 507 -353
rect 271 -356 272 -308
rect 394 -361 395 -355
rect 401 -361 402 -355
rect 415 -356 416 -308
rect 443 -356 444 -308
rect 499 -361 500 -355
rect 292 -361 293 -357
rect 415 -361 416 -357
rect 436 -358 437 -308
rect 443 -361 444 -357
rect 205 -361 206 -359
rect 436 -361 437 -359
rect 2 -416 3 -370
rect 191 -371 192 -369
rect 201 -416 202 -370
rect 331 -416 332 -370
rect 345 -371 346 -369
rect 422 -371 423 -369
rect 485 -371 486 -369
rect 485 -416 486 -370
rect 485 -371 486 -369
rect 485 -416 486 -370
rect 513 -371 514 -369
rect 583 -416 584 -370
rect 9 -373 10 -369
rect 135 -373 136 -369
rect 156 -373 157 -369
rect 163 -373 164 -369
rect 184 -373 185 -369
rect 338 -416 339 -372
rect 348 -373 349 -369
rect 394 -373 395 -369
rect 422 -416 423 -372
rect 478 -373 479 -369
rect 534 -373 535 -369
rect 611 -416 612 -372
rect 16 -375 17 -369
rect 250 -416 251 -374
rect 254 -375 255 -369
rect 285 -375 286 -369
rect 296 -375 297 -369
rect 499 -375 500 -369
rect 555 -416 556 -374
rect 576 -375 577 -369
rect 23 -377 24 -369
rect 149 -377 150 -369
rect 156 -416 157 -376
rect 306 -416 307 -376
rect 313 -377 314 -369
rect 471 -377 472 -369
rect 23 -416 24 -378
rect 33 -416 34 -378
rect 37 -379 38 -369
rect 61 -379 62 -369
rect 65 -379 66 -369
rect 177 -379 178 -369
rect 219 -379 220 -369
rect 327 -379 328 -369
rect 352 -416 353 -378
rect 523 -416 524 -378
rect 30 -381 31 -369
rect 58 -381 59 -369
rect 68 -416 69 -380
rect 177 -416 178 -380
rect 226 -381 227 -369
rect 282 -416 283 -380
rect 296 -416 297 -380
rect 317 -381 318 -369
rect 355 -381 356 -369
rect 548 -381 549 -369
rect 37 -416 38 -382
rect 124 -383 125 -369
rect 149 -416 150 -382
rect 163 -416 164 -382
rect 170 -383 171 -369
rect 184 -416 185 -382
rect 299 -383 300 -369
rect 408 -383 409 -369
rect 443 -383 444 -369
rect 499 -416 500 -382
rect 44 -385 45 -369
rect 271 -385 272 -369
rect 303 -385 304 -369
rect 310 -416 311 -384
rect 366 -385 367 -369
rect 464 -385 465 -369
rect 471 -416 472 -384
rect 520 -385 521 -369
rect 44 -416 45 -386
rect 107 -387 108 -369
rect 121 -416 122 -386
rect 261 -387 262 -369
rect 268 -416 269 -386
rect 366 -416 367 -386
rect 380 -387 381 -369
rect 548 -416 549 -386
rect 51 -389 52 -369
rect 219 -416 220 -388
rect 233 -389 234 -369
rect 261 -416 262 -388
rect 320 -416 321 -388
rect 464 -416 465 -388
rect 51 -416 52 -390
rect 103 -391 104 -369
rect 107 -416 108 -390
rect 114 -391 115 -369
rect 170 -416 171 -390
rect 212 -391 213 -369
rect 233 -416 234 -390
rect 275 -391 276 -369
rect 380 -416 381 -390
rect 527 -391 528 -369
rect 58 -416 59 -392
rect 205 -416 206 -392
rect 212 -416 213 -392
rect 327 -416 328 -392
rect 390 -416 391 -392
rect 576 -416 577 -392
rect 72 -395 73 -369
rect 152 -395 153 -369
rect 191 -416 192 -394
rect 275 -416 276 -394
rect 394 -416 395 -394
rect 401 -395 402 -369
rect 408 -416 409 -394
rect 415 -395 416 -369
rect 443 -416 444 -394
rect 492 -395 493 -369
rect 527 -416 528 -394
rect 569 -395 570 -369
rect 72 -416 73 -396
rect 96 -416 97 -396
rect 100 -416 101 -396
rect 226 -416 227 -396
rect 373 -397 374 -369
rect 401 -416 402 -396
rect 415 -416 416 -396
rect 506 -397 507 -369
rect 558 -397 559 -369
rect 569 -416 570 -396
rect 79 -399 80 -369
rect 208 -399 209 -369
rect 348 -416 349 -398
rect 373 -416 374 -398
rect 387 -399 388 -369
rect 492 -416 493 -398
rect 79 -416 80 -400
rect 142 -401 143 -369
rect 152 -416 153 -400
rect 429 -401 430 -369
rect 450 -401 451 -369
rect 534 -416 535 -400
rect 86 -403 87 -369
rect 243 -403 244 -369
rect 383 -416 384 -402
rect 450 -416 451 -402
rect 457 -403 458 -369
rect 478 -416 479 -402
rect 93 -405 94 -369
rect 131 -405 132 -369
rect 138 -405 139 -369
rect 387 -416 388 -404
rect 411 -416 412 -404
rect 506 -416 507 -404
rect 9 -416 10 -406
rect 138 -416 139 -406
rect 142 -416 143 -406
rect 198 -407 199 -369
rect 243 -416 244 -406
rect 247 -407 248 -369
rect 429 -416 430 -406
rect 541 -407 542 -369
rect 114 -416 115 -408
rect 128 -409 129 -369
rect 247 -416 248 -408
rect 513 -416 514 -408
rect 541 -416 542 -408
rect 562 -409 563 -369
rect 359 -411 360 -369
rect 562 -416 563 -410
rect 436 -413 437 -369
rect 457 -416 458 -412
rect 324 -415 325 -369
rect 436 -416 437 -414
rect 2 -426 3 -424
rect 156 -426 157 -424
rect 198 -426 199 -424
rect 219 -426 220 -424
rect 240 -426 241 -424
rect 520 -493 521 -425
rect 576 -426 577 -424
rect 597 -493 598 -425
rect 611 -426 612 -424
rect 639 -493 640 -425
rect 663 -493 664 -425
rect 674 -493 675 -425
rect 2 -493 3 -427
rect 51 -428 52 -424
rect 79 -428 80 -424
rect 187 -493 188 -427
rect 208 -428 209 -424
rect 352 -428 353 -424
rect 355 -493 356 -427
rect 394 -428 395 -424
rect 464 -428 465 -424
rect 625 -493 626 -427
rect 635 -493 636 -427
rect 667 -493 668 -427
rect 9 -493 10 -429
rect 72 -430 73 -424
rect 79 -493 80 -429
rect 177 -430 178 -424
rect 257 -430 258 -424
rect 338 -430 339 -424
rect 348 -430 349 -424
rect 471 -430 472 -424
rect 506 -430 507 -424
rect 590 -493 591 -429
rect 16 -493 17 -431
rect 114 -432 115 -424
rect 128 -493 129 -431
rect 159 -432 160 -424
rect 170 -432 171 -424
rect 219 -493 220 -431
rect 268 -432 269 -424
rect 268 -493 269 -431
rect 268 -432 269 -424
rect 268 -493 269 -431
rect 271 -432 272 -424
rect 282 -432 283 -424
rect 310 -432 311 -424
rect 383 -432 384 -424
rect 422 -432 423 -424
rect 506 -493 507 -431
rect 513 -432 514 -424
rect 576 -493 577 -431
rect 583 -432 584 -424
rect 604 -493 605 -431
rect 19 -434 20 -424
rect 247 -493 248 -433
rect 275 -434 276 -424
rect 289 -434 290 -424
rect 313 -493 314 -433
rect 415 -434 416 -424
rect 436 -434 437 -424
rect 583 -493 584 -433
rect 30 -493 31 -435
rect 40 -493 41 -435
rect 44 -436 45 -424
rect 205 -436 206 -424
rect 226 -436 227 -424
rect 415 -493 416 -435
rect 492 -436 493 -424
rect 513 -493 514 -435
rect 527 -436 528 -424
rect 611 -493 612 -435
rect 44 -493 45 -437
rect 621 -493 622 -437
rect 47 -493 48 -439
rect 212 -440 213 -424
rect 233 -440 234 -424
rect 289 -493 290 -439
rect 317 -440 318 -424
rect 548 -440 549 -424
rect 51 -493 52 -441
rect 359 -442 360 -424
rect 362 -442 363 -424
rect 555 -442 556 -424
rect 68 -493 69 -443
rect 338 -493 339 -443
rect 373 -444 374 -424
rect 387 -493 388 -443
rect 401 -444 402 -424
rect 436 -493 437 -443
rect 457 -444 458 -424
rect 548 -493 549 -443
rect 72 -493 73 -445
rect 261 -446 262 -424
rect 275 -493 276 -445
rect 397 -493 398 -445
rect 478 -446 479 -424
rect 555 -493 556 -445
rect 86 -448 87 -424
rect 173 -493 174 -447
rect 177 -493 178 -447
rect 191 -448 192 -424
rect 278 -448 279 -424
rect 296 -448 297 -424
rect 303 -493 304 -447
rect 457 -493 458 -447
rect 499 -448 500 -424
rect 527 -493 528 -447
rect 86 -493 87 -449
rect 243 -450 244 -424
rect 282 -493 283 -449
rect 362 -493 363 -449
rect 380 -450 381 -424
rect 429 -450 430 -424
rect 93 -452 94 -424
rect 464 -493 465 -451
rect 93 -493 94 -453
rect 114 -493 115 -453
rect 121 -454 122 -424
rect 212 -493 213 -453
rect 243 -493 244 -453
rect 373 -493 374 -453
rect 429 -493 430 -453
rect 562 -454 563 -424
rect 96 -456 97 -424
rect 117 -493 118 -455
rect 138 -456 139 -424
rect 250 -456 251 -424
rect 296 -493 297 -455
rect 394 -493 395 -455
rect 534 -456 535 -424
rect 562 -493 563 -455
rect 100 -493 101 -457
rect 184 -458 185 -424
rect 191 -493 192 -457
rect 345 -493 346 -457
rect 145 -493 146 -459
rect 226 -493 227 -459
rect 254 -460 255 -424
rect 534 -493 535 -459
rect 149 -493 150 -461
rect 163 -462 164 -424
rect 170 -493 171 -461
rect 401 -493 402 -461
rect 58 -464 59 -424
rect 163 -493 164 -463
rect 254 -493 255 -463
rect 264 -493 265 -463
rect 310 -493 311 -463
rect 478 -493 479 -463
rect 58 -493 59 -465
rect 131 -466 132 -424
rect 156 -493 157 -465
rect 233 -493 234 -465
rect 317 -493 318 -465
rect 352 -493 353 -465
rect 37 -468 38 -424
rect 131 -493 132 -467
rect 320 -468 321 -424
rect 366 -468 367 -424
rect 23 -470 24 -424
rect 37 -493 38 -469
rect 201 -493 202 -469
rect 366 -493 367 -469
rect 23 -493 24 -471
rect 142 -472 143 -424
rect 324 -472 325 -424
rect 471 -493 472 -471
rect 135 -474 136 -424
rect 142 -493 143 -473
rect 324 -493 325 -473
rect 499 -493 500 -473
rect 107 -476 108 -424
rect 135 -493 136 -475
rect 327 -476 328 -424
rect 443 -476 444 -424
rect 107 -493 108 -477
rect 138 -493 139 -477
rect 327 -493 328 -477
rect 646 -493 647 -477
rect 124 -493 125 -479
rect 443 -493 444 -479
rect 331 -482 332 -424
rect 408 -493 409 -481
rect 331 -493 332 -483
rect 541 -484 542 -424
rect 334 -493 335 -485
rect 380 -493 381 -485
rect 450 -486 451 -424
rect 541 -493 542 -485
rect 450 -493 451 -487
rect 569 -488 570 -424
rect 485 -490 486 -424
rect 569 -493 570 -489
rect 422 -493 423 -491
rect 485 -493 486 -491
rect 2 -503 3 -501
rect 47 -503 48 -501
rect 51 -503 52 -501
rect 124 -503 125 -501
rect 128 -503 129 -501
rect 212 -503 213 -501
rect 236 -503 237 -501
rect 457 -503 458 -501
rect 492 -503 493 -501
rect 562 -503 563 -501
rect 597 -503 598 -501
rect 628 -558 629 -502
rect 635 -503 636 -501
rect 674 -503 675 -501
rect 9 -505 10 -501
rect 173 -558 174 -504
rect 205 -505 206 -501
rect 415 -505 416 -501
rect 422 -558 423 -504
rect 464 -505 465 -501
rect 492 -558 493 -504
rect 569 -505 570 -501
rect 597 -558 598 -504
rect 646 -505 647 -501
rect 16 -507 17 -501
rect 191 -507 192 -501
rect 208 -507 209 -501
rect 219 -507 220 -501
rect 240 -507 241 -501
rect 443 -507 444 -501
rect 464 -558 465 -506
rect 548 -507 549 -501
rect 604 -507 605 -501
rect 614 -558 615 -506
rect 618 -507 619 -501
rect 667 -507 668 -501
rect 16 -558 17 -508
rect 75 -558 76 -508
rect 79 -509 80 -501
rect 264 -558 265 -508
rect 289 -509 290 -501
rect 306 -509 307 -501
rect 310 -509 311 -501
rect 415 -558 416 -508
rect 513 -509 514 -501
rect 604 -558 605 -508
rect 639 -509 640 -501
rect 646 -558 647 -508
rect 23 -511 24 -501
rect 198 -511 199 -501
rect 212 -558 213 -510
rect 334 -511 335 -501
rect 345 -511 346 -501
rect 548 -558 549 -510
rect 576 -511 577 -501
rect 618 -558 619 -510
rect 23 -558 24 -512
rect 30 -513 31 -501
rect 37 -558 38 -512
rect 394 -558 395 -512
rect 397 -513 398 -501
rect 527 -513 528 -501
rect 541 -513 542 -501
rect 541 -558 542 -512
rect 541 -513 542 -501
rect 541 -558 542 -512
rect 30 -558 31 -514
rect 72 -515 73 -501
rect 86 -515 87 -501
rect 152 -558 153 -514
rect 170 -515 171 -501
rect 506 -515 507 -501
rect 513 -558 514 -514
rect 555 -515 556 -501
rect 51 -558 52 -516
rect 331 -517 332 -501
rect 334 -558 335 -516
rect 569 -558 570 -516
rect 58 -519 59 -501
rect 208 -558 209 -518
rect 303 -519 304 -501
rect 499 -519 500 -501
rect 527 -558 528 -518
rect 653 -519 654 -501
rect 86 -558 87 -520
rect 282 -521 283 -501
rect 310 -558 311 -520
rect 366 -521 367 -501
rect 369 -558 370 -520
rect 499 -558 500 -520
rect 555 -558 556 -520
rect 590 -521 591 -501
rect 621 -521 622 -501
rect 653 -558 654 -520
rect 93 -523 94 -501
rect 114 -558 115 -522
rect 131 -523 132 -501
rect 562 -558 563 -522
rect 590 -558 591 -522
rect 625 -523 626 -501
rect 93 -558 94 -524
rect 278 -558 279 -524
rect 282 -558 283 -524
rect 352 -558 353 -524
rect 355 -525 356 -501
rect 478 -525 479 -501
rect 495 -525 496 -501
rect 506 -558 507 -524
rect 625 -558 626 -524
rect 642 -558 643 -524
rect 100 -527 101 -501
rect 184 -558 185 -526
rect 191 -558 192 -526
rect 226 -527 227 -501
rect 275 -527 276 -501
rect 303 -558 304 -526
rect 324 -527 325 -501
rect 429 -527 430 -501
rect 478 -558 479 -526
rect 534 -527 535 -501
rect 100 -558 101 -528
rect 163 -529 164 -501
rect 170 -558 171 -528
rect 219 -558 220 -528
rect 226 -558 227 -528
rect 268 -529 269 -501
rect 275 -558 276 -528
rect 471 -529 472 -501
rect 485 -529 486 -501
rect 534 -558 535 -528
rect 107 -531 108 -501
rect 289 -558 290 -530
rect 324 -558 325 -530
rect 390 -558 391 -530
rect 397 -558 398 -530
rect 611 -531 612 -501
rect 107 -558 108 -532
rect 149 -533 150 -501
rect 163 -558 164 -532
rect 611 -558 612 -532
rect 65 -558 66 -534
rect 149 -558 150 -534
rect 177 -535 178 -501
rect 240 -558 241 -534
rect 348 -558 349 -534
rect 443 -558 444 -534
rect 457 -558 458 -534
rect 485 -558 486 -534
rect 61 -558 62 -536
rect 177 -558 178 -536
rect 198 -558 199 -536
rect 254 -537 255 -501
rect 362 -537 363 -501
rect 450 -537 451 -501
rect 121 -558 122 -538
rect 131 -558 132 -538
rect 135 -558 136 -538
rect 156 -539 157 -501
rect 205 -558 206 -538
rect 471 -558 472 -538
rect 142 -541 143 -501
rect 233 -558 234 -540
rect 254 -558 255 -540
rect 313 -541 314 -501
rect 366 -558 367 -540
rect 408 -541 409 -501
rect 429 -558 430 -540
rect 520 -541 521 -501
rect 145 -558 146 -542
rect 632 -543 633 -501
rect 156 -558 157 -544
rect 359 -558 360 -544
rect 373 -545 374 -501
rect 411 -558 412 -544
rect 436 -545 437 -501
rect 450 -558 451 -544
rect 520 -558 521 -544
rect 583 -545 584 -501
rect 632 -558 633 -544
rect 639 -558 640 -544
rect 271 -558 272 -546
rect 583 -558 584 -546
rect 338 -549 339 -501
rect 436 -558 437 -548
rect 296 -551 297 -501
rect 338 -558 339 -550
rect 373 -558 374 -550
rect 401 -551 402 -501
rect 296 -558 297 -552
rect 317 -553 318 -501
rect 380 -553 381 -501
rect 425 -553 426 -501
rect 247 -555 248 -501
rect 317 -558 318 -554
rect 380 -558 381 -554
rect 576 -558 577 -554
rect 247 -558 248 -556
rect 268 -558 269 -556
rect 383 -558 384 -556
rect 387 -557 388 -501
rect 2 -613 3 -567
rect 93 -568 94 -566
rect 100 -568 101 -566
rect 142 -568 143 -566
rect 156 -568 157 -566
rect 240 -568 241 -566
rect 254 -568 255 -566
rect 355 -568 356 -566
rect 369 -568 370 -566
rect 464 -568 465 -566
rect 485 -568 486 -566
rect 555 -568 556 -566
rect 576 -568 577 -566
rect 611 -613 612 -567
rect 618 -568 619 -566
rect 628 -568 629 -566
rect 632 -568 633 -566
rect 632 -613 633 -567
rect 632 -568 633 -566
rect 632 -613 633 -567
rect 642 -568 643 -566
rect 653 -568 654 -566
rect 9 -613 10 -569
rect 100 -613 101 -569
rect 114 -570 115 -566
rect 149 -570 150 -566
rect 170 -570 171 -566
rect 212 -570 213 -566
rect 233 -570 234 -566
rect 268 -570 269 -566
rect 271 -570 272 -566
rect 317 -570 318 -566
rect 352 -570 353 -566
rect 590 -570 591 -566
rect 646 -570 647 -566
rect 653 -613 654 -569
rect 16 -572 17 -566
rect 103 -613 104 -571
rect 114 -613 115 -571
rect 135 -572 136 -566
rect 142 -613 143 -571
rect 205 -572 206 -566
rect 208 -613 209 -571
rect 229 -613 230 -571
rect 261 -572 262 -566
rect 404 -572 405 -566
rect 408 -572 409 -566
rect 604 -572 605 -566
rect 16 -613 17 -573
rect 310 -574 311 -566
rect 331 -613 332 -573
rect 590 -613 591 -573
rect 23 -576 24 -566
rect 79 -576 80 -566
rect 82 -576 83 -566
rect 93 -613 94 -575
rect 135 -613 136 -575
rect 257 -613 258 -575
rect 268 -613 269 -575
rect 324 -576 325 -566
rect 373 -576 374 -566
rect 576 -613 577 -575
rect 583 -576 584 -566
rect 618 -613 619 -575
rect 23 -613 24 -577
rect 191 -578 192 -566
rect 194 -578 195 -566
rect 226 -578 227 -566
rect 278 -613 279 -577
rect 317 -613 318 -577
rect 324 -613 325 -577
rect 450 -578 451 -566
rect 464 -613 465 -577
rect 471 -578 472 -566
rect 544 -613 545 -577
rect 597 -578 598 -566
rect 30 -580 31 -566
rect 380 -613 381 -579
rect 383 -580 384 -566
rect 411 -580 412 -566
rect 429 -580 430 -566
rect 432 -598 433 -579
rect 450 -613 451 -579
rect 625 -613 626 -579
rect 30 -613 31 -581
rect 72 -582 73 -566
rect 79 -613 80 -581
rect 163 -582 164 -566
rect 170 -613 171 -581
rect 184 -582 185 -566
rect 198 -582 199 -566
rect 201 -613 202 -581
rect 205 -613 206 -581
rect 408 -613 409 -581
rect 429 -613 430 -581
rect 478 -582 479 -566
rect 506 -582 507 -566
rect 597 -613 598 -581
rect 51 -584 52 -566
rect 233 -613 234 -583
rect 289 -584 290 -566
rect 289 -613 290 -583
rect 289 -584 290 -566
rect 289 -613 290 -583
rect 303 -584 304 -566
rect 334 -584 335 -566
rect 387 -584 388 -566
rect 520 -584 521 -566
rect 565 -613 566 -583
rect 604 -613 605 -583
rect 51 -613 52 -585
rect 121 -586 122 -566
rect 152 -586 153 -566
rect 163 -613 164 -585
rect 177 -586 178 -566
rect 261 -613 262 -585
rect 296 -586 297 -566
rect 303 -613 304 -585
rect 310 -613 311 -585
rect 436 -586 437 -566
rect 443 -586 444 -566
rect 478 -613 479 -585
rect 506 -613 507 -585
rect 548 -586 549 -566
rect 569 -586 570 -566
rect 583 -613 584 -585
rect 61 -613 62 -587
rect 240 -613 241 -587
rect 264 -588 265 -566
rect 436 -613 437 -587
rect 471 -613 472 -587
rect 499 -588 500 -566
rect 520 -613 521 -587
rect 534 -588 535 -566
rect 548 -613 549 -587
rect 562 -588 563 -566
rect 65 -590 66 -566
rect 296 -613 297 -589
rect 345 -613 346 -589
rect 499 -613 500 -589
rect 527 -590 528 -566
rect 569 -613 570 -589
rect 68 -613 69 -591
rect 128 -613 129 -591
rect 152 -613 153 -591
rect 338 -592 339 -566
rect 394 -592 395 -566
rect 485 -613 486 -591
rect 534 -613 535 -591
rect 541 -592 542 -566
rect 72 -613 73 -593
rect 219 -594 220 -566
rect 226 -613 227 -593
rect 282 -594 283 -566
rect 338 -613 339 -593
rect 362 -613 363 -593
rect 401 -594 402 -566
rect 513 -594 514 -566
rect 58 -596 59 -566
rect 219 -613 220 -595
rect 247 -596 248 -566
rect 394 -613 395 -595
rect 401 -613 402 -595
rect 492 -596 493 -566
rect 86 -598 87 -566
rect 348 -598 349 -566
rect 443 -613 444 -597
rect 457 -598 458 -566
rect 513 -613 514 -597
rect 86 -613 87 -599
rect 191 -613 192 -599
rect 198 -613 199 -599
rect 555 -613 556 -599
rect 107 -602 108 -566
rect 184 -613 185 -601
rect 212 -613 213 -601
rect 352 -613 353 -601
rect 492 -613 493 -601
rect 621 -602 622 -566
rect 37 -604 38 -566
rect 107 -613 108 -603
rect 121 -613 122 -603
rect 373 -613 374 -603
rect 37 -613 38 -605
rect 44 -606 45 -566
rect 156 -613 157 -605
rect 177 -613 178 -605
rect 180 -613 181 -605
rect 247 -613 248 -605
rect 282 -613 283 -605
rect 415 -606 416 -566
rect 44 -613 45 -607
rect 124 -613 125 -607
rect 348 -613 349 -607
rect 366 -613 367 -607
rect 415 -613 416 -607
rect 422 -608 423 -566
rect 359 -610 360 -566
rect 422 -613 423 -609
rect 359 -613 360 -611
rect 387 -613 388 -611
rect 2 -623 3 -621
rect 128 -623 129 -621
rect 131 -623 132 -621
rect 208 -623 209 -621
rect 212 -623 213 -621
rect 334 -623 335 -621
rect 345 -623 346 -621
rect 569 -623 570 -621
rect 625 -623 626 -621
rect 639 -678 640 -622
rect 653 -623 654 -621
rect 653 -678 654 -622
rect 653 -623 654 -621
rect 653 -678 654 -622
rect 2 -678 3 -624
rect 93 -625 94 -621
rect 100 -678 101 -624
rect 152 -625 153 -621
rect 156 -625 157 -621
rect 156 -678 157 -624
rect 156 -625 157 -621
rect 156 -678 157 -624
rect 173 -678 174 -624
rect 583 -625 584 -621
rect 632 -625 633 -621
rect 632 -678 633 -624
rect 632 -625 633 -621
rect 632 -678 633 -624
rect 9 -627 10 -621
rect 205 -627 206 -621
rect 208 -678 209 -626
rect 604 -627 605 -621
rect 9 -678 10 -628
rect 68 -629 69 -621
rect 103 -629 104 -621
rect 194 -629 195 -621
rect 201 -629 202 -621
rect 261 -629 262 -621
rect 296 -629 297 -621
rect 327 -629 328 -621
rect 334 -678 335 -628
rect 562 -678 563 -628
rect 565 -678 566 -628
rect 590 -629 591 -621
rect 16 -631 17 -621
rect 278 -631 279 -621
rect 289 -631 290 -621
rect 296 -678 297 -630
rect 313 -631 314 -621
rect 429 -631 430 -621
rect 443 -631 444 -621
rect 478 -678 479 -630
rect 499 -631 500 -621
rect 499 -678 500 -630
rect 499 -631 500 -621
rect 499 -678 500 -630
rect 513 -631 514 -621
rect 541 -678 542 -630
rect 16 -678 17 -632
rect 131 -678 132 -632
rect 184 -633 185 -621
rect 359 -678 360 -632
rect 362 -633 363 -621
rect 597 -633 598 -621
rect 23 -635 24 -621
rect 177 -635 178 -621
rect 219 -635 220 -621
rect 331 -678 332 -634
rect 348 -635 349 -621
rect 576 -635 577 -621
rect 23 -678 24 -636
rect 96 -678 97 -636
rect 107 -637 108 -621
rect 110 -669 111 -636
rect 114 -637 115 -621
rect 138 -678 139 -636
rect 170 -637 171 -621
rect 184 -678 185 -636
rect 219 -678 220 -636
rect 401 -678 402 -636
rect 415 -637 416 -621
rect 415 -678 416 -636
rect 415 -637 416 -621
rect 415 -678 416 -636
rect 443 -678 444 -636
rect 492 -637 493 -621
rect 520 -637 521 -621
rect 558 -678 559 -636
rect 30 -639 31 -621
rect 152 -678 153 -638
rect 177 -678 178 -638
rect 380 -639 381 -621
rect 429 -678 430 -638
rect 492 -678 493 -638
rect 520 -678 521 -638
rect 548 -639 549 -621
rect 30 -678 31 -640
rect 278 -678 279 -640
rect 324 -641 325 -621
rect 548 -678 549 -640
rect 37 -643 38 -621
rect 65 -643 66 -621
rect 107 -678 108 -642
rect 163 -643 164 -621
rect 222 -678 223 -642
rect 317 -643 318 -621
rect 324 -678 325 -642
rect 404 -643 405 -621
rect 460 -643 461 -621
rect 611 -643 612 -621
rect 37 -678 38 -644
rect 142 -645 143 -621
rect 226 -645 227 -621
rect 387 -645 388 -621
rect 527 -645 528 -621
rect 618 -645 619 -621
rect 44 -647 45 -621
rect 198 -647 199 -621
rect 226 -678 227 -646
rect 247 -647 248 -621
rect 257 -647 258 -621
rect 464 -647 465 -621
rect 44 -678 45 -648
rect 205 -678 206 -648
rect 240 -649 241 -621
rect 289 -678 290 -648
rect 303 -649 304 -621
rect 317 -678 318 -648
rect 338 -649 339 -621
rect 380 -678 381 -648
rect 387 -678 388 -648
rect 394 -649 395 -621
rect 436 -649 437 -621
rect 527 -678 528 -648
rect 51 -651 52 -621
rect 201 -678 202 -650
rect 247 -678 248 -650
rect 457 -651 458 -621
rect 51 -678 52 -652
rect 261 -678 262 -652
rect 275 -678 276 -652
rect 338 -678 339 -652
rect 345 -678 346 -652
rect 404 -678 405 -652
rect 408 -653 409 -621
rect 436 -678 437 -652
rect 58 -678 59 -654
rect 170 -678 171 -654
rect 282 -655 283 -621
rect 303 -678 304 -654
rect 310 -655 311 -621
rect 464 -678 465 -654
rect 61 -657 62 -621
rect 555 -657 556 -621
rect 65 -678 66 -658
rect 229 -659 230 -621
rect 268 -659 269 -621
rect 310 -678 311 -658
rect 313 -678 314 -658
rect 457 -678 458 -658
rect 513 -678 514 -658
rect 555 -678 556 -658
rect 72 -661 73 -621
rect 268 -678 269 -660
rect 352 -678 353 -660
rect 373 -661 374 -621
rect 408 -678 409 -660
rect 450 -661 451 -621
rect 72 -678 73 -662
rect 128 -678 129 -662
rect 135 -663 136 -621
rect 142 -678 143 -662
rect 180 -663 181 -621
rect 450 -678 451 -662
rect 79 -665 80 -621
rect 240 -678 241 -664
rect 355 -665 356 -621
rect 422 -665 423 -621
rect 79 -678 80 -666
rect 135 -678 136 -666
rect 191 -678 192 -666
rect 373 -678 374 -666
rect 422 -678 423 -666
rect 534 -667 535 -621
rect 163 -678 164 -668
rect 366 -669 367 -621
rect 397 -678 398 -668
rect 506 -669 507 -621
rect 534 -678 535 -668
rect 121 -671 122 -621
rect 233 -671 234 -621
rect 369 -678 370 -670
rect 471 -671 472 -621
rect 485 -671 486 -621
rect 506 -678 507 -670
rect 86 -673 87 -621
rect 233 -678 234 -672
rect 257 -678 258 -672
rect 471 -678 472 -672
rect 86 -678 87 -674
rect 149 -678 150 -674
rect 394 -678 395 -674
rect 485 -678 486 -674
rect 121 -678 122 -676
rect 212 -678 213 -676
rect 2 -688 3 -686
rect 205 -688 206 -686
rect 219 -688 220 -686
rect 285 -688 286 -686
rect 289 -745 290 -687
rect 306 -745 307 -687
rect 313 -688 314 -686
rect 415 -688 416 -686
rect 422 -745 423 -687
rect 425 -688 426 -686
rect 429 -745 430 -687
rect 450 -688 451 -686
rect 457 -688 458 -686
rect 611 -745 612 -687
rect 632 -688 633 -686
rect 639 -688 640 -686
rect 653 -688 654 -686
rect 653 -745 654 -687
rect 653 -688 654 -686
rect 653 -745 654 -687
rect 2 -745 3 -689
rect 58 -690 59 -686
rect 65 -690 66 -686
rect 65 -745 66 -689
rect 65 -690 66 -686
rect 65 -745 66 -689
rect 96 -690 97 -686
rect 173 -690 174 -686
rect 177 -690 178 -686
rect 254 -690 255 -686
rect 278 -690 279 -686
rect 296 -690 297 -686
rect 317 -690 318 -686
rect 317 -745 318 -689
rect 317 -690 318 -686
rect 317 -745 318 -689
rect 331 -690 332 -686
rect 457 -745 458 -689
rect 478 -690 479 -686
rect 583 -745 584 -689
rect 9 -692 10 -686
rect 121 -692 122 -686
rect 135 -745 136 -691
rect 156 -692 157 -686
rect 170 -745 171 -691
rect 191 -692 192 -686
rect 194 -745 195 -691
rect 226 -692 227 -686
rect 229 -745 230 -691
rect 590 -745 591 -691
rect 12 -745 13 -693
rect 394 -745 395 -693
rect 397 -694 398 -686
rect 548 -694 549 -686
rect 562 -694 563 -686
rect 663 -745 664 -693
rect 16 -696 17 -686
rect 117 -696 118 -686
rect 121 -745 122 -695
rect 180 -696 181 -686
rect 187 -696 188 -686
rect 562 -745 563 -695
rect 16 -745 17 -697
rect 93 -745 94 -697
rect 114 -698 115 -686
rect 576 -745 577 -697
rect 30 -700 31 -686
rect 128 -700 129 -686
rect 156 -745 157 -699
rect 212 -700 213 -686
rect 219 -745 220 -699
rect 261 -700 262 -686
rect 271 -745 272 -699
rect 331 -745 332 -699
rect 338 -700 339 -686
rect 597 -745 598 -699
rect 30 -745 31 -701
rect 107 -702 108 -686
rect 114 -745 115 -701
rect 478 -745 479 -701
rect 485 -702 486 -686
rect 569 -745 570 -701
rect 37 -704 38 -686
rect 257 -704 258 -686
rect 278 -745 279 -703
rect 401 -745 402 -703
rect 404 -704 405 -686
rect 555 -745 556 -703
rect 37 -745 38 -705
rect 86 -706 87 -686
rect 117 -745 118 -705
rect 296 -745 297 -705
rect 341 -745 342 -705
rect 443 -706 444 -686
rect 464 -706 465 -686
rect 548 -745 549 -705
rect 44 -708 45 -686
rect 47 -745 48 -707
rect 51 -745 52 -707
rect 261 -745 262 -707
rect 345 -708 346 -686
rect 415 -745 416 -707
rect 432 -708 433 -686
rect 506 -708 507 -686
rect 520 -708 521 -686
rect 618 -745 619 -707
rect 54 -710 55 -686
rect 240 -710 241 -686
rect 247 -710 248 -686
rect 285 -745 286 -709
rect 292 -710 293 -686
rect 506 -745 507 -709
rect 527 -710 528 -686
rect 625 -745 626 -709
rect 82 -745 83 -711
rect 212 -745 213 -711
rect 226 -745 227 -711
rect 471 -712 472 -686
rect 492 -712 493 -686
rect 604 -745 605 -711
rect 86 -745 87 -713
rect 142 -714 143 -686
rect 145 -745 146 -713
rect 527 -745 528 -713
rect 100 -716 101 -686
rect 247 -745 248 -715
rect 254 -745 255 -715
rect 373 -745 374 -715
rect 376 -716 377 -686
rect 541 -716 542 -686
rect 128 -745 129 -717
rect 184 -745 185 -717
rect 198 -718 199 -686
rect 324 -718 325 -686
rect 345 -745 346 -717
rect 366 -718 367 -686
rect 376 -745 377 -717
rect 646 -745 647 -717
rect 107 -745 108 -719
rect 198 -745 199 -719
rect 233 -720 234 -686
rect 369 -720 370 -686
rect 380 -720 381 -686
rect 632 -745 633 -719
rect 149 -722 150 -686
rect 338 -745 339 -721
rect 355 -745 356 -721
rect 450 -745 451 -721
rect 499 -722 500 -686
rect 520 -745 521 -721
rect 72 -724 73 -686
rect 499 -745 500 -723
rect 72 -745 73 -725
rect 79 -726 80 -686
rect 149 -745 150 -725
rect 310 -726 311 -686
rect 359 -726 360 -686
rect 485 -745 486 -725
rect 163 -728 164 -686
rect 240 -745 241 -727
rect 268 -728 269 -686
rect 324 -745 325 -727
rect 359 -745 360 -727
rect 534 -728 535 -686
rect 166 -745 167 -729
rect 443 -745 444 -729
rect 513 -730 514 -686
rect 534 -745 535 -729
rect 177 -745 178 -731
rect 201 -732 202 -686
rect 268 -745 269 -731
rect 639 -745 640 -731
rect 191 -745 192 -733
rect 233 -745 234 -733
rect 275 -734 276 -686
rect 541 -745 542 -733
rect 187 -745 188 -735
rect 275 -745 276 -735
rect 303 -736 304 -686
rect 492 -745 493 -735
rect 310 -745 311 -737
rect 352 -738 353 -686
rect 366 -745 367 -737
rect 656 -745 657 -737
rect 352 -745 353 -739
rect 387 -740 388 -686
rect 408 -740 409 -686
rect 464 -745 465 -739
rect 282 -745 283 -741
rect 387 -745 388 -741
rect 436 -742 437 -686
rect 513 -745 514 -741
rect 362 -745 363 -743
rect 436 -745 437 -743
rect 2 -755 3 -753
rect 163 -755 164 -753
rect 184 -818 185 -754
rect 254 -755 255 -753
rect 261 -755 262 -753
rect 362 -755 363 -753
rect 373 -755 374 -753
rect 436 -755 437 -753
rect 471 -755 472 -753
rect 625 -755 626 -753
rect 23 -757 24 -753
rect 387 -757 388 -753
rect 471 -818 472 -756
rect 541 -757 542 -753
rect 558 -818 559 -756
rect 646 -757 647 -753
rect 23 -818 24 -758
rect 100 -759 101 -753
rect 114 -759 115 -753
rect 240 -759 241 -753
rect 243 -818 244 -758
rect 296 -759 297 -753
rect 299 -818 300 -758
rect 597 -759 598 -753
rect 30 -761 31 -753
rect 103 -761 104 -753
rect 114 -818 115 -760
rect 135 -761 136 -753
rect 142 -761 143 -753
rect 604 -761 605 -753
rect 30 -818 31 -762
rect 107 -763 108 -753
rect 117 -763 118 -753
rect 254 -818 255 -762
rect 261 -818 262 -762
rect 345 -763 346 -753
rect 376 -763 377 -753
rect 583 -763 584 -753
rect 597 -818 598 -762
rect 604 -818 605 -762
rect 37 -765 38 -753
rect 149 -765 150 -753
rect 152 -765 153 -753
rect 163 -818 164 -764
rect 187 -765 188 -753
rect 394 -765 395 -753
rect 474 -765 475 -753
rect 555 -765 556 -753
rect 583 -818 584 -764
rect 611 -765 612 -753
rect 54 -818 55 -766
rect 352 -818 353 -766
rect 376 -818 377 -766
rect 618 -767 619 -753
rect 61 -769 62 -753
rect 639 -769 640 -753
rect 65 -771 66 -753
rect 229 -771 230 -753
rect 247 -771 248 -753
rect 247 -818 248 -770
rect 247 -771 248 -753
rect 247 -818 248 -770
rect 268 -771 269 -753
rect 317 -771 318 -753
rect 327 -818 328 -770
rect 415 -771 416 -753
rect 443 -771 444 -753
rect 555 -818 556 -770
rect 618 -818 619 -770
rect 660 -771 661 -753
rect 65 -818 66 -772
rect 156 -773 157 -753
rect 191 -818 192 -772
rect 338 -818 339 -772
rect 345 -818 346 -772
rect 359 -773 360 -753
rect 380 -773 381 -753
rect 513 -773 514 -753
rect 541 -818 542 -772
rect 590 -773 591 -753
rect 79 -818 80 -774
rect 548 -775 549 -753
rect 82 -777 83 -753
rect 492 -777 493 -753
rect 44 -818 45 -778
rect 82 -818 83 -778
rect 86 -779 87 -753
rect 205 -779 206 -753
rect 208 -779 209 -753
rect 576 -779 577 -753
rect 96 -818 97 -780
rect 100 -818 101 -780
rect 107 -818 108 -780
rect 121 -781 122 -753
rect 145 -781 146 -753
rect 170 -781 171 -753
rect 198 -781 199 -753
rect 478 -781 479 -753
rect 93 -783 94 -753
rect 121 -818 122 -782
rect 149 -818 150 -782
rect 205 -818 206 -782
rect 219 -783 220 -753
rect 226 -818 227 -782
rect 268 -818 269 -782
rect 310 -783 311 -753
rect 331 -783 332 -753
rect 513 -818 514 -782
rect 156 -818 157 -784
rect 177 -785 178 -753
rect 219 -818 220 -784
rect 653 -785 654 -753
rect 58 -787 59 -753
rect 177 -818 178 -786
rect 275 -787 276 -753
rect 324 -787 325 -753
rect 359 -818 360 -786
rect 366 -787 367 -753
rect 373 -818 374 -786
rect 590 -818 591 -786
rect 58 -818 59 -788
rect 72 -789 73 -753
rect 170 -818 171 -788
rect 282 -818 283 -788
rect 285 -818 286 -788
rect 499 -789 500 -753
rect 72 -818 73 -790
rect 128 -791 129 -753
rect 275 -818 276 -790
rect 632 -791 633 -753
rect 278 -793 279 -753
rect 464 -793 465 -753
rect 499 -818 500 -792
rect 520 -793 521 -753
rect 198 -818 199 -794
rect 278 -818 279 -794
rect 289 -795 290 -753
rect 408 -795 409 -753
rect 411 -795 412 -753
rect 548 -818 549 -794
rect 212 -797 213 -753
rect 408 -818 409 -796
rect 415 -818 416 -796
rect 527 -797 528 -753
rect 152 -818 153 -798
rect 212 -818 213 -798
rect 233 -799 234 -753
rect 289 -818 290 -798
rect 303 -818 304 -798
rect 331 -818 332 -798
rect 380 -818 381 -798
rect 429 -799 430 -753
rect 443 -818 444 -798
rect 534 -799 535 -753
rect 51 -801 52 -753
rect 233 -818 234 -800
rect 310 -818 311 -800
rect 506 -801 507 -753
rect 527 -818 528 -800
rect 562 -801 563 -753
rect 320 -818 321 -802
rect 366 -818 367 -802
rect 387 -818 388 -802
rect 520 -818 521 -802
rect 562 -818 563 -802
rect 569 -803 570 -753
rect 341 -805 342 -753
rect 506 -818 507 -804
rect 341 -818 342 -806
rect 436 -818 437 -806
rect 450 -807 451 -753
rect 576 -818 577 -806
rect 390 -818 391 -808
rect 492 -818 493 -808
rect 394 -818 395 -810
rect 401 -811 402 -753
rect 422 -811 423 -753
rect 429 -818 430 -810
rect 450 -818 451 -810
rect 485 -811 486 -753
rect 313 -818 314 -812
rect 422 -818 423 -812
rect 457 -813 458 -753
rect 485 -818 486 -812
rect 457 -818 458 -814
rect 537 -818 538 -814
rect 464 -818 465 -816
rect 569 -818 570 -816
rect 9 -861 10 -827
rect 33 -861 34 -827
rect 40 -828 41 -826
rect 96 -828 97 -826
rect 107 -828 108 -826
rect 135 -828 136 -826
rect 149 -861 150 -827
rect 229 -861 230 -827
rect 233 -828 234 -826
rect 373 -828 374 -826
rect 387 -861 388 -827
rect 408 -828 409 -826
rect 415 -828 416 -826
rect 415 -861 416 -827
rect 415 -828 416 -826
rect 415 -861 416 -827
rect 425 -861 426 -827
rect 492 -828 493 -826
rect 513 -861 514 -827
rect 562 -828 563 -826
rect 572 -828 573 -826
rect 618 -828 619 -826
rect 16 -861 17 -829
rect 37 -861 38 -829
rect 54 -830 55 -826
rect 471 -830 472 -826
rect 478 -830 479 -826
rect 541 -830 542 -826
rect 555 -861 556 -829
rect 590 -830 591 -826
rect 30 -832 31 -826
rect 93 -832 94 -826
rect 107 -861 108 -831
rect 184 -832 185 -826
rect 194 -861 195 -831
rect 212 -832 213 -826
rect 222 -861 223 -831
rect 285 -832 286 -826
rect 292 -861 293 -831
rect 492 -861 493 -831
rect 534 -861 535 -831
rect 583 -832 584 -826
rect 58 -834 59 -826
rect 86 -834 87 -826
rect 89 -834 90 -826
rect 100 -834 101 -826
rect 114 -834 115 -826
rect 145 -834 146 -826
rect 170 -834 171 -826
rect 324 -861 325 -833
rect 334 -834 335 -826
rect 548 -834 549 -826
rect 562 -861 563 -833
rect 576 -834 577 -826
rect 23 -836 24 -826
rect 170 -861 171 -835
rect 180 -861 181 -835
rect 240 -861 241 -835
rect 247 -836 248 -826
rect 250 -844 251 -835
rect 268 -836 269 -826
rect 317 -836 318 -826
rect 320 -836 321 -826
rect 436 -836 437 -826
rect 464 -836 465 -826
rect 464 -861 465 -835
rect 464 -836 465 -826
rect 464 -861 465 -835
rect 478 -861 479 -835
rect 506 -836 507 -826
rect 548 -861 549 -835
rect 604 -836 605 -826
rect 23 -861 24 -837
rect 44 -838 45 -826
rect 51 -838 52 -826
rect 100 -861 101 -837
rect 114 -861 115 -837
rect 198 -838 199 -826
rect 226 -838 227 -826
rect 275 -838 276 -826
rect 303 -838 304 -826
rect 373 -861 374 -837
rect 394 -838 395 -826
rect 394 -861 395 -837
rect 394 -838 395 -826
rect 394 -861 395 -837
rect 401 -838 402 -826
rect 450 -838 451 -826
rect 485 -838 486 -826
rect 485 -861 486 -837
rect 485 -838 486 -826
rect 485 -861 486 -837
rect 499 -838 500 -826
rect 506 -861 507 -837
rect 51 -861 52 -839
rect 61 -861 62 -839
rect 65 -840 66 -826
rect 201 -861 202 -839
rect 247 -861 248 -839
rect 289 -840 290 -826
rect 317 -861 318 -839
rect 499 -861 500 -839
rect 65 -861 66 -841
rect 163 -842 164 -826
rect 173 -861 174 -841
rect 268 -861 269 -841
rect 320 -861 321 -841
rect 408 -861 409 -841
rect 422 -842 423 -826
rect 471 -861 472 -841
rect 72 -844 73 -826
rect 128 -844 129 -826
rect 135 -861 136 -843
rect 215 -861 216 -843
rect 289 -861 290 -843
rect 338 -844 339 -826
rect 380 -844 381 -826
rect 404 -844 405 -826
rect 520 -844 521 -826
rect 72 -861 73 -845
rect 82 -846 83 -826
rect 86 -861 87 -845
rect 219 -846 220 -826
rect 254 -846 255 -826
rect 338 -861 339 -845
rect 345 -846 346 -826
rect 516 -861 517 -845
rect 93 -861 94 -847
rect 142 -861 143 -847
rect 163 -861 164 -847
rect 282 -861 283 -847
rect 348 -861 349 -847
rect 457 -848 458 -826
rect 121 -850 122 -826
rect 152 -850 153 -826
rect 177 -850 178 -826
rect 275 -861 276 -849
rect 352 -861 353 -849
rect 359 -850 360 -826
rect 366 -850 367 -826
rect 366 -861 367 -849
rect 366 -850 367 -826
rect 366 -861 367 -849
rect 376 -850 377 -826
rect 401 -861 402 -849
rect 429 -850 430 -826
rect 429 -861 430 -849
rect 429 -850 430 -826
rect 429 -861 430 -849
rect 436 -861 437 -849
rect 443 -850 444 -826
rect 121 -861 122 -851
rect 156 -852 157 -826
rect 184 -861 185 -851
rect 191 -852 192 -826
rect 198 -861 199 -851
rect 310 -861 311 -851
rect 331 -852 332 -826
rect 443 -861 444 -851
rect 2 -861 3 -853
rect 191 -861 192 -853
rect 205 -854 206 -826
rect 254 -861 255 -853
rect 261 -854 262 -826
rect 303 -861 304 -853
rect 345 -861 346 -853
rect 359 -861 360 -853
rect 128 -861 129 -855
rect 278 -856 279 -826
rect 296 -856 297 -826
rect 331 -861 332 -855
rect 355 -856 356 -826
rect 527 -856 528 -826
rect 156 -861 157 -857
rect 205 -861 206 -857
rect 226 -861 227 -857
rect 457 -861 458 -857
rect 520 -861 521 -857
rect 527 -861 528 -857
rect 233 -861 234 -859
rect 261 -861 262 -859
rect 296 -861 297 -859
rect 380 -861 381 -859
rect 2 -871 3 -869
rect 135 -871 136 -869
rect 152 -916 153 -870
rect 387 -871 388 -869
rect 425 -871 426 -869
rect 499 -871 500 -869
rect 516 -871 517 -869
rect 544 -871 545 -869
rect 2 -916 3 -872
rect 114 -873 115 -869
rect 121 -873 122 -869
rect 173 -873 174 -869
rect 205 -873 206 -869
rect 233 -873 234 -869
rect 247 -873 248 -869
rect 320 -873 321 -869
rect 345 -916 346 -872
rect 401 -873 402 -869
rect 443 -873 444 -869
rect 548 -873 549 -869
rect 9 -875 10 -869
rect 44 -875 45 -869
rect 47 -875 48 -869
rect 103 -916 104 -874
rect 135 -916 136 -874
rect 149 -875 150 -869
rect 156 -875 157 -869
rect 233 -916 234 -874
rect 240 -875 241 -869
rect 247 -916 248 -874
rect 261 -916 262 -874
rect 296 -875 297 -869
rect 299 -916 300 -874
rect 387 -916 388 -874
rect 401 -916 402 -874
rect 450 -875 451 -869
rect 453 -875 454 -869
rect 485 -875 486 -869
rect 492 -875 493 -869
rect 492 -916 493 -874
rect 492 -875 493 -869
rect 492 -916 493 -874
rect 520 -875 521 -869
rect 534 -916 535 -874
rect 537 -875 538 -869
rect 541 -916 542 -874
rect 548 -916 549 -874
rect 555 -875 556 -869
rect 16 -877 17 -869
rect 30 -877 31 -869
rect 44 -916 45 -876
rect 51 -877 52 -869
rect 54 -916 55 -876
rect 124 -916 125 -876
rect 142 -916 143 -876
rect 240 -916 241 -876
rect 268 -877 269 -869
rect 499 -916 500 -876
rect 520 -916 521 -876
rect 530 -916 531 -876
rect 16 -916 17 -878
rect 40 -879 41 -869
rect 61 -879 62 -869
rect 72 -879 73 -869
rect 79 -879 80 -869
rect 128 -879 129 -869
rect 173 -916 174 -878
rect 373 -879 374 -869
rect 376 -879 377 -869
rect 464 -879 465 -869
rect 485 -916 486 -878
rect 506 -879 507 -869
rect 527 -879 528 -869
rect 562 -879 563 -869
rect 23 -881 24 -869
rect 37 -881 38 -869
rect 65 -881 66 -869
rect 163 -881 164 -869
rect 191 -881 192 -869
rect 464 -916 465 -880
rect 478 -881 479 -869
rect 506 -916 507 -880
rect 23 -916 24 -882
rect 131 -916 132 -882
rect 163 -916 164 -882
rect 184 -883 185 -869
rect 208 -883 209 -869
rect 338 -883 339 -869
rect 348 -883 349 -869
rect 352 -883 353 -869
rect 380 -883 381 -869
rect 436 -883 437 -869
rect 457 -883 458 -869
rect 457 -916 458 -882
rect 457 -883 458 -869
rect 457 -916 458 -882
rect 68 -916 69 -884
rect 86 -885 87 -869
rect 93 -885 94 -869
rect 201 -916 202 -884
rect 212 -916 213 -884
rect 275 -885 276 -869
rect 282 -885 283 -869
rect 373 -916 374 -884
rect 422 -916 423 -884
rect 527 -916 528 -884
rect 79 -916 80 -886
rect 177 -916 178 -886
rect 194 -916 195 -886
rect 338 -916 339 -886
rect 352 -916 353 -886
rect 366 -887 367 -869
rect 86 -916 87 -888
rect 107 -889 108 -869
rect 121 -916 122 -888
rect 184 -916 185 -888
rect 198 -916 199 -888
rect 380 -916 381 -888
rect 96 -916 97 -890
rect 149 -916 150 -890
rect 219 -891 220 -869
rect 268 -916 269 -890
rect 275 -916 276 -890
rect 289 -891 290 -869
rect 292 -891 293 -869
rect 415 -891 416 -869
rect 100 -893 101 -869
rect 156 -916 157 -892
rect 191 -916 192 -892
rect 219 -916 220 -892
rect 222 -893 223 -869
rect 366 -916 367 -892
rect 415 -916 416 -892
rect 429 -893 430 -869
rect 100 -916 101 -894
rect 114 -916 115 -894
rect 226 -895 227 -869
rect 324 -895 325 -869
rect 331 -895 332 -869
rect 436 -916 437 -894
rect 37 -916 38 -896
rect 331 -916 332 -896
rect 408 -897 409 -869
rect 429 -916 430 -896
rect 229 -916 230 -898
rect 254 -899 255 -869
rect 282 -916 283 -898
rect 513 -899 514 -869
rect 208 -916 209 -900
rect 513 -916 514 -900
rect 243 -916 244 -902
rect 478 -916 479 -902
rect 254 -916 255 -904
rect 289 -916 290 -904
rect 292 -916 293 -904
rect 471 -905 472 -869
rect 303 -907 304 -869
rect 313 -916 314 -906
rect 317 -916 318 -906
rect 359 -907 360 -869
rect 394 -907 395 -869
rect 408 -916 409 -906
rect 65 -916 66 -908
rect 394 -916 395 -908
rect 306 -916 307 -910
rect 446 -916 447 -910
rect 310 -913 311 -869
rect 450 -916 451 -912
rect 324 -916 325 -914
rect 471 -916 472 -914
rect 9 -926 10 -924
rect 394 -926 395 -924
rect 429 -926 430 -924
rect 443 -969 444 -925
rect 450 -926 451 -924
rect 471 -969 472 -925
rect 474 -926 475 -924
rect 485 -926 486 -924
rect 506 -926 507 -924
rect 509 -969 510 -925
rect 530 -926 531 -924
rect 548 -926 549 -924
rect 16 -928 17 -924
rect 30 -928 31 -924
rect 37 -969 38 -927
rect 170 -928 171 -924
rect 173 -928 174 -924
rect 481 -969 482 -927
rect 485 -969 486 -927
rect 520 -928 521 -924
rect 23 -930 24 -924
rect 72 -930 73 -924
rect 79 -930 80 -924
rect 145 -969 146 -929
rect 149 -969 150 -929
rect 331 -930 332 -924
rect 359 -930 360 -924
rect 478 -930 479 -924
rect 506 -969 507 -929
rect 520 -969 521 -929
rect 23 -969 24 -931
rect 117 -969 118 -931
rect 163 -932 164 -924
rect 198 -932 199 -924
rect 201 -969 202 -931
rect 387 -932 388 -924
rect 415 -932 416 -924
rect 429 -969 430 -931
rect 450 -969 451 -931
rect 492 -932 493 -924
rect 44 -969 45 -933
rect 124 -934 125 -924
rect 184 -934 185 -924
rect 247 -934 248 -924
rect 264 -969 265 -933
rect 436 -934 437 -924
rect 457 -934 458 -924
rect 457 -969 458 -933
rect 457 -934 458 -924
rect 457 -969 458 -933
rect 478 -969 479 -933
rect 541 -934 542 -924
rect 54 -969 55 -935
rect 198 -969 199 -935
rect 208 -936 209 -924
rect 212 -936 213 -924
rect 226 -969 227 -935
rect 422 -936 423 -924
rect 436 -969 437 -935
rect 499 -936 500 -924
rect 58 -938 59 -924
rect 86 -938 87 -924
rect 93 -938 94 -924
rect 240 -938 241 -924
rect 268 -938 269 -924
rect 271 -942 272 -937
rect 285 -969 286 -937
rect 383 -969 384 -937
rect 387 -969 388 -937
rect 401 -938 402 -924
rect 499 -969 500 -937
rect 534 -938 535 -924
rect 58 -969 59 -939
rect 142 -940 143 -924
rect 177 -940 178 -924
rect 240 -969 241 -939
rect 268 -969 269 -939
rect 324 -940 325 -924
rect 345 -940 346 -924
rect 415 -969 416 -939
rect 2 -942 3 -924
rect 142 -969 143 -941
rect 152 -942 153 -924
rect 177 -969 178 -941
rect 187 -942 188 -924
rect 212 -969 213 -941
rect 233 -942 234 -924
rect 247 -969 248 -941
rect 324 -969 325 -941
rect 338 -942 339 -924
rect 345 -969 346 -941
rect 359 -969 360 -941
rect 366 -942 367 -924
rect 373 -942 374 -924
rect 401 -969 402 -941
rect 30 -969 31 -943
rect 233 -969 234 -943
rect 243 -944 244 -924
rect 366 -969 367 -943
rect 373 -969 374 -943
rect 467 -969 468 -943
rect 72 -969 73 -945
rect 254 -946 255 -924
rect 299 -969 300 -945
rect 317 -946 318 -924
rect 320 -969 321 -945
rect 394 -969 395 -945
rect 79 -969 80 -947
rect 110 -948 111 -924
rect 114 -948 115 -924
rect 121 -969 122 -947
rect 187 -969 188 -947
rect 464 -948 465 -924
rect 68 -969 69 -949
rect 464 -969 465 -949
rect 86 -969 87 -951
rect 310 -952 311 -924
rect 338 -969 339 -951
rect 411 -969 412 -951
rect 93 -969 94 -953
rect 184 -969 185 -953
rect 191 -969 192 -953
rect 205 -969 206 -953
rect 208 -969 209 -953
rect 513 -954 514 -924
rect 96 -956 97 -924
rect 289 -956 290 -924
rect 303 -956 304 -924
rect 331 -969 332 -955
rect 362 -956 363 -924
rect 408 -956 409 -924
rect 100 -958 101 -924
rect 156 -958 157 -924
rect 194 -958 195 -924
rect 219 -958 220 -924
rect 254 -969 255 -957
rect 261 -958 262 -924
rect 282 -958 283 -924
rect 303 -969 304 -957
rect 306 -958 307 -924
rect 352 -958 353 -924
rect 100 -969 101 -959
rect 152 -969 153 -959
rect 170 -969 171 -959
rect 261 -969 262 -959
rect 289 -969 290 -959
rect 296 -969 297 -959
rect 310 -969 311 -959
rect 380 -960 381 -924
rect 110 -969 111 -961
rect 114 -969 115 -961
rect 128 -962 129 -924
rect 282 -969 283 -961
rect 352 -969 353 -961
rect 492 -969 493 -961
rect 135 -964 136 -924
rect 156 -969 157 -963
rect 219 -969 220 -963
rect 275 -964 276 -924
rect 65 -969 66 -965
rect 275 -969 276 -965
rect 135 -969 136 -967
rect 166 -969 167 -967
rect 16 -1010 17 -978
rect 79 -979 80 -977
rect 107 -979 108 -977
rect 187 -1010 188 -978
rect 219 -979 220 -977
rect 275 -979 276 -977
rect 292 -1010 293 -978
rect 324 -979 325 -977
rect 331 -979 332 -977
rect 485 -979 486 -977
rect 520 -979 521 -977
rect 527 -1010 528 -978
rect 23 -981 24 -977
rect 264 -981 265 -977
rect 320 -981 321 -977
rect 401 -981 402 -977
rect 408 -1010 409 -980
rect 432 -1010 433 -980
rect 464 -981 465 -977
rect 499 -981 500 -977
rect 26 -1010 27 -982
rect 37 -983 38 -977
rect 51 -1010 52 -982
rect 135 -983 136 -977
rect 142 -983 143 -977
rect 142 -1010 143 -982
rect 142 -983 143 -977
rect 142 -1010 143 -982
rect 156 -983 157 -977
rect 208 -983 209 -977
rect 247 -983 248 -977
rect 247 -1010 248 -982
rect 247 -983 248 -977
rect 247 -1010 248 -982
rect 261 -983 262 -977
rect 345 -983 346 -977
rect 352 -983 353 -977
rect 471 -983 472 -977
rect 478 -983 479 -977
rect 478 -1010 479 -982
rect 478 -983 479 -977
rect 478 -1010 479 -982
rect 30 -985 31 -977
rect 229 -985 230 -977
rect 271 -1010 272 -984
rect 352 -1010 353 -984
rect 380 -985 381 -977
rect 443 -985 444 -977
rect 446 -1010 447 -984
rect 464 -1010 465 -984
rect 471 -1010 472 -984
rect 492 -985 493 -977
rect 37 -1010 38 -986
rect 131 -987 132 -977
rect 135 -1010 136 -986
rect 191 -987 192 -977
rect 208 -1010 209 -986
rect 299 -987 300 -977
rect 303 -987 304 -977
rect 345 -1010 346 -986
rect 411 -987 412 -977
rect 429 -987 430 -977
rect 58 -989 59 -977
rect 128 -989 129 -977
rect 131 -1010 132 -988
rect 212 -989 213 -977
rect 229 -1010 230 -988
rect 254 -989 255 -977
rect 278 -989 279 -977
rect 401 -1010 402 -988
rect 422 -989 423 -977
rect 457 -989 458 -977
rect 58 -1010 59 -990
rect 100 -991 101 -977
rect 107 -1010 108 -990
rect 121 -991 122 -977
rect 128 -1010 129 -990
rect 198 -991 199 -977
rect 212 -1010 213 -990
rect 289 -991 290 -977
rect 296 -1010 297 -990
rect 380 -1010 381 -990
rect 390 -1010 391 -990
rect 422 -1010 423 -990
rect 429 -1010 430 -990
rect 509 -991 510 -977
rect 65 -993 66 -977
rect 114 -1010 115 -992
rect 121 -1010 122 -992
rect 184 -993 185 -977
rect 191 -1010 192 -992
rect 261 -1010 262 -992
rect 299 -1010 300 -992
rect 310 -993 311 -977
rect 324 -1010 325 -992
rect 415 -993 416 -977
rect 443 -1010 444 -992
rect 457 -1010 458 -992
rect 65 -1010 66 -994
rect 117 -995 118 -977
rect 156 -1010 157 -994
rect 170 -995 171 -977
rect 173 -1010 174 -994
rect 201 -995 202 -977
rect 233 -1010 234 -994
rect 289 -1010 290 -994
rect 303 -1010 304 -994
rect 338 -995 339 -977
rect 394 -995 395 -977
rect 415 -1010 416 -994
rect 68 -997 69 -977
rect 93 -997 94 -977
rect 100 -1010 101 -996
rect 117 -1010 118 -996
rect 149 -1010 150 -996
rect 170 -1010 171 -996
rect 177 -997 178 -977
rect 226 -1010 227 -996
rect 240 -997 241 -977
rect 310 -1010 311 -996
rect 338 -1010 339 -996
rect 373 -997 374 -977
rect 394 -1010 395 -996
rect 436 -997 437 -977
rect 30 -1010 31 -998
rect 68 -1010 69 -998
rect 72 -999 73 -977
rect 219 -1010 220 -998
rect 236 -1010 237 -998
rect 240 -1010 241 -998
rect 366 -999 367 -977
rect 373 -1010 374 -998
rect 436 -1010 437 -998
rect 450 -999 451 -977
rect 72 -1010 73 -1000
rect 86 -1001 87 -977
rect 110 -1001 111 -977
rect 359 -1001 360 -977
rect 79 -1010 80 -1002
rect 96 -1010 97 -1002
rect 163 -1010 164 -1002
rect 205 -1010 206 -1002
rect 317 -1010 318 -1002
rect 366 -1010 367 -1002
rect 177 -1010 178 -1004
rect 282 -1010 283 -1004
rect 359 -1010 360 -1004
rect 387 -1005 388 -977
rect 198 -1010 199 -1006
rect 331 -1010 332 -1006
rect 201 -1010 202 -1008
rect 254 -1010 255 -1008
rect 268 -1009 269 -977
rect 387 -1010 388 -1008
rect 30 -1020 31 -1018
rect 47 -1020 48 -1018
rect 51 -1020 52 -1018
rect 201 -1020 202 -1018
rect 208 -1020 209 -1018
rect 219 -1020 220 -1018
rect 247 -1020 248 -1018
rect 268 -1020 269 -1018
rect 278 -1020 279 -1018
rect 338 -1020 339 -1018
rect 355 -1047 356 -1019
rect 380 -1020 381 -1018
rect 415 -1020 416 -1018
rect 415 -1047 416 -1019
rect 415 -1020 416 -1018
rect 415 -1047 416 -1019
rect 422 -1020 423 -1018
rect 422 -1047 423 -1019
rect 422 -1020 423 -1018
rect 422 -1047 423 -1019
rect 436 -1020 437 -1018
rect 443 -1020 444 -1018
rect 453 -1020 454 -1018
rect 471 -1020 472 -1018
rect 478 -1020 479 -1018
rect 478 -1047 479 -1019
rect 478 -1020 479 -1018
rect 478 -1047 479 -1019
rect 523 -1020 524 -1018
rect 527 -1020 528 -1018
rect 58 -1022 59 -1018
rect 96 -1022 97 -1018
rect 114 -1022 115 -1018
rect 236 -1047 237 -1021
rect 240 -1022 241 -1018
rect 268 -1047 269 -1021
rect 289 -1047 290 -1021
rect 394 -1022 395 -1018
rect 443 -1047 444 -1021
rect 450 -1047 451 -1021
rect 453 -1047 454 -1021
rect 464 -1022 465 -1018
rect 516 -1047 517 -1021
rect 523 -1047 524 -1021
rect 16 -1024 17 -1018
rect 114 -1047 115 -1023
rect 121 -1024 122 -1018
rect 194 -1024 195 -1018
rect 205 -1047 206 -1023
rect 240 -1047 241 -1023
rect 247 -1047 248 -1023
rect 282 -1047 283 -1023
rect 296 -1047 297 -1023
rect 303 -1024 304 -1018
rect 310 -1024 311 -1018
rect 310 -1047 311 -1023
rect 310 -1024 311 -1018
rect 310 -1047 311 -1023
rect 324 -1024 325 -1018
rect 334 -1047 335 -1023
rect 359 -1024 360 -1018
rect 366 -1047 367 -1023
rect 369 -1024 370 -1018
rect 401 -1024 402 -1018
rect 457 -1024 458 -1018
rect 457 -1047 458 -1023
rect 457 -1024 458 -1018
rect 457 -1047 458 -1023
rect 520 -1024 521 -1018
rect 527 -1047 528 -1023
rect 65 -1047 66 -1025
rect 79 -1026 80 -1018
rect 86 -1026 87 -1018
rect 103 -1047 104 -1025
rect 107 -1026 108 -1018
rect 121 -1047 122 -1025
rect 142 -1026 143 -1018
rect 166 -1047 167 -1025
rect 177 -1026 178 -1018
rect 219 -1047 220 -1025
rect 229 -1026 230 -1018
rect 394 -1047 395 -1025
rect 72 -1028 73 -1018
rect 128 -1047 129 -1027
rect 135 -1028 136 -1018
rect 177 -1047 178 -1027
rect 184 -1028 185 -1018
rect 201 -1047 202 -1027
rect 208 -1047 209 -1027
rect 212 -1028 213 -1018
rect 215 -1047 216 -1027
rect 303 -1047 304 -1027
rect 324 -1047 325 -1027
rect 327 -1028 328 -1018
rect 380 -1047 381 -1027
rect 408 -1028 409 -1018
rect 72 -1047 73 -1029
rect 89 -1030 90 -1018
rect 93 -1047 94 -1029
rect 100 -1030 101 -1018
rect 107 -1047 108 -1029
rect 292 -1030 293 -1018
rect 387 -1030 388 -1018
rect 408 -1047 409 -1029
rect 86 -1047 87 -1031
rect 117 -1032 118 -1018
rect 135 -1047 136 -1031
rect 149 -1032 150 -1018
rect 156 -1032 157 -1018
rect 191 -1047 192 -1031
rect 212 -1047 213 -1031
rect 359 -1047 360 -1031
rect 37 -1034 38 -1018
rect 149 -1047 150 -1033
rect 163 -1034 164 -1018
rect 184 -1047 185 -1033
rect 187 -1034 188 -1018
rect 254 -1034 255 -1018
rect 261 -1034 262 -1018
rect 338 -1047 339 -1033
rect 117 -1047 118 -1035
rect 226 -1036 227 -1018
rect 233 -1036 234 -1018
rect 292 -1047 293 -1035
rect 331 -1036 332 -1018
rect 387 -1047 388 -1035
rect 170 -1047 171 -1037
rect 229 -1047 230 -1037
rect 250 -1047 251 -1037
rect 345 -1038 346 -1018
rect 226 -1047 227 -1039
rect 373 -1040 374 -1018
rect 261 -1047 262 -1041
rect 275 -1042 276 -1018
rect 285 -1042 286 -1018
rect 401 -1047 402 -1041
rect 275 -1047 276 -1043
rect 317 -1044 318 -1018
rect 345 -1047 346 -1043
rect 352 -1044 353 -1018
rect 373 -1047 374 -1043
rect 429 -1047 430 -1043
rect 254 -1047 255 -1045
rect 317 -1047 318 -1045
rect 51 -1092 52 -1056
rect 117 -1057 118 -1055
rect 121 -1057 122 -1055
rect 121 -1092 122 -1056
rect 121 -1057 122 -1055
rect 121 -1092 122 -1056
rect 128 -1057 129 -1055
rect 180 -1092 181 -1056
rect 201 -1057 202 -1055
rect 303 -1057 304 -1055
rect 320 -1092 321 -1056
rect 380 -1057 381 -1055
rect 429 -1057 430 -1055
rect 436 -1092 437 -1056
rect 457 -1057 458 -1055
rect 464 -1092 465 -1056
rect 478 -1057 479 -1055
rect 478 -1092 479 -1056
rect 478 -1057 479 -1055
rect 478 -1092 479 -1056
rect 520 -1057 521 -1055
rect 527 -1057 528 -1055
rect 61 -1092 62 -1058
rect 89 -1059 90 -1055
rect 93 -1059 94 -1055
rect 103 -1059 104 -1055
rect 107 -1059 108 -1055
rect 254 -1059 255 -1055
rect 334 -1059 335 -1055
rect 373 -1059 374 -1055
rect 408 -1059 409 -1055
rect 429 -1092 430 -1058
rect 65 -1061 66 -1055
rect 79 -1061 80 -1055
rect 93 -1092 94 -1060
rect 149 -1061 150 -1055
rect 152 -1061 153 -1055
rect 261 -1061 262 -1055
rect 345 -1061 346 -1055
rect 345 -1092 346 -1060
rect 345 -1061 346 -1055
rect 345 -1092 346 -1060
rect 359 -1061 360 -1055
rect 362 -1061 363 -1055
rect 373 -1092 374 -1060
rect 380 -1092 381 -1060
rect 408 -1092 409 -1060
rect 415 -1061 416 -1055
rect 65 -1092 66 -1062
rect 131 -1092 132 -1062
rect 135 -1063 136 -1055
rect 159 -1063 160 -1055
rect 163 -1063 164 -1055
rect 166 -1077 167 -1062
rect 177 -1063 178 -1055
rect 208 -1063 209 -1055
rect 212 -1063 213 -1055
rect 275 -1063 276 -1055
rect 359 -1092 360 -1062
rect 366 -1063 367 -1055
rect 72 -1065 73 -1055
rect 110 -1092 111 -1064
rect 114 -1065 115 -1055
rect 114 -1092 115 -1064
rect 114 -1065 115 -1055
rect 114 -1092 115 -1064
rect 135 -1092 136 -1064
rect 299 -1092 300 -1064
rect 366 -1092 367 -1064
rect 401 -1065 402 -1055
rect 75 -1092 76 -1066
rect 107 -1092 108 -1066
rect 145 -1067 146 -1055
rect 215 -1067 216 -1055
rect 219 -1067 220 -1055
rect 222 -1092 223 -1066
rect 226 -1092 227 -1066
rect 247 -1067 248 -1055
rect 250 -1067 251 -1055
rect 387 -1067 388 -1055
rect 394 -1067 395 -1055
rect 401 -1092 402 -1066
rect 100 -1092 101 -1068
rect 142 -1069 143 -1055
rect 149 -1092 150 -1068
rect 233 -1092 234 -1068
rect 236 -1069 237 -1055
rect 422 -1092 423 -1068
rect 156 -1092 157 -1070
rect 205 -1071 206 -1055
rect 219 -1092 220 -1070
rect 331 -1092 332 -1070
rect 163 -1092 164 -1072
rect 177 -1092 178 -1072
rect 198 -1092 199 -1072
rect 236 -1092 237 -1072
rect 352 -1092 353 -1072
rect 184 -1075 185 -1055
rect 212 -1092 213 -1074
rect 240 -1075 241 -1055
rect 240 -1092 241 -1074
rect 240 -1075 241 -1055
rect 240 -1092 241 -1074
rect 247 -1092 248 -1074
rect 292 -1075 293 -1055
rect 306 -1092 307 -1074
rect 387 -1092 388 -1074
rect 191 -1077 192 -1055
rect 205 -1092 206 -1076
rect 254 -1092 255 -1076
rect 268 -1077 269 -1055
rect 275 -1092 276 -1076
rect 317 -1077 318 -1055
rect 362 -1092 363 -1076
rect 394 -1092 395 -1076
rect 142 -1092 143 -1078
rect 317 -1092 318 -1078
rect 261 -1092 262 -1080
rect 289 -1081 290 -1055
rect 268 -1092 269 -1082
rect 282 -1083 283 -1055
rect 289 -1092 290 -1082
rect 338 -1083 339 -1055
rect 282 -1092 283 -1084
rect 390 -1092 391 -1084
rect 324 -1087 325 -1055
rect 338 -1092 339 -1086
rect 310 -1089 311 -1055
rect 324 -1092 325 -1088
rect 296 -1091 297 -1055
rect 310 -1092 311 -1090
rect 30 -1129 31 -1101
rect 93 -1102 94 -1100
rect 100 -1102 101 -1100
rect 110 -1102 111 -1100
rect 114 -1102 115 -1100
rect 222 -1102 223 -1100
rect 226 -1102 227 -1100
rect 443 -1129 444 -1101
rect 460 -1102 461 -1100
rect 464 -1102 465 -1100
rect 478 -1102 479 -1100
rect 478 -1129 479 -1101
rect 478 -1102 479 -1100
rect 478 -1129 479 -1101
rect 37 -1129 38 -1103
rect 236 -1104 237 -1100
rect 254 -1104 255 -1100
rect 299 -1104 300 -1100
rect 306 -1104 307 -1100
rect 345 -1104 346 -1100
rect 352 -1104 353 -1100
rect 418 -1104 419 -1100
rect 422 -1104 423 -1100
rect 436 -1129 437 -1103
rect 51 -1106 52 -1100
rect 89 -1106 90 -1100
rect 100 -1129 101 -1105
rect 114 -1129 115 -1105
rect 121 -1106 122 -1100
rect 138 -1106 139 -1100
rect 142 -1106 143 -1100
rect 177 -1129 178 -1105
rect 184 -1106 185 -1100
rect 247 -1106 248 -1100
rect 254 -1129 255 -1105
rect 352 -1129 353 -1105
rect 359 -1106 360 -1100
rect 373 -1106 374 -1100
rect 387 -1106 388 -1100
rect 408 -1106 409 -1100
rect 415 -1106 416 -1100
rect 429 -1106 430 -1100
rect 54 -1129 55 -1107
rect 58 -1129 59 -1107
rect 65 -1108 66 -1100
rect 187 -1108 188 -1100
rect 219 -1129 220 -1107
rect 303 -1108 304 -1100
rect 317 -1129 318 -1107
rect 338 -1108 339 -1100
rect 345 -1129 346 -1107
rect 359 -1129 360 -1107
rect 362 -1129 363 -1107
rect 366 -1108 367 -1100
rect 380 -1108 381 -1100
rect 408 -1129 409 -1107
rect 65 -1129 66 -1109
rect 156 -1110 157 -1100
rect 163 -1110 164 -1100
rect 191 -1110 192 -1100
rect 226 -1129 227 -1109
rect 240 -1110 241 -1100
rect 247 -1129 248 -1109
rect 268 -1110 269 -1100
rect 275 -1110 276 -1100
rect 275 -1129 276 -1109
rect 275 -1110 276 -1100
rect 275 -1129 276 -1109
rect 320 -1110 321 -1100
rect 373 -1129 374 -1109
rect 394 -1110 395 -1100
rect 422 -1129 423 -1109
rect 72 -1112 73 -1100
rect 79 -1112 80 -1100
rect 82 -1129 83 -1111
rect 86 -1129 87 -1111
rect 121 -1129 122 -1111
rect 135 -1112 136 -1100
rect 142 -1129 143 -1111
rect 149 -1112 150 -1100
rect 159 -1129 160 -1111
rect 163 -1129 164 -1111
rect 170 -1112 171 -1100
rect 184 -1129 185 -1111
rect 191 -1129 192 -1111
rect 208 -1129 209 -1111
rect 233 -1129 234 -1111
rect 376 -1112 377 -1100
rect 401 -1112 402 -1100
rect 429 -1129 430 -1111
rect 44 -1129 45 -1113
rect 79 -1129 80 -1113
rect 107 -1114 108 -1100
rect 135 -1129 136 -1113
rect 170 -1129 171 -1113
rect 212 -1114 213 -1100
rect 268 -1129 269 -1113
rect 282 -1114 283 -1100
rect 289 -1129 290 -1113
rect 320 -1129 321 -1113
rect 324 -1114 325 -1100
rect 380 -1129 381 -1113
rect 75 -1129 76 -1115
rect 107 -1129 108 -1115
rect 131 -1129 132 -1115
rect 149 -1129 150 -1115
rect 198 -1116 199 -1100
rect 212 -1129 213 -1115
rect 278 -1129 279 -1115
rect 394 -1129 395 -1115
rect 205 -1118 206 -1100
rect 240 -1129 241 -1117
rect 282 -1129 283 -1117
rect 310 -1118 311 -1100
rect 331 -1118 332 -1100
rect 415 -1129 416 -1117
rect 194 -1129 195 -1119
rect 310 -1129 311 -1119
rect 338 -1129 339 -1119
rect 369 -1129 370 -1119
rect 205 -1129 206 -1121
rect 387 -1129 388 -1121
rect 261 -1124 262 -1100
rect 331 -1129 332 -1123
rect 180 -1126 181 -1100
rect 261 -1129 262 -1125
rect 296 -1126 297 -1100
rect 401 -1129 402 -1125
rect 264 -1129 265 -1127
rect 296 -1129 297 -1127
rect 30 -1139 31 -1137
rect 96 -1139 97 -1137
rect 107 -1139 108 -1137
rect 128 -1139 129 -1137
rect 149 -1139 150 -1137
rect 198 -1139 199 -1137
rect 205 -1139 206 -1137
rect 240 -1139 241 -1137
rect 250 -1172 251 -1138
rect 268 -1139 269 -1137
rect 275 -1139 276 -1137
rect 380 -1139 381 -1137
rect 397 -1172 398 -1138
rect 436 -1139 437 -1137
rect 478 -1139 479 -1137
rect 485 -1139 486 -1137
rect 37 -1141 38 -1137
rect 170 -1141 171 -1137
rect 177 -1141 178 -1137
rect 177 -1172 178 -1140
rect 177 -1141 178 -1137
rect 177 -1172 178 -1140
rect 184 -1141 185 -1137
rect 198 -1172 199 -1140
rect 229 -1141 230 -1137
rect 275 -1172 276 -1140
rect 296 -1141 297 -1137
rect 324 -1172 325 -1140
rect 327 -1141 328 -1137
rect 401 -1141 402 -1137
rect 44 -1143 45 -1137
rect 54 -1172 55 -1142
rect 58 -1143 59 -1137
rect 72 -1172 73 -1142
rect 75 -1143 76 -1137
rect 82 -1172 83 -1142
rect 86 -1172 87 -1142
rect 243 -1172 244 -1142
rect 254 -1143 255 -1137
rect 443 -1143 444 -1137
rect 65 -1145 66 -1137
rect 159 -1145 160 -1137
rect 163 -1145 164 -1137
rect 173 -1172 174 -1144
rect 184 -1172 185 -1144
rect 205 -1172 206 -1144
rect 261 -1145 262 -1137
rect 282 -1145 283 -1137
rect 299 -1172 300 -1144
rect 415 -1145 416 -1137
rect 79 -1147 80 -1137
rect 100 -1147 101 -1137
rect 107 -1172 108 -1146
rect 121 -1147 122 -1137
rect 128 -1172 129 -1146
rect 303 -1147 304 -1137
rect 306 -1147 307 -1137
rect 429 -1147 430 -1137
rect 89 -1149 90 -1137
rect 114 -1172 115 -1148
rect 117 -1149 118 -1137
rect 166 -1172 167 -1148
rect 201 -1149 202 -1137
rect 282 -1172 283 -1148
rect 306 -1172 307 -1148
rect 359 -1172 360 -1148
rect 369 -1149 370 -1137
rect 408 -1149 409 -1137
rect 93 -1172 94 -1150
rect 208 -1151 209 -1137
rect 261 -1172 262 -1150
rect 373 -1151 374 -1137
rect 376 -1172 377 -1150
rect 422 -1151 423 -1137
rect 100 -1172 101 -1152
rect 124 -1172 125 -1152
rect 149 -1172 150 -1152
rect 191 -1153 192 -1137
rect 208 -1172 209 -1152
rect 394 -1153 395 -1137
rect 401 -1172 402 -1152
rect 408 -1172 409 -1152
rect 117 -1172 118 -1154
rect 226 -1155 227 -1137
rect 268 -1172 269 -1154
rect 289 -1155 290 -1137
rect 310 -1155 311 -1137
rect 380 -1172 381 -1154
rect 121 -1172 122 -1156
rect 135 -1157 136 -1137
rect 156 -1172 157 -1156
rect 170 -1172 171 -1156
rect 191 -1172 192 -1156
rect 219 -1157 220 -1137
rect 278 -1157 279 -1137
rect 310 -1172 311 -1156
rect 317 -1172 318 -1156
rect 331 -1157 332 -1137
rect 338 -1157 339 -1137
rect 366 -1172 367 -1156
rect 135 -1172 136 -1158
rect 145 -1172 146 -1158
rect 163 -1172 164 -1158
rect 289 -1172 290 -1158
rect 212 -1161 213 -1137
rect 226 -1172 227 -1160
rect 240 -1172 241 -1160
rect 338 -1172 339 -1160
rect 142 -1163 143 -1137
rect 212 -1172 213 -1162
rect 219 -1172 220 -1162
rect 233 -1163 234 -1137
rect 264 -1163 265 -1137
rect 331 -1172 332 -1162
rect 233 -1172 234 -1164
rect 247 -1165 248 -1137
rect 264 -1172 265 -1164
rect 387 -1165 388 -1137
rect 352 -1167 353 -1137
rect 387 -1172 388 -1166
rect 345 -1169 346 -1137
rect 352 -1172 353 -1168
rect 254 -1172 255 -1170
rect 345 -1172 346 -1170
rect 61 -1182 62 -1180
rect 72 -1182 73 -1180
rect 79 -1203 80 -1181
rect 135 -1182 136 -1180
rect 163 -1203 164 -1181
rect 184 -1182 185 -1180
rect 198 -1182 199 -1180
rect 205 -1182 206 -1180
rect 208 -1182 209 -1180
rect 212 -1182 213 -1180
rect 240 -1182 241 -1180
rect 282 -1182 283 -1180
rect 292 -1203 293 -1181
rect 401 -1182 402 -1180
rect 72 -1203 73 -1183
rect 114 -1184 115 -1180
rect 121 -1184 122 -1180
rect 149 -1184 150 -1180
rect 177 -1184 178 -1180
rect 208 -1203 209 -1183
rect 212 -1203 213 -1183
rect 240 -1203 241 -1183
rect 247 -1184 248 -1180
rect 268 -1184 269 -1180
rect 303 -1184 304 -1180
rect 380 -1184 381 -1180
rect 86 -1186 87 -1180
rect 170 -1186 171 -1180
rect 173 -1203 174 -1185
rect 247 -1203 248 -1185
rect 250 -1186 251 -1180
rect 373 -1203 374 -1185
rect 376 -1186 377 -1180
rect 394 -1203 395 -1185
rect 65 -1203 66 -1187
rect 170 -1203 171 -1187
rect 184 -1203 185 -1187
rect 226 -1188 227 -1180
rect 254 -1203 255 -1187
rect 345 -1188 346 -1180
rect 359 -1188 360 -1180
rect 359 -1203 360 -1187
rect 359 -1188 360 -1180
rect 359 -1203 360 -1187
rect 366 -1188 367 -1180
rect 380 -1203 381 -1187
rect 93 -1203 94 -1189
rect 124 -1190 125 -1180
rect 128 -1190 129 -1180
rect 198 -1203 199 -1189
rect 201 -1190 202 -1180
rect 268 -1203 269 -1189
rect 324 -1190 325 -1180
rect 327 -1198 328 -1189
rect 331 -1190 332 -1180
rect 331 -1203 332 -1189
rect 331 -1190 332 -1180
rect 331 -1203 332 -1189
rect 366 -1203 367 -1189
rect 387 -1190 388 -1180
rect 107 -1192 108 -1180
rect 131 -1203 132 -1191
rect 194 -1203 195 -1191
rect 282 -1203 283 -1191
rect 324 -1203 325 -1191
rect 338 -1192 339 -1180
rect 383 -1203 384 -1191
rect 387 -1203 388 -1191
rect 100 -1194 101 -1180
rect 107 -1203 108 -1193
rect 114 -1203 115 -1193
rect 156 -1194 157 -1180
rect 233 -1194 234 -1180
rect 345 -1203 346 -1193
rect 100 -1203 101 -1195
rect 261 -1196 262 -1180
rect 338 -1203 339 -1195
rect 352 -1196 353 -1180
rect 121 -1203 122 -1197
rect 219 -1198 220 -1180
rect 233 -1203 234 -1197
rect 296 -1198 297 -1180
rect 352 -1203 353 -1197
rect 142 -1203 143 -1199
rect 156 -1203 157 -1199
rect 191 -1200 192 -1180
rect 219 -1203 220 -1199
rect 257 -1200 258 -1180
rect 275 -1200 276 -1180
rect 296 -1203 297 -1199
rect 310 -1200 311 -1180
rect 138 -1203 139 -1201
rect 191 -1203 192 -1201
rect 275 -1203 276 -1201
rect 289 -1202 290 -1180
rect 310 -1203 311 -1201
rect 317 -1202 318 -1180
rect 65 -1213 66 -1211
rect 191 -1213 192 -1211
rect 194 -1232 195 -1212
rect 247 -1213 248 -1211
rect 261 -1213 262 -1211
rect 289 -1232 290 -1212
rect 292 -1213 293 -1211
rect 352 -1213 353 -1211
rect 380 -1232 381 -1212
rect 387 -1213 388 -1211
rect 72 -1215 73 -1211
rect 89 -1215 90 -1211
rect 93 -1215 94 -1211
rect 93 -1232 94 -1214
rect 93 -1215 94 -1211
rect 93 -1232 94 -1214
rect 114 -1215 115 -1211
rect 156 -1232 157 -1214
rect 163 -1215 164 -1211
rect 163 -1232 164 -1214
rect 163 -1215 164 -1211
rect 163 -1232 164 -1214
rect 170 -1232 171 -1214
rect 247 -1232 248 -1214
rect 261 -1232 262 -1214
rect 373 -1215 374 -1211
rect 383 -1215 384 -1211
rect 394 -1215 395 -1211
rect 79 -1217 80 -1211
rect 138 -1217 139 -1211
rect 149 -1217 150 -1211
rect 219 -1217 220 -1211
rect 240 -1217 241 -1211
rect 359 -1217 360 -1211
rect 107 -1219 108 -1211
rect 114 -1232 115 -1218
rect 121 -1219 122 -1211
rect 243 -1219 244 -1211
rect 264 -1219 265 -1211
rect 345 -1219 346 -1211
rect 352 -1232 353 -1218
rect 366 -1219 367 -1211
rect 121 -1232 122 -1220
rect 180 -1221 181 -1211
rect 184 -1232 185 -1220
rect 226 -1232 227 -1220
rect 275 -1221 276 -1211
rect 317 -1221 318 -1211
rect 324 -1232 325 -1220
rect 331 -1221 332 -1211
rect 128 -1223 129 -1211
rect 159 -1223 160 -1211
rect 177 -1223 178 -1211
rect 254 -1223 255 -1211
rect 268 -1223 269 -1211
rect 317 -1232 318 -1222
rect 331 -1232 332 -1222
rect 338 -1223 339 -1211
rect 100 -1225 101 -1211
rect 128 -1232 129 -1224
rect 135 -1232 136 -1224
rect 187 -1225 188 -1211
rect 205 -1232 206 -1224
rect 212 -1225 213 -1211
rect 233 -1225 234 -1211
rect 268 -1232 269 -1224
rect 303 -1225 304 -1211
rect 310 -1225 311 -1211
rect 142 -1227 143 -1211
rect 180 -1232 181 -1226
rect 198 -1227 199 -1211
rect 233 -1232 234 -1226
rect 240 -1232 241 -1226
rect 254 -1232 255 -1226
rect 282 -1227 283 -1211
rect 310 -1232 311 -1226
rect 142 -1232 143 -1228
rect 152 -1232 153 -1228
rect 212 -1232 213 -1228
rect 229 -1229 230 -1211
rect 282 -1232 283 -1228
rect 296 -1229 297 -1211
rect 275 -1232 276 -1230
rect 296 -1232 297 -1230
rect 82 -1253 83 -1241
rect 86 -1253 87 -1241
rect 93 -1242 94 -1240
rect 100 -1242 101 -1240
rect 107 -1253 108 -1241
rect 117 -1253 118 -1241
rect 128 -1242 129 -1240
rect 152 -1242 153 -1240
rect 156 -1242 157 -1240
rect 201 -1242 202 -1240
rect 212 -1242 213 -1240
rect 219 -1242 220 -1240
rect 233 -1242 234 -1240
rect 261 -1242 262 -1240
rect 275 -1242 276 -1240
rect 296 -1253 297 -1241
rect 299 -1242 300 -1240
rect 310 -1242 311 -1240
rect 317 -1242 318 -1240
rect 320 -1253 321 -1241
rect 348 -1242 349 -1240
rect 352 -1242 353 -1240
rect 380 -1242 381 -1240
rect 380 -1253 381 -1241
rect 380 -1242 381 -1240
rect 380 -1253 381 -1241
rect 100 -1253 101 -1243
rect 121 -1253 122 -1243
rect 128 -1253 129 -1243
rect 142 -1244 143 -1240
rect 156 -1253 157 -1243
rect 226 -1244 227 -1240
rect 240 -1244 241 -1240
rect 261 -1253 262 -1243
rect 282 -1244 283 -1240
rect 303 -1253 304 -1243
rect 306 -1244 307 -1240
rect 324 -1244 325 -1240
rect 110 -1246 111 -1240
rect 114 -1246 115 -1240
rect 135 -1246 136 -1240
rect 173 -1253 174 -1245
rect 177 -1253 178 -1245
rect 191 -1246 192 -1240
rect 198 -1253 199 -1245
rect 219 -1253 220 -1245
rect 226 -1253 227 -1245
rect 233 -1253 234 -1245
rect 254 -1253 255 -1245
rect 278 -1253 279 -1245
rect 285 -1253 286 -1245
rect 289 -1246 290 -1240
rect 324 -1253 325 -1245
rect 331 -1246 332 -1240
rect 135 -1253 136 -1247
rect 149 -1253 150 -1247
rect 163 -1248 164 -1240
rect 187 -1248 188 -1240
rect 191 -1253 192 -1247
rect 205 -1248 206 -1240
rect 268 -1253 269 -1247
rect 289 -1253 290 -1247
rect 180 -1250 181 -1240
rect 247 -1250 248 -1240
rect 205 -1253 206 -1251
rect 215 -1253 216 -1251
rect 240 -1253 241 -1251
rect 247 -1253 248 -1251
rect 5 -1263 6 -1261
rect 5 -1268 6 -1262
rect 5 -1263 6 -1261
rect 5 -1268 6 -1262
rect 75 -1263 76 -1261
rect 79 -1263 80 -1261
rect 86 -1263 87 -1261
rect 86 -1268 87 -1262
rect 86 -1263 87 -1261
rect 86 -1268 87 -1262
rect 100 -1263 101 -1261
rect 128 -1263 129 -1261
rect 135 -1263 136 -1261
rect 166 -1263 167 -1261
rect 170 -1268 171 -1262
rect 173 -1263 174 -1261
rect 184 -1263 185 -1261
rect 184 -1268 185 -1262
rect 184 -1263 185 -1261
rect 184 -1268 185 -1262
rect 205 -1263 206 -1261
rect 226 -1268 227 -1262
rect 233 -1263 234 -1261
rect 233 -1268 234 -1262
rect 233 -1263 234 -1261
rect 233 -1268 234 -1262
rect 240 -1263 241 -1261
rect 240 -1268 241 -1262
rect 240 -1263 241 -1261
rect 240 -1268 241 -1262
rect 254 -1263 255 -1261
rect 271 -1268 272 -1262
rect 275 -1263 276 -1261
rect 296 -1263 297 -1261
rect 303 -1263 304 -1261
rect 303 -1268 304 -1262
rect 303 -1263 304 -1261
rect 303 -1268 304 -1262
rect 320 -1263 321 -1261
rect 324 -1263 325 -1261
rect 380 -1263 381 -1261
rect 387 -1268 388 -1262
rect 107 -1265 108 -1261
rect 107 -1268 108 -1264
rect 107 -1265 108 -1261
rect 107 -1268 108 -1264
rect 114 -1265 115 -1261
rect 121 -1265 122 -1261
rect 135 -1268 136 -1264
rect 145 -1265 146 -1261
rect 149 -1265 150 -1261
rect 149 -1268 150 -1264
rect 149 -1265 150 -1261
rect 149 -1268 150 -1264
rect 163 -1265 164 -1261
rect 177 -1265 178 -1261
rect 191 -1265 192 -1261
rect 205 -1268 206 -1264
rect 215 -1268 216 -1264
rect 219 -1265 220 -1261
rect 261 -1265 262 -1261
rect 278 -1265 279 -1261
rect 117 -1268 118 -1266
rect 121 -1268 122 -1266
rect 268 -1267 269 -1261
rect 275 -1268 276 -1266
rect 86 -1278 87 -1276
rect 96 -1278 97 -1276
rect 107 -1278 108 -1276
rect 117 -1278 118 -1276
rect 121 -1278 122 -1276
rect 128 -1278 129 -1276
rect 135 -1278 136 -1276
rect 145 -1278 146 -1276
rect 149 -1278 150 -1276
rect 159 -1278 160 -1276
rect 219 -1278 220 -1276
rect 226 -1278 227 -1276
rect 275 -1278 276 -1276
rect 282 -1278 283 -1276
rect 299 -1278 300 -1276
rect 303 -1278 304 -1276
rect 383 -1278 384 -1276
rect 387 -1278 388 -1276
rect 156 -1280 157 -1276
rect 166 -1280 167 -1276
<< labels >>
rlabel pdiffusion 3 -6 3 -6 0 cellNo=21
rlabel pdiffusion 10 -6 10 -6 0 cellNo=441
rlabel pdiffusion 17 -6 17 -6 0 cellNo=25
rlabel pdiffusion 24 -6 24 -6 0 cellNo=99
rlabel pdiffusion 31 -6 31 -6 0 cellNo=114
rlabel pdiffusion 38 -6 38 -6 0 cellNo=325
rlabel pdiffusion 45 -6 45 -6 0 cellNo=235
rlabel pdiffusion 52 -6 52 -6 0 cellNo=411
rlabel pdiffusion 59 -6 59 -6 0 cellNo=717
rlabel pdiffusion 136 -6 136 -6 0 feedthrough
rlabel pdiffusion 143 -6 143 -6 0 cellNo=490
rlabel pdiffusion 150 -6 150 -6 0 cellNo=111
rlabel pdiffusion 157 -6 157 -6 0 cellNo=280
rlabel pdiffusion 185 -6 185 -6 0 cellNo=383
rlabel pdiffusion 192 -6 192 -6 0 cellNo=137
rlabel pdiffusion 213 -6 213 -6 0 feedthrough
rlabel pdiffusion 220 -6 220 -6 0 cellNo=3
rlabel pdiffusion 255 -6 255 -6 0 cellNo=686
rlabel pdiffusion 3 -21 3 -21 0 cellNo=174
rlabel pdiffusion 10 -21 10 -21 0 cellNo=247
rlabel pdiffusion 17 -21 17 -21 0 cellNo=253
rlabel pdiffusion 24 -21 24 -21 0 cellNo=554
rlabel pdiffusion 31 -21 31 -21 0 cellNo=228
rlabel pdiffusion 38 -21 38 -21 0 cellNo=474
rlabel pdiffusion 45 -21 45 -21 0 cellNo=381
rlabel pdiffusion 52 -21 52 -21 0 cellNo=663
rlabel pdiffusion 143 -21 143 -21 0 cellNo=524
rlabel pdiffusion 150 -21 150 -21 0 feedthrough
rlabel pdiffusion 157 -21 157 -21 0 feedthrough
rlabel pdiffusion 164 -21 164 -21 0 cellNo=639
rlabel pdiffusion 171 -21 171 -21 0 cellNo=315
rlabel pdiffusion 178 -21 178 -21 0 cellNo=263
rlabel pdiffusion 185 -21 185 -21 0 feedthrough
rlabel pdiffusion 192 -21 192 -21 0 cellNo=170
rlabel pdiffusion 199 -21 199 -21 0 feedthrough
rlabel pdiffusion 206 -21 206 -21 0 cellNo=607
rlabel pdiffusion 213 -21 213 -21 0 feedthrough
rlabel pdiffusion 220 -21 220 -21 0 cellNo=589
rlabel pdiffusion 241 -21 241 -21 0 cellNo=193
rlabel pdiffusion 255 -21 255 -21 0 feedthrough
rlabel pdiffusion 262 -21 262 -21 0 cellNo=614
rlabel pdiffusion 269 -21 269 -21 0 cellNo=82
rlabel pdiffusion 311 -21 311 -21 0 cellNo=392
rlabel pdiffusion 3 -40 3 -40 0 cellNo=105
rlabel pdiffusion 10 -40 10 -40 0 cellNo=221
rlabel pdiffusion 17 -40 17 -40 0 cellNo=410
rlabel pdiffusion 24 -40 24 -40 0 cellNo=140
rlabel pdiffusion 31 -40 31 -40 0 cellNo=620
rlabel pdiffusion 38 -40 38 -40 0 cellNo=384
rlabel pdiffusion 45 -40 45 -40 0 cellNo=604
rlabel pdiffusion 52 -40 52 -40 0 cellNo=198
rlabel pdiffusion 101 -40 101 -40 0 cellNo=168
rlabel pdiffusion 143 -40 143 -40 0 cellNo=251
rlabel pdiffusion 150 -40 150 -40 0 feedthrough
rlabel pdiffusion 164 -40 164 -40 0 feedthrough
rlabel pdiffusion 171 -40 171 -40 0 cellNo=92
rlabel pdiffusion 178 -40 178 -40 0 cellNo=573
rlabel pdiffusion 185 -40 185 -40 0 cellNo=159
rlabel pdiffusion 192 -40 192 -40 0 feedthrough
rlabel pdiffusion 199 -40 199 -40 0 cellNo=495
rlabel pdiffusion 206 -40 206 -40 0 cellNo=510
rlabel pdiffusion 213 -40 213 -40 0 feedthrough
rlabel pdiffusion 220 -40 220 -40 0 feedthrough
rlabel pdiffusion 227 -40 227 -40 0 cellNo=120
rlabel pdiffusion 234 -40 234 -40 0 cellNo=59
rlabel pdiffusion 241 -40 241 -40 0 feedthrough
rlabel pdiffusion 248 -40 248 -40 0 feedthrough
rlabel pdiffusion 255 -40 255 -40 0 feedthrough
rlabel pdiffusion 262 -40 262 -40 0 feedthrough
rlabel pdiffusion 269 -40 269 -40 0 cellNo=172
rlabel pdiffusion 311 -40 311 -40 0 feedthrough
rlabel pdiffusion 339 -40 339 -40 0 cellNo=142
rlabel pdiffusion 346 -40 346 -40 0 feedthrough
rlabel pdiffusion 360 -40 360 -40 0 cellNo=426
rlabel pdiffusion 3 -63 3 -63 0 cellNo=88
rlabel pdiffusion 10 -63 10 -63 0 cellNo=100
rlabel pdiffusion 17 -63 17 -63 0 cellNo=310
rlabel pdiffusion 24 -63 24 -63 0 cellNo=336
rlabel pdiffusion 31 -63 31 -63 0 cellNo=339
rlabel pdiffusion 38 -63 38 -63 0 cellNo=591
rlabel pdiffusion 52 -63 52 -63 0 cellNo=64
rlabel pdiffusion 73 -63 73 -63 0 feedthrough
rlabel pdiffusion 94 -63 94 -63 0 cellNo=379
rlabel pdiffusion 101 -63 101 -63 0 feedthrough
rlabel pdiffusion 136 -63 136 -63 0 cellNo=244
rlabel pdiffusion 143 -63 143 -63 0 feedthrough
rlabel pdiffusion 150 -63 150 -63 0 cellNo=701
rlabel pdiffusion 157 -63 157 -63 0 cellNo=74
rlabel pdiffusion 164 -63 164 -63 0 feedthrough
rlabel pdiffusion 171 -63 171 -63 0 feedthrough
rlabel pdiffusion 178 -63 178 -63 0 cellNo=240
rlabel pdiffusion 185 -63 185 -63 0 cellNo=102
rlabel pdiffusion 192 -63 192 -63 0 cellNo=303
rlabel pdiffusion 199 -63 199 -63 0 cellNo=432
rlabel pdiffusion 206 -63 206 -63 0 feedthrough
rlabel pdiffusion 213 -63 213 -63 0 feedthrough
rlabel pdiffusion 220 -63 220 -63 0 feedthrough
rlabel pdiffusion 227 -63 227 -63 0 cellNo=334
rlabel pdiffusion 234 -63 234 -63 0 feedthrough
rlabel pdiffusion 241 -63 241 -63 0 cellNo=702
rlabel pdiffusion 248 -63 248 -63 0 feedthrough
rlabel pdiffusion 255 -63 255 -63 0 feedthrough
rlabel pdiffusion 262 -63 262 -63 0 feedthrough
rlabel pdiffusion 269 -63 269 -63 0 feedthrough
rlabel pdiffusion 276 -63 276 -63 0 cellNo=413
rlabel pdiffusion 283 -63 283 -63 0 cellNo=534
rlabel pdiffusion 290 -63 290 -63 0 feedthrough
rlabel pdiffusion 297 -63 297 -63 0 feedthrough
rlabel pdiffusion 311 -63 311 -63 0 feedthrough
rlabel pdiffusion 318 -63 318 -63 0 cellNo=128
rlabel pdiffusion 339 -63 339 -63 0 feedthrough
rlabel pdiffusion 346 -63 346 -63 0 cellNo=598
rlabel pdiffusion 353 -63 353 -63 0 feedthrough
rlabel pdiffusion 367 -63 367 -63 0 feedthrough
rlabel pdiffusion 3 -94 3 -94 0 cellNo=130
rlabel pdiffusion 10 -94 10 -94 0 cellNo=355
rlabel pdiffusion 17 -94 17 -94 0 cellNo=291
rlabel pdiffusion 24 -94 24 -94 0 cellNo=96
rlabel pdiffusion 31 -94 31 -94 0 cellNo=511
rlabel pdiffusion 52 -94 52 -94 0 cellNo=681
rlabel pdiffusion 59 -94 59 -94 0 feedthrough
rlabel pdiffusion 66 -94 66 -94 0 feedthrough
rlabel pdiffusion 73 -94 73 -94 0 feedthrough
rlabel pdiffusion 80 -94 80 -94 0 feedthrough
rlabel pdiffusion 87 -94 87 -94 0 cellNo=242
rlabel pdiffusion 94 -94 94 -94 0 feedthrough
rlabel pdiffusion 101 -94 101 -94 0 cellNo=577
rlabel pdiffusion 108 -94 108 -94 0 feedthrough
rlabel pdiffusion 115 -94 115 -94 0 feedthrough
rlabel pdiffusion 122 -94 122 -94 0 feedthrough
rlabel pdiffusion 129 -94 129 -94 0 feedthrough
rlabel pdiffusion 136 -94 136 -94 0 cellNo=34
rlabel pdiffusion 143 -94 143 -94 0 cellNo=110
rlabel pdiffusion 150 -94 150 -94 0 feedthrough
rlabel pdiffusion 157 -94 157 -94 0 feedthrough
rlabel pdiffusion 164 -94 164 -94 0 feedthrough
rlabel pdiffusion 171 -94 171 -94 0 cellNo=287
rlabel pdiffusion 178 -94 178 -94 0 cellNo=214
rlabel pdiffusion 185 -94 185 -94 0 cellNo=52
rlabel pdiffusion 192 -94 192 -94 0 cellNo=141
rlabel pdiffusion 199 -94 199 -94 0 cellNo=359
rlabel pdiffusion 206 -94 206 -94 0 cellNo=506
rlabel pdiffusion 213 -94 213 -94 0 feedthrough
rlabel pdiffusion 220 -94 220 -94 0 feedthrough
rlabel pdiffusion 227 -94 227 -94 0 cellNo=365
rlabel pdiffusion 234 -94 234 -94 0 cellNo=90
rlabel pdiffusion 241 -94 241 -94 0 cellNo=719
rlabel pdiffusion 248 -94 248 -94 0 cellNo=552
rlabel pdiffusion 255 -94 255 -94 0 cellNo=553
rlabel pdiffusion 262 -94 262 -94 0 feedthrough
rlabel pdiffusion 269 -94 269 -94 0 feedthrough
rlabel pdiffusion 276 -94 276 -94 0 feedthrough
rlabel pdiffusion 283 -94 283 -94 0 feedthrough
rlabel pdiffusion 290 -94 290 -94 0 feedthrough
rlabel pdiffusion 297 -94 297 -94 0 feedthrough
rlabel pdiffusion 304 -94 304 -94 0 feedthrough
rlabel pdiffusion 311 -94 311 -94 0 feedthrough
rlabel pdiffusion 318 -94 318 -94 0 feedthrough
rlabel pdiffusion 325 -94 325 -94 0 feedthrough
rlabel pdiffusion 332 -94 332 -94 0 feedthrough
rlabel pdiffusion 339 -94 339 -94 0 feedthrough
rlabel pdiffusion 346 -94 346 -94 0 feedthrough
rlabel pdiffusion 353 -94 353 -94 0 feedthrough
rlabel pdiffusion 367 -94 367 -94 0 feedthrough
rlabel pdiffusion 374 -94 374 -94 0 cellNo=375
rlabel pdiffusion 3 -137 3 -137 0 cellNo=180
rlabel pdiffusion 10 -137 10 -137 0 cellNo=276
rlabel pdiffusion 17 -137 17 -137 0 cellNo=331
rlabel pdiffusion 24 -137 24 -137 0 cellNo=496
rlabel pdiffusion 87 -137 87 -137 0 feedthrough
rlabel pdiffusion 94 -137 94 -137 0 feedthrough
rlabel pdiffusion 101 -137 101 -137 0 feedthrough
rlabel pdiffusion 108 -137 108 -137 0 feedthrough
rlabel pdiffusion 115 -137 115 -137 0 cellNo=63
rlabel pdiffusion 122 -137 122 -137 0 cellNo=61
rlabel pdiffusion 129 -137 129 -137 0 feedthrough
rlabel pdiffusion 136 -137 136 -137 0 feedthrough
rlabel pdiffusion 143 -137 143 -137 0 cellNo=65
rlabel pdiffusion 150 -137 150 -137 0 feedthrough
rlabel pdiffusion 157 -137 157 -137 0 cellNo=245
rlabel pdiffusion 164 -137 164 -137 0 feedthrough
rlabel pdiffusion 171 -137 171 -137 0 cellNo=185
rlabel pdiffusion 178 -137 178 -137 0 cellNo=80
rlabel pdiffusion 185 -137 185 -137 0 feedthrough
rlabel pdiffusion 192 -137 192 -137 0 cellNo=94
rlabel pdiffusion 199 -137 199 -137 0 feedthrough
rlabel pdiffusion 206 -137 206 -137 0 cellNo=9
rlabel pdiffusion 213 -137 213 -137 0 feedthrough
rlabel pdiffusion 220 -137 220 -137 0 feedthrough
rlabel pdiffusion 227 -137 227 -137 0 cellNo=138
rlabel pdiffusion 234 -137 234 -137 0 cellNo=684
rlabel pdiffusion 241 -137 241 -137 0 feedthrough
rlabel pdiffusion 248 -137 248 -137 0 cellNo=640
rlabel pdiffusion 255 -137 255 -137 0 feedthrough
rlabel pdiffusion 262 -137 262 -137 0 cellNo=555
rlabel pdiffusion 269 -137 269 -137 0 cellNo=700
rlabel pdiffusion 276 -137 276 -137 0 feedthrough
rlabel pdiffusion 283 -137 283 -137 0 cellNo=660
rlabel pdiffusion 290 -137 290 -137 0 cellNo=516
rlabel pdiffusion 297 -137 297 -137 0 feedthrough
rlabel pdiffusion 304 -137 304 -137 0 feedthrough
rlabel pdiffusion 311 -137 311 -137 0 cellNo=380
rlabel pdiffusion 318 -137 318 -137 0 feedthrough
rlabel pdiffusion 325 -137 325 -137 0 feedthrough
rlabel pdiffusion 332 -137 332 -137 0 feedthrough
rlabel pdiffusion 339 -137 339 -137 0 cellNo=621
rlabel pdiffusion 346 -137 346 -137 0 feedthrough
rlabel pdiffusion 353 -137 353 -137 0 cellNo=14
rlabel pdiffusion 367 -137 367 -137 0 feedthrough
rlabel pdiffusion 381 -137 381 -137 0 feedthrough
rlabel pdiffusion 395 -137 395 -137 0 feedthrough
rlabel pdiffusion 402 -137 402 -137 0 feedthrough
rlabel pdiffusion 3 -172 3 -172 0 cellNo=177
rlabel pdiffusion 10 -172 10 -172 0 cellNo=237
rlabel pdiffusion 17 -172 17 -172 0 cellNo=629
rlabel pdiffusion 66 -172 66 -172 0 feedthrough
rlabel pdiffusion 73 -172 73 -172 0 feedthrough
rlabel pdiffusion 80 -172 80 -172 0 cellNo=543
rlabel pdiffusion 87 -172 87 -172 0 feedthrough
rlabel pdiffusion 94 -172 94 -172 0 feedthrough
rlabel pdiffusion 101 -172 101 -172 0 feedthrough
rlabel pdiffusion 108 -172 108 -172 0 feedthrough
rlabel pdiffusion 115 -172 115 -172 0 cellNo=343
rlabel pdiffusion 122 -172 122 -172 0 feedthrough
rlabel pdiffusion 129 -172 129 -172 0 cellNo=377
rlabel pdiffusion 136 -172 136 -172 0 cellNo=16
rlabel pdiffusion 143 -172 143 -172 0 cellNo=548
rlabel pdiffusion 150 -172 150 -172 0 cellNo=153
rlabel pdiffusion 157 -172 157 -172 0 feedthrough
rlabel pdiffusion 164 -172 164 -172 0 cellNo=67
rlabel pdiffusion 171 -172 171 -172 0 feedthrough
rlabel pdiffusion 178 -172 178 -172 0 cellNo=187
rlabel pdiffusion 185 -172 185 -172 0 feedthrough
rlabel pdiffusion 192 -172 192 -172 0 feedthrough
rlabel pdiffusion 199 -172 199 -172 0 cellNo=590
rlabel pdiffusion 206 -172 206 -172 0 cellNo=51
rlabel pdiffusion 213 -172 213 -172 0 feedthrough
rlabel pdiffusion 220 -172 220 -172 0 cellNo=505
rlabel pdiffusion 227 -172 227 -172 0 cellNo=605
rlabel pdiffusion 234 -172 234 -172 0 feedthrough
rlabel pdiffusion 241 -172 241 -172 0 cellNo=347
rlabel pdiffusion 248 -172 248 -172 0 cellNo=157
rlabel pdiffusion 255 -172 255 -172 0 feedthrough
rlabel pdiffusion 262 -172 262 -172 0 feedthrough
rlabel pdiffusion 269 -172 269 -172 0 feedthrough
rlabel pdiffusion 276 -172 276 -172 0 feedthrough
rlabel pdiffusion 283 -172 283 -172 0 cellNo=583
rlabel pdiffusion 290 -172 290 -172 0 feedthrough
rlabel pdiffusion 297 -172 297 -172 0 feedthrough
rlabel pdiffusion 304 -172 304 -172 0 feedthrough
rlabel pdiffusion 311 -172 311 -172 0 cellNo=45
rlabel pdiffusion 318 -172 318 -172 0 cellNo=649
rlabel pdiffusion 325 -172 325 -172 0 feedthrough
rlabel pdiffusion 332 -172 332 -172 0 feedthrough
rlabel pdiffusion 339 -172 339 -172 0 cellNo=230
rlabel pdiffusion 346 -172 346 -172 0 feedthrough
rlabel pdiffusion 353 -172 353 -172 0 feedthrough
rlabel pdiffusion 360 -172 360 -172 0 feedthrough
rlabel pdiffusion 367 -172 367 -172 0 feedthrough
rlabel pdiffusion 374 -172 374 -172 0 cellNo=612
rlabel pdiffusion 381 -172 381 -172 0 feedthrough
rlabel pdiffusion 388 -172 388 -172 0 cellNo=77
rlabel pdiffusion 395 -172 395 -172 0 feedthrough
rlabel pdiffusion 402 -172 402 -172 0 feedthrough
rlabel pdiffusion 409 -172 409 -172 0 feedthrough
rlabel pdiffusion 416 -172 416 -172 0 feedthrough
rlabel pdiffusion 423 -172 423 -172 0 feedthrough
rlabel pdiffusion 430 -172 430 -172 0 cellNo=458
rlabel pdiffusion 437 -172 437 -172 0 cellNo=600
rlabel pdiffusion 3 -211 3 -211 0 cellNo=402
rlabel pdiffusion 10 -211 10 -211 0 cellNo=439
rlabel pdiffusion 24 -211 24 -211 0 feedthrough
rlabel pdiffusion 31 -211 31 -211 0 feedthrough
rlabel pdiffusion 38 -211 38 -211 0 feedthrough
rlabel pdiffusion 45 -211 45 -211 0 feedthrough
rlabel pdiffusion 52 -211 52 -211 0 feedthrough
rlabel pdiffusion 59 -211 59 -211 0 cellNo=261
rlabel pdiffusion 66 -211 66 -211 0 cellNo=340
rlabel pdiffusion 73 -211 73 -211 0 cellNo=113
rlabel pdiffusion 80 -211 80 -211 0 feedthrough
rlabel pdiffusion 87 -211 87 -211 0 cellNo=536
rlabel pdiffusion 94 -211 94 -211 0 cellNo=156
rlabel pdiffusion 101 -211 101 -211 0 feedthrough
rlabel pdiffusion 108 -211 108 -211 0 feedthrough
rlabel pdiffusion 115 -211 115 -211 0 feedthrough
rlabel pdiffusion 122 -211 122 -211 0 feedthrough
rlabel pdiffusion 129 -211 129 -211 0 feedthrough
rlabel pdiffusion 136 -211 136 -211 0 cellNo=390
rlabel pdiffusion 143 -211 143 -211 0 cellNo=547
rlabel pdiffusion 150 -211 150 -211 0 cellNo=386
rlabel pdiffusion 157 -211 157 -211 0 cellNo=231
rlabel pdiffusion 164 -211 164 -211 0 feedthrough
rlabel pdiffusion 171 -211 171 -211 0 feedthrough
rlabel pdiffusion 178 -211 178 -211 0 feedthrough
rlabel pdiffusion 185 -211 185 -211 0 feedthrough
rlabel pdiffusion 192 -211 192 -211 0 cellNo=165
rlabel pdiffusion 199 -211 199 -211 0 cellNo=714
rlabel pdiffusion 206 -211 206 -211 0 cellNo=529
rlabel pdiffusion 213 -211 213 -211 0 cellNo=476
rlabel pdiffusion 220 -211 220 -211 0 feedthrough
rlabel pdiffusion 227 -211 227 -211 0 feedthrough
rlabel pdiffusion 234 -211 234 -211 0 cellNo=415
rlabel pdiffusion 241 -211 241 -211 0 cellNo=6
rlabel pdiffusion 248 -211 248 -211 0 feedthrough
rlabel pdiffusion 255 -211 255 -211 0 feedthrough
rlabel pdiffusion 262 -211 262 -211 0 feedthrough
rlabel pdiffusion 269 -211 269 -211 0 cellNo=129
rlabel pdiffusion 276 -211 276 -211 0 feedthrough
rlabel pdiffusion 283 -211 283 -211 0 cellNo=403
rlabel pdiffusion 290 -211 290 -211 0 feedthrough
rlabel pdiffusion 297 -211 297 -211 0 cellNo=608
rlabel pdiffusion 304 -211 304 -211 0 feedthrough
rlabel pdiffusion 311 -211 311 -211 0 feedthrough
rlabel pdiffusion 318 -211 318 -211 0 feedthrough
rlabel pdiffusion 325 -211 325 -211 0 cellNo=148
rlabel pdiffusion 332 -211 332 -211 0 feedthrough
rlabel pdiffusion 339 -211 339 -211 0 cellNo=206
rlabel pdiffusion 346 -211 346 -211 0 feedthrough
rlabel pdiffusion 353 -211 353 -211 0 feedthrough
rlabel pdiffusion 360 -211 360 -211 0 feedthrough
rlabel pdiffusion 367 -211 367 -211 0 feedthrough
rlabel pdiffusion 374 -211 374 -211 0 cellNo=126
rlabel pdiffusion 381 -211 381 -211 0 feedthrough
rlabel pdiffusion 388 -211 388 -211 0 feedthrough
rlabel pdiffusion 395 -211 395 -211 0 feedthrough
rlabel pdiffusion 402 -211 402 -211 0 feedthrough
rlabel pdiffusion 409 -211 409 -211 0 cellNo=358
rlabel pdiffusion 416 -211 416 -211 0 feedthrough
rlabel pdiffusion 423 -211 423 -211 0 feedthrough
rlabel pdiffusion 430 -211 430 -211 0 feedthrough
rlabel pdiffusion 437 -211 437 -211 0 feedthrough
rlabel pdiffusion 444 -211 444 -211 0 feedthrough
rlabel pdiffusion 451 -211 451 -211 0 feedthrough
rlabel pdiffusion 458 -211 458 -211 0 feedthrough
rlabel pdiffusion 465 -211 465 -211 0 feedthrough
rlabel pdiffusion 542 -211 542 -211 0 cellNo=603
rlabel pdiffusion 3 -258 3 -258 0 cellNo=412
rlabel pdiffusion 38 -258 38 -258 0 feedthrough
rlabel pdiffusion 45 -258 45 -258 0 feedthrough
rlabel pdiffusion 52 -258 52 -258 0 feedthrough
rlabel pdiffusion 59 -258 59 -258 0 feedthrough
rlabel pdiffusion 66 -258 66 -258 0 feedthrough
rlabel pdiffusion 73 -258 73 -258 0 cellNo=585
rlabel pdiffusion 80 -258 80 -258 0 feedthrough
rlabel pdiffusion 87 -258 87 -258 0 feedthrough
rlabel pdiffusion 94 -258 94 -258 0 feedthrough
rlabel pdiffusion 101 -258 101 -258 0 feedthrough
rlabel pdiffusion 108 -258 108 -258 0 cellNo=8
rlabel pdiffusion 115 -258 115 -258 0 cellNo=32
rlabel pdiffusion 122 -258 122 -258 0 cellNo=219
rlabel pdiffusion 129 -258 129 -258 0 cellNo=83
rlabel pdiffusion 136 -258 136 -258 0 feedthrough
rlabel pdiffusion 143 -258 143 -258 0 cellNo=350
rlabel pdiffusion 150 -258 150 -258 0 cellNo=672
rlabel pdiffusion 157 -258 157 -258 0 feedthrough
rlabel pdiffusion 164 -258 164 -258 0 cellNo=519
rlabel pdiffusion 171 -258 171 -258 0 cellNo=696
rlabel pdiffusion 178 -258 178 -258 0 cellNo=538
rlabel pdiffusion 185 -258 185 -258 0 feedthrough
rlabel pdiffusion 192 -258 192 -258 0 feedthrough
rlabel pdiffusion 199 -258 199 -258 0 cellNo=293
rlabel pdiffusion 206 -258 206 -258 0 cellNo=189
rlabel pdiffusion 213 -258 213 -258 0 feedthrough
rlabel pdiffusion 220 -258 220 -258 0 feedthrough
rlabel pdiffusion 227 -258 227 -258 0 cellNo=447
rlabel pdiffusion 234 -258 234 -258 0 cellNo=107
rlabel pdiffusion 241 -258 241 -258 0 cellNo=387
rlabel pdiffusion 248 -258 248 -258 0 feedthrough
rlabel pdiffusion 255 -258 255 -258 0 feedthrough
rlabel pdiffusion 262 -258 262 -258 0 feedthrough
rlabel pdiffusion 269 -258 269 -258 0 feedthrough
rlabel pdiffusion 276 -258 276 -258 0 feedthrough
rlabel pdiffusion 283 -258 283 -258 0 cellNo=188
rlabel pdiffusion 290 -258 290 -258 0 feedthrough
rlabel pdiffusion 297 -258 297 -258 0 feedthrough
rlabel pdiffusion 304 -258 304 -258 0 cellNo=171
rlabel pdiffusion 311 -258 311 -258 0 feedthrough
rlabel pdiffusion 318 -258 318 -258 0 feedthrough
rlabel pdiffusion 325 -258 325 -258 0 cellNo=89
rlabel pdiffusion 332 -258 332 -258 0 cellNo=55
rlabel pdiffusion 339 -258 339 -258 0 cellNo=256
rlabel pdiffusion 346 -258 346 -258 0 cellNo=123
rlabel pdiffusion 353 -258 353 -258 0 cellNo=345
rlabel pdiffusion 360 -258 360 -258 0 feedthrough
rlabel pdiffusion 367 -258 367 -258 0 feedthrough
rlabel pdiffusion 374 -258 374 -258 0 feedthrough
rlabel pdiffusion 381 -258 381 -258 0 feedthrough
rlabel pdiffusion 388 -258 388 -258 0 feedthrough
rlabel pdiffusion 395 -258 395 -258 0 feedthrough
rlabel pdiffusion 402 -258 402 -258 0 feedthrough
rlabel pdiffusion 409 -258 409 -258 0 feedthrough
rlabel pdiffusion 416 -258 416 -258 0 feedthrough
rlabel pdiffusion 423 -258 423 -258 0 feedthrough
rlabel pdiffusion 430 -258 430 -258 0 feedthrough
rlabel pdiffusion 437 -258 437 -258 0 feedthrough
rlabel pdiffusion 444 -258 444 -258 0 feedthrough
rlabel pdiffusion 451 -258 451 -258 0 feedthrough
rlabel pdiffusion 458 -258 458 -258 0 feedthrough
rlabel pdiffusion 465 -258 465 -258 0 feedthrough
rlabel pdiffusion 472 -258 472 -258 0 feedthrough
rlabel pdiffusion 479 -258 479 -258 0 feedthrough
rlabel pdiffusion 486 -258 486 -258 0 feedthrough
rlabel pdiffusion 493 -258 493 -258 0 feedthrough
rlabel pdiffusion 500 -258 500 -258 0 feedthrough
rlabel pdiffusion 507 -258 507 -258 0 feedthrough
rlabel pdiffusion 514 -258 514 -258 0 feedthrough
rlabel pdiffusion 521 -258 521 -258 0 feedthrough
rlabel pdiffusion 528 -258 528 -258 0 cellNo=616
rlabel pdiffusion 535 -258 535 -258 0 cellNo=501
rlabel pdiffusion 542 -258 542 -258 0 feedthrough
rlabel pdiffusion 3 -305 3 -305 0 cellNo=720
rlabel pdiffusion 38 -305 38 -305 0 feedthrough
rlabel pdiffusion 45 -305 45 -305 0 cellNo=483
rlabel pdiffusion 52 -305 52 -305 0 feedthrough
rlabel pdiffusion 59 -305 59 -305 0 cellNo=190
rlabel pdiffusion 66 -305 66 -305 0 feedthrough
rlabel pdiffusion 73 -305 73 -305 0 feedthrough
rlabel pdiffusion 80 -305 80 -305 0 cellNo=560
rlabel pdiffusion 87 -305 87 -305 0 cellNo=207
rlabel pdiffusion 94 -305 94 -305 0 cellNo=368
rlabel pdiffusion 101 -305 101 -305 0 feedthrough
rlabel pdiffusion 108 -305 108 -305 0 feedthrough
rlabel pdiffusion 115 -305 115 -305 0 cellNo=31
rlabel pdiffusion 122 -305 122 -305 0 feedthrough
rlabel pdiffusion 129 -305 129 -305 0 cellNo=705
rlabel pdiffusion 136 -305 136 -305 0 feedthrough
rlabel pdiffusion 143 -305 143 -305 0 feedthrough
rlabel pdiffusion 150 -305 150 -305 0 feedthrough
rlabel pdiffusion 157 -305 157 -305 0 feedthrough
rlabel pdiffusion 164 -305 164 -305 0 feedthrough
rlabel pdiffusion 171 -305 171 -305 0 feedthrough
rlabel pdiffusion 178 -305 178 -305 0 feedthrough
rlabel pdiffusion 185 -305 185 -305 0 feedthrough
rlabel pdiffusion 192 -305 192 -305 0 cellNo=212
rlabel pdiffusion 199 -305 199 -305 0 feedthrough
rlabel pdiffusion 206 -305 206 -305 0 feedthrough
rlabel pdiffusion 213 -305 213 -305 0 feedthrough
rlabel pdiffusion 220 -305 220 -305 0 feedthrough
rlabel pdiffusion 227 -305 227 -305 0 feedthrough
rlabel pdiffusion 234 -305 234 -305 0 feedthrough
rlabel pdiffusion 241 -305 241 -305 0 feedthrough
rlabel pdiffusion 248 -305 248 -305 0 cellNo=194
rlabel pdiffusion 255 -305 255 -305 0 feedthrough
rlabel pdiffusion 262 -305 262 -305 0 feedthrough
rlabel pdiffusion 269 -305 269 -305 0 cellNo=39
rlabel pdiffusion 276 -305 276 -305 0 feedthrough
rlabel pdiffusion 283 -305 283 -305 0 cellNo=195
rlabel pdiffusion 290 -305 290 -305 0 feedthrough
rlabel pdiffusion 297 -305 297 -305 0 feedthrough
rlabel pdiffusion 304 -305 304 -305 0 cellNo=544
rlabel pdiffusion 311 -305 311 -305 0 feedthrough
rlabel pdiffusion 318 -305 318 -305 0 cellNo=103
rlabel pdiffusion 325 -305 325 -305 0 feedthrough
rlabel pdiffusion 332 -305 332 -305 0 cellNo=707
rlabel pdiffusion 339 -305 339 -305 0 cellNo=42
rlabel pdiffusion 346 -305 346 -305 0 cellNo=30
rlabel pdiffusion 353 -305 353 -305 0 feedthrough
rlabel pdiffusion 360 -305 360 -305 0 cellNo=277
rlabel pdiffusion 367 -305 367 -305 0 cellNo=321
rlabel pdiffusion 374 -305 374 -305 0 feedthrough
rlabel pdiffusion 381 -305 381 -305 0 cellNo=154
rlabel pdiffusion 388 -305 388 -305 0 feedthrough
rlabel pdiffusion 395 -305 395 -305 0 feedthrough
rlabel pdiffusion 402 -305 402 -305 0 feedthrough
rlabel pdiffusion 409 -305 409 -305 0 feedthrough
rlabel pdiffusion 416 -305 416 -305 0 feedthrough
rlabel pdiffusion 423 -305 423 -305 0 feedthrough
rlabel pdiffusion 430 -305 430 -305 0 feedthrough
rlabel pdiffusion 437 -305 437 -305 0 feedthrough
rlabel pdiffusion 444 -305 444 -305 0 feedthrough
rlabel pdiffusion 451 -305 451 -305 0 feedthrough
rlabel pdiffusion 458 -305 458 -305 0 feedthrough
rlabel pdiffusion 465 -305 465 -305 0 cellNo=374
rlabel pdiffusion 472 -305 472 -305 0 feedthrough
rlabel pdiffusion 479 -305 479 -305 0 feedthrough
rlabel pdiffusion 486 -305 486 -305 0 feedthrough
rlabel pdiffusion 493 -305 493 -305 0 feedthrough
rlabel pdiffusion 500 -305 500 -305 0 feedthrough
rlabel pdiffusion 507 -305 507 -305 0 feedthrough
rlabel pdiffusion 514 -305 514 -305 0 feedthrough
rlabel pdiffusion 521 -305 521 -305 0 feedthrough
rlabel pdiffusion 528 -305 528 -305 0 feedthrough
rlabel pdiffusion 535 -305 535 -305 0 feedthrough
rlabel pdiffusion 542 -305 542 -305 0 cellNo=155
rlabel pdiffusion 549 -305 549 -305 0 feedthrough
rlabel pdiffusion 556 -305 556 -305 0 cellNo=18
rlabel pdiffusion 563 -305 563 -305 0 cellNo=192
rlabel pdiffusion 570 -305 570 -305 0 cellNo=201
rlabel pdiffusion 577 -305 577 -305 0 feedthrough
rlabel pdiffusion 10 -366 10 -366 0 feedthrough
rlabel pdiffusion 17 -366 17 -366 0 feedthrough
rlabel pdiffusion 24 -366 24 -366 0 feedthrough
rlabel pdiffusion 31 -366 31 -366 0 feedthrough
rlabel pdiffusion 38 -366 38 -366 0 cellNo=191
rlabel pdiffusion 45 -366 45 -366 0 feedthrough
rlabel pdiffusion 52 -366 52 -366 0 feedthrough
rlabel pdiffusion 59 -366 59 -366 0 cellNo=124
rlabel pdiffusion 66 -366 66 -366 0 feedthrough
rlabel pdiffusion 73 -366 73 -366 0 feedthrough
rlabel pdiffusion 80 -366 80 -366 0 feedthrough
rlabel pdiffusion 87 -366 87 -366 0 feedthrough
rlabel pdiffusion 94 -366 94 -366 0 feedthrough
rlabel pdiffusion 101 -366 101 -366 0 cellNo=408
rlabel pdiffusion 108 -366 108 -366 0 cellNo=394
rlabel pdiffusion 115 -366 115 -366 0 feedthrough
rlabel pdiffusion 122 -366 122 -366 0 cellNo=76
rlabel pdiffusion 129 -366 129 -366 0 cellNo=33
rlabel pdiffusion 136 -366 136 -366 0 cellNo=307
rlabel pdiffusion 143 -366 143 -366 0 feedthrough
rlabel pdiffusion 150 -366 150 -366 0 cellNo=398
rlabel pdiffusion 157 -366 157 -366 0 cellNo=84
rlabel pdiffusion 164 -366 164 -366 0 feedthrough
rlabel pdiffusion 171 -366 171 -366 0 feedthrough
rlabel pdiffusion 178 -366 178 -366 0 cellNo=298
rlabel pdiffusion 185 -366 185 -366 0 feedthrough
rlabel pdiffusion 192 -366 192 -366 0 cellNo=427
rlabel pdiffusion 199 -366 199 -366 0 feedthrough
rlabel pdiffusion 206 -366 206 -366 0 cellNo=182
rlabel pdiffusion 213 -366 213 -366 0 feedthrough
rlabel pdiffusion 220 -366 220 -366 0 feedthrough
rlabel pdiffusion 227 -366 227 -366 0 feedthrough
rlabel pdiffusion 234 -366 234 -366 0 feedthrough
rlabel pdiffusion 241 -366 241 -366 0 cellNo=35
rlabel pdiffusion 248 -366 248 -366 0 feedthrough
rlabel pdiffusion 255 -366 255 -366 0 feedthrough
rlabel pdiffusion 262 -366 262 -366 0 feedthrough
rlabel pdiffusion 269 -366 269 -366 0 cellNo=306
rlabel pdiffusion 276 -366 276 -366 0 feedthrough
rlabel pdiffusion 283 -366 283 -366 0 cellNo=317
rlabel pdiffusion 290 -366 290 -366 0 cellNo=436
rlabel pdiffusion 297 -366 297 -366 0 cellNo=220
rlabel pdiffusion 304 -366 304 -366 0 feedthrough
rlabel pdiffusion 311 -366 311 -366 0 cellNo=19
rlabel pdiffusion 318 -366 318 -366 0 feedthrough
rlabel pdiffusion 325 -366 325 -366 0 cellNo=593
rlabel pdiffusion 332 -366 332 -366 0 cellNo=716
rlabel pdiffusion 339 -366 339 -366 0 cellNo=178
rlabel pdiffusion 346 -366 346 -366 0 cellNo=266
rlabel pdiffusion 353 -366 353 -366 0 cellNo=197
rlabel pdiffusion 360 -366 360 -366 0 feedthrough
rlabel pdiffusion 367 -366 367 -366 0 cellNo=297
rlabel pdiffusion 374 -366 374 -366 0 feedthrough
rlabel pdiffusion 381 -366 381 -366 0 cellNo=367
rlabel pdiffusion 388 -366 388 -366 0 feedthrough
rlabel pdiffusion 395 -366 395 -366 0 feedthrough
rlabel pdiffusion 402 -366 402 -366 0 feedthrough
rlabel pdiffusion 409 -366 409 -366 0 feedthrough
rlabel pdiffusion 416 -366 416 -366 0 feedthrough
rlabel pdiffusion 423 -366 423 -366 0 feedthrough
rlabel pdiffusion 430 -366 430 -366 0 feedthrough
rlabel pdiffusion 437 -366 437 -366 0 feedthrough
rlabel pdiffusion 444 -366 444 -366 0 feedthrough
rlabel pdiffusion 451 -366 451 -366 0 feedthrough
rlabel pdiffusion 458 -366 458 -366 0 feedthrough
rlabel pdiffusion 465 -366 465 -366 0 feedthrough
rlabel pdiffusion 472 -366 472 -366 0 feedthrough
rlabel pdiffusion 479 -366 479 -366 0 feedthrough
rlabel pdiffusion 486 -366 486 -366 0 feedthrough
rlabel pdiffusion 493 -366 493 -366 0 feedthrough
rlabel pdiffusion 500 -366 500 -366 0 feedthrough
rlabel pdiffusion 507 -366 507 -366 0 feedthrough
rlabel pdiffusion 514 -366 514 -366 0 feedthrough
rlabel pdiffusion 521 -366 521 -366 0 feedthrough
rlabel pdiffusion 528 -366 528 -366 0 feedthrough
rlabel pdiffusion 535 -366 535 -366 0 feedthrough
rlabel pdiffusion 542 -366 542 -366 0 feedthrough
rlabel pdiffusion 549 -366 549 -366 0 feedthrough
rlabel pdiffusion 556 -366 556 -366 0 cellNo=227
rlabel pdiffusion 563 -366 563 -366 0 feedthrough
rlabel pdiffusion 570 -366 570 -366 0 feedthrough
rlabel pdiffusion 577 -366 577 -366 0 feedthrough
rlabel pdiffusion 3 -421 3 -421 0 feedthrough
rlabel pdiffusion 10 -421 10 -421 0 cellNo=364
rlabel pdiffusion 17 -421 17 -421 0 cellNo=246
rlabel pdiffusion 24 -421 24 -421 0 feedthrough
rlabel pdiffusion 31 -421 31 -421 0 cellNo=44
rlabel pdiffusion 38 -421 38 -421 0 feedthrough
rlabel pdiffusion 45 -421 45 -421 0 feedthrough
rlabel pdiffusion 52 -421 52 -421 0 feedthrough
rlabel pdiffusion 59 -421 59 -421 0 feedthrough
rlabel pdiffusion 66 -421 66 -421 0 cellNo=622
rlabel pdiffusion 73 -421 73 -421 0 feedthrough
rlabel pdiffusion 80 -421 80 -421 0 feedthrough
rlabel pdiffusion 87 -421 87 -421 0 cellNo=273
rlabel pdiffusion 94 -421 94 -421 0 cellNo=648
rlabel pdiffusion 101 -421 101 -421 0 cellNo=449
rlabel pdiffusion 108 -421 108 -421 0 feedthrough
rlabel pdiffusion 115 -421 115 -421 0 feedthrough
rlabel pdiffusion 122 -421 122 -421 0 feedthrough
rlabel pdiffusion 129 -421 129 -421 0 cellNo=520
rlabel pdiffusion 136 -421 136 -421 0 cellNo=243
rlabel pdiffusion 143 -421 143 -421 0 feedthrough
rlabel pdiffusion 150 -421 150 -421 0 cellNo=709
rlabel pdiffusion 157 -421 157 -421 0 cellNo=41
rlabel pdiffusion 164 -421 164 -421 0 feedthrough
rlabel pdiffusion 171 -421 171 -421 0 feedthrough
rlabel pdiffusion 178 -421 178 -421 0 feedthrough
rlabel pdiffusion 185 -421 185 -421 0 feedthrough
rlabel pdiffusion 192 -421 192 -421 0 feedthrough
rlabel pdiffusion 199 -421 199 -421 0 cellNo=341
rlabel pdiffusion 206 -421 206 -421 0 cellNo=658
rlabel pdiffusion 213 -421 213 -421 0 feedthrough
rlabel pdiffusion 220 -421 220 -421 0 feedthrough
rlabel pdiffusion 227 -421 227 -421 0 feedthrough
rlabel pdiffusion 234 -421 234 -421 0 feedthrough
rlabel pdiffusion 241 -421 241 -421 0 cellNo=249
rlabel pdiffusion 248 -421 248 -421 0 cellNo=482
rlabel pdiffusion 255 -421 255 -421 0 cellNo=270
rlabel pdiffusion 262 -421 262 -421 0 feedthrough
rlabel pdiffusion 269 -421 269 -421 0 cellNo=104
rlabel pdiffusion 276 -421 276 -421 0 cellNo=360
rlabel pdiffusion 283 -421 283 -421 0 feedthrough
rlabel pdiffusion 290 -421 290 -421 0 cellNo=81
rlabel pdiffusion 297 -421 297 -421 0 feedthrough
rlabel pdiffusion 304 -421 304 -421 0 cellNo=499
rlabel pdiffusion 311 -421 311 -421 0 feedthrough
rlabel pdiffusion 318 -421 318 -421 0 cellNo=132
rlabel pdiffusion 325 -421 325 -421 0 cellNo=354
rlabel pdiffusion 332 -421 332 -421 0 feedthrough
rlabel pdiffusion 339 -421 339 -421 0 feedthrough
rlabel pdiffusion 346 -421 346 -421 0 cellNo=289
rlabel pdiffusion 353 -421 353 -421 0 feedthrough
rlabel pdiffusion 360 -421 360 -421 0 cellNo=464
rlabel pdiffusion 367 -421 367 -421 0 feedthrough
rlabel pdiffusion 374 -421 374 -421 0 feedthrough
rlabel pdiffusion 381 -421 381 -421 0 cellNo=642
rlabel pdiffusion 388 -421 388 -421 0 cellNo=631
rlabel pdiffusion 395 -421 395 -421 0 feedthrough
rlabel pdiffusion 402 -421 402 -421 0 feedthrough
rlabel pdiffusion 409 -421 409 -421 0 cellNo=15
rlabel pdiffusion 416 -421 416 -421 0 feedthrough
rlabel pdiffusion 423 -421 423 -421 0 feedthrough
rlabel pdiffusion 430 -421 430 -421 0 feedthrough
rlabel pdiffusion 437 -421 437 -421 0 feedthrough
rlabel pdiffusion 444 -421 444 -421 0 feedthrough
rlabel pdiffusion 451 -421 451 -421 0 feedthrough
rlabel pdiffusion 458 -421 458 -421 0 feedthrough
rlabel pdiffusion 465 -421 465 -421 0 feedthrough
rlabel pdiffusion 472 -421 472 -421 0 feedthrough
rlabel pdiffusion 479 -421 479 -421 0 feedthrough
rlabel pdiffusion 486 -421 486 -421 0 feedthrough
rlabel pdiffusion 493 -421 493 -421 0 feedthrough
rlabel pdiffusion 500 -421 500 -421 0 feedthrough
rlabel pdiffusion 507 -421 507 -421 0 feedthrough
rlabel pdiffusion 514 -421 514 -421 0 feedthrough
rlabel pdiffusion 521 -421 521 -421 0 cellNo=558
rlabel pdiffusion 528 -421 528 -421 0 feedthrough
rlabel pdiffusion 535 -421 535 -421 0 feedthrough
rlabel pdiffusion 542 -421 542 -421 0 feedthrough
rlabel pdiffusion 549 -421 549 -421 0 feedthrough
rlabel pdiffusion 556 -421 556 -421 0 feedthrough
rlabel pdiffusion 563 -421 563 -421 0 feedthrough
rlabel pdiffusion 570 -421 570 -421 0 feedthrough
rlabel pdiffusion 577 -421 577 -421 0 feedthrough
rlabel pdiffusion 584 -421 584 -421 0 feedthrough
rlabel pdiffusion 612 -421 612 -421 0 feedthrough
rlabel pdiffusion 3 -498 3 -498 0 feedthrough
rlabel pdiffusion 10 -498 10 -498 0 feedthrough
rlabel pdiffusion 17 -498 17 -498 0 feedthrough
rlabel pdiffusion 24 -498 24 -498 0 feedthrough
rlabel pdiffusion 31 -498 31 -498 0 feedthrough
rlabel pdiffusion 38 -498 38 -498 0 cellNo=281
rlabel pdiffusion 45 -498 45 -498 0 cellNo=676
rlabel pdiffusion 52 -498 52 -498 0 feedthrough
rlabel pdiffusion 59 -498 59 -498 0 feedthrough
rlabel pdiffusion 66 -498 66 -498 0 cellNo=66
rlabel pdiffusion 73 -498 73 -498 0 feedthrough
rlabel pdiffusion 80 -498 80 -498 0 feedthrough
rlabel pdiffusion 87 -498 87 -498 0 feedthrough
rlabel pdiffusion 94 -498 94 -498 0 feedthrough
rlabel pdiffusion 101 -498 101 -498 0 feedthrough
rlabel pdiffusion 108 -498 108 -498 0 feedthrough
rlabel pdiffusion 115 -498 115 -498 0 cellNo=338
rlabel pdiffusion 122 -498 122 -498 0 cellNo=563
rlabel pdiffusion 129 -498 129 -498 0 cellNo=313
rlabel pdiffusion 136 -498 136 -498 0 cellNo=481
rlabel pdiffusion 143 -498 143 -498 0 cellNo=316
rlabel pdiffusion 150 -498 150 -498 0 feedthrough
rlabel pdiffusion 157 -498 157 -498 0 feedthrough
rlabel pdiffusion 164 -498 164 -498 0 feedthrough
rlabel pdiffusion 171 -498 171 -498 0 cellNo=399
rlabel pdiffusion 178 -498 178 -498 0 feedthrough
rlabel pdiffusion 185 -498 185 -498 0 cellNo=329
rlabel pdiffusion 192 -498 192 -498 0 cellNo=335
rlabel pdiffusion 199 -498 199 -498 0 cellNo=699
rlabel pdiffusion 206 -498 206 -498 0 cellNo=420
rlabel pdiffusion 213 -498 213 -498 0 feedthrough
rlabel pdiffusion 220 -498 220 -498 0 feedthrough
rlabel pdiffusion 227 -498 227 -498 0 feedthrough
rlabel pdiffusion 234 -498 234 -498 0 cellNo=135
rlabel pdiffusion 241 -498 241 -498 0 cellNo=62
rlabel pdiffusion 248 -498 248 -498 0 feedthrough
rlabel pdiffusion 255 -498 255 -498 0 feedthrough
rlabel pdiffusion 262 -498 262 -498 0 cellNo=455
rlabel pdiffusion 269 -498 269 -498 0 feedthrough
rlabel pdiffusion 276 -498 276 -498 0 feedthrough
rlabel pdiffusion 283 -498 283 -498 0 feedthrough
rlabel pdiffusion 290 -498 290 -498 0 feedthrough
rlabel pdiffusion 297 -498 297 -498 0 feedthrough
rlabel pdiffusion 304 -498 304 -498 0 cellNo=211
rlabel pdiffusion 311 -498 311 -498 0 cellNo=255
rlabel pdiffusion 318 -498 318 -498 0 feedthrough
rlabel pdiffusion 325 -498 325 -498 0 cellNo=28
rlabel pdiffusion 332 -498 332 -498 0 cellNo=119
rlabel pdiffusion 339 -498 339 -498 0 feedthrough
rlabel pdiffusion 346 -498 346 -498 0 feedthrough
rlabel pdiffusion 353 -498 353 -498 0 cellNo=186
rlabel pdiffusion 360 -498 360 -498 0 cellNo=467
rlabel pdiffusion 367 -498 367 -498 0 feedthrough
rlabel pdiffusion 374 -498 374 -498 0 feedthrough
rlabel pdiffusion 381 -498 381 -498 0 feedthrough
rlabel pdiffusion 388 -498 388 -498 0 feedthrough
rlabel pdiffusion 395 -498 395 -498 0 cellNo=274
rlabel pdiffusion 402 -498 402 -498 0 feedthrough
rlabel pdiffusion 409 -498 409 -498 0 feedthrough
rlabel pdiffusion 416 -498 416 -498 0 feedthrough
rlabel pdiffusion 423 -498 423 -498 0 cellNo=267
rlabel pdiffusion 430 -498 430 -498 0 feedthrough
rlabel pdiffusion 437 -498 437 -498 0 feedthrough
rlabel pdiffusion 444 -498 444 -498 0 feedthrough
rlabel pdiffusion 451 -498 451 -498 0 feedthrough
rlabel pdiffusion 458 -498 458 -498 0 feedthrough
rlabel pdiffusion 465 -498 465 -498 0 feedthrough
rlabel pdiffusion 472 -498 472 -498 0 feedthrough
rlabel pdiffusion 479 -498 479 -498 0 feedthrough
rlabel pdiffusion 486 -498 486 -498 0 feedthrough
rlabel pdiffusion 493 -498 493 -498 0 cellNo=95
rlabel pdiffusion 500 -498 500 -498 0 feedthrough
rlabel pdiffusion 507 -498 507 -498 0 feedthrough
rlabel pdiffusion 514 -498 514 -498 0 feedthrough
rlabel pdiffusion 521 -498 521 -498 0 feedthrough
rlabel pdiffusion 528 -498 528 -498 0 feedthrough
rlabel pdiffusion 535 -498 535 -498 0 feedthrough
rlabel pdiffusion 542 -498 542 -498 0 feedthrough
rlabel pdiffusion 549 -498 549 -498 0 feedthrough
rlabel pdiffusion 556 -498 556 -498 0 feedthrough
rlabel pdiffusion 563 -498 563 -498 0 feedthrough
rlabel pdiffusion 570 -498 570 -498 0 feedthrough
rlabel pdiffusion 577 -498 577 -498 0 feedthrough
rlabel pdiffusion 584 -498 584 -498 0 feedthrough
rlabel pdiffusion 591 -498 591 -498 0 feedthrough
rlabel pdiffusion 598 -498 598 -498 0 feedthrough
rlabel pdiffusion 605 -498 605 -498 0 feedthrough
rlabel pdiffusion 612 -498 612 -498 0 feedthrough
rlabel pdiffusion 619 -498 619 -498 0 cellNo=363
rlabel pdiffusion 626 -498 626 -498 0 feedthrough
rlabel pdiffusion 633 -498 633 -498 0 cellNo=395
rlabel pdiffusion 640 -498 640 -498 0 feedthrough
rlabel pdiffusion 647 -498 647 -498 0 feedthrough
rlabel pdiffusion 654 -498 654 -498 0 cellNo=53
rlabel pdiffusion 661 -498 661 -498 0 cellNo=302
rlabel pdiffusion 668 -498 668 -498 0 feedthrough
rlabel pdiffusion 675 -498 675 -498 0 feedthrough
rlabel pdiffusion 17 -563 17 -563 0 feedthrough
rlabel pdiffusion 24 -563 24 -563 0 feedthrough
rlabel pdiffusion 31 -563 31 -563 0 feedthrough
rlabel pdiffusion 38 -563 38 -563 0 feedthrough
rlabel pdiffusion 45 -563 45 -563 0 cellNo=86
rlabel pdiffusion 52 -563 52 -563 0 feedthrough
rlabel pdiffusion 59 -563 59 -563 0 cellNo=451
rlabel pdiffusion 66 -563 66 -563 0 feedthrough
rlabel pdiffusion 73 -563 73 -563 0 cellNo=540
rlabel pdiffusion 80 -563 80 -563 0 cellNo=564
rlabel pdiffusion 87 -563 87 -563 0 feedthrough
rlabel pdiffusion 94 -563 94 -563 0 feedthrough
rlabel pdiffusion 101 -563 101 -563 0 feedthrough
rlabel pdiffusion 108 -563 108 -563 0 feedthrough
rlabel pdiffusion 115 -563 115 -563 0 feedthrough
rlabel pdiffusion 122 -563 122 -563 0 feedthrough
rlabel pdiffusion 129 -563 129 -563 0 cellNo=58
rlabel pdiffusion 136 -563 136 -563 0 feedthrough
rlabel pdiffusion 143 -563 143 -563 0 cellNo=122
rlabel pdiffusion 150 -563 150 -563 0 cellNo=498
rlabel pdiffusion 157 -563 157 -563 0 cellNo=258
rlabel pdiffusion 164 -563 164 -563 0 feedthrough
rlabel pdiffusion 171 -563 171 -563 0 cellNo=272
rlabel pdiffusion 178 -563 178 -563 0 feedthrough
rlabel pdiffusion 185 -563 185 -563 0 feedthrough
rlabel pdiffusion 192 -563 192 -563 0 cellNo=393
rlabel pdiffusion 199 -563 199 -563 0 feedthrough
rlabel pdiffusion 206 -563 206 -563 0 cellNo=36
rlabel pdiffusion 213 -563 213 -563 0 feedthrough
rlabel pdiffusion 220 -563 220 -563 0 feedthrough
rlabel pdiffusion 227 -563 227 -563 0 feedthrough
rlabel pdiffusion 234 -563 234 -563 0 feedthrough
rlabel pdiffusion 241 -563 241 -563 0 feedthrough
rlabel pdiffusion 248 -563 248 -563 0 feedthrough
rlabel pdiffusion 255 -563 255 -563 0 feedthrough
rlabel pdiffusion 262 -563 262 -563 0 cellNo=425
rlabel pdiffusion 269 -563 269 -563 0 cellNo=644
rlabel pdiffusion 276 -563 276 -563 0 cellNo=546
rlabel pdiffusion 283 -563 283 -563 0 feedthrough
rlabel pdiffusion 290 -563 290 -563 0 feedthrough
rlabel pdiffusion 297 -563 297 -563 0 feedthrough
rlabel pdiffusion 304 -563 304 -563 0 feedthrough
rlabel pdiffusion 311 -563 311 -563 0 feedthrough
rlabel pdiffusion 318 -563 318 -563 0 feedthrough
rlabel pdiffusion 325 -563 325 -563 0 feedthrough
rlabel pdiffusion 332 -563 332 -563 0 cellNo=685
rlabel pdiffusion 339 -563 339 -563 0 feedthrough
rlabel pdiffusion 346 -563 346 -563 0 cellNo=599
rlabel pdiffusion 353 -563 353 -563 0 cellNo=508
rlabel pdiffusion 360 -563 360 -563 0 feedthrough
rlabel pdiffusion 367 -563 367 -563 0 cellNo=286
rlabel pdiffusion 374 -563 374 -563 0 feedthrough
rlabel pdiffusion 381 -563 381 -563 0 cellNo=606
rlabel pdiffusion 388 -563 388 -563 0 cellNo=473
rlabel pdiffusion 395 -563 395 -563 0 cellNo=290
rlabel pdiffusion 402 -563 402 -563 0 cellNo=423
rlabel pdiffusion 409 -563 409 -563 0 cellNo=98
rlabel pdiffusion 416 -563 416 -563 0 feedthrough
rlabel pdiffusion 423 -563 423 -563 0 feedthrough
rlabel pdiffusion 430 -563 430 -563 0 feedthrough
rlabel pdiffusion 437 -563 437 -563 0 feedthrough
rlabel pdiffusion 444 -563 444 -563 0 feedthrough
rlabel pdiffusion 451 -563 451 -563 0 feedthrough
rlabel pdiffusion 458 -563 458 -563 0 feedthrough
rlabel pdiffusion 465 -563 465 -563 0 feedthrough
rlabel pdiffusion 472 -563 472 -563 0 feedthrough
rlabel pdiffusion 479 -563 479 -563 0 feedthrough
rlabel pdiffusion 486 -563 486 -563 0 cellNo=371
rlabel pdiffusion 493 -563 493 -563 0 feedthrough
rlabel pdiffusion 500 -563 500 -563 0 feedthrough
rlabel pdiffusion 507 -563 507 -563 0 feedthrough
rlabel pdiffusion 514 -563 514 -563 0 feedthrough
rlabel pdiffusion 521 -563 521 -563 0 feedthrough
rlabel pdiffusion 528 -563 528 -563 0 feedthrough
rlabel pdiffusion 535 -563 535 -563 0 feedthrough
rlabel pdiffusion 542 -563 542 -563 0 feedthrough
rlabel pdiffusion 549 -563 549 -563 0 feedthrough
rlabel pdiffusion 556 -563 556 -563 0 feedthrough
rlabel pdiffusion 563 -563 563 -563 0 feedthrough
rlabel pdiffusion 570 -563 570 -563 0 feedthrough
rlabel pdiffusion 577 -563 577 -563 0 feedthrough
rlabel pdiffusion 584 -563 584 -563 0 feedthrough
rlabel pdiffusion 591 -563 591 -563 0 feedthrough
rlabel pdiffusion 598 -563 598 -563 0 feedthrough
rlabel pdiffusion 605 -563 605 -563 0 feedthrough
rlabel pdiffusion 612 -563 612 -563 0 cellNo=305
rlabel pdiffusion 619 -563 619 -563 0 cellNo=710
rlabel pdiffusion 626 -563 626 -563 0 cellNo=703
rlabel pdiffusion 633 -563 633 -563 0 feedthrough
rlabel pdiffusion 640 -563 640 -563 0 cellNo=47
rlabel pdiffusion 647 -563 647 -563 0 feedthrough
rlabel pdiffusion 654 -563 654 -563 0 feedthrough
rlabel pdiffusion 3 -618 3 -618 0 feedthrough
rlabel pdiffusion 10 -618 10 -618 0 feedthrough
rlabel pdiffusion 17 -618 17 -618 0 feedthrough
rlabel pdiffusion 24 -618 24 -618 0 feedthrough
rlabel pdiffusion 31 -618 31 -618 0 feedthrough
rlabel pdiffusion 38 -618 38 -618 0 feedthrough
rlabel pdiffusion 45 -618 45 -618 0 feedthrough
rlabel pdiffusion 52 -618 52 -618 0 feedthrough
rlabel pdiffusion 59 -618 59 -618 0 cellNo=26
rlabel pdiffusion 66 -618 66 -618 0 cellNo=416
rlabel pdiffusion 73 -618 73 -618 0 feedthrough
rlabel pdiffusion 80 -618 80 -618 0 feedthrough
rlabel pdiffusion 87 -618 87 -618 0 feedthrough
rlabel pdiffusion 94 -618 94 -618 0 feedthrough
rlabel pdiffusion 101 -618 101 -618 0 cellNo=602
rlabel pdiffusion 108 -618 108 -618 0 feedthrough
rlabel pdiffusion 115 -618 115 -618 0 feedthrough
rlabel pdiffusion 122 -618 122 -618 0 cellNo=75
rlabel pdiffusion 129 -618 129 -618 0 cellNo=332
rlabel pdiffusion 136 -618 136 -618 0 feedthrough
rlabel pdiffusion 143 -618 143 -618 0 feedthrough
rlabel pdiffusion 150 -618 150 -618 0 cellNo=657
rlabel pdiffusion 157 -618 157 -618 0 feedthrough
rlabel pdiffusion 164 -618 164 -618 0 cellNo=414
rlabel pdiffusion 171 -618 171 -618 0 feedthrough
rlabel pdiffusion 178 -618 178 -618 0 cellNo=610
rlabel pdiffusion 185 -618 185 -618 0 cellNo=144
rlabel pdiffusion 192 -618 192 -618 0 cellNo=271
rlabel pdiffusion 199 -618 199 -618 0 cellNo=692
rlabel pdiffusion 206 -618 206 -618 0 cellNo=163
rlabel pdiffusion 213 -618 213 -618 0 feedthrough
rlabel pdiffusion 220 -618 220 -618 0 feedthrough
rlabel pdiffusion 227 -618 227 -618 0 cellNo=453
rlabel pdiffusion 234 -618 234 -618 0 feedthrough
rlabel pdiffusion 241 -618 241 -618 0 feedthrough
rlabel pdiffusion 248 -618 248 -618 0 feedthrough
rlabel pdiffusion 255 -618 255 -618 0 cellNo=164
rlabel pdiffusion 262 -618 262 -618 0 feedthrough
rlabel pdiffusion 269 -618 269 -618 0 feedthrough
rlabel pdiffusion 276 -618 276 -618 0 cellNo=595
rlabel pdiffusion 283 -618 283 -618 0 feedthrough
rlabel pdiffusion 290 -618 290 -618 0 feedthrough
rlabel pdiffusion 297 -618 297 -618 0 feedthrough
rlabel pdiffusion 304 -618 304 -618 0 feedthrough
rlabel pdiffusion 311 -618 311 -618 0 cellNo=229
rlabel pdiffusion 318 -618 318 -618 0 feedthrough
rlabel pdiffusion 325 -618 325 -618 0 cellNo=79
rlabel pdiffusion 332 -618 332 -618 0 cellNo=152
rlabel pdiffusion 339 -618 339 -618 0 feedthrough
rlabel pdiffusion 346 -618 346 -618 0 cellNo=93
rlabel pdiffusion 353 -618 353 -618 0 cellNo=146
rlabel pdiffusion 360 -618 360 -618 0 cellNo=694
rlabel pdiffusion 367 -618 367 -618 0 feedthrough
rlabel pdiffusion 374 -618 374 -618 0 feedthrough
rlabel pdiffusion 381 -618 381 -618 0 feedthrough
rlabel pdiffusion 388 -618 388 -618 0 feedthrough
rlabel pdiffusion 395 -618 395 -618 0 feedthrough
rlabel pdiffusion 402 -618 402 -618 0 cellNo=238
rlabel pdiffusion 409 -618 409 -618 0 feedthrough
rlabel pdiffusion 416 -618 416 -618 0 feedthrough
rlabel pdiffusion 423 -618 423 -618 0 feedthrough
rlabel pdiffusion 430 -618 430 -618 0 feedthrough
rlabel pdiffusion 437 -618 437 -618 0 feedthrough
rlabel pdiffusion 444 -618 444 -618 0 feedthrough
rlabel pdiffusion 451 -618 451 -618 0 feedthrough
rlabel pdiffusion 458 -618 458 -618 0 cellNo=515
rlabel pdiffusion 465 -618 465 -618 0 feedthrough
rlabel pdiffusion 472 -618 472 -618 0 feedthrough
rlabel pdiffusion 479 -618 479 -618 0 cellNo=635
rlabel pdiffusion 486 -618 486 -618 0 feedthrough
rlabel pdiffusion 493 -618 493 -618 0 feedthrough
rlabel pdiffusion 500 -618 500 -618 0 feedthrough
rlabel pdiffusion 507 -618 507 -618 0 feedthrough
rlabel pdiffusion 514 -618 514 -618 0 feedthrough
rlabel pdiffusion 521 -618 521 -618 0 feedthrough
rlabel pdiffusion 528 -618 528 -618 0 cellNo=442
rlabel pdiffusion 535 -618 535 -618 0 feedthrough
rlabel pdiffusion 542 -618 542 -618 0 cellNo=628
rlabel pdiffusion 549 -618 549 -618 0 feedthrough
rlabel pdiffusion 556 -618 556 -618 0 feedthrough
rlabel pdiffusion 563 -618 563 -618 0 cellNo=424
rlabel pdiffusion 570 -618 570 -618 0 feedthrough
rlabel pdiffusion 577 -618 577 -618 0 feedthrough
rlabel pdiffusion 584 -618 584 -618 0 feedthrough
rlabel pdiffusion 591 -618 591 -618 0 feedthrough
rlabel pdiffusion 598 -618 598 -618 0 feedthrough
rlabel pdiffusion 605 -618 605 -618 0 feedthrough
rlabel pdiffusion 612 -618 612 -618 0 feedthrough
rlabel pdiffusion 619 -618 619 -618 0 feedthrough
rlabel pdiffusion 626 -618 626 -618 0 cellNo=234
rlabel pdiffusion 633 -618 633 -618 0 feedthrough
rlabel pdiffusion 654 -618 654 -618 0 feedthrough
rlabel pdiffusion 3 -683 3 -683 0 feedthrough
rlabel pdiffusion 10 -683 10 -683 0 feedthrough
rlabel pdiffusion 17 -683 17 -683 0 feedthrough
rlabel pdiffusion 24 -683 24 -683 0 cellNo=695
rlabel pdiffusion 31 -683 31 -683 0 feedthrough
rlabel pdiffusion 38 -683 38 -683 0 feedthrough
rlabel pdiffusion 45 -683 45 -683 0 feedthrough
rlabel pdiffusion 52 -683 52 -683 0 cellNo=664
rlabel pdiffusion 59 -683 59 -683 0 feedthrough
rlabel pdiffusion 66 -683 66 -683 0 feedthrough
rlabel pdiffusion 73 -683 73 -683 0 feedthrough
rlabel pdiffusion 80 -683 80 -683 0 feedthrough
rlabel pdiffusion 87 -683 87 -683 0 feedthrough
rlabel pdiffusion 94 -683 94 -683 0 cellNo=647
rlabel pdiffusion 101 -683 101 -683 0 feedthrough
rlabel pdiffusion 108 -683 108 -683 0 feedthrough
rlabel pdiffusion 115 -683 115 -683 0 cellNo=68
rlabel pdiffusion 122 -683 122 -683 0 cellNo=396
rlabel pdiffusion 129 -683 129 -683 0 cellNo=493
rlabel pdiffusion 136 -683 136 -683 0 cellNo=428
rlabel pdiffusion 143 -683 143 -683 0 feedthrough
rlabel pdiffusion 150 -683 150 -683 0 cellNo=502
rlabel pdiffusion 157 -683 157 -683 0 feedthrough
rlabel pdiffusion 164 -683 164 -683 0 feedthrough
rlabel pdiffusion 171 -683 171 -683 0 cellNo=97
rlabel pdiffusion 178 -683 178 -683 0 cellNo=133
rlabel pdiffusion 185 -683 185 -683 0 cellNo=406
rlabel pdiffusion 192 -683 192 -683 0 feedthrough
rlabel pdiffusion 199 -683 199 -683 0 cellNo=149
rlabel pdiffusion 206 -683 206 -683 0 cellNo=407
rlabel pdiffusion 213 -683 213 -683 0 feedthrough
rlabel pdiffusion 220 -683 220 -683 0 cellNo=20
rlabel pdiffusion 227 -683 227 -683 0 feedthrough
rlabel pdiffusion 234 -683 234 -683 0 feedthrough
rlabel pdiffusion 241 -683 241 -683 0 feedthrough
rlabel pdiffusion 248 -683 248 -683 0 feedthrough
rlabel pdiffusion 255 -683 255 -683 0 cellNo=466
rlabel pdiffusion 262 -683 262 -683 0 feedthrough
rlabel pdiffusion 269 -683 269 -683 0 feedthrough
rlabel pdiffusion 276 -683 276 -683 0 cellNo=471
rlabel pdiffusion 283 -683 283 -683 0 cellNo=56
rlabel pdiffusion 290 -683 290 -683 0 cellNo=433
rlabel pdiffusion 297 -683 297 -683 0 feedthrough
rlabel pdiffusion 304 -683 304 -683 0 feedthrough
rlabel pdiffusion 311 -683 311 -683 0 cellNo=40
rlabel pdiffusion 318 -683 318 -683 0 feedthrough
rlabel pdiffusion 325 -683 325 -683 0 feedthrough
rlabel pdiffusion 332 -683 332 -683 0 cellNo=348
rlabel pdiffusion 339 -683 339 -683 0 feedthrough
rlabel pdiffusion 346 -683 346 -683 0 feedthrough
rlabel pdiffusion 353 -683 353 -683 0 feedthrough
rlabel pdiffusion 360 -683 360 -683 0 feedthrough
rlabel pdiffusion 367 -683 367 -683 0 cellNo=656
rlabel pdiffusion 374 -683 374 -683 0 cellNo=328
rlabel pdiffusion 381 -683 381 -683 0 feedthrough
rlabel pdiffusion 388 -683 388 -683 0 feedthrough
rlabel pdiffusion 395 -683 395 -683 0 cellNo=43
rlabel pdiffusion 402 -683 402 -683 0 cellNo=349
rlabel pdiffusion 409 -683 409 -683 0 feedthrough
rlabel pdiffusion 416 -683 416 -683 0 feedthrough
rlabel pdiffusion 423 -683 423 -683 0 cellNo=504
rlabel pdiffusion 430 -683 430 -683 0 cellNo=650
rlabel pdiffusion 437 -683 437 -683 0 feedthrough
rlabel pdiffusion 444 -683 444 -683 0 feedthrough
rlabel pdiffusion 451 -683 451 -683 0 feedthrough
rlabel pdiffusion 458 -683 458 -683 0 feedthrough
rlabel pdiffusion 465 -683 465 -683 0 feedthrough
rlabel pdiffusion 472 -683 472 -683 0 feedthrough
rlabel pdiffusion 479 -683 479 -683 0 feedthrough
rlabel pdiffusion 486 -683 486 -683 0 feedthrough
rlabel pdiffusion 493 -683 493 -683 0 feedthrough
rlabel pdiffusion 500 -683 500 -683 0 feedthrough
rlabel pdiffusion 507 -683 507 -683 0 feedthrough
rlabel pdiffusion 514 -683 514 -683 0 feedthrough
rlabel pdiffusion 521 -683 521 -683 0 feedthrough
rlabel pdiffusion 528 -683 528 -683 0 feedthrough
rlabel pdiffusion 535 -683 535 -683 0 feedthrough
rlabel pdiffusion 542 -683 542 -683 0 feedthrough
rlabel pdiffusion 549 -683 549 -683 0 feedthrough
rlabel pdiffusion 556 -683 556 -683 0 cellNo=609
rlabel pdiffusion 563 -683 563 -683 0 cellNo=13
rlabel pdiffusion 633 -683 633 -683 0 feedthrough
rlabel pdiffusion 640 -683 640 -683 0 cellNo=311
rlabel pdiffusion 654 -683 654 -683 0 feedthrough
rlabel pdiffusion 3 -750 3 -750 0 feedthrough
rlabel pdiffusion 10 -750 10 -750 0 cellNo=541
rlabel pdiffusion 17 -750 17 -750 0 cellNo=217
rlabel pdiffusion 24 -750 24 -750 0 cellNo=419
rlabel pdiffusion 31 -750 31 -750 0 feedthrough
rlabel pdiffusion 38 -750 38 -750 0 feedthrough
rlabel pdiffusion 45 -750 45 -750 0 cellNo=284
rlabel pdiffusion 52 -750 52 -750 0 feedthrough
rlabel pdiffusion 59 -750 59 -750 0 cellNo=351
rlabel pdiffusion 66 -750 66 -750 0 feedthrough
rlabel pdiffusion 73 -750 73 -750 0 feedthrough
rlabel pdiffusion 80 -750 80 -750 0 cellNo=109
rlabel pdiffusion 87 -750 87 -750 0 feedthrough
rlabel pdiffusion 94 -750 94 -750 0 feedthrough
rlabel pdiffusion 101 -750 101 -750 0 cellNo=579
rlabel pdiffusion 108 -750 108 -750 0 feedthrough
rlabel pdiffusion 115 -750 115 -750 0 cellNo=131
rlabel pdiffusion 122 -750 122 -750 0 feedthrough
rlabel pdiffusion 129 -750 129 -750 0 feedthrough
rlabel pdiffusion 136 -750 136 -750 0 feedthrough
rlabel pdiffusion 143 -750 143 -750 0 cellNo=457
rlabel pdiffusion 150 -750 150 -750 0 cellNo=166
rlabel pdiffusion 157 -750 157 -750 0 feedthrough
rlabel pdiffusion 164 -750 164 -750 0 cellNo=233
rlabel pdiffusion 171 -750 171 -750 0 feedthrough
rlabel pdiffusion 178 -750 178 -750 0 feedthrough
rlabel pdiffusion 185 -750 185 -750 0 cellNo=101
rlabel pdiffusion 192 -750 192 -750 0 cellNo=223
rlabel pdiffusion 199 -750 199 -750 0 cellNo=179
rlabel pdiffusion 206 -750 206 -750 0 cellNo=38
rlabel pdiffusion 213 -750 213 -750 0 feedthrough
rlabel pdiffusion 220 -750 220 -750 0 feedthrough
rlabel pdiffusion 227 -750 227 -750 0 cellNo=388
rlabel pdiffusion 234 -750 234 -750 0 feedthrough
rlabel pdiffusion 241 -750 241 -750 0 feedthrough
rlabel pdiffusion 248 -750 248 -750 0 feedthrough
rlabel pdiffusion 255 -750 255 -750 0 feedthrough
rlabel pdiffusion 262 -750 262 -750 0 cellNo=557
rlabel pdiffusion 269 -750 269 -750 0 cellNo=376
rlabel pdiffusion 276 -750 276 -750 0 cellNo=49
rlabel pdiffusion 283 -750 283 -750 0 cellNo=645
rlabel pdiffusion 290 -750 290 -750 0 feedthrough
rlabel pdiffusion 297 -750 297 -750 0 feedthrough
rlabel pdiffusion 304 -750 304 -750 0 cellNo=252
rlabel pdiffusion 311 -750 311 -750 0 feedthrough
rlabel pdiffusion 318 -750 318 -750 0 feedthrough
rlabel pdiffusion 325 -750 325 -750 0 feedthrough
rlabel pdiffusion 332 -750 332 -750 0 feedthrough
rlabel pdiffusion 339 -750 339 -750 0 cellNo=236
rlabel pdiffusion 346 -750 346 -750 0 feedthrough
rlabel pdiffusion 353 -750 353 -750 0 cellNo=382
rlabel pdiffusion 360 -750 360 -750 0 cellNo=151
rlabel pdiffusion 367 -750 367 -750 0 feedthrough
rlabel pdiffusion 374 -750 374 -750 0 cellNo=294
rlabel pdiffusion 381 -750 381 -750 0 cellNo=353
rlabel pdiffusion 388 -750 388 -750 0 feedthrough
rlabel pdiffusion 395 -750 395 -750 0 feedthrough
rlabel pdiffusion 402 -750 402 -750 0 feedthrough
rlabel pdiffusion 409 -750 409 -750 0 cellNo=523
rlabel pdiffusion 416 -750 416 -750 0 feedthrough
rlabel pdiffusion 423 -750 423 -750 0 feedthrough
rlabel pdiffusion 430 -750 430 -750 0 feedthrough
rlabel pdiffusion 437 -750 437 -750 0 feedthrough
rlabel pdiffusion 444 -750 444 -750 0 feedthrough
rlabel pdiffusion 451 -750 451 -750 0 feedthrough
rlabel pdiffusion 458 -750 458 -750 0 feedthrough
rlabel pdiffusion 465 -750 465 -750 0 feedthrough
rlabel pdiffusion 472 -750 472 -750 0 cellNo=680
rlabel pdiffusion 479 -750 479 -750 0 feedthrough
rlabel pdiffusion 486 -750 486 -750 0 feedthrough
rlabel pdiffusion 493 -750 493 -750 0 feedthrough
rlabel pdiffusion 500 -750 500 -750 0 feedthrough
rlabel pdiffusion 507 -750 507 -750 0 feedthrough
rlabel pdiffusion 514 -750 514 -750 0 feedthrough
rlabel pdiffusion 521 -750 521 -750 0 feedthrough
rlabel pdiffusion 528 -750 528 -750 0 feedthrough
rlabel pdiffusion 535 -750 535 -750 0 feedthrough
rlabel pdiffusion 542 -750 542 -750 0 feedthrough
rlabel pdiffusion 549 -750 549 -750 0 feedthrough
rlabel pdiffusion 556 -750 556 -750 0 feedthrough
rlabel pdiffusion 563 -750 563 -750 0 feedthrough
rlabel pdiffusion 570 -750 570 -750 0 feedthrough
rlabel pdiffusion 577 -750 577 -750 0 feedthrough
rlabel pdiffusion 584 -750 584 -750 0 feedthrough
rlabel pdiffusion 591 -750 591 -750 0 feedthrough
rlabel pdiffusion 598 -750 598 -750 0 feedthrough
rlabel pdiffusion 605 -750 605 -750 0 feedthrough
rlabel pdiffusion 612 -750 612 -750 0 feedthrough
rlabel pdiffusion 619 -750 619 -750 0 feedthrough
rlabel pdiffusion 626 -750 626 -750 0 feedthrough
rlabel pdiffusion 633 -750 633 -750 0 feedthrough
rlabel pdiffusion 640 -750 640 -750 0 feedthrough
rlabel pdiffusion 647 -750 647 -750 0 feedthrough
rlabel pdiffusion 654 -750 654 -750 0 cellNo=677
rlabel pdiffusion 661 -750 661 -750 0 cellNo=494
rlabel pdiffusion 24 -823 24 -823 0 feedthrough
rlabel pdiffusion 31 -823 31 -823 0 feedthrough
rlabel pdiffusion 38 -823 38 -823 0 cellNo=202
rlabel pdiffusion 45 -823 45 -823 0 feedthrough
rlabel pdiffusion 52 -823 52 -823 0 cellNo=337
rlabel pdiffusion 59 -823 59 -823 0 feedthrough
rlabel pdiffusion 66 -823 66 -823 0 feedthrough
rlabel pdiffusion 73 -823 73 -823 0 feedthrough
rlabel pdiffusion 80 -823 80 -823 0 cellNo=489
rlabel pdiffusion 87 -823 87 -823 0 cellNo=632
rlabel pdiffusion 94 -823 94 -823 0 cellNo=592
rlabel pdiffusion 101 -823 101 -823 0 feedthrough
rlabel pdiffusion 108 -823 108 -823 0 feedthrough
rlabel pdiffusion 115 -823 115 -823 0 feedthrough
rlabel pdiffusion 122 -823 122 -823 0 feedthrough
rlabel pdiffusion 129 -823 129 -823 0 cellNo=397
rlabel pdiffusion 136 -823 136 -823 0 cellNo=296
rlabel pdiffusion 143 -823 143 -823 0 cellNo=127
rlabel pdiffusion 150 -823 150 -823 0 cellNo=582
rlabel pdiffusion 157 -823 157 -823 0 feedthrough
rlabel pdiffusion 164 -823 164 -823 0 feedthrough
rlabel pdiffusion 171 -823 171 -823 0 feedthrough
rlabel pdiffusion 178 -823 178 -823 0 feedthrough
rlabel pdiffusion 185 -823 185 -823 0 feedthrough
rlabel pdiffusion 192 -823 192 -823 0 feedthrough
rlabel pdiffusion 199 -823 199 -823 0 feedthrough
rlabel pdiffusion 206 -823 206 -823 0 feedthrough
rlabel pdiffusion 213 -823 213 -823 0 feedthrough
rlabel pdiffusion 220 -823 220 -823 0 feedthrough
rlabel pdiffusion 227 -823 227 -823 0 feedthrough
rlabel pdiffusion 234 -823 234 -823 0 feedthrough
rlabel pdiffusion 241 -823 241 -823 0 cellNo=361
rlabel pdiffusion 248 -823 248 -823 0 feedthrough
rlabel pdiffusion 255 -823 255 -823 0 feedthrough
rlabel pdiffusion 262 -823 262 -823 0 feedthrough
rlabel pdiffusion 269 -823 269 -823 0 feedthrough
rlabel pdiffusion 276 -823 276 -823 0 cellNo=260
rlabel pdiffusion 283 -823 283 -823 0 cellNo=485
rlabel pdiffusion 290 -823 290 -823 0 feedthrough
rlabel pdiffusion 297 -823 297 -823 0 cellNo=625
rlabel pdiffusion 304 -823 304 -823 0 feedthrough
rlabel pdiffusion 311 -823 311 -823 0 cellNo=285
rlabel pdiffusion 318 -823 318 -823 0 cellNo=619
rlabel pdiffusion 325 -823 325 -823 0 cellNo=551
rlabel pdiffusion 332 -823 332 -823 0 cellNo=682
rlabel pdiffusion 339 -823 339 -823 0 cellNo=78
rlabel pdiffusion 346 -823 346 -823 0 feedthrough
rlabel pdiffusion 353 -823 353 -823 0 cellNo=434
rlabel pdiffusion 360 -823 360 -823 0 feedthrough
rlabel pdiffusion 367 -823 367 -823 0 feedthrough
rlabel pdiffusion 374 -823 374 -823 0 cellNo=417
rlabel pdiffusion 381 -823 381 -823 0 feedthrough
rlabel pdiffusion 388 -823 388 -823 0 cellNo=668
rlabel pdiffusion 395 -823 395 -823 0 feedthrough
rlabel pdiffusion 402 -823 402 -823 0 cellNo=575
rlabel pdiffusion 409 -823 409 -823 0 feedthrough
rlabel pdiffusion 416 -823 416 -823 0 feedthrough
rlabel pdiffusion 423 -823 423 -823 0 feedthrough
rlabel pdiffusion 430 -823 430 -823 0 feedthrough
rlabel pdiffusion 437 -823 437 -823 0 feedthrough
rlabel pdiffusion 444 -823 444 -823 0 feedthrough
rlabel pdiffusion 451 -823 451 -823 0 feedthrough
rlabel pdiffusion 458 -823 458 -823 0 feedthrough
rlabel pdiffusion 465 -823 465 -823 0 feedthrough
rlabel pdiffusion 472 -823 472 -823 0 feedthrough
rlabel pdiffusion 479 -823 479 -823 0 cellNo=342
rlabel pdiffusion 486 -823 486 -823 0 feedthrough
rlabel pdiffusion 493 -823 493 -823 0 feedthrough
rlabel pdiffusion 500 -823 500 -823 0 feedthrough
rlabel pdiffusion 507 -823 507 -823 0 feedthrough
rlabel pdiffusion 514 -823 514 -823 0 cellNo=115
rlabel pdiffusion 521 -823 521 -823 0 feedthrough
rlabel pdiffusion 528 -823 528 -823 0 feedthrough
rlabel pdiffusion 535 -823 535 -823 0 cellNo=421
rlabel pdiffusion 542 -823 542 -823 0 feedthrough
rlabel pdiffusion 549 -823 549 -823 0 feedthrough
rlabel pdiffusion 556 -823 556 -823 0 cellNo=570
rlabel pdiffusion 563 -823 563 -823 0 feedthrough
rlabel pdiffusion 570 -823 570 -823 0 cellNo=623
rlabel pdiffusion 577 -823 577 -823 0 feedthrough
rlabel pdiffusion 584 -823 584 -823 0 feedthrough
rlabel pdiffusion 591 -823 591 -823 0 feedthrough
rlabel pdiffusion 598 -823 598 -823 0 cellNo=10
rlabel pdiffusion 605 -823 605 -823 0 feedthrough
rlabel pdiffusion 619 -823 619 -823 0 feedthrough
rlabel pdiffusion 3 -866 3 -866 0 feedthrough
rlabel pdiffusion 10 -866 10 -866 0 feedthrough
rlabel pdiffusion 17 -866 17 -866 0 feedthrough
rlabel pdiffusion 24 -866 24 -866 0 feedthrough
rlabel pdiffusion 31 -866 31 -866 0 cellNo=514
rlabel pdiffusion 38 -866 38 -866 0 cellNo=459
rlabel pdiffusion 45 -866 45 -866 0 cellNo=73
rlabel pdiffusion 52 -866 52 -866 0 feedthrough
rlabel pdiffusion 59 -866 59 -866 0 cellNo=121
rlabel pdiffusion 66 -866 66 -866 0 feedthrough
rlabel pdiffusion 73 -866 73 -866 0 feedthrough
rlabel pdiffusion 80 -866 80 -866 0 cellNo=279
rlabel pdiffusion 87 -866 87 -866 0 feedthrough
rlabel pdiffusion 94 -866 94 -866 0 feedthrough
rlabel pdiffusion 101 -866 101 -866 0 feedthrough
rlabel pdiffusion 108 -866 108 -866 0 feedthrough
rlabel pdiffusion 115 -866 115 -866 0 feedthrough
rlabel pdiffusion 122 -866 122 -866 0 feedthrough
rlabel pdiffusion 129 -866 129 -866 0 feedthrough
rlabel pdiffusion 136 -866 136 -866 0 cellNo=478
rlabel pdiffusion 143 -866 143 -866 0 cellNo=669
rlabel pdiffusion 150 -866 150 -866 0 feedthrough
rlabel pdiffusion 157 -866 157 -866 0 feedthrough
rlabel pdiffusion 164 -866 164 -866 0 cellNo=278
rlabel pdiffusion 171 -866 171 -866 0 cellNo=690
rlabel pdiffusion 178 -866 178 -866 0 cellNo=176
rlabel pdiffusion 185 -866 185 -866 0 feedthrough
rlabel pdiffusion 192 -866 192 -866 0 cellNo=627
rlabel pdiffusion 199 -866 199 -866 0 cellNo=643
rlabel pdiffusion 206 -866 206 -866 0 cellNo=674
rlabel pdiffusion 213 -866 213 -866 0 cellNo=509
rlabel pdiffusion 220 -866 220 -866 0 cellNo=319
rlabel pdiffusion 227 -866 227 -866 0 cellNo=162
rlabel pdiffusion 234 -866 234 -866 0 feedthrough
rlabel pdiffusion 241 -866 241 -866 0 feedthrough
rlabel pdiffusion 248 -866 248 -866 0 feedthrough
rlabel pdiffusion 255 -866 255 -866 0 feedthrough
rlabel pdiffusion 262 -866 262 -866 0 cellNo=576
rlabel pdiffusion 269 -866 269 -866 0 feedthrough
rlabel pdiffusion 276 -866 276 -866 0 feedthrough
rlabel pdiffusion 283 -866 283 -866 0 feedthrough
rlabel pdiffusion 290 -866 290 -866 0 cellNo=312
rlabel pdiffusion 297 -866 297 -866 0 feedthrough
rlabel pdiffusion 304 -866 304 -866 0 feedthrough
rlabel pdiffusion 311 -866 311 -866 0 feedthrough
rlabel pdiffusion 318 -866 318 -866 0 cellNo=369
rlabel pdiffusion 325 -866 325 -866 0 feedthrough
rlabel pdiffusion 332 -866 332 -866 0 feedthrough
rlabel pdiffusion 339 -866 339 -866 0 feedthrough
rlabel pdiffusion 346 -866 346 -866 0 cellNo=216
rlabel pdiffusion 353 -866 353 -866 0 feedthrough
rlabel pdiffusion 360 -866 360 -866 0 feedthrough
rlabel pdiffusion 367 -866 367 -866 0 feedthrough
rlabel pdiffusion 374 -866 374 -866 0 cellNo=323
rlabel pdiffusion 381 -866 381 -866 0 cellNo=1
rlabel pdiffusion 388 -866 388 -866 0 feedthrough
rlabel pdiffusion 395 -866 395 -866 0 feedthrough
rlabel pdiffusion 402 -866 402 -866 0 feedthrough
rlabel pdiffusion 409 -866 409 -866 0 feedthrough
rlabel pdiffusion 416 -866 416 -866 0 feedthrough
rlabel pdiffusion 423 -866 423 -866 0 cellNo=326
rlabel pdiffusion 430 -866 430 -866 0 feedthrough
rlabel pdiffusion 437 -866 437 -866 0 feedthrough
rlabel pdiffusion 444 -866 444 -866 0 feedthrough
rlabel pdiffusion 451 -866 451 -866 0 cellNo=268
rlabel pdiffusion 458 -866 458 -866 0 feedthrough
rlabel pdiffusion 465 -866 465 -866 0 feedthrough
rlabel pdiffusion 472 -866 472 -866 0 feedthrough
rlabel pdiffusion 479 -866 479 -866 0 feedthrough
rlabel pdiffusion 486 -866 486 -866 0 feedthrough
rlabel pdiffusion 493 -866 493 -866 0 feedthrough
rlabel pdiffusion 500 -866 500 -866 0 feedthrough
rlabel pdiffusion 507 -866 507 -866 0 feedthrough
rlabel pdiffusion 514 -866 514 -866 0 cellNo=708
rlabel pdiffusion 521 -866 521 -866 0 feedthrough
rlabel pdiffusion 528 -866 528 -866 0 cellNo=262
rlabel pdiffusion 535 -866 535 -866 0 cellNo=418
rlabel pdiffusion 542 -866 542 -866 0 cellNo=477
rlabel pdiffusion 549 -866 549 -866 0 cellNo=465
rlabel pdiffusion 556 -866 556 -866 0 feedthrough
rlabel pdiffusion 563 -866 563 -866 0 feedthrough
rlabel pdiffusion 3 -921 3 -921 0 feedthrough
rlabel pdiffusion 10 -921 10 -921 0 cellNo=588
rlabel pdiffusion 17 -921 17 -921 0 feedthrough
rlabel pdiffusion 24 -921 24 -921 0 feedthrough
rlabel pdiffusion 31 -921 31 -921 0 cellNo=199
rlabel pdiffusion 38 -921 38 -921 0 cellNo=7
rlabel pdiffusion 45 -921 45 -921 0 cellNo=175
rlabel pdiffusion 52 -921 52 -921 0 cellNo=46
rlabel pdiffusion 59 -921 59 -921 0 cellNo=456
rlabel pdiffusion 66 -921 66 -921 0 cellNo=372
rlabel pdiffusion 73 -921 73 -921 0 cellNo=300
rlabel pdiffusion 80 -921 80 -921 0 feedthrough
rlabel pdiffusion 87 -921 87 -921 0 feedthrough
rlabel pdiffusion 94 -921 94 -921 0 cellNo=160
rlabel pdiffusion 101 -921 101 -921 0 cellNo=706
rlabel pdiffusion 108 -921 108 -921 0 cellNo=450
rlabel pdiffusion 115 -921 115 -921 0 feedthrough
rlabel pdiffusion 122 -921 122 -921 0 cellNo=479
rlabel pdiffusion 129 -921 129 -921 0 cellNo=12
rlabel pdiffusion 136 -921 136 -921 0 feedthrough
rlabel pdiffusion 143 -921 143 -921 0 feedthrough
rlabel pdiffusion 150 -921 150 -921 0 cellNo=275
rlabel pdiffusion 157 -921 157 -921 0 feedthrough
rlabel pdiffusion 164 -921 164 -921 0 feedthrough
rlabel pdiffusion 171 -921 171 -921 0 cellNo=27
rlabel pdiffusion 178 -921 178 -921 0 cellNo=259
rlabel pdiffusion 185 -921 185 -921 0 cellNo=400
rlabel pdiffusion 192 -921 192 -921 0 cellNo=48
rlabel pdiffusion 199 -921 199 -921 0 cellNo=693
rlabel pdiffusion 206 -921 206 -921 0 cellNo=378
rlabel pdiffusion 213 -921 213 -921 0 feedthrough
rlabel pdiffusion 220 -921 220 -921 0 feedthrough
rlabel pdiffusion 227 -921 227 -921 0 cellNo=324
rlabel pdiffusion 234 -921 234 -921 0 feedthrough
rlabel pdiffusion 241 -921 241 -921 0 cellNo=468
rlabel pdiffusion 248 -921 248 -921 0 feedthrough
rlabel pdiffusion 255 -921 255 -921 0 feedthrough
rlabel pdiffusion 262 -921 262 -921 0 feedthrough
rlabel pdiffusion 269 -921 269 -921 0 feedthrough
rlabel pdiffusion 276 -921 276 -921 0 feedthrough
rlabel pdiffusion 283 -921 283 -921 0 feedthrough
rlabel pdiffusion 290 -921 290 -921 0 cellNo=527
rlabel pdiffusion 297 -921 297 -921 0 cellNo=469
rlabel pdiffusion 304 -921 304 -921 0 cellNo=327
rlabel pdiffusion 311 -921 311 -921 0 cellNo=173
rlabel pdiffusion 318 -921 318 -921 0 feedthrough
rlabel pdiffusion 325 -921 325 -921 0 feedthrough
rlabel pdiffusion 332 -921 332 -921 0 feedthrough
rlabel pdiffusion 339 -921 339 -921 0 feedthrough
rlabel pdiffusion 346 -921 346 -921 0 feedthrough
rlabel pdiffusion 353 -921 353 -921 0 feedthrough
rlabel pdiffusion 360 -921 360 -921 0 cellNo=673
rlabel pdiffusion 367 -921 367 -921 0 feedthrough
rlabel pdiffusion 374 -921 374 -921 0 feedthrough
rlabel pdiffusion 381 -921 381 -921 0 feedthrough
rlabel pdiffusion 388 -921 388 -921 0 feedthrough
rlabel pdiffusion 395 -921 395 -921 0 feedthrough
rlabel pdiffusion 402 -921 402 -921 0 feedthrough
rlabel pdiffusion 409 -921 409 -921 0 feedthrough
rlabel pdiffusion 416 -921 416 -921 0 feedthrough
rlabel pdiffusion 423 -921 423 -921 0 feedthrough
rlabel pdiffusion 430 -921 430 -921 0 feedthrough
rlabel pdiffusion 437 -921 437 -921 0 feedthrough
rlabel pdiffusion 444 -921 444 -921 0 cellNo=443
rlabel pdiffusion 451 -921 451 -921 0 feedthrough
rlabel pdiffusion 458 -921 458 -921 0 feedthrough
rlabel pdiffusion 465 -921 465 -921 0 feedthrough
rlabel pdiffusion 472 -921 472 -921 0 cellNo=711
rlabel pdiffusion 479 -921 479 -921 0 feedthrough
rlabel pdiffusion 486 -921 486 -921 0 feedthrough
rlabel pdiffusion 493 -921 493 -921 0 feedthrough
rlabel pdiffusion 500 -921 500 -921 0 feedthrough
rlabel pdiffusion 507 -921 507 -921 0 feedthrough
rlabel pdiffusion 514 -921 514 -921 0 feedthrough
rlabel pdiffusion 521 -921 521 -921 0 feedthrough
rlabel pdiffusion 528 -921 528 -921 0 cellNo=431
rlabel pdiffusion 535 -921 535 -921 0 feedthrough
rlabel pdiffusion 542 -921 542 -921 0 feedthrough
rlabel pdiffusion 549 -921 549 -921 0 feedthrough
rlabel pdiffusion 24 -974 24 -974 0 feedthrough
rlabel pdiffusion 31 -974 31 -974 0 feedthrough
rlabel pdiffusion 38 -974 38 -974 0 cellNo=472
rlabel pdiffusion 45 -974 45 -974 0 cellNo=480
rlabel pdiffusion 52 -974 52 -974 0 cellNo=470
rlabel pdiffusion 59 -974 59 -974 0 feedthrough
rlabel pdiffusion 66 -974 66 -974 0 cellNo=401
rlabel pdiffusion 73 -974 73 -974 0 feedthrough
rlabel pdiffusion 80 -974 80 -974 0 feedthrough
rlabel pdiffusion 87 -974 87 -974 0 feedthrough
rlabel pdiffusion 94 -974 94 -974 0 feedthrough
rlabel pdiffusion 101 -974 101 -974 0 feedthrough
rlabel pdiffusion 108 -974 108 -974 0 cellNo=461
rlabel pdiffusion 115 -974 115 -974 0 cellNo=651
rlabel pdiffusion 122 -974 122 -974 0 feedthrough
rlabel pdiffusion 129 -974 129 -974 0 cellNo=578
rlabel pdiffusion 136 -974 136 -974 0 feedthrough
rlabel pdiffusion 143 -974 143 -974 0 cellNo=437
rlabel pdiffusion 150 -974 150 -974 0 cellNo=218
rlabel pdiffusion 157 -974 157 -974 0 feedthrough
rlabel pdiffusion 164 -974 164 -974 0 cellNo=136
rlabel pdiffusion 171 -974 171 -974 0 feedthrough
rlabel pdiffusion 178 -974 178 -974 0 feedthrough
rlabel pdiffusion 185 -974 185 -974 0 cellNo=440
rlabel pdiffusion 192 -974 192 -974 0 feedthrough
rlabel pdiffusion 199 -974 199 -974 0 cellNo=713
rlabel pdiffusion 206 -974 206 -974 0 cellNo=545
rlabel pdiffusion 213 -974 213 -974 0 feedthrough
rlabel pdiffusion 220 -974 220 -974 0 feedthrough
rlabel pdiffusion 227 -974 227 -974 0 cellNo=503
rlabel pdiffusion 234 -974 234 -974 0 cellNo=594
rlabel pdiffusion 241 -974 241 -974 0 feedthrough
rlabel pdiffusion 248 -974 248 -974 0 feedthrough
rlabel pdiffusion 255 -974 255 -974 0 feedthrough
rlabel pdiffusion 262 -974 262 -974 0 cellNo=265
rlabel pdiffusion 269 -974 269 -974 0 feedthrough
rlabel pdiffusion 276 -974 276 -974 0 cellNo=641
rlabel pdiffusion 283 -974 283 -974 0 cellNo=288
rlabel pdiffusion 290 -974 290 -974 0 feedthrough
rlabel pdiffusion 297 -974 297 -974 0 cellNo=597
rlabel pdiffusion 304 -974 304 -974 0 feedthrough
rlabel pdiffusion 311 -974 311 -974 0 feedthrough
rlabel pdiffusion 318 -974 318 -974 0 cellNo=691
rlabel pdiffusion 325 -974 325 -974 0 feedthrough
rlabel pdiffusion 332 -974 332 -974 0 feedthrough
rlabel pdiffusion 339 -974 339 -974 0 feedthrough
rlabel pdiffusion 346 -974 346 -974 0 feedthrough
rlabel pdiffusion 353 -974 353 -974 0 cellNo=512
rlabel pdiffusion 360 -974 360 -974 0 feedthrough
rlabel pdiffusion 367 -974 367 -974 0 feedthrough
rlabel pdiffusion 374 -974 374 -974 0 feedthrough
rlabel pdiffusion 381 -974 381 -974 0 cellNo=435
rlabel pdiffusion 388 -974 388 -974 0 feedthrough
rlabel pdiffusion 395 -974 395 -974 0 feedthrough
rlabel pdiffusion 402 -974 402 -974 0 feedthrough
rlabel pdiffusion 409 -974 409 -974 0 cellNo=147
rlabel pdiffusion 416 -974 416 -974 0 feedthrough
rlabel pdiffusion 423 -974 423 -974 0 cellNo=671
rlabel pdiffusion 430 -974 430 -974 0 feedthrough
rlabel pdiffusion 437 -974 437 -974 0 feedthrough
rlabel pdiffusion 444 -974 444 -974 0 feedthrough
rlabel pdiffusion 451 -974 451 -974 0 feedthrough
rlabel pdiffusion 458 -974 458 -974 0 feedthrough
rlabel pdiffusion 465 -974 465 -974 0 cellNo=167
rlabel pdiffusion 472 -974 472 -974 0 feedthrough
rlabel pdiffusion 479 -974 479 -974 0 cellNo=665
rlabel pdiffusion 486 -974 486 -974 0 cellNo=389
rlabel pdiffusion 493 -974 493 -974 0 feedthrough
rlabel pdiffusion 500 -974 500 -974 0 feedthrough
rlabel pdiffusion 507 -974 507 -974 0 cellNo=385
rlabel pdiffusion 521 -974 521 -974 0 feedthrough
rlabel pdiffusion 17 -1015 17 -1015 0 feedthrough
rlabel pdiffusion 24 -1015 24 -1015 0 cellNo=22
rlabel pdiffusion 31 -1015 31 -1015 0 feedthrough
rlabel pdiffusion 38 -1015 38 -1015 0 feedthrough
rlabel pdiffusion 45 -1015 45 -1015 0 cellNo=241
rlabel pdiffusion 52 -1015 52 -1015 0 feedthrough
rlabel pdiffusion 59 -1015 59 -1015 0 feedthrough
rlabel pdiffusion 66 -1015 66 -1015 0 cellNo=308
rlabel pdiffusion 73 -1015 73 -1015 0 feedthrough
rlabel pdiffusion 80 -1015 80 -1015 0 feedthrough
rlabel pdiffusion 87 -1015 87 -1015 0 cellNo=318
rlabel pdiffusion 94 -1015 94 -1015 0 cellNo=264
rlabel pdiffusion 101 -1015 101 -1015 0 feedthrough
rlabel pdiffusion 108 -1015 108 -1015 0 feedthrough
rlabel pdiffusion 115 -1015 115 -1015 0 cellNo=200
rlabel pdiffusion 122 -1015 122 -1015 0 feedthrough
rlabel pdiffusion 129 -1015 129 -1015 0 cellNo=630
rlabel pdiffusion 136 -1015 136 -1015 0 feedthrough
rlabel pdiffusion 143 -1015 143 -1015 0 feedthrough
rlabel pdiffusion 150 -1015 150 -1015 0 feedthrough
rlabel pdiffusion 157 -1015 157 -1015 0 feedthrough
rlabel pdiffusion 164 -1015 164 -1015 0 feedthrough
rlabel pdiffusion 171 -1015 171 -1015 0 cellNo=526
rlabel pdiffusion 178 -1015 178 -1015 0 feedthrough
rlabel pdiffusion 185 -1015 185 -1015 0 cellNo=203
rlabel pdiffusion 192 -1015 192 -1015 0 cellNo=5
rlabel pdiffusion 199 -1015 199 -1015 0 cellNo=492
rlabel pdiffusion 206 -1015 206 -1015 0 cellNo=531
rlabel pdiffusion 213 -1015 213 -1015 0 feedthrough
rlabel pdiffusion 220 -1015 220 -1015 0 feedthrough
rlabel pdiffusion 227 -1015 227 -1015 0 cellNo=269
rlabel pdiffusion 234 -1015 234 -1015 0 cellNo=430
rlabel pdiffusion 241 -1015 241 -1015 0 feedthrough
rlabel pdiffusion 248 -1015 248 -1015 0 feedthrough
rlabel pdiffusion 255 -1015 255 -1015 0 feedthrough
rlabel pdiffusion 262 -1015 262 -1015 0 feedthrough
rlabel pdiffusion 269 -1015 269 -1015 0 cellNo=125
rlabel pdiffusion 276 -1015 276 -1015 0 cellNo=617
rlabel pdiffusion 283 -1015 283 -1015 0 cellNo=586
rlabel pdiffusion 290 -1015 290 -1015 0 cellNo=601
rlabel pdiffusion 297 -1015 297 -1015 0 cellNo=697
rlabel pdiffusion 304 -1015 304 -1015 0 feedthrough
rlabel pdiffusion 311 -1015 311 -1015 0 feedthrough
rlabel pdiffusion 318 -1015 318 -1015 0 feedthrough
rlabel pdiffusion 325 -1015 325 -1015 0 cellNo=145
rlabel pdiffusion 332 -1015 332 -1015 0 feedthrough
rlabel pdiffusion 339 -1015 339 -1015 0 feedthrough
rlabel pdiffusion 346 -1015 346 -1015 0 feedthrough
rlabel pdiffusion 353 -1015 353 -1015 0 feedthrough
rlabel pdiffusion 360 -1015 360 -1015 0 feedthrough
rlabel pdiffusion 367 -1015 367 -1015 0 cellNo=537
rlabel pdiffusion 374 -1015 374 -1015 0 feedthrough
rlabel pdiffusion 381 -1015 381 -1015 0 feedthrough
rlabel pdiffusion 388 -1015 388 -1015 0 cellNo=444
rlabel pdiffusion 395 -1015 395 -1015 0 feedthrough
rlabel pdiffusion 402 -1015 402 -1015 0 feedthrough
rlabel pdiffusion 409 -1015 409 -1015 0 feedthrough
rlabel pdiffusion 416 -1015 416 -1015 0 feedthrough
rlabel pdiffusion 423 -1015 423 -1015 0 feedthrough
rlabel pdiffusion 430 -1015 430 -1015 0 cellNo=542
rlabel pdiffusion 437 -1015 437 -1015 0 feedthrough
rlabel pdiffusion 444 -1015 444 -1015 0 cellNo=475
rlabel pdiffusion 451 -1015 451 -1015 0 cellNo=646
rlabel pdiffusion 458 -1015 458 -1015 0 feedthrough
rlabel pdiffusion 465 -1015 465 -1015 0 feedthrough
rlabel pdiffusion 472 -1015 472 -1015 0 feedthrough
rlabel pdiffusion 479 -1015 479 -1015 0 feedthrough
rlabel pdiffusion 521 -1015 521 -1015 0 cellNo=226
rlabel pdiffusion 528 -1015 528 -1015 0 feedthrough
rlabel pdiffusion 66 -1052 66 -1052 0 feedthrough
rlabel pdiffusion 73 -1052 73 -1052 0 feedthrough
rlabel pdiffusion 80 -1052 80 -1052 0 cellNo=689
rlabel pdiffusion 87 -1052 87 -1052 0 cellNo=150
rlabel pdiffusion 94 -1052 94 -1052 0 feedthrough
rlabel pdiffusion 101 -1052 101 -1052 0 cellNo=438
rlabel pdiffusion 108 -1052 108 -1052 0 feedthrough
rlabel pdiffusion 115 -1052 115 -1052 0 cellNo=85
rlabel pdiffusion 122 -1052 122 -1052 0 feedthrough
rlabel pdiffusion 129 -1052 129 -1052 0 feedthrough
rlabel pdiffusion 136 -1052 136 -1052 0 feedthrough
rlabel pdiffusion 143 -1052 143 -1052 0 cellNo=295
rlabel pdiffusion 150 -1052 150 -1052 0 cellNo=638
rlabel pdiffusion 157 -1052 157 -1052 0 cellNo=4
rlabel pdiffusion 164 -1052 164 -1052 0 cellNo=484
rlabel pdiffusion 171 -1052 171 -1052 0 feedthrough
rlabel pdiffusion 178 -1052 178 -1052 0 feedthrough
rlabel pdiffusion 185 -1052 185 -1052 0 feedthrough
rlabel pdiffusion 192 -1052 192 -1052 0 feedthrough
rlabel pdiffusion 199 -1052 199 -1052 0 cellNo=181
rlabel pdiffusion 206 -1052 206 -1052 0 cellNo=446
rlabel pdiffusion 213 -1052 213 -1052 0 cellNo=29
rlabel pdiffusion 220 -1052 220 -1052 0 feedthrough
rlabel pdiffusion 227 -1052 227 -1052 0 cellNo=309
rlabel pdiffusion 234 -1052 234 -1052 0 cellNo=373
rlabel pdiffusion 241 -1052 241 -1052 0 feedthrough
rlabel pdiffusion 248 -1052 248 -1052 0 cellNo=232
rlabel pdiffusion 255 -1052 255 -1052 0 cellNo=254
rlabel pdiffusion 262 -1052 262 -1052 0 feedthrough
rlabel pdiffusion 269 -1052 269 -1052 0 feedthrough
rlabel pdiffusion 276 -1052 276 -1052 0 feedthrough
rlabel pdiffusion 283 -1052 283 -1052 0 feedthrough
rlabel pdiffusion 290 -1052 290 -1052 0 cellNo=72
rlabel pdiffusion 297 -1052 297 -1052 0 feedthrough
rlabel pdiffusion 304 -1052 304 -1052 0 feedthrough
rlabel pdiffusion 311 -1052 311 -1052 0 feedthrough
rlabel pdiffusion 318 -1052 318 -1052 0 feedthrough
rlabel pdiffusion 325 -1052 325 -1052 0 feedthrough
rlabel pdiffusion 332 -1052 332 -1052 0 cellNo=532
rlabel pdiffusion 339 -1052 339 -1052 0 feedthrough
rlabel pdiffusion 346 -1052 346 -1052 0 feedthrough
rlabel pdiffusion 353 -1052 353 -1052 0 cellNo=533
rlabel pdiffusion 360 -1052 360 -1052 0 feedthrough
rlabel pdiffusion 367 -1052 367 -1052 0 feedthrough
rlabel pdiffusion 374 -1052 374 -1052 0 feedthrough
rlabel pdiffusion 381 -1052 381 -1052 0 feedthrough
rlabel pdiffusion 388 -1052 388 -1052 0 feedthrough
rlabel pdiffusion 395 -1052 395 -1052 0 feedthrough
rlabel pdiffusion 402 -1052 402 -1052 0 feedthrough
rlabel pdiffusion 409 -1052 409 -1052 0 feedthrough
rlabel pdiffusion 416 -1052 416 -1052 0 feedthrough
rlabel pdiffusion 423 -1052 423 -1052 0 cellNo=580
rlabel pdiffusion 430 -1052 430 -1052 0 cellNo=626
rlabel pdiffusion 444 -1052 444 -1052 0 cellNo=487
rlabel pdiffusion 451 -1052 451 -1052 0 cellNo=391
rlabel pdiffusion 458 -1052 458 -1052 0 feedthrough
rlabel pdiffusion 479 -1052 479 -1052 0 feedthrough
rlabel pdiffusion 514 -1052 514 -1052 0 cellNo=549
rlabel pdiffusion 521 -1052 521 -1052 0 cellNo=108
rlabel pdiffusion 528 -1052 528 -1052 0 feedthrough
rlabel pdiffusion 52 -1097 52 -1097 0 feedthrough
rlabel pdiffusion 59 -1097 59 -1097 0 cellNo=562
rlabel pdiffusion 66 -1097 66 -1097 0 feedthrough
rlabel pdiffusion 73 -1097 73 -1097 0 cellNo=670
rlabel pdiffusion 80 -1097 80 -1097 0 cellNo=139
rlabel pdiffusion 87 -1097 87 -1097 0 cellNo=292
rlabel pdiffusion 94 -1097 94 -1097 0 feedthrough
rlabel pdiffusion 101 -1097 101 -1097 0 feedthrough
rlabel pdiffusion 108 -1097 108 -1097 0 cellNo=633
rlabel pdiffusion 115 -1097 115 -1097 0 feedthrough
rlabel pdiffusion 122 -1097 122 -1097 0 feedthrough
rlabel pdiffusion 129 -1097 129 -1097 0 cellNo=91
rlabel pdiffusion 136 -1097 136 -1097 0 cellNo=539
rlabel pdiffusion 143 -1097 143 -1097 0 feedthrough
rlabel pdiffusion 150 -1097 150 -1097 0 feedthrough
rlabel pdiffusion 157 -1097 157 -1097 0 feedthrough
rlabel pdiffusion 164 -1097 164 -1097 0 feedthrough
rlabel pdiffusion 171 -1097 171 -1097 0 feedthrough
rlabel pdiffusion 178 -1097 178 -1097 0 cellNo=463
rlabel pdiffusion 185 -1097 185 -1097 0 cellNo=667
rlabel pdiffusion 192 -1097 192 -1097 0 cellNo=497
rlabel pdiffusion 199 -1097 199 -1097 0 feedthrough
rlabel pdiffusion 206 -1097 206 -1097 0 feedthrough
rlabel pdiffusion 213 -1097 213 -1097 0 feedthrough
rlabel pdiffusion 220 -1097 220 -1097 0 cellNo=462
rlabel pdiffusion 227 -1097 227 -1097 0 feedthrough
rlabel pdiffusion 234 -1097 234 -1097 0 cellNo=666
rlabel pdiffusion 241 -1097 241 -1097 0 feedthrough
rlabel pdiffusion 248 -1097 248 -1097 0 feedthrough
rlabel pdiffusion 255 -1097 255 -1097 0 feedthrough
rlabel pdiffusion 262 -1097 262 -1097 0 feedthrough
rlabel pdiffusion 269 -1097 269 -1097 0 feedthrough
rlabel pdiffusion 276 -1097 276 -1097 0 feedthrough
rlabel pdiffusion 283 -1097 283 -1097 0 feedthrough
rlabel pdiffusion 290 -1097 290 -1097 0 cellNo=57
rlabel pdiffusion 297 -1097 297 -1097 0 cellNo=250
rlabel pdiffusion 304 -1097 304 -1097 0 cellNo=161
rlabel pdiffusion 311 -1097 311 -1097 0 feedthrough
rlabel pdiffusion 318 -1097 318 -1097 0 cellNo=454
rlabel pdiffusion 325 -1097 325 -1097 0 feedthrough
rlabel pdiffusion 332 -1097 332 -1097 0 feedthrough
rlabel pdiffusion 339 -1097 339 -1097 0 feedthrough
rlabel pdiffusion 346 -1097 346 -1097 0 feedthrough
rlabel pdiffusion 353 -1097 353 -1097 0 feedthrough
rlabel pdiffusion 360 -1097 360 -1097 0 feedthrough
rlabel pdiffusion 367 -1097 367 -1097 0 feedthrough
rlabel pdiffusion 374 -1097 374 -1097 0 cellNo=596
rlabel pdiffusion 381 -1097 381 -1097 0 feedthrough
rlabel pdiffusion 388 -1097 388 -1097 0 cellNo=613
rlabel pdiffusion 395 -1097 395 -1097 0 feedthrough
rlabel pdiffusion 402 -1097 402 -1097 0 feedthrough
rlabel pdiffusion 409 -1097 409 -1097 0 feedthrough
rlabel pdiffusion 416 -1097 416 -1097 0 cellNo=572
rlabel pdiffusion 423 -1097 423 -1097 0 feedthrough
rlabel pdiffusion 430 -1097 430 -1097 0 feedthrough
rlabel pdiffusion 437 -1097 437 -1097 0 cellNo=183
rlabel pdiffusion 458 -1097 458 -1097 0 cellNo=715
rlabel pdiffusion 465 -1097 465 -1097 0 feedthrough
rlabel pdiffusion 479 -1097 479 -1097 0 feedthrough
rlabel pdiffusion 31 -1134 31 -1134 0 feedthrough
rlabel pdiffusion 38 -1134 38 -1134 0 feedthrough
rlabel pdiffusion 45 -1134 45 -1134 0 feedthrough
rlabel pdiffusion 52 -1134 52 -1134 0 cellNo=320
rlabel pdiffusion 59 -1134 59 -1134 0 feedthrough
rlabel pdiffusion 66 -1134 66 -1134 0 feedthrough
rlabel pdiffusion 73 -1134 73 -1134 0 cellNo=486
rlabel pdiffusion 80 -1134 80 -1134 0 cellNo=352
rlabel pdiffusion 87 -1134 87 -1134 0 cellNo=116
rlabel pdiffusion 94 -1134 94 -1134 0 cellNo=634
rlabel pdiffusion 101 -1134 101 -1134 0 feedthrough
rlabel pdiffusion 108 -1134 108 -1134 0 feedthrough
rlabel pdiffusion 115 -1134 115 -1134 0 cellNo=528
rlabel pdiffusion 122 -1134 122 -1134 0 feedthrough
rlabel pdiffusion 129 -1134 129 -1134 0 cellNo=518
rlabel pdiffusion 136 -1134 136 -1134 0 feedthrough
rlabel pdiffusion 143 -1134 143 -1134 0 feedthrough
rlabel pdiffusion 150 -1134 150 -1134 0 feedthrough
rlabel pdiffusion 157 -1134 157 -1134 0 cellNo=333
rlabel pdiffusion 164 -1134 164 -1134 0 feedthrough
rlabel pdiffusion 171 -1134 171 -1134 0 cellNo=118
rlabel pdiffusion 178 -1134 178 -1134 0 feedthrough
rlabel pdiffusion 185 -1134 185 -1134 0 feedthrough
rlabel pdiffusion 192 -1134 192 -1134 0 cellNo=662
rlabel pdiffusion 199 -1134 199 -1134 0 cellNo=11
rlabel pdiffusion 206 -1134 206 -1134 0 cellNo=448
rlabel pdiffusion 213 -1134 213 -1134 0 feedthrough
rlabel pdiffusion 220 -1134 220 -1134 0 feedthrough
rlabel pdiffusion 227 -1134 227 -1134 0 cellNo=653
rlabel pdiffusion 234 -1134 234 -1134 0 feedthrough
rlabel pdiffusion 241 -1134 241 -1134 0 feedthrough
rlabel pdiffusion 248 -1134 248 -1134 0 feedthrough
rlabel pdiffusion 255 -1134 255 -1134 0 cellNo=24
rlabel pdiffusion 262 -1134 262 -1134 0 cellNo=535
rlabel pdiffusion 269 -1134 269 -1134 0 feedthrough
rlabel pdiffusion 276 -1134 276 -1134 0 cellNo=248
rlabel pdiffusion 283 -1134 283 -1134 0 feedthrough
rlabel pdiffusion 290 -1134 290 -1134 0 feedthrough
rlabel pdiffusion 297 -1134 297 -1134 0 feedthrough
rlabel pdiffusion 304 -1134 304 -1134 0 cellNo=143
rlabel pdiffusion 311 -1134 311 -1134 0 feedthrough
rlabel pdiffusion 318 -1134 318 -1134 0 cellNo=718
rlabel pdiffusion 325 -1134 325 -1134 0 cellNo=304
rlabel pdiffusion 332 -1134 332 -1134 0 feedthrough
rlabel pdiffusion 339 -1134 339 -1134 0 feedthrough
rlabel pdiffusion 346 -1134 346 -1134 0 feedthrough
rlabel pdiffusion 353 -1134 353 -1134 0 feedthrough
rlabel pdiffusion 360 -1134 360 -1134 0 cellNo=356
rlabel pdiffusion 367 -1134 367 -1134 0 cellNo=69
rlabel pdiffusion 374 -1134 374 -1134 0 feedthrough
rlabel pdiffusion 381 -1134 381 -1134 0 feedthrough
rlabel pdiffusion 388 -1134 388 -1134 0 feedthrough
rlabel pdiffusion 395 -1134 395 -1134 0 feedthrough
rlabel pdiffusion 402 -1134 402 -1134 0 feedthrough
rlabel pdiffusion 409 -1134 409 -1134 0 feedthrough
rlabel pdiffusion 416 -1134 416 -1134 0 feedthrough
rlabel pdiffusion 423 -1134 423 -1134 0 feedthrough
rlabel pdiffusion 430 -1134 430 -1134 0 feedthrough
rlabel pdiffusion 437 -1134 437 -1134 0 feedthrough
rlabel pdiffusion 444 -1134 444 -1134 0 feedthrough
rlabel pdiffusion 479 -1134 479 -1134 0 feedthrough
rlabel pdiffusion 486 -1134 486 -1134 0 cellNo=460
rlabel pdiffusion 52 -1177 52 -1177 0 cellNo=521
rlabel pdiffusion 59 -1177 59 -1177 0 cellNo=117
rlabel pdiffusion 73 -1177 73 -1177 0 feedthrough
rlabel pdiffusion 80 -1177 80 -1177 0 cellNo=158
rlabel pdiffusion 87 -1177 87 -1177 0 feedthrough
rlabel pdiffusion 94 -1177 94 -1177 0 cellNo=584
rlabel pdiffusion 101 -1177 101 -1177 0 feedthrough
rlabel pdiffusion 108 -1177 108 -1177 0 feedthrough
rlabel pdiffusion 115 -1177 115 -1177 0 cellNo=556
rlabel pdiffusion 122 -1177 122 -1177 0 cellNo=224
rlabel pdiffusion 129 -1177 129 -1177 0 feedthrough
rlabel pdiffusion 136 -1177 136 -1177 0 feedthrough
rlabel pdiffusion 143 -1177 143 -1177 0 cellNo=2
rlabel pdiffusion 150 -1177 150 -1177 0 feedthrough
rlabel pdiffusion 157 -1177 157 -1177 0 feedthrough
rlabel pdiffusion 164 -1177 164 -1177 0 cellNo=712
rlabel pdiffusion 171 -1177 171 -1177 0 cellNo=679
rlabel pdiffusion 178 -1177 178 -1177 0 feedthrough
rlabel pdiffusion 185 -1177 185 -1177 0 feedthrough
rlabel pdiffusion 192 -1177 192 -1177 0 feedthrough
rlabel pdiffusion 199 -1177 199 -1177 0 cellNo=209
rlabel pdiffusion 206 -1177 206 -1177 0 cellNo=659
rlabel pdiffusion 213 -1177 213 -1177 0 feedthrough
rlabel pdiffusion 220 -1177 220 -1177 0 feedthrough
rlabel pdiffusion 227 -1177 227 -1177 0 feedthrough
rlabel pdiffusion 234 -1177 234 -1177 0 feedthrough
rlabel pdiffusion 241 -1177 241 -1177 0 cellNo=654
rlabel pdiffusion 248 -1177 248 -1177 0 cellNo=675
rlabel pdiffusion 255 -1177 255 -1177 0 cellNo=500
rlabel pdiffusion 262 -1177 262 -1177 0 cellNo=71
rlabel pdiffusion 269 -1177 269 -1177 0 feedthrough
rlabel pdiffusion 276 -1177 276 -1177 0 feedthrough
rlabel pdiffusion 283 -1177 283 -1177 0 feedthrough
rlabel pdiffusion 290 -1177 290 -1177 0 feedthrough
rlabel pdiffusion 297 -1177 297 -1177 0 cellNo=357
rlabel pdiffusion 304 -1177 304 -1177 0 cellNo=422
rlabel pdiffusion 311 -1177 311 -1177 0 feedthrough
rlabel pdiffusion 318 -1177 318 -1177 0 feedthrough
rlabel pdiffusion 325 -1177 325 -1177 0 feedthrough
rlabel pdiffusion 332 -1177 332 -1177 0 feedthrough
rlabel pdiffusion 339 -1177 339 -1177 0 feedthrough
rlabel pdiffusion 346 -1177 346 -1177 0 feedthrough
rlabel pdiffusion 353 -1177 353 -1177 0 feedthrough
rlabel pdiffusion 360 -1177 360 -1177 0 feedthrough
rlabel pdiffusion 367 -1177 367 -1177 0 feedthrough
rlabel pdiffusion 374 -1177 374 -1177 0 cellNo=661
rlabel pdiffusion 381 -1177 381 -1177 0 feedthrough
rlabel pdiffusion 388 -1177 388 -1177 0 feedthrough
rlabel pdiffusion 395 -1177 395 -1177 0 cellNo=525
rlabel pdiffusion 402 -1177 402 -1177 0 feedthrough
rlabel pdiffusion 409 -1177 409 -1177 0 cellNo=574
rlabel pdiffusion 66 -1208 66 -1208 0 feedthrough
rlabel pdiffusion 73 -1208 73 -1208 0 feedthrough
rlabel pdiffusion 80 -1208 80 -1208 0 feedthrough
rlabel pdiffusion 87 -1208 87 -1208 0 cellNo=257
rlabel pdiffusion 94 -1208 94 -1208 0 feedthrough
rlabel pdiffusion 101 -1208 101 -1208 0 feedthrough
rlabel pdiffusion 108 -1208 108 -1208 0 cellNo=704
rlabel pdiffusion 115 -1208 115 -1208 0 feedthrough
rlabel pdiffusion 122 -1208 122 -1208 0 feedthrough
rlabel pdiffusion 129 -1208 129 -1208 0 cellNo=60
rlabel pdiffusion 136 -1208 136 -1208 0 cellNo=54
rlabel pdiffusion 143 -1208 143 -1208 0 feedthrough
rlabel pdiffusion 150 -1208 150 -1208 0 cellNo=615
rlabel pdiffusion 157 -1208 157 -1208 0 cellNo=225
rlabel pdiffusion 164 -1208 164 -1208 0 feedthrough
rlabel pdiffusion 171 -1208 171 -1208 0 cellNo=652
rlabel pdiffusion 178 -1208 178 -1208 0 cellNo=106
rlabel pdiffusion 185 -1208 185 -1208 0 cellNo=698
rlabel pdiffusion 192 -1208 192 -1208 0 cellNo=301
rlabel pdiffusion 199 -1208 199 -1208 0 feedthrough
rlabel pdiffusion 206 -1208 206 -1208 0 cellNo=637
rlabel pdiffusion 213 -1208 213 -1208 0 feedthrough
rlabel pdiffusion 220 -1208 220 -1208 0 feedthrough
rlabel pdiffusion 227 -1208 227 -1208 0 cellNo=210
rlabel pdiffusion 234 -1208 234 -1208 0 feedthrough
rlabel pdiffusion 241 -1208 241 -1208 0 cellNo=567
rlabel pdiffusion 248 -1208 248 -1208 0 feedthrough
rlabel pdiffusion 255 -1208 255 -1208 0 feedthrough
rlabel pdiffusion 262 -1208 262 -1208 0 cellNo=678
rlabel pdiffusion 269 -1208 269 -1208 0 feedthrough
rlabel pdiffusion 276 -1208 276 -1208 0 feedthrough
rlabel pdiffusion 283 -1208 283 -1208 0 feedthrough
rlabel pdiffusion 290 -1208 290 -1208 0 cellNo=196
rlabel pdiffusion 297 -1208 297 -1208 0 feedthrough
rlabel pdiffusion 304 -1208 304 -1208 0 cellNo=215
rlabel pdiffusion 311 -1208 311 -1208 0 feedthrough
rlabel pdiffusion 318 -1208 318 -1208 0 cellNo=344
rlabel pdiffusion 325 -1208 325 -1208 0 cellNo=688
rlabel pdiffusion 332 -1208 332 -1208 0 feedthrough
rlabel pdiffusion 339 -1208 339 -1208 0 feedthrough
rlabel pdiffusion 346 -1208 346 -1208 0 feedthrough
rlabel pdiffusion 353 -1208 353 -1208 0 feedthrough
rlabel pdiffusion 360 -1208 360 -1208 0 feedthrough
rlabel pdiffusion 367 -1208 367 -1208 0 feedthrough
rlabel pdiffusion 374 -1208 374 -1208 0 feedthrough
rlabel pdiffusion 381 -1208 381 -1208 0 cellNo=571
rlabel pdiffusion 388 -1208 388 -1208 0 feedthrough
rlabel pdiffusion 395 -1208 395 -1208 0 feedthrough
rlabel pdiffusion 94 -1237 94 -1237 0 feedthrough
rlabel pdiffusion 101 -1237 101 -1237 0 cellNo=370
rlabel pdiffusion 108 -1237 108 -1237 0 cellNo=204
rlabel pdiffusion 115 -1237 115 -1237 0 feedthrough
rlabel pdiffusion 122 -1237 122 -1237 0 cellNo=283
rlabel pdiffusion 129 -1237 129 -1237 0 feedthrough
rlabel pdiffusion 136 -1237 136 -1237 0 feedthrough
rlabel pdiffusion 143 -1237 143 -1237 0 feedthrough
rlabel pdiffusion 150 -1237 150 -1237 0 cellNo=561
rlabel pdiffusion 157 -1237 157 -1237 0 feedthrough
rlabel pdiffusion 164 -1237 164 -1237 0 feedthrough
rlabel pdiffusion 171 -1237 171 -1237 0 cellNo=587
rlabel pdiffusion 178 -1237 178 -1237 0 cellNo=491
rlabel pdiffusion 185 -1237 185 -1237 0 cellNo=205
rlabel pdiffusion 192 -1237 192 -1237 0 cellNo=87
rlabel pdiffusion 199 -1237 199 -1237 0 cellNo=362
rlabel pdiffusion 206 -1237 206 -1237 0 feedthrough
rlabel pdiffusion 213 -1237 213 -1237 0 feedthrough
rlabel pdiffusion 220 -1237 220 -1237 0 cellNo=409
rlabel pdiffusion 227 -1237 227 -1237 0 feedthrough
rlabel pdiffusion 234 -1237 234 -1237 0 feedthrough
rlabel pdiffusion 241 -1237 241 -1237 0 feedthrough
rlabel pdiffusion 248 -1237 248 -1237 0 feedthrough
rlabel pdiffusion 255 -1237 255 -1237 0 cellNo=222
rlabel pdiffusion 262 -1237 262 -1237 0 cellNo=184
rlabel pdiffusion 269 -1237 269 -1237 0 cellNo=239
rlabel pdiffusion 276 -1237 276 -1237 0 feedthrough
rlabel pdiffusion 283 -1237 283 -1237 0 feedthrough
rlabel pdiffusion 290 -1237 290 -1237 0 feedthrough
rlabel pdiffusion 297 -1237 297 -1237 0 cellNo=687
rlabel pdiffusion 304 -1237 304 -1237 0 cellNo=611
rlabel pdiffusion 311 -1237 311 -1237 0 feedthrough
rlabel pdiffusion 318 -1237 318 -1237 0 feedthrough
rlabel pdiffusion 325 -1237 325 -1237 0 feedthrough
rlabel pdiffusion 332 -1237 332 -1237 0 feedthrough
rlabel pdiffusion 346 -1237 346 -1237 0 cellNo=568
rlabel pdiffusion 353 -1237 353 -1237 0 feedthrough
rlabel pdiffusion 381 -1237 381 -1237 0 feedthrough
rlabel pdiffusion 3 -1258 3 -1258 0 cellNo=550
rlabel pdiffusion 73 -1258 73 -1258 0 cellNo=452
rlabel pdiffusion 80 -1258 80 -1258 0 cellNo=50
rlabel pdiffusion 87 -1258 87 -1258 0 feedthrough
rlabel pdiffusion 101 -1258 101 -1258 0 feedthrough
rlabel pdiffusion 108 -1258 108 -1258 0 feedthrough
rlabel pdiffusion 115 -1258 115 -1258 0 cellNo=23
rlabel pdiffusion 122 -1258 122 -1258 0 cellNo=314
rlabel pdiffusion 129 -1258 129 -1258 0 cellNo=112
rlabel pdiffusion 136 -1258 136 -1258 0 feedthrough
rlabel pdiffusion 143 -1258 143 -1258 0 cellNo=581
rlabel pdiffusion 150 -1258 150 -1258 0 cellNo=282
rlabel pdiffusion 157 -1258 157 -1258 0 cellNo=405
rlabel pdiffusion 164 -1258 164 -1258 0 cellNo=346
rlabel pdiffusion 171 -1258 171 -1258 0 cellNo=624
rlabel pdiffusion 178 -1258 178 -1258 0 feedthrough
rlabel pdiffusion 185 -1258 185 -1258 0 cellNo=566
rlabel pdiffusion 192 -1258 192 -1258 0 feedthrough
rlabel pdiffusion 199 -1258 199 -1258 0 cellNo=169
rlabel pdiffusion 206 -1258 206 -1258 0 feedthrough
rlabel pdiffusion 213 -1258 213 -1258 0 cellNo=683
rlabel pdiffusion 220 -1258 220 -1258 0 feedthrough
rlabel pdiffusion 227 -1258 227 -1258 0 cellNo=208
rlabel pdiffusion 234 -1258 234 -1258 0 feedthrough
rlabel pdiffusion 241 -1258 241 -1258 0 feedthrough
rlabel pdiffusion 248 -1258 248 -1258 0 cellNo=213
rlabel pdiffusion 255 -1258 255 -1258 0 feedthrough
rlabel pdiffusion 262 -1258 262 -1258 0 feedthrough
rlabel pdiffusion 269 -1258 269 -1258 0 feedthrough
rlabel pdiffusion 276 -1258 276 -1258 0 cellNo=569
rlabel pdiffusion 283 -1258 283 -1258 0 cellNo=37
rlabel pdiffusion 290 -1258 290 -1258 0 cellNo=299
rlabel pdiffusion 297 -1258 297 -1258 0 feedthrough
rlabel pdiffusion 304 -1258 304 -1258 0 feedthrough
rlabel pdiffusion 318 -1258 318 -1258 0 cellNo=366
rlabel pdiffusion 325 -1258 325 -1258 0 feedthrough
rlabel pdiffusion 381 -1258 381 -1258 0 feedthrough
rlabel pdiffusion 3 -1273 3 -1273 0 cellNo=517
rlabel pdiffusion 87 -1273 87 -1273 0 cellNo=322
rlabel pdiffusion 94 -1273 94 -1273 0 cellNo=513
rlabel pdiffusion 108 -1273 108 -1273 0 feedthrough
rlabel pdiffusion 115 -1273 115 -1273 0 cellNo=488
rlabel pdiffusion 122 -1273 122 -1273 0 feedthrough
rlabel pdiffusion 129 -1273 129 -1273 0 cellNo=530
rlabel pdiffusion 136 -1273 136 -1273 0 feedthrough
rlabel pdiffusion 143 -1273 143 -1273 0 cellNo=636
rlabel pdiffusion 150 -1273 150 -1273 0 feedthrough
rlabel pdiffusion 157 -1273 157 -1273 0 cellNo=522
rlabel pdiffusion 164 -1273 164 -1273 0 cellNo=404
rlabel pdiffusion 171 -1273 171 -1273 0 cellNo=134
rlabel pdiffusion 185 -1273 185 -1273 0 cellNo=70
rlabel pdiffusion 206 -1273 206 -1273 0 cellNo=330
rlabel pdiffusion 213 -1273 213 -1273 0 cellNo=655
rlabel pdiffusion 220 -1273 220 -1273 0 cellNo=445
rlabel pdiffusion 227 -1273 227 -1273 0 feedthrough
rlabel pdiffusion 234 -1273 234 -1273 0 cellNo=559
rlabel pdiffusion 241 -1273 241 -1273 0 cellNo=507
rlabel pdiffusion 269 -1273 269 -1273 0 cellNo=429
rlabel pdiffusion 276 -1273 276 -1273 0 feedthrough
rlabel pdiffusion 283 -1273 283 -1273 0 cellNo=565
rlabel pdiffusion 297 -1273 297 -1273 0 cellNo=618
rlabel pdiffusion 304 -1273 304 -1273 0 feedthrough
rlabel pdiffusion 381 -1273 381 -1273 0 cellNo=17
rlabel pdiffusion 388 -1273 388 -1273 0 feedthrough
rlabel polysilicon 135 -2 135 -2 0 1
rlabel polysilicon 135 -8 135 -8 0 3
rlabel polysilicon 142 -2 142 -2 0 1
rlabel polysilicon 145 -2 145 -2 0 2
rlabel polysilicon 142 -8 142 -8 0 3
rlabel polysilicon 149 -8 149 -8 0 3
rlabel polysilicon 152 -8 152 -8 0 4
rlabel polysilicon 156 -2 156 -2 0 1
rlabel polysilicon 184 -2 184 -2 0 1
rlabel polysilicon 184 -8 184 -8 0 3
rlabel polysilicon 194 -2 194 -2 0 2
rlabel polysilicon 212 -2 212 -2 0 1
rlabel polysilicon 212 -8 212 -8 0 3
rlabel polysilicon 219 -2 219 -2 0 1
rlabel polysilicon 254 -8 254 -8 0 3
rlabel polysilicon 257 -8 257 -8 0 4
rlabel polysilicon 142 -17 142 -17 0 1
rlabel polysilicon 149 -17 149 -17 0 1
rlabel polysilicon 149 -23 149 -23 0 3
rlabel polysilicon 156 -17 156 -17 0 1
rlabel polysilicon 156 -23 156 -23 0 3
rlabel polysilicon 163 -23 163 -23 0 3
rlabel polysilicon 166 -23 166 -23 0 4
rlabel polysilicon 173 -23 173 -23 0 4
rlabel polysilicon 177 -17 177 -17 0 1
rlabel polysilicon 180 -17 180 -17 0 2
rlabel polysilicon 177 -23 177 -23 0 3
rlabel polysilicon 184 -17 184 -17 0 1
rlabel polysilicon 184 -23 184 -23 0 3
rlabel polysilicon 191 -17 191 -17 0 1
rlabel polysilicon 198 -17 198 -17 0 1
rlabel polysilicon 198 -23 198 -23 0 3
rlabel polysilicon 205 -17 205 -17 0 1
rlabel polysilicon 208 -17 208 -17 0 2
rlabel polysilicon 205 -23 205 -23 0 3
rlabel polysilicon 212 -17 212 -17 0 1
rlabel polysilicon 212 -23 212 -23 0 3
rlabel polysilicon 222 -17 222 -17 0 2
rlabel polysilicon 243 -23 243 -23 0 4
rlabel polysilicon 254 -17 254 -17 0 1
rlabel polysilicon 254 -23 254 -23 0 3
rlabel polysilicon 261 -17 261 -17 0 1
rlabel polysilicon 268 -23 268 -23 0 3
rlabel polysilicon 310 -23 310 -23 0 3
rlabel polysilicon 54 -42 54 -42 0 4
rlabel polysilicon 100 -42 100 -42 0 3
rlabel polysilicon 145 -36 145 -36 0 2
rlabel polysilicon 149 -36 149 -36 0 1
rlabel polysilicon 149 -42 149 -42 0 3
rlabel polysilicon 163 -36 163 -36 0 1
rlabel polysilicon 163 -42 163 -42 0 3
rlabel polysilicon 170 -36 170 -36 0 1
rlabel polysilicon 177 -42 177 -42 0 3
rlabel polysilicon 187 -36 187 -36 0 2
rlabel polysilicon 187 -42 187 -42 0 4
rlabel polysilicon 191 -36 191 -36 0 1
rlabel polysilicon 191 -42 191 -42 0 3
rlabel polysilicon 201 -36 201 -36 0 2
rlabel polysilicon 198 -42 198 -42 0 3
rlabel polysilicon 208 -36 208 -36 0 2
rlabel polysilicon 208 -42 208 -42 0 4
rlabel polysilicon 212 -36 212 -36 0 1
rlabel polysilicon 212 -42 212 -42 0 3
rlabel polysilicon 219 -36 219 -36 0 1
rlabel polysilicon 219 -42 219 -42 0 3
rlabel polysilicon 229 -36 229 -36 0 2
rlabel polysilicon 233 -36 233 -36 0 1
rlabel polysilicon 233 -42 233 -42 0 3
rlabel polysilicon 236 -42 236 -42 0 4
rlabel polysilicon 240 -36 240 -36 0 1
rlabel polysilicon 240 -42 240 -42 0 3
rlabel polysilicon 247 -36 247 -36 0 1
rlabel polysilicon 247 -42 247 -42 0 3
rlabel polysilicon 254 -36 254 -36 0 1
rlabel polysilicon 254 -42 254 -42 0 3
rlabel polysilicon 261 -36 261 -36 0 1
rlabel polysilicon 261 -42 261 -42 0 3
rlabel polysilicon 271 -36 271 -36 0 2
rlabel polysilicon 268 -42 268 -42 0 3
rlabel polysilicon 310 -36 310 -36 0 1
rlabel polysilicon 310 -42 310 -42 0 3
rlabel polysilicon 341 -36 341 -36 0 2
rlabel polysilicon 338 -42 338 -42 0 3
rlabel polysilicon 345 -36 345 -36 0 1
rlabel polysilicon 345 -42 345 -42 0 3
rlabel polysilicon 359 -42 359 -42 0 3
rlabel polysilicon 362 -42 362 -42 0 4
rlabel polysilicon 26 -65 26 -65 0 4
rlabel polysilicon 51 -59 51 -59 0 1
rlabel polysilicon 72 -59 72 -59 0 1
rlabel polysilicon 72 -65 72 -65 0 3
rlabel polysilicon 96 -59 96 -59 0 2
rlabel polysilicon 93 -65 93 -65 0 3
rlabel polysilicon 96 -65 96 -65 0 4
rlabel polysilicon 100 -59 100 -59 0 1
rlabel polysilicon 100 -65 100 -65 0 3
rlabel polysilicon 138 -59 138 -59 0 2
rlabel polysilicon 142 -59 142 -59 0 1
rlabel polysilicon 142 -65 142 -65 0 3
rlabel polysilicon 149 -65 149 -65 0 3
rlabel polysilicon 156 -59 156 -59 0 1
rlabel polysilicon 163 -59 163 -59 0 1
rlabel polysilicon 163 -65 163 -65 0 3
rlabel polysilicon 170 -59 170 -59 0 1
rlabel polysilicon 170 -65 170 -65 0 3
rlabel polysilicon 177 -59 177 -59 0 1
rlabel polysilicon 187 -59 187 -59 0 2
rlabel polysilicon 187 -65 187 -65 0 4
rlabel polysilicon 191 -59 191 -59 0 1
rlabel polysilicon 194 -59 194 -59 0 2
rlabel polysilicon 198 -59 198 -59 0 1
rlabel polysilicon 201 -59 201 -59 0 2
rlabel polysilicon 201 -65 201 -65 0 4
rlabel polysilicon 205 -59 205 -59 0 1
rlabel polysilicon 205 -65 205 -65 0 3
rlabel polysilicon 212 -59 212 -59 0 1
rlabel polysilicon 212 -65 212 -65 0 3
rlabel polysilicon 219 -59 219 -59 0 1
rlabel polysilicon 219 -65 219 -65 0 3
rlabel polysilicon 226 -59 226 -59 0 1
rlabel polysilicon 226 -65 226 -65 0 3
rlabel polysilicon 229 -65 229 -65 0 4
rlabel polysilicon 233 -59 233 -59 0 1
rlabel polysilicon 233 -65 233 -65 0 3
rlabel polysilicon 240 -59 240 -59 0 1
rlabel polysilicon 243 -59 243 -59 0 2
rlabel polysilicon 240 -65 240 -65 0 3
rlabel polysilicon 247 -59 247 -59 0 1
rlabel polysilicon 247 -65 247 -65 0 3
rlabel polysilicon 254 -59 254 -59 0 1
rlabel polysilicon 254 -65 254 -65 0 3
rlabel polysilicon 261 -59 261 -59 0 1
rlabel polysilicon 261 -65 261 -65 0 3
rlabel polysilicon 268 -59 268 -59 0 1
rlabel polysilicon 268 -65 268 -65 0 3
rlabel polysilicon 275 -59 275 -59 0 1
rlabel polysilicon 278 -65 278 -65 0 4
rlabel polysilicon 282 -59 282 -59 0 1
rlabel polysilicon 282 -65 282 -65 0 3
rlabel polysilicon 289 -59 289 -59 0 1
rlabel polysilicon 289 -65 289 -65 0 3
rlabel polysilicon 296 -59 296 -59 0 1
rlabel polysilicon 296 -65 296 -65 0 3
rlabel polysilicon 310 -59 310 -59 0 1
rlabel polysilicon 310 -65 310 -65 0 3
rlabel polysilicon 317 -65 317 -65 0 3
rlabel polysilicon 320 -65 320 -65 0 4
rlabel polysilicon 338 -59 338 -59 0 1
rlabel polysilicon 338 -65 338 -65 0 3
rlabel polysilicon 345 -59 345 -59 0 1
rlabel polysilicon 348 -65 348 -65 0 4
rlabel polysilicon 352 -59 352 -59 0 1
rlabel polysilicon 352 -65 352 -65 0 3
rlabel polysilicon 366 -59 366 -59 0 1
rlabel polysilicon 366 -65 366 -65 0 3
rlabel polysilicon 26 -90 26 -90 0 2
rlabel polysilicon 51 -90 51 -90 0 1
rlabel polysilicon 58 -90 58 -90 0 1
rlabel polysilicon 58 -96 58 -96 0 3
rlabel polysilicon 65 -90 65 -90 0 1
rlabel polysilicon 65 -96 65 -96 0 3
rlabel polysilicon 72 -90 72 -90 0 1
rlabel polysilicon 72 -96 72 -96 0 3
rlabel polysilicon 79 -90 79 -90 0 1
rlabel polysilicon 79 -96 79 -96 0 3
rlabel polysilicon 86 -90 86 -90 0 1
rlabel polysilicon 93 -90 93 -90 0 1
rlabel polysilicon 93 -96 93 -96 0 3
rlabel polysilicon 103 -90 103 -90 0 2
rlabel polysilicon 103 -96 103 -96 0 4
rlabel polysilicon 107 -90 107 -90 0 1
rlabel polysilicon 107 -96 107 -96 0 3
rlabel polysilicon 114 -90 114 -90 0 1
rlabel polysilicon 114 -96 114 -96 0 3
rlabel polysilicon 121 -90 121 -90 0 1
rlabel polysilicon 121 -96 121 -96 0 3
rlabel polysilicon 128 -90 128 -90 0 1
rlabel polysilicon 128 -96 128 -96 0 3
rlabel polysilicon 135 -90 135 -90 0 1
rlabel polysilicon 138 -90 138 -90 0 2
rlabel polysilicon 145 -90 145 -90 0 2
rlabel polysilicon 142 -96 142 -96 0 3
rlabel polysilicon 145 -96 145 -96 0 4
rlabel polysilicon 149 -90 149 -90 0 1
rlabel polysilicon 149 -96 149 -96 0 3
rlabel polysilicon 156 -90 156 -90 0 1
rlabel polysilicon 156 -96 156 -96 0 3
rlabel polysilicon 163 -90 163 -90 0 1
rlabel polysilicon 163 -96 163 -96 0 3
rlabel polysilicon 170 -96 170 -96 0 3
rlabel polysilicon 173 -96 173 -96 0 4
rlabel polysilicon 177 -96 177 -96 0 3
rlabel polysilicon 180 -96 180 -96 0 4
rlabel polysilicon 187 -90 187 -90 0 2
rlabel polysilicon 187 -96 187 -96 0 4
rlabel polysilicon 191 -90 191 -90 0 1
rlabel polysilicon 194 -90 194 -90 0 2
rlabel polysilicon 191 -96 191 -96 0 3
rlabel polysilicon 194 -96 194 -96 0 4
rlabel polysilicon 198 -90 198 -90 0 1
rlabel polysilicon 201 -96 201 -96 0 4
rlabel polysilicon 205 -90 205 -90 0 1
rlabel polysilicon 208 -90 208 -90 0 2
rlabel polysilicon 205 -96 205 -96 0 3
rlabel polysilicon 208 -96 208 -96 0 4
rlabel polysilicon 212 -90 212 -90 0 1
rlabel polysilicon 212 -96 212 -96 0 3
rlabel polysilicon 219 -90 219 -90 0 1
rlabel polysilicon 219 -96 219 -96 0 3
rlabel polysilicon 226 -90 226 -90 0 1
rlabel polysilicon 226 -96 226 -96 0 3
rlabel polysilicon 236 -90 236 -90 0 2
rlabel polysilicon 236 -96 236 -96 0 4
rlabel polysilicon 243 -90 243 -90 0 2
rlabel polysilicon 240 -96 240 -96 0 3
rlabel polysilicon 243 -96 243 -96 0 4
rlabel polysilicon 250 -90 250 -90 0 2
rlabel polysilicon 247 -96 247 -96 0 3
rlabel polysilicon 250 -96 250 -96 0 4
rlabel polysilicon 254 -90 254 -90 0 1
rlabel polysilicon 257 -90 257 -90 0 2
rlabel polysilicon 254 -96 254 -96 0 3
rlabel polysilicon 257 -96 257 -96 0 4
rlabel polysilicon 261 -90 261 -90 0 1
rlabel polysilicon 261 -96 261 -96 0 3
rlabel polysilicon 268 -90 268 -90 0 1
rlabel polysilicon 268 -96 268 -96 0 3
rlabel polysilicon 275 -90 275 -90 0 1
rlabel polysilicon 275 -96 275 -96 0 3
rlabel polysilicon 282 -90 282 -90 0 1
rlabel polysilicon 282 -96 282 -96 0 3
rlabel polysilicon 289 -90 289 -90 0 1
rlabel polysilicon 289 -96 289 -96 0 3
rlabel polysilicon 296 -90 296 -90 0 1
rlabel polysilicon 296 -96 296 -96 0 3
rlabel polysilicon 303 -90 303 -90 0 1
rlabel polysilicon 303 -96 303 -96 0 3
rlabel polysilicon 310 -90 310 -90 0 1
rlabel polysilicon 310 -96 310 -96 0 3
rlabel polysilicon 317 -90 317 -90 0 1
rlabel polysilicon 317 -96 317 -96 0 3
rlabel polysilicon 324 -90 324 -90 0 1
rlabel polysilicon 324 -96 324 -96 0 3
rlabel polysilicon 331 -90 331 -90 0 1
rlabel polysilicon 331 -96 331 -96 0 3
rlabel polysilicon 338 -90 338 -90 0 1
rlabel polysilicon 338 -96 338 -96 0 3
rlabel polysilicon 345 -90 345 -90 0 1
rlabel polysilicon 345 -96 345 -96 0 3
rlabel polysilicon 352 -90 352 -90 0 1
rlabel polysilicon 352 -96 352 -96 0 3
rlabel polysilicon 366 -90 366 -90 0 1
rlabel polysilicon 366 -96 366 -96 0 3
rlabel polysilicon 376 -90 376 -90 0 2
rlabel polysilicon 373 -96 373 -96 0 3
rlabel polysilicon 376 -96 376 -96 0 4
rlabel polysilicon 86 -133 86 -133 0 1
rlabel polysilicon 86 -139 86 -139 0 3
rlabel polysilicon 93 -133 93 -133 0 1
rlabel polysilicon 93 -139 93 -139 0 3
rlabel polysilicon 100 -133 100 -133 0 1
rlabel polysilicon 100 -139 100 -139 0 3
rlabel polysilicon 107 -133 107 -133 0 1
rlabel polysilicon 107 -139 107 -139 0 3
rlabel polysilicon 117 -139 117 -139 0 4
rlabel polysilicon 121 -133 121 -133 0 1
rlabel polysilicon 124 -139 124 -139 0 4
rlabel polysilicon 128 -133 128 -133 0 1
rlabel polysilicon 128 -139 128 -139 0 3
rlabel polysilicon 135 -133 135 -133 0 1
rlabel polysilicon 135 -139 135 -139 0 3
rlabel polysilicon 142 -133 142 -133 0 1
rlabel polysilicon 145 -133 145 -133 0 2
rlabel polysilicon 142 -139 142 -139 0 3
rlabel polysilicon 149 -133 149 -133 0 1
rlabel polysilicon 149 -139 149 -139 0 3
rlabel polysilicon 156 -133 156 -133 0 1
rlabel polysilicon 163 -133 163 -133 0 1
rlabel polysilicon 163 -139 163 -139 0 3
rlabel polysilicon 170 -133 170 -133 0 1
rlabel polysilicon 170 -139 170 -139 0 3
rlabel polysilicon 173 -139 173 -139 0 4
rlabel polysilicon 180 -133 180 -133 0 2
rlabel polysilicon 184 -133 184 -133 0 1
rlabel polysilicon 184 -139 184 -139 0 3
rlabel polysilicon 191 -133 191 -133 0 1
rlabel polysilicon 194 -133 194 -133 0 2
rlabel polysilicon 198 -133 198 -133 0 1
rlabel polysilicon 198 -139 198 -139 0 3
rlabel polysilicon 205 -133 205 -133 0 1
rlabel polysilicon 208 -133 208 -133 0 2
rlabel polysilicon 205 -139 205 -139 0 3
rlabel polysilicon 212 -133 212 -133 0 1
rlabel polysilicon 212 -139 212 -139 0 3
rlabel polysilicon 219 -133 219 -133 0 1
rlabel polysilicon 219 -139 219 -139 0 3
rlabel polysilicon 226 -133 226 -133 0 1
rlabel polysilicon 229 -139 229 -139 0 4
rlabel polysilicon 236 -133 236 -133 0 2
rlabel polysilicon 236 -139 236 -139 0 4
rlabel polysilicon 240 -133 240 -133 0 1
rlabel polysilicon 240 -139 240 -139 0 3
rlabel polysilicon 250 -133 250 -133 0 2
rlabel polysilicon 247 -139 247 -139 0 3
rlabel polysilicon 254 -133 254 -133 0 1
rlabel polysilicon 254 -139 254 -139 0 3
rlabel polysilicon 261 -133 261 -133 0 1
rlabel polysilicon 264 -133 264 -133 0 2
rlabel polysilicon 264 -139 264 -139 0 4
rlabel polysilicon 271 -133 271 -133 0 2
rlabel polysilicon 275 -133 275 -133 0 1
rlabel polysilicon 275 -139 275 -139 0 3
rlabel polysilicon 282 -139 282 -139 0 3
rlabel polysilicon 289 -133 289 -133 0 1
rlabel polysilicon 289 -139 289 -139 0 3
rlabel polysilicon 296 -133 296 -133 0 1
rlabel polysilicon 296 -139 296 -139 0 3
rlabel polysilicon 303 -133 303 -133 0 1
rlabel polysilicon 303 -139 303 -139 0 3
rlabel polysilicon 310 -133 310 -133 0 1
rlabel polysilicon 310 -139 310 -139 0 3
rlabel polysilicon 317 -133 317 -133 0 1
rlabel polysilicon 317 -139 317 -139 0 3
rlabel polysilicon 324 -133 324 -133 0 1
rlabel polysilicon 324 -139 324 -139 0 3
rlabel polysilicon 331 -133 331 -133 0 1
rlabel polysilicon 331 -139 331 -139 0 3
rlabel polysilicon 338 -133 338 -133 0 1
rlabel polysilicon 341 -139 341 -139 0 4
rlabel polysilicon 345 -133 345 -133 0 1
rlabel polysilicon 345 -139 345 -139 0 3
rlabel polysilicon 355 -139 355 -139 0 4
rlabel polysilicon 366 -133 366 -133 0 1
rlabel polysilicon 366 -139 366 -139 0 3
rlabel polysilicon 380 -133 380 -133 0 1
rlabel polysilicon 380 -139 380 -139 0 3
rlabel polysilicon 394 -133 394 -133 0 1
rlabel polysilicon 394 -139 394 -139 0 3
rlabel polysilicon 401 -133 401 -133 0 1
rlabel polysilicon 401 -139 401 -139 0 3
rlabel polysilicon 65 -168 65 -168 0 1
rlabel polysilicon 65 -174 65 -174 0 3
rlabel polysilicon 72 -168 72 -168 0 1
rlabel polysilicon 72 -174 72 -174 0 3
rlabel polysilicon 79 -174 79 -174 0 3
rlabel polysilicon 82 -174 82 -174 0 4
rlabel polysilicon 86 -168 86 -168 0 1
rlabel polysilicon 86 -174 86 -174 0 3
rlabel polysilicon 93 -168 93 -168 0 1
rlabel polysilicon 93 -174 93 -174 0 3
rlabel polysilicon 100 -168 100 -168 0 1
rlabel polysilicon 100 -174 100 -174 0 3
rlabel polysilicon 107 -168 107 -168 0 1
rlabel polysilicon 107 -174 107 -174 0 3
rlabel polysilicon 117 -168 117 -168 0 2
rlabel polysilicon 114 -174 114 -174 0 3
rlabel polysilicon 121 -168 121 -168 0 1
rlabel polysilicon 121 -174 121 -174 0 3
rlabel polysilicon 128 -168 128 -168 0 1
rlabel polysilicon 131 -174 131 -174 0 4
rlabel polysilicon 135 -168 135 -168 0 1
rlabel polysilicon 135 -174 135 -174 0 3
rlabel polysilicon 138 -174 138 -174 0 4
rlabel polysilicon 142 -168 142 -168 0 1
rlabel polysilicon 142 -174 142 -174 0 3
rlabel polysilicon 145 -174 145 -174 0 4
rlabel polysilicon 149 -168 149 -168 0 1
rlabel polysilicon 152 -168 152 -168 0 2
rlabel polysilicon 156 -168 156 -168 0 1
rlabel polysilicon 156 -174 156 -174 0 3
rlabel polysilicon 163 -168 163 -168 0 1
rlabel polysilicon 163 -174 163 -174 0 3
rlabel polysilicon 170 -168 170 -168 0 1
rlabel polysilicon 170 -174 170 -174 0 3
rlabel polysilicon 177 -168 177 -168 0 1
rlabel polysilicon 180 -174 180 -174 0 4
rlabel polysilicon 184 -168 184 -168 0 1
rlabel polysilicon 184 -174 184 -174 0 3
rlabel polysilicon 191 -168 191 -168 0 1
rlabel polysilicon 191 -174 191 -174 0 3
rlabel polysilicon 198 -168 198 -168 0 1
rlabel polysilicon 198 -174 198 -174 0 3
rlabel polysilicon 201 -174 201 -174 0 4
rlabel polysilicon 205 -168 205 -168 0 1
rlabel polysilicon 205 -174 205 -174 0 3
rlabel polysilicon 212 -168 212 -168 0 1
rlabel polysilicon 212 -174 212 -174 0 3
rlabel polysilicon 219 -174 219 -174 0 3
rlabel polysilicon 222 -174 222 -174 0 4
rlabel polysilicon 226 -168 226 -168 0 1
rlabel polysilicon 229 -168 229 -168 0 2
rlabel polysilicon 233 -168 233 -168 0 1
rlabel polysilicon 233 -174 233 -174 0 3
rlabel polysilicon 243 -168 243 -168 0 2
rlabel polysilicon 240 -174 240 -174 0 3
rlabel polysilicon 243 -174 243 -174 0 4
rlabel polysilicon 247 -168 247 -168 0 1
rlabel polysilicon 247 -174 247 -174 0 3
rlabel polysilicon 254 -168 254 -168 0 1
rlabel polysilicon 254 -174 254 -174 0 3
rlabel polysilicon 261 -168 261 -168 0 1
rlabel polysilicon 261 -174 261 -174 0 3
rlabel polysilicon 268 -168 268 -168 0 1
rlabel polysilicon 268 -174 268 -174 0 3
rlabel polysilicon 275 -168 275 -168 0 1
rlabel polysilicon 275 -174 275 -174 0 3
rlabel polysilicon 285 -168 285 -168 0 2
rlabel polysilicon 285 -174 285 -174 0 4
rlabel polysilicon 289 -168 289 -168 0 1
rlabel polysilicon 289 -174 289 -174 0 3
rlabel polysilicon 296 -168 296 -168 0 1
rlabel polysilicon 296 -174 296 -174 0 3
rlabel polysilicon 303 -168 303 -168 0 1
rlabel polysilicon 303 -174 303 -174 0 3
rlabel polysilicon 313 -174 313 -174 0 4
rlabel polysilicon 317 -168 317 -168 0 1
rlabel polysilicon 317 -174 317 -174 0 3
rlabel polysilicon 320 -174 320 -174 0 4
rlabel polysilicon 324 -168 324 -168 0 1
rlabel polysilicon 324 -174 324 -174 0 3
rlabel polysilicon 331 -168 331 -168 0 1
rlabel polysilicon 331 -174 331 -174 0 3
rlabel polysilicon 341 -168 341 -168 0 2
rlabel polysilicon 341 -174 341 -174 0 4
rlabel polysilicon 345 -168 345 -168 0 1
rlabel polysilicon 345 -174 345 -174 0 3
rlabel polysilicon 352 -168 352 -168 0 1
rlabel polysilicon 352 -174 352 -174 0 3
rlabel polysilicon 359 -168 359 -168 0 1
rlabel polysilicon 359 -174 359 -174 0 3
rlabel polysilicon 366 -168 366 -168 0 1
rlabel polysilicon 366 -174 366 -174 0 3
rlabel polysilicon 373 -168 373 -168 0 1
rlabel polysilicon 380 -168 380 -168 0 1
rlabel polysilicon 380 -174 380 -174 0 3
rlabel polysilicon 387 -168 387 -168 0 1
rlabel polysilicon 387 -174 387 -174 0 3
rlabel polysilicon 394 -168 394 -168 0 1
rlabel polysilicon 394 -174 394 -174 0 3
rlabel polysilicon 401 -168 401 -168 0 1
rlabel polysilicon 401 -174 401 -174 0 3
rlabel polysilicon 408 -168 408 -168 0 1
rlabel polysilicon 408 -174 408 -174 0 3
rlabel polysilicon 415 -168 415 -168 0 1
rlabel polysilicon 415 -174 415 -174 0 3
rlabel polysilicon 422 -168 422 -168 0 1
rlabel polysilicon 422 -174 422 -174 0 3
rlabel polysilicon 429 -168 429 -168 0 1
rlabel polysilicon 432 -174 432 -174 0 4
rlabel polysilicon 439 -174 439 -174 0 4
rlabel polysilicon 23 -207 23 -207 0 1
rlabel polysilicon 23 -213 23 -213 0 3
rlabel polysilicon 30 -207 30 -207 0 1
rlabel polysilicon 30 -213 30 -213 0 3
rlabel polysilicon 37 -207 37 -207 0 1
rlabel polysilicon 37 -213 37 -213 0 3
rlabel polysilicon 44 -207 44 -207 0 1
rlabel polysilicon 44 -213 44 -213 0 3
rlabel polysilicon 51 -207 51 -207 0 1
rlabel polysilicon 51 -213 51 -213 0 3
rlabel polysilicon 58 -213 58 -213 0 3
rlabel polysilicon 65 -207 65 -207 0 1
rlabel polysilicon 68 -207 68 -207 0 2
rlabel polysilicon 65 -213 65 -213 0 3
rlabel polysilicon 72 -207 72 -207 0 1
rlabel polysilicon 79 -207 79 -207 0 1
rlabel polysilicon 79 -213 79 -213 0 3
rlabel polysilicon 86 -207 86 -207 0 1
rlabel polysilicon 89 -213 89 -213 0 4
rlabel polysilicon 96 -207 96 -207 0 2
rlabel polysilicon 93 -213 93 -213 0 3
rlabel polysilicon 100 -207 100 -207 0 1
rlabel polysilicon 100 -213 100 -213 0 3
rlabel polysilicon 107 -207 107 -207 0 1
rlabel polysilicon 107 -213 107 -213 0 3
rlabel polysilicon 114 -207 114 -207 0 1
rlabel polysilicon 114 -213 114 -213 0 3
rlabel polysilicon 121 -207 121 -207 0 1
rlabel polysilicon 121 -213 121 -213 0 3
rlabel polysilicon 128 -207 128 -207 0 1
rlabel polysilicon 128 -213 128 -213 0 3
rlabel polysilicon 135 -207 135 -207 0 1
rlabel polysilicon 135 -213 135 -213 0 3
rlabel polysilicon 138 -213 138 -213 0 4
rlabel polysilicon 142 -207 142 -207 0 1
rlabel polysilicon 145 -207 145 -207 0 2
rlabel polysilicon 142 -213 142 -213 0 3
rlabel polysilicon 145 -213 145 -213 0 4
rlabel polysilicon 149 -207 149 -207 0 1
rlabel polysilicon 152 -207 152 -207 0 2
rlabel polysilicon 156 -207 156 -207 0 1
rlabel polysilicon 159 -207 159 -207 0 2
rlabel polysilicon 159 -213 159 -213 0 4
rlabel polysilicon 163 -207 163 -207 0 1
rlabel polysilicon 163 -213 163 -213 0 3
rlabel polysilicon 170 -207 170 -207 0 1
rlabel polysilicon 170 -213 170 -213 0 3
rlabel polysilicon 177 -207 177 -207 0 1
rlabel polysilicon 177 -213 177 -213 0 3
rlabel polysilicon 184 -207 184 -207 0 1
rlabel polysilicon 184 -213 184 -213 0 3
rlabel polysilicon 191 -207 191 -207 0 1
rlabel polysilicon 194 -207 194 -207 0 2
rlabel polysilicon 191 -213 191 -213 0 3
rlabel polysilicon 198 -207 198 -207 0 1
rlabel polysilicon 201 -213 201 -213 0 4
rlabel polysilicon 205 -207 205 -207 0 1
rlabel polysilicon 205 -213 205 -213 0 3
rlabel polysilicon 208 -213 208 -213 0 4
rlabel polysilicon 215 -207 215 -207 0 2
rlabel polysilicon 215 -213 215 -213 0 4
rlabel polysilicon 219 -207 219 -207 0 1
rlabel polysilicon 219 -213 219 -213 0 3
rlabel polysilicon 226 -207 226 -207 0 1
rlabel polysilicon 226 -213 226 -213 0 3
rlabel polysilicon 233 -207 233 -207 0 1
rlabel polysilicon 236 -207 236 -207 0 2
rlabel polysilicon 236 -213 236 -213 0 4
rlabel polysilicon 243 -207 243 -207 0 2
rlabel polysilicon 240 -213 240 -213 0 3
rlabel polysilicon 243 -213 243 -213 0 4
rlabel polysilicon 247 -207 247 -207 0 1
rlabel polysilicon 247 -213 247 -213 0 3
rlabel polysilicon 254 -207 254 -207 0 1
rlabel polysilicon 254 -213 254 -213 0 3
rlabel polysilicon 261 -207 261 -207 0 1
rlabel polysilicon 261 -213 261 -213 0 3
rlabel polysilicon 268 -207 268 -207 0 1
rlabel polysilicon 271 -207 271 -207 0 2
rlabel polysilicon 268 -213 268 -213 0 3
rlabel polysilicon 271 -213 271 -213 0 4
rlabel polysilicon 275 -207 275 -207 0 1
rlabel polysilicon 275 -213 275 -213 0 3
rlabel polysilicon 285 -207 285 -207 0 2
rlabel polysilicon 282 -213 282 -213 0 3
rlabel polysilicon 289 -207 289 -207 0 1
rlabel polysilicon 289 -213 289 -213 0 3
rlabel polysilicon 296 -207 296 -207 0 1
rlabel polysilicon 299 -213 299 -213 0 4
rlabel polysilicon 303 -207 303 -207 0 1
rlabel polysilicon 303 -213 303 -213 0 3
rlabel polysilicon 310 -207 310 -207 0 1
rlabel polysilicon 310 -213 310 -213 0 3
rlabel polysilicon 317 -207 317 -207 0 1
rlabel polysilicon 317 -213 317 -213 0 3
rlabel polysilicon 324 -207 324 -207 0 1
rlabel polysilicon 331 -207 331 -207 0 1
rlabel polysilicon 331 -213 331 -213 0 3
rlabel polysilicon 341 -207 341 -207 0 2
rlabel polysilicon 338 -213 338 -213 0 3
rlabel polysilicon 345 -207 345 -207 0 1
rlabel polysilicon 345 -213 345 -213 0 3
rlabel polysilicon 352 -207 352 -207 0 1
rlabel polysilicon 352 -213 352 -213 0 3
rlabel polysilicon 359 -207 359 -207 0 1
rlabel polysilicon 359 -213 359 -213 0 3
rlabel polysilicon 366 -207 366 -207 0 1
rlabel polysilicon 366 -213 366 -213 0 3
rlabel polysilicon 373 -207 373 -207 0 1
rlabel polysilicon 380 -207 380 -207 0 1
rlabel polysilicon 380 -213 380 -213 0 3
rlabel polysilicon 387 -207 387 -207 0 1
rlabel polysilicon 387 -213 387 -213 0 3
rlabel polysilicon 394 -207 394 -207 0 1
rlabel polysilicon 394 -213 394 -213 0 3
rlabel polysilicon 401 -207 401 -207 0 1
rlabel polysilicon 401 -213 401 -213 0 3
rlabel polysilicon 411 -207 411 -207 0 2
rlabel polysilicon 408 -213 408 -213 0 3
rlabel polysilicon 415 -207 415 -207 0 1
rlabel polysilicon 415 -213 415 -213 0 3
rlabel polysilicon 422 -207 422 -207 0 1
rlabel polysilicon 422 -213 422 -213 0 3
rlabel polysilicon 429 -207 429 -207 0 1
rlabel polysilicon 429 -213 429 -213 0 3
rlabel polysilicon 436 -207 436 -207 0 1
rlabel polysilicon 436 -213 436 -213 0 3
rlabel polysilicon 443 -207 443 -207 0 1
rlabel polysilicon 443 -213 443 -213 0 3
rlabel polysilicon 450 -207 450 -207 0 1
rlabel polysilicon 450 -213 450 -213 0 3
rlabel polysilicon 457 -207 457 -207 0 1
rlabel polysilicon 457 -213 457 -213 0 3
rlabel polysilicon 464 -207 464 -207 0 1
rlabel polysilicon 464 -213 464 -213 0 3
rlabel polysilicon 544 -213 544 -213 0 4
rlabel polysilicon 37 -254 37 -254 0 1
rlabel polysilicon 37 -260 37 -260 0 3
rlabel polysilicon 44 -254 44 -254 0 1
rlabel polysilicon 44 -260 44 -260 0 3
rlabel polysilicon 51 -254 51 -254 0 1
rlabel polysilicon 51 -260 51 -260 0 3
rlabel polysilicon 58 -254 58 -254 0 1
rlabel polysilicon 58 -260 58 -260 0 3
rlabel polysilicon 65 -254 65 -254 0 1
rlabel polysilicon 65 -260 65 -260 0 3
rlabel polysilicon 72 -254 72 -254 0 1
rlabel polysilicon 72 -260 72 -260 0 3
rlabel polysilicon 75 -260 75 -260 0 4
rlabel polysilicon 79 -254 79 -254 0 1
rlabel polysilicon 79 -260 79 -260 0 3
rlabel polysilicon 86 -254 86 -254 0 1
rlabel polysilicon 86 -260 86 -260 0 3
rlabel polysilicon 93 -254 93 -254 0 1
rlabel polysilicon 93 -260 93 -260 0 3
rlabel polysilicon 100 -254 100 -254 0 1
rlabel polysilicon 100 -260 100 -260 0 3
rlabel polysilicon 110 -254 110 -254 0 2
rlabel polysilicon 107 -260 107 -260 0 3
rlabel polysilicon 114 -260 114 -260 0 3
rlabel polysilicon 117 -260 117 -260 0 4
rlabel polysilicon 121 -254 121 -254 0 1
rlabel polysilicon 124 -254 124 -254 0 2
rlabel polysilicon 128 -260 128 -260 0 3
rlabel polysilicon 131 -260 131 -260 0 4
rlabel polysilicon 135 -254 135 -254 0 1
rlabel polysilicon 135 -260 135 -260 0 3
rlabel polysilicon 142 -254 142 -254 0 1
rlabel polysilicon 145 -260 145 -260 0 4
rlabel polysilicon 149 -254 149 -254 0 1
rlabel polysilicon 152 -254 152 -254 0 2
rlabel polysilicon 149 -260 149 -260 0 3
rlabel polysilicon 152 -260 152 -260 0 4
rlabel polysilicon 156 -254 156 -254 0 1
rlabel polysilicon 156 -260 156 -260 0 3
rlabel polysilicon 163 -254 163 -254 0 1
rlabel polysilicon 166 -254 166 -254 0 2
rlabel polysilicon 166 -260 166 -260 0 4
rlabel polysilicon 170 -254 170 -254 0 1
rlabel polysilicon 173 -260 173 -260 0 4
rlabel polysilicon 177 -254 177 -254 0 1
rlabel polysilicon 180 -254 180 -254 0 2
rlabel polysilicon 177 -260 177 -260 0 3
rlabel polysilicon 184 -254 184 -254 0 1
rlabel polysilicon 184 -260 184 -260 0 3
rlabel polysilicon 191 -254 191 -254 0 1
rlabel polysilicon 191 -260 191 -260 0 3
rlabel polysilicon 198 -254 198 -254 0 1
rlabel polysilicon 201 -254 201 -254 0 2
rlabel polysilicon 205 -254 205 -254 0 1
rlabel polysilicon 208 -254 208 -254 0 2
rlabel polysilicon 205 -260 205 -260 0 3
rlabel polysilicon 208 -260 208 -260 0 4
rlabel polysilicon 212 -254 212 -254 0 1
rlabel polysilicon 212 -260 212 -260 0 3
rlabel polysilicon 219 -254 219 -254 0 1
rlabel polysilicon 219 -260 219 -260 0 3
rlabel polysilicon 226 -254 226 -254 0 1
rlabel polysilicon 229 -254 229 -254 0 2
rlabel polysilicon 226 -260 226 -260 0 3
rlabel polysilicon 229 -260 229 -260 0 4
rlabel polysilicon 233 -254 233 -254 0 1
rlabel polysilicon 240 -254 240 -254 0 1
rlabel polysilicon 243 -254 243 -254 0 2
rlabel polysilicon 243 -260 243 -260 0 4
rlabel polysilicon 247 -254 247 -254 0 1
rlabel polysilicon 247 -260 247 -260 0 3
rlabel polysilicon 254 -254 254 -254 0 1
rlabel polysilicon 254 -260 254 -260 0 3
rlabel polysilicon 261 -254 261 -254 0 1
rlabel polysilicon 261 -260 261 -260 0 3
rlabel polysilicon 268 -254 268 -254 0 1
rlabel polysilicon 268 -260 268 -260 0 3
rlabel polysilicon 275 -254 275 -254 0 1
rlabel polysilicon 275 -260 275 -260 0 3
rlabel polysilicon 282 -254 282 -254 0 1
rlabel polysilicon 285 -254 285 -254 0 2
rlabel polysilicon 282 -260 282 -260 0 3
rlabel polysilicon 289 -254 289 -254 0 1
rlabel polysilicon 289 -260 289 -260 0 3
rlabel polysilicon 296 -254 296 -254 0 1
rlabel polysilicon 296 -260 296 -260 0 3
rlabel polysilicon 306 -254 306 -254 0 2
rlabel polysilicon 303 -260 303 -260 0 3
rlabel polysilicon 310 -254 310 -254 0 1
rlabel polysilicon 310 -260 310 -260 0 3
rlabel polysilicon 317 -254 317 -254 0 1
rlabel polysilicon 317 -260 317 -260 0 3
rlabel polysilicon 324 -254 324 -254 0 1
rlabel polysilicon 327 -254 327 -254 0 2
rlabel polysilicon 331 -254 331 -254 0 1
rlabel polysilicon 331 -260 331 -260 0 3
rlabel polysilicon 334 -260 334 -260 0 4
rlabel polysilicon 338 -254 338 -254 0 1
rlabel polysilicon 341 -254 341 -254 0 2
rlabel polysilicon 338 -260 338 -260 0 3
rlabel polysilicon 348 -254 348 -254 0 2
rlabel polysilicon 345 -260 345 -260 0 3
rlabel polysilicon 348 -260 348 -260 0 4
rlabel polysilicon 355 -254 355 -254 0 2
rlabel polysilicon 352 -260 352 -260 0 3
rlabel polysilicon 359 -254 359 -254 0 1
rlabel polysilicon 359 -260 359 -260 0 3
rlabel polysilicon 366 -254 366 -254 0 1
rlabel polysilicon 366 -260 366 -260 0 3
rlabel polysilicon 373 -254 373 -254 0 1
rlabel polysilicon 373 -260 373 -260 0 3
rlabel polysilicon 380 -254 380 -254 0 1
rlabel polysilicon 380 -260 380 -260 0 3
rlabel polysilicon 387 -254 387 -254 0 1
rlabel polysilicon 387 -260 387 -260 0 3
rlabel polysilicon 394 -254 394 -254 0 1
rlabel polysilicon 394 -260 394 -260 0 3
rlabel polysilicon 401 -254 401 -254 0 1
rlabel polysilicon 401 -260 401 -260 0 3
rlabel polysilicon 408 -254 408 -254 0 1
rlabel polysilicon 408 -260 408 -260 0 3
rlabel polysilicon 415 -254 415 -254 0 1
rlabel polysilicon 415 -260 415 -260 0 3
rlabel polysilicon 422 -254 422 -254 0 1
rlabel polysilicon 422 -260 422 -260 0 3
rlabel polysilicon 429 -254 429 -254 0 1
rlabel polysilicon 429 -260 429 -260 0 3
rlabel polysilicon 436 -254 436 -254 0 1
rlabel polysilicon 436 -260 436 -260 0 3
rlabel polysilicon 443 -254 443 -254 0 1
rlabel polysilicon 443 -260 443 -260 0 3
rlabel polysilicon 450 -254 450 -254 0 1
rlabel polysilicon 450 -260 450 -260 0 3
rlabel polysilicon 457 -254 457 -254 0 1
rlabel polysilicon 457 -260 457 -260 0 3
rlabel polysilicon 464 -254 464 -254 0 1
rlabel polysilicon 464 -260 464 -260 0 3
rlabel polysilicon 471 -254 471 -254 0 1
rlabel polysilicon 471 -260 471 -260 0 3
rlabel polysilicon 478 -254 478 -254 0 1
rlabel polysilicon 478 -260 478 -260 0 3
rlabel polysilicon 485 -254 485 -254 0 1
rlabel polysilicon 485 -260 485 -260 0 3
rlabel polysilicon 492 -254 492 -254 0 1
rlabel polysilicon 492 -260 492 -260 0 3
rlabel polysilicon 499 -254 499 -254 0 1
rlabel polysilicon 499 -260 499 -260 0 3
rlabel polysilicon 506 -254 506 -254 0 1
rlabel polysilicon 506 -260 506 -260 0 3
rlabel polysilicon 513 -254 513 -254 0 1
rlabel polysilicon 513 -260 513 -260 0 3
rlabel polysilicon 520 -254 520 -254 0 1
rlabel polysilicon 520 -260 520 -260 0 3
rlabel polysilicon 527 -260 527 -260 0 3
rlabel polysilicon 534 -254 534 -254 0 1
rlabel polysilicon 537 -254 537 -254 0 2
rlabel polysilicon 534 -260 534 -260 0 3
rlabel polysilicon 541 -254 541 -254 0 1
rlabel polysilicon 541 -260 541 -260 0 3
rlabel polysilicon 37 -301 37 -301 0 1
rlabel polysilicon 37 -307 37 -307 0 3
rlabel polysilicon 44 -307 44 -307 0 3
rlabel polysilicon 51 -301 51 -301 0 1
rlabel polysilicon 51 -307 51 -307 0 3
rlabel polysilicon 61 -307 61 -307 0 4
rlabel polysilicon 65 -301 65 -301 0 1
rlabel polysilicon 65 -307 65 -307 0 3
rlabel polysilicon 72 -301 72 -301 0 1
rlabel polysilicon 72 -307 72 -307 0 3
rlabel polysilicon 79 -301 79 -301 0 1
rlabel polysilicon 86 -301 86 -301 0 1
rlabel polysilicon 86 -307 86 -307 0 3
rlabel polysilicon 96 -301 96 -301 0 2
rlabel polysilicon 96 -307 96 -307 0 4
rlabel polysilicon 100 -301 100 -301 0 1
rlabel polysilicon 100 -307 100 -307 0 3
rlabel polysilicon 107 -301 107 -301 0 1
rlabel polysilicon 107 -307 107 -307 0 3
rlabel polysilicon 114 -301 114 -301 0 1
rlabel polysilicon 117 -301 117 -301 0 2
rlabel polysilicon 114 -307 114 -307 0 3
rlabel polysilicon 121 -301 121 -301 0 1
rlabel polysilicon 121 -307 121 -307 0 3
rlabel polysilicon 128 -301 128 -301 0 1
rlabel polysilicon 131 -307 131 -307 0 4
rlabel polysilicon 135 -301 135 -301 0 1
rlabel polysilicon 135 -307 135 -307 0 3
rlabel polysilicon 142 -301 142 -301 0 1
rlabel polysilicon 142 -307 142 -307 0 3
rlabel polysilicon 149 -301 149 -301 0 1
rlabel polysilicon 149 -307 149 -307 0 3
rlabel polysilicon 156 -301 156 -301 0 1
rlabel polysilicon 156 -307 156 -307 0 3
rlabel polysilicon 163 -301 163 -301 0 1
rlabel polysilicon 163 -307 163 -307 0 3
rlabel polysilicon 170 -301 170 -301 0 1
rlabel polysilicon 170 -307 170 -307 0 3
rlabel polysilicon 177 -301 177 -301 0 1
rlabel polysilicon 177 -307 177 -307 0 3
rlabel polysilicon 184 -301 184 -301 0 1
rlabel polysilicon 184 -307 184 -307 0 3
rlabel polysilicon 191 -301 191 -301 0 1
rlabel polysilicon 191 -307 191 -307 0 3
rlabel polysilicon 194 -307 194 -307 0 4
rlabel polysilicon 198 -301 198 -301 0 1
rlabel polysilicon 198 -307 198 -307 0 3
rlabel polysilicon 205 -301 205 -301 0 1
rlabel polysilicon 205 -307 205 -307 0 3
rlabel polysilicon 212 -301 212 -301 0 1
rlabel polysilicon 212 -307 212 -307 0 3
rlabel polysilicon 219 -301 219 -301 0 1
rlabel polysilicon 219 -307 219 -307 0 3
rlabel polysilicon 226 -301 226 -301 0 1
rlabel polysilicon 226 -307 226 -307 0 3
rlabel polysilicon 233 -301 233 -301 0 1
rlabel polysilicon 233 -307 233 -307 0 3
rlabel polysilicon 240 -301 240 -301 0 1
rlabel polysilicon 240 -307 240 -307 0 3
rlabel polysilicon 247 -301 247 -301 0 1
rlabel polysilicon 247 -307 247 -307 0 3
rlabel polysilicon 250 -307 250 -307 0 4
rlabel polysilicon 254 -301 254 -301 0 1
rlabel polysilicon 254 -307 254 -307 0 3
rlabel polysilicon 261 -301 261 -301 0 1
rlabel polysilicon 261 -307 261 -307 0 3
rlabel polysilicon 268 -301 268 -301 0 1
rlabel polysilicon 268 -307 268 -307 0 3
rlabel polysilicon 271 -307 271 -307 0 4
rlabel polysilicon 275 -301 275 -301 0 1
rlabel polysilicon 275 -307 275 -307 0 3
rlabel polysilicon 285 -301 285 -301 0 2
rlabel polysilicon 282 -307 282 -307 0 3
rlabel polysilicon 285 -307 285 -307 0 4
rlabel polysilicon 289 -301 289 -301 0 1
rlabel polysilicon 289 -307 289 -307 0 3
rlabel polysilicon 296 -301 296 -301 0 1
rlabel polysilicon 296 -307 296 -307 0 3
rlabel polysilicon 303 -301 303 -301 0 1
rlabel polysilicon 306 -301 306 -301 0 2
rlabel polysilicon 303 -307 303 -307 0 3
rlabel polysilicon 310 -301 310 -301 0 1
rlabel polysilicon 310 -307 310 -307 0 3
rlabel polysilicon 317 -301 317 -301 0 1
rlabel polysilicon 320 -301 320 -301 0 2
rlabel polysilicon 317 -307 317 -307 0 3
rlabel polysilicon 324 -301 324 -301 0 1
rlabel polysilicon 324 -307 324 -307 0 3
rlabel polysilicon 334 -301 334 -301 0 2
rlabel polysilicon 334 -307 334 -307 0 4
rlabel polysilicon 338 -307 338 -307 0 3
rlabel polysilicon 345 -307 345 -307 0 3
rlabel polysilicon 348 -307 348 -307 0 4
rlabel polysilicon 352 -301 352 -301 0 1
rlabel polysilicon 352 -307 352 -307 0 3
rlabel polysilicon 362 -301 362 -301 0 2
rlabel polysilicon 366 -301 366 -301 0 1
rlabel polysilicon 366 -307 366 -307 0 3
rlabel polysilicon 373 -301 373 -301 0 1
rlabel polysilicon 373 -307 373 -307 0 3
rlabel polysilicon 383 -301 383 -301 0 2
rlabel polysilicon 383 -307 383 -307 0 4
rlabel polysilicon 387 -301 387 -301 0 1
rlabel polysilicon 387 -307 387 -307 0 3
rlabel polysilicon 394 -301 394 -301 0 1
rlabel polysilicon 394 -307 394 -307 0 3
rlabel polysilicon 401 -301 401 -301 0 1
rlabel polysilicon 401 -307 401 -307 0 3
rlabel polysilicon 408 -301 408 -301 0 1
rlabel polysilicon 408 -307 408 -307 0 3
rlabel polysilicon 415 -301 415 -301 0 1
rlabel polysilicon 415 -307 415 -307 0 3
rlabel polysilicon 422 -301 422 -301 0 1
rlabel polysilicon 422 -307 422 -307 0 3
rlabel polysilicon 429 -301 429 -301 0 1
rlabel polysilicon 429 -307 429 -307 0 3
rlabel polysilicon 436 -301 436 -301 0 1
rlabel polysilicon 436 -307 436 -307 0 3
rlabel polysilicon 443 -301 443 -301 0 1
rlabel polysilicon 443 -307 443 -307 0 3
rlabel polysilicon 450 -301 450 -301 0 1
rlabel polysilicon 450 -307 450 -307 0 3
rlabel polysilicon 457 -301 457 -301 0 1
rlabel polysilicon 457 -307 457 -307 0 3
rlabel polysilicon 464 -307 464 -307 0 3
rlabel polysilicon 471 -301 471 -301 0 1
rlabel polysilicon 471 -307 471 -307 0 3
rlabel polysilicon 478 -301 478 -301 0 1
rlabel polysilicon 478 -307 478 -307 0 3
rlabel polysilicon 485 -301 485 -301 0 1
rlabel polysilicon 485 -307 485 -307 0 3
rlabel polysilicon 492 -301 492 -301 0 1
rlabel polysilicon 492 -307 492 -307 0 3
rlabel polysilicon 499 -301 499 -301 0 1
rlabel polysilicon 499 -307 499 -307 0 3
rlabel polysilicon 506 -301 506 -301 0 1
rlabel polysilicon 506 -307 506 -307 0 3
rlabel polysilicon 513 -301 513 -301 0 1
rlabel polysilicon 513 -307 513 -307 0 3
rlabel polysilicon 520 -301 520 -301 0 1
rlabel polysilicon 520 -307 520 -307 0 3
rlabel polysilicon 527 -301 527 -301 0 1
rlabel polysilicon 527 -307 527 -307 0 3
rlabel polysilicon 534 -301 534 -301 0 1
rlabel polysilicon 534 -307 534 -307 0 3
rlabel polysilicon 541 -301 541 -301 0 1
rlabel polysilicon 541 -307 541 -307 0 3
rlabel polysilicon 544 -307 544 -307 0 4
rlabel polysilicon 548 -301 548 -301 0 1
rlabel polysilicon 548 -307 548 -307 0 3
rlabel polysilicon 555 -301 555 -301 0 1
rlabel polysilicon 562 -301 562 -301 0 1
rlabel polysilicon 569 -307 569 -307 0 3
rlabel polysilicon 576 -301 576 -301 0 1
rlabel polysilicon 576 -307 576 -307 0 3
rlabel polysilicon 9 -362 9 -362 0 1
rlabel polysilicon 9 -368 9 -368 0 3
rlabel polysilicon 16 -362 16 -362 0 1
rlabel polysilicon 16 -368 16 -368 0 3
rlabel polysilicon 23 -362 23 -362 0 1
rlabel polysilicon 23 -368 23 -368 0 3
rlabel polysilicon 30 -362 30 -362 0 1
rlabel polysilicon 30 -368 30 -368 0 3
rlabel polysilicon 37 -368 37 -368 0 3
rlabel polysilicon 44 -362 44 -362 0 1
rlabel polysilicon 44 -368 44 -368 0 3
rlabel polysilicon 51 -362 51 -362 0 1
rlabel polysilicon 51 -368 51 -368 0 3
rlabel polysilicon 61 -362 61 -362 0 2
rlabel polysilicon 58 -368 58 -368 0 3
rlabel polysilicon 61 -368 61 -368 0 4
rlabel polysilicon 65 -362 65 -362 0 1
rlabel polysilicon 65 -368 65 -368 0 3
rlabel polysilicon 72 -362 72 -362 0 1
rlabel polysilicon 72 -368 72 -368 0 3
rlabel polysilicon 79 -362 79 -362 0 1
rlabel polysilicon 79 -368 79 -368 0 3
rlabel polysilicon 86 -362 86 -362 0 1
rlabel polysilicon 86 -368 86 -368 0 3
rlabel polysilicon 93 -362 93 -362 0 1
rlabel polysilicon 93 -368 93 -368 0 3
rlabel polysilicon 103 -362 103 -362 0 2
rlabel polysilicon 103 -368 103 -368 0 4
rlabel polysilicon 107 -368 107 -368 0 3
rlabel polysilicon 114 -362 114 -362 0 1
rlabel polysilicon 114 -368 114 -368 0 3
rlabel polysilicon 121 -362 121 -362 0 1
rlabel polysilicon 124 -368 124 -368 0 4
rlabel polysilicon 128 -368 128 -368 0 3
rlabel polysilicon 131 -368 131 -368 0 4
rlabel polysilicon 138 -362 138 -362 0 2
rlabel polysilicon 135 -368 135 -368 0 3
rlabel polysilicon 138 -368 138 -368 0 4
rlabel polysilicon 142 -362 142 -362 0 1
rlabel polysilicon 142 -368 142 -368 0 3
rlabel polysilicon 149 -362 149 -362 0 1
rlabel polysilicon 149 -368 149 -368 0 3
rlabel polysilicon 152 -368 152 -368 0 4
rlabel polysilicon 156 -362 156 -362 0 1
rlabel polysilicon 156 -368 156 -368 0 3
rlabel polysilicon 163 -362 163 -362 0 1
rlabel polysilicon 163 -368 163 -368 0 3
rlabel polysilicon 170 -362 170 -362 0 1
rlabel polysilicon 170 -368 170 -368 0 3
rlabel polysilicon 180 -362 180 -362 0 2
rlabel polysilicon 177 -368 177 -368 0 3
rlabel polysilicon 184 -362 184 -362 0 1
rlabel polysilicon 184 -368 184 -368 0 3
rlabel polysilicon 194 -362 194 -362 0 2
rlabel polysilicon 191 -368 191 -368 0 3
rlabel polysilicon 198 -362 198 -362 0 1
rlabel polysilicon 198 -368 198 -368 0 3
rlabel polysilicon 205 -362 205 -362 0 1
rlabel polysilicon 208 -362 208 -362 0 2
rlabel polysilicon 208 -368 208 -368 0 4
rlabel polysilicon 212 -362 212 -362 0 1
rlabel polysilicon 212 -368 212 -368 0 3
rlabel polysilicon 219 -362 219 -362 0 1
rlabel polysilicon 219 -368 219 -368 0 3
rlabel polysilicon 226 -362 226 -362 0 1
rlabel polysilicon 226 -368 226 -368 0 3
rlabel polysilicon 233 -362 233 -362 0 1
rlabel polysilicon 233 -368 233 -368 0 3
rlabel polysilicon 240 -362 240 -362 0 1
rlabel polysilicon 243 -368 243 -368 0 4
rlabel polysilicon 247 -362 247 -362 0 1
rlabel polysilicon 247 -368 247 -368 0 3
rlabel polysilicon 254 -362 254 -362 0 1
rlabel polysilicon 254 -368 254 -368 0 3
rlabel polysilicon 261 -362 261 -362 0 1
rlabel polysilicon 261 -368 261 -368 0 3
rlabel polysilicon 268 -362 268 -362 0 1
rlabel polysilicon 271 -368 271 -368 0 4
rlabel polysilicon 275 -362 275 -362 0 1
rlabel polysilicon 275 -368 275 -368 0 3
rlabel polysilicon 282 -362 282 -362 0 1
rlabel polysilicon 285 -362 285 -362 0 2
rlabel polysilicon 285 -368 285 -368 0 4
rlabel polysilicon 289 -362 289 -362 0 1
rlabel polysilicon 292 -362 292 -362 0 2
rlabel polysilicon 296 -362 296 -362 0 1
rlabel polysilicon 299 -362 299 -362 0 2
rlabel polysilicon 296 -368 296 -368 0 3
rlabel polysilicon 299 -368 299 -368 0 4
rlabel polysilicon 303 -362 303 -362 0 1
rlabel polysilicon 303 -368 303 -368 0 3
rlabel polysilicon 310 -362 310 -362 0 1
rlabel polysilicon 313 -362 313 -362 0 2
rlabel polysilicon 313 -368 313 -368 0 4
rlabel polysilicon 317 -362 317 -362 0 1
rlabel polysilicon 317 -368 317 -368 0 3
rlabel polysilicon 324 -368 324 -368 0 3
rlabel polysilicon 327 -368 327 -368 0 4
rlabel polysilicon 331 -362 331 -362 0 1
rlabel polysilicon 334 -362 334 -362 0 2
rlabel polysilicon 338 -362 338 -362 0 1
rlabel polysilicon 341 -362 341 -362 0 2
rlabel polysilicon 345 -362 345 -362 0 1
rlabel polysilicon 348 -362 348 -362 0 2
rlabel polysilicon 345 -368 345 -368 0 3
rlabel polysilicon 348 -368 348 -368 0 4
rlabel polysilicon 352 -362 352 -362 0 1
rlabel polysilicon 355 -362 355 -362 0 2
rlabel polysilicon 355 -368 355 -368 0 4
rlabel polysilicon 359 -362 359 -362 0 1
rlabel polysilicon 359 -368 359 -368 0 3
rlabel polysilicon 366 -368 366 -368 0 3
rlabel polysilicon 373 -362 373 -362 0 1
rlabel polysilicon 373 -368 373 -368 0 3
rlabel polysilicon 380 -362 380 -362 0 1
rlabel polysilicon 380 -368 380 -368 0 3
rlabel polysilicon 387 -362 387 -362 0 1
rlabel polysilicon 387 -368 387 -368 0 3
rlabel polysilicon 394 -362 394 -362 0 1
rlabel polysilicon 394 -368 394 -368 0 3
rlabel polysilicon 401 -362 401 -362 0 1
rlabel polysilicon 401 -368 401 -368 0 3
rlabel polysilicon 408 -362 408 -362 0 1
rlabel polysilicon 408 -368 408 -368 0 3
rlabel polysilicon 415 -362 415 -362 0 1
rlabel polysilicon 415 -368 415 -368 0 3
rlabel polysilicon 422 -362 422 -362 0 1
rlabel polysilicon 422 -368 422 -368 0 3
rlabel polysilicon 429 -362 429 -362 0 1
rlabel polysilicon 429 -368 429 -368 0 3
rlabel polysilicon 436 -362 436 -362 0 1
rlabel polysilicon 436 -368 436 -368 0 3
rlabel polysilicon 443 -362 443 -362 0 1
rlabel polysilicon 443 -368 443 -368 0 3
rlabel polysilicon 450 -362 450 -362 0 1
rlabel polysilicon 450 -368 450 -368 0 3
rlabel polysilicon 457 -362 457 -362 0 1
rlabel polysilicon 457 -368 457 -368 0 3
rlabel polysilicon 464 -362 464 -362 0 1
rlabel polysilicon 464 -368 464 -368 0 3
rlabel polysilicon 471 -362 471 -362 0 1
rlabel polysilicon 471 -368 471 -368 0 3
rlabel polysilicon 478 -362 478 -362 0 1
rlabel polysilicon 478 -368 478 -368 0 3
rlabel polysilicon 485 -362 485 -362 0 1
rlabel polysilicon 485 -368 485 -368 0 3
rlabel polysilicon 492 -362 492 -362 0 1
rlabel polysilicon 492 -368 492 -368 0 3
rlabel polysilicon 499 -362 499 -362 0 1
rlabel polysilicon 499 -368 499 -368 0 3
rlabel polysilicon 506 -362 506 -362 0 1
rlabel polysilicon 506 -368 506 -368 0 3
rlabel polysilicon 513 -362 513 -362 0 1
rlabel polysilicon 513 -368 513 -368 0 3
rlabel polysilicon 520 -362 520 -362 0 1
rlabel polysilicon 520 -368 520 -368 0 3
rlabel polysilicon 527 -362 527 -362 0 1
rlabel polysilicon 527 -368 527 -368 0 3
rlabel polysilicon 534 -362 534 -362 0 1
rlabel polysilicon 534 -368 534 -368 0 3
rlabel polysilicon 541 -362 541 -362 0 1
rlabel polysilicon 541 -368 541 -368 0 3
rlabel polysilicon 548 -362 548 -362 0 1
rlabel polysilicon 548 -368 548 -368 0 3
rlabel polysilicon 555 -362 555 -362 0 1
rlabel polysilicon 558 -368 558 -368 0 4
rlabel polysilicon 562 -362 562 -362 0 1
rlabel polysilicon 562 -368 562 -368 0 3
rlabel polysilicon 569 -362 569 -362 0 1
rlabel polysilicon 569 -368 569 -368 0 3
rlabel polysilicon 576 -362 576 -362 0 1
rlabel polysilicon 576 -368 576 -368 0 3
rlabel polysilicon 2 -417 2 -417 0 1
rlabel polysilicon 2 -423 2 -423 0 3
rlabel polysilicon 9 -417 9 -417 0 1
rlabel polysilicon 19 -423 19 -423 0 4
rlabel polysilicon 23 -417 23 -417 0 1
rlabel polysilicon 23 -423 23 -423 0 3
rlabel polysilicon 33 -417 33 -417 0 2
rlabel polysilicon 37 -417 37 -417 0 1
rlabel polysilicon 37 -423 37 -423 0 3
rlabel polysilicon 44 -417 44 -417 0 1
rlabel polysilicon 44 -423 44 -423 0 3
rlabel polysilicon 51 -417 51 -417 0 1
rlabel polysilicon 51 -423 51 -423 0 3
rlabel polysilicon 58 -417 58 -417 0 1
rlabel polysilicon 58 -423 58 -423 0 3
rlabel polysilicon 68 -417 68 -417 0 2
rlabel polysilicon 72 -417 72 -417 0 1
rlabel polysilicon 72 -423 72 -423 0 3
rlabel polysilicon 79 -417 79 -417 0 1
rlabel polysilicon 79 -423 79 -423 0 3
rlabel polysilicon 86 -423 86 -423 0 3
rlabel polysilicon 96 -417 96 -417 0 2
rlabel polysilicon 93 -423 93 -423 0 3
rlabel polysilicon 96 -423 96 -423 0 4
rlabel polysilicon 100 -417 100 -417 0 1
rlabel polysilicon 107 -417 107 -417 0 1
rlabel polysilicon 107 -423 107 -423 0 3
rlabel polysilicon 114 -417 114 -417 0 1
rlabel polysilicon 114 -423 114 -423 0 3
rlabel polysilicon 121 -417 121 -417 0 1
rlabel polysilicon 121 -423 121 -423 0 3
rlabel polysilicon 131 -423 131 -423 0 4
rlabel polysilicon 138 -417 138 -417 0 2
rlabel polysilicon 135 -423 135 -423 0 3
rlabel polysilicon 138 -423 138 -423 0 4
rlabel polysilicon 142 -417 142 -417 0 1
rlabel polysilicon 142 -423 142 -423 0 3
rlabel polysilicon 149 -417 149 -417 0 1
rlabel polysilicon 152 -417 152 -417 0 2
rlabel polysilicon 156 -417 156 -417 0 1
rlabel polysilicon 156 -423 156 -423 0 3
rlabel polysilicon 159 -423 159 -423 0 4
rlabel polysilicon 163 -417 163 -417 0 1
rlabel polysilicon 163 -423 163 -423 0 3
rlabel polysilicon 170 -417 170 -417 0 1
rlabel polysilicon 170 -423 170 -423 0 3
rlabel polysilicon 177 -417 177 -417 0 1
rlabel polysilicon 177 -423 177 -423 0 3
rlabel polysilicon 184 -417 184 -417 0 1
rlabel polysilicon 184 -423 184 -423 0 3
rlabel polysilicon 191 -417 191 -417 0 1
rlabel polysilicon 191 -423 191 -423 0 3
rlabel polysilicon 201 -417 201 -417 0 2
rlabel polysilicon 198 -423 198 -423 0 3
rlabel polysilicon 205 -417 205 -417 0 1
rlabel polysilicon 205 -423 205 -423 0 3
rlabel polysilicon 208 -423 208 -423 0 4
rlabel polysilicon 212 -417 212 -417 0 1
rlabel polysilicon 212 -423 212 -423 0 3
rlabel polysilicon 219 -417 219 -417 0 1
rlabel polysilicon 219 -423 219 -423 0 3
rlabel polysilicon 226 -417 226 -417 0 1
rlabel polysilicon 226 -423 226 -423 0 3
rlabel polysilicon 233 -417 233 -417 0 1
rlabel polysilicon 233 -423 233 -423 0 3
rlabel polysilicon 243 -417 243 -417 0 2
rlabel polysilicon 240 -423 240 -423 0 3
rlabel polysilicon 243 -423 243 -423 0 4
rlabel polysilicon 247 -417 247 -417 0 1
rlabel polysilicon 250 -417 250 -417 0 2
rlabel polysilicon 250 -423 250 -423 0 4
rlabel polysilicon 254 -423 254 -423 0 3
rlabel polysilicon 257 -423 257 -423 0 4
rlabel polysilicon 261 -417 261 -417 0 1
rlabel polysilicon 261 -423 261 -423 0 3
rlabel polysilicon 268 -417 268 -417 0 1
rlabel polysilicon 268 -423 268 -423 0 3
rlabel polysilicon 271 -423 271 -423 0 4
rlabel polysilicon 275 -417 275 -417 0 1
rlabel polysilicon 275 -423 275 -423 0 3
rlabel polysilicon 278 -423 278 -423 0 4
rlabel polysilicon 282 -417 282 -417 0 1
rlabel polysilicon 282 -423 282 -423 0 3
rlabel polysilicon 289 -423 289 -423 0 3
rlabel polysilicon 296 -417 296 -417 0 1
rlabel polysilicon 296 -423 296 -423 0 3
rlabel polysilicon 306 -417 306 -417 0 2
rlabel polysilicon 310 -417 310 -417 0 1
rlabel polysilicon 310 -423 310 -423 0 3
rlabel polysilicon 320 -417 320 -417 0 2
rlabel polysilicon 317 -423 317 -423 0 3
rlabel polysilicon 320 -423 320 -423 0 4
rlabel polysilicon 327 -417 327 -417 0 2
rlabel polysilicon 324 -423 324 -423 0 3
rlabel polysilicon 327 -423 327 -423 0 4
rlabel polysilicon 331 -417 331 -417 0 1
rlabel polysilicon 331 -423 331 -423 0 3
rlabel polysilicon 338 -417 338 -417 0 1
rlabel polysilicon 338 -423 338 -423 0 3
rlabel polysilicon 348 -417 348 -417 0 2
rlabel polysilicon 348 -423 348 -423 0 4
rlabel polysilicon 352 -417 352 -417 0 1
rlabel polysilicon 352 -423 352 -423 0 3
rlabel polysilicon 359 -423 359 -423 0 3
rlabel polysilicon 362 -423 362 -423 0 4
rlabel polysilicon 366 -417 366 -417 0 1
rlabel polysilicon 366 -423 366 -423 0 3
rlabel polysilicon 373 -417 373 -417 0 1
rlabel polysilicon 373 -423 373 -423 0 3
rlabel polysilicon 380 -417 380 -417 0 1
rlabel polysilicon 383 -417 383 -417 0 2
rlabel polysilicon 380 -423 380 -423 0 3
rlabel polysilicon 383 -423 383 -423 0 4
rlabel polysilicon 387 -417 387 -417 0 1
rlabel polysilicon 390 -417 390 -417 0 2
rlabel polysilicon 394 -417 394 -417 0 1
rlabel polysilicon 394 -423 394 -423 0 3
rlabel polysilicon 401 -417 401 -417 0 1
rlabel polysilicon 401 -423 401 -423 0 3
rlabel polysilicon 408 -417 408 -417 0 1
rlabel polysilicon 411 -417 411 -417 0 2
rlabel polysilicon 415 -417 415 -417 0 1
rlabel polysilicon 415 -423 415 -423 0 3
rlabel polysilicon 422 -417 422 -417 0 1
rlabel polysilicon 422 -423 422 -423 0 3
rlabel polysilicon 429 -417 429 -417 0 1
rlabel polysilicon 429 -423 429 -423 0 3
rlabel polysilicon 436 -417 436 -417 0 1
rlabel polysilicon 436 -423 436 -423 0 3
rlabel polysilicon 443 -417 443 -417 0 1
rlabel polysilicon 443 -423 443 -423 0 3
rlabel polysilicon 450 -417 450 -417 0 1
rlabel polysilicon 450 -423 450 -423 0 3
rlabel polysilicon 457 -417 457 -417 0 1
rlabel polysilicon 457 -423 457 -423 0 3
rlabel polysilicon 464 -417 464 -417 0 1
rlabel polysilicon 464 -423 464 -423 0 3
rlabel polysilicon 471 -417 471 -417 0 1
rlabel polysilicon 471 -423 471 -423 0 3
rlabel polysilicon 478 -417 478 -417 0 1
rlabel polysilicon 478 -423 478 -423 0 3
rlabel polysilicon 485 -417 485 -417 0 1
rlabel polysilicon 485 -423 485 -423 0 3
rlabel polysilicon 492 -417 492 -417 0 1
rlabel polysilicon 492 -423 492 -423 0 3
rlabel polysilicon 499 -417 499 -417 0 1
rlabel polysilicon 499 -423 499 -423 0 3
rlabel polysilicon 506 -417 506 -417 0 1
rlabel polysilicon 506 -423 506 -423 0 3
rlabel polysilicon 513 -417 513 -417 0 1
rlabel polysilicon 513 -423 513 -423 0 3
rlabel polysilicon 523 -417 523 -417 0 2
rlabel polysilicon 527 -417 527 -417 0 1
rlabel polysilicon 527 -423 527 -423 0 3
rlabel polysilicon 534 -417 534 -417 0 1
rlabel polysilicon 534 -423 534 -423 0 3
rlabel polysilicon 541 -417 541 -417 0 1
rlabel polysilicon 541 -423 541 -423 0 3
rlabel polysilicon 548 -417 548 -417 0 1
rlabel polysilicon 548 -423 548 -423 0 3
rlabel polysilicon 555 -417 555 -417 0 1
rlabel polysilicon 555 -423 555 -423 0 3
rlabel polysilicon 562 -417 562 -417 0 1
rlabel polysilicon 562 -423 562 -423 0 3
rlabel polysilicon 569 -417 569 -417 0 1
rlabel polysilicon 569 -423 569 -423 0 3
rlabel polysilicon 576 -417 576 -417 0 1
rlabel polysilicon 576 -423 576 -423 0 3
rlabel polysilicon 583 -417 583 -417 0 1
rlabel polysilicon 583 -423 583 -423 0 3
rlabel polysilicon 611 -417 611 -417 0 1
rlabel polysilicon 611 -423 611 -423 0 3
rlabel polysilicon 2 -494 2 -494 0 1
rlabel polysilicon 2 -500 2 -500 0 3
rlabel polysilicon 9 -494 9 -494 0 1
rlabel polysilicon 9 -500 9 -500 0 3
rlabel polysilicon 16 -494 16 -494 0 1
rlabel polysilicon 16 -500 16 -500 0 3
rlabel polysilicon 23 -494 23 -494 0 1
rlabel polysilicon 23 -500 23 -500 0 3
rlabel polysilicon 30 -494 30 -494 0 1
rlabel polysilicon 30 -500 30 -500 0 3
rlabel polysilicon 37 -494 37 -494 0 1
rlabel polysilicon 40 -494 40 -494 0 2
rlabel polysilicon 44 -494 44 -494 0 1
rlabel polysilicon 47 -494 47 -494 0 2
rlabel polysilicon 47 -500 47 -500 0 4
rlabel polysilicon 51 -494 51 -494 0 1
rlabel polysilicon 51 -500 51 -500 0 3
rlabel polysilicon 58 -494 58 -494 0 1
rlabel polysilicon 58 -500 58 -500 0 3
rlabel polysilicon 68 -494 68 -494 0 2
rlabel polysilicon 72 -494 72 -494 0 1
rlabel polysilicon 72 -500 72 -500 0 3
rlabel polysilicon 79 -494 79 -494 0 1
rlabel polysilicon 79 -500 79 -500 0 3
rlabel polysilicon 86 -494 86 -494 0 1
rlabel polysilicon 86 -500 86 -500 0 3
rlabel polysilicon 93 -494 93 -494 0 1
rlabel polysilicon 93 -500 93 -500 0 3
rlabel polysilicon 100 -494 100 -494 0 1
rlabel polysilicon 100 -500 100 -500 0 3
rlabel polysilicon 107 -494 107 -494 0 1
rlabel polysilicon 107 -500 107 -500 0 3
rlabel polysilicon 114 -494 114 -494 0 1
rlabel polysilicon 117 -494 117 -494 0 2
rlabel polysilicon 124 -494 124 -494 0 2
rlabel polysilicon 124 -500 124 -500 0 4
rlabel polysilicon 128 -494 128 -494 0 1
rlabel polysilicon 131 -494 131 -494 0 2
rlabel polysilicon 128 -500 128 -500 0 3
rlabel polysilicon 131 -500 131 -500 0 4
rlabel polysilicon 135 -494 135 -494 0 1
rlabel polysilicon 138 -494 138 -494 0 2
rlabel polysilicon 142 -494 142 -494 0 1
rlabel polysilicon 145 -494 145 -494 0 2
rlabel polysilicon 142 -500 142 -500 0 3
rlabel polysilicon 149 -494 149 -494 0 1
rlabel polysilicon 149 -500 149 -500 0 3
rlabel polysilicon 156 -494 156 -494 0 1
rlabel polysilicon 156 -500 156 -500 0 3
rlabel polysilicon 163 -494 163 -494 0 1
rlabel polysilicon 163 -500 163 -500 0 3
rlabel polysilicon 170 -494 170 -494 0 1
rlabel polysilicon 173 -494 173 -494 0 2
rlabel polysilicon 170 -500 170 -500 0 3
rlabel polysilicon 177 -494 177 -494 0 1
rlabel polysilicon 177 -500 177 -500 0 3
rlabel polysilicon 187 -494 187 -494 0 2
rlabel polysilicon 191 -494 191 -494 0 1
rlabel polysilicon 191 -500 191 -500 0 3
rlabel polysilicon 201 -494 201 -494 0 2
rlabel polysilicon 198 -500 198 -500 0 3
rlabel polysilicon 205 -500 205 -500 0 3
rlabel polysilicon 208 -500 208 -500 0 4
rlabel polysilicon 212 -494 212 -494 0 1
rlabel polysilicon 212 -500 212 -500 0 3
rlabel polysilicon 219 -494 219 -494 0 1
rlabel polysilicon 219 -500 219 -500 0 3
rlabel polysilicon 226 -494 226 -494 0 1
rlabel polysilicon 226 -500 226 -500 0 3
rlabel polysilicon 233 -494 233 -494 0 1
rlabel polysilicon 236 -500 236 -500 0 4
rlabel polysilicon 243 -494 243 -494 0 2
rlabel polysilicon 240 -500 240 -500 0 3
rlabel polysilicon 247 -494 247 -494 0 1
rlabel polysilicon 247 -500 247 -500 0 3
rlabel polysilicon 254 -494 254 -494 0 1
rlabel polysilicon 254 -500 254 -500 0 3
rlabel polysilicon 264 -494 264 -494 0 2
rlabel polysilicon 268 -494 268 -494 0 1
rlabel polysilicon 268 -500 268 -500 0 3
rlabel polysilicon 275 -494 275 -494 0 1
rlabel polysilicon 275 -500 275 -500 0 3
rlabel polysilicon 282 -494 282 -494 0 1
rlabel polysilicon 282 -500 282 -500 0 3
rlabel polysilicon 289 -494 289 -494 0 1
rlabel polysilicon 289 -500 289 -500 0 3
rlabel polysilicon 296 -494 296 -494 0 1
rlabel polysilicon 296 -500 296 -500 0 3
rlabel polysilicon 303 -494 303 -494 0 1
rlabel polysilicon 303 -500 303 -500 0 3
rlabel polysilicon 306 -500 306 -500 0 4
rlabel polysilicon 310 -494 310 -494 0 1
rlabel polysilicon 313 -494 313 -494 0 2
rlabel polysilicon 310 -500 310 -500 0 3
rlabel polysilicon 313 -500 313 -500 0 4
rlabel polysilicon 317 -494 317 -494 0 1
rlabel polysilicon 317 -500 317 -500 0 3
rlabel polysilicon 324 -494 324 -494 0 1
rlabel polysilicon 327 -494 327 -494 0 2
rlabel polysilicon 324 -500 324 -500 0 3
rlabel polysilicon 331 -494 331 -494 0 1
rlabel polysilicon 334 -494 334 -494 0 2
rlabel polysilicon 331 -500 331 -500 0 3
rlabel polysilicon 334 -500 334 -500 0 4
rlabel polysilicon 338 -494 338 -494 0 1
rlabel polysilicon 338 -500 338 -500 0 3
rlabel polysilicon 345 -494 345 -494 0 1
rlabel polysilicon 345 -500 345 -500 0 3
rlabel polysilicon 352 -494 352 -494 0 1
rlabel polysilicon 355 -494 355 -494 0 2
rlabel polysilicon 355 -500 355 -500 0 4
rlabel polysilicon 362 -494 362 -494 0 2
rlabel polysilicon 362 -500 362 -500 0 4
rlabel polysilicon 366 -494 366 -494 0 1
rlabel polysilicon 366 -500 366 -500 0 3
rlabel polysilicon 373 -494 373 -494 0 1
rlabel polysilicon 373 -500 373 -500 0 3
rlabel polysilicon 380 -494 380 -494 0 1
rlabel polysilicon 380 -500 380 -500 0 3
rlabel polysilicon 387 -494 387 -494 0 1
rlabel polysilicon 387 -500 387 -500 0 3
rlabel polysilicon 394 -494 394 -494 0 1
rlabel polysilicon 397 -494 397 -494 0 2
rlabel polysilicon 397 -500 397 -500 0 4
rlabel polysilicon 401 -494 401 -494 0 1
rlabel polysilicon 401 -500 401 -500 0 3
rlabel polysilicon 408 -494 408 -494 0 1
rlabel polysilicon 408 -500 408 -500 0 3
rlabel polysilicon 415 -494 415 -494 0 1
rlabel polysilicon 415 -500 415 -500 0 3
rlabel polysilicon 422 -494 422 -494 0 1
rlabel polysilicon 425 -500 425 -500 0 4
rlabel polysilicon 429 -494 429 -494 0 1
rlabel polysilicon 429 -500 429 -500 0 3
rlabel polysilicon 436 -494 436 -494 0 1
rlabel polysilicon 436 -500 436 -500 0 3
rlabel polysilicon 443 -494 443 -494 0 1
rlabel polysilicon 443 -500 443 -500 0 3
rlabel polysilicon 450 -494 450 -494 0 1
rlabel polysilicon 450 -500 450 -500 0 3
rlabel polysilicon 457 -494 457 -494 0 1
rlabel polysilicon 457 -500 457 -500 0 3
rlabel polysilicon 464 -494 464 -494 0 1
rlabel polysilicon 464 -500 464 -500 0 3
rlabel polysilicon 471 -494 471 -494 0 1
rlabel polysilicon 471 -500 471 -500 0 3
rlabel polysilicon 478 -494 478 -494 0 1
rlabel polysilicon 478 -500 478 -500 0 3
rlabel polysilicon 485 -494 485 -494 0 1
rlabel polysilicon 485 -500 485 -500 0 3
rlabel polysilicon 492 -500 492 -500 0 3
rlabel polysilicon 495 -500 495 -500 0 4
rlabel polysilicon 499 -494 499 -494 0 1
rlabel polysilicon 499 -500 499 -500 0 3
rlabel polysilicon 506 -494 506 -494 0 1
rlabel polysilicon 506 -500 506 -500 0 3
rlabel polysilicon 513 -494 513 -494 0 1
rlabel polysilicon 513 -500 513 -500 0 3
rlabel polysilicon 520 -494 520 -494 0 1
rlabel polysilicon 520 -500 520 -500 0 3
rlabel polysilicon 527 -494 527 -494 0 1
rlabel polysilicon 527 -500 527 -500 0 3
rlabel polysilicon 534 -494 534 -494 0 1
rlabel polysilicon 534 -500 534 -500 0 3
rlabel polysilicon 541 -494 541 -494 0 1
rlabel polysilicon 541 -500 541 -500 0 3
rlabel polysilicon 548 -494 548 -494 0 1
rlabel polysilicon 548 -500 548 -500 0 3
rlabel polysilicon 555 -494 555 -494 0 1
rlabel polysilicon 555 -500 555 -500 0 3
rlabel polysilicon 562 -494 562 -494 0 1
rlabel polysilicon 562 -500 562 -500 0 3
rlabel polysilicon 569 -494 569 -494 0 1
rlabel polysilicon 569 -500 569 -500 0 3
rlabel polysilicon 576 -494 576 -494 0 1
rlabel polysilicon 576 -500 576 -500 0 3
rlabel polysilicon 583 -494 583 -494 0 1
rlabel polysilicon 583 -500 583 -500 0 3
rlabel polysilicon 590 -494 590 -494 0 1
rlabel polysilicon 590 -500 590 -500 0 3
rlabel polysilicon 597 -494 597 -494 0 1
rlabel polysilicon 597 -500 597 -500 0 3
rlabel polysilicon 604 -494 604 -494 0 1
rlabel polysilicon 604 -500 604 -500 0 3
rlabel polysilicon 611 -494 611 -494 0 1
rlabel polysilicon 611 -500 611 -500 0 3
rlabel polysilicon 621 -494 621 -494 0 2
rlabel polysilicon 618 -500 618 -500 0 3
rlabel polysilicon 621 -500 621 -500 0 4
rlabel polysilicon 625 -494 625 -494 0 1
rlabel polysilicon 625 -500 625 -500 0 3
rlabel polysilicon 635 -494 635 -494 0 2
rlabel polysilicon 632 -500 632 -500 0 3
rlabel polysilicon 635 -500 635 -500 0 4
rlabel polysilicon 639 -494 639 -494 0 1
rlabel polysilicon 639 -500 639 -500 0 3
rlabel polysilicon 646 -494 646 -494 0 1
rlabel polysilicon 646 -500 646 -500 0 3
rlabel polysilicon 653 -500 653 -500 0 3
rlabel polysilicon 663 -494 663 -494 0 2
rlabel polysilicon 667 -494 667 -494 0 1
rlabel polysilicon 667 -500 667 -500 0 3
rlabel polysilicon 674 -494 674 -494 0 1
rlabel polysilicon 674 -500 674 -500 0 3
rlabel polysilicon 16 -559 16 -559 0 1
rlabel polysilicon 16 -565 16 -565 0 3
rlabel polysilicon 23 -559 23 -559 0 1
rlabel polysilicon 23 -565 23 -565 0 3
rlabel polysilicon 30 -559 30 -559 0 1
rlabel polysilicon 30 -565 30 -565 0 3
rlabel polysilicon 37 -559 37 -559 0 1
rlabel polysilicon 37 -565 37 -565 0 3
rlabel polysilicon 44 -565 44 -565 0 3
rlabel polysilicon 51 -559 51 -559 0 1
rlabel polysilicon 51 -565 51 -565 0 3
rlabel polysilicon 61 -559 61 -559 0 2
rlabel polysilicon 58 -565 58 -565 0 3
rlabel polysilicon 65 -559 65 -559 0 1
rlabel polysilicon 65 -565 65 -565 0 3
rlabel polysilicon 75 -559 75 -559 0 2
rlabel polysilicon 72 -565 72 -565 0 3
rlabel polysilicon 79 -565 79 -565 0 3
rlabel polysilicon 82 -565 82 -565 0 4
rlabel polysilicon 86 -559 86 -559 0 1
rlabel polysilicon 86 -565 86 -565 0 3
rlabel polysilicon 93 -559 93 -559 0 1
rlabel polysilicon 93 -565 93 -565 0 3
rlabel polysilicon 100 -559 100 -559 0 1
rlabel polysilicon 100 -565 100 -565 0 3
rlabel polysilicon 107 -559 107 -559 0 1
rlabel polysilicon 107 -565 107 -565 0 3
rlabel polysilicon 114 -559 114 -559 0 1
rlabel polysilicon 114 -565 114 -565 0 3
rlabel polysilicon 121 -559 121 -559 0 1
rlabel polysilicon 121 -565 121 -565 0 3
rlabel polysilicon 131 -559 131 -559 0 2
rlabel polysilicon 135 -559 135 -559 0 1
rlabel polysilicon 135 -565 135 -565 0 3
rlabel polysilicon 145 -559 145 -559 0 2
rlabel polysilicon 142 -565 142 -565 0 3
rlabel polysilicon 149 -559 149 -559 0 1
rlabel polysilicon 152 -559 152 -559 0 2
rlabel polysilicon 149 -565 149 -565 0 3
rlabel polysilicon 152 -565 152 -565 0 4
rlabel polysilicon 156 -559 156 -559 0 1
rlabel polysilicon 156 -565 156 -565 0 3
rlabel polysilicon 163 -559 163 -559 0 1
rlabel polysilicon 163 -565 163 -565 0 3
rlabel polysilicon 170 -559 170 -559 0 1
rlabel polysilicon 173 -559 173 -559 0 2
rlabel polysilicon 170 -565 170 -565 0 3
rlabel polysilicon 177 -559 177 -559 0 1
rlabel polysilicon 177 -565 177 -565 0 3
rlabel polysilicon 184 -559 184 -559 0 1
rlabel polysilicon 184 -565 184 -565 0 3
rlabel polysilicon 191 -559 191 -559 0 1
rlabel polysilicon 191 -565 191 -565 0 3
rlabel polysilicon 194 -565 194 -565 0 4
rlabel polysilicon 198 -559 198 -559 0 1
rlabel polysilicon 198 -565 198 -565 0 3
rlabel polysilicon 205 -559 205 -559 0 1
rlabel polysilicon 208 -559 208 -559 0 2
rlabel polysilicon 205 -565 205 -565 0 3
rlabel polysilicon 212 -559 212 -559 0 1
rlabel polysilicon 212 -565 212 -565 0 3
rlabel polysilicon 219 -559 219 -559 0 1
rlabel polysilicon 219 -565 219 -565 0 3
rlabel polysilicon 226 -559 226 -559 0 1
rlabel polysilicon 226 -565 226 -565 0 3
rlabel polysilicon 233 -559 233 -559 0 1
rlabel polysilicon 233 -565 233 -565 0 3
rlabel polysilicon 240 -559 240 -559 0 1
rlabel polysilicon 240 -565 240 -565 0 3
rlabel polysilicon 247 -559 247 -559 0 1
rlabel polysilicon 247 -565 247 -565 0 3
rlabel polysilicon 254 -559 254 -559 0 1
rlabel polysilicon 254 -565 254 -565 0 3
rlabel polysilicon 264 -559 264 -559 0 2
rlabel polysilicon 261 -565 261 -565 0 3
rlabel polysilicon 264 -565 264 -565 0 4
rlabel polysilicon 268 -559 268 -559 0 1
rlabel polysilicon 271 -559 271 -559 0 2
rlabel polysilicon 268 -565 268 -565 0 3
rlabel polysilicon 271 -565 271 -565 0 4
rlabel polysilicon 275 -559 275 -559 0 1
rlabel polysilicon 278 -559 278 -559 0 2
rlabel polysilicon 282 -559 282 -559 0 1
rlabel polysilicon 282 -565 282 -565 0 3
rlabel polysilicon 289 -559 289 -559 0 1
rlabel polysilicon 289 -565 289 -565 0 3
rlabel polysilicon 296 -559 296 -559 0 1
rlabel polysilicon 296 -565 296 -565 0 3
rlabel polysilicon 303 -559 303 -559 0 1
rlabel polysilicon 303 -565 303 -565 0 3
rlabel polysilicon 310 -559 310 -559 0 1
rlabel polysilicon 310 -565 310 -565 0 3
rlabel polysilicon 317 -559 317 -559 0 1
rlabel polysilicon 317 -565 317 -565 0 3
rlabel polysilicon 324 -559 324 -559 0 1
rlabel polysilicon 324 -565 324 -565 0 3
rlabel polysilicon 334 -559 334 -559 0 2
rlabel polysilicon 334 -565 334 -565 0 4
rlabel polysilicon 338 -559 338 -559 0 1
rlabel polysilicon 338 -565 338 -565 0 3
rlabel polysilicon 348 -559 348 -559 0 2
rlabel polysilicon 348 -565 348 -565 0 4
rlabel polysilicon 352 -559 352 -559 0 1
rlabel polysilicon 352 -565 352 -565 0 3
rlabel polysilicon 355 -565 355 -565 0 4
rlabel polysilicon 359 -559 359 -559 0 1
rlabel polysilicon 359 -565 359 -565 0 3
rlabel polysilicon 366 -559 366 -559 0 1
rlabel polysilicon 369 -559 369 -559 0 2
rlabel polysilicon 369 -565 369 -565 0 4
rlabel polysilicon 373 -559 373 -559 0 1
rlabel polysilicon 373 -565 373 -565 0 3
rlabel polysilicon 380 -559 380 -559 0 1
rlabel polysilicon 383 -559 383 -559 0 2
rlabel polysilicon 383 -565 383 -565 0 4
rlabel polysilicon 390 -559 390 -559 0 2
rlabel polysilicon 387 -565 387 -565 0 3
rlabel polysilicon 394 -559 394 -559 0 1
rlabel polysilicon 397 -559 397 -559 0 2
rlabel polysilicon 394 -565 394 -565 0 3
rlabel polysilicon 401 -565 401 -565 0 3
rlabel polysilicon 404 -565 404 -565 0 4
rlabel polysilicon 411 -559 411 -559 0 2
rlabel polysilicon 408 -565 408 -565 0 3
rlabel polysilicon 411 -565 411 -565 0 4
rlabel polysilicon 415 -559 415 -559 0 1
rlabel polysilicon 415 -565 415 -565 0 3
rlabel polysilicon 422 -559 422 -559 0 1
rlabel polysilicon 422 -565 422 -565 0 3
rlabel polysilicon 429 -559 429 -559 0 1
rlabel polysilicon 429 -565 429 -565 0 3
rlabel polysilicon 436 -559 436 -559 0 1
rlabel polysilicon 436 -565 436 -565 0 3
rlabel polysilicon 443 -559 443 -559 0 1
rlabel polysilicon 443 -565 443 -565 0 3
rlabel polysilicon 450 -559 450 -559 0 1
rlabel polysilicon 450 -565 450 -565 0 3
rlabel polysilicon 457 -559 457 -559 0 1
rlabel polysilicon 457 -565 457 -565 0 3
rlabel polysilicon 464 -559 464 -559 0 1
rlabel polysilicon 464 -565 464 -565 0 3
rlabel polysilicon 471 -559 471 -559 0 1
rlabel polysilicon 471 -565 471 -565 0 3
rlabel polysilicon 478 -559 478 -559 0 1
rlabel polysilicon 478 -565 478 -565 0 3
rlabel polysilicon 485 -559 485 -559 0 1
rlabel polysilicon 485 -565 485 -565 0 3
rlabel polysilicon 492 -559 492 -559 0 1
rlabel polysilicon 492 -565 492 -565 0 3
rlabel polysilicon 499 -559 499 -559 0 1
rlabel polysilicon 499 -565 499 -565 0 3
rlabel polysilicon 506 -559 506 -559 0 1
rlabel polysilicon 506 -565 506 -565 0 3
rlabel polysilicon 513 -559 513 -559 0 1
rlabel polysilicon 513 -565 513 -565 0 3
rlabel polysilicon 520 -559 520 -559 0 1
rlabel polysilicon 520 -565 520 -565 0 3
rlabel polysilicon 527 -559 527 -559 0 1
rlabel polysilicon 527 -565 527 -565 0 3
rlabel polysilicon 534 -559 534 -559 0 1
rlabel polysilicon 534 -565 534 -565 0 3
rlabel polysilicon 541 -559 541 -559 0 1
rlabel polysilicon 541 -565 541 -565 0 3
rlabel polysilicon 548 -559 548 -559 0 1
rlabel polysilicon 548 -565 548 -565 0 3
rlabel polysilicon 555 -559 555 -559 0 1
rlabel polysilicon 555 -565 555 -565 0 3
rlabel polysilicon 562 -559 562 -559 0 1
rlabel polysilicon 562 -565 562 -565 0 3
rlabel polysilicon 569 -559 569 -559 0 1
rlabel polysilicon 569 -565 569 -565 0 3
rlabel polysilicon 576 -559 576 -559 0 1
rlabel polysilicon 576 -565 576 -565 0 3
rlabel polysilicon 583 -559 583 -559 0 1
rlabel polysilicon 583 -565 583 -565 0 3
rlabel polysilicon 590 -559 590 -559 0 1
rlabel polysilicon 590 -565 590 -565 0 3
rlabel polysilicon 597 -559 597 -559 0 1
rlabel polysilicon 597 -565 597 -565 0 3
rlabel polysilicon 604 -559 604 -559 0 1
rlabel polysilicon 604 -565 604 -565 0 3
rlabel polysilicon 611 -559 611 -559 0 1
rlabel polysilicon 614 -559 614 -559 0 2
rlabel polysilicon 618 -559 618 -559 0 1
rlabel polysilicon 618 -565 618 -565 0 3
rlabel polysilicon 621 -565 621 -565 0 4
rlabel polysilicon 625 -559 625 -559 0 1
rlabel polysilicon 628 -559 628 -559 0 2
rlabel polysilicon 628 -565 628 -565 0 4
rlabel polysilicon 632 -559 632 -559 0 1
rlabel polysilicon 632 -565 632 -565 0 3
rlabel polysilicon 639 -559 639 -559 0 1
rlabel polysilicon 642 -559 642 -559 0 2
rlabel polysilicon 642 -565 642 -565 0 4
rlabel polysilicon 646 -559 646 -559 0 1
rlabel polysilicon 646 -565 646 -565 0 3
rlabel polysilicon 653 -559 653 -559 0 1
rlabel polysilicon 653 -565 653 -565 0 3
rlabel polysilicon 2 -614 2 -614 0 1
rlabel polysilicon 2 -620 2 -620 0 3
rlabel polysilicon 9 -614 9 -614 0 1
rlabel polysilicon 9 -620 9 -620 0 3
rlabel polysilicon 16 -614 16 -614 0 1
rlabel polysilicon 16 -620 16 -620 0 3
rlabel polysilicon 23 -614 23 -614 0 1
rlabel polysilicon 23 -620 23 -620 0 3
rlabel polysilicon 30 -614 30 -614 0 1
rlabel polysilicon 30 -620 30 -620 0 3
rlabel polysilicon 37 -614 37 -614 0 1
rlabel polysilicon 37 -620 37 -620 0 3
rlabel polysilicon 44 -614 44 -614 0 1
rlabel polysilicon 44 -620 44 -620 0 3
rlabel polysilicon 51 -614 51 -614 0 1
rlabel polysilicon 51 -620 51 -620 0 3
rlabel polysilicon 61 -614 61 -614 0 2
rlabel polysilicon 61 -620 61 -620 0 4
rlabel polysilicon 68 -614 68 -614 0 2
rlabel polysilicon 65 -620 65 -620 0 3
rlabel polysilicon 68 -620 68 -620 0 4
rlabel polysilicon 72 -614 72 -614 0 1
rlabel polysilicon 72 -620 72 -620 0 3
rlabel polysilicon 79 -614 79 -614 0 1
rlabel polysilicon 79 -620 79 -620 0 3
rlabel polysilicon 86 -614 86 -614 0 1
rlabel polysilicon 86 -620 86 -620 0 3
rlabel polysilicon 93 -614 93 -614 0 1
rlabel polysilicon 93 -620 93 -620 0 3
rlabel polysilicon 100 -614 100 -614 0 1
rlabel polysilicon 103 -614 103 -614 0 2
rlabel polysilicon 103 -620 103 -620 0 4
rlabel polysilicon 107 -614 107 -614 0 1
rlabel polysilicon 107 -620 107 -620 0 3
rlabel polysilicon 114 -614 114 -614 0 1
rlabel polysilicon 114 -620 114 -620 0 3
rlabel polysilicon 121 -614 121 -614 0 1
rlabel polysilicon 124 -614 124 -614 0 2
rlabel polysilicon 121 -620 121 -620 0 3
rlabel polysilicon 128 -614 128 -614 0 1
rlabel polysilicon 128 -620 128 -620 0 3
rlabel polysilicon 131 -620 131 -620 0 4
rlabel polysilicon 135 -614 135 -614 0 1
rlabel polysilicon 135 -620 135 -620 0 3
rlabel polysilicon 142 -614 142 -614 0 1
rlabel polysilicon 142 -620 142 -620 0 3
rlabel polysilicon 152 -614 152 -614 0 2
rlabel polysilicon 152 -620 152 -620 0 4
rlabel polysilicon 156 -614 156 -614 0 1
rlabel polysilicon 156 -620 156 -620 0 3
rlabel polysilicon 163 -614 163 -614 0 1
rlabel polysilicon 163 -620 163 -620 0 3
rlabel polysilicon 170 -614 170 -614 0 1
rlabel polysilicon 170 -620 170 -620 0 3
rlabel polysilicon 177 -614 177 -614 0 1
rlabel polysilicon 180 -614 180 -614 0 2
rlabel polysilicon 177 -620 177 -620 0 3
rlabel polysilicon 180 -620 180 -620 0 4
rlabel polysilicon 184 -614 184 -614 0 1
rlabel polysilicon 184 -620 184 -620 0 3
rlabel polysilicon 191 -614 191 -614 0 1
rlabel polysilicon 194 -620 194 -620 0 4
rlabel polysilicon 198 -614 198 -614 0 1
rlabel polysilicon 201 -614 201 -614 0 2
rlabel polysilicon 198 -620 198 -620 0 3
rlabel polysilicon 201 -620 201 -620 0 4
rlabel polysilicon 205 -614 205 -614 0 1
rlabel polysilicon 208 -614 208 -614 0 2
rlabel polysilicon 205 -620 205 -620 0 3
rlabel polysilicon 208 -620 208 -620 0 4
rlabel polysilicon 212 -614 212 -614 0 1
rlabel polysilicon 212 -620 212 -620 0 3
rlabel polysilicon 219 -614 219 -614 0 1
rlabel polysilicon 219 -620 219 -620 0 3
rlabel polysilicon 226 -614 226 -614 0 1
rlabel polysilicon 229 -614 229 -614 0 2
rlabel polysilicon 226 -620 226 -620 0 3
rlabel polysilicon 229 -620 229 -620 0 4
rlabel polysilicon 233 -614 233 -614 0 1
rlabel polysilicon 233 -620 233 -620 0 3
rlabel polysilicon 240 -614 240 -614 0 1
rlabel polysilicon 240 -620 240 -620 0 3
rlabel polysilicon 247 -614 247 -614 0 1
rlabel polysilicon 247 -620 247 -620 0 3
rlabel polysilicon 257 -614 257 -614 0 2
rlabel polysilicon 257 -620 257 -620 0 4
rlabel polysilicon 261 -614 261 -614 0 1
rlabel polysilicon 261 -620 261 -620 0 3
rlabel polysilicon 268 -614 268 -614 0 1
rlabel polysilicon 268 -620 268 -620 0 3
rlabel polysilicon 278 -614 278 -614 0 2
rlabel polysilicon 278 -620 278 -620 0 4
rlabel polysilicon 282 -614 282 -614 0 1
rlabel polysilicon 282 -620 282 -620 0 3
rlabel polysilicon 289 -614 289 -614 0 1
rlabel polysilicon 289 -620 289 -620 0 3
rlabel polysilicon 296 -614 296 -614 0 1
rlabel polysilicon 296 -620 296 -620 0 3
rlabel polysilicon 303 -614 303 -614 0 1
rlabel polysilicon 303 -620 303 -620 0 3
rlabel polysilicon 310 -614 310 -614 0 1
rlabel polysilicon 310 -620 310 -620 0 3
rlabel polysilicon 313 -620 313 -620 0 4
rlabel polysilicon 317 -614 317 -614 0 1
rlabel polysilicon 317 -620 317 -620 0 3
rlabel polysilicon 324 -614 324 -614 0 1
rlabel polysilicon 324 -620 324 -620 0 3
rlabel polysilicon 327 -620 327 -620 0 4
rlabel polysilicon 331 -614 331 -614 0 1
rlabel polysilicon 334 -620 334 -620 0 4
rlabel polysilicon 338 -614 338 -614 0 1
rlabel polysilicon 338 -620 338 -620 0 3
rlabel polysilicon 345 -614 345 -614 0 1
rlabel polysilicon 348 -614 348 -614 0 2
rlabel polysilicon 345 -620 345 -620 0 3
rlabel polysilicon 348 -620 348 -620 0 4
rlabel polysilicon 352 -614 352 -614 0 1
rlabel polysilicon 355 -620 355 -620 0 4
rlabel polysilicon 359 -614 359 -614 0 1
rlabel polysilicon 362 -614 362 -614 0 2
rlabel polysilicon 362 -620 362 -620 0 4
rlabel polysilicon 366 -614 366 -614 0 1
rlabel polysilicon 366 -620 366 -620 0 3
rlabel polysilicon 373 -614 373 -614 0 1
rlabel polysilicon 373 -620 373 -620 0 3
rlabel polysilicon 380 -614 380 -614 0 1
rlabel polysilicon 380 -620 380 -620 0 3
rlabel polysilicon 387 -614 387 -614 0 1
rlabel polysilicon 387 -620 387 -620 0 3
rlabel polysilicon 394 -614 394 -614 0 1
rlabel polysilicon 394 -620 394 -620 0 3
rlabel polysilicon 401 -614 401 -614 0 1
rlabel polysilicon 404 -620 404 -620 0 4
rlabel polysilicon 408 -614 408 -614 0 1
rlabel polysilicon 408 -620 408 -620 0 3
rlabel polysilicon 415 -614 415 -614 0 1
rlabel polysilicon 415 -620 415 -620 0 3
rlabel polysilicon 422 -614 422 -614 0 1
rlabel polysilicon 422 -620 422 -620 0 3
rlabel polysilicon 429 -614 429 -614 0 1
rlabel polysilicon 429 -620 429 -620 0 3
rlabel polysilicon 436 -614 436 -614 0 1
rlabel polysilicon 436 -620 436 -620 0 3
rlabel polysilicon 443 -614 443 -614 0 1
rlabel polysilicon 443 -620 443 -620 0 3
rlabel polysilicon 450 -614 450 -614 0 1
rlabel polysilicon 450 -620 450 -620 0 3
rlabel polysilicon 457 -620 457 -620 0 3
rlabel polysilicon 460 -620 460 -620 0 4
rlabel polysilicon 464 -614 464 -614 0 1
rlabel polysilicon 464 -620 464 -620 0 3
rlabel polysilicon 471 -614 471 -614 0 1
rlabel polysilicon 471 -620 471 -620 0 3
rlabel polysilicon 478 -614 478 -614 0 1
rlabel polysilicon 485 -614 485 -614 0 1
rlabel polysilicon 485 -620 485 -620 0 3
rlabel polysilicon 492 -614 492 -614 0 1
rlabel polysilicon 492 -620 492 -620 0 3
rlabel polysilicon 499 -614 499 -614 0 1
rlabel polysilicon 499 -620 499 -620 0 3
rlabel polysilicon 506 -614 506 -614 0 1
rlabel polysilicon 506 -620 506 -620 0 3
rlabel polysilicon 513 -614 513 -614 0 1
rlabel polysilicon 513 -620 513 -620 0 3
rlabel polysilicon 520 -614 520 -614 0 1
rlabel polysilicon 520 -620 520 -620 0 3
rlabel polysilicon 527 -620 527 -620 0 3
rlabel polysilicon 534 -614 534 -614 0 1
rlabel polysilicon 534 -620 534 -620 0 3
rlabel polysilicon 544 -614 544 -614 0 2
rlabel polysilicon 548 -614 548 -614 0 1
rlabel polysilicon 548 -620 548 -620 0 3
rlabel polysilicon 555 -614 555 -614 0 1
rlabel polysilicon 555 -620 555 -620 0 3
rlabel polysilicon 565 -614 565 -614 0 2
rlabel polysilicon 569 -614 569 -614 0 1
rlabel polysilicon 569 -620 569 -620 0 3
rlabel polysilicon 576 -614 576 -614 0 1
rlabel polysilicon 576 -620 576 -620 0 3
rlabel polysilicon 583 -614 583 -614 0 1
rlabel polysilicon 583 -620 583 -620 0 3
rlabel polysilicon 590 -614 590 -614 0 1
rlabel polysilicon 590 -620 590 -620 0 3
rlabel polysilicon 597 -614 597 -614 0 1
rlabel polysilicon 597 -620 597 -620 0 3
rlabel polysilicon 604 -614 604 -614 0 1
rlabel polysilicon 604 -620 604 -620 0 3
rlabel polysilicon 611 -614 611 -614 0 1
rlabel polysilicon 611 -620 611 -620 0 3
rlabel polysilicon 618 -614 618 -614 0 1
rlabel polysilicon 618 -620 618 -620 0 3
rlabel polysilicon 625 -614 625 -614 0 1
rlabel polysilicon 625 -620 625 -620 0 3
rlabel polysilicon 632 -614 632 -614 0 1
rlabel polysilicon 632 -620 632 -620 0 3
rlabel polysilicon 653 -614 653 -614 0 1
rlabel polysilicon 653 -620 653 -620 0 3
rlabel polysilicon 2 -679 2 -679 0 1
rlabel polysilicon 2 -685 2 -685 0 3
rlabel polysilicon 9 -679 9 -679 0 1
rlabel polysilicon 9 -685 9 -685 0 3
rlabel polysilicon 16 -679 16 -679 0 1
rlabel polysilicon 16 -685 16 -685 0 3
rlabel polysilicon 23 -679 23 -679 0 1
rlabel polysilicon 30 -679 30 -679 0 1
rlabel polysilicon 30 -685 30 -685 0 3
rlabel polysilicon 37 -679 37 -679 0 1
rlabel polysilicon 37 -685 37 -685 0 3
rlabel polysilicon 44 -679 44 -679 0 1
rlabel polysilicon 44 -685 44 -685 0 3
rlabel polysilicon 51 -679 51 -679 0 1
rlabel polysilicon 54 -685 54 -685 0 4
rlabel polysilicon 58 -679 58 -679 0 1
rlabel polysilicon 58 -685 58 -685 0 3
rlabel polysilicon 65 -679 65 -679 0 1
rlabel polysilicon 65 -685 65 -685 0 3
rlabel polysilicon 72 -679 72 -679 0 1
rlabel polysilicon 72 -685 72 -685 0 3
rlabel polysilicon 79 -679 79 -679 0 1
rlabel polysilicon 79 -685 79 -685 0 3
rlabel polysilicon 86 -679 86 -679 0 1
rlabel polysilicon 86 -685 86 -685 0 3
rlabel polysilicon 96 -679 96 -679 0 2
rlabel polysilicon 96 -685 96 -685 0 4
rlabel polysilicon 100 -679 100 -679 0 1
rlabel polysilicon 100 -685 100 -685 0 3
rlabel polysilicon 107 -679 107 -679 0 1
rlabel polysilicon 107 -685 107 -685 0 3
rlabel polysilicon 114 -685 114 -685 0 3
rlabel polysilicon 117 -685 117 -685 0 4
rlabel polysilicon 121 -679 121 -679 0 1
rlabel polysilicon 121 -685 121 -685 0 3
rlabel polysilicon 128 -679 128 -679 0 1
rlabel polysilicon 131 -679 131 -679 0 2
rlabel polysilicon 128 -685 128 -685 0 3
rlabel polysilicon 135 -679 135 -679 0 1
rlabel polysilicon 138 -679 138 -679 0 2
rlabel polysilicon 142 -679 142 -679 0 1
rlabel polysilicon 142 -685 142 -685 0 3
rlabel polysilicon 149 -679 149 -679 0 1
rlabel polysilicon 152 -679 152 -679 0 2
rlabel polysilicon 149 -685 149 -685 0 3
rlabel polysilicon 156 -679 156 -679 0 1
rlabel polysilicon 156 -685 156 -685 0 3
rlabel polysilicon 163 -679 163 -679 0 1
rlabel polysilicon 163 -685 163 -685 0 3
rlabel polysilicon 170 -679 170 -679 0 1
rlabel polysilicon 173 -679 173 -679 0 2
rlabel polysilicon 173 -685 173 -685 0 4
rlabel polysilicon 177 -679 177 -679 0 1
rlabel polysilicon 177 -685 177 -685 0 3
rlabel polysilicon 180 -685 180 -685 0 4
rlabel polysilicon 184 -679 184 -679 0 1
rlabel polysilicon 187 -685 187 -685 0 4
rlabel polysilicon 191 -679 191 -679 0 1
rlabel polysilicon 191 -685 191 -685 0 3
rlabel polysilicon 201 -679 201 -679 0 2
rlabel polysilicon 198 -685 198 -685 0 3
rlabel polysilicon 201 -685 201 -685 0 4
rlabel polysilicon 205 -679 205 -679 0 1
rlabel polysilicon 208 -679 208 -679 0 2
rlabel polysilicon 205 -685 205 -685 0 3
rlabel polysilicon 212 -679 212 -679 0 1
rlabel polysilicon 212 -685 212 -685 0 3
rlabel polysilicon 219 -679 219 -679 0 1
rlabel polysilicon 222 -679 222 -679 0 2
rlabel polysilicon 219 -685 219 -685 0 3
rlabel polysilicon 226 -679 226 -679 0 1
rlabel polysilicon 226 -685 226 -685 0 3
rlabel polysilicon 233 -679 233 -679 0 1
rlabel polysilicon 233 -685 233 -685 0 3
rlabel polysilicon 240 -679 240 -679 0 1
rlabel polysilicon 240 -685 240 -685 0 3
rlabel polysilicon 247 -679 247 -679 0 1
rlabel polysilicon 247 -685 247 -685 0 3
rlabel polysilicon 257 -679 257 -679 0 2
rlabel polysilicon 254 -685 254 -685 0 3
rlabel polysilicon 257 -685 257 -685 0 4
rlabel polysilicon 261 -679 261 -679 0 1
rlabel polysilicon 261 -685 261 -685 0 3
rlabel polysilicon 268 -679 268 -679 0 1
rlabel polysilicon 268 -685 268 -685 0 3
rlabel polysilicon 275 -679 275 -679 0 1
rlabel polysilicon 278 -679 278 -679 0 2
rlabel polysilicon 275 -685 275 -685 0 3
rlabel polysilicon 278 -685 278 -685 0 4
rlabel polysilicon 285 -685 285 -685 0 4
rlabel polysilicon 289 -679 289 -679 0 1
rlabel polysilicon 292 -685 292 -685 0 4
rlabel polysilicon 296 -679 296 -679 0 1
rlabel polysilicon 296 -685 296 -685 0 3
rlabel polysilicon 303 -679 303 -679 0 1
rlabel polysilicon 303 -685 303 -685 0 3
rlabel polysilicon 310 -679 310 -679 0 1
rlabel polysilicon 313 -679 313 -679 0 2
rlabel polysilicon 310 -685 310 -685 0 3
rlabel polysilicon 313 -685 313 -685 0 4
rlabel polysilicon 317 -679 317 -679 0 1
rlabel polysilicon 317 -685 317 -685 0 3
rlabel polysilicon 324 -679 324 -679 0 1
rlabel polysilicon 324 -685 324 -685 0 3
rlabel polysilicon 331 -679 331 -679 0 1
rlabel polysilicon 334 -679 334 -679 0 2
rlabel polysilicon 331 -685 331 -685 0 3
rlabel polysilicon 338 -679 338 -679 0 1
rlabel polysilicon 338 -685 338 -685 0 3
rlabel polysilicon 345 -679 345 -679 0 1
rlabel polysilicon 345 -685 345 -685 0 3
rlabel polysilicon 352 -679 352 -679 0 1
rlabel polysilicon 352 -685 352 -685 0 3
rlabel polysilicon 359 -679 359 -679 0 1
rlabel polysilicon 359 -685 359 -685 0 3
rlabel polysilicon 369 -679 369 -679 0 2
rlabel polysilicon 366 -685 366 -685 0 3
rlabel polysilicon 369 -685 369 -685 0 4
rlabel polysilicon 373 -679 373 -679 0 1
rlabel polysilicon 376 -685 376 -685 0 4
rlabel polysilicon 380 -679 380 -679 0 1
rlabel polysilicon 380 -685 380 -685 0 3
rlabel polysilicon 387 -679 387 -679 0 1
rlabel polysilicon 387 -685 387 -685 0 3
rlabel polysilicon 394 -679 394 -679 0 1
rlabel polysilicon 397 -679 397 -679 0 2
rlabel polysilicon 397 -685 397 -685 0 4
rlabel polysilicon 401 -679 401 -679 0 1
rlabel polysilicon 404 -679 404 -679 0 2
rlabel polysilicon 404 -685 404 -685 0 4
rlabel polysilicon 408 -679 408 -679 0 1
rlabel polysilicon 408 -685 408 -685 0 3
rlabel polysilicon 415 -679 415 -679 0 1
rlabel polysilicon 415 -685 415 -685 0 3
rlabel polysilicon 422 -679 422 -679 0 1
rlabel polysilicon 425 -685 425 -685 0 4
rlabel polysilicon 429 -679 429 -679 0 1
rlabel polysilicon 432 -685 432 -685 0 4
rlabel polysilicon 436 -679 436 -679 0 1
rlabel polysilicon 436 -685 436 -685 0 3
rlabel polysilicon 443 -679 443 -679 0 1
rlabel polysilicon 443 -685 443 -685 0 3
rlabel polysilicon 450 -679 450 -679 0 1
rlabel polysilicon 450 -685 450 -685 0 3
rlabel polysilicon 457 -679 457 -679 0 1
rlabel polysilicon 457 -685 457 -685 0 3
rlabel polysilicon 464 -679 464 -679 0 1
rlabel polysilicon 464 -685 464 -685 0 3
rlabel polysilicon 471 -679 471 -679 0 1
rlabel polysilicon 471 -685 471 -685 0 3
rlabel polysilicon 478 -679 478 -679 0 1
rlabel polysilicon 478 -685 478 -685 0 3
rlabel polysilicon 485 -679 485 -679 0 1
rlabel polysilicon 485 -685 485 -685 0 3
rlabel polysilicon 492 -679 492 -679 0 1
rlabel polysilicon 492 -685 492 -685 0 3
rlabel polysilicon 499 -679 499 -679 0 1
rlabel polysilicon 499 -685 499 -685 0 3
rlabel polysilicon 506 -679 506 -679 0 1
rlabel polysilicon 506 -685 506 -685 0 3
rlabel polysilicon 513 -679 513 -679 0 1
rlabel polysilicon 513 -685 513 -685 0 3
rlabel polysilicon 520 -679 520 -679 0 1
rlabel polysilicon 520 -685 520 -685 0 3
rlabel polysilicon 527 -679 527 -679 0 1
rlabel polysilicon 527 -685 527 -685 0 3
rlabel polysilicon 534 -679 534 -679 0 1
rlabel polysilicon 534 -685 534 -685 0 3
rlabel polysilicon 541 -679 541 -679 0 1
rlabel polysilicon 541 -685 541 -685 0 3
rlabel polysilicon 548 -679 548 -679 0 1
rlabel polysilicon 548 -685 548 -685 0 3
rlabel polysilicon 555 -679 555 -679 0 1
rlabel polysilicon 558 -679 558 -679 0 2
rlabel polysilicon 562 -679 562 -679 0 1
rlabel polysilicon 565 -679 565 -679 0 2
rlabel polysilicon 562 -685 562 -685 0 3
rlabel polysilicon 632 -679 632 -679 0 1
rlabel polysilicon 632 -685 632 -685 0 3
rlabel polysilicon 639 -679 639 -679 0 1
rlabel polysilicon 639 -685 639 -685 0 3
rlabel polysilicon 653 -679 653 -679 0 1
rlabel polysilicon 653 -685 653 -685 0 3
rlabel polysilicon 2 -746 2 -746 0 1
rlabel polysilicon 2 -752 2 -752 0 3
rlabel polysilicon 12 -746 12 -746 0 2
rlabel polysilicon 16 -746 16 -746 0 1
rlabel polysilicon 23 -752 23 -752 0 3
rlabel polysilicon 30 -746 30 -746 0 1
rlabel polysilicon 30 -752 30 -752 0 3
rlabel polysilicon 37 -746 37 -746 0 1
rlabel polysilicon 37 -752 37 -752 0 3
rlabel polysilicon 47 -746 47 -746 0 2
rlabel polysilicon 51 -746 51 -746 0 1
rlabel polysilicon 51 -752 51 -752 0 3
rlabel polysilicon 58 -752 58 -752 0 3
rlabel polysilicon 61 -752 61 -752 0 4
rlabel polysilicon 65 -746 65 -746 0 1
rlabel polysilicon 65 -752 65 -752 0 3
rlabel polysilicon 72 -746 72 -746 0 1
rlabel polysilicon 72 -752 72 -752 0 3
rlabel polysilicon 82 -746 82 -746 0 2
rlabel polysilicon 82 -752 82 -752 0 4
rlabel polysilicon 86 -746 86 -746 0 1
rlabel polysilicon 86 -752 86 -752 0 3
rlabel polysilicon 93 -746 93 -746 0 1
rlabel polysilicon 93 -752 93 -752 0 3
rlabel polysilicon 100 -752 100 -752 0 3
rlabel polysilicon 103 -752 103 -752 0 4
rlabel polysilicon 107 -746 107 -746 0 1
rlabel polysilicon 107 -752 107 -752 0 3
rlabel polysilicon 114 -746 114 -746 0 1
rlabel polysilicon 117 -746 117 -746 0 2
rlabel polysilicon 114 -752 114 -752 0 3
rlabel polysilicon 117 -752 117 -752 0 4
rlabel polysilicon 121 -746 121 -746 0 1
rlabel polysilicon 121 -752 121 -752 0 3
rlabel polysilicon 128 -746 128 -746 0 1
rlabel polysilicon 128 -752 128 -752 0 3
rlabel polysilicon 135 -746 135 -746 0 1
rlabel polysilicon 135 -752 135 -752 0 3
rlabel polysilicon 145 -746 145 -746 0 2
rlabel polysilicon 142 -752 142 -752 0 3
rlabel polysilicon 145 -752 145 -752 0 4
rlabel polysilicon 149 -746 149 -746 0 1
rlabel polysilicon 149 -752 149 -752 0 3
rlabel polysilicon 152 -752 152 -752 0 4
rlabel polysilicon 156 -746 156 -746 0 1
rlabel polysilicon 156 -752 156 -752 0 3
rlabel polysilicon 166 -746 166 -746 0 2
rlabel polysilicon 163 -752 163 -752 0 3
rlabel polysilicon 170 -746 170 -746 0 1
rlabel polysilicon 170 -752 170 -752 0 3
rlabel polysilicon 177 -746 177 -746 0 1
rlabel polysilicon 177 -752 177 -752 0 3
rlabel polysilicon 184 -746 184 -746 0 1
rlabel polysilicon 187 -746 187 -746 0 2
rlabel polysilicon 187 -752 187 -752 0 4
rlabel polysilicon 191 -746 191 -746 0 1
rlabel polysilicon 194 -746 194 -746 0 2
rlabel polysilicon 198 -746 198 -746 0 1
rlabel polysilicon 198 -752 198 -752 0 3
rlabel polysilicon 205 -752 205 -752 0 3
rlabel polysilicon 208 -752 208 -752 0 4
rlabel polysilicon 212 -746 212 -746 0 1
rlabel polysilicon 212 -752 212 -752 0 3
rlabel polysilicon 219 -746 219 -746 0 1
rlabel polysilicon 219 -752 219 -752 0 3
rlabel polysilicon 226 -746 226 -746 0 1
rlabel polysilicon 229 -746 229 -746 0 2
rlabel polysilicon 229 -752 229 -752 0 4
rlabel polysilicon 233 -746 233 -746 0 1
rlabel polysilicon 233 -752 233 -752 0 3
rlabel polysilicon 240 -746 240 -746 0 1
rlabel polysilicon 240 -752 240 -752 0 3
rlabel polysilicon 247 -746 247 -746 0 1
rlabel polysilicon 247 -752 247 -752 0 3
rlabel polysilicon 254 -746 254 -746 0 1
rlabel polysilicon 254 -752 254 -752 0 3
rlabel polysilicon 261 -746 261 -746 0 1
rlabel polysilicon 261 -752 261 -752 0 3
rlabel polysilicon 268 -746 268 -746 0 1
rlabel polysilicon 271 -746 271 -746 0 2
rlabel polysilicon 268 -752 268 -752 0 3
rlabel polysilicon 275 -746 275 -746 0 1
rlabel polysilicon 278 -746 278 -746 0 2
rlabel polysilicon 275 -752 275 -752 0 3
rlabel polysilicon 278 -752 278 -752 0 4
rlabel polysilicon 282 -746 282 -746 0 1
rlabel polysilicon 285 -746 285 -746 0 2
rlabel polysilicon 289 -746 289 -746 0 1
rlabel polysilicon 289 -752 289 -752 0 3
rlabel polysilicon 296 -746 296 -746 0 1
rlabel polysilicon 296 -752 296 -752 0 3
rlabel polysilicon 306 -746 306 -746 0 2
rlabel polysilicon 310 -746 310 -746 0 1
rlabel polysilicon 310 -752 310 -752 0 3
rlabel polysilicon 317 -746 317 -746 0 1
rlabel polysilicon 317 -752 317 -752 0 3
rlabel polysilicon 324 -746 324 -746 0 1
rlabel polysilicon 324 -752 324 -752 0 3
rlabel polysilicon 331 -746 331 -746 0 1
rlabel polysilicon 331 -752 331 -752 0 3
rlabel polysilicon 338 -746 338 -746 0 1
rlabel polysilicon 341 -746 341 -746 0 2
rlabel polysilicon 341 -752 341 -752 0 4
rlabel polysilicon 345 -746 345 -746 0 1
rlabel polysilicon 345 -752 345 -752 0 3
rlabel polysilicon 352 -746 352 -746 0 1
rlabel polysilicon 355 -746 355 -746 0 2
rlabel polysilicon 359 -746 359 -746 0 1
rlabel polysilicon 362 -746 362 -746 0 2
rlabel polysilicon 359 -752 359 -752 0 3
rlabel polysilicon 362 -752 362 -752 0 4
rlabel polysilicon 366 -746 366 -746 0 1
rlabel polysilicon 366 -752 366 -752 0 3
rlabel polysilicon 373 -746 373 -746 0 1
rlabel polysilicon 376 -746 376 -746 0 2
rlabel polysilicon 373 -752 373 -752 0 3
rlabel polysilicon 376 -752 376 -752 0 4
rlabel polysilicon 380 -752 380 -752 0 3
rlabel polysilicon 387 -746 387 -746 0 1
rlabel polysilicon 387 -752 387 -752 0 3
rlabel polysilicon 394 -746 394 -746 0 1
rlabel polysilicon 394 -752 394 -752 0 3
rlabel polysilicon 401 -746 401 -746 0 1
rlabel polysilicon 401 -752 401 -752 0 3
rlabel polysilicon 408 -752 408 -752 0 3
rlabel polysilicon 411 -752 411 -752 0 4
rlabel polysilicon 415 -746 415 -746 0 1
rlabel polysilicon 415 -752 415 -752 0 3
rlabel polysilicon 422 -746 422 -746 0 1
rlabel polysilicon 422 -752 422 -752 0 3
rlabel polysilicon 429 -746 429 -746 0 1
rlabel polysilicon 429 -752 429 -752 0 3
rlabel polysilicon 436 -746 436 -746 0 1
rlabel polysilicon 436 -752 436 -752 0 3
rlabel polysilicon 443 -746 443 -746 0 1
rlabel polysilicon 443 -752 443 -752 0 3
rlabel polysilicon 450 -746 450 -746 0 1
rlabel polysilicon 450 -752 450 -752 0 3
rlabel polysilicon 457 -746 457 -746 0 1
rlabel polysilicon 457 -752 457 -752 0 3
rlabel polysilicon 464 -746 464 -746 0 1
rlabel polysilicon 464 -752 464 -752 0 3
rlabel polysilicon 471 -752 471 -752 0 3
rlabel polysilicon 474 -752 474 -752 0 4
rlabel polysilicon 478 -746 478 -746 0 1
rlabel polysilicon 478 -752 478 -752 0 3
rlabel polysilicon 485 -746 485 -746 0 1
rlabel polysilicon 485 -752 485 -752 0 3
rlabel polysilicon 492 -746 492 -746 0 1
rlabel polysilicon 492 -752 492 -752 0 3
rlabel polysilicon 499 -746 499 -746 0 1
rlabel polysilicon 499 -752 499 -752 0 3
rlabel polysilicon 506 -746 506 -746 0 1
rlabel polysilicon 506 -752 506 -752 0 3
rlabel polysilicon 513 -746 513 -746 0 1
rlabel polysilicon 513 -752 513 -752 0 3
rlabel polysilicon 520 -746 520 -746 0 1
rlabel polysilicon 520 -752 520 -752 0 3
rlabel polysilicon 527 -746 527 -746 0 1
rlabel polysilicon 527 -752 527 -752 0 3
rlabel polysilicon 534 -746 534 -746 0 1
rlabel polysilicon 534 -752 534 -752 0 3
rlabel polysilicon 541 -746 541 -746 0 1
rlabel polysilicon 541 -752 541 -752 0 3
rlabel polysilicon 548 -746 548 -746 0 1
rlabel polysilicon 548 -752 548 -752 0 3
rlabel polysilicon 555 -746 555 -746 0 1
rlabel polysilicon 555 -752 555 -752 0 3
rlabel polysilicon 562 -746 562 -746 0 1
rlabel polysilicon 562 -752 562 -752 0 3
rlabel polysilicon 569 -746 569 -746 0 1
rlabel polysilicon 569 -752 569 -752 0 3
rlabel polysilicon 576 -746 576 -746 0 1
rlabel polysilicon 576 -752 576 -752 0 3
rlabel polysilicon 583 -746 583 -746 0 1
rlabel polysilicon 583 -752 583 -752 0 3
rlabel polysilicon 590 -746 590 -746 0 1
rlabel polysilicon 590 -752 590 -752 0 3
rlabel polysilicon 597 -746 597 -746 0 1
rlabel polysilicon 597 -752 597 -752 0 3
rlabel polysilicon 604 -746 604 -746 0 1
rlabel polysilicon 604 -752 604 -752 0 3
rlabel polysilicon 611 -746 611 -746 0 1
rlabel polysilicon 611 -752 611 -752 0 3
rlabel polysilicon 618 -746 618 -746 0 1
rlabel polysilicon 618 -752 618 -752 0 3
rlabel polysilicon 625 -746 625 -746 0 1
rlabel polysilicon 625 -752 625 -752 0 3
rlabel polysilicon 632 -746 632 -746 0 1
rlabel polysilicon 632 -752 632 -752 0 3
rlabel polysilicon 639 -746 639 -746 0 1
rlabel polysilicon 639 -752 639 -752 0 3
rlabel polysilicon 646 -746 646 -746 0 1
rlabel polysilicon 646 -752 646 -752 0 3
rlabel polysilicon 653 -746 653 -746 0 1
rlabel polysilicon 656 -746 656 -746 0 2
rlabel polysilicon 653 -752 653 -752 0 3
rlabel polysilicon 663 -746 663 -746 0 2
rlabel polysilicon 660 -752 660 -752 0 3
rlabel polysilicon 23 -819 23 -819 0 1
rlabel polysilicon 23 -825 23 -825 0 3
rlabel polysilicon 30 -819 30 -819 0 1
rlabel polysilicon 30 -825 30 -825 0 3
rlabel polysilicon 40 -825 40 -825 0 4
rlabel polysilicon 44 -819 44 -819 0 1
rlabel polysilicon 44 -825 44 -825 0 3
rlabel polysilicon 54 -819 54 -819 0 2
rlabel polysilicon 51 -825 51 -825 0 3
rlabel polysilicon 54 -825 54 -825 0 4
rlabel polysilicon 58 -819 58 -819 0 1
rlabel polysilicon 58 -825 58 -825 0 3
rlabel polysilicon 65 -819 65 -819 0 1
rlabel polysilicon 65 -825 65 -825 0 3
rlabel polysilicon 72 -819 72 -819 0 1
rlabel polysilicon 72 -825 72 -825 0 3
rlabel polysilicon 79 -819 79 -819 0 1
rlabel polysilicon 82 -819 82 -819 0 2
rlabel polysilicon 82 -825 82 -825 0 4
rlabel polysilicon 86 -825 86 -825 0 3
rlabel polysilicon 89 -825 89 -825 0 4
rlabel polysilicon 96 -819 96 -819 0 2
rlabel polysilicon 93 -825 93 -825 0 3
rlabel polysilicon 96 -825 96 -825 0 4
rlabel polysilicon 100 -819 100 -819 0 1
rlabel polysilicon 100 -825 100 -825 0 3
rlabel polysilicon 107 -819 107 -819 0 1
rlabel polysilicon 107 -825 107 -825 0 3
rlabel polysilicon 114 -819 114 -819 0 1
rlabel polysilicon 114 -825 114 -825 0 3
rlabel polysilicon 121 -819 121 -819 0 1
rlabel polysilicon 121 -825 121 -825 0 3
rlabel polysilicon 128 -825 128 -825 0 3
rlabel polysilicon 135 -825 135 -825 0 3
rlabel polysilicon 145 -825 145 -825 0 4
rlabel polysilicon 149 -819 149 -819 0 1
rlabel polysilicon 152 -819 152 -819 0 2
rlabel polysilicon 152 -825 152 -825 0 4
rlabel polysilicon 156 -819 156 -819 0 1
rlabel polysilicon 156 -825 156 -825 0 3
rlabel polysilicon 163 -819 163 -819 0 1
rlabel polysilicon 163 -825 163 -825 0 3
rlabel polysilicon 170 -819 170 -819 0 1
rlabel polysilicon 170 -825 170 -825 0 3
rlabel polysilicon 177 -819 177 -819 0 1
rlabel polysilicon 177 -825 177 -825 0 3
rlabel polysilicon 184 -819 184 -819 0 1
rlabel polysilicon 184 -825 184 -825 0 3
rlabel polysilicon 191 -819 191 -819 0 1
rlabel polysilicon 191 -825 191 -825 0 3
rlabel polysilicon 198 -819 198 -819 0 1
rlabel polysilicon 198 -825 198 -825 0 3
rlabel polysilicon 205 -819 205 -819 0 1
rlabel polysilicon 205 -825 205 -825 0 3
rlabel polysilicon 212 -819 212 -819 0 1
rlabel polysilicon 212 -825 212 -825 0 3
rlabel polysilicon 219 -819 219 -819 0 1
rlabel polysilicon 219 -825 219 -825 0 3
rlabel polysilicon 226 -819 226 -819 0 1
rlabel polysilicon 226 -825 226 -825 0 3
rlabel polysilicon 233 -819 233 -819 0 1
rlabel polysilicon 233 -825 233 -825 0 3
rlabel polysilicon 243 -819 243 -819 0 2
rlabel polysilicon 247 -819 247 -819 0 1
rlabel polysilicon 247 -825 247 -825 0 3
rlabel polysilicon 254 -819 254 -819 0 1
rlabel polysilicon 254 -825 254 -825 0 3
rlabel polysilicon 261 -819 261 -819 0 1
rlabel polysilicon 261 -825 261 -825 0 3
rlabel polysilicon 268 -819 268 -819 0 1
rlabel polysilicon 268 -825 268 -825 0 3
rlabel polysilicon 275 -819 275 -819 0 1
rlabel polysilicon 278 -819 278 -819 0 2
rlabel polysilicon 275 -825 275 -825 0 3
rlabel polysilicon 278 -825 278 -825 0 4
rlabel polysilicon 282 -819 282 -819 0 1
rlabel polysilicon 285 -819 285 -819 0 2
rlabel polysilicon 285 -825 285 -825 0 4
rlabel polysilicon 289 -819 289 -819 0 1
rlabel polysilicon 289 -825 289 -825 0 3
rlabel polysilicon 299 -819 299 -819 0 2
rlabel polysilicon 296 -825 296 -825 0 3
rlabel polysilicon 303 -819 303 -819 0 1
rlabel polysilicon 303 -825 303 -825 0 3
rlabel polysilicon 310 -819 310 -819 0 1
rlabel polysilicon 313 -819 313 -819 0 2
rlabel polysilicon 320 -819 320 -819 0 2
rlabel polysilicon 317 -825 317 -825 0 3
rlabel polysilicon 320 -825 320 -825 0 4
rlabel polysilicon 327 -819 327 -819 0 2
rlabel polysilicon 331 -819 331 -819 0 1
rlabel polysilicon 331 -825 331 -825 0 3
rlabel polysilicon 334 -825 334 -825 0 4
rlabel polysilicon 338 -819 338 -819 0 1
rlabel polysilicon 341 -819 341 -819 0 2
rlabel polysilicon 338 -825 338 -825 0 3
rlabel polysilicon 345 -819 345 -819 0 1
rlabel polysilicon 345 -825 345 -825 0 3
rlabel polysilicon 352 -819 352 -819 0 1
rlabel polysilicon 355 -825 355 -825 0 4
rlabel polysilicon 359 -819 359 -819 0 1
rlabel polysilicon 359 -825 359 -825 0 3
rlabel polysilicon 366 -819 366 -819 0 1
rlabel polysilicon 366 -825 366 -825 0 3
rlabel polysilicon 373 -819 373 -819 0 1
rlabel polysilicon 376 -819 376 -819 0 2
rlabel polysilicon 373 -825 373 -825 0 3
rlabel polysilicon 376 -825 376 -825 0 4
rlabel polysilicon 380 -819 380 -819 0 1
rlabel polysilicon 380 -825 380 -825 0 3
rlabel polysilicon 387 -819 387 -819 0 1
rlabel polysilicon 390 -819 390 -819 0 2
rlabel polysilicon 394 -819 394 -819 0 1
rlabel polysilicon 394 -825 394 -825 0 3
rlabel polysilicon 401 -825 401 -825 0 3
rlabel polysilicon 404 -825 404 -825 0 4
rlabel polysilicon 408 -819 408 -819 0 1
rlabel polysilicon 408 -825 408 -825 0 3
rlabel polysilicon 415 -819 415 -819 0 1
rlabel polysilicon 415 -825 415 -825 0 3
rlabel polysilicon 422 -819 422 -819 0 1
rlabel polysilicon 422 -825 422 -825 0 3
rlabel polysilicon 429 -819 429 -819 0 1
rlabel polysilicon 429 -825 429 -825 0 3
rlabel polysilicon 436 -819 436 -819 0 1
rlabel polysilicon 436 -825 436 -825 0 3
rlabel polysilicon 443 -819 443 -819 0 1
rlabel polysilicon 443 -825 443 -825 0 3
rlabel polysilicon 450 -819 450 -819 0 1
rlabel polysilicon 450 -825 450 -825 0 3
rlabel polysilicon 457 -819 457 -819 0 1
rlabel polysilicon 457 -825 457 -825 0 3
rlabel polysilicon 464 -819 464 -819 0 1
rlabel polysilicon 464 -825 464 -825 0 3
rlabel polysilicon 471 -819 471 -819 0 1
rlabel polysilicon 471 -825 471 -825 0 3
rlabel polysilicon 478 -825 478 -825 0 3
rlabel polysilicon 485 -819 485 -819 0 1
rlabel polysilicon 485 -825 485 -825 0 3
rlabel polysilicon 492 -819 492 -819 0 1
rlabel polysilicon 492 -825 492 -825 0 3
rlabel polysilicon 499 -819 499 -819 0 1
rlabel polysilicon 499 -825 499 -825 0 3
rlabel polysilicon 506 -819 506 -819 0 1
rlabel polysilicon 506 -825 506 -825 0 3
rlabel polysilicon 513 -819 513 -819 0 1
rlabel polysilicon 520 -819 520 -819 0 1
rlabel polysilicon 520 -825 520 -825 0 3
rlabel polysilicon 527 -819 527 -819 0 1
rlabel polysilicon 527 -825 527 -825 0 3
rlabel polysilicon 537 -819 537 -819 0 2
rlabel polysilicon 541 -819 541 -819 0 1
rlabel polysilicon 541 -825 541 -825 0 3
rlabel polysilicon 548 -819 548 -819 0 1
rlabel polysilicon 548 -825 548 -825 0 3
rlabel polysilicon 555 -819 555 -819 0 1
rlabel polysilicon 558 -819 558 -819 0 2
rlabel polysilicon 562 -819 562 -819 0 1
rlabel polysilicon 562 -825 562 -825 0 3
rlabel polysilicon 569 -819 569 -819 0 1
rlabel polysilicon 572 -825 572 -825 0 4
rlabel polysilicon 576 -819 576 -819 0 1
rlabel polysilicon 576 -825 576 -825 0 3
rlabel polysilicon 583 -819 583 -819 0 1
rlabel polysilicon 583 -825 583 -825 0 3
rlabel polysilicon 590 -819 590 -819 0 1
rlabel polysilicon 590 -825 590 -825 0 3
rlabel polysilicon 597 -819 597 -819 0 1
rlabel polysilicon 604 -819 604 -819 0 1
rlabel polysilicon 604 -825 604 -825 0 3
rlabel polysilicon 618 -819 618 -819 0 1
rlabel polysilicon 618 -825 618 -825 0 3
rlabel polysilicon 2 -862 2 -862 0 1
rlabel polysilicon 2 -868 2 -868 0 3
rlabel polysilicon 9 -862 9 -862 0 1
rlabel polysilicon 9 -868 9 -868 0 3
rlabel polysilicon 16 -862 16 -862 0 1
rlabel polysilicon 16 -868 16 -868 0 3
rlabel polysilicon 23 -862 23 -862 0 1
rlabel polysilicon 23 -868 23 -868 0 3
rlabel polysilicon 33 -862 33 -862 0 2
rlabel polysilicon 30 -868 30 -868 0 3
rlabel polysilicon 37 -862 37 -862 0 1
rlabel polysilicon 37 -868 37 -868 0 3
rlabel polysilicon 40 -868 40 -868 0 4
rlabel polysilicon 44 -868 44 -868 0 3
rlabel polysilicon 47 -868 47 -868 0 4
rlabel polysilicon 51 -862 51 -862 0 1
rlabel polysilicon 51 -868 51 -868 0 3
rlabel polysilicon 61 -862 61 -862 0 2
rlabel polysilicon 61 -868 61 -868 0 4
rlabel polysilicon 65 -862 65 -862 0 1
rlabel polysilicon 65 -868 65 -868 0 3
rlabel polysilicon 72 -862 72 -862 0 1
rlabel polysilicon 72 -868 72 -868 0 3
rlabel polysilicon 79 -868 79 -868 0 3
rlabel polysilicon 86 -862 86 -862 0 1
rlabel polysilicon 86 -868 86 -868 0 3
rlabel polysilicon 93 -862 93 -862 0 1
rlabel polysilicon 93 -868 93 -868 0 3
rlabel polysilicon 100 -862 100 -862 0 1
rlabel polysilicon 100 -868 100 -868 0 3
rlabel polysilicon 107 -862 107 -862 0 1
rlabel polysilicon 107 -868 107 -868 0 3
rlabel polysilicon 114 -862 114 -862 0 1
rlabel polysilicon 114 -868 114 -868 0 3
rlabel polysilicon 121 -862 121 -862 0 1
rlabel polysilicon 121 -868 121 -868 0 3
rlabel polysilicon 128 -862 128 -862 0 1
rlabel polysilicon 128 -868 128 -868 0 3
rlabel polysilicon 135 -862 135 -862 0 1
rlabel polysilicon 135 -868 135 -868 0 3
rlabel polysilicon 142 -862 142 -862 0 1
rlabel polysilicon 149 -862 149 -862 0 1
rlabel polysilicon 149 -868 149 -868 0 3
rlabel polysilicon 156 -862 156 -862 0 1
rlabel polysilicon 156 -868 156 -868 0 3
rlabel polysilicon 163 -862 163 -862 0 1
rlabel polysilicon 163 -868 163 -868 0 3
rlabel polysilicon 170 -862 170 -862 0 1
rlabel polysilicon 173 -862 173 -862 0 2
rlabel polysilicon 173 -868 173 -868 0 4
rlabel polysilicon 180 -862 180 -862 0 2
rlabel polysilicon 184 -862 184 -862 0 1
rlabel polysilicon 184 -868 184 -868 0 3
rlabel polysilicon 191 -862 191 -862 0 1
rlabel polysilicon 194 -862 194 -862 0 2
rlabel polysilicon 191 -868 191 -868 0 3
rlabel polysilicon 198 -862 198 -862 0 1
rlabel polysilicon 201 -862 201 -862 0 2
rlabel polysilicon 205 -862 205 -862 0 1
rlabel polysilicon 205 -868 205 -868 0 3
rlabel polysilicon 208 -868 208 -868 0 4
rlabel polysilicon 215 -862 215 -862 0 2
rlabel polysilicon 222 -862 222 -862 0 2
rlabel polysilicon 219 -868 219 -868 0 3
rlabel polysilicon 222 -868 222 -868 0 4
rlabel polysilicon 226 -862 226 -862 0 1
rlabel polysilicon 229 -862 229 -862 0 2
rlabel polysilicon 226 -868 226 -868 0 3
rlabel polysilicon 233 -862 233 -862 0 1
rlabel polysilicon 233 -868 233 -868 0 3
rlabel polysilicon 240 -862 240 -862 0 1
rlabel polysilicon 240 -868 240 -868 0 3
rlabel polysilicon 247 -862 247 -862 0 1
rlabel polysilicon 247 -868 247 -868 0 3
rlabel polysilicon 254 -862 254 -862 0 1
rlabel polysilicon 254 -868 254 -868 0 3
rlabel polysilicon 261 -862 261 -862 0 1
rlabel polysilicon 268 -862 268 -862 0 1
rlabel polysilicon 268 -868 268 -868 0 3
rlabel polysilicon 275 -862 275 -862 0 1
rlabel polysilicon 275 -868 275 -868 0 3
rlabel polysilicon 282 -862 282 -862 0 1
rlabel polysilicon 282 -868 282 -868 0 3
rlabel polysilicon 289 -862 289 -862 0 1
rlabel polysilicon 292 -862 292 -862 0 2
rlabel polysilicon 289 -868 289 -868 0 3
rlabel polysilicon 292 -868 292 -868 0 4
rlabel polysilicon 296 -862 296 -862 0 1
rlabel polysilicon 296 -868 296 -868 0 3
rlabel polysilicon 303 -862 303 -862 0 1
rlabel polysilicon 303 -868 303 -868 0 3
rlabel polysilicon 310 -862 310 -862 0 1
rlabel polysilicon 310 -868 310 -868 0 3
rlabel polysilicon 317 -862 317 -862 0 1
rlabel polysilicon 320 -862 320 -862 0 2
rlabel polysilicon 320 -868 320 -868 0 4
rlabel polysilicon 324 -862 324 -862 0 1
rlabel polysilicon 324 -868 324 -868 0 3
rlabel polysilicon 331 -862 331 -862 0 1
rlabel polysilicon 331 -868 331 -868 0 3
rlabel polysilicon 338 -862 338 -862 0 1
rlabel polysilicon 338 -868 338 -868 0 3
rlabel polysilicon 345 -862 345 -862 0 1
rlabel polysilicon 348 -862 348 -862 0 2
rlabel polysilicon 348 -868 348 -868 0 4
rlabel polysilicon 352 -862 352 -862 0 1
rlabel polysilicon 352 -868 352 -868 0 3
rlabel polysilicon 359 -862 359 -862 0 1
rlabel polysilicon 359 -868 359 -868 0 3
rlabel polysilicon 366 -862 366 -862 0 1
rlabel polysilicon 366 -868 366 -868 0 3
rlabel polysilicon 373 -862 373 -862 0 1
rlabel polysilicon 373 -868 373 -868 0 3
rlabel polysilicon 376 -868 376 -868 0 4
rlabel polysilicon 380 -862 380 -862 0 1
rlabel polysilicon 380 -868 380 -868 0 3
rlabel polysilicon 387 -862 387 -862 0 1
rlabel polysilicon 387 -868 387 -868 0 3
rlabel polysilicon 394 -862 394 -862 0 1
rlabel polysilicon 394 -868 394 -868 0 3
rlabel polysilicon 401 -862 401 -862 0 1
rlabel polysilicon 401 -868 401 -868 0 3
rlabel polysilicon 408 -862 408 -862 0 1
rlabel polysilicon 408 -868 408 -868 0 3
rlabel polysilicon 415 -862 415 -862 0 1
rlabel polysilicon 415 -868 415 -868 0 3
rlabel polysilicon 425 -862 425 -862 0 2
rlabel polysilicon 425 -868 425 -868 0 4
rlabel polysilicon 429 -862 429 -862 0 1
rlabel polysilicon 429 -868 429 -868 0 3
rlabel polysilicon 436 -862 436 -862 0 1
rlabel polysilicon 436 -868 436 -868 0 3
rlabel polysilicon 443 -862 443 -862 0 1
rlabel polysilicon 443 -868 443 -868 0 3
rlabel polysilicon 450 -868 450 -868 0 3
rlabel polysilicon 453 -868 453 -868 0 4
rlabel polysilicon 457 -862 457 -862 0 1
rlabel polysilicon 457 -868 457 -868 0 3
rlabel polysilicon 464 -862 464 -862 0 1
rlabel polysilicon 464 -868 464 -868 0 3
rlabel polysilicon 471 -862 471 -862 0 1
rlabel polysilicon 471 -868 471 -868 0 3
rlabel polysilicon 478 -862 478 -862 0 1
rlabel polysilicon 478 -868 478 -868 0 3
rlabel polysilicon 485 -862 485 -862 0 1
rlabel polysilicon 485 -868 485 -868 0 3
rlabel polysilicon 492 -862 492 -862 0 1
rlabel polysilicon 492 -868 492 -868 0 3
rlabel polysilicon 499 -862 499 -862 0 1
rlabel polysilicon 499 -868 499 -868 0 3
rlabel polysilicon 506 -862 506 -862 0 1
rlabel polysilicon 506 -868 506 -868 0 3
rlabel polysilicon 513 -862 513 -862 0 1
rlabel polysilicon 516 -862 516 -862 0 2
rlabel polysilicon 513 -868 513 -868 0 3
rlabel polysilicon 516 -868 516 -868 0 4
rlabel polysilicon 520 -862 520 -862 0 1
rlabel polysilicon 520 -868 520 -868 0 3
rlabel polysilicon 527 -862 527 -862 0 1
rlabel polysilicon 527 -868 527 -868 0 3
rlabel polysilicon 534 -862 534 -862 0 1
rlabel polysilicon 537 -868 537 -868 0 4
rlabel polysilicon 544 -868 544 -868 0 4
rlabel polysilicon 548 -862 548 -862 0 1
rlabel polysilicon 548 -868 548 -868 0 3
rlabel polysilicon 555 -862 555 -862 0 1
rlabel polysilicon 555 -868 555 -868 0 3
rlabel polysilicon 562 -862 562 -862 0 1
rlabel polysilicon 562 -868 562 -868 0 3
rlabel polysilicon 2 -917 2 -917 0 1
rlabel polysilicon 2 -923 2 -923 0 3
rlabel polysilicon 9 -923 9 -923 0 3
rlabel polysilicon 16 -917 16 -917 0 1
rlabel polysilicon 16 -923 16 -923 0 3
rlabel polysilicon 23 -917 23 -917 0 1
rlabel polysilicon 23 -923 23 -923 0 3
rlabel polysilicon 30 -923 30 -923 0 3
rlabel polysilicon 37 -917 37 -917 0 1
rlabel polysilicon 44 -917 44 -917 0 1
rlabel polysilicon 54 -917 54 -917 0 2
rlabel polysilicon 58 -923 58 -923 0 3
rlabel polysilicon 65 -917 65 -917 0 1
rlabel polysilicon 68 -917 68 -917 0 2
rlabel polysilicon 72 -923 72 -923 0 3
rlabel polysilicon 79 -917 79 -917 0 1
rlabel polysilicon 79 -923 79 -923 0 3
rlabel polysilicon 86 -917 86 -917 0 1
rlabel polysilicon 86 -923 86 -923 0 3
rlabel polysilicon 96 -917 96 -917 0 2
rlabel polysilicon 93 -923 93 -923 0 3
rlabel polysilicon 96 -923 96 -923 0 4
rlabel polysilicon 100 -917 100 -917 0 1
rlabel polysilicon 103 -917 103 -917 0 2
rlabel polysilicon 100 -923 100 -923 0 3
rlabel polysilicon 110 -923 110 -923 0 4
rlabel polysilicon 114 -917 114 -917 0 1
rlabel polysilicon 114 -923 114 -923 0 3
rlabel polysilicon 121 -917 121 -917 0 1
rlabel polysilicon 124 -917 124 -917 0 2
rlabel polysilicon 124 -923 124 -923 0 4
rlabel polysilicon 131 -917 131 -917 0 2
rlabel polysilicon 128 -923 128 -923 0 3
rlabel polysilicon 135 -917 135 -917 0 1
rlabel polysilicon 135 -923 135 -923 0 3
rlabel polysilicon 142 -917 142 -917 0 1
rlabel polysilicon 142 -923 142 -923 0 3
rlabel polysilicon 149 -917 149 -917 0 1
rlabel polysilicon 152 -917 152 -917 0 2
rlabel polysilicon 152 -923 152 -923 0 4
rlabel polysilicon 156 -917 156 -917 0 1
rlabel polysilicon 156 -923 156 -923 0 3
rlabel polysilicon 163 -917 163 -917 0 1
rlabel polysilicon 163 -923 163 -923 0 3
rlabel polysilicon 173 -917 173 -917 0 2
rlabel polysilicon 170 -923 170 -923 0 3
rlabel polysilicon 173 -923 173 -923 0 4
rlabel polysilicon 177 -917 177 -917 0 1
rlabel polysilicon 177 -923 177 -923 0 3
rlabel polysilicon 184 -917 184 -917 0 1
rlabel polysilicon 184 -923 184 -923 0 3
rlabel polysilicon 187 -923 187 -923 0 4
rlabel polysilicon 191 -917 191 -917 0 1
rlabel polysilicon 194 -917 194 -917 0 2
rlabel polysilicon 194 -923 194 -923 0 4
rlabel polysilicon 198 -917 198 -917 0 1
rlabel polysilicon 201 -917 201 -917 0 2
rlabel polysilicon 198 -923 198 -923 0 3
rlabel polysilicon 208 -917 208 -917 0 2
rlabel polysilicon 208 -923 208 -923 0 4
rlabel polysilicon 212 -917 212 -917 0 1
rlabel polysilicon 212 -923 212 -923 0 3
rlabel polysilicon 219 -917 219 -917 0 1
rlabel polysilicon 219 -923 219 -923 0 3
rlabel polysilicon 229 -917 229 -917 0 2
rlabel polysilicon 233 -917 233 -917 0 1
rlabel polysilicon 233 -923 233 -923 0 3
rlabel polysilicon 240 -917 240 -917 0 1
rlabel polysilicon 243 -917 243 -917 0 2
rlabel polysilicon 240 -923 240 -923 0 3
rlabel polysilicon 243 -923 243 -923 0 4
rlabel polysilicon 247 -917 247 -917 0 1
rlabel polysilicon 247 -923 247 -923 0 3
rlabel polysilicon 254 -917 254 -917 0 1
rlabel polysilicon 254 -923 254 -923 0 3
rlabel polysilicon 261 -917 261 -917 0 1
rlabel polysilicon 261 -923 261 -923 0 3
rlabel polysilicon 268 -917 268 -917 0 1
rlabel polysilicon 268 -923 268 -923 0 3
rlabel polysilicon 275 -917 275 -917 0 1
rlabel polysilicon 275 -923 275 -923 0 3
rlabel polysilicon 282 -917 282 -917 0 1
rlabel polysilicon 282 -923 282 -923 0 3
rlabel polysilicon 289 -917 289 -917 0 1
rlabel polysilicon 292 -917 292 -917 0 2
rlabel polysilicon 289 -923 289 -923 0 3
rlabel polysilicon 299 -917 299 -917 0 2
rlabel polysilicon 306 -917 306 -917 0 2
rlabel polysilicon 303 -923 303 -923 0 3
rlabel polysilicon 306 -923 306 -923 0 4
rlabel polysilicon 313 -917 313 -917 0 2
rlabel polysilicon 310 -923 310 -923 0 3
rlabel polysilicon 317 -917 317 -917 0 1
rlabel polysilicon 317 -923 317 -923 0 3
rlabel polysilicon 324 -917 324 -917 0 1
rlabel polysilicon 324 -923 324 -923 0 3
rlabel polysilicon 331 -917 331 -917 0 1
rlabel polysilicon 331 -923 331 -923 0 3
rlabel polysilicon 338 -917 338 -917 0 1
rlabel polysilicon 338 -923 338 -923 0 3
rlabel polysilicon 345 -917 345 -917 0 1
rlabel polysilicon 345 -923 345 -923 0 3
rlabel polysilicon 352 -917 352 -917 0 1
rlabel polysilicon 352 -923 352 -923 0 3
rlabel polysilicon 359 -923 359 -923 0 3
rlabel polysilicon 362 -923 362 -923 0 4
rlabel polysilicon 366 -917 366 -917 0 1
rlabel polysilicon 366 -923 366 -923 0 3
rlabel polysilicon 373 -917 373 -917 0 1
rlabel polysilicon 373 -923 373 -923 0 3
rlabel polysilicon 380 -917 380 -917 0 1
rlabel polysilicon 380 -923 380 -923 0 3
rlabel polysilicon 387 -917 387 -917 0 1
rlabel polysilicon 387 -923 387 -923 0 3
rlabel polysilicon 394 -917 394 -917 0 1
rlabel polysilicon 394 -923 394 -923 0 3
rlabel polysilicon 401 -917 401 -917 0 1
rlabel polysilicon 401 -923 401 -923 0 3
rlabel polysilicon 408 -917 408 -917 0 1
rlabel polysilicon 408 -923 408 -923 0 3
rlabel polysilicon 415 -917 415 -917 0 1
rlabel polysilicon 415 -923 415 -923 0 3
rlabel polysilicon 422 -917 422 -917 0 1
rlabel polysilicon 422 -923 422 -923 0 3
rlabel polysilicon 429 -917 429 -917 0 1
rlabel polysilicon 429 -923 429 -923 0 3
rlabel polysilicon 436 -917 436 -917 0 1
rlabel polysilicon 436 -923 436 -923 0 3
rlabel polysilicon 446 -917 446 -917 0 2
rlabel polysilicon 450 -917 450 -917 0 1
rlabel polysilicon 450 -923 450 -923 0 3
rlabel polysilicon 457 -917 457 -917 0 1
rlabel polysilicon 457 -923 457 -923 0 3
rlabel polysilicon 464 -917 464 -917 0 1
rlabel polysilicon 464 -923 464 -923 0 3
rlabel polysilicon 471 -917 471 -917 0 1
rlabel polysilicon 474 -923 474 -923 0 4
rlabel polysilicon 478 -917 478 -917 0 1
rlabel polysilicon 478 -923 478 -923 0 3
rlabel polysilicon 485 -917 485 -917 0 1
rlabel polysilicon 485 -923 485 -923 0 3
rlabel polysilicon 492 -917 492 -917 0 1
rlabel polysilicon 492 -923 492 -923 0 3
rlabel polysilicon 499 -917 499 -917 0 1
rlabel polysilicon 499 -923 499 -923 0 3
rlabel polysilicon 506 -917 506 -917 0 1
rlabel polysilicon 506 -923 506 -923 0 3
rlabel polysilicon 513 -917 513 -917 0 1
rlabel polysilicon 513 -923 513 -923 0 3
rlabel polysilicon 520 -917 520 -917 0 1
rlabel polysilicon 520 -923 520 -923 0 3
rlabel polysilicon 527 -917 527 -917 0 1
rlabel polysilicon 530 -917 530 -917 0 2
rlabel polysilicon 530 -923 530 -923 0 4
rlabel polysilicon 534 -917 534 -917 0 1
rlabel polysilicon 534 -923 534 -923 0 3
rlabel polysilicon 541 -917 541 -917 0 1
rlabel polysilicon 541 -923 541 -923 0 3
rlabel polysilicon 548 -917 548 -917 0 1
rlabel polysilicon 548 -923 548 -923 0 3
rlabel polysilicon 23 -970 23 -970 0 1
rlabel polysilicon 23 -976 23 -976 0 3
rlabel polysilicon 30 -970 30 -970 0 1
rlabel polysilicon 30 -976 30 -976 0 3
rlabel polysilicon 37 -970 37 -970 0 1
rlabel polysilicon 37 -976 37 -976 0 3
rlabel polysilicon 44 -970 44 -970 0 1
rlabel polysilicon 54 -970 54 -970 0 2
rlabel polysilicon 58 -970 58 -970 0 1
rlabel polysilicon 58 -976 58 -976 0 3
rlabel polysilicon 65 -970 65 -970 0 1
rlabel polysilicon 68 -970 68 -970 0 2
rlabel polysilicon 65 -976 65 -976 0 3
rlabel polysilicon 68 -976 68 -976 0 4
rlabel polysilicon 72 -970 72 -970 0 1
rlabel polysilicon 72 -976 72 -976 0 3
rlabel polysilicon 79 -970 79 -970 0 1
rlabel polysilicon 79 -976 79 -976 0 3
rlabel polysilicon 86 -970 86 -970 0 1
rlabel polysilicon 86 -976 86 -976 0 3
rlabel polysilicon 93 -970 93 -970 0 1
rlabel polysilicon 93 -976 93 -976 0 3
rlabel polysilicon 100 -970 100 -970 0 1
rlabel polysilicon 100 -976 100 -976 0 3
rlabel polysilicon 110 -970 110 -970 0 2
rlabel polysilicon 107 -976 107 -976 0 3
rlabel polysilicon 110 -976 110 -976 0 4
rlabel polysilicon 114 -970 114 -970 0 1
rlabel polysilicon 117 -970 117 -970 0 2
rlabel polysilicon 117 -976 117 -976 0 4
rlabel polysilicon 121 -970 121 -970 0 1
rlabel polysilicon 121 -976 121 -976 0 3
rlabel polysilicon 128 -976 128 -976 0 3
rlabel polysilicon 131 -976 131 -976 0 4
rlabel polysilicon 135 -970 135 -970 0 1
rlabel polysilicon 135 -976 135 -976 0 3
rlabel polysilicon 142 -970 142 -970 0 1
rlabel polysilicon 145 -970 145 -970 0 2
rlabel polysilicon 142 -976 142 -976 0 3
rlabel polysilicon 149 -970 149 -970 0 1
rlabel polysilicon 152 -970 152 -970 0 2
rlabel polysilicon 156 -970 156 -970 0 1
rlabel polysilicon 156 -976 156 -976 0 3
rlabel polysilicon 166 -970 166 -970 0 2
rlabel polysilicon 170 -970 170 -970 0 1
rlabel polysilicon 170 -976 170 -976 0 3
rlabel polysilicon 177 -970 177 -970 0 1
rlabel polysilicon 177 -976 177 -976 0 3
rlabel polysilicon 184 -970 184 -970 0 1
rlabel polysilicon 187 -970 187 -970 0 2
rlabel polysilicon 184 -976 184 -976 0 3
rlabel polysilicon 191 -970 191 -970 0 1
rlabel polysilicon 191 -976 191 -976 0 3
rlabel polysilicon 198 -970 198 -970 0 1
rlabel polysilicon 201 -970 201 -970 0 2
rlabel polysilicon 198 -976 198 -976 0 3
rlabel polysilicon 201 -976 201 -976 0 4
rlabel polysilicon 205 -970 205 -970 0 1
rlabel polysilicon 208 -970 208 -970 0 2
rlabel polysilicon 208 -976 208 -976 0 4
rlabel polysilicon 212 -970 212 -970 0 1
rlabel polysilicon 212 -976 212 -976 0 3
rlabel polysilicon 219 -970 219 -970 0 1
rlabel polysilicon 219 -976 219 -976 0 3
rlabel polysilicon 226 -970 226 -970 0 1
rlabel polysilicon 229 -976 229 -976 0 4
rlabel polysilicon 233 -970 233 -970 0 1
rlabel polysilicon 240 -970 240 -970 0 1
rlabel polysilicon 240 -976 240 -976 0 3
rlabel polysilicon 247 -970 247 -970 0 1
rlabel polysilicon 247 -976 247 -976 0 3
rlabel polysilicon 254 -970 254 -970 0 1
rlabel polysilicon 254 -976 254 -976 0 3
rlabel polysilicon 261 -970 261 -970 0 1
rlabel polysilicon 264 -970 264 -970 0 2
rlabel polysilicon 261 -976 261 -976 0 3
rlabel polysilicon 264 -976 264 -976 0 4
rlabel polysilicon 268 -970 268 -970 0 1
rlabel polysilicon 268 -976 268 -976 0 3
rlabel polysilicon 275 -970 275 -970 0 1
rlabel polysilicon 275 -976 275 -976 0 3
rlabel polysilicon 278 -976 278 -976 0 4
rlabel polysilicon 282 -970 282 -970 0 1
rlabel polysilicon 285 -970 285 -970 0 2
rlabel polysilicon 289 -970 289 -970 0 1
rlabel polysilicon 289 -976 289 -976 0 3
rlabel polysilicon 296 -970 296 -970 0 1
rlabel polysilicon 299 -970 299 -970 0 2
rlabel polysilicon 299 -976 299 -976 0 4
rlabel polysilicon 303 -970 303 -970 0 1
rlabel polysilicon 303 -976 303 -976 0 3
rlabel polysilicon 310 -970 310 -970 0 1
rlabel polysilicon 310 -976 310 -976 0 3
rlabel polysilicon 320 -970 320 -970 0 2
rlabel polysilicon 320 -976 320 -976 0 4
rlabel polysilicon 324 -970 324 -970 0 1
rlabel polysilicon 324 -976 324 -976 0 3
rlabel polysilicon 331 -970 331 -970 0 1
rlabel polysilicon 331 -976 331 -976 0 3
rlabel polysilicon 338 -970 338 -970 0 1
rlabel polysilicon 338 -976 338 -976 0 3
rlabel polysilicon 345 -970 345 -970 0 1
rlabel polysilicon 345 -976 345 -976 0 3
rlabel polysilicon 352 -970 352 -970 0 1
rlabel polysilicon 352 -976 352 -976 0 3
rlabel polysilicon 359 -970 359 -970 0 1
rlabel polysilicon 359 -976 359 -976 0 3
rlabel polysilicon 366 -970 366 -970 0 1
rlabel polysilicon 366 -976 366 -976 0 3
rlabel polysilicon 373 -970 373 -970 0 1
rlabel polysilicon 373 -976 373 -976 0 3
rlabel polysilicon 383 -970 383 -970 0 2
rlabel polysilicon 380 -976 380 -976 0 3
rlabel polysilicon 387 -970 387 -970 0 1
rlabel polysilicon 387 -976 387 -976 0 3
rlabel polysilicon 394 -970 394 -970 0 1
rlabel polysilicon 394 -976 394 -976 0 3
rlabel polysilicon 401 -970 401 -970 0 1
rlabel polysilicon 401 -976 401 -976 0 3
rlabel polysilicon 411 -970 411 -970 0 2
rlabel polysilicon 411 -976 411 -976 0 4
rlabel polysilicon 415 -970 415 -970 0 1
rlabel polysilicon 415 -976 415 -976 0 3
rlabel polysilicon 422 -976 422 -976 0 3
rlabel polysilicon 429 -970 429 -970 0 1
rlabel polysilicon 429 -976 429 -976 0 3
rlabel polysilicon 436 -970 436 -970 0 1
rlabel polysilicon 436 -976 436 -976 0 3
rlabel polysilicon 443 -970 443 -970 0 1
rlabel polysilicon 443 -976 443 -976 0 3
rlabel polysilicon 450 -970 450 -970 0 1
rlabel polysilicon 450 -976 450 -976 0 3
rlabel polysilicon 457 -970 457 -970 0 1
rlabel polysilicon 457 -976 457 -976 0 3
rlabel polysilicon 464 -970 464 -970 0 1
rlabel polysilicon 467 -970 467 -970 0 2
rlabel polysilicon 464 -976 464 -976 0 3
rlabel polysilicon 471 -970 471 -970 0 1
rlabel polysilicon 471 -976 471 -976 0 3
rlabel polysilicon 478 -970 478 -970 0 1
rlabel polysilicon 481 -970 481 -970 0 2
rlabel polysilicon 478 -976 478 -976 0 3
rlabel polysilicon 485 -970 485 -970 0 1
rlabel polysilicon 485 -976 485 -976 0 3
rlabel polysilicon 492 -970 492 -970 0 1
rlabel polysilicon 492 -976 492 -976 0 3
rlabel polysilicon 499 -970 499 -970 0 1
rlabel polysilicon 499 -976 499 -976 0 3
rlabel polysilicon 506 -970 506 -970 0 1
rlabel polysilicon 509 -970 509 -970 0 2
rlabel polysilicon 509 -976 509 -976 0 4
rlabel polysilicon 520 -970 520 -970 0 1
rlabel polysilicon 520 -976 520 -976 0 3
rlabel polysilicon 16 -1011 16 -1011 0 1
rlabel polysilicon 16 -1017 16 -1017 0 3
rlabel polysilicon 26 -1011 26 -1011 0 2
rlabel polysilicon 30 -1011 30 -1011 0 1
rlabel polysilicon 30 -1017 30 -1017 0 3
rlabel polysilicon 37 -1011 37 -1011 0 1
rlabel polysilicon 37 -1017 37 -1017 0 3
rlabel polysilicon 47 -1017 47 -1017 0 4
rlabel polysilicon 51 -1011 51 -1011 0 1
rlabel polysilicon 51 -1017 51 -1017 0 3
rlabel polysilicon 58 -1011 58 -1011 0 1
rlabel polysilicon 58 -1017 58 -1017 0 3
rlabel polysilicon 65 -1011 65 -1011 0 1
rlabel polysilicon 68 -1011 68 -1011 0 2
rlabel polysilicon 72 -1011 72 -1011 0 1
rlabel polysilicon 72 -1017 72 -1017 0 3
rlabel polysilicon 79 -1011 79 -1011 0 1
rlabel polysilicon 79 -1017 79 -1017 0 3
rlabel polysilicon 86 -1017 86 -1017 0 3
rlabel polysilicon 89 -1017 89 -1017 0 4
rlabel polysilicon 96 -1011 96 -1011 0 2
rlabel polysilicon 96 -1017 96 -1017 0 4
rlabel polysilicon 100 -1011 100 -1011 0 1
rlabel polysilicon 100 -1017 100 -1017 0 3
rlabel polysilicon 107 -1011 107 -1011 0 1
rlabel polysilicon 107 -1017 107 -1017 0 3
rlabel polysilicon 114 -1011 114 -1011 0 1
rlabel polysilicon 117 -1011 117 -1011 0 2
rlabel polysilicon 114 -1017 114 -1017 0 3
rlabel polysilicon 117 -1017 117 -1017 0 4
rlabel polysilicon 121 -1011 121 -1011 0 1
rlabel polysilicon 121 -1017 121 -1017 0 3
rlabel polysilicon 128 -1011 128 -1011 0 1
rlabel polysilicon 131 -1011 131 -1011 0 2
rlabel polysilicon 135 -1011 135 -1011 0 1
rlabel polysilicon 135 -1017 135 -1017 0 3
rlabel polysilicon 142 -1011 142 -1011 0 1
rlabel polysilicon 142 -1017 142 -1017 0 3
rlabel polysilicon 149 -1011 149 -1011 0 1
rlabel polysilicon 149 -1017 149 -1017 0 3
rlabel polysilicon 156 -1011 156 -1011 0 1
rlabel polysilicon 156 -1017 156 -1017 0 3
rlabel polysilicon 163 -1011 163 -1011 0 1
rlabel polysilicon 163 -1017 163 -1017 0 3
rlabel polysilicon 170 -1011 170 -1011 0 1
rlabel polysilicon 173 -1011 173 -1011 0 2
rlabel polysilicon 177 -1011 177 -1011 0 1
rlabel polysilicon 177 -1017 177 -1017 0 3
rlabel polysilicon 187 -1011 187 -1011 0 2
rlabel polysilicon 184 -1017 184 -1017 0 3
rlabel polysilicon 187 -1017 187 -1017 0 4
rlabel polysilicon 191 -1011 191 -1011 0 1
rlabel polysilicon 194 -1017 194 -1017 0 4
rlabel polysilicon 198 -1011 198 -1011 0 1
rlabel polysilicon 201 -1011 201 -1011 0 2
rlabel polysilicon 201 -1017 201 -1017 0 4
rlabel polysilicon 205 -1011 205 -1011 0 1
rlabel polysilicon 208 -1011 208 -1011 0 2
rlabel polysilicon 208 -1017 208 -1017 0 4
rlabel polysilicon 212 -1011 212 -1011 0 1
rlabel polysilicon 212 -1017 212 -1017 0 3
rlabel polysilicon 219 -1011 219 -1011 0 1
rlabel polysilicon 219 -1017 219 -1017 0 3
rlabel polysilicon 226 -1011 226 -1011 0 1
rlabel polysilicon 229 -1011 229 -1011 0 2
rlabel polysilicon 226 -1017 226 -1017 0 3
rlabel polysilicon 229 -1017 229 -1017 0 4
rlabel polysilicon 233 -1011 233 -1011 0 1
rlabel polysilicon 236 -1011 236 -1011 0 2
rlabel polysilicon 233 -1017 233 -1017 0 3
rlabel polysilicon 240 -1011 240 -1011 0 1
rlabel polysilicon 240 -1017 240 -1017 0 3
rlabel polysilicon 247 -1011 247 -1011 0 1
rlabel polysilicon 247 -1017 247 -1017 0 3
rlabel polysilicon 254 -1011 254 -1011 0 1
rlabel polysilicon 254 -1017 254 -1017 0 3
rlabel polysilicon 261 -1011 261 -1011 0 1
rlabel polysilicon 261 -1017 261 -1017 0 3
rlabel polysilicon 271 -1011 271 -1011 0 2
rlabel polysilicon 268 -1017 268 -1017 0 3
rlabel polysilicon 275 -1017 275 -1017 0 3
rlabel polysilicon 278 -1017 278 -1017 0 4
rlabel polysilicon 282 -1011 282 -1011 0 1
rlabel polysilicon 285 -1017 285 -1017 0 4
rlabel polysilicon 289 -1011 289 -1011 0 1
rlabel polysilicon 292 -1011 292 -1011 0 2
rlabel polysilicon 292 -1017 292 -1017 0 4
rlabel polysilicon 296 -1011 296 -1011 0 1
rlabel polysilicon 299 -1011 299 -1011 0 2
rlabel polysilicon 303 -1011 303 -1011 0 1
rlabel polysilicon 303 -1017 303 -1017 0 3
rlabel polysilicon 310 -1011 310 -1011 0 1
rlabel polysilicon 310 -1017 310 -1017 0 3
rlabel polysilicon 317 -1011 317 -1011 0 1
rlabel polysilicon 317 -1017 317 -1017 0 3
rlabel polysilicon 324 -1011 324 -1011 0 1
rlabel polysilicon 324 -1017 324 -1017 0 3
rlabel polysilicon 327 -1017 327 -1017 0 4
rlabel polysilicon 331 -1011 331 -1011 0 1
rlabel polysilicon 331 -1017 331 -1017 0 3
rlabel polysilicon 338 -1011 338 -1011 0 1
rlabel polysilicon 338 -1017 338 -1017 0 3
rlabel polysilicon 345 -1011 345 -1011 0 1
rlabel polysilicon 345 -1017 345 -1017 0 3
rlabel polysilicon 352 -1011 352 -1011 0 1
rlabel polysilicon 352 -1017 352 -1017 0 3
rlabel polysilicon 359 -1011 359 -1011 0 1
rlabel polysilicon 359 -1017 359 -1017 0 3
rlabel polysilicon 366 -1011 366 -1011 0 1
rlabel polysilicon 369 -1017 369 -1017 0 4
rlabel polysilicon 373 -1011 373 -1011 0 1
rlabel polysilicon 373 -1017 373 -1017 0 3
rlabel polysilicon 380 -1011 380 -1011 0 1
rlabel polysilicon 380 -1017 380 -1017 0 3
rlabel polysilicon 387 -1011 387 -1011 0 1
rlabel polysilicon 390 -1011 390 -1011 0 2
rlabel polysilicon 387 -1017 387 -1017 0 3
rlabel polysilicon 394 -1011 394 -1011 0 1
rlabel polysilicon 394 -1017 394 -1017 0 3
rlabel polysilicon 401 -1011 401 -1011 0 1
rlabel polysilicon 401 -1017 401 -1017 0 3
rlabel polysilicon 408 -1011 408 -1011 0 1
rlabel polysilicon 408 -1017 408 -1017 0 3
rlabel polysilicon 415 -1011 415 -1011 0 1
rlabel polysilicon 415 -1017 415 -1017 0 3
rlabel polysilicon 422 -1011 422 -1011 0 1
rlabel polysilicon 422 -1017 422 -1017 0 3
rlabel polysilicon 429 -1011 429 -1011 0 1
rlabel polysilicon 432 -1011 432 -1011 0 2
rlabel polysilicon 436 -1011 436 -1011 0 1
rlabel polysilicon 436 -1017 436 -1017 0 3
rlabel polysilicon 443 -1011 443 -1011 0 1
rlabel polysilicon 446 -1011 446 -1011 0 2
rlabel polysilicon 443 -1017 443 -1017 0 3
rlabel polysilicon 453 -1017 453 -1017 0 4
rlabel polysilicon 457 -1011 457 -1011 0 1
rlabel polysilicon 457 -1017 457 -1017 0 3
rlabel polysilicon 464 -1011 464 -1011 0 1
rlabel polysilicon 464 -1017 464 -1017 0 3
rlabel polysilicon 471 -1011 471 -1011 0 1
rlabel polysilicon 471 -1017 471 -1017 0 3
rlabel polysilicon 478 -1011 478 -1011 0 1
rlabel polysilicon 478 -1017 478 -1017 0 3
rlabel polysilicon 520 -1017 520 -1017 0 3
rlabel polysilicon 523 -1017 523 -1017 0 4
rlabel polysilicon 527 -1011 527 -1011 0 1
rlabel polysilicon 527 -1017 527 -1017 0 3
rlabel polysilicon 65 -1048 65 -1048 0 1
rlabel polysilicon 65 -1054 65 -1054 0 3
rlabel polysilicon 72 -1048 72 -1048 0 1
rlabel polysilicon 72 -1054 72 -1054 0 3
rlabel polysilicon 79 -1054 79 -1054 0 3
rlabel polysilicon 86 -1048 86 -1048 0 1
rlabel polysilicon 89 -1054 89 -1054 0 4
rlabel polysilicon 93 -1048 93 -1048 0 1
rlabel polysilicon 93 -1054 93 -1054 0 3
rlabel polysilicon 103 -1048 103 -1048 0 2
rlabel polysilicon 103 -1054 103 -1054 0 4
rlabel polysilicon 107 -1048 107 -1048 0 1
rlabel polysilicon 107 -1054 107 -1054 0 3
rlabel polysilicon 114 -1048 114 -1048 0 1
rlabel polysilicon 117 -1048 117 -1048 0 2
rlabel polysilicon 114 -1054 114 -1054 0 3
rlabel polysilicon 117 -1054 117 -1054 0 4
rlabel polysilicon 121 -1048 121 -1048 0 1
rlabel polysilicon 121 -1054 121 -1054 0 3
rlabel polysilicon 128 -1048 128 -1048 0 1
rlabel polysilicon 128 -1054 128 -1054 0 3
rlabel polysilicon 135 -1048 135 -1048 0 1
rlabel polysilicon 135 -1054 135 -1054 0 3
rlabel polysilicon 142 -1054 142 -1054 0 3
rlabel polysilicon 145 -1054 145 -1054 0 4
rlabel polysilicon 149 -1048 149 -1048 0 1
rlabel polysilicon 149 -1054 149 -1054 0 3
rlabel polysilicon 152 -1054 152 -1054 0 4
rlabel polysilicon 159 -1054 159 -1054 0 4
rlabel polysilicon 166 -1048 166 -1048 0 2
rlabel polysilicon 163 -1054 163 -1054 0 3
rlabel polysilicon 170 -1048 170 -1048 0 1
rlabel polysilicon 177 -1048 177 -1048 0 1
rlabel polysilicon 177 -1054 177 -1054 0 3
rlabel polysilicon 184 -1048 184 -1048 0 1
rlabel polysilicon 184 -1054 184 -1054 0 3
rlabel polysilicon 191 -1048 191 -1048 0 1
rlabel polysilicon 191 -1054 191 -1054 0 3
rlabel polysilicon 201 -1048 201 -1048 0 2
rlabel polysilicon 201 -1054 201 -1054 0 4
rlabel polysilicon 205 -1048 205 -1048 0 1
rlabel polysilicon 208 -1048 208 -1048 0 2
rlabel polysilicon 205 -1054 205 -1054 0 3
rlabel polysilicon 208 -1054 208 -1054 0 4
rlabel polysilicon 212 -1048 212 -1048 0 1
rlabel polysilicon 215 -1048 215 -1048 0 2
rlabel polysilicon 212 -1054 212 -1054 0 3
rlabel polysilicon 215 -1054 215 -1054 0 4
rlabel polysilicon 219 -1048 219 -1048 0 1
rlabel polysilicon 219 -1054 219 -1054 0 3
rlabel polysilicon 226 -1048 226 -1048 0 1
rlabel polysilicon 229 -1048 229 -1048 0 2
rlabel polysilicon 236 -1048 236 -1048 0 2
rlabel polysilicon 236 -1054 236 -1054 0 4
rlabel polysilicon 240 -1048 240 -1048 0 1
rlabel polysilicon 240 -1054 240 -1054 0 3
rlabel polysilicon 247 -1048 247 -1048 0 1
rlabel polysilicon 250 -1048 250 -1048 0 2
rlabel polysilicon 247 -1054 247 -1054 0 3
rlabel polysilicon 250 -1054 250 -1054 0 4
rlabel polysilicon 254 -1048 254 -1048 0 1
rlabel polysilicon 254 -1054 254 -1054 0 3
rlabel polysilicon 261 -1048 261 -1048 0 1
rlabel polysilicon 261 -1054 261 -1054 0 3
rlabel polysilicon 268 -1048 268 -1048 0 1
rlabel polysilicon 268 -1054 268 -1054 0 3
rlabel polysilicon 275 -1048 275 -1048 0 1
rlabel polysilicon 275 -1054 275 -1054 0 3
rlabel polysilicon 282 -1048 282 -1048 0 1
rlabel polysilicon 282 -1054 282 -1054 0 3
rlabel polysilicon 289 -1048 289 -1048 0 1
rlabel polysilicon 292 -1048 292 -1048 0 2
rlabel polysilicon 289 -1054 289 -1054 0 3
rlabel polysilicon 292 -1054 292 -1054 0 4
rlabel polysilicon 296 -1048 296 -1048 0 1
rlabel polysilicon 296 -1054 296 -1054 0 3
rlabel polysilicon 303 -1048 303 -1048 0 1
rlabel polysilicon 303 -1054 303 -1054 0 3
rlabel polysilicon 310 -1048 310 -1048 0 1
rlabel polysilicon 310 -1054 310 -1054 0 3
rlabel polysilicon 317 -1048 317 -1048 0 1
rlabel polysilicon 317 -1054 317 -1054 0 3
rlabel polysilicon 324 -1048 324 -1048 0 1
rlabel polysilicon 324 -1054 324 -1054 0 3
rlabel polysilicon 334 -1048 334 -1048 0 2
rlabel polysilicon 334 -1054 334 -1054 0 4
rlabel polysilicon 338 -1048 338 -1048 0 1
rlabel polysilicon 338 -1054 338 -1054 0 3
rlabel polysilicon 345 -1048 345 -1048 0 1
rlabel polysilicon 345 -1054 345 -1054 0 3
rlabel polysilicon 355 -1048 355 -1048 0 2
rlabel polysilicon 359 -1048 359 -1048 0 1
rlabel polysilicon 359 -1054 359 -1054 0 3
rlabel polysilicon 362 -1054 362 -1054 0 4
rlabel polysilicon 366 -1048 366 -1048 0 1
rlabel polysilicon 366 -1054 366 -1054 0 3
rlabel polysilicon 373 -1048 373 -1048 0 1
rlabel polysilicon 373 -1054 373 -1054 0 3
rlabel polysilicon 380 -1048 380 -1048 0 1
rlabel polysilicon 380 -1054 380 -1054 0 3
rlabel polysilicon 387 -1048 387 -1048 0 1
rlabel polysilicon 387 -1054 387 -1054 0 3
rlabel polysilicon 394 -1048 394 -1048 0 1
rlabel polysilicon 394 -1054 394 -1054 0 3
rlabel polysilicon 401 -1048 401 -1048 0 1
rlabel polysilicon 401 -1054 401 -1054 0 3
rlabel polysilicon 408 -1048 408 -1048 0 1
rlabel polysilicon 408 -1054 408 -1054 0 3
rlabel polysilicon 415 -1048 415 -1048 0 1
rlabel polysilicon 415 -1054 415 -1054 0 3
rlabel polysilicon 422 -1048 422 -1048 0 1
rlabel polysilicon 429 -1048 429 -1048 0 1
rlabel polysilicon 429 -1054 429 -1054 0 3
rlabel polysilicon 443 -1048 443 -1048 0 1
rlabel polysilicon 450 -1048 450 -1048 0 1
rlabel polysilicon 453 -1048 453 -1048 0 2
rlabel polysilicon 457 -1048 457 -1048 0 1
rlabel polysilicon 457 -1054 457 -1054 0 3
rlabel polysilicon 478 -1048 478 -1048 0 1
rlabel polysilicon 478 -1054 478 -1054 0 3
rlabel polysilicon 516 -1048 516 -1048 0 2
rlabel polysilicon 523 -1048 523 -1048 0 2
rlabel polysilicon 520 -1054 520 -1054 0 3
rlabel polysilicon 527 -1048 527 -1048 0 1
rlabel polysilicon 527 -1054 527 -1054 0 3
rlabel polysilicon 51 -1093 51 -1093 0 1
rlabel polysilicon 51 -1099 51 -1099 0 3
rlabel polysilicon 61 -1093 61 -1093 0 2
rlabel polysilicon 65 -1093 65 -1093 0 1
rlabel polysilicon 65 -1099 65 -1099 0 3
rlabel polysilicon 75 -1093 75 -1093 0 2
rlabel polysilicon 72 -1099 72 -1099 0 3
rlabel polysilicon 79 -1099 79 -1099 0 3
rlabel polysilicon 89 -1099 89 -1099 0 4
rlabel polysilicon 93 -1093 93 -1093 0 1
rlabel polysilicon 93 -1099 93 -1099 0 3
rlabel polysilicon 100 -1093 100 -1093 0 1
rlabel polysilicon 100 -1099 100 -1099 0 3
rlabel polysilicon 107 -1093 107 -1093 0 1
rlabel polysilicon 110 -1093 110 -1093 0 2
rlabel polysilicon 107 -1099 107 -1099 0 3
rlabel polysilicon 110 -1099 110 -1099 0 4
rlabel polysilicon 114 -1093 114 -1093 0 1
rlabel polysilicon 114 -1099 114 -1099 0 3
rlabel polysilicon 121 -1093 121 -1093 0 1
rlabel polysilicon 121 -1099 121 -1099 0 3
rlabel polysilicon 131 -1093 131 -1093 0 2
rlabel polysilicon 135 -1093 135 -1093 0 1
rlabel polysilicon 135 -1099 135 -1099 0 3
rlabel polysilicon 138 -1099 138 -1099 0 4
rlabel polysilicon 142 -1093 142 -1093 0 1
rlabel polysilicon 142 -1099 142 -1099 0 3
rlabel polysilicon 149 -1093 149 -1093 0 1
rlabel polysilicon 149 -1099 149 -1099 0 3
rlabel polysilicon 156 -1093 156 -1093 0 1
rlabel polysilicon 156 -1099 156 -1099 0 3
rlabel polysilicon 163 -1093 163 -1093 0 1
rlabel polysilicon 163 -1099 163 -1099 0 3
rlabel polysilicon 170 -1099 170 -1099 0 3
rlabel polysilicon 177 -1093 177 -1093 0 1
rlabel polysilicon 180 -1093 180 -1093 0 2
rlabel polysilicon 180 -1099 180 -1099 0 4
rlabel polysilicon 184 -1099 184 -1099 0 3
rlabel polysilicon 187 -1099 187 -1099 0 4
rlabel polysilicon 191 -1099 191 -1099 0 3
rlabel polysilicon 198 -1093 198 -1093 0 1
rlabel polysilicon 198 -1099 198 -1099 0 3
rlabel polysilicon 205 -1093 205 -1093 0 1
rlabel polysilicon 205 -1099 205 -1099 0 3
rlabel polysilicon 212 -1093 212 -1093 0 1
rlabel polysilicon 212 -1099 212 -1099 0 3
rlabel polysilicon 219 -1093 219 -1093 0 1
rlabel polysilicon 222 -1093 222 -1093 0 2
rlabel polysilicon 222 -1099 222 -1099 0 4
rlabel polysilicon 226 -1093 226 -1093 0 1
rlabel polysilicon 226 -1099 226 -1099 0 3
rlabel polysilicon 233 -1093 233 -1093 0 1
rlabel polysilicon 236 -1093 236 -1093 0 2
rlabel polysilicon 236 -1099 236 -1099 0 4
rlabel polysilicon 240 -1093 240 -1093 0 1
rlabel polysilicon 240 -1099 240 -1099 0 3
rlabel polysilicon 247 -1093 247 -1093 0 1
rlabel polysilicon 247 -1099 247 -1099 0 3
rlabel polysilicon 254 -1093 254 -1093 0 1
rlabel polysilicon 254 -1099 254 -1099 0 3
rlabel polysilicon 261 -1093 261 -1093 0 1
rlabel polysilicon 261 -1099 261 -1099 0 3
rlabel polysilicon 268 -1093 268 -1093 0 1
rlabel polysilicon 268 -1099 268 -1099 0 3
rlabel polysilicon 275 -1093 275 -1093 0 1
rlabel polysilicon 275 -1099 275 -1099 0 3
rlabel polysilicon 282 -1093 282 -1093 0 1
rlabel polysilicon 282 -1099 282 -1099 0 3
rlabel polysilicon 289 -1093 289 -1093 0 1
rlabel polysilicon 299 -1093 299 -1093 0 2
rlabel polysilicon 296 -1099 296 -1099 0 3
rlabel polysilicon 299 -1099 299 -1099 0 4
rlabel polysilicon 306 -1093 306 -1093 0 2
rlabel polysilicon 303 -1099 303 -1099 0 3
rlabel polysilicon 306 -1099 306 -1099 0 4
rlabel polysilicon 310 -1093 310 -1093 0 1
rlabel polysilicon 310 -1099 310 -1099 0 3
rlabel polysilicon 317 -1093 317 -1093 0 1
rlabel polysilicon 320 -1093 320 -1093 0 2
rlabel polysilicon 320 -1099 320 -1099 0 4
rlabel polysilicon 324 -1093 324 -1093 0 1
rlabel polysilicon 324 -1099 324 -1099 0 3
rlabel polysilicon 331 -1093 331 -1093 0 1
rlabel polysilicon 331 -1099 331 -1099 0 3
rlabel polysilicon 338 -1093 338 -1093 0 1
rlabel polysilicon 338 -1099 338 -1099 0 3
rlabel polysilicon 345 -1093 345 -1093 0 1
rlabel polysilicon 345 -1099 345 -1099 0 3
rlabel polysilicon 352 -1093 352 -1093 0 1
rlabel polysilicon 352 -1099 352 -1099 0 3
rlabel polysilicon 359 -1093 359 -1093 0 1
rlabel polysilicon 362 -1093 362 -1093 0 2
rlabel polysilicon 359 -1099 359 -1099 0 3
rlabel polysilicon 366 -1093 366 -1093 0 1
rlabel polysilicon 366 -1099 366 -1099 0 3
rlabel polysilicon 373 -1093 373 -1093 0 1
rlabel polysilicon 373 -1099 373 -1099 0 3
rlabel polysilicon 376 -1099 376 -1099 0 4
rlabel polysilicon 380 -1093 380 -1093 0 1
rlabel polysilicon 380 -1099 380 -1099 0 3
rlabel polysilicon 387 -1093 387 -1093 0 1
rlabel polysilicon 390 -1093 390 -1093 0 2
rlabel polysilicon 387 -1099 387 -1099 0 3
rlabel polysilicon 394 -1093 394 -1093 0 1
rlabel polysilicon 394 -1099 394 -1099 0 3
rlabel polysilicon 401 -1093 401 -1093 0 1
rlabel polysilicon 401 -1099 401 -1099 0 3
rlabel polysilicon 408 -1093 408 -1093 0 1
rlabel polysilicon 408 -1099 408 -1099 0 3
rlabel polysilicon 415 -1099 415 -1099 0 3
rlabel polysilicon 418 -1099 418 -1099 0 4
rlabel polysilicon 422 -1093 422 -1093 0 1
rlabel polysilicon 422 -1099 422 -1099 0 3
rlabel polysilicon 429 -1093 429 -1093 0 1
rlabel polysilicon 429 -1099 429 -1099 0 3
rlabel polysilicon 436 -1093 436 -1093 0 1
rlabel polysilicon 460 -1099 460 -1099 0 4
rlabel polysilicon 464 -1093 464 -1093 0 1
rlabel polysilicon 464 -1099 464 -1099 0 3
rlabel polysilicon 478 -1093 478 -1093 0 1
rlabel polysilicon 478 -1099 478 -1099 0 3
rlabel polysilicon 30 -1130 30 -1130 0 1
rlabel polysilicon 30 -1136 30 -1136 0 3
rlabel polysilicon 37 -1130 37 -1130 0 1
rlabel polysilicon 37 -1136 37 -1136 0 3
rlabel polysilicon 44 -1130 44 -1130 0 1
rlabel polysilicon 44 -1136 44 -1136 0 3
rlabel polysilicon 54 -1130 54 -1130 0 2
rlabel polysilicon 58 -1130 58 -1130 0 1
rlabel polysilicon 58 -1136 58 -1136 0 3
rlabel polysilicon 65 -1130 65 -1130 0 1
rlabel polysilicon 65 -1136 65 -1136 0 3
rlabel polysilicon 75 -1130 75 -1130 0 2
rlabel polysilicon 75 -1136 75 -1136 0 4
rlabel polysilicon 79 -1130 79 -1130 0 1
rlabel polysilicon 82 -1130 82 -1130 0 2
rlabel polysilicon 79 -1136 79 -1136 0 3
rlabel polysilicon 86 -1130 86 -1130 0 1
rlabel polysilicon 89 -1136 89 -1136 0 4
rlabel polysilicon 96 -1136 96 -1136 0 4
rlabel polysilicon 100 -1130 100 -1130 0 1
rlabel polysilicon 100 -1136 100 -1136 0 3
rlabel polysilicon 107 -1130 107 -1130 0 1
rlabel polysilicon 107 -1136 107 -1136 0 3
rlabel polysilicon 114 -1130 114 -1130 0 1
rlabel polysilicon 117 -1136 117 -1136 0 4
rlabel polysilicon 121 -1130 121 -1130 0 1
rlabel polysilicon 121 -1136 121 -1136 0 3
rlabel polysilicon 131 -1130 131 -1130 0 2
rlabel polysilicon 128 -1136 128 -1136 0 3
rlabel polysilicon 135 -1130 135 -1130 0 1
rlabel polysilicon 135 -1136 135 -1136 0 3
rlabel polysilicon 142 -1130 142 -1130 0 1
rlabel polysilicon 142 -1136 142 -1136 0 3
rlabel polysilicon 149 -1130 149 -1130 0 1
rlabel polysilicon 149 -1136 149 -1136 0 3
rlabel polysilicon 159 -1130 159 -1130 0 2
rlabel polysilicon 159 -1136 159 -1136 0 4
rlabel polysilicon 163 -1130 163 -1130 0 1
rlabel polysilicon 163 -1136 163 -1136 0 3
rlabel polysilicon 170 -1130 170 -1130 0 1
rlabel polysilicon 170 -1136 170 -1136 0 3
rlabel polysilicon 177 -1130 177 -1130 0 1
rlabel polysilicon 177 -1136 177 -1136 0 3
rlabel polysilicon 184 -1130 184 -1130 0 1
rlabel polysilicon 184 -1136 184 -1136 0 3
rlabel polysilicon 191 -1130 191 -1130 0 1
rlabel polysilicon 194 -1130 194 -1130 0 2
rlabel polysilicon 191 -1136 191 -1136 0 3
rlabel polysilicon 198 -1136 198 -1136 0 3
rlabel polysilicon 201 -1136 201 -1136 0 4
rlabel polysilicon 205 -1130 205 -1130 0 1
rlabel polysilicon 208 -1130 208 -1130 0 2
rlabel polysilicon 205 -1136 205 -1136 0 3
rlabel polysilicon 208 -1136 208 -1136 0 4
rlabel polysilicon 212 -1130 212 -1130 0 1
rlabel polysilicon 212 -1136 212 -1136 0 3
rlabel polysilicon 219 -1130 219 -1130 0 1
rlabel polysilicon 219 -1136 219 -1136 0 3
rlabel polysilicon 226 -1130 226 -1130 0 1
rlabel polysilicon 226 -1136 226 -1136 0 3
rlabel polysilicon 229 -1136 229 -1136 0 4
rlabel polysilicon 233 -1130 233 -1130 0 1
rlabel polysilicon 233 -1136 233 -1136 0 3
rlabel polysilicon 240 -1130 240 -1130 0 1
rlabel polysilicon 240 -1136 240 -1136 0 3
rlabel polysilicon 247 -1130 247 -1130 0 1
rlabel polysilicon 247 -1136 247 -1136 0 3
rlabel polysilicon 254 -1130 254 -1130 0 1
rlabel polysilicon 254 -1136 254 -1136 0 3
rlabel polysilicon 261 -1130 261 -1130 0 1
rlabel polysilicon 264 -1130 264 -1130 0 2
rlabel polysilicon 261 -1136 261 -1136 0 3
rlabel polysilicon 264 -1136 264 -1136 0 4
rlabel polysilicon 268 -1130 268 -1130 0 1
rlabel polysilicon 268 -1136 268 -1136 0 3
rlabel polysilicon 275 -1130 275 -1130 0 1
rlabel polysilicon 278 -1130 278 -1130 0 2
rlabel polysilicon 275 -1136 275 -1136 0 3
rlabel polysilicon 278 -1136 278 -1136 0 4
rlabel polysilicon 282 -1130 282 -1130 0 1
rlabel polysilicon 282 -1136 282 -1136 0 3
rlabel polysilicon 289 -1130 289 -1130 0 1
rlabel polysilicon 289 -1136 289 -1136 0 3
rlabel polysilicon 296 -1130 296 -1130 0 1
rlabel polysilicon 296 -1136 296 -1136 0 3
rlabel polysilicon 303 -1136 303 -1136 0 3
rlabel polysilicon 306 -1136 306 -1136 0 4
rlabel polysilicon 310 -1130 310 -1130 0 1
rlabel polysilicon 310 -1136 310 -1136 0 3
rlabel polysilicon 317 -1130 317 -1130 0 1
rlabel polysilicon 320 -1130 320 -1130 0 2
rlabel polysilicon 327 -1136 327 -1136 0 4
rlabel polysilicon 331 -1130 331 -1130 0 1
rlabel polysilicon 331 -1136 331 -1136 0 3
rlabel polysilicon 338 -1130 338 -1130 0 1
rlabel polysilicon 338 -1136 338 -1136 0 3
rlabel polysilicon 345 -1130 345 -1130 0 1
rlabel polysilicon 345 -1136 345 -1136 0 3
rlabel polysilicon 352 -1130 352 -1130 0 1
rlabel polysilicon 352 -1136 352 -1136 0 3
rlabel polysilicon 359 -1130 359 -1130 0 1
rlabel polysilicon 362 -1130 362 -1130 0 2
rlabel polysilicon 369 -1130 369 -1130 0 2
rlabel polysilicon 369 -1136 369 -1136 0 4
rlabel polysilicon 373 -1130 373 -1130 0 1
rlabel polysilicon 373 -1136 373 -1136 0 3
rlabel polysilicon 380 -1130 380 -1130 0 1
rlabel polysilicon 380 -1136 380 -1136 0 3
rlabel polysilicon 387 -1130 387 -1130 0 1
rlabel polysilicon 387 -1136 387 -1136 0 3
rlabel polysilicon 394 -1130 394 -1130 0 1
rlabel polysilicon 394 -1136 394 -1136 0 3
rlabel polysilicon 401 -1130 401 -1130 0 1
rlabel polysilicon 401 -1136 401 -1136 0 3
rlabel polysilicon 408 -1130 408 -1130 0 1
rlabel polysilicon 408 -1136 408 -1136 0 3
rlabel polysilicon 415 -1130 415 -1130 0 1
rlabel polysilicon 415 -1136 415 -1136 0 3
rlabel polysilicon 422 -1130 422 -1130 0 1
rlabel polysilicon 422 -1136 422 -1136 0 3
rlabel polysilicon 429 -1130 429 -1130 0 1
rlabel polysilicon 429 -1136 429 -1136 0 3
rlabel polysilicon 436 -1130 436 -1130 0 1
rlabel polysilicon 436 -1136 436 -1136 0 3
rlabel polysilicon 443 -1130 443 -1130 0 1
rlabel polysilicon 443 -1136 443 -1136 0 3
rlabel polysilicon 478 -1130 478 -1130 0 1
rlabel polysilicon 478 -1136 478 -1136 0 3
rlabel polysilicon 485 -1136 485 -1136 0 3
rlabel polysilicon 54 -1173 54 -1173 0 2
rlabel polysilicon 61 -1179 61 -1179 0 4
rlabel polysilicon 72 -1173 72 -1173 0 1
rlabel polysilicon 72 -1179 72 -1179 0 3
rlabel polysilicon 82 -1173 82 -1173 0 2
rlabel polysilicon 86 -1173 86 -1173 0 1
rlabel polysilicon 86 -1179 86 -1179 0 3
rlabel polysilicon 93 -1173 93 -1173 0 1
rlabel polysilicon 100 -1173 100 -1173 0 1
rlabel polysilicon 100 -1179 100 -1179 0 3
rlabel polysilicon 107 -1173 107 -1173 0 1
rlabel polysilicon 107 -1179 107 -1179 0 3
rlabel polysilicon 114 -1173 114 -1173 0 1
rlabel polysilicon 117 -1173 117 -1173 0 2
rlabel polysilicon 114 -1179 114 -1179 0 3
rlabel polysilicon 121 -1173 121 -1173 0 1
rlabel polysilicon 124 -1173 124 -1173 0 2
rlabel polysilicon 121 -1179 121 -1179 0 3
rlabel polysilicon 124 -1179 124 -1179 0 4
rlabel polysilicon 128 -1173 128 -1173 0 1
rlabel polysilicon 128 -1179 128 -1179 0 3
rlabel polysilicon 135 -1173 135 -1173 0 1
rlabel polysilicon 135 -1179 135 -1179 0 3
rlabel polysilicon 145 -1173 145 -1173 0 2
rlabel polysilicon 149 -1173 149 -1173 0 1
rlabel polysilicon 149 -1179 149 -1179 0 3
rlabel polysilicon 156 -1173 156 -1173 0 1
rlabel polysilicon 156 -1179 156 -1179 0 3
rlabel polysilicon 163 -1173 163 -1173 0 1
rlabel polysilicon 166 -1173 166 -1173 0 2
rlabel polysilicon 170 -1173 170 -1173 0 1
rlabel polysilicon 173 -1173 173 -1173 0 2
rlabel polysilicon 170 -1179 170 -1179 0 3
rlabel polysilicon 177 -1173 177 -1173 0 1
rlabel polysilicon 177 -1179 177 -1179 0 3
rlabel polysilicon 184 -1173 184 -1173 0 1
rlabel polysilicon 184 -1179 184 -1179 0 3
rlabel polysilicon 191 -1173 191 -1173 0 1
rlabel polysilicon 191 -1179 191 -1179 0 3
rlabel polysilicon 198 -1173 198 -1173 0 1
rlabel polysilicon 198 -1179 198 -1179 0 3
rlabel polysilicon 201 -1179 201 -1179 0 4
rlabel polysilicon 205 -1173 205 -1173 0 1
rlabel polysilicon 208 -1173 208 -1173 0 2
rlabel polysilicon 205 -1179 205 -1179 0 3
rlabel polysilicon 208 -1179 208 -1179 0 4
rlabel polysilicon 212 -1173 212 -1173 0 1
rlabel polysilicon 212 -1179 212 -1179 0 3
rlabel polysilicon 219 -1173 219 -1173 0 1
rlabel polysilicon 219 -1179 219 -1179 0 3
rlabel polysilicon 226 -1173 226 -1173 0 1
rlabel polysilicon 226 -1179 226 -1179 0 3
rlabel polysilicon 233 -1173 233 -1173 0 1
rlabel polysilicon 233 -1179 233 -1179 0 3
rlabel polysilicon 240 -1173 240 -1173 0 1
rlabel polysilicon 243 -1173 243 -1173 0 2
rlabel polysilicon 240 -1179 240 -1179 0 3
rlabel polysilicon 250 -1173 250 -1173 0 2
rlabel polysilicon 247 -1179 247 -1179 0 3
rlabel polysilicon 250 -1179 250 -1179 0 4
rlabel polysilicon 254 -1173 254 -1173 0 1
rlabel polysilicon 257 -1179 257 -1179 0 4
rlabel polysilicon 261 -1173 261 -1173 0 1
rlabel polysilicon 264 -1173 264 -1173 0 2
rlabel polysilicon 261 -1179 261 -1179 0 3
rlabel polysilicon 268 -1173 268 -1173 0 1
rlabel polysilicon 268 -1179 268 -1179 0 3
rlabel polysilicon 275 -1173 275 -1173 0 1
rlabel polysilicon 275 -1179 275 -1179 0 3
rlabel polysilicon 282 -1173 282 -1173 0 1
rlabel polysilicon 282 -1179 282 -1179 0 3
rlabel polysilicon 289 -1173 289 -1173 0 1
rlabel polysilicon 289 -1179 289 -1179 0 3
rlabel polysilicon 299 -1173 299 -1173 0 2
rlabel polysilicon 296 -1179 296 -1179 0 3
rlabel polysilicon 306 -1173 306 -1173 0 2
rlabel polysilicon 303 -1179 303 -1179 0 3
rlabel polysilicon 310 -1173 310 -1173 0 1
rlabel polysilicon 310 -1179 310 -1179 0 3
rlabel polysilicon 317 -1173 317 -1173 0 1
rlabel polysilicon 317 -1179 317 -1179 0 3
rlabel polysilicon 324 -1173 324 -1173 0 1
rlabel polysilicon 324 -1179 324 -1179 0 3
rlabel polysilicon 331 -1173 331 -1173 0 1
rlabel polysilicon 331 -1179 331 -1179 0 3
rlabel polysilicon 338 -1173 338 -1173 0 1
rlabel polysilicon 338 -1179 338 -1179 0 3
rlabel polysilicon 345 -1173 345 -1173 0 1
rlabel polysilicon 345 -1179 345 -1179 0 3
rlabel polysilicon 352 -1173 352 -1173 0 1
rlabel polysilicon 352 -1179 352 -1179 0 3
rlabel polysilicon 359 -1173 359 -1173 0 1
rlabel polysilicon 359 -1179 359 -1179 0 3
rlabel polysilicon 366 -1173 366 -1173 0 1
rlabel polysilicon 366 -1179 366 -1179 0 3
rlabel polysilicon 376 -1173 376 -1173 0 2
rlabel polysilicon 376 -1179 376 -1179 0 4
rlabel polysilicon 380 -1173 380 -1173 0 1
rlabel polysilicon 380 -1179 380 -1179 0 3
rlabel polysilicon 387 -1173 387 -1173 0 1
rlabel polysilicon 387 -1179 387 -1179 0 3
rlabel polysilicon 397 -1173 397 -1173 0 2
rlabel polysilicon 401 -1173 401 -1173 0 1
rlabel polysilicon 401 -1179 401 -1179 0 3
rlabel polysilicon 408 -1173 408 -1173 0 1
rlabel polysilicon 65 -1204 65 -1204 0 1
rlabel polysilicon 65 -1210 65 -1210 0 3
rlabel polysilicon 72 -1204 72 -1204 0 1
rlabel polysilicon 72 -1210 72 -1210 0 3
rlabel polysilicon 79 -1204 79 -1204 0 1
rlabel polysilicon 79 -1210 79 -1210 0 3
rlabel polysilicon 89 -1210 89 -1210 0 4
rlabel polysilicon 93 -1204 93 -1204 0 1
rlabel polysilicon 93 -1210 93 -1210 0 3
rlabel polysilicon 100 -1204 100 -1204 0 1
rlabel polysilicon 100 -1210 100 -1210 0 3
rlabel polysilicon 107 -1204 107 -1204 0 1
rlabel polysilicon 107 -1210 107 -1210 0 3
rlabel polysilicon 114 -1204 114 -1204 0 1
rlabel polysilicon 114 -1210 114 -1210 0 3
rlabel polysilicon 121 -1204 121 -1204 0 1
rlabel polysilicon 121 -1210 121 -1210 0 3
rlabel polysilicon 131 -1204 131 -1204 0 2
rlabel polysilicon 128 -1210 128 -1210 0 3
rlabel polysilicon 138 -1204 138 -1204 0 2
rlabel polysilicon 138 -1210 138 -1210 0 4
rlabel polysilicon 142 -1204 142 -1204 0 1
rlabel polysilicon 142 -1210 142 -1210 0 3
rlabel polysilicon 149 -1210 149 -1210 0 3
rlabel polysilicon 156 -1204 156 -1204 0 1
rlabel polysilicon 159 -1210 159 -1210 0 4
rlabel polysilicon 163 -1204 163 -1204 0 1
rlabel polysilicon 163 -1210 163 -1210 0 3
rlabel polysilicon 170 -1204 170 -1204 0 1
rlabel polysilicon 173 -1204 173 -1204 0 2
rlabel polysilicon 177 -1210 177 -1210 0 3
rlabel polysilicon 180 -1210 180 -1210 0 4
rlabel polysilicon 184 -1204 184 -1204 0 1
rlabel polysilicon 187 -1210 187 -1210 0 4
rlabel polysilicon 191 -1204 191 -1204 0 1
rlabel polysilicon 194 -1204 194 -1204 0 2
rlabel polysilicon 191 -1210 191 -1210 0 3
rlabel polysilicon 198 -1204 198 -1204 0 1
rlabel polysilicon 198 -1210 198 -1210 0 3
rlabel polysilicon 208 -1204 208 -1204 0 2
rlabel polysilicon 212 -1204 212 -1204 0 1
rlabel polysilicon 212 -1210 212 -1210 0 3
rlabel polysilicon 219 -1204 219 -1204 0 1
rlabel polysilicon 219 -1210 219 -1210 0 3
rlabel polysilicon 229 -1210 229 -1210 0 4
rlabel polysilicon 233 -1204 233 -1204 0 1
rlabel polysilicon 233 -1210 233 -1210 0 3
rlabel polysilicon 240 -1204 240 -1204 0 1
rlabel polysilicon 240 -1210 240 -1210 0 3
rlabel polysilicon 243 -1210 243 -1210 0 4
rlabel polysilicon 247 -1204 247 -1204 0 1
rlabel polysilicon 247 -1210 247 -1210 0 3
rlabel polysilicon 254 -1204 254 -1204 0 1
rlabel polysilicon 254 -1210 254 -1210 0 3
rlabel polysilicon 261 -1210 261 -1210 0 3
rlabel polysilicon 264 -1210 264 -1210 0 4
rlabel polysilicon 268 -1204 268 -1204 0 1
rlabel polysilicon 268 -1210 268 -1210 0 3
rlabel polysilicon 275 -1204 275 -1204 0 1
rlabel polysilicon 275 -1210 275 -1210 0 3
rlabel polysilicon 282 -1204 282 -1204 0 1
rlabel polysilicon 282 -1210 282 -1210 0 3
rlabel polysilicon 292 -1204 292 -1204 0 2
rlabel polysilicon 292 -1210 292 -1210 0 4
rlabel polysilicon 296 -1204 296 -1204 0 1
rlabel polysilicon 296 -1210 296 -1210 0 3
rlabel polysilicon 303 -1210 303 -1210 0 3
rlabel polysilicon 310 -1204 310 -1204 0 1
rlabel polysilicon 310 -1210 310 -1210 0 3
rlabel polysilicon 317 -1210 317 -1210 0 3
rlabel polysilicon 324 -1204 324 -1204 0 1
rlabel polysilicon 331 -1204 331 -1204 0 1
rlabel polysilicon 331 -1210 331 -1210 0 3
rlabel polysilicon 338 -1204 338 -1204 0 1
rlabel polysilicon 338 -1210 338 -1210 0 3
rlabel polysilicon 345 -1204 345 -1204 0 1
rlabel polysilicon 345 -1210 345 -1210 0 3
rlabel polysilicon 352 -1204 352 -1204 0 1
rlabel polysilicon 352 -1210 352 -1210 0 3
rlabel polysilicon 359 -1204 359 -1204 0 1
rlabel polysilicon 359 -1210 359 -1210 0 3
rlabel polysilicon 366 -1204 366 -1204 0 1
rlabel polysilicon 366 -1210 366 -1210 0 3
rlabel polysilicon 373 -1204 373 -1204 0 1
rlabel polysilicon 373 -1210 373 -1210 0 3
rlabel polysilicon 380 -1204 380 -1204 0 1
rlabel polysilicon 383 -1204 383 -1204 0 2
rlabel polysilicon 383 -1210 383 -1210 0 4
rlabel polysilicon 387 -1204 387 -1204 0 1
rlabel polysilicon 387 -1210 387 -1210 0 3
rlabel polysilicon 394 -1204 394 -1204 0 1
rlabel polysilicon 394 -1210 394 -1210 0 3
rlabel polysilicon 93 -1233 93 -1233 0 1
rlabel polysilicon 93 -1239 93 -1239 0 3
rlabel polysilicon 100 -1239 100 -1239 0 3
rlabel polysilicon 110 -1239 110 -1239 0 4
rlabel polysilicon 114 -1233 114 -1233 0 1
rlabel polysilicon 114 -1239 114 -1239 0 3
rlabel polysilicon 121 -1233 121 -1233 0 1
rlabel polysilicon 128 -1233 128 -1233 0 1
rlabel polysilicon 128 -1239 128 -1239 0 3
rlabel polysilicon 135 -1233 135 -1233 0 1
rlabel polysilicon 135 -1239 135 -1239 0 3
rlabel polysilicon 142 -1233 142 -1233 0 1
rlabel polysilicon 142 -1239 142 -1239 0 3
rlabel polysilicon 152 -1233 152 -1233 0 2
rlabel polysilicon 152 -1239 152 -1239 0 4
rlabel polysilicon 156 -1233 156 -1233 0 1
rlabel polysilicon 156 -1239 156 -1239 0 3
rlabel polysilicon 163 -1233 163 -1233 0 1
rlabel polysilicon 163 -1239 163 -1239 0 3
rlabel polysilicon 170 -1233 170 -1233 0 1
rlabel polysilicon 180 -1233 180 -1233 0 2
rlabel polysilicon 180 -1239 180 -1239 0 4
rlabel polysilicon 184 -1233 184 -1233 0 1
rlabel polysilicon 187 -1239 187 -1239 0 4
rlabel polysilicon 194 -1233 194 -1233 0 2
rlabel polysilicon 191 -1239 191 -1239 0 3
rlabel polysilicon 201 -1239 201 -1239 0 4
rlabel polysilicon 205 -1233 205 -1233 0 1
rlabel polysilicon 205 -1239 205 -1239 0 3
rlabel polysilicon 212 -1233 212 -1233 0 1
rlabel polysilicon 212 -1239 212 -1239 0 3
rlabel polysilicon 219 -1239 219 -1239 0 3
rlabel polysilicon 226 -1233 226 -1233 0 1
rlabel polysilicon 226 -1239 226 -1239 0 3
rlabel polysilicon 233 -1233 233 -1233 0 1
rlabel polysilicon 233 -1239 233 -1239 0 3
rlabel polysilicon 240 -1233 240 -1233 0 1
rlabel polysilicon 240 -1239 240 -1239 0 3
rlabel polysilicon 247 -1233 247 -1233 0 1
rlabel polysilicon 247 -1239 247 -1239 0 3
rlabel polysilicon 254 -1233 254 -1233 0 1
rlabel polysilicon 261 -1233 261 -1233 0 1
rlabel polysilicon 261 -1239 261 -1239 0 3
rlabel polysilicon 268 -1233 268 -1233 0 1
rlabel polysilicon 275 -1233 275 -1233 0 1
rlabel polysilicon 275 -1239 275 -1239 0 3
rlabel polysilicon 282 -1233 282 -1233 0 1
rlabel polysilicon 282 -1239 282 -1239 0 3
rlabel polysilicon 289 -1233 289 -1233 0 1
rlabel polysilicon 289 -1239 289 -1239 0 3
rlabel polysilicon 296 -1233 296 -1233 0 1
rlabel polysilicon 299 -1239 299 -1239 0 4
rlabel polysilicon 306 -1239 306 -1239 0 4
rlabel polysilicon 310 -1233 310 -1233 0 1
rlabel polysilicon 310 -1239 310 -1239 0 3
rlabel polysilicon 317 -1233 317 -1233 0 1
rlabel polysilicon 317 -1239 317 -1239 0 3
rlabel polysilicon 324 -1233 324 -1233 0 1
rlabel polysilicon 324 -1239 324 -1239 0 3
rlabel polysilicon 331 -1233 331 -1233 0 1
rlabel polysilicon 331 -1239 331 -1239 0 3
rlabel polysilicon 348 -1239 348 -1239 0 4
rlabel polysilicon 352 -1233 352 -1233 0 1
rlabel polysilicon 352 -1239 352 -1239 0 3
rlabel polysilicon 380 -1233 380 -1233 0 1
rlabel polysilicon 380 -1239 380 -1239 0 3
rlabel polysilicon 5 -1260 5 -1260 0 4
rlabel polysilicon 75 -1260 75 -1260 0 4
rlabel polysilicon 82 -1254 82 -1254 0 2
rlabel polysilicon 79 -1260 79 -1260 0 3
rlabel polysilicon 86 -1254 86 -1254 0 1
rlabel polysilicon 86 -1260 86 -1260 0 3
rlabel polysilicon 100 -1254 100 -1254 0 1
rlabel polysilicon 100 -1260 100 -1260 0 3
rlabel polysilicon 107 -1254 107 -1254 0 1
rlabel polysilicon 107 -1260 107 -1260 0 3
rlabel polysilicon 117 -1254 117 -1254 0 2
rlabel polysilicon 114 -1260 114 -1260 0 3
rlabel polysilicon 121 -1254 121 -1254 0 1
rlabel polysilicon 121 -1260 121 -1260 0 3
rlabel polysilicon 128 -1254 128 -1254 0 1
rlabel polysilicon 128 -1260 128 -1260 0 3
rlabel polysilicon 135 -1254 135 -1254 0 1
rlabel polysilicon 135 -1260 135 -1260 0 3
rlabel polysilicon 145 -1260 145 -1260 0 4
rlabel polysilicon 149 -1254 149 -1254 0 1
rlabel polysilicon 149 -1260 149 -1260 0 3
rlabel polysilicon 156 -1254 156 -1254 0 1
rlabel polysilicon 163 -1260 163 -1260 0 3
rlabel polysilicon 166 -1260 166 -1260 0 4
rlabel polysilicon 173 -1254 173 -1254 0 2
rlabel polysilicon 173 -1260 173 -1260 0 4
rlabel polysilicon 177 -1254 177 -1254 0 1
rlabel polysilicon 177 -1260 177 -1260 0 3
rlabel polysilicon 184 -1260 184 -1260 0 3
rlabel polysilicon 191 -1254 191 -1254 0 1
rlabel polysilicon 191 -1260 191 -1260 0 3
rlabel polysilicon 198 -1254 198 -1254 0 1
rlabel polysilicon 205 -1254 205 -1254 0 1
rlabel polysilicon 205 -1260 205 -1260 0 3
rlabel polysilicon 215 -1254 215 -1254 0 2
rlabel polysilicon 219 -1254 219 -1254 0 1
rlabel polysilicon 219 -1260 219 -1260 0 3
rlabel polysilicon 226 -1254 226 -1254 0 1
rlabel polysilicon 233 -1254 233 -1254 0 1
rlabel polysilicon 233 -1260 233 -1260 0 3
rlabel polysilicon 240 -1254 240 -1254 0 1
rlabel polysilicon 240 -1260 240 -1260 0 3
rlabel polysilicon 247 -1254 247 -1254 0 1
rlabel polysilicon 254 -1254 254 -1254 0 1
rlabel polysilicon 254 -1260 254 -1260 0 3
rlabel polysilicon 261 -1254 261 -1254 0 1
rlabel polysilicon 261 -1260 261 -1260 0 3
rlabel polysilicon 268 -1254 268 -1254 0 1
rlabel polysilicon 268 -1260 268 -1260 0 3
rlabel polysilicon 278 -1254 278 -1254 0 2
rlabel polysilicon 275 -1260 275 -1260 0 3
rlabel polysilicon 278 -1260 278 -1260 0 4
rlabel polysilicon 285 -1254 285 -1254 0 2
rlabel polysilicon 289 -1254 289 -1254 0 1
rlabel polysilicon 296 -1254 296 -1254 0 1
rlabel polysilicon 296 -1260 296 -1260 0 3
rlabel polysilicon 303 -1254 303 -1254 0 1
rlabel polysilicon 303 -1260 303 -1260 0 3
rlabel polysilicon 320 -1254 320 -1254 0 2
rlabel polysilicon 320 -1260 320 -1260 0 4
rlabel polysilicon 324 -1254 324 -1254 0 1
rlabel polysilicon 324 -1260 324 -1260 0 3
rlabel polysilicon 380 -1254 380 -1254 0 1
rlabel polysilicon 380 -1260 380 -1260 0 3
rlabel polysilicon 5 -1269 5 -1269 0 2
rlabel polysilicon 86 -1269 86 -1269 0 1
rlabel polysilicon 86 -1275 86 -1275 0 3
rlabel polysilicon 96 -1275 96 -1275 0 4
rlabel polysilicon 107 -1269 107 -1269 0 1
rlabel polysilicon 107 -1275 107 -1275 0 3
rlabel polysilicon 117 -1269 117 -1269 0 2
rlabel polysilicon 117 -1275 117 -1275 0 4
rlabel polysilicon 121 -1269 121 -1269 0 1
rlabel polysilicon 121 -1275 121 -1275 0 3
rlabel polysilicon 128 -1275 128 -1275 0 3
rlabel polysilicon 135 -1269 135 -1269 0 1
rlabel polysilicon 135 -1275 135 -1275 0 3
rlabel polysilicon 145 -1275 145 -1275 0 4
rlabel polysilicon 149 -1269 149 -1269 0 1
rlabel polysilicon 149 -1275 149 -1275 0 3
rlabel polysilicon 156 -1275 156 -1275 0 3
rlabel polysilicon 159 -1275 159 -1275 0 4
rlabel polysilicon 166 -1275 166 -1275 0 4
rlabel polysilicon 170 -1269 170 -1269 0 1
rlabel polysilicon 184 -1269 184 -1269 0 1
rlabel polysilicon 205 -1269 205 -1269 0 1
rlabel polysilicon 215 -1269 215 -1269 0 2
rlabel polysilicon 219 -1275 219 -1275 0 3
rlabel polysilicon 226 -1269 226 -1269 0 1
rlabel polysilicon 226 -1275 226 -1275 0 3
rlabel polysilicon 233 -1269 233 -1269 0 1
rlabel polysilicon 240 -1269 240 -1269 0 1
rlabel polysilicon 271 -1269 271 -1269 0 2
rlabel polysilicon 275 -1269 275 -1269 0 1
rlabel polysilicon 275 -1275 275 -1275 0 3
rlabel polysilicon 282 -1275 282 -1275 0 3
rlabel polysilicon 299 -1275 299 -1275 0 4
rlabel polysilicon 303 -1269 303 -1269 0 1
rlabel polysilicon 303 -1275 303 -1275 0 3
rlabel polysilicon 383 -1275 383 -1275 0 4
rlabel polysilicon 387 -1269 387 -1269 0 1
rlabel polysilicon 387 -1275 387 -1275 0 3
rlabel metal2 135 1 135 1 0 net=1299
rlabel metal2 145 1 145 1 0 net=616
rlabel metal2 184 1 184 1 0 net=608
rlabel metal2 212 1 212 1 0 net=2777
rlabel metal2 135 -10 135 -10 0 net=1300
rlabel metal2 156 -10 156 -10 0 net=2031
rlabel metal2 191 -10 191 -10 0 net=2749
rlabel metal2 208 -10 208 -10 0 net=2778
rlabel metal2 254 -10 254 -10 0 net=1853
rlabel metal2 254 -10 254 -10 0 net=1853
rlabel metal2 257 -10 257 -10 0 net=179
rlabel metal2 142 -12 142 -12 0 net=170
rlabel metal2 142 -12 142 -12 0 net=170
rlabel metal2 149 -12 149 -12 0 net=2607
rlabel metal2 177 -12 177 -12 0 net=421
rlabel metal2 212 -12 212 -12 0 net=1763
rlabel metal2 184 -14 184 -14 0 net=1965
rlabel metal2 149 -25 149 -25 0 net=2608
rlabel metal2 170 -25 170 -25 0 net=1966
rlabel metal2 187 -25 187 -25 0 net=1317
rlabel metal2 198 -25 198 -25 0 net=2751
rlabel metal2 229 -25 229 -25 0 net=2097
rlabel metal2 268 -25 268 -25 0 net=319
rlabel metal2 310 -25 310 -25 0 net=2521
rlabel metal2 310 -25 310 -25 0 net=2521
rlabel metal2 341 -25 341 -25 0 net=2813
rlabel metal2 145 -27 145 -27 0 net=1661
rlabel metal2 156 -27 156 -27 0 net=2032
rlabel metal2 177 -27 177 -27 0 net=283
rlabel metal2 243 -27 243 -27 0 net=2993
rlabel metal2 254 -27 254 -27 0 net=1855
rlabel metal2 254 -27 254 -27 0 net=1855
rlabel metal2 163 -29 163 -29 0 net=1359
rlabel metal2 163 -29 163 -29 0 net=1359
rlabel metal2 201 -29 201 -29 0 net=1764
rlabel metal2 205 -31 205 -31 0 net=1529
rlabel metal2 212 -33 212 -33 0 net=2017
rlabel metal2 51 -44 51 -44 0 net=591
rlabel metal2 72 -44 72 -44 0 net=1401
rlabel metal2 100 -44 100 -44 0 net=2309
rlabel metal2 100 -44 100 -44 0 net=2309
rlabel metal2 138 -44 138 -44 0 net=1662
rlabel metal2 156 -44 156 -44 0 net=674
rlabel metal2 201 -44 201 -44 0 net=2752
rlabel metal2 233 -44 233 -44 0 net=1831
rlabel metal2 233 -44 233 -44 0 net=1831
rlabel metal2 236 -44 236 -44 0 net=2994
rlabel metal2 282 -44 282 -44 0 net=2545
rlabel metal2 310 -44 310 -44 0 net=2523
rlabel metal2 310 -44 310 -44 0 net=2523
rlabel metal2 338 -44 338 -44 0 net=2299
rlabel metal2 338 -44 338 -44 0 net=2299
rlabel metal2 345 -44 345 -44 0 net=2815
rlabel metal2 359 -44 359 -44 0 net=2413
rlabel metal2 142 -46 142 -46 0 net=1369
rlabel metal2 208 -46 208 -46 0 net=2018
rlabel metal2 240 -46 240 -46 0 net=1530
rlabel metal2 247 -46 247 -46 0 net=2099
rlabel metal2 345 -46 345 -46 0 net=513
rlabel metal2 163 -48 163 -48 0 net=1360
rlabel metal2 191 -48 191 -48 0 net=1319
rlabel metal2 240 -48 240 -48 0 net=2741
rlabel metal2 170 -50 170 -50 0 net=963
rlabel metal2 177 -52 177 -52 0 net=445
rlabel metal2 194 -52 194 -52 0 net=1569
rlabel metal2 261 -52 261 -52 0 net=2019
rlabel metal2 163 -54 163 -54 0 net=953
rlabel metal2 187 -54 187 -54 0 net=1255
rlabel metal2 254 -54 254 -54 0 net=1857
rlabel metal2 226 -56 226 -56 0 net=1851
rlabel metal2 26 -67 26 -67 0 net=527
rlabel metal2 26 -67 26 -67 0 net=527
rlabel metal2 51 -67 51 -67 0 net=1402
rlabel metal2 79 -67 79 -67 0 net=1371
rlabel metal2 149 -67 149 -67 0 net=221
rlabel metal2 194 -67 194 -67 0 net=1256
rlabel metal2 219 -67 219 -67 0 net=1571
rlabel metal2 282 -67 282 -67 0 net=465
rlabel metal2 58 -69 58 -69 0 net=2531
rlabel metal2 149 -69 149 -69 0 net=1011
rlabel metal2 247 -69 247 -69 0 net=2101
rlabel metal2 310 -69 310 -69 0 net=2524
rlabel metal2 320 -69 320 -69 0 net=2171
rlabel metal2 338 -69 338 -69 0 net=2300
rlabel metal2 366 -69 366 -69 0 net=2415
rlabel metal2 366 -69 366 -69 0 net=2415
rlabel metal2 65 -71 65 -71 0 net=965
rlabel metal2 198 -71 198 -71 0 net=1591
rlabel metal2 289 -71 289 -71 0 net=2547
rlabel metal2 345 -71 345 -71 0 net=2817
rlabel metal2 72 -73 72 -73 0 net=1929
rlabel metal2 93 -73 93 -73 0 net=522
rlabel metal2 156 -73 156 -73 0 net=1539
rlabel metal2 201 -73 201 -73 0 net=1852
rlabel metal2 257 -73 257 -73 0 net=2375
rlabel metal2 93 -75 93 -75 0 net=1179
rlabel metal2 229 -75 229 -75 0 net=2717
rlabel metal2 96 -77 96 -77 0 net=2310
rlabel metal2 103 -77 103 -77 0 net=1301
rlabel metal2 121 -77 121 -77 0 net=1533
rlabel metal2 254 -77 254 -77 0 net=1858
rlabel metal2 278 -77 278 -77 0 net=1843
rlabel metal2 107 -79 107 -79 0 net=1021
rlabel metal2 163 -79 163 -79 0 net=955
rlabel metal2 163 -79 163 -79 0 net=955
rlabel metal2 205 -79 205 -79 0 net=1321
rlabel metal2 226 -79 226 -79 0 net=1715
rlabel metal2 296 -79 296 -79 0 net=2743
rlabel metal2 128 -81 128 -81 0 net=2333
rlabel metal2 205 -81 205 -81 0 net=1497
rlabel metal2 212 -83 212 -83 0 net=1093
rlabel metal2 261 -83 261 -83 0 net=2021
rlabel metal2 208 -85 208 -85 0 net=1389
rlabel metal2 233 -87 233 -87 0 net=1832
rlabel metal2 58 -98 58 -98 0 net=2532
rlabel metal2 173 -98 173 -98 0 net=1390
rlabel metal2 345 -98 345 -98 0 net=2819
rlabel metal2 345 -98 345 -98 0 net=2819
rlabel metal2 352 -98 352 -98 0 net=1845
rlabel metal2 65 -100 65 -100 0 net=966
rlabel metal2 184 -100 184 -100 0 net=1095
rlabel metal2 236 -100 236 -100 0 net=1592
rlabel metal2 366 -100 366 -100 0 net=2416
rlabel metal2 376 -100 376 -100 0 net=2259
rlabel metal2 72 -102 72 -102 0 net=1930
rlabel metal2 107 -102 107 -102 0 net=1022
rlabel metal2 205 -102 205 -102 0 net=1322
rlabel metal2 243 -102 243 -102 0 net=2744
rlabel metal2 100 -104 100 -104 0 net=1303
rlabel metal2 135 -104 135 -104 0 net=869
rlabel metal2 187 -104 187 -104 0 net=2102
rlabel metal2 324 -104 324 -104 0 net=2377
rlabel metal2 107 -106 107 -106 0 net=1535
rlabel metal2 145 -106 145 -106 0 net=471
rlabel metal2 198 -106 198 -106 0 net=1237
rlabel metal2 338 -106 338 -106 0 net=2423
rlabel metal2 86 -108 86 -108 0 net=2551
rlabel metal2 142 -108 142 -108 0 net=262
rlabel metal2 149 -108 149 -108 0 net=1012
rlabel metal2 236 -108 236 -108 0 net=2009
rlabel metal2 79 -110 79 -110 0 net=1372
rlabel metal2 149 -110 149 -110 0 net=1541
rlabel metal2 163 -110 163 -110 0 net=957
rlabel metal2 247 -110 247 -110 0 net=2022
rlabel metal2 93 -112 93 -112 0 net=1180
rlabel metal2 163 -112 163 -112 0 net=1503
rlabel metal2 250 -112 250 -112 0 net=1827
rlabel metal2 93 -114 93 -114 0 net=2335
rlabel metal2 177 -114 177 -114 0 net=268
rlabel metal2 254 -114 254 -114 0 net=2718
rlabel metal2 128 -116 128 -116 0 net=1601
rlabel metal2 191 -116 191 -116 0 net=2548
rlabel metal2 317 -116 317 -116 0 net=2173
rlabel metal2 191 -118 191 -118 0 net=1572
rlabel metal2 310 -118 310 -118 0 net=2947
rlabel metal2 194 -120 194 -120 0 net=2467
rlabel metal2 254 -120 254 -120 0 net=1547
rlabel metal2 205 -122 205 -122 0 net=1507
rlabel metal2 208 -124 208 -124 0 net=710
rlabel metal2 208 -126 208 -126 0 net=1498
rlabel metal2 219 -128 219 -128 0 net=1653
rlabel metal2 257 -128 257 -128 0 net=1716
rlabel metal2 289 -130 289 -130 0 net=2925
rlabel metal2 65 -141 65 -141 0 net=1097
rlabel metal2 191 -141 191 -141 0 net=977
rlabel metal2 380 -141 380 -141 0 net=1847
rlabel metal2 93 -143 93 -143 0 net=2336
rlabel metal2 142 -143 142 -143 0 net=751
rlabel metal2 170 -143 170 -143 0 net=2468
rlabel metal2 243 -143 243 -143 0 net=2961
rlabel metal2 93 -145 93 -145 0 net=2735
rlabel metal2 121 -145 121 -145 0 net=1543
rlabel metal2 163 -145 163 -145 0 net=1505
rlabel metal2 184 -145 184 -145 0 net=1063
rlabel metal2 264 -145 264 -145 0 net=2549
rlabel metal2 380 -145 380 -145 0 net=2921
rlabel metal2 401 -145 401 -145 0 net=2260
rlabel metal2 72 -147 72 -147 0 net=1567
rlabel metal2 152 -147 152 -147 0 net=671
rlabel metal2 205 -147 205 -147 0 net=958
rlabel metal2 226 -147 226 -147 0 net=1439
rlabel metal2 275 -147 275 -147 0 net=1509
rlabel metal2 275 -147 275 -147 0 net=1509
rlabel metal2 289 -147 289 -147 0 net=3043
rlabel metal2 86 -149 86 -149 0 net=2552
rlabel metal2 177 -149 177 -149 0 net=1177
rlabel metal2 233 -149 233 -149 0 net=1549
rlabel metal2 289 -149 289 -149 0 net=1829
rlabel metal2 310 -149 310 -149 0 net=2174
rlabel metal2 331 -149 331 -149 0 net=2949
rlabel metal2 394 -149 394 -149 0 net=2425
rlabel metal2 86 -151 86 -151 0 net=1603
rlabel metal2 229 -151 229 -151 0 net=1795
rlabel metal2 285 -151 285 -151 0 net=1577
rlabel metal2 317 -151 317 -151 0 net=663
rlabel metal2 107 -153 107 -153 0 net=1536
rlabel metal2 331 -153 331 -153 0 net=1721
rlabel metal2 366 -153 366 -153 0 net=2379
rlabel metal2 107 -155 107 -155 0 net=871
rlabel metal2 142 -155 142 -155 0 net=223
rlabel metal2 324 -155 324 -155 0 net=2011
rlabel metal2 100 -157 100 -157 0 net=1304
rlabel metal2 219 -157 219 -157 0 net=1655
rlabel metal2 341 -157 341 -157 0 net=2820
rlabel metal2 100 -159 100 -159 0 net=1239
rlabel metal2 303 -159 303 -159 0 net=2927
rlabel metal2 128 -161 128 -161 0 net=565
rlabel metal2 247 -161 247 -161 0 net=1993
rlabel metal2 198 -163 198 -163 0 net=1563
rlabel metal2 247 -165 247 -165 0 net=309
rlabel metal2 23 -176 23 -176 0 net=1257
rlabel metal2 72 -176 72 -176 0 net=1568
rlabel metal2 205 -176 205 -176 0 net=1215
rlabel metal2 219 -176 219 -176 0 net=1994
rlabel metal2 313 -176 313 -176 0 net=2550
rlabel metal2 387 -176 387 -176 0 net=1848
rlabel metal2 411 -176 411 -176 0 net=2779
rlabel metal2 37 -178 37 -178 0 net=1871
rlabel metal2 261 -178 261 -178 0 net=1441
rlabel metal2 261 -178 261 -178 0 net=1441
rlabel metal2 285 -178 285 -178 0 net=1722
rlabel metal2 341 -178 341 -178 0 net=2877
rlabel metal2 44 -180 44 -180 0 net=1385
rlabel metal2 82 -180 82 -180 0 net=611
rlabel metal2 149 -180 149 -180 0 net=752
rlabel metal2 170 -180 170 -180 0 net=1506
rlabel metal2 184 -180 184 -180 0 net=1065
rlabel metal2 184 -180 184 -180 0 net=1065
rlabel metal2 191 -180 191 -180 0 net=979
rlabel metal2 236 -180 236 -180 0 net=264
rlabel metal2 296 -180 296 -180 0 net=1579
rlabel metal2 317 -180 317 -180 0 net=2933
rlabel metal2 51 -182 51 -182 0 net=873
rlabel metal2 114 -182 114 -182 0 net=1605
rlabel metal2 114 -182 114 -182 0 net=1605
rlabel metal2 128 -182 128 -182 0 net=767
rlabel metal2 198 -182 198 -182 0 net=1550
rlabel metal2 240 -182 240 -182 0 net=1830
rlabel metal2 303 -182 303 -182 0 net=1657
rlabel metal2 352 -182 352 -182 0 net=2013
rlabel metal2 380 -182 380 -182 0 net=2923
rlabel metal2 394 -182 394 -182 0 net=2381
rlabel metal2 65 -184 65 -184 0 net=1099
rlabel metal2 243 -184 243 -184 0 net=1987
rlabel metal2 401 -184 401 -184 0 net=2426
rlabel metal2 72 -186 72 -186 0 net=1663
rlabel metal2 86 -186 86 -186 0 net=1604
rlabel metal2 156 -186 156 -186 0 net=278
rlabel metal2 247 -186 247 -186 0 net=1615
rlabel metal2 359 -186 359 -186 0 net=2951
rlabel metal2 415 -186 415 -186 0 net=2963
rlabel metal2 65 -188 65 -188 0 net=572
rlabel metal2 93 -188 93 -188 0 net=2736
rlabel metal2 177 -188 177 -188 0 net=757
rlabel metal2 268 -188 268 -188 0 net=1564
rlabel metal2 373 -188 373 -188 0 net=2023
rlabel metal2 415 -188 415 -188 0 net=2043
rlabel metal2 100 -190 100 -190 0 net=1240
rlabel metal2 275 -190 275 -190 0 net=1511
rlabel metal2 320 -190 320 -190 0 net=2721
rlabel metal2 422 -190 422 -190 0 net=3045
rlabel metal2 96 -192 96 -192 0 net=907
rlabel metal2 107 -192 107 -192 0 net=1679
rlabel metal2 191 -192 191 -192 0 net=1027
rlabel metal2 268 -192 268 -192 0 net=2133
rlabel metal2 121 -194 121 -194 0 net=1544
rlabel metal2 159 -194 159 -194 0 net=1105
rlabel metal2 285 -194 285 -194 0 net=1595
rlabel metal2 324 -194 324 -194 0 net=2657
rlabel metal2 121 -196 121 -196 0 net=1133
rlabel metal2 138 -196 138 -196 0 net=1033
rlabel metal2 198 -196 198 -196 0 net=1178
rlabel metal2 135 -198 135 -198 0 net=193
rlabel metal2 163 -198 163 -198 0 net=1619
rlabel metal2 30 -200 30 -200 0 net=1995
rlabel metal2 205 -200 205 -200 0 net=2928
rlabel metal2 254 -202 254 -202 0 net=1797
rlabel metal2 23 -215 23 -215 0 net=1258
rlabel metal2 100 -215 100 -215 0 net=908
rlabel metal2 152 -215 152 -215 0 net=3046
rlabel metal2 457 -215 457 -215 0 net=2879
rlabel metal2 541 -215 541 -215 0 net=2653
rlabel metal2 30 -217 30 -217 0 net=1996
rlabel metal2 215 -217 215 -217 0 net=234
rlabel metal2 380 -217 380 -217 0 net=1989
rlabel metal2 380 -217 380 -217 0 net=1989
rlabel metal2 408 -217 408 -217 0 net=2583
rlabel metal2 485 -217 485 -217 0 net=2569
rlabel metal2 37 -219 37 -219 0 net=1872
rlabel metal2 156 -219 156 -219 0 net=759
rlabel metal2 184 -219 184 -219 0 net=1067
rlabel metal2 226 -219 226 -219 0 net=1100
rlabel metal2 271 -219 271 -219 0 net=2952
rlabel metal2 422 -219 422 -219 0 net=2135
rlabel metal2 422 -219 422 -219 0 net=2135
rlabel metal2 436 -219 436 -219 0 net=2781
rlabel metal2 37 -221 37 -221 0 net=2519
rlabel metal2 149 -221 149 -221 0 net=721
rlabel metal2 191 -221 191 -221 0 net=1658
rlabel metal2 317 -221 317 -221 0 net=1512
rlabel metal2 345 -221 345 -221 0 net=1799
rlabel metal2 44 -223 44 -223 0 net=1386
rlabel metal2 65 -223 65 -223 0 net=1664
rlabel metal2 100 -223 100 -223 0 net=1607
rlabel metal2 142 -223 142 -223 0 net=322
rlabel metal2 229 -223 229 -223 0 net=2924
rlabel metal2 429 -223 429 -223 0 net=2383
rlabel metal2 450 -223 450 -223 0 net=2273
rlabel metal2 44 -225 44 -225 0 net=2959
rlabel metal2 107 -225 107 -225 0 net=1680
rlabel metal2 247 -225 247 -225 0 net=1029
rlabel metal2 247 -225 247 -225 0 net=1029
rlabel metal2 261 -225 261 -225 0 net=1443
rlabel metal2 299 -225 299 -225 0 net=2722
rlabel metal2 464 -225 464 -225 0 net=2935
rlabel metal2 51 -227 51 -227 0 net=874
rlabel metal2 159 -227 159 -227 0 net=122
rlabel metal2 236 -227 236 -227 0 net=1765
rlabel metal2 275 -227 275 -227 0 net=1106
rlabel metal2 327 -227 327 -227 0 net=2797
rlabel metal2 443 -227 443 -227 0 net=2965
rlabel metal2 58 -229 58 -229 0 net=783
rlabel metal2 240 -229 240 -229 0 net=1216
rlabel metal2 275 -229 275 -229 0 net=1617
rlabel metal2 338 -229 338 -229 0 net=3041
rlabel metal2 65 -231 65 -231 0 net=769
rlabel metal2 163 -231 163 -231 0 net=1620
rlabel metal2 205 -231 205 -231 0 net=1209
rlabel metal2 285 -231 285 -231 0 net=1873
rlabel metal2 51 -233 51 -233 0 net=1723
rlabel metal2 219 -233 219 -233 0 net=981
rlabel metal2 306 -233 306 -233 0 net=2005
rlabel metal2 79 -235 79 -235 0 net=1483
rlabel metal2 142 -235 142 -235 0 net=1289
rlabel metal2 310 -235 310 -235 0 net=1581
rlabel metal2 331 -235 331 -235 0 net=2791
rlabel metal2 86 -237 86 -237 0 net=959
rlabel metal2 166 -237 166 -237 0 net=1379
rlabel metal2 198 -237 198 -237 0 net=659
rlabel metal2 289 -237 289 -237 0 net=1597
rlabel metal2 338 -237 338 -237 0 net=2599
rlabel metal2 93 -239 93 -239 0 net=1135
rlabel metal2 135 -239 135 -239 0 net=1129
rlabel metal2 352 -239 352 -239 0 net=2015
rlabel metal2 89 -241 89 -241 0 net=188
rlabel metal2 170 -241 170 -241 0 net=1034
rlabel metal2 355 -241 355 -241 0 net=2361
rlabel metal2 170 -243 170 -243 0 net=1777
rlabel metal2 366 -243 366 -243 0 net=2025
rlabel metal2 208 -245 208 -245 0 net=2658
rlabel metal2 394 -245 394 -245 0 net=2045
rlabel metal2 243 -247 243 -247 0 net=1805
rlabel metal2 282 -249 282 -249 0 net=2111
rlabel metal2 282 -251 282 -251 0 net=2311
rlabel metal2 37 -262 37 -262 0 net=2520
rlabel metal2 240 -262 240 -262 0 net=1767
rlabel metal2 282 -262 282 -262 0 net=2016
rlabel metal2 443 -262 443 -262 0 net=2312
rlabel metal2 562 -262 562 -262 0 net=2237
rlabel metal2 37 -264 37 -264 0 net=2865
rlabel metal2 142 -264 142 -264 0 net=1069
rlabel metal2 285 -264 285 -264 0 net=1444
rlabel metal2 303 -264 303 -264 0 net=1582
rlabel metal2 320 -264 320 -264 0 net=1800
rlabel metal2 527 -264 527 -264 0 net=529
rlabel metal2 44 -266 44 -266 0 net=2960
rlabel metal2 152 -266 152 -266 0 net=1639
rlabel metal2 296 -266 296 -266 0 net=2137
rlabel metal2 464 -266 464 -266 0 net=2967
rlabel metal2 65 -268 65 -268 0 net=770
rlabel metal2 156 -268 156 -268 0 net=761
rlabel metal2 156 -268 156 -268 0 net=761
rlabel metal2 163 -268 163 -268 0 net=1291
rlabel metal2 306 -268 306 -268 0 net=3042
rlabel metal2 65 -270 65 -270 0 net=2305
rlabel metal2 145 -270 145 -270 0 net=1351
rlabel metal2 310 -270 310 -270 0 net=1599
rlabel metal2 310 -270 310 -270 0 net=1599
rlabel metal2 324 -270 324 -270 0 net=1991
rlabel metal2 383 -270 383 -270 0 net=2983
rlabel metal2 75 -272 75 -272 0 net=684
rlabel metal2 170 -272 170 -272 0 net=1381
rlabel metal2 198 -272 198 -272 0 net=1779
rlabel metal2 331 -272 331 -272 0 net=2026
rlabel metal2 373 -272 373 -272 0 net=1875
rlabel metal2 373 -272 373 -272 0 net=1875
rlabel metal2 408 -272 408 -272 0 net=2799
rlabel metal2 86 -274 86 -274 0 net=960
rlabel metal2 149 -274 149 -274 0 net=1057
rlabel metal2 289 -274 289 -274 0 net=2007
rlabel metal2 408 -274 408 -274 0 net=2113
rlabel metal2 422 -274 422 -274 0 net=2363
rlabel metal2 485 -274 485 -274 0 net=2571
rlabel metal2 485 -274 485 -274 0 net=2571
rlabel metal2 492 -274 492 -274 0 net=2793
rlabel metal2 492 -274 492 -274 0 net=2793
rlabel metal2 499 -274 499 -274 0 net=2881
rlabel metal2 86 -276 86 -276 0 net=711
rlabel metal2 173 -276 173 -276 0 net=2213
rlabel metal2 226 -276 226 -276 0 net=1211
rlabel metal2 334 -276 334 -276 0 net=2584
rlabel metal2 520 -276 520 -276 0 net=2655
rlabel metal2 79 -278 79 -278 0 net=1485
rlabel metal2 338 -278 338 -278 0 net=2477
rlabel metal2 394 -278 394 -278 0 net=2047
rlabel metal2 93 -280 93 -280 0 net=1136
rlabel metal2 191 -280 191 -280 0 net=502
rlabel metal2 345 -280 345 -280 0 net=2936
rlabel metal2 96 -282 96 -282 0 net=117
rlabel metal2 208 -282 208 -282 0 net=1618
rlabel metal2 317 -282 317 -282 0 net=2737
rlabel metal2 100 -284 100 -284 0 net=1609
rlabel metal2 275 -284 275 -284 0 net=1807
rlabel metal2 362 -284 362 -284 0 net=175
rlabel metal2 415 -284 415 -284 0 net=2275
rlabel metal2 471 -284 471 -284 0 net=2783
rlabel metal2 51 -286 51 -286 0 net=1725
rlabel metal2 107 -286 107 -286 0 net=1131
rlabel metal2 243 -286 243 -286 0 net=2389
rlabel metal2 457 -286 457 -286 0 net=2601
rlabel metal2 51 -288 51 -288 0 net=2559
rlabel metal2 135 -288 135 -288 0 net=1139
rlabel metal2 205 -288 205 -288 0 net=2419
rlabel metal2 72 -290 72 -290 0 net=1631
rlabel metal2 184 -290 184 -290 0 net=723
rlabel metal2 348 -290 348 -290 0 net=2661
rlabel metal2 429 -290 429 -290 0 net=2385
rlabel metal2 443 -290 443 -290 0 net=2301
rlabel metal2 58 -292 58 -292 0 net=785
rlabel metal2 303 -292 303 -292 0 net=2645
rlabel metal2 177 -294 177 -294 0 net=1031
rlabel metal2 352 -294 352 -294 0 net=2057
rlabel metal2 247 -296 247 -296 0 net=982
rlabel metal2 334 -296 334 -296 0 net=1773
rlabel metal2 79 -298 79 -298 0 net=1197
rlabel metal2 9 -309 9 -309 0 net=2481
rlabel metal2 93 -309 93 -309 0 net=1059
rlabel metal2 177 -309 177 -309 0 net=1032
rlabel metal2 334 -309 334 -309 0 net=500
rlabel metal2 366 -309 366 -309 0 net=2784
rlabel metal2 485 -309 485 -309 0 net=2573
rlabel metal2 485 -309 485 -309 0 net=2573
rlabel metal2 520 -309 520 -309 0 net=2656
rlabel metal2 548 -309 548 -309 0 net=2985
rlabel metal2 16 -311 16 -311 0 net=1809
rlabel metal2 285 -311 285 -311 0 net=1600
rlabel metal2 334 -311 334 -311 0 net=2238
rlabel metal2 23 -313 23 -313 0 net=2719
rlabel metal2 100 -313 100 -313 0 net=1726
rlabel metal2 338 -313 338 -313 0 net=2420
rlabel metal2 464 -313 464 -313 0 net=2794
rlabel metal2 527 -313 527 -313 0 net=2801
rlabel metal2 30 -315 30 -315 0 net=805
rlabel metal2 51 -315 51 -315 0 net=2560
rlabel metal2 65 -315 65 -315 0 net=2306
rlabel metal2 250 -315 250 -315 0 net=2503
rlabel metal2 471 -315 471 -315 0 net=2602
rlabel metal2 37 -317 37 -317 0 net=2866
rlabel metal2 240 -317 240 -317 0 net=1768
rlabel metal2 285 -317 285 -317 0 net=3037
rlabel metal2 44 -319 44 -319 0 net=1641
rlabel metal2 240 -319 240 -319 0 net=2364
rlabel metal2 429 -319 429 -319 0 net=2387
rlabel metal2 51 -321 51 -321 0 net=1141
rlabel metal2 180 -321 180 -321 0 net=861
rlabel metal2 289 -321 289 -321 0 net=2008
rlabel metal2 289 -321 289 -321 0 net=2008
rlabel metal2 296 -321 296 -321 0 net=2139
rlabel metal2 450 -321 450 -321 0 net=2390
rlabel metal2 61 -323 61 -323 0 net=533
rlabel metal2 184 -323 184 -323 0 net=787
rlabel metal2 254 -323 254 -323 0 net=1198
rlabel metal2 373 -323 373 -323 0 net=1877
rlabel metal2 471 -323 471 -323 0 net=2739
rlabel metal2 65 -325 65 -325 0 net=1633
rlabel metal2 79 -325 79 -325 0 net=1781
rlabel metal2 226 -325 226 -325 0 net=1213
rlabel metal2 268 -325 268 -325 0 net=1992
rlabel metal2 348 -325 348 -325 0 net=2727
rlabel metal2 72 -327 72 -327 0 net=1071
rlabel metal2 184 -327 184 -327 0 net=725
rlabel metal2 219 -327 219 -327 0 net=1353
rlabel metal2 282 -327 282 -327 0 net=2999
rlabel metal2 86 -329 86 -329 0 net=1383
rlabel metal2 194 -329 194 -329 0 net=2214
rlabel metal2 219 -329 219 -329 0 net=1487
rlabel metal2 299 -329 299 -329 0 net=2707
rlabel metal2 103 -331 103 -331 0 net=1727
rlabel metal2 261 -331 261 -331 0 net=1811
rlabel metal2 310 -331 310 -331 0 net=2825
rlabel metal2 107 -333 107 -333 0 net=1132
rlabel metal2 142 -333 142 -333 0 net=1493
rlabel metal2 348 -333 348 -333 0 net=295
rlabel metal2 114 -335 114 -335 0 net=2114
rlabel metal2 534 -335 534 -335 0 net=2883
rlabel metal2 114 -337 114 -337 0 net=1611
rlabel metal2 149 -337 149 -337 0 net=737
rlabel metal2 194 -337 194 -337 0 net=2039
rlabel metal2 317 -337 317 -337 0 net=2593
rlabel metal2 121 -339 121 -339 0 net=265
rlabel metal2 198 -339 198 -339 0 net=1275
rlabel metal2 317 -339 317 -339 0 net=2081
rlabel metal2 345 -339 345 -339 0 net=2533
rlabel metal2 163 -341 163 -341 0 net=1293
rlabel metal2 352 -341 352 -341 0 net=1775
rlabel metal2 156 -343 156 -343 0 net=763
rlabel metal2 352 -343 352 -343 0 net=2511
rlabel metal2 156 -345 156 -345 0 net=1673
rlabel metal2 373 -345 373 -345 0 net=2059
rlabel metal2 380 -347 380 -347 0 net=2968
rlabel metal2 383 -349 383 -349 0 net=2048
rlabel metal2 387 -351 387 -351 0 net=2479
rlabel metal2 341 -353 341 -353 0 net=2891
rlabel metal2 394 -353 394 -353 0 net=2663
rlabel metal2 271 -355 271 -355 0 net=1357
rlabel metal2 401 -355 401 -355 0 net=2277
rlabel metal2 443 -355 443 -355 0 net=2303
rlabel metal2 292 -357 292 -357 0 net=1447
rlabel metal2 436 -357 436 -357 0 net=2647
rlabel metal2 205 -359 205 -359 0 net=2441
rlabel metal2 2 -370 2 -370 0 net=2323
rlabel metal2 201 -370 201 -370 0 net=1769
rlabel metal2 345 -370 345 -370 0 net=1878
rlabel metal2 485 -370 485 -370 0 net=2575
rlabel metal2 485 -370 485 -370 0 net=2575
rlabel metal2 513 -370 513 -370 0 net=2709
rlabel metal2 9 -372 9 -372 0 net=2482
rlabel metal2 156 -372 156 -372 0 net=764
rlabel metal2 184 -372 184 -372 0 net=727
rlabel metal2 348 -372 348 -372 0 net=1358
rlabel metal2 422 -372 422 -372 0 net=2513
rlabel metal2 534 -372 534 -372 0 net=2535
rlabel metal2 16 -374 16 -374 0 net=1810
rlabel metal2 254 -374 254 -374 0 net=1214
rlabel metal2 296 -374 296 -374 0 net=2304
rlabel metal2 555 -374 555 -374 0 net=3039
rlabel metal2 23 -376 23 -376 0 net=2720
rlabel metal2 156 -376 156 -376 0 net=85
rlabel metal2 313 -376 313 -376 0 net=2740
rlabel metal2 23 -378 23 -378 0 net=1387
rlabel metal2 37 -378 37 -378 0 net=274
rlabel metal2 65 -378 65 -378 0 net=1634
rlabel metal2 219 -378 219 -378 0 net=1488
rlabel metal2 352 -378 352 -378 0 net=2899
rlabel metal2 30 -380 30 -380 0 net=806
rlabel metal2 68 -380 68 -380 0 net=779
rlabel metal2 226 -380 226 -380 0 net=1355
rlabel metal2 296 -380 296 -380 0 net=2083
rlabel metal2 355 -380 355 -380 0 net=2802
rlabel metal2 37 -382 37 -382 0 net=2437
rlabel metal2 149 -382 149 -382 0 net=1431
rlabel metal2 170 -382 170 -382 0 net=739
rlabel metal2 299 -382 299 -382 0 net=1776
rlabel metal2 443 -382 443 -382 0 net=2649
rlabel metal2 44 -384 44 -384 0 net=1642
rlabel metal2 303 -384 303 -384 0 net=2041
rlabel metal2 366 -384 366 -384 0 net=2480
rlabel metal2 471 -384 471 -384 0 net=2729
rlabel metal2 44 -386 44 -386 0 net=1345
rlabel metal2 121 -386 121 -386 0 net=1813
rlabel metal2 268 -386 268 -386 0 net=2901
rlabel metal2 380 -386 380 -386 0 net=1201
rlabel metal2 51 -388 51 -388 0 net=1143
rlabel metal2 233 -388 233 -388 0 net=1729
rlabel metal2 320 -388 320 -388 0 net=2837
rlabel metal2 51 -390 51 -390 0 net=2121
rlabel metal2 107 -390 107 -390 0 net=1613
rlabel metal2 170 -390 170 -390 0 net=1295
rlabel metal2 233 -390 233 -390 0 net=863
rlabel metal2 380 -390 380 -390 0 net=2388
rlabel metal2 58 -392 58 -392 0 net=1463
rlabel metal2 212 -392 212 -392 0 net=1887
rlabel metal2 390 -392 390 -392 0 net=2125
rlabel metal2 72 -394 72 -394 0 net=1072
rlabel metal2 191 -394 191 -394 0 net=1189
rlabel metal2 394 -394 394 -394 0 net=2279
rlabel metal2 408 -394 408 -394 0 net=1448
rlabel metal2 443 -394 443 -394 0 net=2595
rlabel metal2 527 -394 527 -394 0 net=3001
rlabel metal2 72 -396 72 -396 0 net=1783
rlabel metal2 100 -396 100 -396 0 net=1897
rlabel metal2 373 -396 373 -396 0 net=2061
rlabel metal2 415 -396 415 -396 0 net=2665
rlabel metal2 558 -396 558 -396 0 net=1971
rlabel metal2 79 -398 79 -398 0 net=1782
rlabel metal2 348 -398 348 -398 0 net=1697
rlabel metal2 387 -398 387 -398 0 net=2893
rlabel metal2 79 -400 79 -400 0 net=1495
rlabel metal2 152 -400 152 -400 0 net=2140
rlabel metal2 450 -400 450 -400 0 net=2827
rlabel metal2 86 -402 86 -402 0 net=1384
rlabel metal2 383 -402 383 -402 0 net=2391
rlabel metal2 457 -402 457 -402 0 net=2505
rlabel metal2 93 -404 93 -404 0 net=1060
rlabel metal2 138 -404 138 -404 0 net=217
rlabel metal2 411 -404 411 -404 0 net=2753
rlabel metal2 9 -406 9 -406 0 net=196
rlabel metal2 142 -406 142 -406 0 net=1277
rlabel metal2 243 -406 243 -406 0 net=788
rlabel metal2 429 -406 429 -406 0 net=2885
rlabel metal2 114 -408 114 -408 0 net=1573
rlabel metal2 247 -408 247 -408 0 net=2713
rlabel metal2 541 -408 541 -408 0 net=2987
rlabel metal2 359 -410 359 -410 0 net=1675
rlabel metal2 436 -412 436 -412 0 net=2443
rlabel metal2 324 -414 324 -414 0 net=2621
rlabel metal2 2 -425 2 -425 0 net=2324
rlabel metal2 198 -425 198 -425 0 net=1144
rlabel metal2 240 -425 240 -425 0 net=2349
rlabel metal2 576 -425 576 -425 0 net=2127
rlabel metal2 611 -425 611 -425 0 net=2537
rlabel metal2 663 -425 663 -425 0 net=2641
rlabel metal2 2 -427 2 -427 0 net=2123
rlabel metal2 79 -427 79 -427 0 net=1496
rlabel metal2 208 -427 208 -427 0 net=2900
rlabel metal2 355 -427 355 -427 0 net=2280
rlabel metal2 464 -427 464 -427 0 net=2839
rlabel metal2 635 -427 635 -427 0 net=2627
rlabel metal2 9 -429 9 -429 0 net=1785
rlabel metal2 79 -429 79 -429 0 net=781
rlabel metal2 257 -429 257 -429 0 net=728
rlabel metal2 348 -429 348 -429 0 net=2730
rlabel metal2 506 -429 506 -429 0 net=2755
rlabel metal2 16 -431 16 -431 0 net=1575
rlabel metal2 128 -431 128 -431 0 net=50
rlabel metal2 170 -431 170 -431 0 net=1297
rlabel metal2 268 -431 268 -431 0 net=1625
rlabel metal2 268 -431 268 -431 0 net=1625
rlabel metal2 271 -431 271 -431 0 net=1356
rlabel metal2 310 -431 310 -431 0 net=2042
rlabel metal2 422 -431 422 -431 0 net=2515
rlabel metal2 513 -431 513 -431 0 net=2715
rlabel metal2 583 -431 583 -431 0 net=2711
rlabel metal2 19 -433 19 -433 0 net=2163
rlabel metal2 275 -433 275 -433 0 net=667
rlabel metal2 313 -433 313 -433 0 net=2666
rlabel metal2 436 -433 436 -433 0 net=2623
rlabel metal2 30 -435 30 -435 0 net=897
rlabel metal2 44 -435 44 -435 0 net=1346
rlabel metal2 226 -435 226 -435 0 net=1899
rlabel metal2 492 -435 492 -435 0 net=2895
rlabel metal2 527 -435 527 -435 0 net=3003
rlabel metal2 44 -437 44 -437 0 net=224
rlabel metal2 47 -439 47 -439 0 net=1888
rlabel metal2 233 -439 233 -439 0 net=865
rlabel metal2 317 -439 317 -439 0 net=1202
rlabel metal2 51 -441 51 -441 0 net=1115
rlabel metal2 362 -441 362 -441 0 net=3040
rlabel metal2 68 -443 68 -443 0 net=1499
rlabel metal2 373 -443 373 -443 0 net=1699
rlabel metal2 401 -443 401 -443 0 net=2063
rlabel metal2 457 -443 457 -443 0 net=2445
rlabel metal2 72 -445 72 -445 0 net=1731
rlabel metal2 275 -445 275 -445 0 net=1621
rlabel metal2 478 -445 478 -445 0 net=2507
rlabel metal2 86 -447 86 -447 0 net=535
rlabel metal2 177 -447 177 -447 0 net=1191
rlabel metal2 278 -447 278 -447 0 net=2084
rlabel metal2 303 -447 303 -447 0 net=2217
rlabel metal2 499 -447 499 -447 0 net=2651
rlabel metal2 86 -449 86 -449 0 net=1013
rlabel metal2 282 -449 282 -449 0 net=1833
rlabel metal2 380 -449 380 -449 0 net=2886
rlabel metal2 93 -451 93 -451 0 net=2197
rlabel metal2 93 -453 93 -453 0 net=1865
rlabel metal2 121 -453 121 -453 0 net=1815
rlabel metal2 243 -453 243 -453 0 net=1671
rlabel metal2 429 -453 429 -453 0 net=1677
rlabel metal2 96 -455 96 -455 0 net=695
rlabel metal2 138 -455 138 -455 0 net=567
rlabel metal2 296 -455 296 -455 0 net=2325
rlabel metal2 534 -455 534 -455 0 net=2829
rlabel metal2 100 -457 100 -457 0 net=741
rlabel metal2 191 -457 191 -457 0 net=2667
rlabel metal2 145 -459 145 -459 0 net=919
rlabel metal2 254 -459 254 -459 0 net=2369
rlabel metal2 149 -461 149 -461 0 net=1433
rlabel metal2 170 -461 170 -461 0 net=1753
rlabel metal2 58 -463 58 -463 0 net=1465
rlabel metal2 254 -463 254 -463 0 net=1173
rlabel metal2 310 -463 310 -463 0 net=2347
rlabel metal2 58 -465 58 -465 0 net=1061
rlabel metal2 156 -465 156 -465 0 net=1119
rlabel metal2 317 -465 317 -465 0 net=1331
rlabel metal2 37 -467 37 -467 0 net=2438
rlabel metal2 320 -467 320 -467 0 net=2902
rlabel metal2 23 -469 23 -469 0 net=1388
rlabel metal2 201 -469 201 -469 0 net=1647
rlabel metal2 23 -471 23 -471 0 net=1279
rlabel metal2 324 -471 324 -471 0 net=2263
rlabel metal2 135 -473 135 -473 0 net=263
rlabel metal2 324 -473 324 -473 0 net=2453
rlabel metal2 107 -475 107 -475 0 net=1614
rlabel metal2 327 -475 327 -475 0 net=2596
rlabel metal2 107 -477 107 -477 0 net=1323
rlabel metal2 327 -477 327 -477 0 net=2887
rlabel metal2 124 -479 124 -479 0 net=2161
rlabel metal2 331 -481 331 -481 0 net=1771
rlabel metal2 331 -483 331 -483 0 net=2988
rlabel metal2 334 -485 334 -485 0 net=1181
rlabel metal2 450 -485 450 -485 0 net=2393
rlabel metal2 450 -487 450 -487 0 net=1973
rlabel metal2 485 -489 485 -489 0 net=2577
rlabel metal2 422 -491 422 -491 0 net=2103
rlabel metal2 2 -502 2 -502 0 net=2124
rlabel metal2 51 -502 51 -502 0 net=1116
rlabel metal2 128 -502 128 -502 0 net=1816
rlabel metal2 236 -502 236 -502 0 net=2218
rlabel metal2 492 -502 492 -502 0 net=2830
rlabel metal2 597 -502 597 -502 0 net=2128
rlabel metal2 635 -502 635 -502 0 net=2642
rlabel metal2 9 -504 9 -504 0 net=1786
rlabel metal2 205 -504 205 -504 0 net=1900
rlabel metal2 422 -504 422 -504 0 net=2199
rlabel metal2 492 -504 492 -504 0 net=2579
rlabel metal2 597 -504 597 -504 0 net=2889
rlabel metal2 16 -506 16 -506 0 net=1576
rlabel metal2 208 -506 208 -506 0 net=1298
rlabel metal2 240 -506 240 -506 0 net=2162
rlabel metal2 464 -506 464 -506 0 net=2447
rlabel metal2 604 -506 604 -506 0 net=2712
rlabel metal2 618 -506 618 -506 0 net=2628
rlabel metal2 16 -508 16 -508 0 net=2257
rlabel metal2 79 -508 79 -508 0 net=782
rlabel metal2 289 -508 289 -508 0 net=866
rlabel metal2 310 -508 310 -508 0 net=2085
rlabel metal2 513 -508 513 -508 0 net=2897
rlabel metal2 639 -508 639 -508 0 net=2539
rlabel metal2 23 -510 23 -510 0 net=1280
rlabel metal2 212 -510 212 -510 0 net=1841
rlabel metal2 345 -510 345 -510 0 net=2669
rlabel metal2 576 -510 576 -510 0 net=2716
rlabel metal2 23 -512 23 -512 0 net=899
rlabel metal2 37 -512 37 -512 0 net=1449
rlabel metal2 397 -512 397 -512 0 net=2652
rlabel metal2 541 -512 541 -512 0 net=2395
rlabel metal2 541 -512 541 -512 0 net=2395
rlabel metal2 30 -514 30 -514 0 net=1733
rlabel metal2 86 -514 86 -514 0 net=1014
rlabel metal2 170 -514 170 -514 0 net=2516
rlabel metal2 513 -514 513 -514 0 net=2509
rlabel metal2 51 -516 51 -516 0 net=2027
rlabel metal2 334 -516 334 -516 0 net=2929
rlabel metal2 58 -518 58 -518 0 net=1062
rlabel metal2 303 -518 303 -518 0 net=2454
rlabel metal2 527 -518 527 -518 0 net=2745
rlabel metal2 86 -520 86 -520 0 net=1835
rlabel metal2 310 -520 310 -520 0 net=1649
rlabel metal2 369 -520 369 -520 0 net=2629
rlabel metal2 555 -520 555 -520 0 net=2757
rlabel metal2 621 -520 621 -520 0 net=2517
rlabel metal2 93 -522 93 -522 0 net=1867
rlabel metal2 131 -522 131 -522 0 net=2683
rlabel metal2 590 -522 590 -522 0 net=2841
rlabel metal2 93 -524 93 -524 0 net=2603
rlabel metal2 282 -524 282 -524 0 net=1263
rlabel metal2 355 -524 355 -524 0 net=2348
rlabel metal2 495 -524 495 -524 0 net=2561
rlabel metal2 625 -524 625 -524 0 net=432
rlabel metal2 100 -526 100 -526 0 net=743
rlabel metal2 191 -526 191 -526 0 net=920
rlabel metal2 275 -526 275 -526 0 net=1623
rlabel metal2 324 -526 324 -526 0 net=1678
rlabel metal2 478 -526 478 -526 0 net=2371
rlabel metal2 100 -528 100 -528 0 net=1467
rlabel metal2 170 -528 170 -528 0 net=1471
rlabel metal2 226 -528 226 -528 0 net=1627
rlabel metal2 275 -528 275 -528 0 net=2264
rlabel metal2 485 -528 485 -528 0 net=2105
rlabel metal2 107 -530 107 -530 0 net=1325
rlabel metal2 324 -530 324 -530 0 net=831
rlabel metal2 397 -530 397 -530 0 net=3004
rlabel metal2 107 -532 107 -532 0 net=1435
rlabel metal2 163 -532 163 -532 0 net=1109
rlabel metal2 65 -534 65 -534 0 net=1245
rlabel metal2 177 -534 177 -534 0 net=1193
rlabel metal2 348 -534 348 -534 0 net=2763
rlabel metal2 457 -534 457 -534 0 net=2691
rlabel metal2 61 -536 61 -536 0 net=1587
rlabel metal2 198 -536 198 -536 0 net=1175
rlabel metal2 362 -536 362 -536 0 net=1974
rlabel metal2 121 -538 121 -538 0 net=1489
rlabel metal2 135 -538 135 -538 0 net=1121
rlabel metal2 205 -538 205 -538 0 net=2365
rlabel metal2 142 -540 142 -540 0 net=1035
rlabel metal2 254 -540 254 -540 0 net=1165
rlabel metal2 366 -540 366 -540 0 net=1772
rlabel metal2 429 -540 429 -540 0 net=2351
rlabel metal2 145 -542 145 -542 0 net=355
rlabel metal2 156 -544 156 -544 0 net=2409
rlabel metal2 373 -544 373 -544 0 net=1672
rlabel metal2 436 -544 436 -544 0 net=2065
rlabel metal2 520 -544 520 -544 0 net=2625
rlabel metal2 632 -544 632 -544 0 net=2635
rlabel metal2 271 -546 271 -546 0 net=3029
rlabel metal2 338 -548 338 -548 0 net=1501
rlabel metal2 296 -550 296 -550 0 net=2327
rlabel metal2 373 -550 373 -550 0 net=1755
rlabel metal2 296 -552 296 -552 0 net=1333
rlabel metal2 380 -552 380 -552 0 net=1182
rlabel metal2 247 -554 247 -554 0 net=2165
rlabel metal2 380 -554 380 -554 0 net=3025
rlabel metal2 247 -556 247 -556 0 net=1981
rlabel metal2 383 -556 383 -556 0 net=1700
rlabel metal2 2 -567 2 -567 0 net=2605
rlabel metal2 100 -567 100 -567 0 net=1468
rlabel metal2 156 -567 156 -567 0 net=1194
rlabel metal2 254 -567 254 -567 0 net=1166
rlabel metal2 369 -567 369 -567 0 net=2448
rlabel metal2 485 -567 485 -567 0 net=2758
rlabel metal2 576 -567 576 -567 0 net=3027
rlabel metal2 618 -567 618 -567 0 net=679
rlabel metal2 632 -567 632 -567 0 net=2637
rlabel metal2 632 -567 632 -567 0 net=2637
rlabel metal2 642 -567 642 -567 0 net=2518
rlabel metal2 9 -569 9 -569 0 net=2175
rlabel metal2 114 -569 114 -569 0 net=1868
rlabel metal2 170 -569 170 -569 0 net=1842
rlabel metal2 233 -569 233 -569 0 net=1036
rlabel metal2 271 -569 271 -569 0 net=2166
rlabel metal2 352 -569 352 -569 0 net=2842
rlabel metal2 646 -569 646 -569 0 net=2541
rlabel metal2 16 -571 16 -571 0 net=2258
rlabel metal2 114 -571 114 -571 0 net=1123
rlabel metal2 142 -571 142 -571 0 net=1931
rlabel metal2 208 -571 208 -571 0 net=512
rlabel metal2 261 -571 261 -571 0 net=449
rlabel metal2 408 -571 408 -571 0 net=2898
rlabel metal2 16 -573 16 -573 0 net=1651
rlabel metal2 331 -573 331 -573 0 net=2945
rlabel metal2 23 -575 23 -575 0 net=900
rlabel metal2 82 -575 82 -575 0 net=1787
rlabel metal2 135 -575 135 -575 0 net=901
rlabel metal2 268 -575 268 -575 0 net=833
rlabel metal2 373 -575 373 -575 0 net=1757
rlabel metal2 583 -575 583 -575 0 net=3031
rlabel metal2 23 -577 23 -577 0 net=1019
rlabel metal2 194 -577 194 -577 0 net=1628
rlabel metal2 278 -577 278 -577 0 net=1315
rlabel metal2 324 -577 324 -577 0 net=2066
rlabel metal2 464 -577 464 -577 0 net=2367
rlabel metal2 544 -577 544 -577 0 net=2890
rlabel metal2 30 -579 30 -579 0 net=1735
rlabel metal2 383 -579 383 -579 0 net=378
rlabel metal2 429 -579 429 -579 0 net=2353
rlabel metal2 450 -579 450 -579 0 net=1953
rlabel metal2 30 -581 30 -581 0 net=1593
rlabel metal2 79 -581 79 -581 0 net=1111
rlabel metal2 170 -581 170 -581 0 net=745
rlabel metal2 198 -581 198 -581 0 net=1176
rlabel metal2 205 -581 205 -581 0 net=2189
rlabel metal2 429 -581 429 -581 0 net=2373
rlabel metal2 506 -581 506 -581 0 net=2563
rlabel metal2 51 -583 51 -583 0 net=2029
rlabel metal2 289 -583 289 -583 0 net=1327
rlabel metal2 289 -583 289 -583 0 net=1327
rlabel metal2 303 -583 303 -583 0 net=1624
rlabel metal2 387 -583 387 -583 0 net=2626
rlabel metal2 565 -583 565 -583 0 net=2991
rlabel metal2 51 -585 51 -585 0 net=1491
rlabel metal2 152 -585 152 -585 0 net=507
rlabel metal2 177 -585 177 -585 0 net=1589
rlabel metal2 296 -585 296 -585 0 net=1335
rlabel metal2 310 -585 310 -585 0 net=1502
rlabel metal2 443 -585 443 -585 0 net=2764
rlabel metal2 506 -585 506 -585 0 net=2671
rlabel metal2 569 -585 569 -585 0 net=2931
rlabel metal2 61 -587 61 -587 0 net=1205
rlabel metal2 264 -587 264 -587 0 net=2697
rlabel metal2 471 -587 471 -587 0 net=2631
rlabel metal2 520 -587 520 -587 0 net=2107
rlabel metal2 548 -587 548 -587 0 net=2685
rlabel metal2 65 -589 65 -589 0 net=1247
rlabel metal2 345 -589 345 -589 0 net=2609
rlabel metal2 527 -589 527 -589 0 net=2747
rlabel metal2 68 -591 68 -591 0 net=143
rlabel metal2 152 -591 152 -591 0 net=2328
rlabel metal2 394 -591 394 -591 0 net=2565
rlabel metal2 534 -591 534 -591 0 net=2397
rlabel metal2 72 -593 72 -593 0 net=1473
rlabel metal2 226 -593 226 -593 0 net=1264
rlabel metal2 338 -593 338 -593 0 net=1935
rlabel metal2 401 -593 401 -593 0 net=2510
rlabel metal2 58 -595 58 -595 0 net=789
rlabel metal2 247 -595 247 -595 0 net=1983
rlabel metal2 401 -595 401 -595 0 net=2580
rlabel metal2 86 -597 86 -597 0 net=1836
rlabel metal2 457 -597 457 -597 0 net=2693
rlabel metal2 86 -599 86 -599 0 net=2129
rlabel metal2 198 -599 198 -599 0 net=2723
rlabel metal2 107 -601 107 -601 0 net=1436
rlabel metal2 212 -601 212 -601 0 net=1849
rlabel metal2 492 -601 492 -601 0 net=2219
rlabel metal2 37 -603 37 -603 0 net=1451
rlabel metal2 121 -603 121 -603 0 net=1705
rlabel metal2 37 -605 37 -605 0 net=1551
rlabel metal2 156 -605 156 -605 0 net=909
rlabel metal2 180 -605 180 -605 0 net=1259
rlabel metal2 282 -605 282 -605 0 net=2087
rlabel metal2 44 -607 44 -607 0 net=1037
rlabel metal2 348 -607 348 -607 0 net=1151
rlabel metal2 415 -607 415 -607 0 net=2201
rlabel metal2 359 -609 359 -609 0 net=2411
rlabel metal2 359 -611 359 -611 0 net=2145
rlabel metal2 2 -622 2 -622 0 net=2606
rlabel metal2 131 -622 131 -622 0 net=76
rlabel metal2 212 -622 212 -622 0 net=1850
rlabel metal2 345 -622 345 -622 0 net=2748
rlabel metal2 625 -622 625 -622 0 net=220
rlabel metal2 653 -622 653 -622 0 net=2543
rlabel metal2 653 -622 653 -622 0 net=2543
rlabel metal2 2 -624 2 -624 0 net=1789
rlabel metal2 100 -624 100 -624 0 net=771
rlabel metal2 156 -624 156 -624 0 net=911
rlabel metal2 156 -624 156 -624 0 net=911
rlabel metal2 173 -624 173 -624 0 net=2932
rlabel metal2 632 -624 632 -624 0 net=2639
rlabel metal2 632 -624 632 -624 0 net=2639
rlabel metal2 9 -626 9 -626 0 net=2176
rlabel metal2 208 -626 208 -626 0 net=2992
rlabel metal2 9 -628 9 -628 0 net=893
rlabel metal2 103 -628 103 -628 0 net=327
rlabel metal2 201 -628 201 -628 0 net=1590
rlabel metal2 296 -628 296 -628 0 net=1248
rlabel metal2 334 -628 334 -628 0 net=517
rlabel metal2 565 -628 565 -628 0 net=2946
rlabel metal2 16 -630 16 -630 0 net=1652
rlabel metal2 289 -630 289 -630 0 net=1329
rlabel metal2 313 -630 313 -630 0 net=2374
rlabel metal2 443 -630 443 -630 0 net=2355
rlabel metal2 499 -630 499 -630 0 net=2611
rlabel metal2 499 -630 499 -630 0 net=2611
rlabel metal2 513 -630 513 -630 0 net=2695
rlabel metal2 16 -632 16 -632 0 net=917
rlabel metal2 184 -632 184 -632 0 net=2115
rlabel metal2 362 -632 362 -632 0 net=2564
rlabel metal2 23 -634 23 -634 0 net=1020
rlabel metal2 219 -634 219 -634 0 net=790
rlabel metal2 348 -634 348 -634 0 net=1758
rlabel metal2 23 -636 23 -636 0 net=593
rlabel metal2 107 -636 107 -636 0 net=1453
rlabel metal2 114 -636 114 -636 0 net=1124
rlabel metal2 170 -636 170 -636 0 net=746
rlabel metal2 219 -636 219 -636 0 net=433
rlabel metal2 415 -636 415 -636 0 net=2203
rlabel metal2 415 -636 415 -636 0 net=2203
rlabel metal2 443 -636 443 -636 0 net=2221
rlabel metal2 520 -636 520 -636 0 net=2108
rlabel metal2 30 -638 30 -638 0 net=1594
rlabel metal2 177 -638 177 -638 0 net=1736
rlabel metal2 429 -638 429 -638 0 net=2525
rlabel metal2 520 -638 520 -638 0 net=2687
rlabel metal2 30 -640 30 -640 0 net=1077
rlabel metal2 324 -640 324 -640 0 net=2981
rlabel metal2 37 -642 37 -642 0 net=1552
rlabel metal2 107 -642 107 -642 0 net=1073
rlabel metal2 222 -642 222 -642 0 net=1316
rlabel metal2 324 -642 324 -642 0 net=2109
rlabel metal2 460 -642 460 -642 0 net=3028
rlabel metal2 37 -644 37 -644 0 net=1933
rlabel metal2 226 -644 226 -644 0 net=2146
rlabel metal2 527 -644 527 -644 0 net=3032
rlabel metal2 44 -646 44 -646 0 net=1038
rlabel metal2 226 -646 226 -646 0 net=1261
rlabel metal2 257 -646 257 -646 0 net=2368
rlabel metal2 44 -648 44 -648 0 net=813
rlabel metal2 240 -648 240 -648 0 net=1206
rlabel metal2 303 -648 303 -648 0 net=1337
rlabel metal2 338 -648 338 -648 0 net=1937
rlabel metal2 387 -648 387 -648 0 net=1985
rlabel metal2 436 -648 436 -648 0 net=2699
rlabel metal2 51 -650 51 -650 0 net=1492
rlabel metal2 247 -650 247 -650 0 net=1281
rlabel metal2 51 -652 51 -652 0 net=1283
rlabel metal2 275 -652 275 -652 0 net=2205
rlabel metal2 345 -652 345 -652 0 net=1397
rlabel metal2 408 -652 408 -652 0 net=2191
rlabel metal2 58 -654 58 -654 0 net=1265
rlabel metal2 282 -654 282 -654 0 net=2089
rlabel metal2 310 -654 310 -654 0 net=2283
rlabel metal2 61 -656 61 -656 0 net=2724
rlabel metal2 65 -658 65 -658 0 net=973
rlabel metal2 268 -658 268 -658 0 net=834
rlabel metal2 313 -658 313 -658 0 net=2765
rlabel metal2 513 -658 513 -658 0 net=2313
rlabel metal2 72 -660 72 -660 0 net=1475
rlabel metal2 352 -660 352 -660 0 net=1707
rlabel metal2 408 -660 408 -660 0 net=1955
rlabel metal2 72 -662 72 -662 0 net=1717
rlabel metal2 135 -662 135 -662 0 net=903
rlabel metal2 180 -662 180 -662 0 net=2229
rlabel metal2 79 -664 79 -664 0 net=1113
rlabel metal2 355 -664 355 -664 0 net=2412
rlabel metal2 79 -666 79 -666 0 net=937
rlabel metal2 191 -666 191 -666 0 net=815
rlabel metal2 422 -666 422 -666 0 net=2398
rlabel metal2 366 -668 366 -668 0 net=1152
rlabel metal2 506 -668 506 -668 0 net=2673
rlabel metal2 121 -670 121 -670 0 net=2030
rlabel metal2 369 -670 369 -670 0 net=2632
rlabel metal2 485 -670 485 -670 0 net=2567
rlabel metal2 86 -672 86 -672 0 net=2131
rlabel metal2 257 -672 257 -672 0 net=2431
rlabel metal2 86 -674 86 -674 0 net=1053
rlabel metal2 394 -674 394 -674 0 net=2461
rlabel metal2 121 -676 121 -676 0 net=1153
rlabel metal2 2 -687 2 -687 0 net=1790
rlabel metal2 219 -687 219 -687 0 net=160
rlabel metal2 289 -687 289 -687 0 net=1559
rlabel metal2 313 -687 313 -687 0 net=2204
rlabel metal2 422 -687 422 -687 0 net=2067
rlabel metal2 429 -687 429 -687 0 net=2231
rlabel metal2 457 -687 457 -687 0 net=2767
rlabel metal2 632 -687 632 -687 0 net=2640
rlabel metal2 653 -687 653 -687 0 net=2544
rlabel metal2 653 -687 653 -687 0 net=2544
rlabel metal2 2 -689 2 -689 0 net=1267
rlabel metal2 65 -689 65 -689 0 net=975
rlabel metal2 65 -689 65 -689 0 net=975
rlabel metal2 96 -689 96 -689 0 net=46
rlabel metal2 177 -689 177 -689 0 net=532
rlabel metal2 278 -689 278 -689 0 net=1330
rlabel metal2 317 -689 317 -689 0 net=1339
rlabel metal2 317 -689 317 -689 0 net=1339
rlabel metal2 331 -689 331 -689 0 net=2849
rlabel metal2 478 -689 478 -689 0 net=2357
rlabel metal2 9 -691 9 -691 0 net=894
rlabel metal2 135 -691 135 -691 0 net=913
rlabel metal2 170 -691 170 -691 0 net=817
rlabel metal2 194 -691 194 -691 0 net=1262
rlabel metal2 229 -691 229 -691 0 net=2759
rlabel metal2 12 -693 12 -693 0 net=1521
rlabel metal2 397 -693 397 -693 0 net=2982
rlabel metal2 562 -693 562 -693 0 net=70
rlabel metal2 16 -695 16 -695 0 net=918
rlabel metal2 121 -695 121 -695 0 net=1341
rlabel metal2 187 -695 187 -695 0 net=2449
rlabel metal2 16 -697 16 -697 0 net=1513
rlabel metal2 114 -697 114 -697 0 net=2337
rlabel metal2 30 -699 30 -699 0 net=1078
rlabel metal2 156 -699 156 -699 0 net=1155
rlabel metal2 219 -699 219 -699 0 net=1285
rlabel metal2 271 -699 271 -699 0 net=1373
rlabel metal2 338 -699 338 -699 0 net=2207
rlabel metal2 30 -701 30 -701 0 net=1075
rlabel metal2 114 -701 114 -701 0 net=2003
rlabel metal2 485 -701 485 -701 0 net=2463
rlabel metal2 37 -703 37 -703 0 net=1934
rlabel metal2 278 -703 278 -703 0 net=1879
rlabel metal2 404 -703 404 -703 0 net=2287
rlabel metal2 37 -705 37 -705 0 net=1055
rlabel metal2 117 -705 117 -705 0 net=1425
rlabel metal2 341 -705 341 -705 0 net=2222
rlabel metal2 464 -705 464 -705 0 net=2285
rlabel metal2 44 -707 44 -707 0 net=814
rlabel metal2 51 -707 51 -707 0 net=1407
rlabel metal2 345 -707 345 -707 0 net=1399
rlabel metal2 432 -707 432 -707 0 net=2568
rlabel metal2 520 -707 520 -707 0 net=2689
rlabel metal2 54 -709 54 -709 0 net=1114
rlabel metal2 247 -709 247 -709 0 net=1282
rlabel metal2 292 -709 292 -709 0 net=2159
rlabel metal2 527 -709 527 -709 0 net=2701
rlabel metal2 82 -711 82 -711 0 net=2241
rlabel metal2 226 -711 226 -711 0 net=2432
rlabel metal2 492 -711 492 -711 0 net=2527
rlabel metal2 86 -713 86 -713 0 net=905
rlabel metal2 145 -713 145 -713 0 net=2247
rlabel metal2 100 -715 100 -715 0 net=773
rlabel metal2 254 -715 254 -715 0 net=983
rlabel metal2 376 -715 376 -715 0 net=2696
rlabel metal2 128 -717 128 -717 0 net=1007
rlabel metal2 198 -717 198 -717 0 net=2110
rlabel metal2 345 -717 345 -717 0 net=1413
rlabel metal2 376 -717 376 -717 0 net=2989
rlabel metal2 107 -719 107 -719 0 net=1967
rlabel metal2 233 -719 233 -719 0 net=2132
rlabel metal2 380 -719 380 -719 0 net=1939
rlabel metal2 149 -721 149 -721 0 net=599
rlabel metal2 355 -721 355 -721 0 net=1523
rlabel metal2 499 -721 499 -721 0 net=2613
rlabel metal2 72 -723 72 -723 0 net=1719
rlabel metal2 72 -725 72 -725 0 net=939
rlabel metal2 149 -725 149 -725 0 net=81
rlabel metal2 359 -725 359 -725 0 net=2117
rlabel metal2 163 -727 163 -727 0 net=1455
rlabel metal2 268 -727 268 -727 0 net=1477
rlabel metal2 359 -727 359 -727 0 net=2674
rlabel metal2 166 -729 166 -729 0 net=1713
rlabel metal2 513 -729 513 -729 0 net=2315
rlabel metal2 177 -731 177 -731 0 net=851
rlabel metal2 268 -731 268 -731 0 net=2811
rlabel metal2 191 -733 191 -733 0 net=885
rlabel metal2 275 -733 275 -733 0 net=2329
rlabel metal2 187 -735 187 -735 0 net=669
rlabel metal2 303 -735 303 -735 0 net=2091
rlabel metal2 310 -737 310 -737 0 net=1709
rlabel metal2 366 -737 366 -737 0 net=1419
rlabel metal2 352 -739 352 -739 0 net=1986
rlabel metal2 408 -739 408 -739 0 net=1957
rlabel metal2 282 -741 282 -741 0 net=1891
rlabel metal2 436 -741 436 -741 0 net=2193
rlabel metal2 362 -743 362 -743 0 net=1869
rlabel metal2 2 -754 2 -754 0 net=1268
rlabel metal2 184 -754 184 -754 0 net=985
rlabel metal2 261 -754 261 -754 0 net=77
rlabel metal2 373 -754 373 -754 0 net=1870
rlabel metal2 471 -754 471 -754 0 net=2702
rlabel metal2 23 -756 23 -756 0 net=1892
rlabel metal2 471 -756 471 -756 0 net=2331
rlabel metal2 558 -756 558 -756 0 net=2990
rlabel metal2 23 -758 23 -758 0 net=2399
rlabel metal2 114 -758 114 -758 0 net=1456
rlabel metal2 243 -758 243 -758 0 net=1426
rlabel metal2 299 -758 299 -758 0 net=2208
rlabel metal2 30 -760 30 -760 0 net=1076
rlabel metal2 114 -760 114 -760 0 net=915
rlabel metal2 142 -760 142 -760 0 net=2528
rlabel metal2 30 -762 30 -762 0 net=1969
rlabel metal2 117 -762 117 -762 0 net=2141
rlabel metal2 261 -762 261 -762 0 net=1415
rlabel metal2 376 -762 376 -762 0 net=2358
rlabel metal2 597 -762 597 -762 0 net=1079
rlabel metal2 37 -764 37 -764 0 net=1056
rlabel metal2 152 -764 152 -764 0 net=753
rlabel metal2 187 -764 187 -764 0 net=1522
rlabel metal2 474 -764 474 -764 0 net=2288
rlabel metal2 583 -764 583 -764 0 net=2769
rlabel metal2 54 -766 54 -766 0 net=373
rlabel metal2 376 -766 376 -766 0 net=2690
rlabel metal2 61 -768 61 -768 0 net=2812
rlabel metal2 65 -770 65 -770 0 net=976
rlabel metal2 247 -770 247 -770 0 net=775
rlabel metal2 247 -770 247 -770 0 net=775
rlabel metal2 268 -770 268 -770 0 net=1340
rlabel metal2 327 -770 327 -770 0 net=1400
rlabel metal2 443 -770 443 -770 0 net=1714
rlabel metal2 618 -770 618 -770 0 net=2079
rlabel metal2 65 -772 65 -772 0 net=1157
rlabel metal2 191 -772 191 -772 0 net=1361
rlabel metal2 345 -772 345 -772 0 net=1445
rlabel metal2 380 -772 380 -772 0 net=2194
rlabel metal2 541 -772 541 -772 0 net=2761
rlabel metal2 79 -774 79 -774 0 net=2286
rlabel metal2 82 -776 82 -776 0 net=2092
rlabel metal2 44 -778 44 -778 0 net=2209
rlabel metal2 86 -778 86 -778 0 net=906
rlabel metal2 208 -778 208 -778 0 net=2338
rlabel metal2 96 -780 96 -780 0 net=951
rlabel metal2 107 -780 107 -780 0 net=1343
rlabel metal2 145 -780 145 -780 0 net=818
rlabel metal2 198 -780 198 -780 0 net=2004
rlabel metal2 93 -782 93 -782 0 net=1515
rlabel metal2 149 -782 149 -782 0 net=1003
rlabel metal2 219 -782 219 -782 0 net=1287
rlabel metal2 268 -782 268 -782 0 net=1711
rlabel metal2 331 -782 331 -782 0 net=1374
rlabel metal2 156 -784 156 -784 0 net=853
rlabel metal2 219 -784 219 -784 0 net=1427
rlabel metal2 58 -786 58 -786 0 net=1249
rlabel metal2 275 -786 275 -786 0 net=1478
rlabel metal2 359 -786 359 -786 0 net=1421
rlabel metal2 373 -786 373 -786 0 net=1553
rlabel metal2 58 -788 58 -788 0 net=941
rlabel metal2 170 -788 170 -788 0 net=1921
rlabel metal2 285 -788 285 -788 0 net=1720
rlabel metal2 72 -790 72 -790 0 net=1009
rlabel metal2 275 -790 275 -790 0 net=1940
rlabel metal2 278 -792 278 -792 0 net=1958
rlabel metal2 499 -792 499 -792 0 net=2615
rlabel metal2 198 -794 198 -794 0 net=1391
rlabel metal2 289 -794 289 -794 0 net=1560
rlabel metal2 411 -794 411 -794 0 net=2957
rlabel metal2 212 -796 212 -796 0 net=2243
rlabel metal2 415 -796 415 -796 0 net=2249
rlabel metal2 152 -798 152 -798 0 net=1145
rlabel metal2 233 -798 233 -798 0 net=887
rlabel metal2 303 -798 303 -798 0 net=1203
rlabel metal2 380 -798 380 -798 0 net=2233
rlabel metal2 443 -798 443 -798 0 net=2317
rlabel metal2 51 -800 51 -800 0 net=1409
rlabel metal2 310 -800 310 -800 0 net=2160
rlabel metal2 527 -800 527 -800 0 net=2451
rlabel metal2 320 -802 320 -802 0 net=1747
rlabel metal2 387 -802 387 -802 0 net=2439
rlabel metal2 562 -802 562 -802 0 net=2465
rlabel metal2 341 -804 341 -804 0 net=2771
rlabel metal2 341 -806 341 -806 0 net=2169
rlabel metal2 450 -806 450 -806 0 net=1525
rlabel metal2 390 -808 390 -808 0 net=1919
rlabel metal2 394 -810 394 -810 0 net=1881
rlabel metal2 422 -810 422 -810 0 net=2069
rlabel metal2 450 -810 450 -810 0 net=2119
rlabel metal2 313 -812 313 -812 0 net=2491
rlabel metal2 457 -812 457 -812 0 net=2851
rlabel metal2 457 -814 457 -814 0 net=2261
rlabel metal2 464 -816 464 -816 0 net=2427
rlabel metal2 9 -827 9 -827 0 net=2581
rlabel metal2 40 -827 40 -827 0 net=643
rlabel metal2 107 -827 107 -827 0 net=1344
rlabel metal2 149 -827 149 -827 0 net=1081
rlabel metal2 233 -827 233 -827 0 net=1410
rlabel metal2 387 -827 387 -827 0 net=2245
rlabel metal2 415 -827 415 -827 0 net=2251
rlabel metal2 415 -827 415 -827 0 net=2251
rlabel metal2 425 -827 425 -827 0 net=1920
rlabel metal2 513 -827 513 -827 0 net=2466
rlabel metal2 572 -827 572 -827 0 net=2080
rlabel metal2 16 -829 16 -829 0 net=2321
rlabel metal2 54 -829 54 -829 0 net=2332
rlabel metal2 478 -829 478 -829 0 net=2762
rlabel metal2 555 -829 555 -829 0 net=1555
rlabel metal2 30 -831 30 -831 0 net=1970
rlabel metal2 107 -831 107 -831 0 net=987
rlabel metal2 194 -831 194 -831 0 net=1146
rlabel metal2 222 -831 222 -831 0 net=259
rlabel metal2 292 -831 292 -831 0 net=2585
rlabel metal2 534 -831 534 -831 0 net=2770
rlabel metal2 58 -833 58 -833 0 net=942
rlabel metal2 89 -833 89 -833 0 net=952
rlabel metal2 114 -833 114 -833 0 net=916
rlabel metal2 170 -833 170 -833 0 net=1923
rlabel metal2 334 -833 334 -833 0 net=2958
rlabel metal2 562 -833 562 -833 0 net=1527
rlabel metal2 23 -835 23 -835 0 net=2400
rlabel metal2 180 -835 180 -835 0 net=995
rlabel metal2 247 -835 247 -835 0 net=776
rlabel metal2 268 -835 268 -835 0 net=1712
rlabel metal2 320 -835 320 -835 0 net=2170
rlabel metal2 464 -835 464 -835 0 net=2429
rlabel metal2 464 -835 464 -835 0 net=2429
rlabel metal2 478 -835 478 -835 0 net=2773
rlabel metal2 548 -835 548 -835 0 net=1080
rlabel metal2 23 -837 23 -837 0 net=2211
rlabel metal2 51 -837 51 -837 0 net=1403
rlabel metal2 114 -837 114 -837 0 net=1393
rlabel metal2 226 -837 226 -837 0 net=1288
rlabel metal2 303 -837 303 -837 0 net=1204
rlabel metal2 394 -837 394 -837 0 net=1883
rlabel metal2 394 -837 394 -837 0 net=1883
rlabel metal2 401 -837 401 -837 0 net=2120
rlabel metal2 485 -837 485 -837 0 net=2853
rlabel metal2 485 -837 485 -837 0 net=2853
rlabel metal2 499 -837 499 -837 0 net=2617
rlabel metal2 51 -839 51 -839 0 net=791
rlabel metal2 65 -839 65 -839 0 net=1158
rlabel metal2 247 -839 247 -839 0 net=889
rlabel metal2 317 -839 317 -839 0 net=2979
rlabel metal2 65 -841 65 -841 0 net=755
rlabel metal2 173 -841 173 -841 0 net=2903
rlabel metal2 320 -841 320 -841 0 net=2483
rlabel metal2 422 -841 422 -841 0 net=2493
rlabel metal2 72 -843 72 -843 0 net=1010
rlabel metal2 135 -843 135 -843 0 net=69
rlabel metal2 338 -843 338 -843 0 net=2234
rlabel metal2 404 -843 404 -843 0 net=2440
rlabel metal2 72 -845 72 -845 0 net=1669
rlabel metal2 86 -845 86 -845 0 net=1429
rlabel metal2 254 -845 254 -845 0 net=2143
rlabel metal2 345 -845 345 -845 0 net=1446
rlabel metal2 93 -847 93 -847 0 net=1313
rlabel metal2 163 -847 163 -847 0 net=1307
rlabel metal2 348 -847 348 -847 0 net=2262
rlabel metal2 121 -849 121 -849 0 net=1516
rlabel metal2 177 -849 177 -849 0 net=1251
rlabel metal2 352 -849 352 -849 0 net=1423
rlabel metal2 366 -849 366 -849 0 net=1749
rlabel metal2 366 -849 366 -849 0 net=1749
rlabel metal2 376 -849 376 -849 0 net=2267
rlabel metal2 429 -849 429 -849 0 net=2071
rlabel metal2 429 -849 429 -849 0 net=2071
rlabel metal2 436 -849 436 -849 0 net=2319
rlabel metal2 121 -851 121 -851 0 net=855
rlabel metal2 184 -851 184 -851 0 net=1363
rlabel metal2 198 -851 198 -851 0 net=2151
rlabel metal2 331 -851 331 -851 0 net=2417
rlabel metal2 2 -853 2 -853 0 net=2725
rlabel metal2 205 -853 205 -853 0 net=1005
rlabel metal2 261 -853 261 -853 0 net=1417
rlabel metal2 345 -853 345 -853 0 net=1665
rlabel metal2 128 -855 128 -855 0 net=2265
rlabel metal2 296 -855 296 -855 0 net=2033
rlabel metal2 355 -855 355 -855 0 net=2452
rlabel metal2 156 -857 156 -857 0 net=877
rlabel metal2 226 -857 226 -857 0 net=2495
rlabel metal2 520 -857 520 -857 0 net=2785
rlabel metal2 233 -859 233 -859 0 net=867
rlabel metal2 296 -859 296 -859 0 net=1231
rlabel metal2 2 -870 2 -870 0 net=2726
rlabel metal2 152 -870 152 -870 0 net=2246
rlabel metal2 425 -870 425 -870 0 net=2980
rlabel metal2 516 -870 516 -870 0 net=182
rlabel metal2 2 -872 2 -872 0 net=1395
rlabel metal2 121 -872 121 -872 0 net=856
rlabel metal2 205 -872 205 -872 0 net=868
rlabel metal2 247 -872 247 -872 0 net=890
rlabel metal2 345 -872 345 -872 0 net=2269
rlabel metal2 443 -872 443 -872 0 net=2418
rlabel metal2 9 -874 9 -874 0 net=2582
rlabel metal2 47 -874 47 -874 0 net=98
rlabel metal2 135 -874 135 -874 0 net=1083
rlabel metal2 156 -874 156 -874 0 net=879
rlabel metal2 240 -874 240 -874 0 net=997
rlabel metal2 261 -874 261 -874 0 net=1233
rlabel metal2 299 -874 299 -874 0 net=1859
rlabel metal2 401 -874 401 -874 0 net=2289
rlabel metal2 453 -874 453 -874 0 net=2854
rlabel metal2 492 -874 492 -874 0 net=2587
rlabel metal2 492 -874 492 -874 0 net=2587
rlabel metal2 520 -874 520 -874 0 net=2787
rlabel metal2 537 -874 537 -874 0 net=797
rlabel metal2 548 -874 548 -874 0 net=1557
rlabel metal2 16 -876 16 -876 0 net=2322
rlabel metal2 44 -876 44 -876 0 net=792
rlabel metal2 54 -876 54 -876 0 net=162
rlabel metal2 142 -876 142 -876 0 net=1041
rlabel metal2 268 -876 268 -876 0 net=2905
rlabel metal2 520 -876 520 -876 0 net=2703
rlabel metal2 16 -878 16 -878 0 net=1207
rlabel metal2 61 -878 61 -878 0 net=1670
rlabel metal2 79 -878 79 -878 0 net=2266
rlabel metal2 173 -878 173 -878 0 net=416
rlabel metal2 376 -878 376 -878 0 net=2430
rlabel metal2 485 -878 485 -878 0 net=2619
rlabel metal2 527 -878 527 -878 0 net=1528
rlabel metal2 23 -880 23 -880 0 net=2212
rlabel metal2 65 -880 65 -880 0 net=756
rlabel metal2 191 -880 191 -880 0 net=2195
rlabel metal2 478 -880 478 -880 0 net=2775
rlabel metal2 23 -882 23 -882 0 net=1199
rlabel metal2 163 -882 163 -882 0 net=1365
rlabel metal2 208 -882 208 -882 0 net=2144
rlabel metal2 348 -882 348 -882 0 net=1424
rlabel metal2 380 -882 380 -882 0 net=2320
rlabel metal2 457 -882 457 -882 0 net=2497
rlabel metal2 457 -882 457 -882 0 net=2497
rlabel metal2 68 -884 68 -884 0 net=1430
rlabel metal2 93 -884 93 -884 0 net=1314
rlabel metal2 212 -884 212 -884 0 net=1253
rlabel metal2 282 -884 282 -884 0 net=1309
rlabel metal2 422 -884 422 -884 0 net=1959
rlabel metal2 79 -886 79 -886 0 net=1863
rlabel metal2 194 -886 194 -886 0 net=1517
rlabel metal2 352 -886 352 -886 0 net=1751
rlabel metal2 86 -888 86 -888 0 net=989
rlabel metal2 121 -888 121 -888 0 net=213
rlabel metal2 198 -888 198 -888 0 net=2093
rlabel metal2 96 -890 96 -890 0 net=222
rlabel metal2 219 -890 219 -890 0 net=1045
rlabel metal2 275 -890 275 -890 0 net=1347
rlabel metal2 292 -890 292 -890 0 net=2252
rlabel metal2 100 -892 100 -892 0 net=1405
rlabel metal2 191 -892 191 -892 0 net=829
rlabel metal2 222 -892 222 -892 0 net=1583
rlabel metal2 415 -892 415 -892 0 net=2073
rlabel metal2 100 -894 100 -894 0 net=921
rlabel metal2 226 -894 226 -894 0 net=1924
rlabel metal2 331 -894 331 -894 0 net=2035
rlabel metal2 37 -896 37 -896 0 net=1411
rlabel metal2 408 -896 408 -896 0 net=2485
rlabel metal2 229 -898 229 -898 0 net=1006
rlabel metal2 282 -898 282 -898 0 net=1167
rlabel metal2 208 -900 208 -900 0 net=3007
rlabel metal2 243 -902 243 -902 0 net=2659
rlabel metal2 254 -904 254 -904 0 net=967
rlabel metal2 292 -904 292 -904 0 net=2494
rlabel metal2 303 -906 303 -906 0 net=1418
rlabel metal2 317 -906 317 -906 0 net=1667
rlabel metal2 394 -906 394 -906 0 net=1885
rlabel metal2 65 -908 65 -908 0 net=1861
rlabel metal2 306 -910 306 -910 0 net=490
rlabel metal2 310 -912 310 -912 0 net=2153
rlabel metal2 324 -914 324 -914 0 net=1459
rlabel metal2 9 -925 9 -925 0 net=1862
rlabel metal2 429 -925 429 -925 0 net=2487
rlabel metal2 450 -925 450 -925 0 net=2155
rlabel metal2 474 -925 474 -925 0 net=2620
rlabel metal2 506 -925 506 -925 0 net=2776
rlabel metal2 530 -925 530 -925 0 net=1558
rlabel metal2 16 -927 16 -927 0 net=1208
rlabel metal2 37 -927 37 -927 0 net=362
rlabel metal2 173 -927 173 -927 0 net=713
rlabel metal2 485 -927 485 -927 0 net=2704
rlabel metal2 23 -929 23 -929 0 net=1200
rlabel metal2 79 -929 79 -929 0 net=1864
rlabel metal2 149 -929 149 -929 0 net=1412
rlabel metal2 359 -929 359 -929 0 net=2660
rlabel metal2 506 -929 506 -929 0 net=2953
rlabel metal2 23 -931 23 -931 0 net=2239
rlabel metal2 163 -931 163 -931 0 net=1366
rlabel metal2 201 -931 201 -931 0 net=1860
rlabel metal2 415 -931 415 -931 0 net=2075
rlabel metal2 450 -931 450 -931 0 net=2589
rlabel metal2 44 -933 44 -933 0 net=227
rlabel metal2 184 -933 184 -933 0 net=998
rlabel metal2 264 -933 264 -933 0 net=2036
rlabel metal2 457 -933 457 -933 0 net=2499
rlabel metal2 457 -933 457 -933 0 net=2499
rlabel metal2 478 -933 478 -933 0 net=798
rlabel metal2 54 -935 54 -935 0 net=366
rlabel metal2 208 -935 208 -935 0 net=1254
rlabel metal2 226 -935 226 -935 0 net=1960
rlabel metal2 436 -935 436 -935 0 net=2907
rlabel metal2 58 -937 58 -937 0 net=990
rlabel metal2 93 -937 93 -937 0 net=447
rlabel metal2 268 -937 268 -937 0 net=1047
rlabel metal2 285 -937 285 -937 0 net=641
rlabel metal2 387 -937 387 -937 0 net=2291
rlabel metal2 499 -937 499 -937 0 net=2789
rlabel metal2 58 -939 58 -939 0 net=1043
rlabel metal2 177 -939 177 -939 0 net=1907
rlabel metal2 268 -939 268 -939 0 net=1461
rlabel metal2 345 -939 345 -939 0 net=2271
rlabel metal2 2 -941 2 -941 0 net=1396
rlabel metal2 152 -941 152 -941 0 net=943
rlabel metal2 187 -941 187 -941 0 net=1531
rlabel metal2 233 -941 233 -941 0 net=881
rlabel metal2 338 -941 338 -941 0 net=1519
rlabel metal2 359 -941 359 -941 0 net=1585
rlabel metal2 373 -941 373 -941 0 net=1311
rlabel metal2 30 -943 30 -943 0 net=1107
rlabel metal2 243 -943 243 -943 0 net=1925
rlabel metal2 373 -943 373 -943 0 net=1801
rlabel metal2 72 -945 72 -945 0 net=969
rlabel metal2 299 -945 299 -945 0 net=1668
rlabel metal2 320 -945 320 -945 0 net=3013
rlabel metal2 79 -947 79 -947 0 net=2181
rlabel metal2 114 -947 114 -947 0 net=923
rlabel metal2 187 -947 187 -947 0 net=2196
rlabel metal2 68 -949 68 -949 0 net=439
rlabel metal2 86 -951 86 -951 0 net=1159
rlabel metal2 338 -951 338 -951 0 net=1817
rlabel metal2 93 -953 93 -953 0 net=1039
rlabel metal2 191 -953 191 -953 0 net=729
rlabel metal2 208 -953 208 -953 0 net=3008
rlabel metal2 96 -955 96 -955 0 net=267
rlabel metal2 303 -955 303 -955 0 net=1437
rlabel metal2 362 -955 362 -955 0 net=1886
rlabel metal2 100 -957 100 -957 0 net=1406
rlabel metal2 194 -957 194 -957 0 net=830
rlabel metal2 254 -957 254 -957 0 net=1235
rlabel metal2 282 -957 282 -957 0 net=1169
rlabel metal2 306 -957 306 -957 0 net=1752
rlabel metal2 100 -959 100 -959 0 net=991
rlabel metal2 170 -959 170 -959 0 net=819
rlabel metal2 289 -959 289 -959 0 net=1997
rlabel metal2 310 -959 310 -959 0 net=2095
rlabel metal2 110 -961 110 -961 0 net=660
rlabel metal2 128 -961 128 -961 0 net=339
rlabel metal2 352 -961 352 -961 0 net=2731
rlabel metal2 135 -963 135 -963 0 net=1085
rlabel metal2 219 -963 219 -963 0 net=1349
rlabel metal2 65 -965 65 -965 0 net=231
rlabel metal2 135 -967 135 -967 0 net=2177
rlabel metal2 16 -978 16 -978 0 net=2183
rlabel metal2 107 -978 107 -978 0 net=130
rlabel metal2 219 -978 219 -978 0 net=1350
rlabel metal2 292 -978 292 -978 0 net=1048
rlabel metal2 331 -978 331 -978 0 net=1438
rlabel metal2 520 -978 520 -978 0 net=2955
rlabel metal2 23 -980 23 -980 0 net=2240
rlabel metal2 320 -980 320 -980 0 net=1312
rlabel metal2 408 -980 408 -980 0 net=2807
rlabel metal2 464 -980 464 -980 0 net=2790
rlabel metal2 26 -982 26 -982 0 net=54
rlabel metal2 51 -982 51 -982 0 net=2179
rlabel metal2 142 -982 142 -982 0 net=765
rlabel metal2 142 -982 142 -982 0 net=765
rlabel metal2 156 -982 156 -982 0 net=1086
rlabel metal2 247 -982 247 -982 0 net=883
rlabel metal2 247 -982 247 -982 0 net=883
rlabel metal2 261 -982 261 -982 0 net=1520
rlabel metal2 352 -982 352 -982 0 net=2156
rlabel metal2 478 -982 478 -982 0 net=2339
rlabel metal2 478 -982 478 -982 0 net=2339
rlabel metal2 30 -984 30 -984 0 net=1108
rlabel metal2 271 -984 271 -984 0 net=2455
rlabel metal2 380 -984 380 -984 0 net=2488
rlabel metal2 446 -984 446 -984 0 net=2501
rlabel metal2 471 -984 471 -984 0 net=2733
rlabel metal2 37 -986 37 -986 0 net=2407
rlabel metal2 135 -986 135 -986 0 net=731
rlabel metal2 208 -986 208 -986 0 net=367
rlabel metal2 303 -986 303 -986 0 net=1171
rlabel metal2 411 -986 411 -986 0 net=2076
rlabel metal2 58 -988 58 -988 0 net=1044
rlabel metal2 131 -988 131 -988 0 net=1532
rlabel metal2 229 -988 229 -988 0 net=1236
rlabel metal2 278 -988 278 -988 0 net=2969
rlabel metal2 422 -988 422 -988 0 net=2500
rlabel metal2 58 -990 58 -990 0 net=993
rlabel metal2 107 -990 107 -990 0 net=925
rlabel metal2 128 -990 128 -990 0 net=452
rlabel metal2 212 -990 212 -990 0 net=1999
rlabel metal2 296 -990 296 -990 0 net=2215
rlabel metal2 390 -990 390 -990 0 net=793
rlabel metal2 429 -990 429 -990 0 net=551
rlabel metal2 65 -992 65 -992 0 net=209
rlabel metal2 121 -992 121 -992 0 net=1793
rlabel metal2 191 -992 191 -992 0 net=1961
rlabel metal2 299 -992 299 -992 0 net=2096
rlabel metal2 324 -992 324 -992 0 net=2272
rlabel metal2 443 -992 443 -992 0 net=2843
rlabel metal2 65 -994 65 -994 0 net=602
rlabel metal2 156 -994 156 -994 0 net=821
rlabel metal2 173 -994 173 -994 0 net=4
rlabel metal2 233 -994 233 -994 0 net=115
rlabel metal2 303 -994 303 -994 0 net=1819
rlabel metal2 394 -994 394 -994 0 net=3015
rlabel metal2 68 -996 68 -996 0 net=1040
rlabel metal2 100 -996 100 -996 0 net=1903
rlabel metal2 149 -996 149 -996 0 net=1479
rlabel metal2 177 -996 177 -996 0 net=944
rlabel metal2 240 -996 240 -996 0 net=1909
rlabel metal2 338 -996 338 -996 0 net=1803
rlabel metal2 394 -996 394 -996 0 net=2909
rlabel metal2 30 -998 30 -998 0 net=1117
rlabel metal2 72 -998 72 -998 0 net=971
rlabel metal2 236 -998 236 -998 0 net=1225
rlabel metal2 366 -998 366 -998 0 net=1927
rlabel metal2 436 -998 436 -998 0 net=2591
rlabel metal2 72 -1000 72 -1000 0 net=1161
rlabel metal2 110 -1000 110 -1000 0 net=1586
rlabel metal2 79 -1002 79 -1002 0 net=841
rlabel metal2 163 -1002 163 -1002 0 net=1087
rlabel metal2 317 -1002 317 -1002 0 net=1241
rlabel metal2 177 -1004 177 -1004 0 net=1049
rlabel metal2 359 -1004 359 -1004 0 net=2293
rlabel metal2 198 -1006 198 -1006 0 net=2401
rlabel metal2 201 -1008 201 -1008 0 net=2405
rlabel metal2 268 -1008 268 -1008 0 net=1462
rlabel metal2 30 -1019 30 -1019 0 net=1118
rlabel metal2 51 -1019 51 -1019 0 net=2180
rlabel metal2 208 -1019 208 -1019 0 net=972
rlabel metal2 247 -1019 247 -1019 0 net=884
rlabel metal2 278 -1019 278 -1019 0 net=1804
rlabel metal2 355 -1019 355 -1019 0 net=2216
rlabel metal2 415 -1019 415 -1019 0 net=3017
rlabel metal2 415 -1019 415 -1019 0 net=3017
rlabel metal2 422 -1019 422 -1019 0 net=794
rlabel metal2 422 -1019 422 -1019 0 net=794
rlabel metal2 436 -1019 436 -1019 0 net=2592
rlabel metal2 453 -1019 453 -1019 0 net=2734
rlabel metal2 478 -1019 478 -1019 0 net=2341
rlabel metal2 478 -1019 478 -1019 0 net=2341
rlabel metal2 523 -1019 523 -1019 0 net=2956
rlabel metal2 58 -1021 58 -1021 0 net=994
rlabel metal2 114 -1021 114 -1021 0 net=665
rlabel metal2 240 -1021 240 -1021 0 net=1227
rlabel metal2 289 -1021 289 -1021 0 net=2910
rlabel metal2 443 -1021 443 -1021 0 net=401
rlabel metal2 453 -1021 453 -1021 0 net=2502
rlabel metal2 516 -1021 516 -1021 0 net=692
rlabel metal2 16 -1023 16 -1023 0 net=2184
rlabel metal2 121 -1023 121 -1023 0 net=1794
rlabel metal2 205 -1023 205 -1023 0 net=1893
rlabel metal2 247 -1023 247 -1023 0 net=1681
rlabel metal2 296 -1023 296 -1023 0 net=1821
rlabel metal2 310 -1023 310 -1023 0 net=1911
rlabel metal2 310 -1023 310 -1023 0 net=1911
rlabel metal2 324 -1023 324 -1023 0 net=184
rlabel metal2 359 -1023 359 -1023 0 net=2295
rlabel metal2 369 -1023 369 -1023 0 net=2970
rlabel metal2 457 -1023 457 -1023 0 net=2845
rlabel metal2 457 -1023 457 -1023 0 net=2845
rlabel metal2 520 -1023 520 -1023 0 net=3023
rlabel metal2 65 -1025 65 -1025 0 net=843
rlabel metal2 86 -1025 86 -1025 0 net=408
rlabel metal2 107 -1025 107 -1025 0 net=927
rlabel metal2 142 -1025 142 -1025 0 net=766
rlabel metal2 177 -1025 177 -1025 0 net=1051
rlabel metal2 229 -1025 229 -1025 0 net=2915
rlabel metal2 72 -1027 72 -1027 0 net=1163
rlabel metal2 135 -1027 135 -1027 0 net=733
rlabel metal2 184 -1027 184 -1027 0 net=387
rlabel metal2 208 -1027 208 -1027 0 net=2000
rlabel metal2 215 -1027 215 -1027 0 net=1791
rlabel metal2 324 -1027 324 -1027 0 net=2185
rlabel metal2 380 -1027 380 -1027 0 net=2809
rlabel metal2 72 -1029 72 -1029 0 net=2705
rlabel metal2 93 -1029 93 -1029 0 net=1905
rlabel metal2 107 -1029 107 -1029 0 net=2157
rlabel metal2 387 -1029 387 -1029 0 net=2675
rlabel metal2 86 -1031 86 -1031 0 net=330
rlabel metal2 135 -1031 135 -1031 0 net=1481
rlabel metal2 156 -1031 156 -1031 0 net=823
rlabel metal2 212 -1031 212 -1031 0 net=2831
rlabel metal2 37 -1033 37 -1033 0 net=2408
rlabel metal2 163 -1033 163 -1033 0 net=1089
rlabel metal2 187 -1033 187 -1033 0 net=2406
rlabel metal2 261 -1033 261 -1033 0 net=1963
rlabel metal2 117 -1035 117 -1035 0 net=462
rlabel metal2 233 -1035 233 -1035 0 net=550
rlabel metal2 331 -1035 331 -1035 0 net=2403
rlabel metal2 170 -1037 170 -1037 0 net=1221
rlabel metal2 250 -1037 250 -1037 0 net=1172
rlabel metal2 226 -1039 226 -1039 0 net=1928
rlabel metal2 261 -1041 261 -1041 0 net=1537
rlabel metal2 285 -1041 285 -1041 0 net=3009
rlabel metal2 275 -1043 275 -1043 0 net=1243
rlabel metal2 345 -1043 345 -1043 0 net=2457
rlabel metal2 373 -1043 373 -1043 0 net=2307
rlabel metal2 254 -1045 254 -1045 0 net=2147
rlabel metal2 51 -1056 51 -1056 0 net=2421
rlabel metal2 121 -1056 121 -1056 0 net=929
rlabel metal2 121 -1056 121 -1056 0 net=929
rlabel metal2 128 -1056 128 -1056 0 net=1164
rlabel metal2 201 -1056 201 -1056 0 net=1792
rlabel metal2 320 -1056 320 -1056 0 net=2810
rlabel metal2 429 -1056 429 -1056 0 net=661
rlabel metal2 457 -1056 457 -1056 0 net=2847
rlabel metal2 478 -1056 478 -1056 0 net=2343
rlabel metal2 478 -1056 478 -1056 0 net=2343
rlabel metal2 520 -1056 520 -1056 0 net=3024
rlabel metal2 61 -1058 61 -1058 0 net=390
rlabel metal2 93 -1058 93 -1058 0 net=1906
rlabel metal2 107 -1058 107 -1058 0 net=2158
rlabel metal2 334 -1058 334 -1058 0 net=2308
rlabel metal2 408 -1058 408 -1058 0 net=2677
rlabel metal2 65 -1060 65 -1060 0 net=844
rlabel metal2 93 -1060 93 -1060 0 net=857
rlabel metal2 152 -1060 152 -1060 0 net=1538
rlabel metal2 345 -1060 345 -1060 0 net=2459
rlabel metal2 345 -1060 345 -1060 0 net=2459
rlabel metal2 359 -1060 359 -1060 0 net=2833
rlabel metal2 373 -1060 373 -1060 0 net=2911
rlabel metal2 408 -1060 408 -1060 0 net=3019
rlabel metal2 65 -1062 65 -1062 0 net=2037
rlabel metal2 135 -1062 135 -1062 0 net=1482
rlabel metal2 163 -1062 163 -1062 0 net=1147
rlabel metal2 177 -1062 177 -1062 0 net=734
rlabel metal2 212 -1062 212 -1062 0 net=1244
rlabel metal2 359 -1062 359 -1062 0 net=2297
rlabel metal2 72 -1064 72 -1064 0 net=2706
rlabel metal2 114 -1064 114 -1064 0 net=2597
rlabel metal2 114 -1064 114 -1064 0 net=2597
rlabel metal2 135 -1064 135 -1064 0 net=275
rlabel metal2 366 -1064 366 -1064 0 net=3011
rlabel metal2 75 -1066 75 -1066 0 net=686
rlabel metal2 145 -1066 145 -1066 0 net=559
rlabel metal2 219 -1066 219 -1066 0 net=1052
rlabel metal2 226 -1066 226 -1066 0 net=1759
rlabel metal2 250 -1066 250 -1066 0 net=2404
rlabel metal2 394 -1066 394 -1066 0 net=2917
rlabel metal2 100 -1068 100 -1068 0 net=2359
rlabel metal2 149 -1068 149 -1068 0 net=945
rlabel metal2 236 -1068 236 -1068 0 net=2971
rlabel metal2 156 -1070 156 -1070 0 net=1217
rlabel metal2 219 -1070 219 -1070 0 net=2803
rlabel metal2 163 -1072 163 -1072 0 net=1223
rlabel metal2 177 -1072 177 -1072 0 net=1269
rlabel metal2 236 -1072 236 -1072 0 net=2529
rlabel metal2 184 -1074 184 -1074 0 net=1091
rlabel metal2 240 -1074 240 -1074 0 net=1895
rlabel metal2 240 -1074 240 -1074 0 net=1895
rlabel metal2 247 -1074 247 -1074 0 net=1889
rlabel metal2 306 -1074 306 -1074 0 net=157
rlabel metal2 191 -1076 191 -1076 0 net=825
rlabel metal2 254 -1076 254 -1076 0 net=1229
rlabel metal2 275 -1076 275 -1076 0 net=2149
rlabel metal2 362 -1076 362 -1076 0 net=1
rlabel metal2 142 -1078 142 -1078 0 net=835
rlabel metal2 261 -1080 261 -1080 0 net=1737
rlabel metal2 268 -1082 268 -1082 0 net=1683
rlabel metal2 289 -1082 289 -1082 0 net=1964
rlabel metal2 282 -1084 282 -1084 0 net=999
rlabel metal2 324 -1086 324 -1086 0 net=2187
rlabel metal2 310 -1088 310 -1088 0 net=1913
rlabel metal2 296 -1090 296 -1090 0 net=1823
rlabel metal2 30 -1101 30 -1101 0 net=859
rlabel metal2 100 -1101 100 -1101 0 net=2360
rlabel metal2 114 -1101 114 -1101 0 net=2598
rlabel metal2 226 -1101 226 -1101 0 net=1761
rlabel metal2 460 -1101 460 -1101 0 net=2848
rlabel metal2 478 -1101 478 -1101 0 net=2345
rlabel metal2 478 -1101 478 -1101 0 net=2345
rlabel metal2 37 -1103 37 -1103 0 net=2223
rlabel metal2 254 -1103 254 -1103 0 net=1230
rlabel metal2 306 -1103 306 -1103 0 net=2460
rlabel metal2 352 -1103 352 -1103 0 net=2530
rlabel metal2 422 -1103 422 -1103 0 net=2973
rlabel metal2 51 -1105 51 -1105 0 net=2422
rlabel metal2 100 -1105 100 -1105 0 net=777
rlabel metal2 121 -1105 121 -1105 0 net=930
rlabel metal2 142 -1105 142 -1105 0 net=837
rlabel metal2 184 -1105 184 -1105 0 net=1890
rlabel metal2 254 -1105 254 -1105 0 net=2937
rlabel metal2 359 -1105 359 -1105 0 net=2298
rlabel metal2 387 -1105 387 -1105 0 net=3020
rlabel metal2 415 -1105 415 -1105 0 net=2678
rlabel metal2 54 -1107 54 -1107 0 net=747
rlabel metal2 65 -1107 65 -1107 0 net=2038
rlabel metal2 219 -1107 219 -1107 0 net=1183
rlabel metal2 317 -1107 317 -1107 0 net=2188
rlabel metal2 345 -1107 345 -1107 0 net=2867
rlabel metal2 362 -1107 362 -1107 0 net=3012
rlabel metal2 380 -1107 380 -1107 0 net=2913
rlabel metal2 65 -1109 65 -1109 0 net=1219
rlabel metal2 163 -1109 163 -1109 0 net=1224
rlabel metal2 226 -1109 226 -1109 0 net=1896
rlabel metal2 247 -1109 247 -1109 0 net=1685
rlabel metal2 275 -1109 275 -1109 0 net=2150
rlabel metal2 275 -1109 275 -1109 0 net=2150
rlabel metal2 320 -1109 320 -1109 0 net=1901
rlabel metal2 394 -1109 394 -1109 0 net=2835
rlabel metal2 72 -1111 72 -1111 0 net=80
rlabel metal2 82 -1111 82 -1111 0 net=459
rlabel metal2 121 -1111 121 -1111 0 net=1701
rlabel metal2 142 -1111 142 -1111 0 net=947
rlabel metal2 159 -1111 159 -1111 0 net=895
rlabel metal2 170 -1111 170 -1111 0 net=1149
rlabel metal2 191 -1111 191 -1111 0 net=144
rlabel metal2 233 -1111 233 -1111 0 net=807
rlabel metal2 401 -1111 401 -1111 0 net=2919
rlabel metal2 44 -1113 44 -1113 0 net=1745
rlabel metal2 107 -1113 107 -1113 0 net=1561
rlabel metal2 170 -1113 170 -1113 0 net=1092
rlabel metal2 268 -1113 268 -1113 0 net=1001
rlabel metal2 289 -1113 289 -1113 0 net=1101
rlabel metal2 324 -1113 324 -1113 0 net=1915
rlabel metal2 75 -1115 75 -1115 0 net=875
rlabel metal2 131 -1115 131 -1115 0 net=795
rlabel metal2 198 -1115 198 -1115 0 net=1271
rlabel metal2 278 -1115 278 -1115 0 net=2235
rlabel metal2 205 -1117 205 -1117 0 net=827
rlabel metal2 282 -1117 282 -1117 0 net=1825
rlabel metal2 331 -1117 331 -1117 0 net=2805
rlabel metal2 194 -1119 194 -1119 0 net=2253
rlabel metal2 338 -1119 338 -1119 0 net=2225
rlabel metal2 205 -1121 205 -1121 0 net=2167
rlabel metal2 261 -1123 261 -1123 0 net=1739
rlabel metal2 180 -1125 180 -1125 0 net=25
rlabel metal2 296 -1125 296 -1125 0 net=2643
rlabel metal2 264 -1127 264 -1127 0 net=2049
rlabel metal2 30 -1138 30 -1138 0 net=860
rlabel metal2 107 -1138 107 -1138 0 net=876
rlabel metal2 149 -1138 149 -1138 0 net=796
rlabel metal2 205 -1138 205 -1138 0 net=828
rlabel metal2 250 -1138 250 -1138 0 net=1002
rlabel metal2 275 -1138 275 -1138 0 net=1916
rlabel metal2 397 -1138 397 -1138 0 net=2974
rlabel metal2 478 -1138 478 -1138 0 net=2346
rlabel metal2 37 -1140 37 -1140 0 net=2224
rlabel metal2 177 -1140 177 -1140 0 net=839
rlabel metal2 177 -1140 177 -1140 0 net=839
rlabel metal2 184 -1140 184 -1140 0 net=1150
rlabel metal2 229 -1140 229 -1140 0 net=1565
rlabel metal2 296 -1140 296 -1140 0 net=2051
rlabel metal2 327 -1140 327 -1140 0 net=2644
rlabel metal2 44 -1142 44 -1142 0 net=1746
rlabel metal2 58 -1142 58 -1142 0 net=749
rlabel metal2 75 -1142 75 -1142 0 net=315
rlabel metal2 86 -1142 86 -1142 0 net=3021
rlabel metal2 254 -1142 254 -1142 0 net=1762
rlabel metal2 65 -1144 65 -1144 0 net=1220
rlabel metal2 163 -1144 163 -1144 0 net=896
rlabel metal2 184 -1144 184 -1144 0 net=931
rlabel metal2 261 -1144 261 -1144 0 net=1826
rlabel metal2 299 -1144 299 -1144 0 net=2806
rlabel metal2 79 -1146 79 -1146 0 net=778
rlabel metal2 107 -1146 107 -1146 0 net=1703
rlabel metal2 128 -1146 128 -1146 0 net=845
rlabel metal2 306 -1146 306 -1146 0 net=2920
rlabel metal2 89 -1148 89 -1148 0 net=359
rlabel metal2 117 -1148 117 -1148 0 net=670
rlabel metal2 201 -1148 201 -1148 0 net=2995
rlabel metal2 306 -1148 306 -1148 0 net=3033
rlabel metal2 369 -1148 369 -1148 0 net=2914
rlabel metal2 93 -1150 93 -1150 0 net=293
rlabel metal2 261 -1150 261 -1150 0 net=1902
rlabel metal2 376 -1150 376 -1150 0 net=2836
rlabel metal2 100 -1152 100 -1152 0 net=1979
rlabel metal2 149 -1152 149 -1152 0 net=1195
rlabel metal2 208 -1152 208 -1152 0 net=2236
rlabel metal2 401 -1152 401 -1152 0 net=1629
rlabel metal2 117 -1154 117 -1154 0 net=7
rlabel metal2 268 -1154 268 -1154 0 net=1103
rlabel metal2 310 -1154 310 -1154 0 net=2255
rlabel metal2 121 -1156 121 -1156 0 net=1562
rlabel metal2 156 -1156 156 -1156 0 net=1691
rlabel metal2 191 -1156 191 -1156 0 net=1185
rlabel metal2 278 -1156 278 -1156 0 net=1943
rlabel metal2 317 -1156 317 -1156 0 net=1741
rlabel metal2 338 -1156 338 -1156 0 net=2227
rlabel metal2 135 -1158 135 -1158 0 net=1643
rlabel metal2 163 -1158 163 -1158 0 net=2975
rlabel metal2 212 -1160 212 -1160 0 net=1273
rlabel metal2 240 -1160 240 -1160 0 net=2997
rlabel metal2 142 -1162 142 -1162 0 net=949
rlabel metal2 219 -1162 219 -1162 0 net=809
rlabel metal2 264 -1162 264 -1162 0 net=2855
rlabel metal2 233 -1164 233 -1164 0 net=1687
rlabel metal2 264 -1164 264 -1164 0 net=2168
rlabel metal2 352 -1166 352 -1166 0 net=2939
rlabel metal2 345 -1168 345 -1168 0 net=2869
rlabel metal2 254 -1170 254 -1170 0 net=2861
rlabel metal2 61 -1181 61 -1181 0 net=750
rlabel metal2 79 -1181 79 -1181 0 net=1645
rlabel metal2 163 -1181 163 -1181 0 net=933
rlabel metal2 198 -1181 198 -1181 0 net=197
rlabel metal2 208 -1181 208 -1181 0 net=950
rlabel metal2 240 -1181 240 -1181 0 net=2996
rlabel metal2 292 -1181 292 -1181 0 net=1630
rlabel metal2 72 -1183 72 -1183 0 net=961
rlabel metal2 121 -1183 121 -1183 0 net=1196
rlabel metal2 177 -1183 177 -1183 0 net=840
rlabel metal2 212 -1183 212 -1183 0 net=799
rlabel metal2 247 -1183 247 -1183 0 net=1104
rlabel metal2 303 -1183 303 -1183 0 net=2256
rlabel metal2 86 -1185 86 -1185 0 net=3022
rlabel metal2 173 -1185 173 -1185 0 net=2795
rlabel metal2 250 -1185 250 -1185 0 net=1917
rlabel metal2 376 -1185 376 -1185 0 net=1127
rlabel metal2 65 -1187 65 -1187 0 net=1015
rlabel metal2 184 -1187 184 -1187 0 net=1274
rlabel metal2 254 -1187 254 -1187 0 net=2863
rlabel metal2 359 -1187 359 -1187 0 net=3035
rlabel metal2 359 -1187 359 -1187 0 net=3035
rlabel metal2 366 -1187 366 -1187 0 net=2228
rlabel metal2 93 -1189 93 -1189 0 net=2821
rlabel metal2 128 -1189 128 -1189 0 net=847
rlabel metal2 201 -1189 201 -1189 0 net=2679
rlabel metal2 324 -1189 324 -1189 0 net=2053
rlabel metal2 331 -1189 331 -1189 0 net=2857
rlabel metal2 331 -1189 331 -1189 0 net=2857
rlabel metal2 366 -1189 366 -1189 0 net=2941
rlabel metal2 107 -1191 107 -1191 0 net=1704
rlabel metal2 194 -1191 194 -1191 0 net=1375
rlabel metal2 324 -1191 324 -1191 0 net=2998
rlabel metal2 383 -1191 383 -1191 0 net=2469
rlabel metal2 100 -1193 100 -1193 0 net=1980
rlabel metal2 114 -1193 114 -1193 0 net=1693
rlabel metal2 233 -1193 233 -1193 0 net=1689
rlabel metal2 100 -1195 100 -1195 0 net=1635
rlabel metal2 338 -1195 338 -1195 0 net=2871
rlabel metal2 121 -1197 121 -1197 0 net=811
rlabel metal2 233 -1197 233 -1197 0 net=891
rlabel metal2 142 -1199 142 -1199 0 net=1305
rlabel metal2 191 -1199 191 -1199 0 net=1187
rlabel metal2 257 -1199 257 -1199 0 net=1566
rlabel metal2 296 -1199 296 -1199 0 net=1945
rlabel metal2 138 -1201 138 -1201 0 net=600
rlabel metal2 275 -1201 275 -1201 0 net=2977
rlabel metal2 310 -1201 310 -1201 0 net=1743
rlabel metal2 65 -1212 65 -1212 0 net=1016
rlabel metal2 194 -1212 194 -1212 0 net=2796
rlabel metal2 261 -1212 261 -1212 0 net=735
rlabel metal2 292 -1212 292 -1212 0 net=2054
rlabel metal2 380 -1212 380 -1212 0 net=2471
rlabel metal2 72 -1214 72 -1214 0 net=962
rlabel metal2 93 -1214 93 -1214 0 net=2823
rlabel metal2 93 -1214 93 -1214 0 net=2823
rlabel metal2 114 -1214 114 -1214 0 net=1695
rlabel metal2 163 -1214 163 -1214 0 net=935
rlabel metal2 163 -1214 163 -1214 0 net=935
rlabel metal2 170 -1214 170 -1214 0 net=2055
rlabel metal2 261 -1214 261 -1214 0 net=1918
rlabel metal2 383 -1214 383 -1214 0 net=1128
rlabel metal2 79 -1216 79 -1216 0 net=1646
rlabel metal2 149 -1216 149 -1216 0 net=1188
rlabel metal2 240 -1216 240 -1216 0 net=3036
rlabel metal2 107 -1218 107 -1218 0 net=2077
rlabel metal2 121 -1218 121 -1218 0 net=812
rlabel metal2 264 -1218 264 -1218 0 net=1690
rlabel metal2 352 -1218 352 -1218 0 net=2943
rlabel metal2 121 -1220 121 -1220 0 net=210
rlabel metal2 184 -1220 184 -1220 0 net=2633
rlabel metal2 275 -1220 275 -1220 0 net=2978
rlabel metal2 324 -1220 324 -1220 0 net=2859
rlabel metal2 128 -1222 128 -1222 0 net=254
rlabel metal2 177 -1222 177 -1222 0 net=2864
rlabel metal2 268 -1222 268 -1222 0 net=2681
rlabel metal2 331 -1222 331 -1222 0 net=2873
rlabel metal2 100 -1224 100 -1224 0 net=1637
rlabel metal2 135 -1224 135 -1224 0 net=1659
rlabel metal2 205 -1224 205 -1224 0 net=801
rlabel metal2 233 -1224 233 -1224 0 net=892
rlabel metal2 303 -1224 303 -1224 0 net=1744
rlabel metal2 142 -1226 142 -1226 0 net=1306
rlabel metal2 198 -1226 198 -1226 0 net=849
rlabel metal2 240 -1226 240 -1226 0 net=1975
rlabel metal2 282 -1226 282 -1226 0 net=1377
rlabel metal2 142 -1228 142 -1228 0 net=2281
rlabel metal2 212 -1228 212 -1228 0 net=1367
rlabel metal2 282 -1228 282 -1228 0 net=1947
rlabel metal2 275 -1230 275 -1230 0 net=1837
rlabel metal2 82 -1241 82 -1241 0 net=1545
rlabel metal2 93 -1241 93 -1241 0 net=2824
rlabel metal2 107 -1241 107 -1241 0 net=2433
rlabel metal2 128 -1241 128 -1241 0 net=1638
rlabel metal2 156 -1241 156 -1241 0 net=1696
rlabel metal2 212 -1241 212 -1241 0 net=1368
rlabel metal2 233 -1241 233 -1241 0 net=850
rlabel metal2 275 -1241 275 -1241 0 net=1839
rlabel metal2 299 -1241 299 -1241 0 net=1378
rlabel metal2 317 -1241 317 -1241 0 net=2682
rlabel metal2 348 -1241 348 -1241 0 net=2944
rlabel metal2 380 -1241 380 -1241 0 net=2473
rlabel metal2 380 -1241 380 -1241 0 net=2473
rlabel metal2 100 -1243 100 -1243 0 net=3005
rlabel metal2 128 -1243 128 -1243 0 net=2282
rlabel metal2 156 -1243 156 -1243 0 net=2634
rlabel metal2 240 -1243 240 -1243 0 net=1977
rlabel metal2 282 -1243 282 -1243 0 net=1949
rlabel metal2 306 -1243 306 -1243 0 net=2860
rlabel metal2 110 -1245 110 -1245 0 net=2078
rlabel metal2 135 -1245 135 -1245 0 net=1660
rlabel metal2 177 -1245 177 -1245 0 net=1457
rlabel metal2 198 -1245 198 -1245 0 net=1125
rlabel metal2 226 -1245 226 -1245 0 net=2001
rlabel metal2 254 -1245 254 -1245 0 net=2553
rlabel metal2 285 -1245 285 -1245 0 net=736
rlabel metal2 324 -1245 324 -1245 0 net=2875
rlabel metal2 135 -1247 135 -1247 0 net=1017
rlabel metal2 163 -1247 163 -1247 0 net=936
rlabel metal2 191 -1247 191 -1247 0 net=803
rlabel metal2 268 -1247 268 -1247 0 net=2555
rlabel metal2 180 -1249 180 -1249 0 net=2056
rlabel metal2 205 -1251 205 -1251 0 net=1023
rlabel metal2 240 -1251 240 -1251 0 net=1941
rlabel metal2 5 -1262 5 -1262 0 net=718
rlabel metal2 5 -1262 5 -1262 0 net=718
rlabel metal2 75 -1262 75 -1262 0 net=438
rlabel metal2 86 -1262 86 -1262 0 net=1546
rlabel metal2 86 -1262 86 -1262 0 net=1546
rlabel metal2 100 -1262 100 -1262 0 net=3006
rlabel metal2 135 -1262 135 -1262 0 net=1018
rlabel metal2 170 -1262 170 -1262 0 net=11
rlabel metal2 184 -1262 184 -1262 0 net=342
rlabel metal2 184 -1262 184 -1262 0 net=342
rlabel metal2 205 -1262 205 -1262 0 net=1025
rlabel metal2 233 -1262 233 -1262 0 net=2002
rlabel metal2 233 -1262 233 -1262 0 net=2002
rlabel metal2 240 -1262 240 -1262 0 net=1942
rlabel metal2 240 -1262 240 -1262 0 net=1942
rlabel metal2 254 -1262 254 -1262 0 net=2554
rlabel metal2 275 -1262 275 -1262 0 net=1840
rlabel metal2 303 -1262 303 -1262 0 net=1951
rlabel metal2 303 -1262 303 -1262 0 net=1951
rlabel metal2 320 -1262 320 -1262 0 net=2876
rlabel metal2 380 -1262 380 -1262 0 net=2475
rlabel metal2 107 -1264 107 -1264 0 net=2435
rlabel metal2 107 -1264 107 -1264 0 net=2435
rlabel metal2 114 -1264 114 -1264 0 net=288
rlabel metal2 135 -1264 135 -1264 0 net=2489
rlabel metal2 149 -1264 149 -1264 0 net=1469
rlabel metal2 149 -1264 149 -1264 0 net=1469
rlabel metal2 163 -1264 163 -1264 0 net=1458
rlabel metal2 191 -1264 191 -1264 0 net=804
rlabel metal2 215 -1264 215 -1264 0 net=1126
rlabel metal2 261 -1264 261 -1264 0 net=1978
rlabel metal2 117 -1266 117 -1266 0 net=1137
rlabel metal2 268 -1266 268 -1266 0 net=2557
rlabel metal2 86 -1277 86 -1277 0 net=172
rlabel metal2 107 -1277 107 -1277 0 net=2436
rlabel metal2 121 -1277 121 -1277 0 net=1138
rlabel metal2 135 -1277 135 -1277 0 net=2490
rlabel metal2 149 -1277 149 -1277 0 net=1470
rlabel metal2 219 -1277 219 -1277 0 net=1026
rlabel metal2 275 -1277 275 -1277 0 net=2558
rlabel metal2 299 -1277 299 -1277 0 net=1952
rlabel metal2 383 -1277 383 -1277 0 net=2476
rlabel metal2 156 -1279 156 -1279 0 net=127
<< end >>
